magic
tech sky130B
timestamp 1662168084
<< metal1 >>
rect 0 7990 8000 8000
rect 0 7955 75 7990
rect 175 7955 325 7990
rect 425 7955 575 7990
rect 675 7955 825 7990
rect 925 7955 1075 7990
rect 1175 7955 1325 7990
rect 1425 7955 1575 7990
rect 1675 7955 1825 7990
rect 1925 7955 2075 7990
rect 2175 7955 2325 7990
rect 2425 7955 2575 7990
rect 2675 7955 2825 7990
rect 2925 7955 3075 7990
rect 3175 7955 3325 7990
rect 3425 7955 3575 7990
rect 3675 7955 3825 7990
rect 3925 7955 4075 7990
rect 4175 7955 4325 7990
rect 4425 7955 4575 7990
rect 4675 7955 4825 7990
rect 4925 7955 5075 7990
rect 5175 7955 5325 7990
rect 5425 7955 5575 7990
rect 5675 7955 5825 7990
rect 5925 7955 6075 7990
rect 6175 7955 6325 7990
rect 6425 7955 6575 7990
rect 6675 7955 6825 7990
rect 6925 7955 7075 7990
rect 7175 7955 7325 7990
rect 7425 7955 7575 7990
rect 7675 7955 7825 7990
rect 7925 7955 8000 7990
rect 0 7950 8000 7955
rect 0 7940 60 7950
rect 190 7940 310 7950
rect 440 7940 560 7950
rect 690 7940 810 7950
rect 940 7940 1060 7950
rect 1190 7940 1310 7950
rect 1440 7940 1560 7950
rect 1690 7940 1810 7950
rect 1940 7940 2060 7950
rect 2190 7940 2310 7950
rect 2440 7940 2560 7950
rect 2690 7940 2810 7950
rect 2940 7940 3060 7950
rect 3190 7940 3310 7950
rect 3440 7940 3560 7950
rect 3690 7940 3810 7950
rect 3940 7940 4060 7950
rect 4190 7940 4310 7950
rect 4440 7940 4560 7950
rect 4690 7940 4810 7950
rect 4940 7940 5060 7950
rect 5190 7940 5310 7950
rect 5440 7940 5560 7950
rect 5690 7940 5810 7950
rect 5940 7940 6060 7950
rect 6190 7940 6310 7950
rect 6440 7940 6560 7950
rect 6690 7940 6810 7950
rect 6940 7940 7060 7950
rect 7190 7940 7310 7950
rect 7440 7940 7560 7950
rect 7690 7940 7810 7950
rect 7940 7940 8000 7950
rect 0 7925 50 7940
rect 0 7825 10 7925
rect 45 7825 50 7925
rect 0 7810 50 7825
rect 200 7925 300 7940
rect 200 7825 205 7925
rect 240 7825 260 7925
rect 295 7825 300 7925
rect 200 7810 300 7825
rect 450 7925 550 7940
rect 450 7825 455 7925
rect 490 7825 510 7925
rect 545 7825 550 7925
rect 450 7810 550 7825
rect 700 7925 800 7940
rect 700 7825 705 7925
rect 740 7825 760 7925
rect 795 7825 800 7925
rect 700 7810 800 7825
rect 950 7925 1050 7940
rect 950 7825 955 7925
rect 990 7825 1010 7925
rect 1045 7825 1050 7925
rect 950 7810 1050 7825
rect 1200 7925 1300 7940
rect 1200 7825 1205 7925
rect 1240 7825 1260 7925
rect 1295 7825 1300 7925
rect 1200 7810 1300 7825
rect 1450 7925 1550 7940
rect 1450 7825 1455 7925
rect 1490 7825 1510 7925
rect 1545 7825 1550 7925
rect 1450 7810 1550 7825
rect 1700 7925 1800 7940
rect 1700 7825 1705 7925
rect 1740 7825 1760 7925
rect 1795 7825 1800 7925
rect 1700 7810 1800 7825
rect 1950 7925 2050 7940
rect 1950 7825 1955 7925
rect 1990 7825 2010 7925
rect 2045 7825 2050 7925
rect 1950 7810 2050 7825
rect 2200 7925 2300 7940
rect 2200 7825 2205 7925
rect 2240 7825 2260 7925
rect 2295 7825 2300 7925
rect 2200 7810 2300 7825
rect 2450 7925 2550 7940
rect 2450 7825 2455 7925
rect 2490 7825 2510 7925
rect 2545 7825 2550 7925
rect 2450 7810 2550 7825
rect 2700 7925 2800 7940
rect 2700 7825 2705 7925
rect 2740 7825 2760 7925
rect 2795 7825 2800 7925
rect 2700 7810 2800 7825
rect 2950 7925 3050 7940
rect 2950 7825 2955 7925
rect 2990 7825 3010 7925
rect 3045 7825 3050 7925
rect 2950 7810 3050 7825
rect 3200 7925 3300 7940
rect 3200 7825 3205 7925
rect 3240 7825 3260 7925
rect 3295 7825 3300 7925
rect 3200 7810 3300 7825
rect 3450 7925 3550 7940
rect 3450 7825 3455 7925
rect 3490 7825 3510 7925
rect 3545 7825 3550 7925
rect 3450 7810 3550 7825
rect 3700 7925 3800 7940
rect 3700 7825 3705 7925
rect 3740 7825 3760 7925
rect 3795 7825 3800 7925
rect 3700 7810 3800 7825
rect 3950 7925 4050 7940
rect 3950 7825 3955 7925
rect 3990 7825 4010 7925
rect 4045 7825 4050 7925
rect 3950 7810 4050 7825
rect 4200 7925 4300 7940
rect 4200 7825 4205 7925
rect 4240 7825 4260 7925
rect 4295 7825 4300 7925
rect 4200 7810 4300 7825
rect 4450 7925 4550 7940
rect 4450 7825 4455 7925
rect 4490 7825 4510 7925
rect 4545 7825 4550 7925
rect 4450 7810 4550 7825
rect 4700 7925 4800 7940
rect 4700 7825 4705 7925
rect 4740 7825 4760 7925
rect 4795 7825 4800 7925
rect 4700 7810 4800 7825
rect 4950 7925 5050 7940
rect 4950 7825 4955 7925
rect 4990 7825 5010 7925
rect 5045 7825 5050 7925
rect 4950 7810 5050 7825
rect 5200 7925 5300 7940
rect 5200 7825 5205 7925
rect 5240 7825 5260 7925
rect 5295 7825 5300 7925
rect 5200 7810 5300 7825
rect 5450 7925 5550 7940
rect 5450 7825 5455 7925
rect 5490 7825 5510 7925
rect 5545 7825 5550 7925
rect 5450 7810 5550 7825
rect 5700 7925 5800 7940
rect 5700 7825 5705 7925
rect 5740 7825 5760 7925
rect 5795 7825 5800 7925
rect 5700 7810 5800 7825
rect 5950 7925 6050 7940
rect 5950 7825 5955 7925
rect 5990 7825 6010 7925
rect 6045 7825 6050 7925
rect 5950 7810 6050 7825
rect 6200 7925 6300 7940
rect 6200 7825 6205 7925
rect 6240 7825 6260 7925
rect 6295 7825 6300 7925
rect 6200 7810 6300 7825
rect 6450 7925 6550 7940
rect 6450 7825 6455 7925
rect 6490 7825 6510 7925
rect 6545 7825 6550 7925
rect 6450 7810 6550 7825
rect 6700 7925 6800 7940
rect 6700 7825 6705 7925
rect 6740 7825 6760 7925
rect 6795 7825 6800 7925
rect 6700 7810 6800 7825
rect 6950 7925 7050 7940
rect 6950 7825 6955 7925
rect 6990 7825 7010 7925
rect 7045 7825 7050 7925
rect 6950 7810 7050 7825
rect 7200 7925 7300 7940
rect 7200 7825 7205 7925
rect 7240 7825 7260 7925
rect 7295 7825 7300 7925
rect 7200 7810 7300 7825
rect 7450 7925 7550 7940
rect 7450 7825 7455 7925
rect 7490 7825 7510 7925
rect 7545 7825 7550 7925
rect 7450 7810 7550 7825
rect 7700 7925 7800 7940
rect 7700 7825 7705 7925
rect 7740 7825 7760 7925
rect 7795 7825 7800 7925
rect 7700 7810 7800 7825
rect 7950 7925 8000 7940
rect 7950 7825 7955 7925
rect 7990 7825 8000 7925
rect 7950 7810 8000 7825
rect 0 7800 60 7810
rect 190 7800 310 7810
rect 440 7800 560 7810
rect 690 7800 810 7810
rect 940 7800 1060 7810
rect 1190 7800 1310 7810
rect 1440 7800 1560 7810
rect 1690 7800 1810 7810
rect 1940 7800 2060 7810
rect 2190 7800 2310 7810
rect 2440 7800 2560 7810
rect 2690 7800 2810 7810
rect 2940 7800 3060 7810
rect 3190 7800 3310 7810
rect 3440 7800 3560 7810
rect 3690 7800 3810 7810
rect 3940 7800 4060 7810
rect 4190 7800 4310 7810
rect 4440 7800 4560 7810
rect 4690 7800 4810 7810
rect 4940 7800 5060 7810
rect 5190 7800 5310 7810
rect 5440 7800 5560 7810
rect 5690 7800 5810 7810
rect 5940 7800 6060 7810
rect 6190 7800 6310 7810
rect 6440 7800 6560 7810
rect 6690 7800 6810 7810
rect 6940 7800 7060 7810
rect 7190 7800 7310 7810
rect 7440 7800 7560 7810
rect 7690 7800 7810 7810
rect 7940 7800 8000 7810
rect 0 7795 8000 7800
rect 0 7760 75 7795
rect 175 7760 325 7795
rect 425 7760 575 7795
rect 675 7760 825 7795
rect 925 7760 1075 7795
rect 1175 7760 1325 7795
rect 1425 7760 1575 7795
rect 1675 7760 1825 7795
rect 1925 7760 2075 7795
rect 2175 7760 2325 7795
rect 2425 7760 2575 7795
rect 2675 7760 2825 7795
rect 2925 7760 3075 7795
rect 3175 7760 3325 7795
rect 3425 7760 3575 7795
rect 3675 7760 3825 7795
rect 3925 7760 4075 7795
rect 4175 7760 4325 7795
rect 4425 7760 4575 7795
rect 4675 7760 4825 7795
rect 4925 7760 5075 7795
rect 5175 7760 5325 7795
rect 5425 7760 5575 7795
rect 5675 7760 5825 7795
rect 5925 7760 6075 7795
rect 6175 7760 6325 7795
rect 6425 7760 6575 7795
rect 6675 7760 6825 7795
rect 6925 7760 7075 7795
rect 7175 7760 7325 7795
rect 7425 7760 7575 7795
rect 7675 7760 7825 7795
rect 7925 7760 8000 7795
rect 0 7740 8000 7760
rect 0 7705 75 7740
rect 175 7705 325 7740
rect 425 7705 575 7740
rect 675 7705 825 7740
rect 925 7705 1075 7740
rect 1175 7705 1325 7740
rect 1425 7705 1575 7740
rect 1675 7705 1825 7740
rect 1925 7705 2075 7740
rect 2175 7705 2325 7740
rect 2425 7705 2575 7740
rect 2675 7705 2825 7740
rect 2925 7705 3075 7740
rect 3175 7705 3325 7740
rect 3425 7705 3575 7740
rect 3675 7705 3825 7740
rect 3925 7705 4075 7740
rect 4175 7705 4325 7740
rect 4425 7705 4575 7740
rect 4675 7705 4825 7740
rect 4925 7705 5075 7740
rect 5175 7705 5325 7740
rect 5425 7705 5575 7740
rect 5675 7705 5825 7740
rect 5925 7705 6075 7740
rect 6175 7705 6325 7740
rect 6425 7705 6575 7740
rect 6675 7705 6825 7740
rect 6925 7705 7075 7740
rect 7175 7705 7325 7740
rect 7425 7705 7575 7740
rect 7675 7705 7825 7740
rect 7925 7705 8000 7740
rect 0 7700 8000 7705
rect 0 7690 60 7700
rect 190 7690 310 7700
rect 440 7690 560 7700
rect 690 7690 810 7700
rect 940 7690 1060 7700
rect 1190 7690 1310 7700
rect 1440 7690 1560 7700
rect 1690 7690 1810 7700
rect 1940 7690 2060 7700
rect 2190 7690 2310 7700
rect 2440 7690 2560 7700
rect 2690 7690 2810 7700
rect 2940 7690 3060 7700
rect 3190 7690 3310 7700
rect 3440 7690 3560 7700
rect 3690 7690 3810 7700
rect 3940 7690 4060 7700
rect 4190 7690 4310 7700
rect 4440 7690 4560 7700
rect 4690 7690 4810 7700
rect 4940 7690 5060 7700
rect 5190 7690 5310 7700
rect 5440 7690 5560 7700
rect 5690 7690 5810 7700
rect 5940 7690 6060 7700
rect 6190 7690 6310 7700
rect 6440 7690 6560 7700
rect 6690 7690 6810 7700
rect 6940 7690 7060 7700
rect 7190 7690 7310 7700
rect 7440 7690 7560 7700
rect 7690 7690 7810 7700
rect 7940 7690 8000 7700
rect 0 7675 50 7690
rect 0 7575 10 7675
rect 45 7575 50 7675
rect 0 7560 50 7575
rect 200 7675 300 7690
rect 200 7575 205 7675
rect 240 7575 260 7675
rect 295 7575 300 7675
rect 200 7560 300 7575
rect 450 7675 550 7690
rect 450 7575 455 7675
rect 490 7575 510 7675
rect 545 7575 550 7675
rect 450 7560 550 7575
rect 700 7675 800 7690
rect 700 7575 705 7675
rect 740 7575 760 7675
rect 795 7575 800 7675
rect 700 7560 800 7575
rect 950 7675 1050 7690
rect 950 7575 955 7675
rect 990 7575 1010 7675
rect 1045 7575 1050 7675
rect 950 7560 1050 7575
rect 1200 7675 1300 7690
rect 1200 7575 1205 7675
rect 1240 7575 1260 7675
rect 1295 7575 1300 7675
rect 1200 7560 1300 7575
rect 1450 7675 1550 7690
rect 1450 7575 1455 7675
rect 1490 7575 1510 7675
rect 1545 7575 1550 7675
rect 1450 7560 1550 7575
rect 1700 7675 1800 7690
rect 1700 7575 1705 7675
rect 1740 7575 1760 7675
rect 1795 7575 1800 7675
rect 1700 7560 1800 7575
rect 1950 7675 2050 7690
rect 1950 7575 1955 7675
rect 1990 7575 2010 7675
rect 2045 7575 2050 7675
rect 1950 7560 2050 7575
rect 2200 7675 2300 7690
rect 2200 7575 2205 7675
rect 2240 7575 2260 7675
rect 2295 7575 2300 7675
rect 2200 7560 2300 7575
rect 2450 7675 2550 7690
rect 2450 7575 2455 7675
rect 2490 7575 2510 7675
rect 2545 7575 2550 7675
rect 2450 7560 2550 7575
rect 2700 7675 2800 7690
rect 2700 7575 2705 7675
rect 2740 7575 2760 7675
rect 2795 7575 2800 7675
rect 2700 7560 2800 7575
rect 2950 7675 3050 7690
rect 2950 7575 2955 7675
rect 2990 7575 3010 7675
rect 3045 7575 3050 7675
rect 2950 7560 3050 7575
rect 3200 7675 3300 7690
rect 3200 7575 3205 7675
rect 3240 7575 3260 7675
rect 3295 7575 3300 7675
rect 3200 7560 3300 7575
rect 3450 7675 3550 7690
rect 3450 7575 3455 7675
rect 3490 7575 3510 7675
rect 3545 7575 3550 7675
rect 3450 7560 3550 7575
rect 3700 7675 3800 7690
rect 3700 7575 3705 7675
rect 3740 7575 3760 7675
rect 3795 7575 3800 7675
rect 3700 7560 3800 7575
rect 3950 7675 4050 7690
rect 3950 7575 3955 7675
rect 3990 7575 4010 7675
rect 4045 7575 4050 7675
rect 3950 7560 4050 7575
rect 4200 7675 4300 7690
rect 4200 7575 4205 7675
rect 4240 7575 4260 7675
rect 4295 7575 4300 7675
rect 4200 7560 4300 7575
rect 4450 7675 4550 7690
rect 4450 7575 4455 7675
rect 4490 7575 4510 7675
rect 4545 7575 4550 7675
rect 4450 7560 4550 7575
rect 4700 7675 4800 7690
rect 4700 7575 4705 7675
rect 4740 7575 4760 7675
rect 4795 7575 4800 7675
rect 4700 7560 4800 7575
rect 4950 7675 5050 7690
rect 4950 7575 4955 7675
rect 4990 7575 5010 7675
rect 5045 7575 5050 7675
rect 4950 7560 5050 7575
rect 5200 7675 5300 7690
rect 5200 7575 5205 7675
rect 5240 7575 5260 7675
rect 5295 7575 5300 7675
rect 5200 7560 5300 7575
rect 5450 7675 5550 7690
rect 5450 7575 5455 7675
rect 5490 7575 5510 7675
rect 5545 7575 5550 7675
rect 5450 7560 5550 7575
rect 5700 7675 5800 7690
rect 5700 7575 5705 7675
rect 5740 7575 5760 7675
rect 5795 7575 5800 7675
rect 5700 7560 5800 7575
rect 5950 7675 6050 7690
rect 5950 7575 5955 7675
rect 5990 7575 6010 7675
rect 6045 7575 6050 7675
rect 5950 7560 6050 7575
rect 6200 7675 6300 7690
rect 6200 7575 6205 7675
rect 6240 7575 6260 7675
rect 6295 7575 6300 7675
rect 6200 7560 6300 7575
rect 6450 7675 6550 7690
rect 6450 7575 6455 7675
rect 6490 7575 6510 7675
rect 6545 7575 6550 7675
rect 6450 7560 6550 7575
rect 6700 7675 6800 7690
rect 6700 7575 6705 7675
rect 6740 7575 6760 7675
rect 6795 7575 6800 7675
rect 6700 7560 6800 7575
rect 6950 7675 7050 7690
rect 6950 7575 6955 7675
rect 6990 7575 7010 7675
rect 7045 7575 7050 7675
rect 6950 7560 7050 7575
rect 7200 7675 7300 7690
rect 7200 7575 7205 7675
rect 7240 7575 7260 7675
rect 7295 7575 7300 7675
rect 7200 7560 7300 7575
rect 7450 7675 7550 7690
rect 7450 7575 7455 7675
rect 7490 7575 7510 7675
rect 7545 7575 7550 7675
rect 7450 7560 7550 7575
rect 7700 7675 7800 7690
rect 7700 7575 7705 7675
rect 7740 7575 7760 7675
rect 7795 7575 7800 7675
rect 7700 7560 7800 7575
rect 7950 7675 8000 7690
rect 7950 7575 7955 7675
rect 7990 7575 8000 7675
rect 7950 7560 8000 7575
rect 0 7550 60 7560
rect 190 7550 310 7560
rect 440 7550 560 7560
rect 690 7550 810 7560
rect 940 7550 1060 7560
rect 1190 7550 1310 7560
rect 1440 7550 1560 7560
rect 1690 7550 1810 7560
rect 1940 7550 2060 7560
rect 2190 7550 2310 7560
rect 2440 7550 2560 7560
rect 2690 7550 2810 7560
rect 2940 7550 3060 7560
rect 3190 7550 3310 7560
rect 3440 7550 3560 7560
rect 3690 7550 3810 7560
rect 3940 7550 4060 7560
rect 4190 7550 4310 7560
rect 4440 7550 4560 7560
rect 4690 7550 4810 7560
rect 4940 7550 5060 7560
rect 5190 7550 5310 7560
rect 5440 7550 5560 7560
rect 5690 7550 5810 7560
rect 5940 7550 6060 7560
rect 6190 7550 6310 7560
rect 6440 7550 6560 7560
rect 6690 7550 6810 7560
rect 6940 7550 7060 7560
rect 7190 7550 7310 7560
rect 7440 7550 7560 7560
rect 7690 7550 7810 7560
rect 7940 7550 8000 7560
rect 0 7545 8000 7550
rect 0 7510 75 7545
rect 175 7510 325 7545
rect 425 7510 575 7545
rect 675 7510 825 7545
rect 925 7510 1075 7545
rect 1175 7510 1325 7545
rect 1425 7510 1575 7545
rect 1675 7510 1825 7545
rect 1925 7510 2075 7545
rect 2175 7510 2325 7545
rect 2425 7510 2575 7545
rect 2675 7510 2825 7545
rect 2925 7510 3075 7545
rect 3175 7510 3325 7545
rect 3425 7510 3575 7545
rect 3675 7510 3825 7545
rect 3925 7510 4075 7545
rect 4175 7510 4325 7545
rect 4425 7510 4575 7545
rect 4675 7510 4825 7545
rect 4925 7510 5075 7545
rect 5175 7510 5325 7545
rect 5425 7510 5575 7545
rect 5675 7510 5825 7545
rect 5925 7510 6075 7545
rect 6175 7510 6325 7545
rect 6425 7510 6575 7545
rect 6675 7510 6825 7545
rect 6925 7510 7075 7545
rect 7175 7510 7325 7545
rect 7425 7510 7575 7545
rect 7675 7510 7825 7545
rect 7925 7510 8000 7545
rect 0 7490 8000 7510
rect 0 7455 75 7490
rect 175 7455 325 7490
rect 425 7455 575 7490
rect 675 7455 825 7490
rect 925 7455 1075 7490
rect 1175 7455 1325 7490
rect 1425 7455 1575 7490
rect 1675 7455 1825 7490
rect 1925 7455 2075 7490
rect 2175 7455 2325 7490
rect 2425 7455 2575 7490
rect 2675 7455 2825 7490
rect 2925 7455 3075 7490
rect 3175 7455 3325 7490
rect 3425 7455 3575 7490
rect 3675 7455 3825 7490
rect 3925 7455 4075 7490
rect 4175 7455 4325 7490
rect 4425 7455 4575 7490
rect 4675 7455 4825 7490
rect 4925 7455 5075 7490
rect 5175 7455 5325 7490
rect 5425 7455 5575 7490
rect 5675 7455 5825 7490
rect 5925 7455 6075 7490
rect 6175 7455 6325 7490
rect 6425 7455 6575 7490
rect 6675 7455 6825 7490
rect 6925 7455 7075 7490
rect 7175 7455 7325 7490
rect 7425 7455 7575 7490
rect 7675 7455 7825 7490
rect 7925 7455 8000 7490
rect 0 7450 8000 7455
rect 0 7440 60 7450
rect 190 7440 310 7450
rect 440 7440 560 7450
rect 690 7440 810 7450
rect 940 7440 1060 7450
rect 1190 7440 1310 7450
rect 1440 7440 1560 7450
rect 1690 7440 1810 7450
rect 1940 7440 2060 7450
rect 2190 7440 2310 7450
rect 2440 7440 2560 7450
rect 2690 7440 2810 7450
rect 2940 7440 3060 7450
rect 3190 7440 3310 7450
rect 3440 7440 3560 7450
rect 3690 7440 3810 7450
rect 3940 7440 4060 7450
rect 4190 7440 4310 7450
rect 4440 7440 4560 7450
rect 4690 7440 4810 7450
rect 4940 7440 5060 7450
rect 5190 7440 5310 7450
rect 5440 7440 5560 7450
rect 5690 7440 5810 7450
rect 5940 7440 6060 7450
rect 6190 7440 6310 7450
rect 6440 7440 6560 7450
rect 6690 7440 6810 7450
rect 6940 7440 7060 7450
rect 7190 7440 7310 7450
rect 7440 7440 7560 7450
rect 7690 7440 7810 7450
rect 7940 7440 8000 7450
rect 0 7425 50 7440
rect 0 7325 10 7425
rect 45 7325 50 7425
rect 0 7310 50 7325
rect 200 7425 300 7440
rect 200 7325 205 7425
rect 240 7325 260 7425
rect 295 7325 300 7425
rect 200 7310 300 7325
rect 450 7425 550 7440
rect 450 7325 455 7425
rect 490 7325 510 7425
rect 545 7325 550 7425
rect 450 7310 550 7325
rect 700 7425 800 7440
rect 700 7325 705 7425
rect 740 7325 760 7425
rect 795 7325 800 7425
rect 700 7310 800 7325
rect 950 7425 1050 7440
rect 950 7325 955 7425
rect 990 7325 1010 7425
rect 1045 7325 1050 7425
rect 950 7310 1050 7325
rect 1200 7425 1300 7440
rect 1200 7325 1205 7425
rect 1240 7325 1260 7425
rect 1295 7325 1300 7425
rect 1200 7310 1300 7325
rect 1450 7425 1550 7440
rect 1450 7325 1455 7425
rect 1490 7325 1510 7425
rect 1545 7325 1550 7425
rect 1450 7310 1550 7325
rect 1700 7425 1800 7440
rect 1700 7325 1705 7425
rect 1740 7325 1760 7425
rect 1795 7325 1800 7425
rect 1700 7310 1800 7325
rect 1950 7425 2050 7440
rect 1950 7325 1955 7425
rect 1990 7325 2010 7425
rect 2045 7325 2050 7425
rect 1950 7310 2050 7325
rect 2200 7425 2300 7440
rect 2200 7325 2205 7425
rect 2240 7325 2260 7425
rect 2295 7325 2300 7425
rect 2200 7310 2300 7325
rect 2450 7425 2550 7440
rect 2450 7325 2455 7425
rect 2490 7325 2510 7425
rect 2545 7325 2550 7425
rect 2450 7310 2550 7325
rect 2700 7425 2800 7440
rect 2700 7325 2705 7425
rect 2740 7325 2760 7425
rect 2795 7325 2800 7425
rect 2700 7310 2800 7325
rect 2950 7425 3050 7440
rect 2950 7325 2955 7425
rect 2990 7325 3010 7425
rect 3045 7325 3050 7425
rect 2950 7310 3050 7325
rect 3200 7425 3300 7440
rect 3200 7325 3205 7425
rect 3240 7325 3260 7425
rect 3295 7325 3300 7425
rect 3200 7310 3300 7325
rect 3450 7425 3550 7440
rect 3450 7325 3455 7425
rect 3490 7325 3510 7425
rect 3545 7325 3550 7425
rect 3450 7310 3550 7325
rect 3700 7425 3800 7440
rect 3700 7325 3705 7425
rect 3740 7325 3760 7425
rect 3795 7325 3800 7425
rect 3700 7310 3800 7325
rect 3950 7425 4050 7440
rect 3950 7325 3955 7425
rect 3990 7325 4010 7425
rect 4045 7325 4050 7425
rect 3950 7310 4050 7325
rect 4200 7425 4300 7440
rect 4200 7325 4205 7425
rect 4240 7325 4260 7425
rect 4295 7325 4300 7425
rect 4200 7310 4300 7325
rect 4450 7425 4550 7440
rect 4450 7325 4455 7425
rect 4490 7325 4510 7425
rect 4545 7325 4550 7425
rect 4450 7310 4550 7325
rect 4700 7425 4800 7440
rect 4700 7325 4705 7425
rect 4740 7325 4760 7425
rect 4795 7325 4800 7425
rect 4700 7310 4800 7325
rect 4950 7425 5050 7440
rect 4950 7325 4955 7425
rect 4990 7325 5010 7425
rect 5045 7325 5050 7425
rect 4950 7310 5050 7325
rect 5200 7425 5300 7440
rect 5200 7325 5205 7425
rect 5240 7325 5260 7425
rect 5295 7325 5300 7425
rect 5200 7310 5300 7325
rect 5450 7425 5550 7440
rect 5450 7325 5455 7425
rect 5490 7325 5510 7425
rect 5545 7325 5550 7425
rect 5450 7310 5550 7325
rect 5700 7425 5800 7440
rect 5700 7325 5705 7425
rect 5740 7325 5760 7425
rect 5795 7325 5800 7425
rect 5700 7310 5800 7325
rect 5950 7425 6050 7440
rect 5950 7325 5955 7425
rect 5990 7325 6010 7425
rect 6045 7325 6050 7425
rect 5950 7310 6050 7325
rect 6200 7425 6300 7440
rect 6200 7325 6205 7425
rect 6240 7325 6260 7425
rect 6295 7325 6300 7425
rect 6200 7310 6300 7325
rect 6450 7425 6550 7440
rect 6450 7325 6455 7425
rect 6490 7325 6510 7425
rect 6545 7325 6550 7425
rect 6450 7310 6550 7325
rect 6700 7425 6800 7440
rect 6700 7325 6705 7425
rect 6740 7325 6760 7425
rect 6795 7325 6800 7425
rect 6700 7310 6800 7325
rect 6950 7425 7050 7440
rect 6950 7325 6955 7425
rect 6990 7325 7010 7425
rect 7045 7325 7050 7425
rect 6950 7310 7050 7325
rect 7200 7425 7300 7440
rect 7200 7325 7205 7425
rect 7240 7325 7260 7425
rect 7295 7325 7300 7425
rect 7200 7310 7300 7325
rect 7450 7425 7550 7440
rect 7450 7325 7455 7425
rect 7490 7325 7510 7425
rect 7545 7325 7550 7425
rect 7450 7310 7550 7325
rect 7700 7425 7800 7440
rect 7700 7325 7705 7425
rect 7740 7325 7760 7425
rect 7795 7325 7800 7425
rect 7700 7310 7800 7325
rect 7950 7425 8000 7440
rect 7950 7325 7955 7425
rect 7990 7325 8000 7425
rect 7950 7310 8000 7325
rect 0 7300 60 7310
rect 190 7300 310 7310
rect 440 7300 560 7310
rect 690 7300 810 7310
rect 940 7300 1060 7310
rect 1190 7300 1310 7310
rect 1440 7300 1560 7310
rect 1690 7300 1810 7310
rect 1940 7300 2060 7310
rect 2190 7300 2310 7310
rect 2440 7300 2560 7310
rect 2690 7300 2810 7310
rect 2940 7300 3060 7310
rect 3190 7300 3310 7310
rect 3440 7300 3560 7310
rect 3690 7300 3810 7310
rect 3940 7300 4060 7310
rect 4190 7300 4310 7310
rect 4440 7300 4560 7310
rect 4690 7300 4810 7310
rect 4940 7300 5060 7310
rect 5190 7300 5310 7310
rect 5440 7300 5560 7310
rect 5690 7300 5810 7310
rect 5940 7300 6060 7310
rect 6190 7300 6310 7310
rect 6440 7300 6560 7310
rect 6690 7300 6810 7310
rect 6940 7300 7060 7310
rect 7190 7300 7310 7310
rect 7440 7300 7560 7310
rect 7690 7300 7810 7310
rect 7940 7300 8000 7310
rect 0 7295 8000 7300
rect 0 7260 75 7295
rect 175 7260 325 7295
rect 425 7260 575 7295
rect 675 7260 825 7295
rect 925 7260 1075 7295
rect 1175 7260 1325 7295
rect 1425 7260 1575 7295
rect 1675 7260 1825 7295
rect 1925 7260 2075 7295
rect 2175 7260 2325 7295
rect 2425 7260 2575 7295
rect 2675 7260 2825 7295
rect 2925 7260 3075 7295
rect 3175 7260 3325 7295
rect 3425 7260 3575 7295
rect 3675 7260 3825 7295
rect 3925 7260 4075 7295
rect 4175 7260 4325 7295
rect 4425 7260 4575 7295
rect 4675 7260 4825 7295
rect 4925 7260 5075 7295
rect 5175 7260 5325 7295
rect 5425 7260 5575 7295
rect 5675 7260 5825 7295
rect 5925 7260 6075 7295
rect 6175 7260 6325 7295
rect 6425 7260 6575 7295
rect 6675 7260 6825 7295
rect 6925 7260 7075 7295
rect 7175 7260 7325 7295
rect 7425 7260 7575 7295
rect 7675 7260 7825 7295
rect 7925 7260 8000 7295
rect 0 7240 8000 7260
rect 0 7205 75 7240
rect 175 7205 325 7240
rect 425 7205 575 7240
rect 675 7205 825 7240
rect 925 7205 1075 7240
rect 1175 7205 1325 7240
rect 1425 7205 1575 7240
rect 1675 7205 1825 7240
rect 1925 7205 2075 7240
rect 2175 7205 2325 7240
rect 2425 7205 2575 7240
rect 2675 7205 2825 7240
rect 2925 7205 3075 7240
rect 3175 7205 3325 7240
rect 3425 7205 3575 7240
rect 3675 7205 3825 7240
rect 3925 7205 4075 7240
rect 4175 7205 4325 7240
rect 4425 7205 4575 7240
rect 4675 7205 4825 7240
rect 4925 7205 5075 7240
rect 5175 7205 5325 7240
rect 5425 7205 5575 7240
rect 5675 7205 5825 7240
rect 5925 7205 6075 7240
rect 6175 7205 6325 7240
rect 6425 7205 6575 7240
rect 6675 7205 6825 7240
rect 6925 7205 7075 7240
rect 7175 7205 7325 7240
rect 7425 7205 7575 7240
rect 7675 7205 7825 7240
rect 7925 7205 8000 7240
rect 0 7200 8000 7205
rect 0 7190 60 7200
rect 190 7190 310 7200
rect 440 7190 560 7200
rect 690 7190 810 7200
rect 940 7190 1060 7200
rect 1190 7190 1310 7200
rect 1440 7190 1560 7200
rect 1690 7190 1810 7200
rect 1940 7190 2060 7200
rect 2190 7190 2310 7200
rect 2440 7190 2560 7200
rect 2690 7190 2810 7200
rect 2940 7190 3060 7200
rect 3190 7190 3310 7200
rect 3440 7190 3560 7200
rect 3690 7190 3810 7200
rect 3940 7190 4060 7200
rect 4190 7190 4310 7200
rect 4440 7190 4560 7200
rect 4690 7190 4810 7200
rect 4940 7190 5060 7200
rect 5190 7190 5310 7200
rect 5440 7190 5560 7200
rect 5690 7190 5810 7200
rect 5940 7190 6060 7200
rect 6190 7190 6310 7200
rect 6440 7190 6560 7200
rect 6690 7190 6810 7200
rect 6940 7190 7060 7200
rect 7190 7190 7310 7200
rect 7440 7190 7560 7200
rect 7690 7190 7810 7200
rect 7940 7190 8000 7200
rect 0 7175 50 7190
rect 0 7075 10 7175
rect 45 7075 50 7175
rect 0 7060 50 7075
rect 200 7175 300 7190
rect 200 7075 205 7175
rect 240 7075 260 7175
rect 295 7075 300 7175
rect 200 7060 300 7075
rect 450 7175 550 7190
rect 450 7075 455 7175
rect 490 7075 510 7175
rect 545 7075 550 7175
rect 450 7060 550 7075
rect 700 7175 800 7190
rect 700 7075 705 7175
rect 740 7075 760 7175
rect 795 7075 800 7175
rect 700 7060 800 7075
rect 950 7175 1050 7190
rect 950 7075 955 7175
rect 990 7075 1010 7175
rect 1045 7075 1050 7175
rect 950 7060 1050 7075
rect 1200 7175 1300 7190
rect 1200 7075 1205 7175
rect 1240 7075 1260 7175
rect 1295 7075 1300 7175
rect 1200 7060 1300 7075
rect 1450 7175 1550 7190
rect 1450 7075 1455 7175
rect 1490 7075 1510 7175
rect 1545 7075 1550 7175
rect 1450 7060 1550 7075
rect 1700 7175 1800 7190
rect 1700 7075 1705 7175
rect 1740 7075 1760 7175
rect 1795 7075 1800 7175
rect 1700 7060 1800 7075
rect 1950 7175 2050 7190
rect 1950 7075 1955 7175
rect 1990 7075 2010 7175
rect 2045 7075 2050 7175
rect 1950 7060 2050 7075
rect 2200 7175 2300 7190
rect 2200 7075 2205 7175
rect 2240 7075 2260 7175
rect 2295 7075 2300 7175
rect 2200 7060 2300 7075
rect 2450 7175 2550 7190
rect 2450 7075 2455 7175
rect 2490 7075 2510 7175
rect 2545 7075 2550 7175
rect 2450 7060 2550 7075
rect 2700 7175 2800 7190
rect 2700 7075 2705 7175
rect 2740 7075 2760 7175
rect 2795 7075 2800 7175
rect 2700 7060 2800 7075
rect 2950 7175 3050 7190
rect 2950 7075 2955 7175
rect 2990 7075 3010 7175
rect 3045 7075 3050 7175
rect 2950 7060 3050 7075
rect 3200 7175 3300 7190
rect 3200 7075 3205 7175
rect 3240 7075 3260 7175
rect 3295 7075 3300 7175
rect 3200 7060 3300 7075
rect 3450 7175 3550 7190
rect 3450 7075 3455 7175
rect 3490 7075 3510 7175
rect 3545 7075 3550 7175
rect 3450 7060 3550 7075
rect 3700 7175 3800 7190
rect 3700 7075 3705 7175
rect 3740 7075 3760 7175
rect 3795 7075 3800 7175
rect 3700 7060 3800 7075
rect 3950 7175 4050 7190
rect 3950 7075 3955 7175
rect 3990 7075 4010 7175
rect 4045 7075 4050 7175
rect 3950 7060 4050 7075
rect 4200 7175 4300 7190
rect 4200 7075 4205 7175
rect 4240 7075 4260 7175
rect 4295 7075 4300 7175
rect 4200 7060 4300 7075
rect 4450 7175 4550 7190
rect 4450 7075 4455 7175
rect 4490 7075 4510 7175
rect 4545 7075 4550 7175
rect 4450 7060 4550 7075
rect 4700 7175 4800 7190
rect 4700 7075 4705 7175
rect 4740 7075 4760 7175
rect 4795 7075 4800 7175
rect 4700 7060 4800 7075
rect 4950 7175 5050 7190
rect 4950 7075 4955 7175
rect 4990 7075 5010 7175
rect 5045 7075 5050 7175
rect 4950 7060 5050 7075
rect 5200 7175 5300 7190
rect 5200 7075 5205 7175
rect 5240 7075 5260 7175
rect 5295 7075 5300 7175
rect 5200 7060 5300 7075
rect 5450 7175 5550 7190
rect 5450 7075 5455 7175
rect 5490 7075 5510 7175
rect 5545 7075 5550 7175
rect 5450 7060 5550 7075
rect 5700 7175 5800 7190
rect 5700 7075 5705 7175
rect 5740 7075 5760 7175
rect 5795 7075 5800 7175
rect 5700 7060 5800 7075
rect 5950 7175 6050 7190
rect 5950 7075 5955 7175
rect 5990 7075 6010 7175
rect 6045 7075 6050 7175
rect 5950 7060 6050 7075
rect 6200 7175 6300 7190
rect 6200 7075 6205 7175
rect 6240 7075 6260 7175
rect 6295 7075 6300 7175
rect 6200 7060 6300 7075
rect 6450 7175 6550 7190
rect 6450 7075 6455 7175
rect 6490 7075 6510 7175
rect 6545 7075 6550 7175
rect 6450 7060 6550 7075
rect 6700 7175 6800 7190
rect 6700 7075 6705 7175
rect 6740 7075 6760 7175
rect 6795 7075 6800 7175
rect 6700 7060 6800 7075
rect 6950 7175 7050 7190
rect 6950 7075 6955 7175
rect 6990 7075 7010 7175
rect 7045 7075 7050 7175
rect 6950 7060 7050 7075
rect 7200 7175 7300 7190
rect 7200 7075 7205 7175
rect 7240 7075 7260 7175
rect 7295 7075 7300 7175
rect 7200 7060 7300 7075
rect 7450 7175 7550 7190
rect 7450 7075 7455 7175
rect 7490 7075 7510 7175
rect 7545 7075 7550 7175
rect 7450 7060 7550 7075
rect 7700 7175 7800 7190
rect 7700 7075 7705 7175
rect 7740 7075 7760 7175
rect 7795 7075 7800 7175
rect 7700 7060 7800 7075
rect 7950 7175 8000 7190
rect 7950 7075 7955 7175
rect 7990 7075 8000 7175
rect 7950 7060 8000 7075
rect 0 7050 60 7060
rect 190 7050 310 7060
rect 440 7050 560 7060
rect 690 7050 810 7060
rect 940 7050 1060 7060
rect 1190 7050 1310 7060
rect 1440 7050 1560 7060
rect 1690 7050 1810 7060
rect 1940 7050 2060 7060
rect 2190 7050 2310 7060
rect 2440 7050 2560 7060
rect 2690 7050 2810 7060
rect 2940 7050 3060 7060
rect 3190 7050 3310 7060
rect 3440 7050 3560 7060
rect 3690 7050 3810 7060
rect 3940 7050 4060 7060
rect 4190 7050 4310 7060
rect 4440 7050 4560 7060
rect 4690 7050 4810 7060
rect 4940 7050 5060 7060
rect 5190 7050 5310 7060
rect 5440 7050 5560 7060
rect 5690 7050 5810 7060
rect 5940 7050 6060 7060
rect 6190 7050 6310 7060
rect 6440 7050 6560 7060
rect 6690 7050 6810 7060
rect 6940 7050 7060 7060
rect 7190 7050 7310 7060
rect 7440 7050 7560 7060
rect 7690 7050 7810 7060
rect 7940 7050 8000 7060
rect 0 7045 8000 7050
rect 0 7010 75 7045
rect 175 7010 325 7045
rect 425 7010 575 7045
rect 675 7010 825 7045
rect 925 7010 1075 7045
rect 1175 7010 1325 7045
rect 1425 7010 1575 7045
rect 1675 7010 1825 7045
rect 1925 7010 2075 7045
rect 2175 7010 2325 7045
rect 2425 7010 2575 7045
rect 2675 7010 2825 7045
rect 2925 7010 3075 7045
rect 3175 7010 3325 7045
rect 3425 7010 3575 7045
rect 3675 7010 3825 7045
rect 3925 7010 4075 7045
rect 4175 7010 4325 7045
rect 4425 7010 4575 7045
rect 4675 7010 4825 7045
rect 4925 7010 5075 7045
rect 5175 7010 5325 7045
rect 5425 7010 5575 7045
rect 5675 7010 5825 7045
rect 5925 7010 6075 7045
rect 6175 7010 6325 7045
rect 6425 7010 6575 7045
rect 6675 7010 6825 7045
rect 6925 7010 7075 7045
rect 7175 7010 7325 7045
rect 7425 7010 7575 7045
rect 7675 7010 7825 7045
rect 7925 7010 8000 7045
rect 0 6990 8000 7010
rect 0 6955 75 6990
rect 175 6955 325 6990
rect 425 6955 575 6990
rect 675 6955 825 6990
rect 925 6955 1075 6990
rect 1175 6955 1325 6990
rect 1425 6955 1575 6990
rect 1675 6955 1825 6990
rect 1925 6955 2075 6990
rect 2175 6955 2325 6990
rect 2425 6955 2575 6990
rect 2675 6955 2825 6990
rect 2925 6955 3075 6990
rect 3175 6955 3325 6990
rect 3425 6955 3575 6990
rect 3675 6955 3825 6990
rect 3925 6955 4075 6990
rect 4175 6955 4325 6990
rect 4425 6955 4575 6990
rect 4675 6955 4825 6990
rect 4925 6955 5075 6990
rect 5175 6955 5325 6990
rect 5425 6955 5575 6990
rect 5675 6955 5825 6990
rect 5925 6955 6075 6990
rect 6175 6955 6325 6990
rect 6425 6955 6575 6990
rect 6675 6955 6825 6990
rect 6925 6955 7075 6990
rect 7175 6955 7325 6990
rect 7425 6955 7575 6990
rect 7675 6955 7825 6990
rect 7925 6955 8000 6990
rect 0 6950 8000 6955
rect 0 6940 60 6950
rect 190 6940 310 6950
rect 440 6940 560 6950
rect 690 6940 810 6950
rect 940 6940 1060 6950
rect 1190 6940 1310 6950
rect 1440 6940 1560 6950
rect 1690 6940 1810 6950
rect 1940 6940 2060 6950
rect 2190 6940 2310 6950
rect 2440 6940 2560 6950
rect 2690 6940 2810 6950
rect 2940 6940 3060 6950
rect 3190 6940 3310 6950
rect 3440 6940 3560 6950
rect 3690 6940 3810 6950
rect 3940 6940 4060 6950
rect 4190 6940 4310 6950
rect 4440 6940 4560 6950
rect 4690 6940 4810 6950
rect 4940 6940 5060 6950
rect 5190 6940 5310 6950
rect 5440 6940 5560 6950
rect 5690 6940 5810 6950
rect 5940 6940 6060 6950
rect 6190 6940 6310 6950
rect 6440 6940 6560 6950
rect 6690 6940 6810 6950
rect 6940 6940 7060 6950
rect 7190 6940 7310 6950
rect 7440 6940 7560 6950
rect 7690 6940 7810 6950
rect 7940 6940 8000 6950
rect 0 6925 50 6940
rect 0 6825 10 6925
rect 45 6825 50 6925
rect 0 6810 50 6825
rect 200 6925 300 6940
rect 200 6825 205 6925
rect 240 6825 260 6925
rect 295 6825 300 6925
rect 200 6810 300 6825
rect 450 6925 550 6940
rect 450 6825 455 6925
rect 490 6825 510 6925
rect 545 6825 550 6925
rect 450 6810 550 6825
rect 700 6925 800 6940
rect 700 6825 705 6925
rect 740 6825 760 6925
rect 795 6825 800 6925
rect 700 6810 800 6825
rect 950 6925 1050 6940
rect 950 6825 955 6925
rect 990 6825 1010 6925
rect 1045 6825 1050 6925
rect 950 6810 1050 6825
rect 1200 6925 1300 6940
rect 1200 6825 1205 6925
rect 1240 6825 1260 6925
rect 1295 6825 1300 6925
rect 1200 6810 1300 6825
rect 1450 6925 1550 6940
rect 1450 6825 1455 6925
rect 1490 6825 1510 6925
rect 1545 6825 1550 6925
rect 1450 6810 1550 6825
rect 1700 6925 1800 6940
rect 1700 6825 1705 6925
rect 1740 6825 1760 6925
rect 1795 6825 1800 6925
rect 1700 6810 1800 6825
rect 1950 6925 2050 6940
rect 1950 6825 1955 6925
rect 1990 6825 2010 6925
rect 2045 6825 2050 6925
rect 1950 6810 2050 6825
rect 2200 6925 2300 6940
rect 2200 6825 2205 6925
rect 2240 6825 2260 6925
rect 2295 6825 2300 6925
rect 2200 6810 2300 6825
rect 2450 6925 2550 6940
rect 2450 6825 2455 6925
rect 2490 6825 2510 6925
rect 2545 6825 2550 6925
rect 2450 6810 2550 6825
rect 2700 6925 2800 6940
rect 2700 6825 2705 6925
rect 2740 6825 2760 6925
rect 2795 6825 2800 6925
rect 2700 6810 2800 6825
rect 2950 6925 3050 6940
rect 2950 6825 2955 6925
rect 2990 6825 3010 6925
rect 3045 6825 3050 6925
rect 2950 6810 3050 6825
rect 3200 6925 3300 6940
rect 3200 6825 3205 6925
rect 3240 6825 3260 6925
rect 3295 6825 3300 6925
rect 3200 6810 3300 6825
rect 3450 6925 3550 6940
rect 3450 6825 3455 6925
rect 3490 6825 3510 6925
rect 3545 6825 3550 6925
rect 3450 6810 3550 6825
rect 3700 6925 3800 6940
rect 3700 6825 3705 6925
rect 3740 6825 3760 6925
rect 3795 6825 3800 6925
rect 3700 6810 3800 6825
rect 3950 6925 4050 6940
rect 3950 6825 3955 6925
rect 3990 6825 4010 6925
rect 4045 6825 4050 6925
rect 3950 6810 4050 6825
rect 4200 6925 4300 6940
rect 4200 6825 4205 6925
rect 4240 6825 4260 6925
rect 4295 6825 4300 6925
rect 4200 6810 4300 6825
rect 4450 6925 4550 6940
rect 4450 6825 4455 6925
rect 4490 6825 4510 6925
rect 4545 6825 4550 6925
rect 4450 6810 4550 6825
rect 4700 6925 4800 6940
rect 4700 6825 4705 6925
rect 4740 6825 4760 6925
rect 4795 6825 4800 6925
rect 4700 6810 4800 6825
rect 4950 6925 5050 6940
rect 4950 6825 4955 6925
rect 4990 6825 5010 6925
rect 5045 6825 5050 6925
rect 4950 6810 5050 6825
rect 5200 6925 5300 6940
rect 5200 6825 5205 6925
rect 5240 6825 5260 6925
rect 5295 6825 5300 6925
rect 5200 6810 5300 6825
rect 5450 6925 5550 6940
rect 5450 6825 5455 6925
rect 5490 6825 5510 6925
rect 5545 6825 5550 6925
rect 5450 6810 5550 6825
rect 5700 6925 5800 6940
rect 5700 6825 5705 6925
rect 5740 6825 5760 6925
rect 5795 6825 5800 6925
rect 5700 6810 5800 6825
rect 5950 6925 6050 6940
rect 5950 6825 5955 6925
rect 5990 6825 6010 6925
rect 6045 6825 6050 6925
rect 5950 6810 6050 6825
rect 6200 6925 6300 6940
rect 6200 6825 6205 6925
rect 6240 6825 6260 6925
rect 6295 6825 6300 6925
rect 6200 6810 6300 6825
rect 6450 6925 6550 6940
rect 6450 6825 6455 6925
rect 6490 6825 6510 6925
rect 6545 6825 6550 6925
rect 6450 6810 6550 6825
rect 6700 6925 6800 6940
rect 6700 6825 6705 6925
rect 6740 6825 6760 6925
rect 6795 6825 6800 6925
rect 6700 6810 6800 6825
rect 6950 6925 7050 6940
rect 6950 6825 6955 6925
rect 6990 6825 7010 6925
rect 7045 6825 7050 6925
rect 6950 6810 7050 6825
rect 7200 6925 7300 6940
rect 7200 6825 7205 6925
rect 7240 6825 7260 6925
rect 7295 6825 7300 6925
rect 7200 6810 7300 6825
rect 7450 6925 7550 6940
rect 7450 6825 7455 6925
rect 7490 6825 7510 6925
rect 7545 6825 7550 6925
rect 7450 6810 7550 6825
rect 7700 6925 7800 6940
rect 7700 6825 7705 6925
rect 7740 6825 7760 6925
rect 7795 6825 7800 6925
rect 7700 6810 7800 6825
rect 7950 6925 8000 6940
rect 7950 6825 7955 6925
rect 7990 6825 8000 6925
rect 7950 6810 8000 6825
rect 0 6800 60 6810
rect 190 6800 310 6810
rect 440 6800 560 6810
rect 690 6800 810 6810
rect 940 6800 1060 6810
rect 1190 6800 1310 6810
rect 1440 6800 1560 6810
rect 1690 6800 1810 6810
rect 1940 6800 2060 6810
rect 2190 6800 2310 6810
rect 2440 6800 2560 6810
rect 2690 6800 2810 6810
rect 2940 6800 3060 6810
rect 3190 6800 3310 6810
rect 3440 6800 3560 6810
rect 3690 6800 3810 6810
rect 3940 6800 4060 6810
rect 4190 6800 4310 6810
rect 4440 6800 4560 6810
rect 4690 6800 4810 6810
rect 4940 6800 5060 6810
rect 5190 6800 5310 6810
rect 5440 6800 5560 6810
rect 5690 6800 5810 6810
rect 5940 6800 6060 6810
rect 6190 6800 6310 6810
rect 6440 6800 6560 6810
rect 6690 6800 6810 6810
rect 6940 6800 7060 6810
rect 7190 6800 7310 6810
rect 7440 6800 7560 6810
rect 7690 6800 7810 6810
rect 7940 6800 8000 6810
rect 0 6795 8000 6800
rect 0 6760 75 6795
rect 175 6760 325 6795
rect 425 6760 575 6795
rect 675 6760 825 6795
rect 925 6760 1075 6795
rect 1175 6760 1325 6795
rect 1425 6760 1575 6795
rect 1675 6760 1825 6795
rect 1925 6760 2075 6795
rect 2175 6760 2325 6795
rect 2425 6760 2575 6795
rect 2675 6760 2825 6795
rect 2925 6760 3075 6795
rect 3175 6760 3325 6795
rect 3425 6760 3575 6795
rect 3675 6760 3825 6795
rect 3925 6760 4075 6795
rect 4175 6760 4325 6795
rect 4425 6760 4575 6795
rect 4675 6760 4825 6795
rect 4925 6760 5075 6795
rect 5175 6760 5325 6795
rect 5425 6760 5575 6795
rect 5675 6760 5825 6795
rect 5925 6760 6075 6795
rect 6175 6760 6325 6795
rect 6425 6760 6575 6795
rect 6675 6760 6825 6795
rect 6925 6760 7075 6795
rect 7175 6760 7325 6795
rect 7425 6760 7575 6795
rect 7675 6760 7825 6795
rect 7925 6760 8000 6795
rect 0 6740 8000 6760
rect 0 6705 75 6740
rect 175 6705 325 6740
rect 425 6705 575 6740
rect 675 6705 825 6740
rect 925 6705 1075 6740
rect 1175 6705 1325 6740
rect 1425 6705 1575 6740
rect 1675 6705 1825 6740
rect 1925 6705 2075 6740
rect 2175 6705 2325 6740
rect 2425 6705 2575 6740
rect 2675 6705 2825 6740
rect 2925 6705 3075 6740
rect 3175 6705 3325 6740
rect 3425 6705 3575 6740
rect 3675 6705 3825 6740
rect 3925 6705 4075 6740
rect 4175 6705 4325 6740
rect 4425 6705 4575 6740
rect 4675 6705 4825 6740
rect 4925 6705 5075 6740
rect 5175 6705 5325 6740
rect 5425 6705 5575 6740
rect 5675 6705 5825 6740
rect 5925 6705 6075 6740
rect 6175 6705 6325 6740
rect 6425 6705 6575 6740
rect 6675 6705 6825 6740
rect 6925 6705 7075 6740
rect 7175 6705 7325 6740
rect 7425 6705 7575 6740
rect 7675 6705 7825 6740
rect 7925 6705 8000 6740
rect 0 6700 8000 6705
rect 0 6690 60 6700
rect 190 6690 310 6700
rect 440 6690 560 6700
rect 690 6690 810 6700
rect 940 6690 1060 6700
rect 1190 6690 1310 6700
rect 1440 6690 1560 6700
rect 1690 6690 1810 6700
rect 1940 6690 2060 6700
rect 2190 6690 2310 6700
rect 2440 6690 2560 6700
rect 2690 6690 2810 6700
rect 2940 6690 3060 6700
rect 3190 6690 3310 6700
rect 3440 6690 3560 6700
rect 3690 6690 3810 6700
rect 3940 6690 4060 6700
rect 4190 6690 4310 6700
rect 4440 6690 4560 6700
rect 4690 6690 4810 6700
rect 4940 6690 5060 6700
rect 5190 6690 5310 6700
rect 5440 6690 5560 6700
rect 5690 6690 5810 6700
rect 5940 6690 6060 6700
rect 6190 6690 6310 6700
rect 6440 6690 6560 6700
rect 6690 6690 6810 6700
rect 6940 6690 7060 6700
rect 7190 6690 7310 6700
rect 7440 6690 7560 6700
rect 7690 6690 7810 6700
rect 7940 6690 8000 6700
rect 0 6675 50 6690
rect 0 6575 10 6675
rect 45 6575 50 6675
rect 0 6560 50 6575
rect 200 6675 300 6690
rect 200 6575 205 6675
rect 240 6575 260 6675
rect 295 6575 300 6675
rect 200 6560 300 6575
rect 450 6675 550 6690
rect 450 6575 455 6675
rect 490 6575 510 6675
rect 545 6575 550 6675
rect 450 6560 550 6575
rect 700 6675 800 6690
rect 700 6575 705 6675
rect 740 6575 760 6675
rect 795 6575 800 6675
rect 700 6560 800 6575
rect 950 6675 1050 6690
rect 950 6575 955 6675
rect 990 6575 1010 6675
rect 1045 6575 1050 6675
rect 950 6560 1050 6575
rect 1200 6675 1300 6690
rect 1200 6575 1205 6675
rect 1240 6575 1260 6675
rect 1295 6575 1300 6675
rect 1200 6560 1300 6575
rect 1450 6675 1550 6690
rect 1450 6575 1455 6675
rect 1490 6575 1510 6675
rect 1545 6575 1550 6675
rect 1450 6560 1550 6575
rect 1700 6675 1800 6690
rect 1700 6575 1705 6675
rect 1740 6575 1760 6675
rect 1795 6575 1800 6675
rect 1700 6560 1800 6575
rect 1950 6675 2050 6690
rect 1950 6575 1955 6675
rect 1990 6575 2010 6675
rect 2045 6575 2050 6675
rect 1950 6560 2050 6575
rect 2200 6675 2300 6690
rect 2200 6575 2205 6675
rect 2240 6575 2260 6675
rect 2295 6575 2300 6675
rect 2200 6560 2300 6575
rect 2450 6675 2550 6690
rect 2450 6575 2455 6675
rect 2490 6575 2510 6675
rect 2545 6575 2550 6675
rect 2450 6560 2550 6575
rect 2700 6675 2800 6690
rect 2700 6575 2705 6675
rect 2740 6575 2760 6675
rect 2795 6575 2800 6675
rect 2700 6560 2800 6575
rect 2950 6675 3050 6690
rect 2950 6575 2955 6675
rect 2990 6575 3010 6675
rect 3045 6575 3050 6675
rect 2950 6560 3050 6575
rect 3200 6675 3300 6690
rect 3200 6575 3205 6675
rect 3240 6575 3260 6675
rect 3295 6575 3300 6675
rect 3200 6560 3300 6575
rect 3450 6675 3550 6690
rect 3450 6575 3455 6675
rect 3490 6575 3510 6675
rect 3545 6575 3550 6675
rect 3450 6560 3550 6575
rect 3700 6675 3800 6690
rect 3700 6575 3705 6675
rect 3740 6575 3760 6675
rect 3795 6575 3800 6675
rect 3700 6560 3800 6575
rect 3950 6675 4050 6690
rect 3950 6575 3955 6675
rect 3990 6575 4010 6675
rect 4045 6575 4050 6675
rect 3950 6560 4050 6575
rect 4200 6675 4300 6690
rect 4200 6575 4205 6675
rect 4240 6575 4260 6675
rect 4295 6575 4300 6675
rect 4200 6560 4300 6575
rect 4450 6675 4550 6690
rect 4450 6575 4455 6675
rect 4490 6575 4510 6675
rect 4545 6575 4550 6675
rect 4450 6560 4550 6575
rect 4700 6675 4800 6690
rect 4700 6575 4705 6675
rect 4740 6575 4760 6675
rect 4795 6575 4800 6675
rect 4700 6560 4800 6575
rect 4950 6675 5050 6690
rect 4950 6575 4955 6675
rect 4990 6575 5010 6675
rect 5045 6575 5050 6675
rect 4950 6560 5050 6575
rect 5200 6675 5300 6690
rect 5200 6575 5205 6675
rect 5240 6575 5260 6675
rect 5295 6575 5300 6675
rect 5200 6560 5300 6575
rect 5450 6675 5550 6690
rect 5450 6575 5455 6675
rect 5490 6575 5510 6675
rect 5545 6575 5550 6675
rect 5450 6560 5550 6575
rect 5700 6675 5800 6690
rect 5700 6575 5705 6675
rect 5740 6575 5760 6675
rect 5795 6575 5800 6675
rect 5700 6560 5800 6575
rect 5950 6675 6050 6690
rect 5950 6575 5955 6675
rect 5990 6575 6010 6675
rect 6045 6575 6050 6675
rect 5950 6560 6050 6575
rect 6200 6675 6300 6690
rect 6200 6575 6205 6675
rect 6240 6575 6260 6675
rect 6295 6575 6300 6675
rect 6200 6560 6300 6575
rect 6450 6675 6550 6690
rect 6450 6575 6455 6675
rect 6490 6575 6510 6675
rect 6545 6575 6550 6675
rect 6450 6560 6550 6575
rect 6700 6675 6800 6690
rect 6700 6575 6705 6675
rect 6740 6575 6760 6675
rect 6795 6575 6800 6675
rect 6700 6560 6800 6575
rect 6950 6675 7050 6690
rect 6950 6575 6955 6675
rect 6990 6575 7010 6675
rect 7045 6575 7050 6675
rect 6950 6560 7050 6575
rect 7200 6675 7300 6690
rect 7200 6575 7205 6675
rect 7240 6575 7260 6675
rect 7295 6575 7300 6675
rect 7200 6560 7300 6575
rect 7450 6675 7550 6690
rect 7450 6575 7455 6675
rect 7490 6575 7510 6675
rect 7545 6575 7550 6675
rect 7450 6560 7550 6575
rect 7700 6675 7800 6690
rect 7700 6575 7705 6675
rect 7740 6575 7760 6675
rect 7795 6575 7800 6675
rect 7700 6560 7800 6575
rect 7950 6675 8000 6690
rect 7950 6575 7955 6675
rect 7990 6575 8000 6675
rect 7950 6560 8000 6575
rect 0 6550 60 6560
rect 190 6550 310 6560
rect 440 6550 560 6560
rect 690 6550 810 6560
rect 940 6550 1060 6560
rect 1190 6550 1310 6560
rect 1440 6550 1560 6560
rect 1690 6550 1810 6560
rect 1940 6550 2060 6560
rect 2190 6550 2310 6560
rect 2440 6550 2560 6560
rect 2690 6550 2810 6560
rect 2940 6550 3060 6560
rect 3190 6550 3310 6560
rect 3440 6550 3560 6560
rect 3690 6550 3810 6560
rect 3940 6550 4060 6560
rect 4190 6550 4310 6560
rect 4440 6550 4560 6560
rect 4690 6550 4810 6560
rect 4940 6550 5060 6560
rect 5190 6550 5310 6560
rect 5440 6550 5560 6560
rect 5690 6550 5810 6560
rect 5940 6550 6060 6560
rect 6190 6550 6310 6560
rect 6440 6550 6560 6560
rect 6690 6550 6810 6560
rect 6940 6550 7060 6560
rect 7190 6550 7310 6560
rect 7440 6550 7560 6560
rect 7690 6550 7810 6560
rect 7940 6550 8000 6560
rect 0 6545 8000 6550
rect 0 6510 75 6545
rect 175 6510 325 6545
rect 425 6510 575 6545
rect 675 6510 825 6545
rect 925 6510 1075 6545
rect 1175 6510 1325 6545
rect 1425 6510 1575 6545
rect 1675 6510 1825 6545
rect 1925 6510 2075 6545
rect 2175 6510 2325 6545
rect 2425 6510 2575 6545
rect 2675 6510 2825 6545
rect 2925 6510 3075 6545
rect 3175 6510 3325 6545
rect 3425 6510 3575 6545
rect 3675 6510 3825 6545
rect 3925 6510 4075 6545
rect 4175 6510 4325 6545
rect 4425 6510 4575 6545
rect 4675 6510 4825 6545
rect 4925 6510 5075 6545
rect 5175 6510 5325 6545
rect 5425 6510 5575 6545
rect 5675 6510 5825 6545
rect 5925 6510 6075 6545
rect 6175 6510 6325 6545
rect 6425 6510 6575 6545
rect 6675 6510 6825 6545
rect 6925 6510 7075 6545
rect 7175 6510 7325 6545
rect 7425 6510 7575 6545
rect 7675 6510 7825 6545
rect 7925 6510 8000 6545
rect 0 6490 8000 6510
rect 0 6455 75 6490
rect 175 6455 325 6490
rect 425 6455 575 6490
rect 675 6455 825 6490
rect 925 6455 1075 6490
rect 1175 6455 1325 6490
rect 1425 6455 1575 6490
rect 1675 6455 1825 6490
rect 1925 6455 2075 6490
rect 2175 6455 2325 6490
rect 2425 6455 2575 6490
rect 2675 6455 2825 6490
rect 2925 6455 3075 6490
rect 3175 6455 3325 6490
rect 3425 6455 3575 6490
rect 3675 6455 3825 6490
rect 3925 6455 4075 6490
rect 4175 6455 4325 6490
rect 4425 6455 4575 6490
rect 4675 6455 4825 6490
rect 4925 6455 5075 6490
rect 5175 6455 5325 6490
rect 5425 6455 5575 6490
rect 5675 6455 5825 6490
rect 5925 6455 6075 6490
rect 6175 6455 6325 6490
rect 6425 6455 6575 6490
rect 6675 6455 6825 6490
rect 6925 6455 7075 6490
rect 7175 6455 7325 6490
rect 7425 6455 7575 6490
rect 7675 6455 7825 6490
rect 7925 6455 8000 6490
rect 0 6450 8000 6455
rect 0 6440 60 6450
rect 190 6440 310 6450
rect 440 6440 560 6450
rect 690 6440 810 6450
rect 940 6440 1060 6450
rect 1190 6440 1310 6450
rect 1440 6440 1560 6450
rect 1690 6440 1810 6450
rect 1940 6440 2060 6450
rect 2190 6440 2310 6450
rect 2440 6440 2560 6450
rect 2690 6440 2810 6450
rect 2940 6440 3060 6450
rect 3190 6440 3310 6450
rect 3440 6440 3560 6450
rect 3690 6440 3810 6450
rect 3940 6440 4060 6450
rect 4190 6440 4310 6450
rect 4440 6440 4560 6450
rect 4690 6440 4810 6450
rect 4940 6440 5060 6450
rect 5190 6440 5310 6450
rect 5440 6440 5560 6450
rect 5690 6440 5810 6450
rect 5940 6440 6060 6450
rect 6190 6440 6310 6450
rect 6440 6440 6560 6450
rect 6690 6440 6810 6450
rect 6940 6440 7060 6450
rect 7190 6440 7310 6450
rect 7440 6440 7560 6450
rect 7690 6440 7810 6450
rect 7940 6440 8000 6450
rect 0 6425 50 6440
rect 0 6325 10 6425
rect 45 6325 50 6425
rect 0 6310 50 6325
rect 200 6425 300 6440
rect 200 6325 205 6425
rect 240 6325 260 6425
rect 295 6325 300 6425
rect 200 6310 300 6325
rect 450 6425 550 6440
rect 450 6325 455 6425
rect 490 6325 510 6425
rect 545 6325 550 6425
rect 450 6310 550 6325
rect 700 6425 800 6440
rect 700 6325 705 6425
rect 740 6325 760 6425
rect 795 6325 800 6425
rect 700 6310 800 6325
rect 950 6425 1050 6440
rect 950 6325 955 6425
rect 990 6325 1010 6425
rect 1045 6325 1050 6425
rect 950 6310 1050 6325
rect 1200 6425 1300 6440
rect 1200 6325 1205 6425
rect 1240 6325 1260 6425
rect 1295 6325 1300 6425
rect 1200 6310 1300 6325
rect 1450 6425 1550 6440
rect 1450 6325 1455 6425
rect 1490 6325 1510 6425
rect 1545 6325 1550 6425
rect 1450 6310 1550 6325
rect 1700 6425 1800 6440
rect 1700 6325 1705 6425
rect 1740 6325 1760 6425
rect 1795 6325 1800 6425
rect 1700 6310 1800 6325
rect 1950 6425 2050 6440
rect 1950 6325 1955 6425
rect 1990 6325 2010 6425
rect 2045 6325 2050 6425
rect 1950 6310 2050 6325
rect 2200 6425 2300 6440
rect 2200 6325 2205 6425
rect 2240 6325 2260 6425
rect 2295 6325 2300 6425
rect 2200 6310 2300 6325
rect 2450 6425 2550 6440
rect 2450 6325 2455 6425
rect 2490 6325 2510 6425
rect 2545 6325 2550 6425
rect 2450 6310 2550 6325
rect 2700 6425 2800 6440
rect 2700 6325 2705 6425
rect 2740 6325 2760 6425
rect 2795 6325 2800 6425
rect 2700 6310 2800 6325
rect 2950 6425 3050 6440
rect 2950 6325 2955 6425
rect 2990 6325 3010 6425
rect 3045 6325 3050 6425
rect 2950 6310 3050 6325
rect 3200 6425 3300 6440
rect 3200 6325 3205 6425
rect 3240 6325 3260 6425
rect 3295 6325 3300 6425
rect 3200 6310 3300 6325
rect 3450 6425 3550 6440
rect 3450 6325 3455 6425
rect 3490 6325 3510 6425
rect 3545 6325 3550 6425
rect 3450 6310 3550 6325
rect 3700 6425 3800 6440
rect 3700 6325 3705 6425
rect 3740 6325 3760 6425
rect 3795 6325 3800 6425
rect 3700 6310 3800 6325
rect 3950 6425 4050 6440
rect 3950 6325 3955 6425
rect 3990 6325 4010 6425
rect 4045 6325 4050 6425
rect 3950 6310 4050 6325
rect 4200 6425 4300 6440
rect 4200 6325 4205 6425
rect 4240 6325 4260 6425
rect 4295 6325 4300 6425
rect 4200 6310 4300 6325
rect 4450 6425 4550 6440
rect 4450 6325 4455 6425
rect 4490 6325 4510 6425
rect 4545 6325 4550 6425
rect 4450 6310 4550 6325
rect 4700 6425 4800 6440
rect 4700 6325 4705 6425
rect 4740 6325 4760 6425
rect 4795 6325 4800 6425
rect 4700 6310 4800 6325
rect 4950 6425 5050 6440
rect 4950 6325 4955 6425
rect 4990 6325 5010 6425
rect 5045 6325 5050 6425
rect 4950 6310 5050 6325
rect 5200 6425 5300 6440
rect 5200 6325 5205 6425
rect 5240 6325 5260 6425
rect 5295 6325 5300 6425
rect 5200 6310 5300 6325
rect 5450 6425 5550 6440
rect 5450 6325 5455 6425
rect 5490 6325 5510 6425
rect 5545 6325 5550 6425
rect 5450 6310 5550 6325
rect 5700 6425 5800 6440
rect 5700 6325 5705 6425
rect 5740 6325 5760 6425
rect 5795 6325 5800 6425
rect 5700 6310 5800 6325
rect 5950 6425 6050 6440
rect 5950 6325 5955 6425
rect 5990 6325 6010 6425
rect 6045 6325 6050 6425
rect 5950 6310 6050 6325
rect 6200 6425 6300 6440
rect 6200 6325 6205 6425
rect 6240 6325 6260 6425
rect 6295 6325 6300 6425
rect 6200 6310 6300 6325
rect 6450 6425 6550 6440
rect 6450 6325 6455 6425
rect 6490 6325 6510 6425
rect 6545 6325 6550 6425
rect 6450 6310 6550 6325
rect 6700 6425 6800 6440
rect 6700 6325 6705 6425
rect 6740 6325 6760 6425
rect 6795 6325 6800 6425
rect 6700 6310 6800 6325
rect 6950 6425 7050 6440
rect 6950 6325 6955 6425
rect 6990 6325 7010 6425
rect 7045 6325 7050 6425
rect 6950 6310 7050 6325
rect 7200 6425 7300 6440
rect 7200 6325 7205 6425
rect 7240 6325 7260 6425
rect 7295 6325 7300 6425
rect 7200 6310 7300 6325
rect 7450 6425 7550 6440
rect 7450 6325 7455 6425
rect 7490 6325 7510 6425
rect 7545 6325 7550 6425
rect 7450 6310 7550 6325
rect 7700 6425 7800 6440
rect 7700 6325 7705 6425
rect 7740 6325 7760 6425
rect 7795 6325 7800 6425
rect 7700 6310 7800 6325
rect 7950 6425 8000 6440
rect 7950 6325 7955 6425
rect 7990 6325 8000 6425
rect 7950 6310 8000 6325
rect 0 6300 60 6310
rect 190 6300 310 6310
rect 440 6300 560 6310
rect 690 6300 810 6310
rect 940 6300 1060 6310
rect 1190 6300 1310 6310
rect 1440 6300 1560 6310
rect 1690 6300 1810 6310
rect 1940 6300 2060 6310
rect 2190 6300 2310 6310
rect 2440 6300 2560 6310
rect 2690 6300 2810 6310
rect 2940 6300 3060 6310
rect 3190 6300 3310 6310
rect 3440 6300 3560 6310
rect 3690 6300 3810 6310
rect 3940 6300 4060 6310
rect 4190 6300 4310 6310
rect 4440 6300 4560 6310
rect 4690 6300 4810 6310
rect 4940 6300 5060 6310
rect 5190 6300 5310 6310
rect 5440 6300 5560 6310
rect 5690 6300 5810 6310
rect 5940 6300 6060 6310
rect 6190 6300 6310 6310
rect 6440 6300 6560 6310
rect 6690 6300 6810 6310
rect 6940 6300 7060 6310
rect 7190 6300 7310 6310
rect 7440 6300 7560 6310
rect 7690 6300 7810 6310
rect 7940 6300 8000 6310
rect 0 6295 8000 6300
rect 0 6260 75 6295
rect 175 6260 325 6295
rect 425 6260 575 6295
rect 675 6260 825 6295
rect 925 6260 1075 6295
rect 1175 6260 1325 6295
rect 1425 6260 1575 6295
rect 1675 6260 1825 6295
rect 1925 6260 2075 6295
rect 2175 6260 2325 6295
rect 2425 6260 2575 6295
rect 2675 6260 2825 6295
rect 2925 6260 3075 6295
rect 3175 6260 3325 6295
rect 3425 6260 3575 6295
rect 3675 6260 3825 6295
rect 3925 6260 4075 6295
rect 4175 6260 4325 6295
rect 4425 6260 4575 6295
rect 4675 6260 4825 6295
rect 4925 6260 5075 6295
rect 5175 6260 5325 6295
rect 5425 6260 5575 6295
rect 5675 6260 5825 6295
rect 5925 6260 6075 6295
rect 6175 6260 6325 6295
rect 6425 6260 6575 6295
rect 6675 6260 6825 6295
rect 6925 6260 7075 6295
rect 7175 6260 7325 6295
rect 7425 6260 7575 6295
rect 7675 6260 7825 6295
rect 7925 6260 8000 6295
rect 0 6240 8000 6260
rect 0 6205 75 6240
rect 175 6205 325 6240
rect 425 6205 575 6240
rect 675 6205 825 6240
rect 925 6205 1075 6240
rect 1175 6205 1325 6240
rect 1425 6205 1575 6240
rect 1675 6205 1825 6240
rect 1925 6205 2075 6240
rect 2175 6205 2325 6240
rect 2425 6205 2575 6240
rect 2675 6205 2825 6240
rect 2925 6205 3075 6240
rect 3175 6205 3325 6240
rect 3425 6205 3575 6240
rect 3675 6205 3825 6240
rect 3925 6205 4075 6240
rect 4175 6205 4325 6240
rect 4425 6205 4575 6240
rect 4675 6205 4825 6240
rect 4925 6205 5075 6240
rect 5175 6205 5325 6240
rect 5425 6205 5575 6240
rect 5675 6205 5825 6240
rect 5925 6205 6075 6240
rect 6175 6205 6325 6240
rect 6425 6205 6575 6240
rect 6675 6205 6825 6240
rect 6925 6205 7075 6240
rect 7175 6205 7325 6240
rect 7425 6205 7575 6240
rect 7675 6205 7825 6240
rect 7925 6205 8000 6240
rect 0 6200 8000 6205
rect 0 6190 60 6200
rect 190 6190 310 6200
rect 440 6190 560 6200
rect 690 6190 810 6200
rect 940 6190 1060 6200
rect 1190 6190 1310 6200
rect 1440 6190 1560 6200
rect 1690 6190 1810 6200
rect 1940 6190 2060 6200
rect 2190 6190 2310 6200
rect 2440 6190 2560 6200
rect 2690 6190 2810 6200
rect 2940 6190 3060 6200
rect 3190 6190 3310 6200
rect 3440 6190 3560 6200
rect 3690 6190 3810 6200
rect 3940 6190 4060 6200
rect 4190 6190 4310 6200
rect 4440 6190 4560 6200
rect 4690 6190 4810 6200
rect 4940 6190 5060 6200
rect 5190 6190 5310 6200
rect 5440 6190 5560 6200
rect 5690 6190 5810 6200
rect 5940 6190 6060 6200
rect 6190 6190 6310 6200
rect 6440 6190 6560 6200
rect 6690 6190 6810 6200
rect 6940 6190 7060 6200
rect 7190 6190 7310 6200
rect 7440 6190 7560 6200
rect 7690 6190 7810 6200
rect 7940 6190 8000 6200
rect 0 6175 50 6190
rect 0 6075 10 6175
rect 45 6075 50 6175
rect 0 6060 50 6075
rect 200 6175 300 6190
rect 200 6075 205 6175
rect 240 6075 260 6175
rect 295 6075 300 6175
rect 200 6060 300 6075
rect 450 6175 550 6190
rect 450 6075 455 6175
rect 490 6075 510 6175
rect 545 6075 550 6175
rect 450 6060 550 6075
rect 700 6175 800 6190
rect 700 6075 705 6175
rect 740 6075 760 6175
rect 795 6075 800 6175
rect 700 6060 800 6075
rect 950 6175 1050 6190
rect 950 6075 955 6175
rect 990 6075 1010 6175
rect 1045 6075 1050 6175
rect 950 6060 1050 6075
rect 1200 6175 1300 6190
rect 1200 6075 1205 6175
rect 1240 6075 1260 6175
rect 1295 6075 1300 6175
rect 1200 6060 1300 6075
rect 1450 6175 1550 6190
rect 1450 6075 1455 6175
rect 1490 6075 1510 6175
rect 1545 6075 1550 6175
rect 1450 6060 1550 6075
rect 1700 6175 1800 6190
rect 1700 6075 1705 6175
rect 1740 6075 1760 6175
rect 1795 6075 1800 6175
rect 1700 6060 1800 6075
rect 1950 6175 2050 6190
rect 1950 6075 1955 6175
rect 1990 6075 2010 6175
rect 2045 6075 2050 6175
rect 1950 6060 2050 6075
rect 2200 6175 2300 6190
rect 2200 6075 2205 6175
rect 2240 6075 2260 6175
rect 2295 6075 2300 6175
rect 2200 6060 2300 6075
rect 2450 6175 2550 6190
rect 2450 6075 2455 6175
rect 2490 6075 2510 6175
rect 2545 6075 2550 6175
rect 2450 6060 2550 6075
rect 2700 6175 2800 6190
rect 2700 6075 2705 6175
rect 2740 6075 2760 6175
rect 2795 6075 2800 6175
rect 2700 6060 2800 6075
rect 2950 6175 3050 6190
rect 2950 6075 2955 6175
rect 2990 6075 3010 6175
rect 3045 6075 3050 6175
rect 2950 6060 3050 6075
rect 3200 6175 3300 6190
rect 3200 6075 3205 6175
rect 3240 6075 3260 6175
rect 3295 6075 3300 6175
rect 3200 6060 3300 6075
rect 3450 6175 3550 6190
rect 3450 6075 3455 6175
rect 3490 6075 3510 6175
rect 3545 6075 3550 6175
rect 3450 6060 3550 6075
rect 3700 6175 3800 6190
rect 3700 6075 3705 6175
rect 3740 6075 3760 6175
rect 3795 6075 3800 6175
rect 3700 6060 3800 6075
rect 3950 6175 4050 6190
rect 3950 6075 3955 6175
rect 3990 6075 4010 6175
rect 4045 6075 4050 6175
rect 3950 6060 4050 6075
rect 4200 6175 4300 6190
rect 4200 6075 4205 6175
rect 4240 6075 4260 6175
rect 4295 6075 4300 6175
rect 4200 6060 4300 6075
rect 4450 6175 4550 6190
rect 4450 6075 4455 6175
rect 4490 6075 4510 6175
rect 4545 6075 4550 6175
rect 4450 6060 4550 6075
rect 4700 6175 4800 6190
rect 4700 6075 4705 6175
rect 4740 6075 4760 6175
rect 4795 6075 4800 6175
rect 4700 6060 4800 6075
rect 4950 6175 5050 6190
rect 4950 6075 4955 6175
rect 4990 6075 5010 6175
rect 5045 6075 5050 6175
rect 4950 6060 5050 6075
rect 5200 6175 5300 6190
rect 5200 6075 5205 6175
rect 5240 6075 5260 6175
rect 5295 6075 5300 6175
rect 5200 6060 5300 6075
rect 5450 6175 5550 6190
rect 5450 6075 5455 6175
rect 5490 6075 5510 6175
rect 5545 6075 5550 6175
rect 5450 6060 5550 6075
rect 5700 6175 5800 6190
rect 5700 6075 5705 6175
rect 5740 6075 5760 6175
rect 5795 6075 5800 6175
rect 5700 6060 5800 6075
rect 5950 6175 6050 6190
rect 5950 6075 5955 6175
rect 5990 6075 6010 6175
rect 6045 6075 6050 6175
rect 5950 6060 6050 6075
rect 6200 6175 6300 6190
rect 6200 6075 6205 6175
rect 6240 6075 6260 6175
rect 6295 6075 6300 6175
rect 6200 6060 6300 6075
rect 6450 6175 6550 6190
rect 6450 6075 6455 6175
rect 6490 6075 6510 6175
rect 6545 6075 6550 6175
rect 6450 6060 6550 6075
rect 6700 6175 6800 6190
rect 6700 6075 6705 6175
rect 6740 6075 6760 6175
rect 6795 6075 6800 6175
rect 6700 6060 6800 6075
rect 6950 6175 7050 6190
rect 6950 6075 6955 6175
rect 6990 6075 7010 6175
rect 7045 6075 7050 6175
rect 6950 6060 7050 6075
rect 7200 6175 7300 6190
rect 7200 6075 7205 6175
rect 7240 6075 7260 6175
rect 7295 6075 7300 6175
rect 7200 6060 7300 6075
rect 7450 6175 7550 6190
rect 7450 6075 7455 6175
rect 7490 6075 7510 6175
rect 7545 6075 7550 6175
rect 7450 6060 7550 6075
rect 7700 6175 7800 6190
rect 7700 6075 7705 6175
rect 7740 6075 7760 6175
rect 7795 6075 7800 6175
rect 7700 6060 7800 6075
rect 7950 6175 8000 6190
rect 7950 6075 7955 6175
rect 7990 6075 8000 6175
rect 7950 6060 8000 6075
rect 0 6050 60 6060
rect 190 6050 310 6060
rect 440 6050 560 6060
rect 690 6050 810 6060
rect 940 6050 1060 6060
rect 1190 6050 1310 6060
rect 1440 6050 1560 6060
rect 1690 6050 1810 6060
rect 1940 6050 2060 6060
rect 2190 6050 2310 6060
rect 2440 6050 2560 6060
rect 2690 6050 2810 6060
rect 2940 6050 3060 6060
rect 3190 6050 3310 6060
rect 3440 6050 3560 6060
rect 3690 6050 3810 6060
rect 3940 6050 4060 6060
rect 4190 6050 4310 6060
rect 4440 6050 4560 6060
rect 4690 6050 4810 6060
rect 4940 6050 5060 6060
rect 5190 6050 5310 6060
rect 5440 6050 5560 6060
rect 5690 6050 5810 6060
rect 5940 6050 6060 6060
rect 6190 6050 6310 6060
rect 6440 6050 6560 6060
rect 6690 6050 6810 6060
rect 6940 6050 7060 6060
rect 7190 6050 7310 6060
rect 7440 6050 7560 6060
rect 7690 6050 7810 6060
rect 7940 6050 8000 6060
rect 0 6045 8000 6050
rect 0 6010 75 6045
rect 175 6010 325 6045
rect 425 6010 575 6045
rect 675 6010 825 6045
rect 925 6010 1075 6045
rect 1175 6010 1325 6045
rect 1425 6010 1575 6045
rect 1675 6010 1825 6045
rect 1925 6010 2075 6045
rect 2175 6010 2325 6045
rect 2425 6010 2575 6045
rect 2675 6010 2825 6045
rect 2925 6010 3075 6045
rect 3175 6010 3325 6045
rect 3425 6010 3575 6045
rect 3675 6010 3825 6045
rect 3925 6010 4075 6045
rect 4175 6010 4325 6045
rect 4425 6010 4575 6045
rect 4675 6010 4825 6045
rect 4925 6010 5075 6045
rect 5175 6010 5325 6045
rect 5425 6010 5575 6045
rect 5675 6010 5825 6045
rect 5925 6010 6075 6045
rect 6175 6010 6325 6045
rect 6425 6010 6575 6045
rect 6675 6010 6825 6045
rect 6925 6010 7075 6045
rect 7175 6010 7325 6045
rect 7425 6010 7575 6045
rect 7675 6010 7825 6045
rect 7925 6010 8000 6045
rect 0 5990 8000 6010
rect 0 5955 75 5990
rect 175 5955 325 5990
rect 425 5955 575 5990
rect 675 5955 825 5990
rect 925 5955 1075 5990
rect 1175 5955 1325 5990
rect 1425 5955 1575 5990
rect 1675 5955 1825 5990
rect 1925 5955 2075 5990
rect 2175 5955 2325 5990
rect 2425 5955 2575 5990
rect 2675 5955 2825 5990
rect 2925 5955 3075 5990
rect 3175 5955 3325 5990
rect 3425 5955 3575 5990
rect 3675 5955 3825 5990
rect 3925 5955 4075 5990
rect 4175 5955 4325 5990
rect 4425 5955 4575 5990
rect 4675 5955 4825 5990
rect 4925 5955 5075 5990
rect 5175 5955 5325 5990
rect 5425 5955 5575 5990
rect 5675 5955 5825 5990
rect 5925 5955 6075 5990
rect 6175 5955 6325 5990
rect 6425 5955 6575 5990
rect 6675 5955 6825 5990
rect 6925 5955 7075 5990
rect 7175 5955 7325 5990
rect 7425 5955 7575 5990
rect 7675 5955 7825 5990
rect 7925 5955 8000 5990
rect 0 5950 8000 5955
rect 0 5940 60 5950
rect 190 5940 310 5950
rect 440 5940 560 5950
rect 690 5940 810 5950
rect 940 5940 1060 5950
rect 1190 5940 1310 5950
rect 1440 5940 1560 5950
rect 1690 5940 1810 5950
rect 1940 5940 2060 5950
rect 2190 5940 2310 5950
rect 2440 5940 2560 5950
rect 2690 5940 2810 5950
rect 2940 5940 3060 5950
rect 3190 5940 3310 5950
rect 3440 5940 3560 5950
rect 3690 5940 3810 5950
rect 3940 5940 4060 5950
rect 4190 5940 4310 5950
rect 4440 5940 4560 5950
rect 4690 5940 4810 5950
rect 4940 5940 5060 5950
rect 5190 5940 5310 5950
rect 5440 5940 5560 5950
rect 5690 5940 5810 5950
rect 5940 5940 6060 5950
rect 6190 5940 6310 5950
rect 6440 5940 6560 5950
rect 6690 5940 6810 5950
rect 6940 5940 7060 5950
rect 7190 5940 7310 5950
rect 7440 5940 7560 5950
rect 7690 5940 7810 5950
rect 7940 5940 8000 5950
rect 0 5925 50 5940
rect 0 5825 10 5925
rect 45 5825 50 5925
rect 0 5810 50 5825
rect 200 5925 300 5940
rect 200 5825 205 5925
rect 240 5825 260 5925
rect 295 5825 300 5925
rect 200 5810 300 5825
rect 450 5925 550 5940
rect 450 5825 455 5925
rect 490 5825 510 5925
rect 545 5825 550 5925
rect 450 5810 550 5825
rect 700 5925 800 5940
rect 700 5825 705 5925
rect 740 5825 760 5925
rect 795 5825 800 5925
rect 700 5810 800 5825
rect 950 5925 1050 5940
rect 950 5825 955 5925
rect 990 5825 1010 5925
rect 1045 5825 1050 5925
rect 950 5810 1050 5825
rect 1200 5925 1300 5940
rect 1200 5825 1205 5925
rect 1240 5825 1260 5925
rect 1295 5825 1300 5925
rect 1200 5810 1300 5825
rect 1450 5925 1550 5940
rect 1450 5825 1455 5925
rect 1490 5825 1510 5925
rect 1545 5825 1550 5925
rect 1450 5810 1550 5825
rect 1700 5925 1800 5940
rect 1700 5825 1705 5925
rect 1740 5825 1760 5925
rect 1795 5825 1800 5925
rect 1700 5810 1800 5825
rect 1950 5925 2050 5940
rect 1950 5825 1955 5925
rect 1990 5825 2010 5925
rect 2045 5825 2050 5925
rect 1950 5810 2050 5825
rect 2200 5925 2300 5940
rect 2200 5825 2205 5925
rect 2240 5825 2260 5925
rect 2295 5825 2300 5925
rect 2200 5810 2300 5825
rect 2450 5925 2550 5940
rect 2450 5825 2455 5925
rect 2490 5825 2510 5925
rect 2545 5825 2550 5925
rect 2450 5810 2550 5825
rect 2700 5925 2800 5940
rect 2700 5825 2705 5925
rect 2740 5825 2760 5925
rect 2795 5825 2800 5925
rect 2700 5810 2800 5825
rect 2950 5925 3050 5940
rect 2950 5825 2955 5925
rect 2990 5825 3010 5925
rect 3045 5825 3050 5925
rect 2950 5810 3050 5825
rect 3200 5925 3300 5940
rect 3200 5825 3205 5925
rect 3240 5825 3260 5925
rect 3295 5825 3300 5925
rect 3200 5810 3300 5825
rect 3450 5925 3550 5940
rect 3450 5825 3455 5925
rect 3490 5825 3510 5925
rect 3545 5825 3550 5925
rect 3450 5810 3550 5825
rect 3700 5925 3800 5940
rect 3700 5825 3705 5925
rect 3740 5825 3760 5925
rect 3795 5825 3800 5925
rect 3700 5810 3800 5825
rect 3950 5925 4050 5940
rect 3950 5825 3955 5925
rect 3990 5825 4010 5925
rect 4045 5825 4050 5925
rect 3950 5810 4050 5825
rect 4200 5925 4300 5940
rect 4200 5825 4205 5925
rect 4240 5825 4260 5925
rect 4295 5825 4300 5925
rect 4200 5810 4300 5825
rect 4450 5925 4550 5940
rect 4450 5825 4455 5925
rect 4490 5825 4510 5925
rect 4545 5825 4550 5925
rect 4450 5810 4550 5825
rect 4700 5925 4800 5940
rect 4700 5825 4705 5925
rect 4740 5825 4760 5925
rect 4795 5825 4800 5925
rect 4700 5810 4800 5825
rect 4950 5925 5050 5940
rect 4950 5825 4955 5925
rect 4990 5825 5010 5925
rect 5045 5825 5050 5925
rect 4950 5810 5050 5825
rect 5200 5925 5300 5940
rect 5200 5825 5205 5925
rect 5240 5825 5260 5925
rect 5295 5825 5300 5925
rect 5200 5810 5300 5825
rect 5450 5925 5550 5940
rect 5450 5825 5455 5925
rect 5490 5825 5510 5925
rect 5545 5825 5550 5925
rect 5450 5810 5550 5825
rect 5700 5925 5800 5940
rect 5700 5825 5705 5925
rect 5740 5825 5760 5925
rect 5795 5825 5800 5925
rect 5700 5810 5800 5825
rect 5950 5925 6050 5940
rect 5950 5825 5955 5925
rect 5990 5825 6010 5925
rect 6045 5825 6050 5925
rect 5950 5810 6050 5825
rect 6200 5925 6300 5940
rect 6200 5825 6205 5925
rect 6240 5825 6260 5925
rect 6295 5825 6300 5925
rect 6200 5810 6300 5825
rect 6450 5925 6550 5940
rect 6450 5825 6455 5925
rect 6490 5825 6510 5925
rect 6545 5825 6550 5925
rect 6450 5810 6550 5825
rect 6700 5925 6800 5940
rect 6700 5825 6705 5925
rect 6740 5825 6760 5925
rect 6795 5825 6800 5925
rect 6700 5810 6800 5825
rect 6950 5925 7050 5940
rect 6950 5825 6955 5925
rect 6990 5825 7010 5925
rect 7045 5825 7050 5925
rect 6950 5810 7050 5825
rect 7200 5925 7300 5940
rect 7200 5825 7205 5925
rect 7240 5825 7260 5925
rect 7295 5825 7300 5925
rect 7200 5810 7300 5825
rect 7450 5925 7550 5940
rect 7450 5825 7455 5925
rect 7490 5825 7510 5925
rect 7545 5825 7550 5925
rect 7450 5810 7550 5825
rect 7700 5925 7800 5940
rect 7700 5825 7705 5925
rect 7740 5825 7760 5925
rect 7795 5825 7800 5925
rect 7700 5810 7800 5825
rect 7950 5925 8000 5940
rect 7950 5825 7955 5925
rect 7990 5825 8000 5925
rect 7950 5810 8000 5825
rect 0 5800 60 5810
rect 190 5800 310 5810
rect 440 5800 560 5810
rect 690 5800 810 5810
rect 940 5800 1060 5810
rect 1190 5800 1310 5810
rect 1440 5800 1560 5810
rect 1690 5800 1810 5810
rect 1940 5800 2060 5810
rect 2190 5800 2310 5810
rect 2440 5800 2560 5810
rect 2690 5800 2810 5810
rect 2940 5800 3060 5810
rect 3190 5800 3310 5810
rect 3440 5800 3560 5810
rect 3690 5800 3810 5810
rect 3940 5800 4060 5810
rect 4190 5800 4310 5810
rect 4440 5800 4560 5810
rect 4690 5800 4810 5810
rect 4940 5800 5060 5810
rect 5190 5800 5310 5810
rect 5440 5800 5560 5810
rect 5690 5800 5810 5810
rect 5940 5800 6060 5810
rect 6190 5800 6310 5810
rect 6440 5800 6560 5810
rect 6690 5800 6810 5810
rect 6940 5800 7060 5810
rect 7190 5800 7310 5810
rect 7440 5800 7560 5810
rect 7690 5800 7810 5810
rect 7940 5800 8000 5810
rect 0 5795 8000 5800
rect 0 5760 75 5795
rect 175 5760 325 5795
rect 425 5760 575 5795
rect 675 5760 825 5795
rect 925 5760 1075 5795
rect 1175 5760 1325 5795
rect 1425 5760 1575 5795
rect 1675 5760 1825 5795
rect 1925 5760 2075 5795
rect 2175 5760 2325 5795
rect 2425 5760 2575 5795
rect 2675 5760 2825 5795
rect 2925 5760 3075 5795
rect 3175 5760 3325 5795
rect 3425 5760 3575 5795
rect 3675 5760 3825 5795
rect 3925 5760 4075 5795
rect 4175 5760 4325 5795
rect 4425 5760 4575 5795
rect 4675 5760 4825 5795
rect 4925 5760 5075 5795
rect 5175 5760 5325 5795
rect 5425 5760 5575 5795
rect 5675 5760 5825 5795
rect 5925 5760 6075 5795
rect 6175 5760 6325 5795
rect 6425 5760 6575 5795
rect 6675 5760 6825 5795
rect 6925 5760 7075 5795
rect 7175 5760 7325 5795
rect 7425 5760 7575 5795
rect 7675 5760 7825 5795
rect 7925 5760 8000 5795
rect 0 5740 8000 5760
rect 0 5705 75 5740
rect 175 5705 325 5740
rect 425 5705 575 5740
rect 675 5705 825 5740
rect 925 5705 1075 5740
rect 1175 5705 1325 5740
rect 1425 5705 1575 5740
rect 1675 5705 1825 5740
rect 1925 5705 2075 5740
rect 2175 5705 2325 5740
rect 2425 5705 2575 5740
rect 2675 5705 2825 5740
rect 2925 5705 3075 5740
rect 3175 5705 3325 5740
rect 3425 5705 3575 5740
rect 3675 5705 3825 5740
rect 3925 5705 4075 5740
rect 4175 5705 4325 5740
rect 4425 5705 4575 5740
rect 4675 5705 4825 5740
rect 4925 5705 5075 5740
rect 5175 5705 5325 5740
rect 5425 5705 5575 5740
rect 5675 5705 5825 5740
rect 5925 5705 6075 5740
rect 6175 5705 6325 5740
rect 6425 5705 6575 5740
rect 6675 5705 6825 5740
rect 6925 5705 7075 5740
rect 7175 5705 7325 5740
rect 7425 5705 7575 5740
rect 7675 5705 7825 5740
rect 7925 5705 8000 5740
rect 0 5700 8000 5705
rect 0 5690 60 5700
rect 190 5690 310 5700
rect 440 5690 560 5700
rect 690 5690 810 5700
rect 940 5690 1060 5700
rect 1190 5690 1310 5700
rect 1440 5690 1560 5700
rect 1690 5690 1810 5700
rect 1940 5690 2060 5700
rect 2190 5690 2310 5700
rect 2440 5690 2560 5700
rect 2690 5690 2810 5700
rect 2940 5690 3060 5700
rect 3190 5690 3310 5700
rect 3440 5690 3560 5700
rect 3690 5690 3810 5700
rect 3940 5690 4060 5700
rect 4190 5690 4310 5700
rect 4440 5690 4560 5700
rect 4690 5690 4810 5700
rect 4940 5690 5060 5700
rect 5190 5690 5310 5700
rect 5440 5690 5560 5700
rect 5690 5690 5810 5700
rect 5940 5690 6060 5700
rect 6190 5690 6310 5700
rect 6440 5690 6560 5700
rect 6690 5690 6810 5700
rect 6940 5690 7060 5700
rect 7190 5690 7310 5700
rect 7440 5690 7560 5700
rect 7690 5690 7810 5700
rect 7940 5690 8000 5700
rect 0 5675 50 5690
rect 0 5575 10 5675
rect 45 5575 50 5675
rect 0 5560 50 5575
rect 200 5675 300 5690
rect 200 5575 205 5675
rect 240 5575 260 5675
rect 295 5575 300 5675
rect 200 5560 300 5575
rect 450 5675 550 5690
rect 450 5575 455 5675
rect 490 5575 510 5675
rect 545 5575 550 5675
rect 450 5560 550 5575
rect 700 5675 800 5690
rect 700 5575 705 5675
rect 740 5575 760 5675
rect 795 5575 800 5675
rect 700 5560 800 5575
rect 950 5675 1050 5690
rect 950 5575 955 5675
rect 990 5575 1010 5675
rect 1045 5575 1050 5675
rect 950 5560 1050 5575
rect 1200 5675 1300 5690
rect 1200 5575 1205 5675
rect 1240 5575 1260 5675
rect 1295 5575 1300 5675
rect 1200 5560 1300 5575
rect 1450 5675 1550 5690
rect 1450 5575 1455 5675
rect 1490 5575 1510 5675
rect 1545 5575 1550 5675
rect 1450 5560 1550 5575
rect 1700 5675 1800 5690
rect 1700 5575 1705 5675
rect 1740 5575 1760 5675
rect 1795 5575 1800 5675
rect 1700 5560 1800 5575
rect 1950 5675 2050 5690
rect 1950 5575 1955 5675
rect 1990 5575 2010 5675
rect 2045 5575 2050 5675
rect 1950 5560 2050 5575
rect 2200 5675 2300 5690
rect 2200 5575 2205 5675
rect 2240 5575 2260 5675
rect 2295 5575 2300 5675
rect 2200 5560 2300 5575
rect 2450 5675 2550 5690
rect 2450 5575 2455 5675
rect 2490 5575 2510 5675
rect 2545 5575 2550 5675
rect 2450 5560 2550 5575
rect 2700 5675 2800 5690
rect 2700 5575 2705 5675
rect 2740 5575 2760 5675
rect 2795 5575 2800 5675
rect 2700 5560 2800 5575
rect 2950 5675 3050 5690
rect 2950 5575 2955 5675
rect 2990 5575 3010 5675
rect 3045 5575 3050 5675
rect 2950 5560 3050 5575
rect 3200 5675 3300 5690
rect 3200 5575 3205 5675
rect 3240 5575 3260 5675
rect 3295 5575 3300 5675
rect 3200 5560 3300 5575
rect 3450 5675 3550 5690
rect 3450 5575 3455 5675
rect 3490 5575 3510 5675
rect 3545 5575 3550 5675
rect 3450 5560 3550 5575
rect 3700 5675 3800 5690
rect 3700 5575 3705 5675
rect 3740 5575 3760 5675
rect 3795 5575 3800 5675
rect 3700 5560 3800 5575
rect 3950 5675 4050 5690
rect 3950 5575 3955 5675
rect 3990 5575 4010 5675
rect 4045 5575 4050 5675
rect 3950 5560 4050 5575
rect 4200 5675 4300 5690
rect 4200 5575 4205 5675
rect 4240 5575 4260 5675
rect 4295 5575 4300 5675
rect 4200 5560 4300 5575
rect 4450 5675 4550 5690
rect 4450 5575 4455 5675
rect 4490 5575 4510 5675
rect 4545 5575 4550 5675
rect 4450 5560 4550 5575
rect 4700 5675 4800 5690
rect 4700 5575 4705 5675
rect 4740 5575 4760 5675
rect 4795 5575 4800 5675
rect 4700 5560 4800 5575
rect 4950 5675 5050 5690
rect 4950 5575 4955 5675
rect 4990 5575 5010 5675
rect 5045 5575 5050 5675
rect 4950 5560 5050 5575
rect 5200 5675 5300 5690
rect 5200 5575 5205 5675
rect 5240 5575 5260 5675
rect 5295 5575 5300 5675
rect 5200 5560 5300 5575
rect 5450 5675 5550 5690
rect 5450 5575 5455 5675
rect 5490 5575 5510 5675
rect 5545 5575 5550 5675
rect 5450 5560 5550 5575
rect 5700 5675 5800 5690
rect 5700 5575 5705 5675
rect 5740 5575 5760 5675
rect 5795 5575 5800 5675
rect 5700 5560 5800 5575
rect 5950 5675 6050 5690
rect 5950 5575 5955 5675
rect 5990 5575 6010 5675
rect 6045 5575 6050 5675
rect 5950 5560 6050 5575
rect 6200 5675 6300 5690
rect 6200 5575 6205 5675
rect 6240 5575 6260 5675
rect 6295 5575 6300 5675
rect 6200 5560 6300 5575
rect 6450 5675 6550 5690
rect 6450 5575 6455 5675
rect 6490 5575 6510 5675
rect 6545 5575 6550 5675
rect 6450 5560 6550 5575
rect 6700 5675 6800 5690
rect 6700 5575 6705 5675
rect 6740 5575 6760 5675
rect 6795 5575 6800 5675
rect 6700 5560 6800 5575
rect 6950 5675 7050 5690
rect 6950 5575 6955 5675
rect 6990 5575 7010 5675
rect 7045 5575 7050 5675
rect 6950 5560 7050 5575
rect 7200 5675 7300 5690
rect 7200 5575 7205 5675
rect 7240 5575 7260 5675
rect 7295 5575 7300 5675
rect 7200 5560 7300 5575
rect 7450 5675 7550 5690
rect 7450 5575 7455 5675
rect 7490 5575 7510 5675
rect 7545 5575 7550 5675
rect 7450 5560 7550 5575
rect 7700 5675 7800 5690
rect 7700 5575 7705 5675
rect 7740 5575 7760 5675
rect 7795 5575 7800 5675
rect 7700 5560 7800 5575
rect 7950 5675 8000 5690
rect 7950 5575 7955 5675
rect 7990 5575 8000 5675
rect 7950 5560 8000 5575
rect 0 5550 60 5560
rect 190 5550 310 5560
rect 440 5550 560 5560
rect 690 5550 810 5560
rect 940 5550 1060 5560
rect 1190 5550 1310 5560
rect 1440 5550 1560 5560
rect 1690 5550 1810 5560
rect 1940 5550 2060 5560
rect 2190 5550 2310 5560
rect 2440 5550 2560 5560
rect 2690 5550 2810 5560
rect 2940 5550 3060 5560
rect 3190 5550 3310 5560
rect 3440 5550 3560 5560
rect 3690 5550 3810 5560
rect 3940 5550 4060 5560
rect 4190 5550 4310 5560
rect 4440 5550 4560 5560
rect 4690 5550 4810 5560
rect 4940 5550 5060 5560
rect 5190 5550 5310 5560
rect 5440 5550 5560 5560
rect 5690 5550 5810 5560
rect 5940 5550 6060 5560
rect 6190 5550 6310 5560
rect 6440 5550 6560 5560
rect 6690 5550 6810 5560
rect 6940 5550 7060 5560
rect 7190 5550 7310 5560
rect 7440 5550 7560 5560
rect 7690 5550 7810 5560
rect 7940 5550 8000 5560
rect 0 5545 8000 5550
rect 0 5510 75 5545
rect 175 5510 325 5545
rect 425 5510 575 5545
rect 675 5510 825 5545
rect 925 5510 1075 5545
rect 1175 5510 1325 5545
rect 1425 5510 1575 5545
rect 1675 5510 1825 5545
rect 1925 5510 2075 5545
rect 2175 5510 2325 5545
rect 2425 5510 2575 5545
rect 2675 5510 2825 5545
rect 2925 5510 3075 5545
rect 3175 5510 3325 5545
rect 3425 5510 3575 5545
rect 3675 5510 3825 5545
rect 3925 5510 4075 5545
rect 4175 5510 4325 5545
rect 4425 5510 4575 5545
rect 4675 5510 4825 5545
rect 4925 5510 5075 5545
rect 5175 5510 5325 5545
rect 5425 5510 5575 5545
rect 5675 5510 5825 5545
rect 5925 5510 6075 5545
rect 6175 5510 6325 5545
rect 6425 5510 6575 5545
rect 6675 5510 6825 5545
rect 6925 5510 7075 5545
rect 7175 5510 7325 5545
rect 7425 5510 7575 5545
rect 7675 5510 7825 5545
rect 7925 5510 8000 5545
rect 0 5490 8000 5510
rect 0 5455 75 5490
rect 175 5455 325 5490
rect 425 5455 575 5490
rect 675 5455 825 5490
rect 925 5455 1075 5490
rect 1175 5455 1325 5490
rect 1425 5455 1575 5490
rect 1675 5455 1825 5490
rect 1925 5455 2075 5490
rect 2175 5455 2325 5490
rect 2425 5455 2575 5490
rect 2675 5455 2825 5490
rect 2925 5455 3075 5490
rect 3175 5455 3325 5490
rect 3425 5455 3575 5490
rect 3675 5455 3825 5490
rect 3925 5455 4075 5490
rect 4175 5455 4325 5490
rect 4425 5455 4575 5490
rect 4675 5455 4825 5490
rect 4925 5455 5075 5490
rect 5175 5455 5325 5490
rect 5425 5455 5575 5490
rect 5675 5455 5825 5490
rect 5925 5455 6075 5490
rect 6175 5455 6325 5490
rect 6425 5455 6575 5490
rect 6675 5455 6825 5490
rect 6925 5455 7075 5490
rect 7175 5455 7325 5490
rect 7425 5455 7575 5490
rect 7675 5455 7825 5490
rect 7925 5455 8000 5490
rect 0 5450 8000 5455
rect 0 5440 60 5450
rect 190 5440 310 5450
rect 440 5440 560 5450
rect 690 5440 810 5450
rect 940 5440 1060 5450
rect 1190 5440 1310 5450
rect 1440 5440 1560 5450
rect 1690 5440 1810 5450
rect 1940 5440 2060 5450
rect 2190 5440 2310 5450
rect 2440 5440 2560 5450
rect 2690 5440 2810 5450
rect 2940 5440 3060 5450
rect 3190 5440 3310 5450
rect 3440 5440 3560 5450
rect 3690 5440 3810 5450
rect 3940 5440 4060 5450
rect 4190 5440 4310 5450
rect 4440 5440 4560 5450
rect 4690 5440 4810 5450
rect 4940 5440 5060 5450
rect 5190 5440 5310 5450
rect 5440 5440 5560 5450
rect 5690 5440 5810 5450
rect 5940 5440 6060 5450
rect 6190 5440 6310 5450
rect 6440 5440 6560 5450
rect 6690 5440 6810 5450
rect 6940 5440 7060 5450
rect 7190 5440 7310 5450
rect 7440 5440 7560 5450
rect 7690 5440 7810 5450
rect 7940 5440 8000 5450
rect 0 5425 50 5440
rect 0 5325 10 5425
rect 45 5325 50 5425
rect 0 5310 50 5325
rect 200 5425 300 5440
rect 200 5325 205 5425
rect 240 5325 260 5425
rect 295 5325 300 5425
rect 200 5310 300 5325
rect 450 5425 550 5440
rect 450 5325 455 5425
rect 490 5325 510 5425
rect 545 5325 550 5425
rect 450 5310 550 5325
rect 700 5425 800 5440
rect 700 5325 705 5425
rect 740 5325 760 5425
rect 795 5325 800 5425
rect 700 5310 800 5325
rect 950 5425 1050 5440
rect 950 5325 955 5425
rect 990 5325 1010 5425
rect 1045 5325 1050 5425
rect 950 5310 1050 5325
rect 1200 5425 1300 5440
rect 1200 5325 1205 5425
rect 1240 5325 1260 5425
rect 1295 5325 1300 5425
rect 1200 5310 1300 5325
rect 1450 5425 1550 5440
rect 1450 5325 1455 5425
rect 1490 5325 1510 5425
rect 1545 5325 1550 5425
rect 1450 5310 1550 5325
rect 1700 5425 1800 5440
rect 1700 5325 1705 5425
rect 1740 5325 1760 5425
rect 1795 5325 1800 5425
rect 1700 5310 1800 5325
rect 1950 5425 2050 5440
rect 1950 5325 1955 5425
rect 1990 5325 2010 5425
rect 2045 5325 2050 5425
rect 1950 5310 2050 5325
rect 2200 5425 2300 5440
rect 2200 5325 2205 5425
rect 2240 5325 2260 5425
rect 2295 5325 2300 5425
rect 2200 5310 2300 5325
rect 2450 5425 2550 5440
rect 2450 5325 2455 5425
rect 2490 5325 2510 5425
rect 2545 5325 2550 5425
rect 2450 5310 2550 5325
rect 2700 5425 2800 5440
rect 2700 5325 2705 5425
rect 2740 5325 2760 5425
rect 2795 5325 2800 5425
rect 2700 5310 2800 5325
rect 2950 5425 3050 5440
rect 2950 5325 2955 5425
rect 2990 5325 3010 5425
rect 3045 5325 3050 5425
rect 2950 5310 3050 5325
rect 3200 5425 3300 5440
rect 3200 5325 3205 5425
rect 3240 5325 3260 5425
rect 3295 5325 3300 5425
rect 3200 5310 3300 5325
rect 3450 5425 3550 5440
rect 3450 5325 3455 5425
rect 3490 5325 3510 5425
rect 3545 5325 3550 5425
rect 3450 5310 3550 5325
rect 3700 5425 3800 5440
rect 3700 5325 3705 5425
rect 3740 5325 3760 5425
rect 3795 5325 3800 5425
rect 3700 5310 3800 5325
rect 3950 5425 4050 5440
rect 3950 5325 3955 5425
rect 3990 5325 4010 5425
rect 4045 5325 4050 5425
rect 3950 5310 4050 5325
rect 4200 5425 4300 5440
rect 4200 5325 4205 5425
rect 4240 5325 4260 5425
rect 4295 5325 4300 5425
rect 4200 5310 4300 5325
rect 4450 5425 4550 5440
rect 4450 5325 4455 5425
rect 4490 5325 4510 5425
rect 4545 5325 4550 5425
rect 4450 5310 4550 5325
rect 4700 5425 4800 5440
rect 4700 5325 4705 5425
rect 4740 5325 4760 5425
rect 4795 5325 4800 5425
rect 4700 5310 4800 5325
rect 4950 5425 5050 5440
rect 4950 5325 4955 5425
rect 4990 5325 5010 5425
rect 5045 5325 5050 5425
rect 4950 5310 5050 5325
rect 5200 5425 5300 5440
rect 5200 5325 5205 5425
rect 5240 5325 5260 5425
rect 5295 5325 5300 5425
rect 5200 5310 5300 5325
rect 5450 5425 5550 5440
rect 5450 5325 5455 5425
rect 5490 5325 5510 5425
rect 5545 5325 5550 5425
rect 5450 5310 5550 5325
rect 5700 5425 5800 5440
rect 5700 5325 5705 5425
rect 5740 5325 5760 5425
rect 5795 5325 5800 5425
rect 5700 5310 5800 5325
rect 5950 5425 6050 5440
rect 5950 5325 5955 5425
rect 5990 5325 6010 5425
rect 6045 5325 6050 5425
rect 5950 5310 6050 5325
rect 6200 5425 6300 5440
rect 6200 5325 6205 5425
rect 6240 5325 6260 5425
rect 6295 5325 6300 5425
rect 6200 5310 6300 5325
rect 6450 5425 6550 5440
rect 6450 5325 6455 5425
rect 6490 5325 6510 5425
rect 6545 5325 6550 5425
rect 6450 5310 6550 5325
rect 6700 5425 6800 5440
rect 6700 5325 6705 5425
rect 6740 5325 6760 5425
rect 6795 5325 6800 5425
rect 6700 5310 6800 5325
rect 6950 5425 7050 5440
rect 6950 5325 6955 5425
rect 6990 5325 7010 5425
rect 7045 5325 7050 5425
rect 6950 5310 7050 5325
rect 7200 5425 7300 5440
rect 7200 5325 7205 5425
rect 7240 5325 7260 5425
rect 7295 5325 7300 5425
rect 7200 5310 7300 5325
rect 7450 5425 7550 5440
rect 7450 5325 7455 5425
rect 7490 5325 7510 5425
rect 7545 5325 7550 5425
rect 7450 5310 7550 5325
rect 7700 5425 7800 5440
rect 7700 5325 7705 5425
rect 7740 5325 7760 5425
rect 7795 5325 7800 5425
rect 7700 5310 7800 5325
rect 7950 5425 8000 5440
rect 7950 5325 7955 5425
rect 7990 5325 8000 5425
rect 7950 5310 8000 5325
rect 0 5300 60 5310
rect 190 5300 310 5310
rect 440 5300 560 5310
rect 690 5300 810 5310
rect 940 5300 1060 5310
rect 1190 5300 1310 5310
rect 1440 5300 1560 5310
rect 1690 5300 1810 5310
rect 1940 5300 2060 5310
rect 2190 5300 2310 5310
rect 2440 5300 2560 5310
rect 2690 5300 2810 5310
rect 2940 5300 3060 5310
rect 3190 5300 3310 5310
rect 3440 5300 3560 5310
rect 3690 5300 3810 5310
rect 3940 5300 4060 5310
rect 4190 5300 4310 5310
rect 4440 5300 4560 5310
rect 4690 5300 4810 5310
rect 4940 5300 5060 5310
rect 5190 5300 5310 5310
rect 5440 5300 5560 5310
rect 5690 5300 5810 5310
rect 5940 5300 6060 5310
rect 6190 5300 6310 5310
rect 6440 5300 6560 5310
rect 6690 5300 6810 5310
rect 6940 5300 7060 5310
rect 7190 5300 7310 5310
rect 7440 5300 7560 5310
rect 7690 5300 7810 5310
rect 7940 5300 8000 5310
rect 0 5295 8000 5300
rect 0 5260 75 5295
rect 175 5260 325 5295
rect 425 5260 575 5295
rect 675 5260 825 5295
rect 925 5260 1075 5295
rect 1175 5260 1325 5295
rect 1425 5260 1575 5295
rect 1675 5260 1825 5295
rect 1925 5260 2075 5295
rect 2175 5260 2325 5295
rect 2425 5260 2575 5295
rect 2675 5260 2825 5295
rect 2925 5260 3075 5295
rect 3175 5260 3325 5295
rect 3425 5260 3575 5295
rect 3675 5260 3825 5295
rect 3925 5260 4075 5295
rect 4175 5260 4325 5295
rect 4425 5260 4575 5295
rect 4675 5260 4825 5295
rect 4925 5260 5075 5295
rect 5175 5260 5325 5295
rect 5425 5260 5575 5295
rect 5675 5260 5825 5295
rect 5925 5260 6075 5295
rect 6175 5260 6325 5295
rect 6425 5260 6575 5295
rect 6675 5260 6825 5295
rect 6925 5260 7075 5295
rect 7175 5260 7325 5295
rect 7425 5260 7575 5295
rect 7675 5260 7825 5295
rect 7925 5260 8000 5295
rect 0 5240 8000 5260
rect 0 5205 75 5240
rect 175 5205 325 5240
rect 425 5205 575 5240
rect 675 5205 825 5240
rect 925 5205 1075 5240
rect 1175 5205 1325 5240
rect 1425 5205 1575 5240
rect 1675 5205 1825 5240
rect 1925 5205 2075 5240
rect 2175 5205 2325 5240
rect 2425 5205 2575 5240
rect 2675 5205 2825 5240
rect 2925 5205 3075 5240
rect 3175 5205 3325 5240
rect 3425 5205 3575 5240
rect 3675 5205 3825 5240
rect 3925 5205 4075 5240
rect 4175 5205 4325 5240
rect 4425 5205 4575 5240
rect 4675 5205 4825 5240
rect 4925 5205 5075 5240
rect 5175 5205 5325 5240
rect 5425 5205 5575 5240
rect 5675 5205 5825 5240
rect 5925 5205 6075 5240
rect 6175 5205 6325 5240
rect 6425 5205 6575 5240
rect 6675 5205 6825 5240
rect 6925 5205 7075 5240
rect 7175 5205 7325 5240
rect 7425 5205 7575 5240
rect 7675 5205 7825 5240
rect 7925 5205 8000 5240
rect 0 5200 8000 5205
rect 0 5190 60 5200
rect 190 5190 310 5200
rect 440 5190 560 5200
rect 690 5190 810 5200
rect 940 5190 1060 5200
rect 1190 5190 1310 5200
rect 1440 5190 1560 5200
rect 1690 5190 1810 5200
rect 1940 5190 2060 5200
rect 2190 5190 2310 5200
rect 2440 5190 2560 5200
rect 2690 5190 2810 5200
rect 2940 5190 3060 5200
rect 3190 5190 3310 5200
rect 3440 5190 3560 5200
rect 3690 5190 3810 5200
rect 3940 5190 4060 5200
rect 4190 5190 4310 5200
rect 4440 5190 4560 5200
rect 4690 5190 4810 5200
rect 4940 5190 5060 5200
rect 5190 5190 5310 5200
rect 5440 5190 5560 5200
rect 5690 5190 5810 5200
rect 5940 5190 6060 5200
rect 6190 5190 6310 5200
rect 6440 5190 6560 5200
rect 6690 5190 6810 5200
rect 6940 5190 7060 5200
rect 7190 5190 7310 5200
rect 7440 5190 7560 5200
rect 7690 5190 7810 5200
rect 7940 5190 8000 5200
rect 0 5175 50 5190
rect 0 5075 10 5175
rect 45 5075 50 5175
rect 0 5060 50 5075
rect 200 5175 300 5190
rect 200 5075 205 5175
rect 240 5075 260 5175
rect 295 5075 300 5175
rect 200 5060 300 5075
rect 450 5175 550 5190
rect 450 5075 455 5175
rect 490 5075 510 5175
rect 545 5075 550 5175
rect 450 5060 550 5075
rect 700 5175 800 5190
rect 700 5075 705 5175
rect 740 5075 760 5175
rect 795 5075 800 5175
rect 700 5060 800 5075
rect 950 5175 1050 5190
rect 950 5075 955 5175
rect 990 5075 1010 5175
rect 1045 5075 1050 5175
rect 950 5060 1050 5075
rect 1200 5175 1300 5190
rect 1200 5075 1205 5175
rect 1240 5075 1260 5175
rect 1295 5075 1300 5175
rect 1200 5060 1300 5075
rect 1450 5175 1550 5190
rect 1450 5075 1455 5175
rect 1490 5075 1510 5175
rect 1545 5075 1550 5175
rect 1450 5060 1550 5075
rect 1700 5175 1800 5190
rect 1700 5075 1705 5175
rect 1740 5075 1760 5175
rect 1795 5075 1800 5175
rect 1700 5060 1800 5075
rect 1950 5175 2050 5190
rect 1950 5075 1955 5175
rect 1990 5075 2010 5175
rect 2045 5075 2050 5175
rect 1950 5060 2050 5075
rect 2200 5175 2300 5190
rect 2200 5075 2205 5175
rect 2240 5075 2260 5175
rect 2295 5075 2300 5175
rect 2200 5060 2300 5075
rect 2450 5175 2550 5190
rect 2450 5075 2455 5175
rect 2490 5075 2510 5175
rect 2545 5075 2550 5175
rect 2450 5060 2550 5075
rect 2700 5175 2800 5190
rect 2700 5075 2705 5175
rect 2740 5075 2760 5175
rect 2795 5075 2800 5175
rect 2700 5060 2800 5075
rect 2950 5175 3050 5190
rect 2950 5075 2955 5175
rect 2990 5075 3010 5175
rect 3045 5075 3050 5175
rect 2950 5060 3050 5075
rect 3200 5175 3300 5190
rect 3200 5075 3205 5175
rect 3240 5075 3260 5175
rect 3295 5075 3300 5175
rect 3200 5060 3300 5075
rect 3450 5175 3550 5190
rect 3450 5075 3455 5175
rect 3490 5075 3510 5175
rect 3545 5075 3550 5175
rect 3450 5060 3550 5075
rect 3700 5175 3800 5190
rect 3700 5075 3705 5175
rect 3740 5075 3760 5175
rect 3795 5075 3800 5175
rect 3700 5060 3800 5075
rect 3950 5175 4050 5190
rect 3950 5075 3955 5175
rect 3990 5075 4010 5175
rect 4045 5075 4050 5175
rect 3950 5060 4050 5075
rect 4200 5175 4300 5190
rect 4200 5075 4205 5175
rect 4240 5075 4260 5175
rect 4295 5075 4300 5175
rect 4200 5060 4300 5075
rect 4450 5175 4550 5190
rect 4450 5075 4455 5175
rect 4490 5075 4510 5175
rect 4545 5075 4550 5175
rect 4450 5060 4550 5075
rect 4700 5175 4800 5190
rect 4700 5075 4705 5175
rect 4740 5075 4760 5175
rect 4795 5075 4800 5175
rect 4700 5060 4800 5075
rect 4950 5175 5050 5190
rect 4950 5075 4955 5175
rect 4990 5075 5010 5175
rect 5045 5075 5050 5175
rect 4950 5060 5050 5075
rect 5200 5175 5300 5190
rect 5200 5075 5205 5175
rect 5240 5075 5260 5175
rect 5295 5075 5300 5175
rect 5200 5060 5300 5075
rect 5450 5175 5550 5190
rect 5450 5075 5455 5175
rect 5490 5075 5510 5175
rect 5545 5075 5550 5175
rect 5450 5060 5550 5075
rect 5700 5175 5800 5190
rect 5700 5075 5705 5175
rect 5740 5075 5760 5175
rect 5795 5075 5800 5175
rect 5700 5060 5800 5075
rect 5950 5175 6050 5190
rect 5950 5075 5955 5175
rect 5990 5075 6010 5175
rect 6045 5075 6050 5175
rect 5950 5060 6050 5075
rect 6200 5175 6300 5190
rect 6200 5075 6205 5175
rect 6240 5075 6260 5175
rect 6295 5075 6300 5175
rect 6200 5060 6300 5075
rect 6450 5175 6550 5190
rect 6450 5075 6455 5175
rect 6490 5075 6510 5175
rect 6545 5075 6550 5175
rect 6450 5060 6550 5075
rect 6700 5175 6800 5190
rect 6700 5075 6705 5175
rect 6740 5075 6760 5175
rect 6795 5075 6800 5175
rect 6700 5060 6800 5075
rect 6950 5175 7050 5190
rect 6950 5075 6955 5175
rect 6990 5075 7010 5175
rect 7045 5075 7050 5175
rect 6950 5060 7050 5075
rect 7200 5175 7300 5190
rect 7200 5075 7205 5175
rect 7240 5075 7260 5175
rect 7295 5075 7300 5175
rect 7200 5060 7300 5075
rect 7450 5175 7550 5190
rect 7450 5075 7455 5175
rect 7490 5075 7510 5175
rect 7545 5075 7550 5175
rect 7450 5060 7550 5075
rect 7700 5175 7800 5190
rect 7700 5075 7705 5175
rect 7740 5075 7760 5175
rect 7795 5075 7800 5175
rect 7700 5060 7800 5075
rect 7950 5175 8000 5190
rect 7950 5075 7955 5175
rect 7990 5075 8000 5175
rect 7950 5060 8000 5075
rect 0 5050 60 5060
rect 190 5050 310 5060
rect 440 5050 560 5060
rect 690 5050 810 5060
rect 940 5050 1060 5060
rect 1190 5050 1310 5060
rect 1440 5050 1560 5060
rect 1690 5050 1810 5060
rect 1940 5050 2060 5060
rect 2190 5050 2310 5060
rect 2440 5050 2560 5060
rect 2690 5050 2810 5060
rect 2940 5050 3060 5060
rect 3190 5050 3310 5060
rect 3440 5050 3560 5060
rect 3690 5050 3810 5060
rect 3940 5050 4060 5060
rect 4190 5050 4310 5060
rect 4440 5050 4560 5060
rect 4690 5050 4810 5060
rect 4940 5050 5060 5060
rect 5190 5050 5310 5060
rect 5440 5050 5560 5060
rect 5690 5050 5810 5060
rect 5940 5050 6060 5060
rect 6190 5050 6310 5060
rect 6440 5050 6560 5060
rect 6690 5050 6810 5060
rect 6940 5050 7060 5060
rect 7190 5050 7310 5060
rect 7440 5050 7560 5060
rect 7690 5050 7810 5060
rect 7940 5050 8000 5060
rect 0 5045 8000 5050
rect 0 5010 75 5045
rect 175 5010 325 5045
rect 425 5010 575 5045
rect 675 5010 825 5045
rect 925 5010 1075 5045
rect 1175 5010 1325 5045
rect 1425 5010 1575 5045
rect 1675 5010 1825 5045
rect 1925 5010 2075 5045
rect 2175 5010 2325 5045
rect 2425 5010 2575 5045
rect 2675 5010 2825 5045
rect 2925 5010 3075 5045
rect 3175 5010 3325 5045
rect 3425 5010 3575 5045
rect 3675 5010 3825 5045
rect 3925 5010 4075 5045
rect 4175 5010 4325 5045
rect 4425 5010 4575 5045
rect 4675 5010 4825 5045
rect 4925 5010 5075 5045
rect 5175 5010 5325 5045
rect 5425 5010 5575 5045
rect 5675 5010 5825 5045
rect 5925 5010 6075 5045
rect 6175 5010 6325 5045
rect 6425 5010 6575 5045
rect 6675 5010 6825 5045
rect 6925 5010 7075 5045
rect 7175 5010 7325 5045
rect 7425 5010 7575 5045
rect 7675 5010 7825 5045
rect 7925 5010 8000 5045
rect 0 4990 8000 5010
rect 0 4955 75 4990
rect 175 4955 325 4990
rect 425 4955 575 4990
rect 675 4955 825 4990
rect 925 4955 1075 4990
rect 1175 4955 1325 4990
rect 1425 4955 1575 4990
rect 1675 4955 1825 4990
rect 1925 4955 2075 4990
rect 2175 4955 2325 4990
rect 2425 4955 2575 4990
rect 2675 4955 2825 4990
rect 2925 4955 3075 4990
rect 3175 4955 3325 4990
rect 3425 4955 3575 4990
rect 3675 4955 3825 4990
rect 3925 4955 4075 4990
rect 4175 4955 4325 4990
rect 4425 4955 4575 4990
rect 4675 4955 4825 4990
rect 4925 4955 5075 4990
rect 5175 4955 5325 4990
rect 5425 4955 5575 4990
rect 5675 4955 5825 4990
rect 5925 4955 6075 4990
rect 6175 4955 6325 4990
rect 6425 4955 6575 4990
rect 6675 4955 6825 4990
rect 6925 4955 7075 4990
rect 7175 4955 7325 4990
rect 7425 4955 7575 4990
rect 7675 4955 7825 4990
rect 7925 4955 8000 4990
rect 0 4950 8000 4955
rect 0 4940 60 4950
rect 190 4940 310 4950
rect 440 4940 560 4950
rect 690 4940 810 4950
rect 940 4940 1060 4950
rect 1190 4940 1310 4950
rect 1440 4940 1560 4950
rect 1690 4940 1810 4950
rect 1940 4940 2060 4950
rect 2190 4940 2310 4950
rect 2440 4940 2560 4950
rect 2690 4940 2810 4950
rect 2940 4940 3060 4950
rect 3190 4940 3310 4950
rect 3440 4940 3560 4950
rect 3690 4940 3810 4950
rect 3940 4940 4060 4950
rect 4190 4940 4310 4950
rect 4440 4940 4560 4950
rect 4690 4940 4810 4950
rect 4940 4940 5060 4950
rect 5190 4940 5310 4950
rect 5440 4940 5560 4950
rect 5690 4940 5810 4950
rect 5940 4940 6060 4950
rect 6190 4940 6310 4950
rect 6440 4940 6560 4950
rect 6690 4940 6810 4950
rect 6940 4940 7060 4950
rect 7190 4940 7310 4950
rect 7440 4940 7560 4950
rect 7690 4940 7810 4950
rect 7940 4940 8000 4950
rect 0 4925 50 4940
rect 0 4825 10 4925
rect 45 4825 50 4925
rect 0 4810 50 4825
rect 200 4925 300 4940
rect 200 4825 205 4925
rect 240 4825 260 4925
rect 295 4825 300 4925
rect 200 4810 300 4825
rect 450 4925 550 4940
rect 450 4825 455 4925
rect 490 4825 510 4925
rect 545 4825 550 4925
rect 450 4810 550 4825
rect 700 4925 800 4940
rect 700 4825 705 4925
rect 740 4825 760 4925
rect 795 4825 800 4925
rect 700 4810 800 4825
rect 950 4925 1050 4940
rect 950 4825 955 4925
rect 990 4825 1010 4925
rect 1045 4825 1050 4925
rect 950 4810 1050 4825
rect 1200 4925 1300 4940
rect 1200 4825 1205 4925
rect 1240 4825 1260 4925
rect 1295 4825 1300 4925
rect 1200 4810 1300 4825
rect 1450 4925 1550 4940
rect 1450 4825 1455 4925
rect 1490 4825 1510 4925
rect 1545 4825 1550 4925
rect 1450 4810 1550 4825
rect 1700 4925 1800 4940
rect 1700 4825 1705 4925
rect 1740 4825 1760 4925
rect 1795 4825 1800 4925
rect 1700 4810 1800 4825
rect 1950 4925 2050 4940
rect 1950 4825 1955 4925
rect 1990 4825 2010 4925
rect 2045 4825 2050 4925
rect 1950 4810 2050 4825
rect 2200 4925 2300 4940
rect 2200 4825 2205 4925
rect 2240 4825 2260 4925
rect 2295 4825 2300 4925
rect 2200 4810 2300 4825
rect 2450 4925 2550 4940
rect 2450 4825 2455 4925
rect 2490 4825 2510 4925
rect 2545 4825 2550 4925
rect 2450 4810 2550 4825
rect 2700 4925 2800 4940
rect 2700 4825 2705 4925
rect 2740 4825 2760 4925
rect 2795 4825 2800 4925
rect 2700 4810 2800 4825
rect 2950 4925 3050 4940
rect 2950 4825 2955 4925
rect 2990 4825 3010 4925
rect 3045 4825 3050 4925
rect 2950 4810 3050 4825
rect 3200 4925 3300 4940
rect 3200 4825 3205 4925
rect 3240 4825 3260 4925
rect 3295 4825 3300 4925
rect 3200 4810 3300 4825
rect 3450 4925 3550 4940
rect 3450 4825 3455 4925
rect 3490 4825 3510 4925
rect 3545 4825 3550 4925
rect 3450 4810 3550 4825
rect 3700 4925 3800 4940
rect 3700 4825 3705 4925
rect 3740 4825 3760 4925
rect 3795 4825 3800 4925
rect 3700 4810 3800 4825
rect 3950 4925 4050 4940
rect 3950 4825 3955 4925
rect 3990 4825 4010 4925
rect 4045 4825 4050 4925
rect 3950 4810 4050 4825
rect 4200 4925 4300 4940
rect 4200 4825 4205 4925
rect 4240 4825 4260 4925
rect 4295 4825 4300 4925
rect 4200 4810 4300 4825
rect 4450 4925 4550 4940
rect 4450 4825 4455 4925
rect 4490 4825 4510 4925
rect 4545 4825 4550 4925
rect 4450 4810 4550 4825
rect 4700 4925 4800 4940
rect 4700 4825 4705 4925
rect 4740 4825 4760 4925
rect 4795 4825 4800 4925
rect 4700 4810 4800 4825
rect 4950 4925 5050 4940
rect 4950 4825 4955 4925
rect 4990 4825 5010 4925
rect 5045 4825 5050 4925
rect 4950 4810 5050 4825
rect 5200 4925 5300 4940
rect 5200 4825 5205 4925
rect 5240 4825 5260 4925
rect 5295 4825 5300 4925
rect 5200 4810 5300 4825
rect 5450 4925 5550 4940
rect 5450 4825 5455 4925
rect 5490 4825 5510 4925
rect 5545 4825 5550 4925
rect 5450 4810 5550 4825
rect 5700 4925 5800 4940
rect 5700 4825 5705 4925
rect 5740 4825 5760 4925
rect 5795 4825 5800 4925
rect 5700 4810 5800 4825
rect 5950 4925 6050 4940
rect 5950 4825 5955 4925
rect 5990 4825 6010 4925
rect 6045 4825 6050 4925
rect 5950 4810 6050 4825
rect 6200 4925 6300 4940
rect 6200 4825 6205 4925
rect 6240 4825 6260 4925
rect 6295 4825 6300 4925
rect 6200 4810 6300 4825
rect 6450 4925 6550 4940
rect 6450 4825 6455 4925
rect 6490 4825 6510 4925
rect 6545 4825 6550 4925
rect 6450 4810 6550 4825
rect 6700 4925 6800 4940
rect 6700 4825 6705 4925
rect 6740 4825 6760 4925
rect 6795 4825 6800 4925
rect 6700 4810 6800 4825
rect 6950 4925 7050 4940
rect 6950 4825 6955 4925
rect 6990 4825 7010 4925
rect 7045 4825 7050 4925
rect 6950 4810 7050 4825
rect 7200 4925 7300 4940
rect 7200 4825 7205 4925
rect 7240 4825 7260 4925
rect 7295 4825 7300 4925
rect 7200 4810 7300 4825
rect 7450 4925 7550 4940
rect 7450 4825 7455 4925
rect 7490 4825 7510 4925
rect 7545 4825 7550 4925
rect 7450 4810 7550 4825
rect 7700 4925 7800 4940
rect 7700 4825 7705 4925
rect 7740 4825 7760 4925
rect 7795 4825 7800 4925
rect 7700 4810 7800 4825
rect 7950 4925 8000 4940
rect 7950 4825 7955 4925
rect 7990 4825 8000 4925
rect 7950 4810 8000 4825
rect 0 4800 60 4810
rect 190 4800 310 4810
rect 440 4800 560 4810
rect 690 4800 810 4810
rect 940 4800 1060 4810
rect 1190 4800 1310 4810
rect 1440 4800 1560 4810
rect 1690 4800 1810 4810
rect 1940 4800 2060 4810
rect 2190 4800 2310 4810
rect 2440 4800 2560 4810
rect 2690 4800 2810 4810
rect 2940 4800 3060 4810
rect 3190 4800 3310 4810
rect 3440 4800 3560 4810
rect 3690 4800 3810 4810
rect 3940 4800 4060 4810
rect 4190 4800 4310 4810
rect 4440 4800 4560 4810
rect 4690 4800 4810 4810
rect 4940 4800 5060 4810
rect 5190 4800 5310 4810
rect 5440 4800 5560 4810
rect 5690 4800 5810 4810
rect 5940 4800 6060 4810
rect 6190 4800 6310 4810
rect 6440 4800 6560 4810
rect 6690 4800 6810 4810
rect 6940 4800 7060 4810
rect 7190 4800 7310 4810
rect 7440 4800 7560 4810
rect 7690 4800 7810 4810
rect 7940 4800 8000 4810
rect 0 4795 8000 4800
rect 0 4760 75 4795
rect 175 4760 325 4795
rect 425 4760 575 4795
rect 675 4760 825 4795
rect 925 4760 1075 4795
rect 1175 4760 1325 4795
rect 1425 4760 1575 4795
rect 1675 4760 1825 4795
rect 1925 4760 2075 4795
rect 2175 4760 2325 4795
rect 2425 4760 2575 4795
rect 2675 4760 2825 4795
rect 2925 4760 3075 4795
rect 3175 4760 3325 4795
rect 3425 4760 3575 4795
rect 3675 4760 3825 4795
rect 3925 4760 4075 4795
rect 4175 4760 4325 4795
rect 4425 4760 4575 4795
rect 4675 4760 4825 4795
rect 4925 4760 5075 4795
rect 5175 4760 5325 4795
rect 5425 4760 5575 4795
rect 5675 4760 5825 4795
rect 5925 4760 6075 4795
rect 6175 4760 6325 4795
rect 6425 4760 6575 4795
rect 6675 4760 6825 4795
rect 6925 4760 7075 4795
rect 7175 4760 7325 4795
rect 7425 4760 7575 4795
rect 7675 4760 7825 4795
rect 7925 4760 8000 4795
rect 0 4740 8000 4760
rect 0 4705 75 4740
rect 175 4705 325 4740
rect 425 4705 575 4740
rect 675 4705 825 4740
rect 925 4705 1075 4740
rect 1175 4705 1325 4740
rect 1425 4705 1575 4740
rect 1675 4705 1825 4740
rect 1925 4705 2075 4740
rect 2175 4705 2325 4740
rect 2425 4705 2575 4740
rect 2675 4705 2825 4740
rect 2925 4705 3075 4740
rect 3175 4705 3325 4740
rect 3425 4705 3575 4740
rect 3675 4705 3825 4740
rect 3925 4705 4075 4740
rect 4175 4705 4325 4740
rect 4425 4705 4575 4740
rect 4675 4705 4825 4740
rect 4925 4705 5075 4740
rect 5175 4705 5325 4740
rect 5425 4705 5575 4740
rect 5675 4705 5825 4740
rect 5925 4705 6075 4740
rect 6175 4705 6325 4740
rect 6425 4705 6575 4740
rect 6675 4705 6825 4740
rect 6925 4705 7075 4740
rect 7175 4705 7325 4740
rect 7425 4705 7575 4740
rect 7675 4705 7825 4740
rect 7925 4705 8000 4740
rect 0 4700 8000 4705
rect 0 4690 60 4700
rect 190 4690 310 4700
rect 440 4690 560 4700
rect 690 4690 810 4700
rect 940 4690 1060 4700
rect 1190 4690 1310 4700
rect 1440 4690 1560 4700
rect 1690 4690 1810 4700
rect 1940 4690 2060 4700
rect 2190 4690 2310 4700
rect 2440 4690 2560 4700
rect 2690 4690 2810 4700
rect 2940 4690 3060 4700
rect 3190 4690 3310 4700
rect 3440 4690 3560 4700
rect 3690 4690 3810 4700
rect 3940 4690 4060 4700
rect 4190 4690 4310 4700
rect 4440 4690 4560 4700
rect 4690 4690 4810 4700
rect 4940 4690 5060 4700
rect 5190 4690 5310 4700
rect 5440 4690 5560 4700
rect 5690 4690 5810 4700
rect 5940 4690 6060 4700
rect 6190 4690 6310 4700
rect 6440 4690 6560 4700
rect 6690 4690 6810 4700
rect 6940 4690 7060 4700
rect 7190 4690 7310 4700
rect 7440 4690 7560 4700
rect 7690 4690 7810 4700
rect 7940 4690 8000 4700
rect 0 4675 50 4690
rect 0 4575 10 4675
rect 45 4575 50 4675
rect 0 4560 50 4575
rect 200 4675 300 4690
rect 200 4575 205 4675
rect 240 4575 260 4675
rect 295 4575 300 4675
rect 200 4560 300 4575
rect 450 4675 550 4690
rect 450 4575 455 4675
rect 490 4575 510 4675
rect 545 4575 550 4675
rect 450 4560 550 4575
rect 700 4675 800 4690
rect 700 4575 705 4675
rect 740 4575 760 4675
rect 795 4575 800 4675
rect 700 4560 800 4575
rect 950 4675 1050 4690
rect 950 4575 955 4675
rect 990 4575 1010 4675
rect 1045 4575 1050 4675
rect 950 4560 1050 4575
rect 1200 4675 1300 4690
rect 1200 4575 1205 4675
rect 1240 4575 1260 4675
rect 1295 4575 1300 4675
rect 1200 4560 1300 4575
rect 1450 4675 1550 4690
rect 1450 4575 1455 4675
rect 1490 4575 1510 4675
rect 1545 4575 1550 4675
rect 1450 4560 1550 4575
rect 1700 4675 1800 4690
rect 1700 4575 1705 4675
rect 1740 4575 1760 4675
rect 1795 4575 1800 4675
rect 1700 4560 1800 4575
rect 1950 4675 2050 4690
rect 1950 4575 1955 4675
rect 1990 4575 2010 4675
rect 2045 4575 2050 4675
rect 1950 4560 2050 4575
rect 2200 4675 2300 4690
rect 2200 4575 2205 4675
rect 2240 4575 2260 4675
rect 2295 4575 2300 4675
rect 2200 4560 2300 4575
rect 2450 4675 2550 4690
rect 2450 4575 2455 4675
rect 2490 4575 2510 4675
rect 2545 4575 2550 4675
rect 2450 4560 2550 4575
rect 2700 4675 2800 4690
rect 2700 4575 2705 4675
rect 2740 4575 2760 4675
rect 2795 4575 2800 4675
rect 2700 4560 2800 4575
rect 2950 4675 3050 4690
rect 2950 4575 2955 4675
rect 2990 4575 3010 4675
rect 3045 4575 3050 4675
rect 2950 4560 3050 4575
rect 3200 4675 3300 4690
rect 3200 4575 3205 4675
rect 3240 4575 3260 4675
rect 3295 4575 3300 4675
rect 3200 4560 3300 4575
rect 3450 4675 3550 4690
rect 3450 4575 3455 4675
rect 3490 4575 3510 4675
rect 3545 4575 3550 4675
rect 3450 4560 3550 4575
rect 3700 4675 3800 4690
rect 3700 4575 3705 4675
rect 3740 4575 3760 4675
rect 3795 4575 3800 4675
rect 3700 4560 3800 4575
rect 3950 4675 4050 4690
rect 3950 4575 3955 4675
rect 3990 4575 4010 4675
rect 4045 4575 4050 4675
rect 3950 4560 4050 4575
rect 4200 4675 4300 4690
rect 4200 4575 4205 4675
rect 4240 4575 4260 4675
rect 4295 4575 4300 4675
rect 4200 4560 4300 4575
rect 4450 4675 4550 4690
rect 4450 4575 4455 4675
rect 4490 4575 4510 4675
rect 4545 4575 4550 4675
rect 4450 4560 4550 4575
rect 4700 4675 4800 4690
rect 4700 4575 4705 4675
rect 4740 4575 4760 4675
rect 4795 4575 4800 4675
rect 4700 4560 4800 4575
rect 4950 4675 5050 4690
rect 4950 4575 4955 4675
rect 4990 4575 5010 4675
rect 5045 4575 5050 4675
rect 4950 4560 5050 4575
rect 5200 4675 5300 4690
rect 5200 4575 5205 4675
rect 5240 4575 5260 4675
rect 5295 4575 5300 4675
rect 5200 4560 5300 4575
rect 5450 4675 5550 4690
rect 5450 4575 5455 4675
rect 5490 4575 5510 4675
rect 5545 4575 5550 4675
rect 5450 4560 5550 4575
rect 5700 4675 5800 4690
rect 5700 4575 5705 4675
rect 5740 4575 5760 4675
rect 5795 4575 5800 4675
rect 5700 4560 5800 4575
rect 5950 4675 6050 4690
rect 5950 4575 5955 4675
rect 5990 4575 6010 4675
rect 6045 4575 6050 4675
rect 5950 4560 6050 4575
rect 6200 4675 6300 4690
rect 6200 4575 6205 4675
rect 6240 4575 6260 4675
rect 6295 4575 6300 4675
rect 6200 4560 6300 4575
rect 6450 4675 6550 4690
rect 6450 4575 6455 4675
rect 6490 4575 6510 4675
rect 6545 4575 6550 4675
rect 6450 4560 6550 4575
rect 6700 4675 6800 4690
rect 6700 4575 6705 4675
rect 6740 4575 6760 4675
rect 6795 4575 6800 4675
rect 6700 4560 6800 4575
rect 6950 4675 7050 4690
rect 6950 4575 6955 4675
rect 6990 4575 7010 4675
rect 7045 4575 7050 4675
rect 6950 4560 7050 4575
rect 7200 4675 7300 4690
rect 7200 4575 7205 4675
rect 7240 4575 7260 4675
rect 7295 4575 7300 4675
rect 7200 4560 7300 4575
rect 7450 4675 7550 4690
rect 7450 4575 7455 4675
rect 7490 4575 7510 4675
rect 7545 4575 7550 4675
rect 7450 4560 7550 4575
rect 7700 4675 7800 4690
rect 7700 4575 7705 4675
rect 7740 4575 7760 4675
rect 7795 4575 7800 4675
rect 7700 4560 7800 4575
rect 7950 4675 8000 4690
rect 7950 4575 7955 4675
rect 7990 4575 8000 4675
rect 7950 4560 8000 4575
rect 0 4550 60 4560
rect 190 4550 310 4560
rect 440 4550 560 4560
rect 690 4550 810 4560
rect 940 4550 1060 4560
rect 1190 4550 1310 4560
rect 1440 4550 1560 4560
rect 1690 4550 1810 4560
rect 1940 4550 2060 4560
rect 2190 4550 2310 4560
rect 2440 4550 2560 4560
rect 2690 4550 2810 4560
rect 2940 4550 3060 4560
rect 3190 4550 3310 4560
rect 3440 4550 3560 4560
rect 3690 4550 3810 4560
rect 3940 4550 4060 4560
rect 4190 4550 4310 4560
rect 4440 4550 4560 4560
rect 4690 4550 4810 4560
rect 4940 4550 5060 4560
rect 5190 4550 5310 4560
rect 5440 4550 5560 4560
rect 5690 4550 5810 4560
rect 5940 4550 6060 4560
rect 6190 4550 6310 4560
rect 6440 4550 6560 4560
rect 6690 4550 6810 4560
rect 6940 4550 7060 4560
rect 7190 4550 7310 4560
rect 7440 4550 7560 4560
rect 7690 4550 7810 4560
rect 7940 4550 8000 4560
rect 0 4545 8000 4550
rect 0 4510 75 4545
rect 175 4510 325 4545
rect 425 4510 575 4545
rect 675 4510 825 4545
rect 925 4510 1075 4545
rect 1175 4510 1325 4545
rect 1425 4510 1575 4545
rect 1675 4510 1825 4545
rect 1925 4510 2075 4545
rect 2175 4510 2325 4545
rect 2425 4510 2575 4545
rect 2675 4510 2825 4545
rect 2925 4510 3075 4545
rect 3175 4510 3325 4545
rect 3425 4510 3575 4545
rect 3675 4510 3825 4545
rect 3925 4510 4075 4545
rect 4175 4510 4325 4545
rect 4425 4510 4575 4545
rect 4675 4510 4825 4545
rect 4925 4510 5075 4545
rect 5175 4510 5325 4545
rect 5425 4510 5575 4545
rect 5675 4510 5825 4545
rect 5925 4510 6075 4545
rect 6175 4510 6325 4545
rect 6425 4510 6575 4545
rect 6675 4510 6825 4545
rect 6925 4510 7075 4545
rect 7175 4510 7325 4545
rect 7425 4510 7575 4545
rect 7675 4510 7825 4545
rect 7925 4510 8000 4545
rect 0 4490 8000 4510
rect 0 4455 75 4490
rect 175 4455 325 4490
rect 425 4455 575 4490
rect 675 4455 825 4490
rect 925 4455 1075 4490
rect 1175 4455 1325 4490
rect 1425 4455 1575 4490
rect 1675 4455 1825 4490
rect 1925 4455 2075 4490
rect 2175 4455 2325 4490
rect 2425 4455 2575 4490
rect 2675 4455 2825 4490
rect 2925 4455 3075 4490
rect 3175 4455 3325 4490
rect 3425 4455 3575 4490
rect 3675 4455 3825 4490
rect 3925 4455 4075 4490
rect 4175 4455 4325 4490
rect 4425 4455 4575 4490
rect 4675 4455 4825 4490
rect 4925 4455 5075 4490
rect 5175 4455 5325 4490
rect 5425 4455 5575 4490
rect 5675 4455 5825 4490
rect 5925 4455 6075 4490
rect 6175 4455 6325 4490
rect 6425 4455 6575 4490
rect 6675 4455 6825 4490
rect 6925 4455 7075 4490
rect 7175 4455 7325 4490
rect 7425 4455 7575 4490
rect 7675 4455 7825 4490
rect 7925 4455 8000 4490
rect 0 4450 8000 4455
rect 0 4440 60 4450
rect 190 4440 310 4450
rect 440 4440 560 4450
rect 690 4440 810 4450
rect 940 4440 1060 4450
rect 1190 4440 1310 4450
rect 1440 4440 1560 4450
rect 1690 4440 1810 4450
rect 1940 4440 2060 4450
rect 2190 4440 2310 4450
rect 2440 4440 2560 4450
rect 2690 4440 2810 4450
rect 2940 4440 3060 4450
rect 3190 4440 3310 4450
rect 3440 4440 3560 4450
rect 3690 4440 3810 4450
rect 3940 4440 4060 4450
rect 4190 4440 4310 4450
rect 4440 4440 4560 4450
rect 4690 4440 4810 4450
rect 4940 4440 5060 4450
rect 5190 4440 5310 4450
rect 5440 4440 5560 4450
rect 5690 4440 5810 4450
rect 5940 4440 6060 4450
rect 6190 4440 6310 4450
rect 6440 4440 6560 4450
rect 6690 4440 6810 4450
rect 6940 4440 7060 4450
rect 7190 4440 7310 4450
rect 7440 4440 7560 4450
rect 7690 4440 7810 4450
rect 7940 4440 8000 4450
rect 0 4425 50 4440
rect 0 4325 10 4425
rect 45 4325 50 4425
rect 0 4310 50 4325
rect 200 4425 300 4440
rect 200 4325 205 4425
rect 240 4325 260 4425
rect 295 4325 300 4425
rect 200 4310 300 4325
rect 450 4425 550 4440
rect 450 4325 455 4425
rect 490 4325 510 4425
rect 545 4325 550 4425
rect 450 4310 550 4325
rect 700 4425 800 4440
rect 700 4325 705 4425
rect 740 4325 760 4425
rect 795 4325 800 4425
rect 700 4310 800 4325
rect 950 4425 1050 4440
rect 950 4325 955 4425
rect 990 4325 1010 4425
rect 1045 4325 1050 4425
rect 950 4310 1050 4325
rect 1200 4425 1300 4440
rect 1200 4325 1205 4425
rect 1240 4325 1260 4425
rect 1295 4325 1300 4425
rect 1200 4310 1300 4325
rect 1450 4425 1550 4440
rect 1450 4325 1455 4425
rect 1490 4325 1510 4425
rect 1545 4325 1550 4425
rect 1450 4310 1550 4325
rect 1700 4425 1800 4440
rect 1700 4325 1705 4425
rect 1740 4325 1760 4425
rect 1795 4325 1800 4425
rect 1700 4310 1800 4325
rect 1950 4425 2050 4440
rect 1950 4325 1955 4425
rect 1990 4325 2010 4425
rect 2045 4325 2050 4425
rect 1950 4310 2050 4325
rect 2200 4425 2300 4440
rect 2200 4325 2205 4425
rect 2240 4325 2260 4425
rect 2295 4325 2300 4425
rect 2200 4310 2300 4325
rect 2450 4425 2550 4440
rect 2450 4325 2455 4425
rect 2490 4325 2510 4425
rect 2545 4325 2550 4425
rect 2450 4310 2550 4325
rect 2700 4425 2800 4440
rect 2700 4325 2705 4425
rect 2740 4325 2760 4425
rect 2795 4325 2800 4425
rect 2700 4310 2800 4325
rect 2950 4425 3050 4440
rect 2950 4325 2955 4425
rect 2990 4325 3010 4425
rect 3045 4325 3050 4425
rect 2950 4310 3050 4325
rect 3200 4425 3300 4440
rect 3200 4325 3205 4425
rect 3240 4325 3260 4425
rect 3295 4325 3300 4425
rect 3200 4310 3300 4325
rect 3450 4425 3550 4440
rect 3450 4325 3455 4425
rect 3490 4325 3510 4425
rect 3545 4325 3550 4425
rect 3450 4310 3550 4325
rect 3700 4425 3800 4440
rect 3700 4325 3705 4425
rect 3740 4325 3760 4425
rect 3795 4325 3800 4425
rect 3700 4310 3800 4325
rect 3950 4425 4050 4440
rect 3950 4325 3955 4425
rect 3990 4325 4010 4425
rect 4045 4325 4050 4425
rect 3950 4310 4050 4325
rect 4200 4425 4300 4440
rect 4200 4325 4205 4425
rect 4240 4325 4260 4425
rect 4295 4325 4300 4425
rect 4200 4310 4300 4325
rect 4450 4425 4550 4440
rect 4450 4325 4455 4425
rect 4490 4325 4510 4425
rect 4545 4325 4550 4425
rect 4450 4310 4550 4325
rect 4700 4425 4800 4440
rect 4700 4325 4705 4425
rect 4740 4325 4760 4425
rect 4795 4325 4800 4425
rect 4700 4310 4800 4325
rect 4950 4425 5050 4440
rect 4950 4325 4955 4425
rect 4990 4325 5010 4425
rect 5045 4325 5050 4425
rect 4950 4310 5050 4325
rect 5200 4425 5300 4440
rect 5200 4325 5205 4425
rect 5240 4325 5260 4425
rect 5295 4325 5300 4425
rect 5200 4310 5300 4325
rect 5450 4425 5550 4440
rect 5450 4325 5455 4425
rect 5490 4325 5510 4425
rect 5545 4325 5550 4425
rect 5450 4310 5550 4325
rect 5700 4425 5800 4440
rect 5700 4325 5705 4425
rect 5740 4325 5760 4425
rect 5795 4325 5800 4425
rect 5700 4310 5800 4325
rect 5950 4425 6050 4440
rect 5950 4325 5955 4425
rect 5990 4325 6010 4425
rect 6045 4325 6050 4425
rect 5950 4310 6050 4325
rect 6200 4425 6300 4440
rect 6200 4325 6205 4425
rect 6240 4325 6260 4425
rect 6295 4325 6300 4425
rect 6200 4310 6300 4325
rect 6450 4425 6550 4440
rect 6450 4325 6455 4425
rect 6490 4325 6510 4425
rect 6545 4325 6550 4425
rect 6450 4310 6550 4325
rect 6700 4425 6800 4440
rect 6700 4325 6705 4425
rect 6740 4325 6760 4425
rect 6795 4325 6800 4425
rect 6700 4310 6800 4325
rect 6950 4425 7050 4440
rect 6950 4325 6955 4425
rect 6990 4325 7010 4425
rect 7045 4325 7050 4425
rect 6950 4310 7050 4325
rect 7200 4425 7300 4440
rect 7200 4325 7205 4425
rect 7240 4325 7260 4425
rect 7295 4325 7300 4425
rect 7200 4310 7300 4325
rect 7450 4425 7550 4440
rect 7450 4325 7455 4425
rect 7490 4325 7510 4425
rect 7545 4325 7550 4425
rect 7450 4310 7550 4325
rect 7700 4425 7800 4440
rect 7700 4325 7705 4425
rect 7740 4325 7760 4425
rect 7795 4325 7800 4425
rect 7700 4310 7800 4325
rect 7950 4425 8000 4440
rect 7950 4325 7955 4425
rect 7990 4325 8000 4425
rect 7950 4310 8000 4325
rect 0 4300 60 4310
rect 190 4300 310 4310
rect 440 4300 560 4310
rect 690 4300 810 4310
rect 940 4300 1060 4310
rect 1190 4300 1310 4310
rect 1440 4300 1560 4310
rect 1690 4300 1810 4310
rect 1940 4300 2060 4310
rect 2190 4300 2310 4310
rect 2440 4300 2560 4310
rect 2690 4300 2810 4310
rect 2940 4300 3060 4310
rect 3190 4300 3310 4310
rect 3440 4300 3560 4310
rect 3690 4300 3810 4310
rect 3940 4300 4060 4310
rect 4190 4300 4310 4310
rect 4440 4300 4560 4310
rect 4690 4300 4810 4310
rect 4940 4300 5060 4310
rect 5190 4300 5310 4310
rect 5440 4300 5560 4310
rect 5690 4300 5810 4310
rect 5940 4300 6060 4310
rect 6190 4300 6310 4310
rect 6440 4300 6560 4310
rect 6690 4300 6810 4310
rect 6940 4300 7060 4310
rect 7190 4300 7310 4310
rect 7440 4300 7560 4310
rect 7690 4300 7810 4310
rect 7940 4300 8000 4310
rect 0 4295 8000 4300
rect 0 4260 75 4295
rect 175 4260 325 4295
rect 425 4260 575 4295
rect 675 4260 825 4295
rect 925 4260 1075 4295
rect 1175 4260 1325 4295
rect 1425 4260 1575 4295
rect 1675 4260 1825 4295
rect 1925 4260 2075 4295
rect 2175 4260 2325 4295
rect 2425 4260 2575 4295
rect 2675 4260 2825 4295
rect 2925 4260 3075 4295
rect 3175 4260 3325 4295
rect 3425 4260 3575 4295
rect 3675 4260 3825 4295
rect 3925 4260 4075 4295
rect 4175 4260 4325 4295
rect 4425 4260 4575 4295
rect 4675 4260 4825 4295
rect 4925 4260 5075 4295
rect 5175 4260 5325 4295
rect 5425 4260 5575 4295
rect 5675 4260 5825 4295
rect 5925 4260 6075 4295
rect 6175 4260 6325 4295
rect 6425 4260 6575 4295
rect 6675 4260 6825 4295
rect 6925 4260 7075 4295
rect 7175 4260 7325 4295
rect 7425 4260 7575 4295
rect 7675 4260 7825 4295
rect 7925 4260 8000 4295
rect 0 4240 8000 4260
rect 0 4205 75 4240
rect 175 4205 325 4240
rect 425 4205 575 4240
rect 675 4205 825 4240
rect 925 4205 1075 4240
rect 1175 4205 1325 4240
rect 1425 4205 1575 4240
rect 1675 4205 1825 4240
rect 1925 4205 2075 4240
rect 2175 4205 2325 4240
rect 2425 4205 2575 4240
rect 2675 4205 2825 4240
rect 2925 4205 3075 4240
rect 3175 4205 3325 4240
rect 3425 4205 3575 4240
rect 3675 4205 3825 4240
rect 3925 4205 4075 4240
rect 4175 4205 4325 4240
rect 4425 4205 4575 4240
rect 4675 4205 4825 4240
rect 4925 4205 5075 4240
rect 5175 4205 5325 4240
rect 5425 4205 5575 4240
rect 5675 4205 5825 4240
rect 5925 4205 6075 4240
rect 6175 4205 6325 4240
rect 6425 4205 6575 4240
rect 6675 4205 6825 4240
rect 6925 4205 7075 4240
rect 7175 4205 7325 4240
rect 7425 4205 7575 4240
rect 7675 4205 7825 4240
rect 7925 4205 8000 4240
rect 0 4200 8000 4205
rect 0 4190 60 4200
rect 190 4190 310 4200
rect 440 4190 560 4200
rect 690 4190 810 4200
rect 940 4190 1060 4200
rect 1190 4190 1310 4200
rect 1440 4190 1560 4200
rect 1690 4190 1810 4200
rect 1940 4190 2060 4200
rect 2190 4190 2310 4200
rect 2440 4190 2560 4200
rect 2690 4190 2810 4200
rect 2940 4190 3060 4200
rect 3190 4190 3310 4200
rect 3440 4190 3560 4200
rect 3690 4190 3810 4200
rect 3940 4190 4060 4200
rect 4190 4190 4310 4200
rect 4440 4190 4560 4200
rect 4690 4190 4810 4200
rect 4940 4190 5060 4200
rect 5190 4190 5310 4200
rect 5440 4190 5560 4200
rect 5690 4190 5810 4200
rect 5940 4190 6060 4200
rect 6190 4190 6310 4200
rect 6440 4190 6560 4200
rect 6690 4190 6810 4200
rect 6940 4190 7060 4200
rect 7190 4190 7310 4200
rect 7440 4190 7560 4200
rect 7690 4190 7810 4200
rect 7940 4190 8000 4200
rect 0 4175 50 4190
rect 0 4075 10 4175
rect 45 4075 50 4175
rect 0 4060 50 4075
rect 200 4175 300 4190
rect 200 4075 205 4175
rect 240 4075 260 4175
rect 295 4075 300 4175
rect 200 4060 300 4075
rect 450 4175 550 4190
rect 450 4075 455 4175
rect 490 4075 510 4175
rect 545 4075 550 4175
rect 450 4060 550 4075
rect 700 4175 800 4190
rect 700 4075 705 4175
rect 740 4075 760 4175
rect 795 4075 800 4175
rect 700 4060 800 4075
rect 950 4175 1050 4190
rect 950 4075 955 4175
rect 990 4075 1010 4175
rect 1045 4075 1050 4175
rect 950 4060 1050 4075
rect 1200 4175 1300 4190
rect 1200 4075 1205 4175
rect 1240 4075 1260 4175
rect 1295 4075 1300 4175
rect 1200 4060 1300 4075
rect 1450 4175 1550 4190
rect 1450 4075 1455 4175
rect 1490 4075 1510 4175
rect 1545 4075 1550 4175
rect 1450 4060 1550 4075
rect 1700 4175 1800 4190
rect 1700 4075 1705 4175
rect 1740 4075 1760 4175
rect 1795 4075 1800 4175
rect 1700 4060 1800 4075
rect 1950 4175 2050 4190
rect 1950 4075 1955 4175
rect 1990 4075 2010 4175
rect 2045 4075 2050 4175
rect 1950 4060 2050 4075
rect 2200 4175 2300 4190
rect 2200 4075 2205 4175
rect 2240 4075 2260 4175
rect 2295 4075 2300 4175
rect 2200 4060 2300 4075
rect 2450 4175 2550 4190
rect 2450 4075 2455 4175
rect 2490 4075 2510 4175
rect 2545 4075 2550 4175
rect 2450 4060 2550 4075
rect 2700 4175 2800 4190
rect 2700 4075 2705 4175
rect 2740 4075 2760 4175
rect 2795 4075 2800 4175
rect 2700 4060 2800 4075
rect 2950 4175 3050 4190
rect 2950 4075 2955 4175
rect 2990 4075 3010 4175
rect 3045 4075 3050 4175
rect 2950 4060 3050 4075
rect 3200 4175 3300 4190
rect 3200 4075 3205 4175
rect 3240 4075 3260 4175
rect 3295 4075 3300 4175
rect 3200 4060 3300 4075
rect 3450 4175 3550 4190
rect 3450 4075 3455 4175
rect 3490 4075 3510 4175
rect 3545 4075 3550 4175
rect 3450 4060 3550 4075
rect 3700 4175 3800 4190
rect 3700 4075 3705 4175
rect 3740 4075 3760 4175
rect 3795 4075 3800 4175
rect 3700 4060 3800 4075
rect 3950 4175 4050 4190
rect 3950 4075 3955 4175
rect 3990 4075 4010 4175
rect 4045 4075 4050 4175
rect 3950 4060 4050 4075
rect 4200 4175 4300 4190
rect 4200 4075 4205 4175
rect 4240 4075 4260 4175
rect 4295 4075 4300 4175
rect 4200 4060 4300 4075
rect 4450 4175 4550 4190
rect 4450 4075 4455 4175
rect 4490 4075 4510 4175
rect 4545 4075 4550 4175
rect 4450 4060 4550 4075
rect 4700 4175 4800 4190
rect 4700 4075 4705 4175
rect 4740 4075 4760 4175
rect 4795 4075 4800 4175
rect 4700 4060 4800 4075
rect 4950 4175 5050 4190
rect 4950 4075 4955 4175
rect 4990 4075 5010 4175
rect 5045 4075 5050 4175
rect 4950 4060 5050 4075
rect 5200 4175 5300 4190
rect 5200 4075 5205 4175
rect 5240 4075 5260 4175
rect 5295 4075 5300 4175
rect 5200 4060 5300 4075
rect 5450 4175 5550 4190
rect 5450 4075 5455 4175
rect 5490 4075 5510 4175
rect 5545 4075 5550 4175
rect 5450 4060 5550 4075
rect 5700 4175 5800 4190
rect 5700 4075 5705 4175
rect 5740 4075 5760 4175
rect 5795 4075 5800 4175
rect 5700 4060 5800 4075
rect 5950 4175 6050 4190
rect 5950 4075 5955 4175
rect 5990 4075 6010 4175
rect 6045 4075 6050 4175
rect 5950 4060 6050 4075
rect 6200 4175 6300 4190
rect 6200 4075 6205 4175
rect 6240 4075 6260 4175
rect 6295 4075 6300 4175
rect 6200 4060 6300 4075
rect 6450 4175 6550 4190
rect 6450 4075 6455 4175
rect 6490 4075 6510 4175
rect 6545 4075 6550 4175
rect 6450 4060 6550 4075
rect 6700 4175 6800 4190
rect 6700 4075 6705 4175
rect 6740 4075 6760 4175
rect 6795 4075 6800 4175
rect 6700 4060 6800 4075
rect 6950 4175 7050 4190
rect 6950 4075 6955 4175
rect 6990 4075 7010 4175
rect 7045 4075 7050 4175
rect 6950 4060 7050 4075
rect 7200 4175 7300 4190
rect 7200 4075 7205 4175
rect 7240 4075 7260 4175
rect 7295 4075 7300 4175
rect 7200 4060 7300 4075
rect 7450 4175 7550 4190
rect 7450 4075 7455 4175
rect 7490 4075 7510 4175
rect 7545 4075 7550 4175
rect 7450 4060 7550 4075
rect 7700 4175 7800 4190
rect 7700 4075 7705 4175
rect 7740 4075 7760 4175
rect 7795 4075 7800 4175
rect 7700 4060 7800 4075
rect 7950 4175 8000 4190
rect 7950 4075 7955 4175
rect 7990 4075 8000 4175
rect 7950 4060 8000 4075
rect 0 4050 60 4060
rect 190 4050 310 4060
rect 440 4050 560 4060
rect 690 4050 810 4060
rect 940 4050 1060 4060
rect 1190 4050 1310 4060
rect 1440 4050 1560 4060
rect 1690 4050 1810 4060
rect 1940 4050 2060 4060
rect 2190 4050 2310 4060
rect 2440 4050 2560 4060
rect 2690 4050 2810 4060
rect 2940 4050 3060 4060
rect 3190 4050 3310 4060
rect 3440 4050 3560 4060
rect 3690 4050 3810 4060
rect 3940 4050 4060 4060
rect 4190 4050 4310 4060
rect 4440 4050 4560 4060
rect 4690 4050 4810 4060
rect 4940 4050 5060 4060
rect 5190 4050 5310 4060
rect 5440 4050 5560 4060
rect 5690 4050 5810 4060
rect 5940 4050 6060 4060
rect 6190 4050 6310 4060
rect 6440 4050 6560 4060
rect 6690 4050 6810 4060
rect 6940 4050 7060 4060
rect 7190 4050 7310 4060
rect 7440 4050 7560 4060
rect 7690 4050 7810 4060
rect 7940 4050 8000 4060
rect 0 4045 8000 4050
rect 0 4010 75 4045
rect 175 4010 325 4045
rect 425 4010 575 4045
rect 675 4010 825 4045
rect 925 4010 1075 4045
rect 1175 4010 1325 4045
rect 1425 4010 1575 4045
rect 1675 4010 1825 4045
rect 1925 4010 2075 4045
rect 2175 4010 2325 4045
rect 2425 4010 2575 4045
rect 2675 4010 2825 4045
rect 2925 4010 3075 4045
rect 3175 4010 3325 4045
rect 3425 4010 3575 4045
rect 3675 4010 3825 4045
rect 3925 4010 4075 4045
rect 4175 4010 4325 4045
rect 4425 4010 4575 4045
rect 4675 4010 4825 4045
rect 4925 4010 5075 4045
rect 5175 4010 5325 4045
rect 5425 4010 5575 4045
rect 5675 4010 5825 4045
rect 5925 4010 6075 4045
rect 6175 4010 6325 4045
rect 6425 4010 6575 4045
rect 6675 4010 6825 4045
rect 6925 4010 7075 4045
rect 7175 4010 7325 4045
rect 7425 4010 7575 4045
rect 7675 4010 7825 4045
rect 7925 4010 8000 4045
rect 0 3990 8000 4010
rect 0 3955 75 3990
rect 175 3955 325 3990
rect 425 3955 575 3990
rect 675 3955 825 3990
rect 925 3955 1075 3990
rect 1175 3955 1325 3990
rect 1425 3955 1575 3990
rect 1675 3955 1825 3990
rect 1925 3955 2075 3990
rect 2175 3955 2325 3990
rect 2425 3955 2575 3990
rect 2675 3955 2825 3990
rect 2925 3955 3075 3990
rect 3175 3955 3325 3990
rect 3425 3955 3575 3990
rect 3675 3955 3825 3990
rect 3925 3955 4075 3990
rect 4175 3955 4325 3990
rect 4425 3955 4575 3990
rect 4675 3955 4825 3990
rect 4925 3955 5075 3990
rect 5175 3955 5325 3990
rect 5425 3955 5575 3990
rect 5675 3955 5825 3990
rect 5925 3955 6075 3990
rect 6175 3955 6325 3990
rect 6425 3955 6575 3990
rect 6675 3955 6825 3990
rect 6925 3955 7075 3990
rect 7175 3955 7325 3990
rect 7425 3955 7575 3990
rect 7675 3955 7825 3990
rect 7925 3955 8000 3990
rect 0 3950 8000 3955
rect 0 3940 60 3950
rect 190 3940 310 3950
rect 440 3940 560 3950
rect 690 3940 810 3950
rect 940 3940 1060 3950
rect 1190 3940 1310 3950
rect 1440 3940 1560 3950
rect 1690 3940 1810 3950
rect 1940 3940 2060 3950
rect 2190 3940 2310 3950
rect 2440 3940 2560 3950
rect 2690 3940 2810 3950
rect 2940 3940 3060 3950
rect 3190 3940 3310 3950
rect 3440 3940 3560 3950
rect 3690 3940 3810 3950
rect 3940 3940 4060 3950
rect 4190 3940 4310 3950
rect 4440 3940 4560 3950
rect 4690 3940 4810 3950
rect 4940 3940 5060 3950
rect 5190 3940 5310 3950
rect 5440 3940 5560 3950
rect 5690 3940 5810 3950
rect 5940 3940 6060 3950
rect 6190 3940 6310 3950
rect 6440 3940 6560 3950
rect 6690 3940 6810 3950
rect 6940 3940 7060 3950
rect 7190 3940 7310 3950
rect 7440 3940 7560 3950
rect 7690 3940 7810 3950
rect 7940 3940 8000 3950
rect 0 3925 50 3940
rect 0 3825 10 3925
rect 45 3825 50 3925
rect 0 3810 50 3825
rect 200 3925 300 3940
rect 200 3825 205 3925
rect 240 3825 260 3925
rect 295 3825 300 3925
rect 200 3810 300 3825
rect 450 3925 550 3940
rect 450 3825 455 3925
rect 490 3825 510 3925
rect 545 3825 550 3925
rect 450 3810 550 3825
rect 700 3925 800 3940
rect 700 3825 705 3925
rect 740 3825 760 3925
rect 795 3825 800 3925
rect 700 3810 800 3825
rect 950 3925 1050 3940
rect 950 3825 955 3925
rect 990 3825 1010 3925
rect 1045 3825 1050 3925
rect 950 3810 1050 3825
rect 1200 3925 1300 3940
rect 1200 3825 1205 3925
rect 1240 3825 1260 3925
rect 1295 3825 1300 3925
rect 1200 3810 1300 3825
rect 1450 3925 1550 3940
rect 1450 3825 1455 3925
rect 1490 3825 1510 3925
rect 1545 3825 1550 3925
rect 1450 3810 1550 3825
rect 1700 3925 1800 3940
rect 1700 3825 1705 3925
rect 1740 3825 1760 3925
rect 1795 3825 1800 3925
rect 1700 3810 1800 3825
rect 1950 3925 2050 3940
rect 1950 3825 1955 3925
rect 1990 3825 2010 3925
rect 2045 3825 2050 3925
rect 1950 3810 2050 3825
rect 2200 3925 2300 3940
rect 2200 3825 2205 3925
rect 2240 3825 2260 3925
rect 2295 3825 2300 3925
rect 2200 3810 2300 3825
rect 2450 3925 2550 3940
rect 2450 3825 2455 3925
rect 2490 3825 2510 3925
rect 2545 3825 2550 3925
rect 2450 3810 2550 3825
rect 2700 3925 2800 3940
rect 2700 3825 2705 3925
rect 2740 3825 2760 3925
rect 2795 3825 2800 3925
rect 2700 3810 2800 3825
rect 2950 3925 3050 3940
rect 2950 3825 2955 3925
rect 2990 3825 3010 3925
rect 3045 3825 3050 3925
rect 2950 3810 3050 3825
rect 3200 3925 3300 3940
rect 3200 3825 3205 3925
rect 3240 3825 3260 3925
rect 3295 3825 3300 3925
rect 3200 3810 3300 3825
rect 3450 3925 3550 3940
rect 3450 3825 3455 3925
rect 3490 3825 3510 3925
rect 3545 3825 3550 3925
rect 3450 3810 3550 3825
rect 3700 3925 3800 3940
rect 3700 3825 3705 3925
rect 3740 3825 3760 3925
rect 3795 3825 3800 3925
rect 3700 3810 3800 3825
rect 3950 3925 4050 3940
rect 3950 3825 3955 3925
rect 3990 3825 4010 3925
rect 4045 3825 4050 3925
rect 3950 3810 4050 3825
rect 4200 3925 4300 3940
rect 4200 3825 4205 3925
rect 4240 3825 4260 3925
rect 4295 3825 4300 3925
rect 4200 3810 4300 3825
rect 4450 3925 4550 3940
rect 4450 3825 4455 3925
rect 4490 3825 4510 3925
rect 4545 3825 4550 3925
rect 4450 3810 4550 3825
rect 4700 3925 4800 3940
rect 4700 3825 4705 3925
rect 4740 3825 4760 3925
rect 4795 3825 4800 3925
rect 4700 3810 4800 3825
rect 4950 3925 5050 3940
rect 4950 3825 4955 3925
rect 4990 3825 5010 3925
rect 5045 3825 5050 3925
rect 4950 3810 5050 3825
rect 5200 3925 5300 3940
rect 5200 3825 5205 3925
rect 5240 3825 5260 3925
rect 5295 3825 5300 3925
rect 5200 3810 5300 3825
rect 5450 3925 5550 3940
rect 5450 3825 5455 3925
rect 5490 3825 5510 3925
rect 5545 3825 5550 3925
rect 5450 3810 5550 3825
rect 5700 3925 5800 3940
rect 5700 3825 5705 3925
rect 5740 3825 5760 3925
rect 5795 3825 5800 3925
rect 5700 3810 5800 3825
rect 5950 3925 6050 3940
rect 5950 3825 5955 3925
rect 5990 3825 6010 3925
rect 6045 3825 6050 3925
rect 5950 3810 6050 3825
rect 6200 3925 6300 3940
rect 6200 3825 6205 3925
rect 6240 3825 6260 3925
rect 6295 3825 6300 3925
rect 6200 3810 6300 3825
rect 6450 3925 6550 3940
rect 6450 3825 6455 3925
rect 6490 3825 6510 3925
rect 6545 3825 6550 3925
rect 6450 3810 6550 3825
rect 6700 3925 6800 3940
rect 6700 3825 6705 3925
rect 6740 3825 6760 3925
rect 6795 3825 6800 3925
rect 6700 3810 6800 3825
rect 6950 3925 7050 3940
rect 6950 3825 6955 3925
rect 6990 3825 7010 3925
rect 7045 3825 7050 3925
rect 6950 3810 7050 3825
rect 7200 3925 7300 3940
rect 7200 3825 7205 3925
rect 7240 3825 7260 3925
rect 7295 3825 7300 3925
rect 7200 3810 7300 3825
rect 7450 3925 7550 3940
rect 7450 3825 7455 3925
rect 7490 3825 7510 3925
rect 7545 3825 7550 3925
rect 7450 3810 7550 3825
rect 7700 3925 7800 3940
rect 7700 3825 7705 3925
rect 7740 3825 7760 3925
rect 7795 3825 7800 3925
rect 7700 3810 7800 3825
rect 7950 3925 8000 3940
rect 7950 3825 7955 3925
rect 7990 3825 8000 3925
rect 7950 3810 8000 3825
rect 0 3800 60 3810
rect 190 3800 310 3810
rect 440 3800 560 3810
rect 690 3800 810 3810
rect 940 3800 1060 3810
rect 1190 3800 1310 3810
rect 1440 3800 1560 3810
rect 1690 3800 1810 3810
rect 1940 3800 2060 3810
rect 2190 3800 2310 3810
rect 2440 3800 2560 3810
rect 2690 3800 2810 3810
rect 2940 3800 3060 3810
rect 3190 3800 3310 3810
rect 3440 3800 3560 3810
rect 3690 3800 3810 3810
rect 3940 3800 4060 3810
rect 4190 3800 4310 3810
rect 4440 3800 4560 3810
rect 4690 3800 4810 3810
rect 4940 3800 5060 3810
rect 5190 3800 5310 3810
rect 5440 3800 5560 3810
rect 5690 3800 5810 3810
rect 5940 3800 6060 3810
rect 6190 3800 6310 3810
rect 6440 3800 6560 3810
rect 6690 3800 6810 3810
rect 6940 3800 7060 3810
rect 7190 3800 7310 3810
rect 7440 3800 7560 3810
rect 7690 3800 7810 3810
rect 7940 3800 8000 3810
rect 0 3795 8000 3800
rect 0 3760 75 3795
rect 175 3760 325 3795
rect 425 3760 575 3795
rect 675 3760 825 3795
rect 925 3760 1075 3795
rect 1175 3760 1325 3795
rect 1425 3760 1575 3795
rect 1675 3760 1825 3795
rect 1925 3760 2075 3795
rect 2175 3760 2325 3795
rect 2425 3760 2575 3795
rect 2675 3760 2825 3795
rect 2925 3760 3075 3795
rect 3175 3760 3325 3795
rect 3425 3760 3575 3795
rect 3675 3760 3825 3795
rect 3925 3760 4075 3795
rect 4175 3760 4325 3795
rect 4425 3760 4575 3795
rect 4675 3760 4825 3795
rect 4925 3760 5075 3795
rect 5175 3760 5325 3795
rect 5425 3760 5575 3795
rect 5675 3760 5825 3795
rect 5925 3760 6075 3795
rect 6175 3760 6325 3795
rect 6425 3760 6575 3795
rect 6675 3760 6825 3795
rect 6925 3760 7075 3795
rect 7175 3760 7325 3795
rect 7425 3760 7575 3795
rect 7675 3760 7825 3795
rect 7925 3760 8000 3795
rect 0 3740 8000 3760
rect 0 3705 75 3740
rect 175 3705 325 3740
rect 425 3705 575 3740
rect 675 3705 825 3740
rect 925 3705 1075 3740
rect 1175 3705 1325 3740
rect 1425 3705 1575 3740
rect 1675 3705 1825 3740
rect 1925 3705 2075 3740
rect 2175 3705 2325 3740
rect 2425 3705 2575 3740
rect 2675 3705 2825 3740
rect 2925 3705 3075 3740
rect 3175 3705 3325 3740
rect 3425 3705 3575 3740
rect 3675 3705 3825 3740
rect 3925 3705 4075 3740
rect 4175 3705 4325 3740
rect 4425 3705 4575 3740
rect 4675 3705 4825 3740
rect 4925 3705 5075 3740
rect 5175 3705 5325 3740
rect 5425 3705 5575 3740
rect 5675 3705 5825 3740
rect 5925 3705 6075 3740
rect 6175 3705 6325 3740
rect 6425 3705 6575 3740
rect 6675 3705 6825 3740
rect 6925 3705 7075 3740
rect 7175 3705 7325 3740
rect 7425 3705 7575 3740
rect 7675 3705 7825 3740
rect 7925 3705 8000 3740
rect 0 3700 8000 3705
rect 0 3690 60 3700
rect 190 3690 310 3700
rect 440 3690 560 3700
rect 690 3690 810 3700
rect 940 3690 1060 3700
rect 1190 3690 1310 3700
rect 1440 3690 1560 3700
rect 1690 3690 1810 3700
rect 1940 3690 2060 3700
rect 2190 3690 2310 3700
rect 2440 3690 2560 3700
rect 2690 3690 2810 3700
rect 2940 3690 3060 3700
rect 3190 3690 3310 3700
rect 3440 3690 3560 3700
rect 3690 3690 3810 3700
rect 3940 3690 4060 3700
rect 4190 3690 4310 3700
rect 4440 3690 4560 3700
rect 4690 3690 4810 3700
rect 4940 3690 5060 3700
rect 5190 3690 5310 3700
rect 5440 3690 5560 3700
rect 5690 3690 5810 3700
rect 5940 3690 6060 3700
rect 6190 3690 6310 3700
rect 6440 3690 6560 3700
rect 6690 3690 6810 3700
rect 6940 3690 7060 3700
rect 7190 3690 7310 3700
rect 7440 3690 7560 3700
rect 7690 3690 7810 3700
rect 7940 3690 8000 3700
rect 0 3675 50 3690
rect 0 3575 10 3675
rect 45 3575 50 3675
rect 0 3560 50 3575
rect 200 3675 300 3690
rect 200 3575 205 3675
rect 240 3575 260 3675
rect 295 3575 300 3675
rect 200 3560 300 3575
rect 450 3675 550 3690
rect 450 3575 455 3675
rect 490 3575 510 3675
rect 545 3575 550 3675
rect 450 3560 550 3575
rect 700 3675 800 3690
rect 700 3575 705 3675
rect 740 3575 760 3675
rect 795 3575 800 3675
rect 700 3560 800 3575
rect 950 3675 1050 3690
rect 950 3575 955 3675
rect 990 3575 1010 3675
rect 1045 3575 1050 3675
rect 950 3560 1050 3575
rect 1200 3675 1300 3690
rect 1200 3575 1205 3675
rect 1240 3575 1260 3675
rect 1295 3575 1300 3675
rect 1200 3560 1300 3575
rect 1450 3675 1550 3690
rect 1450 3575 1455 3675
rect 1490 3575 1510 3675
rect 1545 3575 1550 3675
rect 1450 3560 1550 3575
rect 1700 3675 1800 3690
rect 1700 3575 1705 3675
rect 1740 3575 1760 3675
rect 1795 3575 1800 3675
rect 1700 3560 1800 3575
rect 1950 3675 2050 3690
rect 1950 3575 1955 3675
rect 1990 3575 2010 3675
rect 2045 3575 2050 3675
rect 1950 3560 2050 3575
rect 2200 3675 2300 3690
rect 2200 3575 2205 3675
rect 2240 3575 2260 3675
rect 2295 3575 2300 3675
rect 2200 3560 2300 3575
rect 2450 3675 2550 3690
rect 2450 3575 2455 3675
rect 2490 3575 2510 3675
rect 2545 3575 2550 3675
rect 2450 3560 2550 3575
rect 2700 3675 2800 3690
rect 2700 3575 2705 3675
rect 2740 3575 2760 3675
rect 2795 3575 2800 3675
rect 2700 3560 2800 3575
rect 2950 3675 3050 3690
rect 2950 3575 2955 3675
rect 2990 3575 3010 3675
rect 3045 3575 3050 3675
rect 2950 3560 3050 3575
rect 3200 3675 3300 3690
rect 3200 3575 3205 3675
rect 3240 3575 3260 3675
rect 3295 3575 3300 3675
rect 3200 3560 3300 3575
rect 3450 3675 3550 3690
rect 3450 3575 3455 3675
rect 3490 3575 3510 3675
rect 3545 3575 3550 3675
rect 3450 3560 3550 3575
rect 3700 3675 3800 3690
rect 3700 3575 3705 3675
rect 3740 3575 3760 3675
rect 3795 3575 3800 3675
rect 3700 3560 3800 3575
rect 3950 3675 4050 3690
rect 3950 3575 3955 3675
rect 3990 3575 4010 3675
rect 4045 3575 4050 3675
rect 3950 3560 4050 3575
rect 4200 3675 4300 3690
rect 4200 3575 4205 3675
rect 4240 3575 4260 3675
rect 4295 3575 4300 3675
rect 4200 3560 4300 3575
rect 4450 3675 4550 3690
rect 4450 3575 4455 3675
rect 4490 3575 4510 3675
rect 4545 3575 4550 3675
rect 4450 3560 4550 3575
rect 4700 3675 4800 3690
rect 4700 3575 4705 3675
rect 4740 3575 4760 3675
rect 4795 3575 4800 3675
rect 4700 3560 4800 3575
rect 4950 3675 5050 3690
rect 4950 3575 4955 3675
rect 4990 3575 5010 3675
rect 5045 3575 5050 3675
rect 4950 3560 5050 3575
rect 5200 3675 5300 3690
rect 5200 3575 5205 3675
rect 5240 3575 5260 3675
rect 5295 3575 5300 3675
rect 5200 3560 5300 3575
rect 5450 3675 5550 3690
rect 5450 3575 5455 3675
rect 5490 3575 5510 3675
rect 5545 3575 5550 3675
rect 5450 3560 5550 3575
rect 5700 3675 5800 3690
rect 5700 3575 5705 3675
rect 5740 3575 5760 3675
rect 5795 3575 5800 3675
rect 5700 3560 5800 3575
rect 5950 3675 6050 3690
rect 5950 3575 5955 3675
rect 5990 3575 6010 3675
rect 6045 3575 6050 3675
rect 5950 3560 6050 3575
rect 6200 3675 6300 3690
rect 6200 3575 6205 3675
rect 6240 3575 6260 3675
rect 6295 3575 6300 3675
rect 6200 3560 6300 3575
rect 6450 3675 6550 3690
rect 6450 3575 6455 3675
rect 6490 3575 6510 3675
rect 6545 3575 6550 3675
rect 6450 3560 6550 3575
rect 6700 3675 6800 3690
rect 6700 3575 6705 3675
rect 6740 3575 6760 3675
rect 6795 3575 6800 3675
rect 6700 3560 6800 3575
rect 6950 3675 7050 3690
rect 6950 3575 6955 3675
rect 6990 3575 7010 3675
rect 7045 3575 7050 3675
rect 6950 3560 7050 3575
rect 7200 3675 7300 3690
rect 7200 3575 7205 3675
rect 7240 3575 7260 3675
rect 7295 3575 7300 3675
rect 7200 3560 7300 3575
rect 7450 3675 7550 3690
rect 7450 3575 7455 3675
rect 7490 3575 7510 3675
rect 7545 3575 7550 3675
rect 7450 3560 7550 3575
rect 7700 3675 7800 3690
rect 7700 3575 7705 3675
rect 7740 3575 7760 3675
rect 7795 3575 7800 3675
rect 7700 3560 7800 3575
rect 7950 3675 8000 3690
rect 7950 3575 7955 3675
rect 7990 3575 8000 3675
rect 7950 3560 8000 3575
rect 0 3550 60 3560
rect 190 3550 310 3560
rect 440 3550 560 3560
rect 690 3550 810 3560
rect 940 3550 1060 3560
rect 1190 3550 1310 3560
rect 1440 3550 1560 3560
rect 1690 3550 1810 3560
rect 1940 3550 2060 3560
rect 2190 3550 2310 3560
rect 2440 3550 2560 3560
rect 2690 3550 2810 3560
rect 2940 3550 3060 3560
rect 3190 3550 3310 3560
rect 3440 3550 3560 3560
rect 3690 3550 3810 3560
rect 3940 3550 4060 3560
rect 4190 3550 4310 3560
rect 4440 3550 4560 3560
rect 4690 3550 4810 3560
rect 4940 3550 5060 3560
rect 5190 3550 5310 3560
rect 5440 3550 5560 3560
rect 5690 3550 5810 3560
rect 5940 3550 6060 3560
rect 6190 3550 6310 3560
rect 6440 3550 6560 3560
rect 6690 3550 6810 3560
rect 6940 3550 7060 3560
rect 7190 3550 7310 3560
rect 7440 3550 7560 3560
rect 7690 3550 7810 3560
rect 7940 3550 8000 3560
rect 0 3545 8000 3550
rect 0 3510 75 3545
rect 175 3510 325 3545
rect 425 3510 575 3545
rect 675 3510 825 3545
rect 925 3510 1075 3545
rect 1175 3510 1325 3545
rect 1425 3510 1575 3545
rect 1675 3510 1825 3545
rect 1925 3510 2075 3545
rect 2175 3510 2325 3545
rect 2425 3510 2575 3545
rect 2675 3510 2825 3545
rect 2925 3510 3075 3545
rect 3175 3510 3325 3545
rect 3425 3510 3575 3545
rect 3675 3510 3825 3545
rect 3925 3510 4075 3545
rect 4175 3510 4325 3545
rect 4425 3510 4575 3545
rect 4675 3510 4825 3545
rect 4925 3510 5075 3545
rect 5175 3510 5325 3545
rect 5425 3510 5575 3545
rect 5675 3510 5825 3545
rect 5925 3510 6075 3545
rect 6175 3510 6325 3545
rect 6425 3510 6575 3545
rect 6675 3510 6825 3545
rect 6925 3510 7075 3545
rect 7175 3510 7325 3545
rect 7425 3510 7575 3545
rect 7675 3510 7825 3545
rect 7925 3510 8000 3545
rect 0 3490 8000 3510
rect 0 3455 75 3490
rect 175 3455 325 3490
rect 425 3455 575 3490
rect 675 3455 825 3490
rect 925 3455 1075 3490
rect 1175 3455 1325 3490
rect 1425 3455 1575 3490
rect 1675 3455 1825 3490
rect 1925 3455 2075 3490
rect 2175 3455 2325 3490
rect 2425 3455 2575 3490
rect 2675 3455 2825 3490
rect 2925 3455 3075 3490
rect 3175 3455 3325 3490
rect 3425 3455 3575 3490
rect 3675 3455 3825 3490
rect 3925 3455 4075 3490
rect 4175 3455 4325 3490
rect 4425 3455 4575 3490
rect 4675 3455 4825 3490
rect 4925 3455 5075 3490
rect 5175 3455 5325 3490
rect 5425 3455 5575 3490
rect 5675 3455 5825 3490
rect 5925 3455 6075 3490
rect 6175 3455 6325 3490
rect 6425 3455 6575 3490
rect 6675 3455 6825 3490
rect 6925 3455 7075 3490
rect 7175 3455 7325 3490
rect 7425 3455 7575 3490
rect 7675 3455 7825 3490
rect 7925 3455 8000 3490
rect 0 3450 8000 3455
rect 0 3440 60 3450
rect 190 3440 310 3450
rect 440 3440 560 3450
rect 690 3440 810 3450
rect 940 3440 1060 3450
rect 1190 3440 1310 3450
rect 1440 3440 1560 3450
rect 1690 3440 1810 3450
rect 1940 3440 2060 3450
rect 2190 3440 2310 3450
rect 2440 3440 2560 3450
rect 2690 3440 2810 3450
rect 2940 3440 3060 3450
rect 3190 3440 3310 3450
rect 3440 3440 3560 3450
rect 3690 3440 3810 3450
rect 3940 3440 4060 3450
rect 4190 3440 4310 3450
rect 4440 3440 4560 3450
rect 4690 3440 4810 3450
rect 4940 3440 5060 3450
rect 5190 3440 5310 3450
rect 5440 3440 5560 3450
rect 5690 3440 5810 3450
rect 5940 3440 6060 3450
rect 6190 3440 6310 3450
rect 6440 3440 6560 3450
rect 6690 3440 6810 3450
rect 6940 3440 7060 3450
rect 7190 3440 7310 3450
rect 7440 3440 7560 3450
rect 7690 3440 7810 3450
rect 7940 3440 8000 3450
rect 0 3425 50 3440
rect 0 3325 10 3425
rect 45 3325 50 3425
rect 0 3310 50 3325
rect 200 3425 300 3440
rect 200 3325 205 3425
rect 240 3325 260 3425
rect 295 3325 300 3425
rect 200 3310 300 3325
rect 450 3425 550 3440
rect 450 3325 455 3425
rect 490 3325 510 3425
rect 545 3325 550 3425
rect 450 3310 550 3325
rect 700 3425 800 3440
rect 700 3325 705 3425
rect 740 3325 760 3425
rect 795 3325 800 3425
rect 700 3310 800 3325
rect 950 3425 1050 3440
rect 950 3325 955 3425
rect 990 3325 1010 3425
rect 1045 3325 1050 3425
rect 950 3310 1050 3325
rect 1200 3425 1300 3440
rect 1200 3325 1205 3425
rect 1240 3325 1260 3425
rect 1295 3325 1300 3425
rect 1200 3310 1300 3325
rect 1450 3425 1550 3440
rect 1450 3325 1455 3425
rect 1490 3325 1510 3425
rect 1545 3325 1550 3425
rect 1450 3310 1550 3325
rect 1700 3425 1800 3440
rect 1700 3325 1705 3425
rect 1740 3325 1760 3425
rect 1795 3325 1800 3425
rect 1700 3310 1800 3325
rect 1950 3425 2050 3440
rect 1950 3325 1955 3425
rect 1990 3325 2010 3425
rect 2045 3325 2050 3425
rect 1950 3310 2050 3325
rect 2200 3425 2300 3440
rect 2200 3325 2205 3425
rect 2240 3325 2260 3425
rect 2295 3325 2300 3425
rect 2200 3310 2300 3325
rect 2450 3425 2550 3440
rect 2450 3325 2455 3425
rect 2490 3325 2510 3425
rect 2545 3325 2550 3425
rect 2450 3310 2550 3325
rect 2700 3425 2800 3440
rect 2700 3325 2705 3425
rect 2740 3325 2760 3425
rect 2795 3325 2800 3425
rect 2700 3310 2800 3325
rect 2950 3425 3050 3440
rect 2950 3325 2955 3425
rect 2990 3325 3010 3425
rect 3045 3325 3050 3425
rect 2950 3310 3050 3325
rect 3200 3425 3300 3440
rect 3200 3325 3205 3425
rect 3240 3325 3260 3425
rect 3295 3325 3300 3425
rect 3200 3310 3300 3325
rect 3450 3425 3550 3440
rect 3450 3325 3455 3425
rect 3490 3325 3510 3425
rect 3545 3325 3550 3425
rect 3450 3310 3550 3325
rect 3700 3425 3800 3440
rect 3700 3325 3705 3425
rect 3740 3325 3760 3425
rect 3795 3325 3800 3425
rect 3700 3310 3800 3325
rect 3950 3425 4050 3440
rect 3950 3325 3955 3425
rect 3990 3325 4010 3425
rect 4045 3325 4050 3425
rect 3950 3310 4050 3325
rect 4200 3425 4300 3440
rect 4200 3325 4205 3425
rect 4240 3325 4260 3425
rect 4295 3325 4300 3425
rect 4200 3310 4300 3325
rect 4450 3425 4550 3440
rect 4450 3325 4455 3425
rect 4490 3325 4510 3425
rect 4545 3325 4550 3425
rect 4450 3310 4550 3325
rect 4700 3425 4800 3440
rect 4700 3325 4705 3425
rect 4740 3325 4760 3425
rect 4795 3325 4800 3425
rect 4700 3310 4800 3325
rect 4950 3425 5050 3440
rect 4950 3325 4955 3425
rect 4990 3325 5010 3425
rect 5045 3325 5050 3425
rect 4950 3310 5050 3325
rect 5200 3425 5300 3440
rect 5200 3325 5205 3425
rect 5240 3325 5260 3425
rect 5295 3325 5300 3425
rect 5200 3310 5300 3325
rect 5450 3425 5550 3440
rect 5450 3325 5455 3425
rect 5490 3325 5510 3425
rect 5545 3325 5550 3425
rect 5450 3310 5550 3325
rect 5700 3425 5800 3440
rect 5700 3325 5705 3425
rect 5740 3325 5760 3425
rect 5795 3325 5800 3425
rect 5700 3310 5800 3325
rect 5950 3425 6050 3440
rect 5950 3325 5955 3425
rect 5990 3325 6010 3425
rect 6045 3325 6050 3425
rect 5950 3310 6050 3325
rect 6200 3425 6300 3440
rect 6200 3325 6205 3425
rect 6240 3325 6260 3425
rect 6295 3325 6300 3425
rect 6200 3310 6300 3325
rect 6450 3425 6550 3440
rect 6450 3325 6455 3425
rect 6490 3325 6510 3425
rect 6545 3325 6550 3425
rect 6450 3310 6550 3325
rect 6700 3425 6800 3440
rect 6700 3325 6705 3425
rect 6740 3325 6760 3425
rect 6795 3325 6800 3425
rect 6700 3310 6800 3325
rect 6950 3425 7050 3440
rect 6950 3325 6955 3425
rect 6990 3325 7010 3425
rect 7045 3325 7050 3425
rect 6950 3310 7050 3325
rect 7200 3425 7300 3440
rect 7200 3325 7205 3425
rect 7240 3325 7260 3425
rect 7295 3325 7300 3425
rect 7200 3310 7300 3325
rect 7450 3425 7550 3440
rect 7450 3325 7455 3425
rect 7490 3325 7510 3425
rect 7545 3325 7550 3425
rect 7450 3310 7550 3325
rect 7700 3425 7800 3440
rect 7700 3325 7705 3425
rect 7740 3325 7760 3425
rect 7795 3325 7800 3425
rect 7700 3310 7800 3325
rect 7950 3425 8000 3440
rect 7950 3325 7955 3425
rect 7990 3325 8000 3425
rect 7950 3310 8000 3325
rect 0 3300 60 3310
rect 190 3300 310 3310
rect 440 3300 560 3310
rect 690 3300 810 3310
rect 940 3300 1060 3310
rect 1190 3300 1310 3310
rect 1440 3300 1560 3310
rect 1690 3300 1810 3310
rect 1940 3300 2060 3310
rect 2190 3300 2310 3310
rect 2440 3300 2560 3310
rect 2690 3300 2810 3310
rect 2940 3300 3060 3310
rect 3190 3300 3310 3310
rect 3440 3300 3560 3310
rect 3690 3300 3810 3310
rect 3940 3300 4060 3310
rect 4190 3300 4310 3310
rect 4440 3300 4560 3310
rect 4690 3300 4810 3310
rect 4940 3300 5060 3310
rect 5190 3300 5310 3310
rect 5440 3300 5560 3310
rect 5690 3300 5810 3310
rect 5940 3300 6060 3310
rect 6190 3300 6310 3310
rect 6440 3300 6560 3310
rect 6690 3300 6810 3310
rect 6940 3300 7060 3310
rect 7190 3300 7310 3310
rect 7440 3300 7560 3310
rect 7690 3300 7810 3310
rect 7940 3300 8000 3310
rect 0 3295 8000 3300
rect 0 3260 75 3295
rect 175 3260 325 3295
rect 425 3260 575 3295
rect 675 3260 825 3295
rect 925 3260 1075 3295
rect 1175 3260 1325 3295
rect 1425 3260 1575 3295
rect 1675 3260 1825 3295
rect 1925 3260 2075 3295
rect 2175 3260 2325 3295
rect 2425 3260 2575 3295
rect 2675 3260 2825 3295
rect 2925 3260 3075 3295
rect 3175 3260 3325 3295
rect 3425 3260 3575 3295
rect 3675 3260 3825 3295
rect 3925 3260 4075 3295
rect 4175 3260 4325 3295
rect 4425 3260 4575 3295
rect 4675 3260 4825 3295
rect 4925 3260 5075 3295
rect 5175 3260 5325 3295
rect 5425 3260 5575 3295
rect 5675 3260 5825 3295
rect 5925 3260 6075 3295
rect 6175 3260 6325 3295
rect 6425 3260 6575 3295
rect 6675 3260 6825 3295
rect 6925 3260 7075 3295
rect 7175 3260 7325 3295
rect 7425 3260 7575 3295
rect 7675 3260 7825 3295
rect 7925 3260 8000 3295
rect 0 3240 8000 3260
rect 0 3205 75 3240
rect 175 3205 325 3240
rect 425 3205 575 3240
rect 675 3205 825 3240
rect 925 3205 1075 3240
rect 1175 3205 1325 3240
rect 1425 3205 1575 3240
rect 1675 3205 1825 3240
rect 1925 3205 2075 3240
rect 2175 3205 2325 3240
rect 2425 3205 2575 3240
rect 2675 3205 2825 3240
rect 2925 3205 3075 3240
rect 3175 3205 3325 3240
rect 3425 3205 3575 3240
rect 3675 3205 3825 3240
rect 3925 3205 4075 3240
rect 4175 3205 4325 3240
rect 4425 3205 4575 3240
rect 4675 3205 4825 3240
rect 4925 3205 5075 3240
rect 5175 3205 5325 3240
rect 5425 3205 5575 3240
rect 5675 3205 5825 3240
rect 5925 3205 6075 3240
rect 6175 3205 6325 3240
rect 6425 3205 6575 3240
rect 6675 3205 6825 3240
rect 6925 3205 7075 3240
rect 7175 3205 7325 3240
rect 7425 3205 7575 3240
rect 7675 3205 7825 3240
rect 7925 3205 8000 3240
rect 0 3200 8000 3205
rect 0 3190 60 3200
rect 190 3190 310 3200
rect 440 3190 560 3200
rect 690 3190 810 3200
rect 940 3190 1060 3200
rect 1190 3190 1310 3200
rect 1440 3190 1560 3200
rect 1690 3190 1810 3200
rect 1940 3190 2060 3200
rect 2190 3190 2310 3200
rect 2440 3190 2560 3200
rect 2690 3190 2810 3200
rect 2940 3190 3060 3200
rect 3190 3190 3310 3200
rect 3440 3190 3560 3200
rect 3690 3190 3810 3200
rect 3940 3190 4060 3200
rect 4190 3190 4310 3200
rect 4440 3190 4560 3200
rect 4690 3190 4810 3200
rect 4940 3190 5060 3200
rect 5190 3190 5310 3200
rect 5440 3190 5560 3200
rect 5690 3190 5810 3200
rect 5940 3190 6060 3200
rect 6190 3190 6310 3200
rect 6440 3190 6560 3200
rect 6690 3190 6810 3200
rect 6940 3190 7060 3200
rect 7190 3190 7310 3200
rect 7440 3190 7560 3200
rect 7690 3190 7810 3200
rect 7940 3190 8000 3200
rect 0 3175 50 3190
rect 0 3075 10 3175
rect 45 3075 50 3175
rect 0 3060 50 3075
rect 200 3175 300 3190
rect 200 3075 205 3175
rect 240 3075 260 3175
rect 295 3075 300 3175
rect 200 3060 300 3075
rect 450 3175 550 3190
rect 450 3075 455 3175
rect 490 3075 510 3175
rect 545 3075 550 3175
rect 450 3060 550 3075
rect 700 3175 800 3190
rect 700 3075 705 3175
rect 740 3075 760 3175
rect 795 3075 800 3175
rect 700 3060 800 3075
rect 950 3175 1050 3190
rect 950 3075 955 3175
rect 990 3075 1010 3175
rect 1045 3075 1050 3175
rect 950 3060 1050 3075
rect 1200 3175 1300 3190
rect 1200 3075 1205 3175
rect 1240 3075 1260 3175
rect 1295 3075 1300 3175
rect 1200 3060 1300 3075
rect 1450 3175 1550 3190
rect 1450 3075 1455 3175
rect 1490 3075 1510 3175
rect 1545 3075 1550 3175
rect 1450 3060 1550 3075
rect 1700 3175 1800 3190
rect 1700 3075 1705 3175
rect 1740 3075 1760 3175
rect 1795 3075 1800 3175
rect 1700 3060 1800 3075
rect 1950 3175 2050 3190
rect 1950 3075 1955 3175
rect 1990 3075 2010 3175
rect 2045 3075 2050 3175
rect 1950 3060 2050 3075
rect 2200 3175 2300 3190
rect 2200 3075 2205 3175
rect 2240 3075 2260 3175
rect 2295 3075 2300 3175
rect 2200 3060 2300 3075
rect 2450 3175 2550 3190
rect 2450 3075 2455 3175
rect 2490 3075 2510 3175
rect 2545 3075 2550 3175
rect 2450 3060 2550 3075
rect 2700 3175 2800 3190
rect 2700 3075 2705 3175
rect 2740 3075 2760 3175
rect 2795 3075 2800 3175
rect 2700 3060 2800 3075
rect 2950 3175 3050 3190
rect 2950 3075 2955 3175
rect 2990 3075 3010 3175
rect 3045 3075 3050 3175
rect 2950 3060 3050 3075
rect 3200 3175 3300 3190
rect 3200 3075 3205 3175
rect 3240 3075 3260 3175
rect 3295 3075 3300 3175
rect 3200 3060 3300 3075
rect 3450 3175 3550 3190
rect 3450 3075 3455 3175
rect 3490 3075 3510 3175
rect 3545 3075 3550 3175
rect 3450 3060 3550 3075
rect 3700 3175 3800 3190
rect 3700 3075 3705 3175
rect 3740 3075 3760 3175
rect 3795 3075 3800 3175
rect 3700 3060 3800 3075
rect 3950 3175 4050 3190
rect 3950 3075 3955 3175
rect 3990 3075 4010 3175
rect 4045 3075 4050 3175
rect 3950 3060 4050 3075
rect 4200 3175 4300 3190
rect 4200 3075 4205 3175
rect 4240 3075 4260 3175
rect 4295 3075 4300 3175
rect 4200 3060 4300 3075
rect 4450 3175 4550 3190
rect 4450 3075 4455 3175
rect 4490 3075 4510 3175
rect 4545 3075 4550 3175
rect 4450 3060 4550 3075
rect 4700 3175 4800 3190
rect 4700 3075 4705 3175
rect 4740 3075 4760 3175
rect 4795 3075 4800 3175
rect 4700 3060 4800 3075
rect 4950 3175 5050 3190
rect 4950 3075 4955 3175
rect 4990 3075 5010 3175
rect 5045 3075 5050 3175
rect 4950 3060 5050 3075
rect 5200 3175 5300 3190
rect 5200 3075 5205 3175
rect 5240 3075 5260 3175
rect 5295 3075 5300 3175
rect 5200 3060 5300 3075
rect 5450 3175 5550 3190
rect 5450 3075 5455 3175
rect 5490 3075 5510 3175
rect 5545 3075 5550 3175
rect 5450 3060 5550 3075
rect 5700 3175 5800 3190
rect 5700 3075 5705 3175
rect 5740 3075 5760 3175
rect 5795 3075 5800 3175
rect 5700 3060 5800 3075
rect 5950 3175 6050 3190
rect 5950 3075 5955 3175
rect 5990 3075 6010 3175
rect 6045 3075 6050 3175
rect 5950 3060 6050 3075
rect 6200 3175 6300 3190
rect 6200 3075 6205 3175
rect 6240 3075 6260 3175
rect 6295 3075 6300 3175
rect 6200 3060 6300 3075
rect 6450 3175 6550 3190
rect 6450 3075 6455 3175
rect 6490 3075 6510 3175
rect 6545 3075 6550 3175
rect 6450 3060 6550 3075
rect 6700 3175 6800 3190
rect 6700 3075 6705 3175
rect 6740 3075 6760 3175
rect 6795 3075 6800 3175
rect 6700 3060 6800 3075
rect 6950 3175 7050 3190
rect 6950 3075 6955 3175
rect 6990 3075 7010 3175
rect 7045 3075 7050 3175
rect 6950 3060 7050 3075
rect 7200 3175 7300 3190
rect 7200 3075 7205 3175
rect 7240 3075 7260 3175
rect 7295 3075 7300 3175
rect 7200 3060 7300 3075
rect 7450 3175 7550 3190
rect 7450 3075 7455 3175
rect 7490 3075 7510 3175
rect 7545 3075 7550 3175
rect 7450 3060 7550 3075
rect 7700 3175 7800 3190
rect 7700 3075 7705 3175
rect 7740 3075 7760 3175
rect 7795 3075 7800 3175
rect 7700 3060 7800 3075
rect 7950 3175 8000 3190
rect 7950 3075 7955 3175
rect 7990 3075 8000 3175
rect 7950 3060 8000 3075
rect 0 3050 60 3060
rect 190 3050 310 3060
rect 440 3050 560 3060
rect 690 3050 810 3060
rect 940 3050 1060 3060
rect 1190 3050 1310 3060
rect 1440 3050 1560 3060
rect 1690 3050 1810 3060
rect 1940 3050 2060 3060
rect 2190 3050 2310 3060
rect 2440 3050 2560 3060
rect 2690 3050 2810 3060
rect 2940 3050 3060 3060
rect 3190 3050 3310 3060
rect 3440 3050 3560 3060
rect 3690 3050 3810 3060
rect 3940 3050 4060 3060
rect 4190 3050 4310 3060
rect 4440 3050 4560 3060
rect 4690 3050 4810 3060
rect 4940 3050 5060 3060
rect 5190 3050 5310 3060
rect 5440 3050 5560 3060
rect 5690 3050 5810 3060
rect 5940 3050 6060 3060
rect 6190 3050 6310 3060
rect 6440 3050 6560 3060
rect 6690 3050 6810 3060
rect 6940 3050 7060 3060
rect 7190 3050 7310 3060
rect 7440 3050 7560 3060
rect 7690 3050 7810 3060
rect 7940 3050 8000 3060
rect 0 3045 8000 3050
rect 0 3010 75 3045
rect 175 3010 325 3045
rect 425 3010 575 3045
rect 675 3010 825 3045
rect 925 3010 1075 3045
rect 1175 3010 1325 3045
rect 1425 3010 1575 3045
rect 1675 3010 1825 3045
rect 1925 3010 2075 3045
rect 2175 3010 2325 3045
rect 2425 3010 2575 3045
rect 2675 3010 2825 3045
rect 2925 3010 3075 3045
rect 3175 3010 3325 3045
rect 3425 3010 3575 3045
rect 3675 3010 3825 3045
rect 3925 3010 4075 3045
rect 4175 3010 4325 3045
rect 4425 3010 4575 3045
rect 4675 3010 4825 3045
rect 4925 3010 5075 3045
rect 5175 3010 5325 3045
rect 5425 3010 5575 3045
rect 5675 3010 5825 3045
rect 5925 3010 6075 3045
rect 6175 3010 6325 3045
rect 6425 3010 6575 3045
rect 6675 3010 6825 3045
rect 6925 3010 7075 3045
rect 7175 3010 7325 3045
rect 7425 3010 7575 3045
rect 7675 3010 7825 3045
rect 7925 3010 8000 3045
rect 0 2990 8000 3010
rect 0 2955 75 2990
rect 175 2955 325 2990
rect 425 2955 575 2990
rect 675 2955 825 2990
rect 925 2955 1075 2990
rect 1175 2955 1325 2990
rect 1425 2955 1575 2990
rect 1675 2955 1825 2990
rect 1925 2955 2075 2990
rect 2175 2955 2325 2990
rect 2425 2955 2575 2990
rect 2675 2955 2825 2990
rect 2925 2955 3075 2990
rect 3175 2955 3325 2990
rect 3425 2955 3575 2990
rect 3675 2955 3825 2990
rect 3925 2955 4075 2990
rect 4175 2955 4325 2990
rect 4425 2955 4575 2990
rect 4675 2955 4825 2990
rect 4925 2955 5075 2990
rect 5175 2955 5325 2990
rect 5425 2955 5575 2990
rect 5675 2955 5825 2990
rect 5925 2955 6075 2990
rect 6175 2955 6325 2990
rect 6425 2955 6575 2990
rect 6675 2955 6825 2990
rect 6925 2955 7075 2990
rect 7175 2955 7325 2990
rect 7425 2955 7575 2990
rect 7675 2955 7825 2990
rect 7925 2955 8000 2990
rect 0 2950 8000 2955
rect 0 2940 60 2950
rect 190 2940 310 2950
rect 440 2940 560 2950
rect 690 2940 810 2950
rect 940 2940 1060 2950
rect 1190 2940 1310 2950
rect 1440 2940 1560 2950
rect 1690 2940 1810 2950
rect 1940 2940 2060 2950
rect 2190 2940 2310 2950
rect 2440 2940 2560 2950
rect 2690 2940 2810 2950
rect 2940 2940 3060 2950
rect 3190 2940 3310 2950
rect 3440 2940 3560 2950
rect 3690 2940 3810 2950
rect 3940 2940 4060 2950
rect 4190 2940 4310 2950
rect 4440 2940 4560 2950
rect 4690 2940 4810 2950
rect 4940 2940 5060 2950
rect 5190 2940 5310 2950
rect 5440 2940 5560 2950
rect 5690 2940 5810 2950
rect 5940 2940 6060 2950
rect 6190 2940 6310 2950
rect 6440 2940 6560 2950
rect 6690 2940 6810 2950
rect 6940 2940 7060 2950
rect 7190 2940 7310 2950
rect 7440 2940 7560 2950
rect 7690 2940 7810 2950
rect 7940 2940 8000 2950
rect 0 2925 50 2940
rect 0 2825 10 2925
rect 45 2825 50 2925
rect 0 2810 50 2825
rect 200 2925 300 2940
rect 200 2825 205 2925
rect 240 2825 260 2925
rect 295 2825 300 2925
rect 200 2810 300 2825
rect 450 2925 550 2940
rect 450 2825 455 2925
rect 490 2825 510 2925
rect 545 2825 550 2925
rect 450 2810 550 2825
rect 700 2925 800 2940
rect 700 2825 705 2925
rect 740 2825 760 2925
rect 795 2825 800 2925
rect 700 2810 800 2825
rect 950 2925 1050 2940
rect 950 2825 955 2925
rect 990 2825 1010 2925
rect 1045 2825 1050 2925
rect 950 2810 1050 2825
rect 1200 2925 1300 2940
rect 1200 2825 1205 2925
rect 1240 2825 1260 2925
rect 1295 2825 1300 2925
rect 1200 2810 1300 2825
rect 1450 2925 1550 2940
rect 1450 2825 1455 2925
rect 1490 2825 1510 2925
rect 1545 2825 1550 2925
rect 1450 2810 1550 2825
rect 1700 2925 1800 2940
rect 1700 2825 1705 2925
rect 1740 2825 1760 2925
rect 1795 2825 1800 2925
rect 1700 2810 1800 2825
rect 1950 2925 2050 2940
rect 1950 2825 1955 2925
rect 1990 2825 2010 2925
rect 2045 2825 2050 2925
rect 1950 2810 2050 2825
rect 2200 2925 2300 2940
rect 2200 2825 2205 2925
rect 2240 2825 2260 2925
rect 2295 2825 2300 2925
rect 2200 2810 2300 2825
rect 2450 2925 2550 2940
rect 2450 2825 2455 2925
rect 2490 2825 2510 2925
rect 2545 2825 2550 2925
rect 2450 2810 2550 2825
rect 2700 2925 2800 2940
rect 2700 2825 2705 2925
rect 2740 2825 2760 2925
rect 2795 2825 2800 2925
rect 2700 2810 2800 2825
rect 2950 2925 3050 2940
rect 2950 2825 2955 2925
rect 2990 2825 3010 2925
rect 3045 2825 3050 2925
rect 2950 2810 3050 2825
rect 3200 2925 3300 2940
rect 3200 2825 3205 2925
rect 3240 2825 3260 2925
rect 3295 2825 3300 2925
rect 3200 2810 3300 2825
rect 3450 2925 3550 2940
rect 3450 2825 3455 2925
rect 3490 2825 3510 2925
rect 3545 2825 3550 2925
rect 3450 2810 3550 2825
rect 3700 2925 3800 2940
rect 3700 2825 3705 2925
rect 3740 2825 3760 2925
rect 3795 2825 3800 2925
rect 3700 2810 3800 2825
rect 3950 2925 4050 2940
rect 3950 2825 3955 2925
rect 3990 2825 4010 2925
rect 4045 2825 4050 2925
rect 3950 2810 4050 2825
rect 4200 2925 4300 2940
rect 4200 2825 4205 2925
rect 4240 2825 4260 2925
rect 4295 2825 4300 2925
rect 4200 2810 4300 2825
rect 4450 2925 4550 2940
rect 4450 2825 4455 2925
rect 4490 2825 4510 2925
rect 4545 2825 4550 2925
rect 4450 2810 4550 2825
rect 4700 2925 4800 2940
rect 4700 2825 4705 2925
rect 4740 2825 4760 2925
rect 4795 2825 4800 2925
rect 4700 2810 4800 2825
rect 4950 2925 5050 2940
rect 4950 2825 4955 2925
rect 4990 2825 5010 2925
rect 5045 2825 5050 2925
rect 4950 2810 5050 2825
rect 5200 2925 5300 2940
rect 5200 2825 5205 2925
rect 5240 2825 5260 2925
rect 5295 2825 5300 2925
rect 5200 2810 5300 2825
rect 5450 2925 5550 2940
rect 5450 2825 5455 2925
rect 5490 2825 5510 2925
rect 5545 2825 5550 2925
rect 5450 2810 5550 2825
rect 5700 2925 5800 2940
rect 5700 2825 5705 2925
rect 5740 2825 5760 2925
rect 5795 2825 5800 2925
rect 5700 2810 5800 2825
rect 5950 2925 6050 2940
rect 5950 2825 5955 2925
rect 5990 2825 6010 2925
rect 6045 2825 6050 2925
rect 5950 2810 6050 2825
rect 6200 2925 6300 2940
rect 6200 2825 6205 2925
rect 6240 2825 6260 2925
rect 6295 2825 6300 2925
rect 6200 2810 6300 2825
rect 6450 2925 6550 2940
rect 6450 2825 6455 2925
rect 6490 2825 6510 2925
rect 6545 2825 6550 2925
rect 6450 2810 6550 2825
rect 6700 2925 6800 2940
rect 6700 2825 6705 2925
rect 6740 2825 6760 2925
rect 6795 2825 6800 2925
rect 6700 2810 6800 2825
rect 6950 2925 7050 2940
rect 6950 2825 6955 2925
rect 6990 2825 7010 2925
rect 7045 2825 7050 2925
rect 6950 2810 7050 2825
rect 7200 2925 7300 2940
rect 7200 2825 7205 2925
rect 7240 2825 7260 2925
rect 7295 2825 7300 2925
rect 7200 2810 7300 2825
rect 7450 2925 7550 2940
rect 7450 2825 7455 2925
rect 7490 2825 7510 2925
rect 7545 2825 7550 2925
rect 7450 2810 7550 2825
rect 7700 2925 7800 2940
rect 7700 2825 7705 2925
rect 7740 2825 7760 2925
rect 7795 2825 7800 2925
rect 7700 2810 7800 2825
rect 7950 2925 8000 2940
rect 7950 2825 7955 2925
rect 7990 2825 8000 2925
rect 7950 2810 8000 2825
rect 0 2800 60 2810
rect 190 2800 310 2810
rect 440 2800 560 2810
rect 690 2800 810 2810
rect 940 2800 1060 2810
rect 1190 2800 1310 2810
rect 1440 2800 1560 2810
rect 1690 2800 1810 2810
rect 1940 2800 2060 2810
rect 2190 2800 2310 2810
rect 2440 2800 2560 2810
rect 2690 2800 2810 2810
rect 2940 2800 3060 2810
rect 3190 2800 3310 2810
rect 3440 2800 3560 2810
rect 3690 2800 3810 2810
rect 3940 2800 4060 2810
rect 4190 2800 4310 2810
rect 4440 2800 4560 2810
rect 4690 2800 4810 2810
rect 4940 2800 5060 2810
rect 5190 2800 5310 2810
rect 5440 2800 5560 2810
rect 5690 2800 5810 2810
rect 5940 2800 6060 2810
rect 6190 2800 6310 2810
rect 6440 2800 6560 2810
rect 6690 2800 6810 2810
rect 6940 2800 7060 2810
rect 7190 2800 7310 2810
rect 7440 2800 7560 2810
rect 7690 2800 7810 2810
rect 7940 2800 8000 2810
rect 0 2795 8000 2800
rect 0 2760 75 2795
rect 175 2760 325 2795
rect 425 2760 575 2795
rect 675 2760 825 2795
rect 925 2760 1075 2795
rect 1175 2760 1325 2795
rect 1425 2760 1575 2795
rect 1675 2760 1825 2795
rect 1925 2760 2075 2795
rect 2175 2760 2325 2795
rect 2425 2760 2575 2795
rect 2675 2760 2825 2795
rect 2925 2760 3075 2795
rect 3175 2760 3325 2795
rect 3425 2760 3575 2795
rect 3675 2760 3825 2795
rect 3925 2760 4075 2795
rect 4175 2760 4325 2795
rect 4425 2760 4575 2795
rect 4675 2760 4825 2795
rect 4925 2760 5075 2795
rect 5175 2760 5325 2795
rect 5425 2760 5575 2795
rect 5675 2760 5825 2795
rect 5925 2760 6075 2795
rect 6175 2760 6325 2795
rect 6425 2760 6575 2795
rect 6675 2760 6825 2795
rect 6925 2760 7075 2795
rect 7175 2760 7325 2795
rect 7425 2760 7575 2795
rect 7675 2760 7825 2795
rect 7925 2760 8000 2795
rect 0 2740 8000 2760
rect 0 2705 75 2740
rect 175 2705 325 2740
rect 425 2705 575 2740
rect 675 2705 825 2740
rect 925 2705 1075 2740
rect 1175 2705 1325 2740
rect 1425 2705 1575 2740
rect 1675 2705 1825 2740
rect 1925 2705 2075 2740
rect 2175 2705 2325 2740
rect 2425 2705 2575 2740
rect 2675 2705 2825 2740
rect 2925 2705 3075 2740
rect 3175 2705 3325 2740
rect 3425 2705 3575 2740
rect 3675 2705 3825 2740
rect 3925 2705 4075 2740
rect 4175 2705 4325 2740
rect 4425 2705 4575 2740
rect 4675 2705 4825 2740
rect 4925 2705 5075 2740
rect 5175 2705 5325 2740
rect 5425 2705 5575 2740
rect 5675 2705 5825 2740
rect 5925 2705 6075 2740
rect 6175 2705 6325 2740
rect 6425 2705 6575 2740
rect 6675 2705 6825 2740
rect 6925 2705 7075 2740
rect 7175 2705 7325 2740
rect 7425 2705 7575 2740
rect 7675 2705 7825 2740
rect 7925 2705 8000 2740
rect 0 2700 8000 2705
rect 0 2690 60 2700
rect 190 2690 310 2700
rect 440 2690 560 2700
rect 690 2690 810 2700
rect 940 2690 1060 2700
rect 1190 2690 1310 2700
rect 1440 2690 1560 2700
rect 1690 2690 1810 2700
rect 1940 2690 2060 2700
rect 2190 2690 2310 2700
rect 2440 2690 2560 2700
rect 2690 2690 2810 2700
rect 2940 2690 3060 2700
rect 3190 2690 3310 2700
rect 3440 2690 3560 2700
rect 3690 2690 3810 2700
rect 3940 2690 4060 2700
rect 4190 2690 4310 2700
rect 4440 2690 4560 2700
rect 4690 2690 4810 2700
rect 4940 2690 5060 2700
rect 5190 2690 5310 2700
rect 5440 2690 5560 2700
rect 5690 2690 5810 2700
rect 5940 2690 6060 2700
rect 6190 2690 6310 2700
rect 6440 2690 6560 2700
rect 6690 2690 6810 2700
rect 6940 2690 7060 2700
rect 7190 2690 7310 2700
rect 7440 2690 7560 2700
rect 7690 2690 7810 2700
rect 7940 2690 8000 2700
rect 0 2675 50 2690
rect 0 2575 10 2675
rect 45 2575 50 2675
rect 0 2560 50 2575
rect 200 2675 300 2690
rect 200 2575 205 2675
rect 240 2575 260 2675
rect 295 2575 300 2675
rect 200 2560 300 2575
rect 450 2675 550 2690
rect 450 2575 455 2675
rect 490 2575 510 2675
rect 545 2575 550 2675
rect 450 2560 550 2575
rect 700 2675 800 2690
rect 700 2575 705 2675
rect 740 2575 760 2675
rect 795 2575 800 2675
rect 700 2560 800 2575
rect 950 2675 1050 2690
rect 950 2575 955 2675
rect 990 2575 1010 2675
rect 1045 2575 1050 2675
rect 950 2560 1050 2575
rect 1200 2675 1300 2690
rect 1200 2575 1205 2675
rect 1240 2575 1260 2675
rect 1295 2575 1300 2675
rect 1200 2560 1300 2575
rect 1450 2675 1550 2690
rect 1450 2575 1455 2675
rect 1490 2575 1510 2675
rect 1545 2575 1550 2675
rect 1450 2560 1550 2575
rect 1700 2675 1800 2690
rect 1700 2575 1705 2675
rect 1740 2575 1760 2675
rect 1795 2575 1800 2675
rect 1700 2560 1800 2575
rect 1950 2675 2050 2690
rect 1950 2575 1955 2675
rect 1990 2575 2010 2675
rect 2045 2575 2050 2675
rect 1950 2560 2050 2575
rect 2200 2675 2300 2690
rect 2200 2575 2205 2675
rect 2240 2575 2260 2675
rect 2295 2575 2300 2675
rect 2200 2560 2300 2575
rect 2450 2675 2550 2690
rect 2450 2575 2455 2675
rect 2490 2575 2510 2675
rect 2545 2575 2550 2675
rect 2450 2560 2550 2575
rect 2700 2675 2800 2690
rect 2700 2575 2705 2675
rect 2740 2575 2760 2675
rect 2795 2575 2800 2675
rect 2700 2560 2800 2575
rect 2950 2675 3050 2690
rect 2950 2575 2955 2675
rect 2990 2575 3010 2675
rect 3045 2575 3050 2675
rect 2950 2560 3050 2575
rect 3200 2675 3300 2690
rect 3200 2575 3205 2675
rect 3240 2575 3260 2675
rect 3295 2575 3300 2675
rect 3200 2560 3300 2575
rect 3450 2675 3550 2690
rect 3450 2575 3455 2675
rect 3490 2575 3510 2675
rect 3545 2575 3550 2675
rect 3450 2560 3550 2575
rect 3700 2675 3800 2690
rect 3700 2575 3705 2675
rect 3740 2575 3760 2675
rect 3795 2575 3800 2675
rect 3700 2560 3800 2575
rect 3950 2675 4050 2690
rect 3950 2575 3955 2675
rect 3990 2575 4010 2675
rect 4045 2575 4050 2675
rect 3950 2560 4050 2575
rect 4200 2675 4300 2690
rect 4200 2575 4205 2675
rect 4240 2575 4260 2675
rect 4295 2575 4300 2675
rect 4200 2560 4300 2575
rect 4450 2675 4550 2690
rect 4450 2575 4455 2675
rect 4490 2575 4510 2675
rect 4545 2575 4550 2675
rect 4450 2560 4550 2575
rect 4700 2675 4800 2690
rect 4700 2575 4705 2675
rect 4740 2575 4760 2675
rect 4795 2575 4800 2675
rect 4700 2560 4800 2575
rect 4950 2675 5050 2690
rect 4950 2575 4955 2675
rect 4990 2575 5010 2675
rect 5045 2575 5050 2675
rect 4950 2560 5050 2575
rect 5200 2675 5300 2690
rect 5200 2575 5205 2675
rect 5240 2575 5260 2675
rect 5295 2575 5300 2675
rect 5200 2560 5300 2575
rect 5450 2675 5550 2690
rect 5450 2575 5455 2675
rect 5490 2575 5510 2675
rect 5545 2575 5550 2675
rect 5450 2560 5550 2575
rect 5700 2675 5800 2690
rect 5700 2575 5705 2675
rect 5740 2575 5760 2675
rect 5795 2575 5800 2675
rect 5700 2560 5800 2575
rect 5950 2675 6050 2690
rect 5950 2575 5955 2675
rect 5990 2575 6010 2675
rect 6045 2575 6050 2675
rect 5950 2560 6050 2575
rect 6200 2675 6300 2690
rect 6200 2575 6205 2675
rect 6240 2575 6260 2675
rect 6295 2575 6300 2675
rect 6200 2560 6300 2575
rect 6450 2675 6550 2690
rect 6450 2575 6455 2675
rect 6490 2575 6510 2675
rect 6545 2575 6550 2675
rect 6450 2560 6550 2575
rect 6700 2675 6800 2690
rect 6700 2575 6705 2675
rect 6740 2575 6760 2675
rect 6795 2575 6800 2675
rect 6700 2560 6800 2575
rect 6950 2675 7050 2690
rect 6950 2575 6955 2675
rect 6990 2575 7010 2675
rect 7045 2575 7050 2675
rect 6950 2560 7050 2575
rect 7200 2675 7300 2690
rect 7200 2575 7205 2675
rect 7240 2575 7260 2675
rect 7295 2575 7300 2675
rect 7200 2560 7300 2575
rect 7450 2675 7550 2690
rect 7450 2575 7455 2675
rect 7490 2575 7510 2675
rect 7545 2575 7550 2675
rect 7450 2560 7550 2575
rect 7700 2675 7800 2690
rect 7700 2575 7705 2675
rect 7740 2575 7760 2675
rect 7795 2575 7800 2675
rect 7700 2560 7800 2575
rect 7950 2675 8000 2690
rect 7950 2575 7955 2675
rect 7990 2575 8000 2675
rect 7950 2560 8000 2575
rect 0 2550 60 2560
rect 190 2550 310 2560
rect 440 2550 560 2560
rect 690 2550 810 2560
rect 940 2550 1060 2560
rect 1190 2550 1310 2560
rect 1440 2550 1560 2560
rect 1690 2550 1810 2560
rect 1940 2550 2060 2560
rect 2190 2550 2310 2560
rect 2440 2550 2560 2560
rect 2690 2550 2810 2560
rect 2940 2550 3060 2560
rect 3190 2550 3310 2560
rect 3440 2550 3560 2560
rect 3690 2550 3810 2560
rect 3940 2550 4060 2560
rect 4190 2550 4310 2560
rect 4440 2550 4560 2560
rect 4690 2550 4810 2560
rect 4940 2550 5060 2560
rect 5190 2550 5310 2560
rect 5440 2550 5560 2560
rect 5690 2550 5810 2560
rect 5940 2550 6060 2560
rect 6190 2550 6310 2560
rect 6440 2550 6560 2560
rect 6690 2550 6810 2560
rect 6940 2550 7060 2560
rect 7190 2550 7310 2560
rect 7440 2550 7560 2560
rect 7690 2550 7810 2560
rect 7940 2550 8000 2560
rect 0 2545 8000 2550
rect 0 2510 75 2545
rect 175 2510 325 2545
rect 425 2510 575 2545
rect 675 2510 825 2545
rect 925 2510 1075 2545
rect 1175 2510 1325 2545
rect 1425 2510 1575 2545
rect 1675 2510 1825 2545
rect 1925 2510 2075 2545
rect 2175 2510 2325 2545
rect 2425 2510 2575 2545
rect 2675 2510 2825 2545
rect 2925 2510 3075 2545
rect 3175 2510 3325 2545
rect 3425 2510 3575 2545
rect 3675 2510 3825 2545
rect 3925 2510 4075 2545
rect 4175 2510 4325 2545
rect 4425 2510 4575 2545
rect 4675 2510 4825 2545
rect 4925 2510 5075 2545
rect 5175 2510 5325 2545
rect 5425 2510 5575 2545
rect 5675 2510 5825 2545
rect 5925 2510 6075 2545
rect 6175 2510 6325 2545
rect 6425 2510 6575 2545
rect 6675 2510 6825 2545
rect 6925 2510 7075 2545
rect 7175 2510 7325 2545
rect 7425 2510 7575 2545
rect 7675 2510 7825 2545
rect 7925 2510 8000 2545
rect 0 2490 8000 2510
rect 0 2455 75 2490
rect 175 2455 325 2490
rect 425 2455 575 2490
rect 675 2455 825 2490
rect 925 2455 1075 2490
rect 1175 2455 1325 2490
rect 1425 2455 1575 2490
rect 1675 2455 1825 2490
rect 1925 2455 2075 2490
rect 2175 2455 2325 2490
rect 2425 2455 2575 2490
rect 2675 2455 2825 2490
rect 2925 2455 3075 2490
rect 3175 2455 3325 2490
rect 3425 2455 3575 2490
rect 3675 2455 3825 2490
rect 3925 2455 4075 2490
rect 4175 2455 4325 2490
rect 4425 2455 4575 2490
rect 4675 2455 4825 2490
rect 4925 2455 5075 2490
rect 5175 2455 5325 2490
rect 5425 2455 5575 2490
rect 5675 2455 5825 2490
rect 5925 2455 6075 2490
rect 6175 2455 6325 2490
rect 6425 2455 6575 2490
rect 6675 2455 6825 2490
rect 6925 2455 7075 2490
rect 7175 2455 7325 2490
rect 7425 2455 7575 2490
rect 7675 2455 7825 2490
rect 7925 2455 8000 2490
rect 0 2450 8000 2455
rect 0 2440 60 2450
rect 190 2440 310 2450
rect 440 2440 560 2450
rect 690 2440 810 2450
rect 940 2440 1060 2450
rect 1190 2440 1310 2450
rect 1440 2440 1560 2450
rect 1690 2440 1810 2450
rect 1940 2440 2060 2450
rect 2190 2440 2310 2450
rect 2440 2440 2560 2450
rect 2690 2440 2810 2450
rect 2940 2440 3060 2450
rect 3190 2440 3310 2450
rect 3440 2440 3560 2450
rect 3690 2440 3810 2450
rect 3940 2440 4060 2450
rect 4190 2440 4310 2450
rect 4440 2440 4560 2450
rect 4690 2440 4810 2450
rect 4940 2440 5060 2450
rect 5190 2440 5310 2450
rect 5440 2440 5560 2450
rect 5690 2440 5810 2450
rect 5940 2440 6060 2450
rect 6190 2440 6310 2450
rect 6440 2440 6560 2450
rect 6690 2440 6810 2450
rect 6940 2440 7060 2450
rect 7190 2440 7310 2450
rect 7440 2440 7560 2450
rect 7690 2440 7810 2450
rect 7940 2440 8000 2450
rect 0 2425 50 2440
rect 0 2325 10 2425
rect 45 2325 50 2425
rect 0 2310 50 2325
rect 200 2425 300 2440
rect 200 2325 205 2425
rect 240 2325 260 2425
rect 295 2325 300 2425
rect 200 2310 300 2325
rect 450 2425 550 2440
rect 450 2325 455 2425
rect 490 2325 510 2425
rect 545 2325 550 2425
rect 450 2310 550 2325
rect 700 2425 800 2440
rect 700 2325 705 2425
rect 740 2325 760 2425
rect 795 2325 800 2425
rect 700 2310 800 2325
rect 950 2425 1050 2440
rect 950 2325 955 2425
rect 990 2325 1010 2425
rect 1045 2325 1050 2425
rect 950 2310 1050 2325
rect 1200 2425 1300 2440
rect 1200 2325 1205 2425
rect 1240 2325 1260 2425
rect 1295 2325 1300 2425
rect 1200 2310 1300 2325
rect 1450 2425 1550 2440
rect 1450 2325 1455 2425
rect 1490 2325 1510 2425
rect 1545 2325 1550 2425
rect 1450 2310 1550 2325
rect 1700 2425 1800 2440
rect 1700 2325 1705 2425
rect 1740 2325 1760 2425
rect 1795 2325 1800 2425
rect 1700 2310 1800 2325
rect 1950 2425 2050 2440
rect 1950 2325 1955 2425
rect 1990 2325 2010 2425
rect 2045 2325 2050 2425
rect 1950 2310 2050 2325
rect 2200 2425 2300 2440
rect 2200 2325 2205 2425
rect 2240 2325 2260 2425
rect 2295 2325 2300 2425
rect 2200 2310 2300 2325
rect 2450 2425 2550 2440
rect 2450 2325 2455 2425
rect 2490 2325 2510 2425
rect 2545 2325 2550 2425
rect 2450 2310 2550 2325
rect 2700 2425 2800 2440
rect 2700 2325 2705 2425
rect 2740 2325 2760 2425
rect 2795 2325 2800 2425
rect 2700 2310 2800 2325
rect 2950 2425 3050 2440
rect 2950 2325 2955 2425
rect 2990 2325 3010 2425
rect 3045 2325 3050 2425
rect 2950 2310 3050 2325
rect 3200 2425 3300 2440
rect 3200 2325 3205 2425
rect 3240 2325 3260 2425
rect 3295 2325 3300 2425
rect 3200 2310 3300 2325
rect 3450 2425 3550 2440
rect 3450 2325 3455 2425
rect 3490 2325 3510 2425
rect 3545 2325 3550 2425
rect 3450 2310 3550 2325
rect 3700 2425 3800 2440
rect 3700 2325 3705 2425
rect 3740 2325 3760 2425
rect 3795 2325 3800 2425
rect 3700 2310 3800 2325
rect 3950 2425 4050 2440
rect 3950 2325 3955 2425
rect 3990 2325 4010 2425
rect 4045 2325 4050 2425
rect 3950 2310 4050 2325
rect 4200 2425 4300 2440
rect 4200 2325 4205 2425
rect 4240 2325 4260 2425
rect 4295 2325 4300 2425
rect 4200 2310 4300 2325
rect 4450 2425 4550 2440
rect 4450 2325 4455 2425
rect 4490 2325 4510 2425
rect 4545 2325 4550 2425
rect 4450 2310 4550 2325
rect 4700 2425 4800 2440
rect 4700 2325 4705 2425
rect 4740 2325 4760 2425
rect 4795 2325 4800 2425
rect 4700 2310 4800 2325
rect 4950 2425 5050 2440
rect 4950 2325 4955 2425
rect 4990 2325 5010 2425
rect 5045 2325 5050 2425
rect 4950 2310 5050 2325
rect 5200 2425 5300 2440
rect 5200 2325 5205 2425
rect 5240 2325 5260 2425
rect 5295 2325 5300 2425
rect 5200 2310 5300 2325
rect 5450 2425 5550 2440
rect 5450 2325 5455 2425
rect 5490 2325 5510 2425
rect 5545 2325 5550 2425
rect 5450 2310 5550 2325
rect 5700 2425 5800 2440
rect 5700 2325 5705 2425
rect 5740 2325 5760 2425
rect 5795 2325 5800 2425
rect 5700 2310 5800 2325
rect 5950 2425 6050 2440
rect 5950 2325 5955 2425
rect 5990 2325 6010 2425
rect 6045 2325 6050 2425
rect 5950 2310 6050 2325
rect 6200 2425 6300 2440
rect 6200 2325 6205 2425
rect 6240 2325 6260 2425
rect 6295 2325 6300 2425
rect 6200 2310 6300 2325
rect 6450 2425 6550 2440
rect 6450 2325 6455 2425
rect 6490 2325 6510 2425
rect 6545 2325 6550 2425
rect 6450 2310 6550 2325
rect 6700 2425 6800 2440
rect 6700 2325 6705 2425
rect 6740 2325 6760 2425
rect 6795 2325 6800 2425
rect 6700 2310 6800 2325
rect 6950 2425 7050 2440
rect 6950 2325 6955 2425
rect 6990 2325 7010 2425
rect 7045 2325 7050 2425
rect 6950 2310 7050 2325
rect 7200 2425 7300 2440
rect 7200 2325 7205 2425
rect 7240 2325 7260 2425
rect 7295 2325 7300 2425
rect 7200 2310 7300 2325
rect 7450 2425 7550 2440
rect 7450 2325 7455 2425
rect 7490 2325 7510 2425
rect 7545 2325 7550 2425
rect 7450 2310 7550 2325
rect 7700 2425 7800 2440
rect 7700 2325 7705 2425
rect 7740 2325 7760 2425
rect 7795 2325 7800 2425
rect 7700 2310 7800 2325
rect 7950 2425 8000 2440
rect 7950 2325 7955 2425
rect 7990 2325 8000 2425
rect 7950 2310 8000 2325
rect 0 2300 60 2310
rect 190 2300 310 2310
rect 440 2300 560 2310
rect 690 2300 810 2310
rect 940 2300 1060 2310
rect 1190 2300 1310 2310
rect 1440 2300 1560 2310
rect 1690 2300 1810 2310
rect 1940 2300 2060 2310
rect 2190 2300 2310 2310
rect 2440 2300 2560 2310
rect 2690 2300 2810 2310
rect 2940 2300 3060 2310
rect 3190 2300 3310 2310
rect 3440 2300 3560 2310
rect 3690 2300 3810 2310
rect 3940 2300 4060 2310
rect 4190 2300 4310 2310
rect 4440 2300 4560 2310
rect 4690 2300 4810 2310
rect 4940 2300 5060 2310
rect 5190 2300 5310 2310
rect 5440 2300 5560 2310
rect 5690 2300 5810 2310
rect 5940 2300 6060 2310
rect 6190 2300 6310 2310
rect 6440 2300 6560 2310
rect 6690 2300 6810 2310
rect 6940 2300 7060 2310
rect 7190 2300 7310 2310
rect 7440 2300 7560 2310
rect 7690 2300 7810 2310
rect 7940 2300 8000 2310
rect 0 2295 8000 2300
rect 0 2260 75 2295
rect 175 2260 325 2295
rect 425 2260 575 2295
rect 675 2260 825 2295
rect 925 2260 1075 2295
rect 1175 2260 1325 2295
rect 1425 2260 1575 2295
rect 1675 2260 1825 2295
rect 1925 2260 2075 2295
rect 2175 2260 2325 2295
rect 2425 2260 2575 2295
rect 2675 2260 2825 2295
rect 2925 2260 3075 2295
rect 3175 2260 3325 2295
rect 3425 2260 3575 2295
rect 3675 2260 3825 2295
rect 3925 2260 4075 2295
rect 4175 2260 4325 2295
rect 4425 2260 4575 2295
rect 4675 2260 4825 2295
rect 4925 2260 5075 2295
rect 5175 2260 5325 2295
rect 5425 2260 5575 2295
rect 5675 2260 5825 2295
rect 5925 2260 6075 2295
rect 6175 2260 6325 2295
rect 6425 2260 6575 2295
rect 6675 2260 6825 2295
rect 6925 2260 7075 2295
rect 7175 2260 7325 2295
rect 7425 2260 7575 2295
rect 7675 2260 7825 2295
rect 7925 2260 8000 2295
rect 0 2240 8000 2260
rect 0 2205 75 2240
rect 175 2205 325 2240
rect 425 2205 575 2240
rect 675 2205 825 2240
rect 925 2205 1075 2240
rect 1175 2205 1325 2240
rect 1425 2205 1575 2240
rect 1675 2205 1825 2240
rect 1925 2205 2075 2240
rect 2175 2205 2325 2240
rect 2425 2205 2575 2240
rect 2675 2205 2825 2240
rect 2925 2205 3075 2240
rect 3175 2205 3325 2240
rect 3425 2205 3575 2240
rect 3675 2205 3825 2240
rect 3925 2205 4075 2240
rect 4175 2205 4325 2240
rect 4425 2205 4575 2240
rect 4675 2205 4825 2240
rect 4925 2205 5075 2240
rect 5175 2205 5325 2240
rect 5425 2205 5575 2240
rect 5675 2205 5825 2240
rect 5925 2205 6075 2240
rect 6175 2205 6325 2240
rect 6425 2205 6575 2240
rect 6675 2205 6825 2240
rect 6925 2205 7075 2240
rect 7175 2205 7325 2240
rect 7425 2205 7575 2240
rect 7675 2205 7825 2240
rect 7925 2205 8000 2240
rect 0 2200 8000 2205
rect 0 2190 60 2200
rect 190 2190 310 2200
rect 440 2190 560 2200
rect 690 2190 810 2200
rect 940 2190 1060 2200
rect 1190 2190 1310 2200
rect 1440 2190 1560 2200
rect 1690 2190 1810 2200
rect 1940 2190 2060 2200
rect 2190 2190 2310 2200
rect 2440 2190 2560 2200
rect 2690 2190 2810 2200
rect 2940 2190 3060 2200
rect 3190 2190 3310 2200
rect 3440 2190 3560 2200
rect 3690 2190 3810 2200
rect 3940 2190 4060 2200
rect 4190 2190 4310 2200
rect 4440 2190 4560 2200
rect 4690 2190 4810 2200
rect 4940 2190 5060 2200
rect 5190 2190 5310 2200
rect 5440 2190 5560 2200
rect 5690 2190 5810 2200
rect 5940 2190 6060 2200
rect 6190 2190 6310 2200
rect 6440 2190 6560 2200
rect 6690 2190 6810 2200
rect 6940 2190 7060 2200
rect 7190 2190 7310 2200
rect 7440 2190 7560 2200
rect 7690 2190 7810 2200
rect 7940 2190 8000 2200
rect 0 2175 50 2190
rect 0 2075 10 2175
rect 45 2075 50 2175
rect 0 2060 50 2075
rect 200 2175 300 2190
rect 200 2075 205 2175
rect 240 2075 260 2175
rect 295 2075 300 2175
rect 200 2060 300 2075
rect 450 2175 550 2190
rect 450 2075 455 2175
rect 490 2075 510 2175
rect 545 2075 550 2175
rect 450 2060 550 2075
rect 700 2175 800 2190
rect 700 2075 705 2175
rect 740 2075 760 2175
rect 795 2075 800 2175
rect 700 2060 800 2075
rect 950 2175 1050 2190
rect 950 2075 955 2175
rect 990 2075 1010 2175
rect 1045 2075 1050 2175
rect 950 2060 1050 2075
rect 1200 2175 1300 2190
rect 1200 2075 1205 2175
rect 1240 2075 1260 2175
rect 1295 2075 1300 2175
rect 1200 2060 1300 2075
rect 1450 2175 1550 2190
rect 1450 2075 1455 2175
rect 1490 2075 1510 2175
rect 1545 2075 1550 2175
rect 1450 2060 1550 2075
rect 1700 2175 1800 2190
rect 1700 2075 1705 2175
rect 1740 2075 1760 2175
rect 1795 2075 1800 2175
rect 1700 2060 1800 2075
rect 1950 2175 2050 2190
rect 1950 2075 1955 2175
rect 1990 2075 2010 2175
rect 2045 2075 2050 2175
rect 1950 2060 2050 2075
rect 2200 2175 2300 2190
rect 2200 2075 2205 2175
rect 2240 2075 2260 2175
rect 2295 2075 2300 2175
rect 2200 2060 2300 2075
rect 2450 2175 2550 2190
rect 2450 2075 2455 2175
rect 2490 2075 2510 2175
rect 2545 2075 2550 2175
rect 2450 2060 2550 2075
rect 2700 2175 2800 2190
rect 2700 2075 2705 2175
rect 2740 2075 2760 2175
rect 2795 2075 2800 2175
rect 2700 2060 2800 2075
rect 2950 2175 3050 2190
rect 2950 2075 2955 2175
rect 2990 2075 3010 2175
rect 3045 2075 3050 2175
rect 2950 2060 3050 2075
rect 3200 2175 3300 2190
rect 3200 2075 3205 2175
rect 3240 2075 3260 2175
rect 3295 2075 3300 2175
rect 3200 2060 3300 2075
rect 3450 2175 3550 2190
rect 3450 2075 3455 2175
rect 3490 2075 3510 2175
rect 3545 2075 3550 2175
rect 3450 2060 3550 2075
rect 3700 2175 3800 2190
rect 3700 2075 3705 2175
rect 3740 2075 3760 2175
rect 3795 2075 3800 2175
rect 3700 2060 3800 2075
rect 3950 2175 4050 2190
rect 3950 2075 3955 2175
rect 3990 2075 4010 2175
rect 4045 2075 4050 2175
rect 3950 2060 4050 2075
rect 4200 2175 4300 2190
rect 4200 2075 4205 2175
rect 4240 2075 4260 2175
rect 4295 2075 4300 2175
rect 4200 2060 4300 2075
rect 4450 2175 4550 2190
rect 4450 2075 4455 2175
rect 4490 2075 4510 2175
rect 4545 2075 4550 2175
rect 4450 2060 4550 2075
rect 4700 2175 4800 2190
rect 4700 2075 4705 2175
rect 4740 2075 4760 2175
rect 4795 2075 4800 2175
rect 4700 2060 4800 2075
rect 4950 2175 5050 2190
rect 4950 2075 4955 2175
rect 4990 2075 5010 2175
rect 5045 2075 5050 2175
rect 4950 2060 5050 2075
rect 5200 2175 5300 2190
rect 5200 2075 5205 2175
rect 5240 2075 5260 2175
rect 5295 2075 5300 2175
rect 5200 2060 5300 2075
rect 5450 2175 5550 2190
rect 5450 2075 5455 2175
rect 5490 2075 5510 2175
rect 5545 2075 5550 2175
rect 5450 2060 5550 2075
rect 5700 2175 5800 2190
rect 5700 2075 5705 2175
rect 5740 2075 5760 2175
rect 5795 2075 5800 2175
rect 5700 2060 5800 2075
rect 5950 2175 6050 2190
rect 5950 2075 5955 2175
rect 5990 2075 6010 2175
rect 6045 2075 6050 2175
rect 5950 2060 6050 2075
rect 6200 2175 6300 2190
rect 6200 2075 6205 2175
rect 6240 2075 6260 2175
rect 6295 2075 6300 2175
rect 6200 2060 6300 2075
rect 6450 2175 6550 2190
rect 6450 2075 6455 2175
rect 6490 2075 6510 2175
rect 6545 2075 6550 2175
rect 6450 2060 6550 2075
rect 6700 2175 6800 2190
rect 6700 2075 6705 2175
rect 6740 2075 6760 2175
rect 6795 2075 6800 2175
rect 6700 2060 6800 2075
rect 6950 2175 7050 2190
rect 6950 2075 6955 2175
rect 6990 2075 7010 2175
rect 7045 2075 7050 2175
rect 6950 2060 7050 2075
rect 7200 2175 7300 2190
rect 7200 2075 7205 2175
rect 7240 2075 7260 2175
rect 7295 2075 7300 2175
rect 7200 2060 7300 2075
rect 7450 2175 7550 2190
rect 7450 2075 7455 2175
rect 7490 2075 7510 2175
rect 7545 2075 7550 2175
rect 7450 2060 7550 2075
rect 7700 2175 7800 2190
rect 7700 2075 7705 2175
rect 7740 2075 7760 2175
rect 7795 2075 7800 2175
rect 7700 2060 7800 2075
rect 7950 2175 8000 2190
rect 7950 2075 7955 2175
rect 7990 2075 8000 2175
rect 7950 2060 8000 2075
rect 0 2050 60 2060
rect 190 2050 310 2060
rect 440 2050 560 2060
rect 690 2050 810 2060
rect 940 2050 1060 2060
rect 1190 2050 1310 2060
rect 1440 2050 1560 2060
rect 1690 2050 1810 2060
rect 1940 2050 2060 2060
rect 2190 2050 2310 2060
rect 2440 2050 2560 2060
rect 2690 2050 2810 2060
rect 2940 2050 3060 2060
rect 3190 2050 3310 2060
rect 3440 2050 3560 2060
rect 3690 2050 3810 2060
rect 3940 2050 4060 2060
rect 4190 2050 4310 2060
rect 4440 2050 4560 2060
rect 4690 2050 4810 2060
rect 4940 2050 5060 2060
rect 5190 2050 5310 2060
rect 5440 2050 5560 2060
rect 5690 2050 5810 2060
rect 5940 2050 6060 2060
rect 6190 2050 6310 2060
rect 6440 2050 6560 2060
rect 6690 2050 6810 2060
rect 6940 2050 7060 2060
rect 7190 2050 7310 2060
rect 7440 2050 7560 2060
rect 7690 2050 7810 2060
rect 7940 2050 8000 2060
rect 0 2045 8000 2050
rect 0 2010 75 2045
rect 175 2010 325 2045
rect 425 2010 575 2045
rect 675 2010 825 2045
rect 925 2010 1075 2045
rect 1175 2010 1325 2045
rect 1425 2010 1575 2045
rect 1675 2010 1825 2045
rect 1925 2010 2075 2045
rect 2175 2010 2325 2045
rect 2425 2010 2575 2045
rect 2675 2010 2825 2045
rect 2925 2010 3075 2045
rect 3175 2010 3325 2045
rect 3425 2010 3575 2045
rect 3675 2010 3825 2045
rect 3925 2010 4075 2045
rect 4175 2010 4325 2045
rect 4425 2010 4575 2045
rect 4675 2010 4825 2045
rect 4925 2010 5075 2045
rect 5175 2010 5325 2045
rect 5425 2010 5575 2045
rect 5675 2010 5825 2045
rect 5925 2010 6075 2045
rect 6175 2010 6325 2045
rect 6425 2010 6575 2045
rect 6675 2010 6825 2045
rect 6925 2010 7075 2045
rect 7175 2010 7325 2045
rect 7425 2010 7575 2045
rect 7675 2010 7825 2045
rect 7925 2010 8000 2045
rect 0 1990 8000 2010
rect 0 1955 75 1990
rect 175 1955 325 1990
rect 425 1955 575 1990
rect 675 1955 825 1990
rect 925 1955 1075 1990
rect 1175 1955 1325 1990
rect 1425 1955 1575 1990
rect 1675 1955 1825 1990
rect 1925 1955 2075 1990
rect 2175 1955 2325 1990
rect 2425 1955 2575 1990
rect 2675 1955 2825 1990
rect 2925 1955 3075 1990
rect 3175 1955 3325 1990
rect 3425 1955 3575 1990
rect 3675 1955 3825 1990
rect 3925 1955 4075 1990
rect 4175 1955 4325 1990
rect 4425 1955 4575 1990
rect 4675 1955 4825 1990
rect 4925 1955 5075 1990
rect 5175 1955 5325 1990
rect 5425 1955 5575 1990
rect 5675 1955 5825 1990
rect 5925 1955 6075 1990
rect 6175 1955 6325 1990
rect 6425 1955 6575 1990
rect 6675 1955 6825 1990
rect 6925 1955 7075 1990
rect 7175 1955 7325 1990
rect 7425 1955 7575 1990
rect 7675 1955 7825 1990
rect 7925 1955 8000 1990
rect 0 1950 8000 1955
rect 0 1940 60 1950
rect 190 1940 310 1950
rect 440 1940 560 1950
rect 690 1940 810 1950
rect 940 1940 1060 1950
rect 1190 1940 1310 1950
rect 1440 1940 1560 1950
rect 1690 1940 1810 1950
rect 1940 1940 2060 1950
rect 2190 1940 2310 1950
rect 2440 1940 2560 1950
rect 2690 1940 2810 1950
rect 2940 1940 3060 1950
rect 3190 1940 3310 1950
rect 3440 1940 3560 1950
rect 3690 1940 3810 1950
rect 3940 1940 4060 1950
rect 4190 1940 4310 1950
rect 4440 1940 4560 1950
rect 4690 1940 4810 1950
rect 4940 1940 5060 1950
rect 5190 1940 5310 1950
rect 5440 1940 5560 1950
rect 5690 1940 5810 1950
rect 5940 1940 6060 1950
rect 6190 1940 6310 1950
rect 6440 1940 6560 1950
rect 6690 1940 6810 1950
rect 6940 1940 7060 1950
rect 7190 1940 7310 1950
rect 7440 1940 7560 1950
rect 7690 1940 7810 1950
rect 7940 1940 8000 1950
rect 0 1925 50 1940
rect 0 1825 10 1925
rect 45 1825 50 1925
rect 0 1810 50 1825
rect 200 1925 300 1940
rect 200 1825 205 1925
rect 240 1825 260 1925
rect 295 1825 300 1925
rect 200 1810 300 1825
rect 450 1925 550 1940
rect 450 1825 455 1925
rect 490 1825 510 1925
rect 545 1825 550 1925
rect 450 1810 550 1825
rect 700 1925 800 1940
rect 700 1825 705 1925
rect 740 1825 760 1925
rect 795 1825 800 1925
rect 700 1810 800 1825
rect 950 1925 1050 1940
rect 950 1825 955 1925
rect 990 1825 1010 1925
rect 1045 1825 1050 1925
rect 950 1810 1050 1825
rect 1200 1925 1300 1940
rect 1200 1825 1205 1925
rect 1240 1825 1260 1925
rect 1295 1825 1300 1925
rect 1200 1810 1300 1825
rect 1450 1925 1550 1940
rect 1450 1825 1455 1925
rect 1490 1825 1510 1925
rect 1545 1825 1550 1925
rect 1450 1810 1550 1825
rect 1700 1925 1800 1940
rect 1700 1825 1705 1925
rect 1740 1825 1760 1925
rect 1795 1825 1800 1925
rect 1700 1810 1800 1825
rect 1950 1925 2050 1940
rect 1950 1825 1955 1925
rect 1990 1825 2010 1925
rect 2045 1825 2050 1925
rect 1950 1810 2050 1825
rect 2200 1925 2300 1940
rect 2200 1825 2205 1925
rect 2240 1825 2260 1925
rect 2295 1825 2300 1925
rect 2200 1810 2300 1825
rect 2450 1925 2550 1940
rect 2450 1825 2455 1925
rect 2490 1825 2510 1925
rect 2545 1825 2550 1925
rect 2450 1810 2550 1825
rect 2700 1925 2800 1940
rect 2700 1825 2705 1925
rect 2740 1825 2760 1925
rect 2795 1825 2800 1925
rect 2700 1810 2800 1825
rect 2950 1925 3050 1940
rect 2950 1825 2955 1925
rect 2990 1825 3010 1925
rect 3045 1825 3050 1925
rect 2950 1810 3050 1825
rect 3200 1925 3300 1940
rect 3200 1825 3205 1925
rect 3240 1825 3260 1925
rect 3295 1825 3300 1925
rect 3200 1810 3300 1825
rect 3450 1925 3550 1940
rect 3450 1825 3455 1925
rect 3490 1825 3510 1925
rect 3545 1825 3550 1925
rect 3450 1810 3550 1825
rect 3700 1925 3800 1940
rect 3700 1825 3705 1925
rect 3740 1825 3760 1925
rect 3795 1825 3800 1925
rect 3700 1810 3800 1825
rect 3950 1925 4050 1940
rect 3950 1825 3955 1925
rect 3990 1825 4010 1925
rect 4045 1825 4050 1925
rect 3950 1810 4050 1825
rect 4200 1925 4300 1940
rect 4200 1825 4205 1925
rect 4240 1825 4260 1925
rect 4295 1825 4300 1925
rect 4200 1810 4300 1825
rect 4450 1925 4550 1940
rect 4450 1825 4455 1925
rect 4490 1825 4510 1925
rect 4545 1825 4550 1925
rect 4450 1810 4550 1825
rect 4700 1925 4800 1940
rect 4700 1825 4705 1925
rect 4740 1825 4760 1925
rect 4795 1825 4800 1925
rect 4700 1810 4800 1825
rect 4950 1925 5050 1940
rect 4950 1825 4955 1925
rect 4990 1825 5010 1925
rect 5045 1825 5050 1925
rect 4950 1810 5050 1825
rect 5200 1925 5300 1940
rect 5200 1825 5205 1925
rect 5240 1825 5260 1925
rect 5295 1825 5300 1925
rect 5200 1810 5300 1825
rect 5450 1925 5550 1940
rect 5450 1825 5455 1925
rect 5490 1825 5510 1925
rect 5545 1825 5550 1925
rect 5450 1810 5550 1825
rect 5700 1925 5800 1940
rect 5700 1825 5705 1925
rect 5740 1825 5760 1925
rect 5795 1825 5800 1925
rect 5700 1810 5800 1825
rect 5950 1925 6050 1940
rect 5950 1825 5955 1925
rect 5990 1825 6010 1925
rect 6045 1825 6050 1925
rect 5950 1810 6050 1825
rect 6200 1925 6300 1940
rect 6200 1825 6205 1925
rect 6240 1825 6260 1925
rect 6295 1825 6300 1925
rect 6200 1810 6300 1825
rect 6450 1925 6550 1940
rect 6450 1825 6455 1925
rect 6490 1825 6510 1925
rect 6545 1825 6550 1925
rect 6450 1810 6550 1825
rect 6700 1925 6800 1940
rect 6700 1825 6705 1925
rect 6740 1825 6760 1925
rect 6795 1825 6800 1925
rect 6700 1810 6800 1825
rect 6950 1925 7050 1940
rect 6950 1825 6955 1925
rect 6990 1825 7010 1925
rect 7045 1825 7050 1925
rect 6950 1810 7050 1825
rect 7200 1925 7300 1940
rect 7200 1825 7205 1925
rect 7240 1825 7260 1925
rect 7295 1825 7300 1925
rect 7200 1810 7300 1825
rect 7450 1925 7550 1940
rect 7450 1825 7455 1925
rect 7490 1825 7510 1925
rect 7545 1825 7550 1925
rect 7450 1810 7550 1825
rect 7700 1925 7800 1940
rect 7700 1825 7705 1925
rect 7740 1825 7760 1925
rect 7795 1825 7800 1925
rect 7700 1810 7800 1825
rect 7950 1925 8000 1940
rect 7950 1825 7955 1925
rect 7990 1825 8000 1925
rect 7950 1810 8000 1825
rect 0 1800 60 1810
rect 190 1800 310 1810
rect 440 1800 560 1810
rect 690 1800 810 1810
rect 940 1800 1060 1810
rect 1190 1800 1310 1810
rect 1440 1800 1560 1810
rect 1690 1800 1810 1810
rect 1940 1800 2060 1810
rect 2190 1800 2310 1810
rect 2440 1800 2560 1810
rect 2690 1800 2810 1810
rect 2940 1800 3060 1810
rect 3190 1800 3310 1810
rect 3440 1800 3560 1810
rect 3690 1800 3810 1810
rect 3940 1800 4060 1810
rect 4190 1800 4310 1810
rect 4440 1800 4560 1810
rect 4690 1800 4810 1810
rect 4940 1800 5060 1810
rect 5190 1800 5310 1810
rect 5440 1800 5560 1810
rect 5690 1800 5810 1810
rect 5940 1800 6060 1810
rect 6190 1800 6310 1810
rect 6440 1800 6560 1810
rect 6690 1800 6810 1810
rect 6940 1800 7060 1810
rect 7190 1800 7310 1810
rect 7440 1800 7560 1810
rect 7690 1800 7810 1810
rect 7940 1800 8000 1810
rect 0 1795 8000 1800
rect 0 1760 75 1795
rect 175 1760 325 1795
rect 425 1760 575 1795
rect 675 1760 825 1795
rect 925 1760 1075 1795
rect 1175 1760 1325 1795
rect 1425 1760 1575 1795
rect 1675 1760 1825 1795
rect 1925 1760 2075 1795
rect 2175 1760 2325 1795
rect 2425 1760 2575 1795
rect 2675 1760 2825 1795
rect 2925 1760 3075 1795
rect 3175 1760 3325 1795
rect 3425 1760 3575 1795
rect 3675 1760 3825 1795
rect 3925 1760 4075 1795
rect 4175 1760 4325 1795
rect 4425 1760 4575 1795
rect 4675 1760 4825 1795
rect 4925 1760 5075 1795
rect 5175 1760 5325 1795
rect 5425 1760 5575 1795
rect 5675 1760 5825 1795
rect 5925 1760 6075 1795
rect 6175 1760 6325 1795
rect 6425 1760 6575 1795
rect 6675 1760 6825 1795
rect 6925 1760 7075 1795
rect 7175 1760 7325 1795
rect 7425 1760 7575 1795
rect 7675 1760 7825 1795
rect 7925 1760 8000 1795
rect 0 1740 8000 1760
rect 0 1705 75 1740
rect 175 1705 325 1740
rect 425 1705 575 1740
rect 675 1705 825 1740
rect 925 1705 1075 1740
rect 1175 1705 1325 1740
rect 1425 1705 1575 1740
rect 1675 1705 1825 1740
rect 1925 1705 2075 1740
rect 2175 1705 2325 1740
rect 2425 1705 2575 1740
rect 2675 1705 2825 1740
rect 2925 1705 3075 1740
rect 3175 1705 3325 1740
rect 3425 1705 3575 1740
rect 3675 1705 3825 1740
rect 3925 1705 4075 1740
rect 4175 1705 4325 1740
rect 4425 1705 4575 1740
rect 4675 1705 4825 1740
rect 4925 1705 5075 1740
rect 5175 1705 5325 1740
rect 5425 1705 5575 1740
rect 5675 1705 5825 1740
rect 5925 1705 6075 1740
rect 6175 1705 6325 1740
rect 6425 1705 6575 1740
rect 6675 1705 6825 1740
rect 6925 1705 7075 1740
rect 7175 1705 7325 1740
rect 7425 1705 7575 1740
rect 7675 1705 7825 1740
rect 7925 1705 8000 1740
rect 0 1700 8000 1705
rect 0 1690 60 1700
rect 190 1690 310 1700
rect 440 1690 560 1700
rect 690 1690 810 1700
rect 940 1690 1060 1700
rect 1190 1690 1310 1700
rect 1440 1690 1560 1700
rect 1690 1690 1810 1700
rect 1940 1690 2060 1700
rect 2190 1690 2310 1700
rect 2440 1690 2560 1700
rect 2690 1690 2810 1700
rect 2940 1690 3060 1700
rect 3190 1690 3310 1700
rect 3440 1690 3560 1700
rect 3690 1690 3810 1700
rect 3940 1690 4060 1700
rect 4190 1690 4310 1700
rect 4440 1690 4560 1700
rect 4690 1690 4810 1700
rect 4940 1690 5060 1700
rect 5190 1690 5310 1700
rect 5440 1690 5560 1700
rect 5690 1690 5810 1700
rect 5940 1690 6060 1700
rect 6190 1690 6310 1700
rect 6440 1690 6560 1700
rect 6690 1690 6810 1700
rect 6940 1690 7060 1700
rect 7190 1690 7310 1700
rect 7440 1690 7560 1700
rect 7690 1690 7810 1700
rect 7940 1690 8000 1700
rect 0 1675 50 1690
rect 0 1575 10 1675
rect 45 1575 50 1675
rect 0 1560 50 1575
rect 200 1675 300 1690
rect 200 1575 205 1675
rect 240 1575 260 1675
rect 295 1575 300 1675
rect 200 1560 300 1575
rect 450 1675 550 1690
rect 450 1575 455 1675
rect 490 1575 510 1675
rect 545 1575 550 1675
rect 450 1560 550 1575
rect 700 1675 800 1690
rect 700 1575 705 1675
rect 740 1575 760 1675
rect 795 1575 800 1675
rect 700 1560 800 1575
rect 950 1675 1050 1690
rect 950 1575 955 1675
rect 990 1575 1010 1675
rect 1045 1575 1050 1675
rect 950 1560 1050 1575
rect 1200 1675 1300 1690
rect 1200 1575 1205 1675
rect 1240 1575 1260 1675
rect 1295 1575 1300 1675
rect 1200 1560 1300 1575
rect 1450 1675 1550 1690
rect 1450 1575 1455 1675
rect 1490 1575 1510 1675
rect 1545 1575 1550 1675
rect 1450 1560 1550 1575
rect 1700 1675 1800 1690
rect 1700 1575 1705 1675
rect 1740 1575 1760 1675
rect 1795 1575 1800 1675
rect 1700 1560 1800 1575
rect 1950 1675 2050 1690
rect 1950 1575 1955 1675
rect 1990 1575 2010 1675
rect 2045 1575 2050 1675
rect 1950 1560 2050 1575
rect 2200 1675 2300 1690
rect 2200 1575 2205 1675
rect 2240 1575 2260 1675
rect 2295 1575 2300 1675
rect 2200 1560 2300 1575
rect 2450 1675 2550 1690
rect 2450 1575 2455 1675
rect 2490 1575 2510 1675
rect 2545 1575 2550 1675
rect 2450 1560 2550 1575
rect 2700 1675 2800 1690
rect 2700 1575 2705 1675
rect 2740 1575 2760 1675
rect 2795 1575 2800 1675
rect 2700 1560 2800 1575
rect 2950 1675 3050 1690
rect 2950 1575 2955 1675
rect 2990 1575 3010 1675
rect 3045 1575 3050 1675
rect 2950 1560 3050 1575
rect 3200 1675 3300 1690
rect 3200 1575 3205 1675
rect 3240 1575 3260 1675
rect 3295 1575 3300 1675
rect 3200 1560 3300 1575
rect 3450 1675 3550 1690
rect 3450 1575 3455 1675
rect 3490 1575 3510 1675
rect 3545 1575 3550 1675
rect 3450 1560 3550 1575
rect 3700 1675 3800 1690
rect 3700 1575 3705 1675
rect 3740 1575 3760 1675
rect 3795 1575 3800 1675
rect 3700 1560 3800 1575
rect 3950 1675 4050 1690
rect 3950 1575 3955 1675
rect 3990 1575 4010 1675
rect 4045 1575 4050 1675
rect 3950 1560 4050 1575
rect 4200 1675 4300 1690
rect 4200 1575 4205 1675
rect 4240 1575 4260 1675
rect 4295 1575 4300 1675
rect 4200 1560 4300 1575
rect 4450 1675 4550 1690
rect 4450 1575 4455 1675
rect 4490 1575 4510 1675
rect 4545 1575 4550 1675
rect 4450 1560 4550 1575
rect 4700 1675 4800 1690
rect 4700 1575 4705 1675
rect 4740 1575 4760 1675
rect 4795 1575 4800 1675
rect 4700 1560 4800 1575
rect 4950 1675 5050 1690
rect 4950 1575 4955 1675
rect 4990 1575 5010 1675
rect 5045 1575 5050 1675
rect 4950 1560 5050 1575
rect 5200 1675 5300 1690
rect 5200 1575 5205 1675
rect 5240 1575 5260 1675
rect 5295 1575 5300 1675
rect 5200 1560 5300 1575
rect 5450 1675 5550 1690
rect 5450 1575 5455 1675
rect 5490 1575 5510 1675
rect 5545 1575 5550 1675
rect 5450 1560 5550 1575
rect 5700 1675 5800 1690
rect 5700 1575 5705 1675
rect 5740 1575 5760 1675
rect 5795 1575 5800 1675
rect 5700 1560 5800 1575
rect 5950 1675 6050 1690
rect 5950 1575 5955 1675
rect 5990 1575 6010 1675
rect 6045 1575 6050 1675
rect 5950 1560 6050 1575
rect 6200 1675 6300 1690
rect 6200 1575 6205 1675
rect 6240 1575 6260 1675
rect 6295 1575 6300 1675
rect 6200 1560 6300 1575
rect 6450 1675 6550 1690
rect 6450 1575 6455 1675
rect 6490 1575 6510 1675
rect 6545 1575 6550 1675
rect 6450 1560 6550 1575
rect 6700 1675 6800 1690
rect 6700 1575 6705 1675
rect 6740 1575 6760 1675
rect 6795 1575 6800 1675
rect 6700 1560 6800 1575
rect 6950 1675 7050 1690
rect 6950 1575 6955 1675
rect 6990 1575 7010 1675
rect 7045 1575 7050 1675
rect 6950 1560 7050 1575
rect 7200 1675 7300 1690
rect 7200 1575 7205 1675
rect 7240 1575 7260 1675
rect 7295 1575 7300 1675
rect 7200 1560 7300 1575
rect 7450 1675 7550 1690
rect 7450 1575 7455 1675
rect 7490 1575 7510 1675
rect 7545 1575 7550 1675
rect 7450 1560 7550 1575
rect 7700 1675 7800 1690
rect 7700 1575 7705 1675
rect 7740 1575 7760 1675
rect 7795 1575 7800 1675
rect 7700 1560 7800 1575
rect 7950 1675 8000 1690
rect 7950 1575 7955 1675
rect 7990 1575 8000 1675
rect 7950 1560 8000 1575
rect 0 1550 60 1560
rect 190 1550 310 1560
rect 440 1550 560 1560
rect 690 1550 810 1560
rect 940 1550 1060 1560
rect 1190 1550 1310 1560
rect 1440 1550 1560 1560
rect 1690 1550 1810 1560
rect 1940 1550 2060 1560
rect 2190 1550 2310 1560
rect 2440 1550 2560 1560
rect 2690 1550 2810 1560
rect 2940 1550 3060 1560
rect 3190 1550 3310 1560
rect 3440 1550 3560 1560
rect 3690 1550 3810 1560
rect 3940 1550 4060 1560
rect 4190 1550 4310 1560
rect 4440 1550 4560 1560
rect 4690 1550 4810 1560
rect 4940 1550 5060 1560
rect 5190 1550 5310 1560
rect 5440 1550 5560 1560
rect 5690 1550 5810 1560
rect 5940 1550 6060 1560
rect 6190 1550 6310 1560
rect 6440 1550 6560 1560
rect 6690 1550 6810 1560
rect 6940 1550 7060 1560
rect 7190 1550 7310 1560
rect 7440 1550 7560 1560
rect 7690 1550 7810 1560
rect 7940 1550 8000 1560
rect 0 1545 8000 1550
rect 0 1510 75 1545
rect 175 1510 325 1545
rect 425 1510 575 1545
rect 675 1510 825 1545
rect 925 1510 1075 1545
rect 1175 1510 1325 1545
rect 1425 1510 1575 1545
rect 1675 1510 1825 1545
rect 1925 1510 2075 1545
rect 2175 1510 2325 1545
rect 2425 1510 2575 1545
rect 2675 1510 2825 1545
rect 2925 1510 3075 1545
rect 3175 1510 3325 1545
rect 3425 1510 3575 1545
rect 3675 1510 3825 1545
rect 3925 1510 4075 1545
rect 4175 1510 4325 1545
rect 4425 1510 4575 1545
rect 4675 1510 4825 1545
rect 4925 1510 5075 1545
rect 5175 1510 5325 1545
rect 5425 1510 5575 1545
rect 5675 1510 5825 1545
rect 5925 1510 6075 1545
rect 6175 1510 6325 1545
rect 6425 1510 6575 1545
rect 6675 1510 6825 1545
rect 6925 1510 7075 1545
rect 7175 1510 7325 1545
rect 7425 1510 7575 1545
rect 7675 1510 7825 1545
rect 7925 1510 8000 1545
rect 0 1490 8000 1510
rect 0 1455 75 1490
rect 175 1455 325 1490
rect 425 1455 575 1490
rect 675 1455 825 1490
rect 925 1455 1075 1490
rect 1175 1455 1325 1490
rect 1425 1455 1575 1490
rect 1675 1455 1825 1490
rect 1925 1455 2075 1490
rect 2175 1455 2325 1490
rect 2425 1455 2575 1490
rect 2675 1455 2825 1490
rect 2925 1455 3075 1490
rect 3175 1455 3325 1490
rect 3425 1455 3575 1490
rect 3675 1455 3825 1490
rect 3925 1455 4075 1490
rect 4175 1455 4325 1490
rect 4425 1455 4575 1490
rect 4675 1455 4825 1490
rect 4925 1455 5075 1490
rect 5175 1455 5325 1490
rect 5425 1455 5575 1490
rect 5675 1455 5825 1490
rect 5925 1455 6075 1490
rect 6175 1455 6325 1490
rect 6425 1455 6575 1490
rect 6675 1455 6825 1490
rect 6925 1455 7075 1490
rect 7175 1455 7325 1490
rect 7425 1455 7575 1490
rect 7675 1455 7825 1490
rect 7925 1455 8000 1490
rect 0 1450 8000 1455
rect 0 1440 60 1450
rect 190 1440 310 1450
rect 440 1440 560 1450
rect 690 1440 810 1450
rect 940 1440 1060 1450
rect 1190 1440 1310 1450
rect 1440 1440 1560 1450
rect 1690 1440 1810 1450
rect 1940 1440 2060 1450
rect 2190 1440 2310 1450
rect 2440 1440 2560 1450
rect 2690 1440 2810 1450
rect 2940 1440 3060 1450
rect 3190 1440 3310 1450
rect 3440 1440 3560 1450
rect 3690 1440 3810 1450
rect 3940 1440 4060 1450
rect 4190 1440 4310 1450
rect 4440 1440 4560 1450
rect 4690 1440 4810 1450
rect 4940 1440 5060 1450
rect 5190 1440 5310 1450
rect 5440 1440 5560 1450
rect 5690 1440 5810 1450
rect 5940 1440 6060 1450
rect 6190 1440 6310 1450
rect 6440 1440 6560 1450
rect 6690 1440 6810 1450
rect 6940 1440 7060 1450
rect 7190 1440 7310 1450
rect 7440 1440 7560 1450
rect 7690 1440 7810 1450
rect 7940 1440 8000 1450
rect 0 1425 50 1440
rect 0 1325 10 1425
rect 45 1325 50 1425
rect 0 1310 50 1325
rect 200 1425 300 1440
rect 200 1325 205 1425
rect 240 1325 260 1425
rect 295 1325 300 1425
rect 200 1310 300 1325
rect 450 1425 550 1440
rect 450 1325 455 1425
rect 490 1325 510 1425
rect 545 1325 550 1425
rect 450 1310 550 1325
rect 700 1425 800 1440
rect 700 1325 705 1425
rect 740 1325 760 1425
rect 795 1325 800 1425
rect 700 1310 800 1325
rect 950 1425 1050 1440
rect 950 1325 955 1425
rect 990 1325 1010 1425
rect 1045 1325 1050 1425
rect 950 1310 1050 1325
rect 1200 1425 1300 1440
rect 1200 1325 1205 1425
rect 1240 1325 1260 1425
rect 1295 1325 1300 1425
rect 1200 1310 1300 1325
rect 1450 1425 1550 1440
rect 1450 1325 1455 1425
rect 1490 1325 1510 1425
rect 1545 1325 1550 1425
rect 1450 1310 1550 1325
rect 1700 1425 1800 1440
rect 1700 1325 1705 1425
rect 1740 1325 1760 1425
rect 1795 1325 1800 1425
rect 1700 1310 1800 1325
rect 1950 1425 2050 1440
rect 1950 1325 1955 1425
rect 1990 1325 2010 1425
rect 2045 1325 2050 1425
rect 1950 1310 2050 1325
rect 2200 1425 2300 1440
rect 2200 1325 2205 1425
rect 2240 1325 2260 1425
rect 2295 1325 2300 1425
rect 2200 1310 2300 1325
rect 2450 1425 2550 1440
rect 2450 1325 2455 1425
rect 2490 1325 2510 1425
rect 2545 1325 2550 1425
rect 2450 1310 2550 1325
rect 2700 1425 2800 1440
rect 2700 1325 2705 1425
rect 2740 1325 2760 1425
rect 2795 1325 2800 1425
rect 2700 1310 2800 1325
rect 2950 1425 3050 1440
rect 2950 1325 2955 1425
rect 2990 1325 3010 1425
rect 3045 1325 3050 1425
rect 2950 1310 3050 1325
rect 3200 1425 3300 1440
rect 3200 1325 3205 1425
rect 3240 1325 3260 1425
rect 3295 1325 3300 1425
rect 3200 1310 3300 1325
rect 3450 1425 3550 1440
rect 3450 1325 3455 1425
rect 3490 1325 3510 1425
rect 3545 1325 3550 1425
rect 3450 1310 3550 1325
rect 3700 1425 3800 1440
rect 3700 1325 3705 1425
rect 3740 1325 3760 1425
rect 3795 1325 3800 1425
rect 3700 1310 3800 1325
rect 3950 1425 4050 1440
rect 3950 1325 3955 1425
rect 3990 1325 4010 1425
rect 4045 1325 4050 1425
rect 3950 1310 4050 1325
rect 4200 1425 4300 1440
rect 4200 1325 4205 1425
rect 4240 1325 4260 1425
rect 4295 1325 4300 1425
rect 4200 1310 4300 1325
rect 4450 1425 4550 1440
rect 4450 1325 4455 1425
rect 4490 1325 4510 1425
rect 4545 1325 4550 1425
rect 4450 1310 4550 1325
rect 4700 1425 4800 1440
rect 4700 1325 4705 1425
rect 4740 1325 4760 1425
rect 4795 1325 4800 1425
rect 4700 1310 4800 1325
rect 4950 1425 5050 1440
rect 4950 1325 4955 1425
rect 4990 1325 5010 1425
rect 5045 1325 5050 1425
rect 4950 1310 5050 1325
rect 5200 1425 5300 1440
rect 5200 1325 5205 1425
rect 5240 1325 5260 1425
rect 5295 1325 5300 1425
rect 5200 1310 5300 1325
rect 5450 1425 5550 1440
rect 5450 1325 5455 1425
rect 5490 1325 5510 1425
rect 5545 1325 5550 1425
rect 5450 1310 5550 1325
rect 5700 1425 5800 1440
rect 5700 1325 5705 1425
rect 5740 1325 5760 1425
rect 5795 1325 5800 1425
rect 5700 1310 5800 1325
rect 5950 1425 6050 1440
rect 5950 1325 5955 1425
rect 5990 1325 6010 1425
rect 6045 1325 6050 1425
rect 5950 1310 6050 1325
rect 6200 1425 6300 1440
rect 6200 1325 6205 1425
rect 6240 1325 6260 1425
rect 6295 1325 6300 1425
rect 6200 1310 6300 1325
rect 6450 1425 6550 1440
rect 6450 1325 6455 1425
rect 6490 1325 6510 1425
rect 6545 1325 6550 1425
rect 6450 1310 6550 1325
rect 6700 1425 6800 1440
rect 6700 1325 6705 1425
rect 6740 1325 6760 1425
rect 6795 1325 6800 1425
rect 6700 1310 6800 1325
rect 6950 1425 7050 1440
rect 6950 1325 6955 1425
rect 6990 1325 7010 1425
rect 7045 1325 7050 1425
rect 6950 1310 7050 1325
rect 7200 1425 7300 1440
rect 7200 1325 7205 1425
rect 7240 1325 7260 1425
rect 7295 1325 7300 1425
rect 7200 1310 7300 1325
rect 7450 1425 7550 1440
rect 7450 1325 7455 1425
rect 7490 1325 7510 1425
rect 7545 1325 7550 1425
rect 7450 1310 7550 1325
rect 7700 1425 7800 1440
rect 7700 1325 7705 1425
rect 7740 1325 7760 1425
rect 7795 1325 7800 1425
rect 7700 1310 7800 1325
rect 7950 1425 8000 1440
rect 7950 1325 7955 1425
rect 7990 1325 8000 1425
rect 7950 1310 8000 1325
rect 0 1300 60 1310
rect 190 1300 310 1310
rect 440 1300 560 1310
rect 690 1300 810 1310
rect 940 1300 1060 1310
rect 1190 1300 1310 1310
rect 1440 1300 1560 1310
rect 1690 1300 1810 1310
rect 1940 1300 2060 1310
rect 2190 1300 2310 1310
rect 2440 1300 2560 1310
rect 2690 1300 2810 1310
rect 2940 1300 3060 1310
rect 3190 1300 3310 1310
rect 3440 1300 3560 1310
rect 3690 1300 3810 1310
rect 3940 1300 4060 1310
rect 4190 1300 4310 1310
rect 4440 1300 4560 1310
rect 4690 1300 4810 1310
rect 4940 1300 5060 1310
rect 5190 1300 5310 1310
rect 5440 1300 5560 1310
rect 5690 1300 5810 1310
rect 5940 1300 6060 1310
rect 6190 1300 6310 1310
rect 6440 1300 6560 1310
rect 6690 1300 6810 1310
rect 6940 1300 7060 1310
rect 7190 1300 7310 1310
rect 7440 1300 7560 1310
rect 7690 1300 7810 1310
rect 7940 1300 8000 1310
rect 0 1295 8000 1300
rect 0 1260 75 1295
rect 175 1260 325 1295
rect 425 1260 575 1295
rect 675 1260 825 1295
rect 925 1260 1075 1295
rect 1175 1260 1325 1295
rect 1425 1260 1575 1295
rect 1675 1260 1825 1295
rect 1925 1260 2075 1295
rect 2175 1260 2325 1295
rect 2425 1260 2575 1295
rect 2675 1260 2825 1295
rect 2925 1260 3075 1295
rect 3175 1260 3325 1295
rect 3425 1260 3575 1295
rect 3675 1260 3825 1295
rect 3925 1260 4075 1295
rect 4175 1260 4325 1295
rect 4425 1260 4575 1295
rect 4675 1260 4825 1295
rect 4925 1260 5075 1295
rect 5175 1260 5325 1295
rect 5425 1260 5575 1295
rect 5675 1260 5825 1295
rect 5925 1260 6075 1295
rect 6175 1260 6325 1295
rect 6425 1260 6575 1295
rect 6675 1260 6825 1295
rect 6925 1260 7075 1295
rect 7175 1260 7325 1295
rect 7425 1260 7575 1295
rect 7675 1260 7825 1295
rect 7925 1260 8000 1295
rect 0 1240 8000 1260
rect 0 1205 75 1240
rect 175 1205 325 1240
rect 425 1205 575 1240
rect 675 1205 825 1240
rect 925 1205 1075 1240
rect 1175 1205 1325 1240
rect 1425 1205 1575 1240
rect 1675 1205 1825 1240
rect 1925 1205 2075 1240
rect 2175 1205 2325 1240
rect 2425 1205 2575 1240
rect 2675 1205 2825 1240
rect 2925 1205 3075 1240
rect 3175 1205 3325 1240
rect 3425 1205 3575 1240
rect 3675 1205 3825 1240
rect 3925 1205 4075 1240
rect 4175 1205 4325 1240
rect 4425 1205 4575 1240
rect 4675 1205 4825 1240
rect 4925 1205 5075 1240
rect 5175 1205 5325 1240
rect 5425 1205 5575 1240
rect 5675 1205 5825 1240
rect 5925 1205 6075 1240
rect 6175 1205 6325 1240
rect 6425 1205 6575 1240
rect 6675 1205 6825 1240
rect 6925 1205 7075 1240
rect 7175 1205 7325 1240
rect 7425 1205 7575 1240
rect 7675 1205 7825 1240
rect 7925 1205 8000 1240
rect 0 1200 8000 1205
rect 0 1190 60 1200
rect 190 1190 310 1200
rect 440 1190 560 1200
rect 690 1190 810 1200
rect 940 1190 1060 1200
rect 1190 1190 1310 1200
rect 1440 1190 1560 1200
rect 1690 1190 1810 1200
rect 1940 1190 2060 1200
rect 2190 1190 2310 1200
rect 2440 1190 2560 1200
rect 2690 1190 2810 1200
rect 2940 1190 3060 1200
rect 3190 1190 3310 1200
rect 3440 1190 3560 1200
rect 3690 1190 3810 1200
rect 3940 1190 4060 1200
rect 4190 1190 4310 1200
rect 4440 1190 4560 1200
rect 4690 1190 4810 1200
rect 4940 1190 5060 1200
rect 5190 1190 5310 1200
rect 5440 1190 5560 1200
rect 5690 1190 5810 1200
rect 5940 1190 6060 1200
rect 6190 1190 6310 1200
rect 6440 1190 6560 1200
rect 6690 1190 6810 1200
rect 6940 1190 7060 1200
rect 7190 1190 7310 1200
rect 7440 1190 7560 1200
rect 7690 1190 7810 1200
rect 7940 1190 8000 1200
rect 0 1175 50 1190
rect 0 1075 10 1175
rect 45 1075 50 1175
rect 0 1060 50 1075
rect 200 1175 300 1190
rect 200 1075 205 1175
rect 240 1075 260 1175
rect 295 1075 300 1175
rect 200 1060 300 1075
rect 450 1175 550 1190
rect 450 1075 455 1175
rect 490 1075 510 1175
rect 545 1075 550 1175
rect 450 1060 550 1075
rect 700 1175 800 1190
rect 700 1075 705 1175
rect 740 1075 760 1175
rect 795 1075 800 1175
rect 700 1060 800 1075
rect 950 1175 1050 1190
rect 950 1075 955 1175
rect 990 1075 1010 1175
rect 1045 1075 1050 1175
rect 950 1060 1050 1075
rect 1200 1175 1300 1190
rect 1200 1075 1205 1175
rect 1240 1075 1260 1175
rect 1295 1075 1300 1175
rect 1200 1060 1300 1075
rect 1450 1175 1550 1190
rect 1450 1075 1455 1175
rect 1490 1075 1510 1175
rect 1545 1075 1550 1175
rect 1450 1060 1550 1075
rect 1700 1175 1800 1190
rect 1700 1075 1705 1175
rect 1740 1075 1760 1175
rect 1795 1075 1800 1175
rect 1700 1060 1800 1075
rect 1950 1175 2050 1190
rect 1950 1075 1955 1175
rect 1990 1075 2010 1175
rect 2045 1075 2050 1175
rect 1950 1060 2050 1075
rect 2200 1175 2300 1190
rect 2200 1075 2205 1175
rect 2240 1075 2260 1175
rect 2295 1075 2300 1175
rect 2200 1060 2300 1075
rect 2450 1175 2550 1190
rect 2450 1075 2455 1175
rect 2490 1075 2510 1175
rect 2545 1075 2550 1175
rect 2450 1060 2550 1075
rect 2700 1175 2800 1190
rect 2700 1075 2705 1175
rect 2740 1075 2760 1175
rect 2795 1075 2800 1175
rect 2700 1060 2800 1075
rect 2950 1175 3050 1190
rect 2950 1075 2955 1175
rect 2990 1075 3010 1175
rect 3045 1075 3050 1175
rect 2950 1060 3050 1075
rect 3200 1175 3300 1190
rect 3200 1075 3205 1175
rect 3240 1075 3260 1175
rect 3295 1075 3300 1175
rect 3200 1060 3300 1075
rect 3450 1175 3550 1190
rect 3450 1075 3455 1175
rect 3490 1075 3510 1175
rect 3545 1075 3550 1175
rect 3450 1060 3550 1075
rect 3700 1175 3800 1190
rect 3700 1075 3705 1175
rect 3740 1075 3760 1175
rect 3795 1075 3800 1175
rect 3700 1060 3800 1075
rect 3950 1175 4050 1190
rect 3950 1075 3955 1175
rect 3990 1075 4010 1175
rect 4045 1075 4050 1175
rect 3950 1060 4050 1075
rect 4200 1175 4300 1190
rect 4200 1075 4205 1175
rect 4240 1075 4260 1175
rect 4295 1075 4300 1175
rect 4200 1060 4300 1075
rect 4450 1175 4550 1190
rect 4450 1075 4455 1175
rect 4490 1075 4510 1175
rect 4545 1075 4550 1175
rect 4450 1060 4550 1075
rect 4700 1175 4800 1190
rect 4700 1075 4705 1175
rect 4740 1075 4760 1175
rect 4795 1075 4800 1175
rect 4700 1060 4800 1075
rect 4950 1175 5050 1190
rect 4950 1075 4955 1175
rect 4990 1075 5010 1175
rect 5045 1075 5050 1175
rect 4950 1060 5050 1075
rect 5200 1175 5300 1190
rect 5200 1075 5205 1175
rect 5240 1075 5260 1175
rect 5295 1075 5300 1175
rect 5200 1060 5300 1075
rect 5450 1175 5550 1190
rect 5450 1075 5455 1175
rect 5490 1075 5510 1175
rect 5545 1075 5550 1175
rect 5450 1060 5550 1075
rect 5700 1175 5800 1190
rect 5700 1075 5705 1175
rect 5740 1075 5760 1175
rect 5795 1075 5800 1175
rect 5700 1060 5800 1075
rect 5950 1175 6050 1190
rect 5950 1075 5955 1175
rect 5990 1075 6010 1175
rect 6045 1075 6050 1175
rect 5950 1060 6050 1075
rect 6200 1175 6300 1190
rect 6200 1075 6205 1175
rect 6240 1075 6260 1175
rect 6295 1075 6300 1175
rect 6200 1060 6300 1075
rect 6450 1175 6550 1190
rect 6450 1075 6455 1175
rect 6490 1075 6510 1175
rect 6545 1075 6550 1175
rect 6450 1060 6550 1075
rect 6700 1175 6800 1190
rect 6700 1075 6705 1175
rect 6740 1075 6760 1175
rect 6795 1075 6800 1175
rect 6700 1060 6800 1075
rect 6950 1175 7050 1190
rect 6950 1075 6955 1175
rect 6990 1075 7010 1175
rect 7045 1075 7050 1175
rect 6950 1060 7050 1075
rect 7200 1175 7300 1190
rect 7200 1075 7205 1175
rect 7240 1075 7260 1175
rect 7295 1075 7300 1175
rect 7200 1060 7300 1075
rect 7450 1175 7550 1190
rect 7450 1075 7455 1175
rect 7490 1075 7510 1175
rect 7545 1075 7550 1175
rect 7450 1060 7550 1075
rect 7700 1175 7800 1190
rect 7700 1075 7705 1175
rect 7740 1075 7760 1175
rect 7795 1075 7800 1175
rect 7700 1060 7800 1075
rect 7950 1175 8000 1190
rect 7950 1075 7955 1175
rect 7990 1075 8000 1175
rect 7950 1060 8000 1075
rect 0 1050 60 1060
rect 190 1050 310 1060
rect 440 1050 560 1060
rect 690 1050 810 1060
rect 940 1050 1060 1060
rect 1190 1050 1310 1060
rect 1440 1050 1560 1060
rect 1690 1050 1810 1060
rect 1940 1050 2060 1060
rect 2190 1050 2310 1060
rect 2440 1050 2560 1060
rect 2690 1050 2810 1060
rect 2940 1050 3060 1060
rect 3190 1050 3310 1060
rect 3440 1050 3560 1060
rect 3690 1050 3810 1060
rect 3940 1050 4060 1060
rect 4190 1050 4310 1060
rect 4440 1050 4560 1060
rect 4690 1050 4810 1060
rect 4940 1050 5060 1060
rect 5190 1050 5310 1060
rect 5440 1050 5560 1060
rect 5690 1050 5810 1060
rect 5940 1050 6060 1060
rect 6190 1050 6310 1060
rect 6440 1050 6560 1060
rect 6690 1050 6810 1060
rect 6940 1050 7060 1060
rect 7190 1050 7310 1060
rect 7440 1050 7560 1060
rect 7690 1050 7810 1060
rect 7940 1050 8000 1060
rect 0 1045 8000 1050
rect 0 1010 75 1045
rect 175 1010 325 1045
rect 425 1010 575 1045
rect 675 1010 825 1045
rect 925 1010 1075 1045
rect 1175 1010 1325 1045
rect 1425 1010 1575 1045
rect 1675 1010 1825 1045
rect 1925 1010 2075 1045
rect 2175 1010 2325 1045
rect 2425 1010 2575 1045
rect 2675 1010 2825 1045
rect 2925 1010 3075 1045
rect 3175 1010 3325 1045
rect 3425 1010 3575 1045
rect 3675 1010 3825 1045
rect 3925 1010 4075 1045
rect 4175 1010 4325 1045
rect 4425 1010 4575 1045
rect 4675 1010 4825 1045
rect 4925 1010 5075 1045
rect 5175 1010 5325 1045
rect 5425 1010 5575 1045
rect 5675 1010 5825 1045
rect 5925 1010 6075 1045
rect 6175 1010 6325 1045
rect 6425 1010 6575 1045
rect 6675 1010 6825 1045
rect 6925 1010 7075 1045
rect 7175 1010 7325 1045
rect 7425 1010 7575 1045
rect 7675 1010 7825 1045
rect 7925 1010 8000 1045
rect 0 990 8000 1010
rect 0 955 75 990
rect 175 955 325 990
rect 425 955 575 990
rect 675 955 825 990
rect 925 955 1075 990
rect 1175 955 1325 990
rect 1425 955 1575 990
rect 1675 955 1825 990
rect 1925 955 2075 990
rect 2175 955 2325 990
rect 2425 955 2575 990
rect 2675 955 2825 990
rect 2925 955 3075 990
rect 3175 955 3325 990
rect 3425 955 3575 990
rect 3675 955 3825 990
rect 3925 955 4075 990
rect 4175 955 4325 990
rect 4425 955 4575 990
rect 4675 955 4825 990
rect 4925 955 5075 990
rect 5175 955 5325 990
rect 5425 955 5575 990
rect 5675 955 5825 990
rect 5925 955 6075 990
rect 6175 955 6325 990
rect 6425 955 6575 990
rect 6675 955 6825 990
rect 6925 955 7075 990
rect 7175 955 7325 990
rect 7425 955 7575 990
rect 7675 955 7825 990
rect 7925 955 8000 990
rect 0 950 8000 955
rect 0 940 60 950
rect 190 940 310 950
rect 440 940 560 950
rect 690 940 810 950
rect 940 940 1060 950
rect 1190 940 1310 950
rect 1440 940 1560 950
rect 1690 940 1810 950
rect 1940 940 2060 950
rect 2190 940 2310 950
rect 2440 940 2560 950
rect 2690 940 2810 950
rect 2940 940 3060 950
rect 3190 940 3310 950
rect 3440 940 3560 950
rect 3690 940 3810 950
rect 3940 940 4060 950
rect 4190 940 4310 950
rect 4440 940 4560 950
rect 4690 940 4810 950
rect 4940 940 5060 950
rect 5190 940 5310 950
rect 5440 940 5560 950
rect 5690 940 5810 950
rect 5940 940 6060 950
rect 6190 940 6310 950
rect 6440 940 6560 950
rect 6690 940 6810 950
rect 6940 940 7060 950
rect 7190 940 7310 950
rect 7440 940 7560 950
rect 7690 940 7810 950
rect 7940 940 8000 950
rect 0 925 50 940
rect 0 825 10 925
rect 45 825 50 925
rect 0 810 50 825
rect 200 925 300 940
rect 200 825 205 925
rect 240 825 260 925
rect 295 825 300 925
rect 200 810 300 825
rect 450 925 550 940
rect 450 825 455 925
rect 490 825 510 925
rect 545 825 550 925
rect 450 810 550 825
rect 700 925 800 940
rect 700 825 705 925
rect 740 825 760 925
rect 795 825 800 925
rect 700 810 800 825
rect 950 925 1050 940
rect 950 825 955 925
rect 990 825 1010 925
rect 1045 825 1050 925
rect 950 810 1050 825
rect 1200 925 1300 940
rect 1200 825 1205 925
rect 1240 825 1260 925
rect 1295 825 1300 925
rect 1200 810 1300 825
rect 1450 925 1550 940
rect 1450 825 1455 925
rect 1490 825 1510 925
rect 1545 825 1550 925
rect 1450 810 1550 825
rect 1700 925 1800 940
rect 1700 825 1705 925
rect 1740 825 1760 925
rect 1795 825 1800 925
rect 1700 810 1800 825
rect 1950 925 2050 940
rect 1950 825 1955 925
rect 1990 825 2010 925
rect 2045 825 2050 925
rect 1950 810 2050 825
rect 2200 925 2300 940
rect 2200 825 2205 925
rect 2240 825 2260 925
rect 2295 825 2300 925
rect 2200 810 2300 825
rect 2450 925 2550 940
rect 2450 825 2455 925
rect 2490 825 2510 925
rect 2545 825 2550 925
rect 2450 810 2550 825
rect 2700 925 2800 940
rect 2700 825 2705 925
rect 2740 825 2760 925
rect 2795 825 2800 925
rect 2700 810 2800 825
rect 2950 925 3050 940
rect 2950 825 2955 925
rect 2990 825 3010 925
rect 3045 825 3050 925
rect 2950 810 3050 825
rect 3200 925 3300 940
rect 3200 825 3205 925
rect 3240 825 3260 925
rect 3295 825 3300 925
rect 3200 810 3300 825
rect 3450 925 3550 940
rect 3450 825 3455 925
rect 3490 825 3510 925
rect 3545 825 3550 925
rect 3450 810 3550 825
rect 3700 925 3800 940
rect 3700 825 3705 925
rect 3740 825 3760 925
rect 3795 825 3800 925
rect 3700 810 3800 825
rect 3950 925 4050 940
rect 3950 825 3955 925
rect 3990 825 4010 925
rect 4045 825 4050 925
rect 3950 810 4050 825
rect 4200 925 4300 940
rect 4200 825 4205 925
rect 4240 825 4260 925
rect 4295 825 4300 925
rect 4200 810 4300 825
rect 4450 925 4550 940
rect 4450 825 4455 925
rect 4490 825 4510 925
rect 4545 825 4550 925
rect 4450 810 4550 825
rect 4700 925 4800 940
rect 4700 825 4705 925
rect 4740 825 4760 925
rect 4795 825 4800 925
rect 4700 810 4800 825
rect 4950 925 5050 940
rect 4950 825 4955 925
rect 4990 825 5010 925
rect 5045 825 5050 925
rect 4950 810 5050 825
rect 5200 925 5300 940
rect 5200 825 5205 925
rect 5240 825 5260 925
rect 5295 825 5300 925
rect 5200 810 5300 825
rect 5450 925 5550 940
rect 5450 825 5455 925
rect 5490 825 5510 925
rect 5545 825 5550 925
rect 5450 810 5550 825
rect 5700 925 5800 940
rect 5700 825 5705 925
rect 5740 825 5760 925
rect 5795 825 5800 925
rect 5700 810 5800 825
rect 5950 925 6050 940
rect 5950 825 5955 925
rect 5990 825 6010 925
rect 6045 825 6050 925
rect 5950 810 6050 825
rect 6200 925 6300 940
rect 6200 825 6205 925
rect 6240 825 6260 925
rect 6295 825 6300 925
rect 6200 810 6300 825
rect 6450 925 6550 940
rect 6450 825 6455 925
rect 6490 825 6510 925
rect 6545 825 6550 925
rect 6450 810 6550 825
rect 6700 925 6800 940
rect 6700 825 6705 925
rect 6740 825 6760 925
rect 6795 825 6800 925
rect 6700 810 6800 825
rect 6950 925 7050 940
rect 6950 825 6955 925
rect 6990 825 7010 925
rect 7045 825 7050 925
rect 6950 810 7050 825
rect 7200 925 7300 940
rect 7200 825 7205 925
rect 7240 825 7260 925
rect 7295 825 7300 925
rect 7200 810 7300 825
rect 7450 925 7550 940
rect 7450 825 7455 925
rect 7490 825 7510 925
rect 7545 825 7550 925
rect 7450 810 7550 825
rect 7700 925 7800 940
rect 7700 825 7705 925
rect 7740 825 7760 925
rect 7795 825 7800 925
rect 7700 810 7800 825
rect 7950 925 8000 940
rect 7950 825 7955 925
rect 7990 825 8000 925
rect 7950 810 8000 825
rect 0 800 60 810
rect 190 800 310 810
rect 440 800 560 810
rect 690 800 810 810
rect 940 800 1060 810
rect 1190 800 1310 810
rect 1440 800 1560 810
rect 1690 800 1810 810
rect 1940 800 2060 810
rect 2190 800 2310 810
rect 2440 800 2560 810
rect 2690 800 2810 810
rect 2940 800 3060 810
rect 3190 800 3310 810
rect 3440 800 3560 810
rect 3690 800 3810 810
rect 3940 800 4060 810
rect 4190 800 4310 810
rect 4440 800 4560 810
rect 4690 800 4810 810
rect 4940 800 5060 810
rect 5190 800 5310 810
rect 5440 800 5560 810
rect 5690 800 5810 810
rect 5940 800 6060 810
rect 6190 800 6310 810
rect 6440 800 6560 810
rect 6690 800 6810 810
rect 6940 800 7060 810
rect 7190 800 7310 810
rect 7440 800 7560 810
rect 7690 800 7810 810
rect 7940 800 8000 810
rect 0 795 8000 800
rect 0 760 75 795
rect 175 760 325 795
rect 425 760 575 795
rect 675 760 825 795
rect 925 760 1075 795
rect 1175 760 1325 795
rect 1425 760 1575 795
rect 1675 760 1825 795
rect 1925 760 2075 795
rect 2175 760 2325 795
rect 2425 760 2575 795
rect 2675 760 2825 795
rect 2925 760 3075 795
rect 3175 760 3325 795
rect 3425 760 3575 795
rect 3675 760 3825 795
rect 3925 760 4075 795
rect 4175 760 4325 795
rect 4425 760 4575 795
rect 4675 760 4825 795
rect 4925 760 5075 795
rect 5175 760 5325 795
rect 5425 760 5575 795
rect 5675 760 5825 795
rect 5925 760 6075 795
rect 6175 760 6325 795
rect 6425 760 6575 795
rect 6675 760 6825 795
rect 6925 760 7075 795
rect 7175 760 7325 795
rect 7425 760 7575 795
rect 7675 760 7825 795
rect 7925 760 8000 795
rect 0 740 8000 760
rect 0 705 75 740
rect 175 705 325 740
rect 425 705 575 740
rect 675 705 825 740
rect 925 705 1075 740
rect 1175 705 1325 740
rect 1425 705 1575 740
rect 1675 705 1825 740
rect 1925 705 2075 740
rect 2175 705 2325 740
rect 2425 705 2575 740
rect 2675 705 2825 740
rect 2925 705 3075 740
rect 3175 705 3325 740
rect 3425 705 3575 740
rect 3675 705 3825 740
rect 3925 705 4075 740
rect 4175 705 4325 740
rect 4425 705 4575 740
rect 4675 705 4825 740
rect 4925 705 5075 740
rect 5175 705 5325 740
rect 5425 705 5575 740
rect 5675 705 5825 740
rect 5925 705 6075 740
rect 6175 705 6325 740
rect 6425 705 6575 740
rect 6675 705 6825 740
rect 6925 705 7075 740
rect 7175 705 7325 740
rect 7425 705 7575 740
rect 7675 705 7825 740
rect 7925 705 8000 740
rect 0 700 8000 705
rect 0 690 60 700
rect 190 690 310 700
rect 440 690 560 700
rect 690 690 810 700
rect 940 690 1060 700
rect 1190 690 1310 700
rect 1440 690 1560 700
rect 1690 690 1810 700
rect 1940 690 2060 700
rect 2190 690 2310 700
rect 2440 690 2560 700
rect 2690 690 2810 700
rect 2940 690 3060 700
rect 3190 690 3310 700
rect 3440 690 3560 700
rect 3690 690 3810 700
rect 3940 690 4060 700
rect 4190 690 4310 700
rect 4440 690 4560 700
rect 4690 690 4810 700
rect 4940 690 5060 700
rect 5190 690 5310 700
rect 5440 690 5560 700
rect 5690 690 5810 700
rect 5940 690 6060 700
rect 6190 690 6310 700
rect 6440 690 6560 700
rect 6690 690 6810 700
rect 6940 690 7060 700
rect 7190 690 7310 700
rect 7440 690 7560 700
rect 7690 690 7810 700
rect 7940 690 8000 700
rect 0 675 50 690
rect 0 575 10 675
rect 45 575 50 675
rect 0 560 50 575
rect 200 675 300 690
rect 200 575 205 675
rect 240 575 260 675
rect 295 575 300 675
rect 200 560 300 575
rect 450 675 550 690
rect 450 575 455 675
rect 490 575 510 675
rect 545 575 550 675
rect 450 560 550 575
rect 700 675 800 690
rect 700 575 705 675
rect 740 575 760 675
rect 795 575 800 675
rect 700 560 800 575
rect 950 675 1050 690
rect 950 575 955 675
rect 990 575 1010 675
rect 1045 575 1050 675
rect 950 560 1050 575
rect 1200 675 1300 690
rect 1200 575 1205 675
rect 1240 575 1260 675
rect 1295 575 1300 675
rect 1200 560 1300 575
rect 1450 675 1550 690
rect 1450 575 1455 675
rect 1490 575 1510 675
rect 1545 575 1550 675
rect 1450 560 1550 575
rect 1700 675 1800 690
rect 1700 575 1705 675
rect 1740 575 1760 675
rect 1795 575 1800 675
rect 1700 560 1800 575
rect 1950 675 2050 690
rect 1950 575 1955 675
rect 1990 575 2010 675
rect 2045 575 2050 675
rect 1950 560 2050 575
rect 2200 675 2300 690
rect 2200 575 2205 675
rect 2240 575 2260 675
rect 2295 575 2300 675
rect 2200 560 2300 575
rect 2450 675 2550 690
rect 2450 575 2455 675
rect 2490 575 2510 675
rect 2545 575 2550 675
rect 2450 560 2550 575
rect 2700 675 2800 690
rect 2700 575 2705 675
rect 2740 575 2760 675
rect 2795 575 2800 675
rect 2700 560 2800 575
rect 2950 675 3050 690
rect 2950 575 2955 675
rect 2990 575 3010 675
rect 3045 575 3050 675
rect 2950 560 3050 575
rect 3200 675 3300 690
rect 3200 575 3205 675
rect 3240 575 3260 675
rect 3295 575 3300 675
rect 3200 560 3300 575
rect 3450 675 3550 690
rect 3450 575 3455 675
rect 3490 575 3510 675
rect 3545 575 3550 675
rect 3450 560 3550 575
rect 3700 675 3800 690
rect 3700 575 3705 675
rect 3740 575 3760 675
rect 3795 575 3800 675
rect 3700 560 3800 575
rect 3950 675 4050 690
rect 3950 575 3955 675
rect 3990 575 4010 675
rect 4045 575 4050 675
rect 3950 560 4050 575
rect 4200 675 4300 690
rect 4200 575 4205 675
rect 4240 575 4260 675
rect 4295 575 4300 675
rect 4200 560 4300 575
rect 4450 675 4550 690
rect 4450 575 4455 675
rect 4490 575 4510 675
rect 4545 575 4550 675
rect 4450 560 4550 575
rect 4700 675 4800 690
rect 4700 575 4705 675
rect 4740 575 4760 675
rect 4795 575 4800 675
rect 4700 560 4800 575
rect 4950 675 5050 690
rect 4950 575 4955 675
rect 4990 575 5010 675
rect 5045 575 5050 675
rect 4950 560 5050 575
rect 5200 675 5300 690
rect 5200 575 5205 675
rect 5240 575 5260 675
rect 5295 575 5300 675
rect 5200 560 5300 575
rect 5450 675 5550 690
rect 5450 575 5455 675
rect 5490 575 5510 675
rect 5545 575 5550 675
rect 5450 560 5550 575
rect 5700 675 5800 690
rect 5700 575 5705 675
rect 5740 575 5760 675
rect 5795 575 5800 675
rect 5700 560 5800 575
rect 5950 675 6050 690
rect 5950 575 5955 675
rect 5990 575 6010 675
rect 6045 575 6050 675
rect 5950 560 6050 575
rect 6200 675 6300 690
rect 6200 575 6205 675
rect 6240 575 6260 675
rect 6295 575 6300 675
rect 6200 560 6300 575
rect 6450 675 6550 690
rect 6450 575 6455 675
rect 6490 575 6510 675
rect 6545 575 6550 675
rect 6450 560 6550 575
rect 6700 675 6800 690
rect 6700 575 6705 675
rect 6740 575 6760 675
rect 6795 575 6800 675
rect 6700 560 6800 575
rect 6950 675 7050 690
rect 6950 575 6955 675
rect 6990 575 7010 675
rect 7045 575 7050 675
rect 6950 560 7050 575
rect 7200 675 7300 690
rect 7200 575 7205 675
rect 7240 575 7260 675
rect 7295 575 7300 675
rect 7200 560 7300 575
rect 7450 675 7550 690
rect 7450 575 7455 675
rect 7490 575 7510 675
rect 7545 575 7550 675
rect 7450 560 7550 575
rect 7700 675 7800 690
rect 7700 575 7705 675
rect 7740 575 7760 675
rect 7795 575 7800 675
rect 7700 560 7800 575
rect 7950 675 8000 690
rect 7950 575 7955 675
rect 7990 575 8000 675
rect 7950 560 8000 575
rect 0 550 60 560
rect 190 550 310 560
rect 440 550 560 560
rect 690 550 810 560
rect 940 550 1060 560
rect 1190 550 1310 560
rect 1440 550 1560 560
rect 1690 550 1810 560
rect 1940 550 2060 560
rect 2190 550 2310 560
rect 2440 550 2560 560
rect 2690 550 2810 560
rect 2940 550 3060 560
rect 3190 550 3310 560
rect 3440 550 3560 560
rect 3690 550 3810 560
rect 3940 550 4060 560
rect 4190 550 4310 560
rect 4440 550 4560 560
rect 4690 550 4810 560
rect 4940 550 5060 560
rect 5190 550 5310 560
rect 5440 550 5560 560
rect 5690 550 5810 560
rect 5940 550 6060 560
rect 6190 550 6310 560
rect 6440 550 6560 560
rect 6690 550 6810 560
rect 6940 550 7060 560
rect 7190 550 7310 560
rect 7440 550 7560 560
rect 7690 550 7810 560
rect 7940 550 8000 560
rect 0 545 8000 550
rect 0 510 75 545
rect 175 510 325 545
rect 425 510 575 545
rect 675 510 825 545
rect 925 510 1075 545
rect 1175 510 1325 545
rect 1425 510 1575 545
rect 1675 510 1825 545
rect 1925 510 2075 545
rect 2175 510 2325 545
rect 2425 510 2575 545
rect 2675 510 2825 545
rect 2925 510 3075 545
rect 3175 510 3325 545
rect 3425 510 3575 545
rect 3675 510 3825 545
rect 3925 510 4075 545
rect 4175 510 4325 545
rect 4425 510 4575 545
rect 4675 510 4825 545
rect 4925 510 5075 545
rect 5175 510 5325 545
rect 5425 510 5575 545
rect 5675 510 5825 545
rect 5925 510 6075 545
rect 6175 510 6325 545
rect 6425 510 6575 545
rect 6675 510 6825 545
rect 6925 510 7075 545
rect 7175 510 7325 545
rect 7425 510 7575 545
rect 7675 510 7825 545
rect 7925 510 8000 545
rect 0 490 8000 510
rect 0 455 75 490
rect 175 455 325 490
rect 425 455 575 490
rect 675 455 825 490
rect 925 455 1075 490
rect 1175 455 1325 490
rect 1425 455 1575 490
rect 1675 455 1825 490
rect 1925 455 2075 490
rect 2175 455 2325 490
rect 2425 455 2575 490
rect 2675 455 2825 490
rect 2925 455 3075 490
rect 3175 455 3325 490
rect 3425 455 3575 490
rect 3675 455 3825 490
rect 3925 455 4075 490
rect 4175 455 4325 490
rect 4425 455 4575 490
rect 4675 455 4825 490
rect 4925 455 5075 490
rect 5175 455 5325 490
rect 5425 455 5575 490
rect 5675 455 5825 490
rect 5925 455 6075 490
rect 6175 455 6325 490
rect 6425 455 6575 490
rect 6675 455 6825 490
rect 6925 455 7075 490
rect 7175 455 7325 490
rect 7425 455 7575 490
rect 7675 455 7825 490
rect 7925 455 8000 490
rect 0 450 8000 455
rect 0 440 60 450
rect 190 440 310 450
rect 440 440 560 450
rect 690 440 810 450
rect 940 440 1060 450
rect 1190 440 1310 450
rect 1440 440 1560 450
rect 1690 440 1810 450
rect 1940 440 2060 450
rect 2190 440 2310 450
rect 2440 440 2560 450
rect 2690 440 2810 450
rect 2940 440 3060 450
rect 3190 440 3310 450
rect 3440 440 3560 450
rect 3690 440 3810 450
rect 3940 440 4060 450
rect 4190 440 4310 450
rect 4440 440 4560 450
rect 4690 440 4810 450
rect 4940 440 5060 450
rect 5190 440 5310 450
rect 5440 440 5560 450
rect 5690 440 5810 450
rect 5940 440 6060 450
rect 6190 440 6310 450
rect 6440 440 6560 450
rect 6690 440 6810 450
rect 6940 440 7060 450
rect 7190 440 7310 450
rect 7440 440 7560 450
rect 7690 440 7810 450
rect 7940 440 8000 450
rect 0 425 50 440
rect 0 325 10 425
rect 45 325 50 425
rect 0 310 50 325
rect 200 425 300 440
rect 200 325 205 425
rect 240 325 260 425
rect 295 325 300 425
rect 200 310 300 325
rect 450 425 550 440
rect 450 325 455 425
rect 490 325 510 425
rect 545 325 550 425
rect 450 310 550 325
rect 700 425 800 440
rect 700 325 705 425
rect 740 325 760 425
rect 795 325 800 425
rect 700 310 800 325
rect 950 425 1050 440
rect 950 325 955 425
rect 990 325 1010 425
rect 1045 325 1050 425
rect 950 310 1050 325
rect 1200 425 1300 440
rect 1200 325 1205 425
rect 1240 325 1260 425
rect 1295 325 1300 425
rect 1200 310 1300 325
rect 1450 425 1550 440
rect 1450 325 1455 425
rect 1490 325 1510 425
rect 1545 325 1550 425
rect 1450 310 1550 325
rect 1700 425 1800 440
rect 1700 325 1705 425
rect 1740 325 1760 425
rect 1795 325 1800 425
rect 1700 310 1800 325
rect 1950 425 2050 440
rect 1950 325 1955 425
rect 1990 325 2010 425
rect 2045 325 2050 425
rect 1950 310 2050 325
rect 2200 425 2300 440
rect 2200 325 2205 425
rect 2240 325 2260 425
rect 2295 325 2300 425
rect 2200 310 2300 325
rect 2450 425 2550 440
rect 2450 325 2455 425
rect 2490 325 2510 425
rect 2545 325 2550 425
rect 2450 310 2550 325
rect 2700 425 2800 440
rect 2700 325 2705 425
rect 2740 325 2760 425
rect 2795 325 2800 425
rect 2700 310 2800 325
rect 2950 425 3050 440
rect 2950 325 2955 425
rect 2990 325 3010 425
rect 3045 325 3050 425
rect 2950 310 3050 325
rect 3200 425 3300 440
rect 3200 325 3205 425
rect 3240 325 3260 425
rect 3295 325 3300 425
rect 3200 310 3300 325
rect 3450 425 3550 440
rect 3450 325 3455 425
rect 3490 325 3510 425
rect 3545 325 3550 425
rect 3450 310 3550 325
rect 3700 425 3800 440
rect 3700 325 3705 425
rect 3740 325 3760 425
rect 3795 325 3800 425
rect 3700 310 3800 325
rect 3950 425 4050 440
rect 3950 325 3955 425
rect 3990 325 4010 425
rect 4045 325 4050 425
rect 3950 310 4050 325
rect 4200 425 4300 440
rect 4200 325 4205 425
rect 4240 325 4260 425
rect 4295 325 4300 425
rect 4200 310 4300 325
rect 4450 425 4550 440
rect 4450 325 4455 425
rect 4490 325 4510 425
rect 4545 325 4550 425
rect 4450 310 4550 325
rect 4700 425 4800 440
rect 4700 325 4705 425
rect 4740 325 4760 425
rect 4795 325 4800 425
rect 4700 310 4800 325
rect 4950 425 5050 440
rect 4950 325 4955 425
rect 4990 325 5010 425
rect 5045 325 5050 425
rect 4950 310 5050 325
rect 5200 425 5300 440
rect 5200 325 5205 425
rect 5240 325 5260 425
rect 5295 325 5300 425
rect 5200 310 5300 325
rect 5450 425 5550 440
rect 5450 325 5455 425
rect 5490 325 5510 425
rect 5545 325 5550 425
rect 5450 310 5550 325
rect 5700 425 5800 440
rect 5700 325 5705 425
rect 5740 325 5760 425
rect 5795 325 5800 425
rect 5700 310 5800 325
rect 5950 425 6050 440
rect 5950 325 5955 425
rect 5990 325 6010 425
rect 6045 325 6050 425
rect 5950 310 6050 325
rect 6200 425 6300 440
rect 6200 325 6205 425
rect 6240 325 6260 425
rect 6295 325 6300 425
rect 6200 310 6300 325
rect 6450 425 6550 440
rect 6450 325 6455 425
rect 6490 325 6510 425
rect 6545 325 6550 425
rect 6450 310 6550 325
rect 6700 425 6800 440
rect 6700 325 6705 425
rect 6740 325 6760 425
rect 6795 325 6800 425
rect 6700 310 6800 325
rect 6950 425 7050 440
rect 6950 325 6955 425
rect 6990 325 7010 425
rect 7045 325 7050 425
rect 6950 310 7050 325
rect 7200 425 7300 440
rect 7200 325 7205 425
rect 7240 325 7260 425
rect 7295 325 7300 425
rect 7200 310 7300 325
rect 7450 425 7550 440
rect 7450 325 7455 425
rect 7490 325 7510 425
rect 7545 325 7550 425
rect 7450 310 7550 325
rect 7700 425 7800 440
rect 7700 325 7705 425
rect 7740 325 7760 425
rect 7795 325 7800 425
rect 7700 310 7800 325
rect 7950 425 8000 440
rect 7950 325 7955 425
rect 7990 325 8000 425
rect 7950 310 8000 325
rect 0 300 60 310
rect 190 300 310 310
rect 440 300 560 310
rect 690 300 810 310
rect 940 300 1060 310
rect 1190 300 1310 310
rect 1440 300 1560 310
rect 1690 300 1810 310
rect 1940 300 2060 310
rect 2190 300 2310 310
rect 2440 300 2560 310
rect 2690 300 2810 310
rect 2940 300 3060 310
rect 3190 300 3310 310
rect 3440 300 3560 310
rect 3690 300 3810 310
rect 3940 300 4060 310
rect 4190 300 4310 310
rect 4440 300 4560 310
rect 4690 300 4810 310
rect 4940 300 5060 310
rect 5190 300 5310 310
rect 5440 300 5560 310
rect 5690 300 5810 310
rect 5940 300 6060 310
rect 6190 300 6310 310
rect 6440 300 6560 310
rect 6690 300 6810 310
rect 6940 300 7060 310
rect 7190 300 7310 310
rect 7440 300 7560 310
rect 7690 300 7810 310
rect 7940 300 8000 310
rect 0 295 8000 300
rect 0 260 75 295
rect 175 260 325 295
rect 425 260 575 295
rect 675 260 825 295
rect 925 260 1075 295
rect 1175 260 1325 295
rect 1425 260 1575 295
rect 1675 260 1825 295
rect 1925 260 2075 295
rect 2175 260 2325 295
rect 2425 260 2575 295
rect 2675 260 2825 295
rect 2925 260 3075 295
rect 3175 260 3325 295
rect 3425 260 3575 295
rect 3675 260 3825 295
rect 3925 260 4075 295
rect 4175 260 4325 295
rect 4425 260 4575 295
rect 4675 260 4825 295
rect 4925 260 5075 295
rect 5175 260 5325 295
rect 5425 260 5575 295
rect 5675 260 5825 295
rect 5925 260 6075 295
rect 6175 260 6325 295
rect 6425 260 6575 295
rect 6675 260 6825 295
rect 6925 260 7075 295
rect 7175 260 7325 295
rect 7425 260 7575 295
rect 7675 260 7825 295
rect 7925 260 8000 295
rect 0 240 8000 260
rect 0 205 75 240
rect 175 205 325 240
rect 425 205 575 240
rect 675 205 825 240
rect 925 205 1075 240
rect 1175 205 1325 240
rect 1425 205 1575 240
rect 1675 205 1825 240
rect 1925 205 2075 240
rect 2175 205 2325 240
rect 2425 205 2575 240
rect 2675 205 2825 240
rect 2925 205 3075 240
rect 3175 205 3325 240
rect 3425 205 3575 240
rect 3675 205 3825 240
rect 3925 205 4075 240
rect 4175 205 4325 240
rect 4425 205 4575 240
rect 4675 205 4825 240
rect 4925 205 5075 240
rect 5175 205 5325 240
rect 5425 205 5575 240
rect 5675 205 5825 240
rect 5925 205 6075 240
rect 6175 205 6325 240
rect 6425 205 6575 240
rect 6675 205 6825 240
rect 6925 205 7075 240
rect 7175 205 7325 240
rect 7425 205 7575 240
rect 7675 205 7825 240
rect 7925 205 8000 240
rect 0 200 8000 205
rect 0 190 60 200
rect 190 190 310 200
rect 440 190 560 200
rect 690 190 810 200
rect 940 190 1060 200
rect 1190 190 1310 200
rect 1440 190 1560 200
rect 1690 190 1810 200
rect 1940 190 2060 200
rect 2190 190 2310 200
rect 2440 190 2560 200
rect 2690 190 2810 200
rect 2940 190 3060 200
rect 3190 190 3310 200
rect 3440 190 3560 200
rect 3690 190 3810 200
rect 3940 190 4060 200
rect 4190 190 4310 200
rect 4440 190 4560 200
rect 4690 190 4810 200
rect 4940 190 5060 200
rect 5190 190 5310 200
rect 5440 190 5560 200
rect 5690 190 5810 200
rect 5940 190 6060 200
rect 6190 190 6310 200
rect 6440 190 6560 200
rect 6690 190 6810 200
rect 6940 190 7060 200
rect 7190 190 7310 200
rect 7440 190 7560 200
rect 7690 190 7810 200
rect 7940 190 8000 200
rect 0 175 50 190
rect 0 75 10 175
rect 45 75 50 175
rect 0 60 50 75
rect 200 175 300 190
rect 200 75 205 175
rect 240 75 260 175
rect 295 75 300 175
rect 200 60 300 75
rect 450 175 550 190
rect 450 75 455 175
rect 490 75 510 175
rect 545 75 550 175
rect 450 60 550 75
rect 700 175 800 190
rect 700 75 705 175
rect 740 75 760 175
rect 795 75 800 175
rect 700 60 800 75
rect 950 175 1050 190
rect 950 75 955 175
rect 990 75 1010 175
rect 1045 75 1050 175
rect 950 60 1050 75
rect 1200 175 1300 190
rect 1200 75 1205 175
rect 1240 75 1260 175
rect 1295 75 1300 175
rect 1200 60 1300 75
rect 1450 175 1550 190
rect 1450 75 1455 175
rect 1490 75 1510 175
rect 1545 75 1550 175
rect 1450 60 1550 75
rect 1700 175 1800 190
rect 1700 75 1705 175
rect 1740 75 1760 175
rect 1795 75 1800 175
rect 1700 60 1800 75
rect 1950 175 2050 190
rect 1950 75 1955 175
rect 1990 75 2010 175
rect 2045 75 2050 175
rect 1950 60 2050 75
rect 2200 175 2300 190
rect 2200 75 2205 175
rect 2240 75 2260 175
rect 2295 75 2300 175
rect 2200 60 2300 75
rect 2450 175 2550 190
rect 2450 75 2455 175
rect 2490 75 2510 175
rect 2545 75 2550 175
rect 2450 60 2550 75
rect 2700 175 2800 190
rect 2700 75 2705 175
rect 2740 75 2760 175
rect 2795 75 2800 175
rect 2700 60 2800 75
rect 2950 175 3050 190
rect 2950 75 2955 175
rect 2990 75 3010 175
rect 3045 75 3050 175
rect 2950 60 3050 75
rect 3200 175 3300 190
rect 3200 75 3205 175
rect 3240 75 3260 175
rect 3295 75 3300 175
rect 3200 60 3300 75
rect 3450 175 3550 190
rect 3450 75 3455 175
rect 3490 75 3510 175
rect 3545 75 3550 175
rect 3450 60 3550 75
rect 3700 175 3800 190
rect 3700 75 3705 175
rect 3740 75 3760 175
rect 3795 75 3800 175
rect 3700 60 3800 75
rect 3950 175 4050 190
rect 3950 75 3955 175
rect 3990 75 4010 175
rect 4045 75 4050 175
rect 3950 60 4050 75
rect 4200 175 4300 190
rect 4200 75 4205 175
rect 4240 75 4260 175
rect 4295 75 4300 175
rect 4200 60 4300 75
rect 4450 175 4550 190
rect 4450 75 4455 175
rect 4490 75 4510 175
rect 4545 75 4550 175
rect 4450 60 4550 75
rect 4700 175 4800 190
rect 4700 75 4705 175
rect 4740 75 4760 175
rect 4795 75 4800 175
rect 4700 60 4800 75
rect 4950 175 5050 190
rect 4950 75 4955 175
rect 4990 75 5010 175
rect 5045 75 5050 175
rect 4950 60 5050 75
rect 5200 175 5300 190
rect 5200 75 5205 175
rect 5240 75 5260 175
rect 5295 75 5300 175
rect 5200 60 5300 75
rect 5450 175 5550 190
rect 5450 75 5455 175
rect 5490 75 5510 175
rect 5545 75 5550 175
rect 5450 60 5550 75
rect 5700 175 5800 190
rect 5700 75 5705 175
rect 5740 75 5760 175
rect 5795 75 5800 175
rect 5700 60 5800 75
rect 5950 175 6050 190
rect 5950 75 5955 175
rect 5990 75 6010 175
rect 6045 75 6050 175
rect 5950 60 6050 75
rect 6200 175 6300 190
rect 6200 75 6205 175
rect 6240 75 6260 175
rect 6295 75 6300 175
rect 6200 60 6300 75
rect 6450 175 6550 190
rect 6450 75 6455 175
rect 6490 75 6510 175
rect 6545 75 6550 175
rect 6450 60 6550 75
rect 6700 175 6800 190
rect 6700 75 6705 175
rect 6740 75 6760 175
rect 6795 75 6800 175
rect 6700 60 6800 75
rect 6950 175 7050 190
rect 6950 75 6955 175
rect 6990 75 7010 175
rect 7045 75 7050 175
rect 6950 60 7050 75
rect 7200 175 7300 190
rect 7200 75 7205 175
rect 7240 75 7260 175
rect 7295 75 7300 175
rect 7200 60 7300 75
rect 7450 175 7550 190
rect 7450 75 7455 175
rect 7490 75 7510 175
rect 7545 75 7550 175
rect 7450 60 7550 75
rect 7700 175 7800 190
rect 7700 75 7705 175
rect 7740 75 7760 175
rect 7795 75 7800 175
rect 7700 60 7800 75
rect 7950 175 8000 190
rect 7950 75 7955 175
rect 7990 75 8000 175
rect 7950 60 8000 75
rect 0 50 60 60
rect 190 50 310 60
rect 440 50 560 60
rect 690 50 810 60
rect 940 50 1060 60
rect 1190 50 1310 60
rect 1440 50 1560 60
rect 1690 50 1810 60
rect 1940 50 2060 60
rect 2190 50 2310 60
rect 2440 50 2560 60
rect 2690 50 2810 60
rect 2940 50 3060 60
rect 3190 50 3310 60
rect 3440 50 3560 60
rect 3690 50 3810 60
rect 3940 50 4060 60
rect 4190 50 4310 60
rect 4440 50 4560 60
rect 4690 50 4810 60
rect 4940 50 5060 60
rect 5190 50 5310 60
rect 5440 50 5560 60
rect 5690 50 5810 60
rect 5940 50 6060 60
rect 6190 50 6310 60
rect 6440 50 6560 60
rect 6690 50 6810 60
rect 6940 50 7060 60
rect 7190 50 7310 60
rect 7440 50 7560 60
rect 7690 50 7810 60
rect 7940 50 8000 60
rect 0 45 8000 50
rect 0 10 75 45
rect 175 10 325 45
rect 425 10 575 45
rect 675 10 825 45
rect 925 10 1075 45
rect 1175 10 1325 45
rect 1425 10 1575 45
rect 1675 10 1825 45
rect 1925 10 2075 45
rect 2175 10 2325 45
rect 2425 10 2575 45
rect 2675 10 2825 45
rect 2925 10 3075 45
rect 3175 10 3325 45
rect 3425 10 3575 45
rect 3675 10 3825 45
rect 3925 10 4075 45
rect 4175 10 4325 45
rect 4425 10 4575 45
rect 4675 10 4825 45
rect 4925 10 5075 45
rect 5175 10 5325 45
rect 5425 10 5575 45
rect 5675 10 5825 45
rect 5925 10 6075 45
rect 6175 10 6325 45
rect 6425 10 6575 45
rect 6675 10 6825 45
rect 6925 10 7075 45
rect 7175 10 7325 45
rect 7425 10 7575 45
rect 7675 10 7825 45
rect 7925 10 8000 45
rect 0 0 8000 10
<< via1 >>
rect 75 7955 175 7990
rect 325 7955 425 7990
rect 575 7955 675 7990
rect 825 7955 925 7990
rect 1075 7955 1175 7990
rect 1325 7955 1425 7990
rect 1575 7955 1675 7990
rect 1825 7955 1925 7990
rect 2075 7955 2175 7990
rect 2325 7955 2425 7990
rect 2575 7955 2675 7990
rect 2825 7955 2925 7990
rect 3075 7955 3175 7990
rect 3325 7955 3425 7990
rect 3575 7955 3675 7990
rect 3825 7955 3925 7990
rect 4075 7955 4175 7990
rect 4325 7955 4425 7990
rect 4575 7955 4675 7990
rect 4825 7955 4925 7990
rect 5075 7955 5175 7990
rect 5325 7955 5425 7990
rect 5575 7955 5675 7990
rect 5825 7955 5925 7990
rect 6075 7955 6175 7990
rect 6325 7955 6425 7990
rect 6575 7955 6675 7990
rect 6825 7955 6925 7990
rect 7075 7955 7175 7990
rect 7325 7955 7425 7990
rect 7575 7955 7675 7990
rect 7825 7955 7925 7990
rect 10 7825 45 7925
rect 205 7825 240 7925
rect 260 7825 295 7925
rect 455 7825 490 7925
rect 510 7825 545 7925
rect 705 7825 740 7925
rect 760 7825 795 7925
rect 955 7825 990 7925
rect 1010 7825 1045 7925
rect 1205 7825 1240 7925
rect 1260 7825 1295 7925
rect 1455 7825 1490 7925
rect 1510 7825 1545 7925
rect 1705 7825 1740 7925
rect 1760 7825 1795 7925
rect 1955 7825 1990 7925
rect 2010 7825 2045 7925
rect 2205 7825 2240 7925
rect 2260 7825 2295 7925
rect 2455 7825 2490 7925
rect 2510 7825 2545 7925
rect 2705 7825 2740 7925
rect 2760 7825 2795 7925
rect 2955 7825 2990 7925
rect 3010 7825 3045 7925
rect 3205 7825 3240 7925
rect 3260 7825 3295 7925
rect 3455 7825 3490 7925
rect 3510 7825 3545 7925
rect 3705 7825 3740 7925
rect 3760 7825 3795 7925
rect 3955 7825 3990 7925
rect 4010 7825 4045 7925
rect 4205 7825 4240 7925
rect 4260 7825 4295 7925
rect 4455 7825 4490 7925
rect 4510 7825 4545 7925
rect 4705 7825 4740 7925
rect 4760 7825 4795 7925
rect 4955 7825 4990 7925
rect 5010 7825 5045 7925
rect 5205 7825 5240 7925
rect 5260 7825 5295 7925
rect 5455 7825 5490 7925
rect 5510 7825 5545 7925
rect 5705 7825 5740 7925
rect 5760 7825 5795 7925
rect 5955 7825 5990 7925
rect 6010 7825 6045 7925
rect 6205 7825 6240 7925
rect 6260 7825 6295 7925
rect 6455 7825 6490 7925
rect 6510 7825 6545 7925
rect 6705 7825 6740 7925
rect 6760 7825 6795 7925
rect 6955 7825 6990 7925
rect 7010 7825 7045 7925
rect 7205 7825 7240 7925
rect 7260 7825 7295 7925
rect 7455 7825 7490 7925
rect 7510 7825 7545 7925
rect 7705 7825 7740 7925
rect 7760 7825 7795 7925
rect 7955 7825 7990 7925
rect 75 7760 175 7795
rect 325 7760 425 7795
rect 575 7760 675 7795
rect 825 7760 925 7795
rect 1075 7760 1175 7795
rect 1325 7760 1425 7795
rect 1575 7760 1675 7795
rect 1825 7760 1925 7795
rect 2075 7760 2175 7795
rect 2325 7760 2425 7795
rect 2575 7760 2675 7795
rect 2825 7760 2925 7795
rect 3075 7760 3175 7795
rect 3325 7760 3425 7795
rect 3575 7760 3675 7795
rect 3825 7760 3925 7795
rect 4075 7760 4175 7795
rect 4325 7760 4425 7795
rect 4575 7760 4675 7795
rect 4825 7760 4925 7795
rect 5075 7760 5175 7795
rect 5325 7760 5425 7795
rect 5575 7760 5675 7795
rect 5825 7760 5925 7795
rect 6075 7760 6175 7795
rect 6325 7760 6425 7795
rect 6575 7760 6675 7795
rect 6825 7760 6925 7795
rect 7075 7760 7175 7795
rect 7325 7760 7425 7795
rect 7575 7760 7675 7795
rect 7825 7760 7925 7795
rect 75 7705 175 7740
rect 325 7705 425 7740
rect 575 7705 675 7740
rect 825 7705 925 7740
rect 1075 7705 1175 7740
rect 1325 7705 1425 7740
rect 1575 7705 1675 7740
rect 1825 7705 1925 7740
rect 2075 7705 2175 7740
rect 2325 7705 2425 7740
rect 2575 7705 2675 7740
rect 2825 7705 2925 7740
rect 3075 7705 3175 7740
rect 3325 7705 3425 7740
rect 3575 7705 3675 7740
rect 3825 7705 3925 7740
rect 4075 7705 4175 7740
rect 4325 7705 4425 7740
rect 4575 7705 4675 7740
rect 4825 7705 4925 7740
rect 5075 7705 5175 7740
rect 5325 7705 5425 7740
rect 5575 7705 5675 7740
rect 5825 7705 5925 7740
rect 6075 7705 6175 7740
rect 6325 7705 6425 7740
rect 6575 7705 6675 7740
rect 6825 7705 6925 7740
rect 7075 7705 7175 7740
rect 7325 7705 7425 7740
rect 7575 7705 7675 7740
rect 7825 7705 7925 7740
rect 10 7575 45 7675
rect 205 7575 240 7675
rect 260 7575 295 7675
rect 455 7575 490 7675
rect 510 7575 545 7675
rect 705 7575 740 7675
rect 760 7575 795 7675
rect 955 7575 990 7675
rect 1010 7575 1045 7675
rect 1205 7575 1240 7675
rect 1260 7575 1295 7675
rect 1455 7575 1490 7675
rect 1510 7575 1545 7675
rect 1705 7575 1740 7675
rect 1760 7575 1795 7675
rect 1955 7575 1990 7675
rect 2010 7575 2045 7675
rect 2205 7575 2240 7675
rect 2260 7575 2295 7675
rect 2455 7575 2490 7675
rect 2510 7575 2545 7675
rect 2705 7575 2740 7675
rect 2760 7575 2795 7675
rect 2955 7575 2990 7675
rect 3010 7575 3045 7675
rect 3205 7575 3240 7675
rect 3260 7575 3295 7675
rect 3455 7575 3490 7675
rect 3510 7575 3545 7675
rect 3705 7575 3740 7675
rect 3760 7575 3795 7675
rect 3955 7575 3990 7675
rect 4010 7575 4045 7675
rect 4205 7575 4240 7675
rect 4260 7575 4295 7675
rect 4455 7575 4490 7675
rect 4510 7575 4545 7675
rect 4705 7575 4740 7675
rect 4760 7575 4795 7675
rect 4955 7575 4990 7675
rect 5010 7575 5045 7675
rect 5205 7575 5240 7675
rect 5260 7575 5295 7675
rect 5455 7575 5490 7675
rect 5510 7575 5545 7675
rect 5705 7575 5740 7675
rect 5760 7575 5795 7675
rect 5955 7575 5990 7675
rect 6010 7575 6045 7675
rect 6205 7575 6240 7675
rect 6260 7575 6295 7675
rect 6455 7575 6490 7675
rect 6510 7575 6545 7675
rect 6705 7575 6740 7675
rect 6760 7575 6795 7675
rect 6955 7575 6990 7675
rect 7010 7575 7045 7675
rect 7205 7575 7240 7675
rect 7260 7575 7295 7675
rect 7455 7575 7490 7675
rect 7510 7575 7545 7675
rect 7705 7575 7740 7675
rect 7760 7575 7795 7675
rect 7955 7575 7990 7675
rect 75 7510 175 7545
rect 325 7510 425 7545
rect 575 7510 675 7545
rect 825 7510 925 7545
rect 1075 7510 1175 7545
rect 1325 7510 1425 7545
rect 1575 7510 1675 7545
rect 1825 7510 1925 7545
rect 2075 7510 2175 7545
rect 2325 7510 2425 7545
rect 2575 7510 2675 7545
rect 2825 7510 2925 7545
rect 3075 7510 3175 7545
rect 3325 7510 3425 7545
rect 3575 7510 3675 7545
rect 3825 7510 3925 7545
rect 4075 7510 4175 7545
rect 4325 7510 4425 7545
rect 4575 7510 4675 7545
rect 4825 7510 4925 7545
rect 5075 7510 5175 7545
rect 5325 7510 5425 7545
rect 5575 7510 5675 7545
rect 5825 7510 5925 7545
rect 6075 7510 6175 7545
rect 6325 7510 6425 7545
rect 6575 7510 6675 7545
rect 6825 7510 6925 7545
rect 7075 7510 7175 7545
rect 7325 7510 7425 7545
rect 7575 7510 7675 7545
rect 7825 7510 7925 7545
rect 75 7455 175 7490
rect 325 7455 425 7490
rect 575 7455 675 7490
rect 825 7455 925 7490
rect 1075 7455 1175 7490
rect 1325 7455 1425 7490
rect 1575 7455 1675 7490
rect 1825 7455 1925 7490
rect 2075 7455 2175 7490
rect 2325 7455 2425 7490
rect 2575 7455 2675 7490
rect 2825 7455 2925 7490
rect 3075 7455 3175 7490
rect 3325 7455 3425 7490
rect 3575 7455 3675 7490
rect 3825 7455 3925 7490
rect 4075 7455 4175 7490
rect 4325 7455 4425 7490
rect 4575 7455 4675 7490
rect 4825 7455 4925 7490
rect 5075 7455 5175 7490
rect 5325 7455 5425 7490
rect 5575 7455 5675 7490
rect 5825 7455 5925 7490
rect 6075 7455 6175 7490
rect 6325 7455 6425 7490
rect 6575 7455 6675 7490
rect 6825 7455 6925 7490
rect 7075 7455 7175 7490
rect 7325 7455 7425 7490
rect 7575 7455 7675 7490
rect 7825 7455 7925 7490
rect 10 7325 45 7425
rect 205 7325 240 7425
rect 260 7325 295 7425
rect 455 7325 490 7425
rect 510 7325 545 7425
rect 705 7325 740 7425
rect 760 7325 795 7425
rect 955 7325 990 7425
rect 1010 7325 1045 7425
rect 1205 7325 1240 7425
rect 1260 7325 1295 7425
rect 1455 7325 1490 7425
rect 1510 7325 1545 7425
rect 1705 7325 1740 7425
rect 1760 7325 1795 7425
rect 1955 7325 1990 7425
rect 2010 7325 2045 7425
rect 2205 7325 2240 7425
rect 2260 7325 2295 7425
rect 2455 7325 2490 7425
rect 2510 7325 2545 7425
rect 2705 7325 2740 7425
rect 2760 7325 2795 7425
rect 2955 7325 2990 7425
rect 3010 7325 3045 7425
rect 3205 7325 3240 7425
rect 3260 7325 3295 7425
rect 3455 7325 3490 7425
rect 3510 7325 3545 7425
rect 3705 7325 3740 7425
rect 3760 7325 3795 7425
rect 3955 7325 3990 7425
rect 4010 7325 4045 7425
rect 4205 7325 4240 7425
rect 4260 7325 4295 7425
rect 4455 7325 4490 7425
rect 4510 7325 4545 7425
rect 4705 7325 4740 7425
rect 4760 7325 4795 7425
rect 4955 7325 4990 7425
rect 5010 7325 5045 7425
rect 5205 7325 5240 7425
rect 5260 7325 5295 7425
rect 5455 7325 5490 7425
rect 5510 7325 5545 7425
rect 5705 7325 5740 7425
rect 5760 7325 5795 7425
rect 5955 7325 5990 7425
rect 6010 7325 6045 7425
rect 6205 7325 6240 7425
rect 6260 7325 6295 7425
rect 6455 7325 6490 7425
rect 6510 7325 6545 7425
rect 6705 7325 6740 7425
rect 6760 7325 6795 7425
rect 6955 7325 6990 7425
rect 7010 7325 7045 7425
rect 7205 7325 7240 7425
rect 7260 7325 7295 7425
rect 7455 7325 7490 7425
rect 7510 7325 7545 7425
rect 7705 7325 7740 7425
rect 7760 7325 7795 7425
rect 7955 7325 7990 7425
rect 75 7260 175 7295
rect 325 7260 425 7295
rect 575 7260 675 7295
rect 825 7260 925 7295
rect 1075 7260 1175 7295
rect 1325 7260 1425 7295
rect 1575 7260 1675 7295
rect 1825 7260 1925 7295
rect 2075 7260 2175 7295
rect 2325 7260 2425 7295
rect 2575 7260 2675 7295
rect 2825 7260 2925 7295
rect 3075 7260 3175 7295
rect 3325 7260 3425 7295
rect 3575 7260 3675 7295
rect 3825 7260 3925 7295
rect 4075 7260 4175 7295
rect 4325 7260 4425 7295
rect 4575 7260 4675 7295
rect 4825 7260 4925 7295
rect 5075 7260 5175 7295
rect 5325 7260 5425 7295
rect 5575 7260 5675 7295
rect 5825 7260 5925 7295
rect 6075 7260 6175 7295
rect 6325 7260 6425 7295
rect 6575 7260 6675 7295
rect 6825 7260 6925 7295
rect 7075 7260 7175 7295
rect 7325 7260 7425 7295
rect 7575 7260 7675 7295
rect 7825 7260 7925 7295
rect 75 7205 175 7240
rect 325 7205 425 7240
rect 575 7205 675 7240
rect 825 7205 925 7240
rect 1075 7205 1175 7240
rect 1325 7205 1425 7240
rect 1575 7205 1675 7240
rect 1825 7205 1925 7240
rect 2075 7205 2175 7240
rect 2325 7205 2425 7240
rect 2575 7205 2675 7240
rect 2825 7205 2925 7240
rect 3075 7205 3175 7240
rect 3325 7205 3425 7240
rect 3575 7205 3675 7240
rect 3825 7205 3925 7240
rect 4075 7205 4175 7240
rect 4325 7205 4425 7240
rect 4575 7205 4675 7240
rect 4825 7205 4925 7240
rect 5075 7205 5175 7240
rect 5325 7205 5425 7240
rect 5575 7205 5675 7240
rect 5825 7205 5925 7240
rect 6075 7205 6175 7240
rect 6325 7205 6425 7240
rect 6575 7205 6675 7240
rect 6825 7205 6925 7240
rect 7075 7205 7175 7240
rect 7325 7205 7425 7240
rect 7575 7205 7675 7240
rect 7825 7205 7925 7240
rect 10 7075 45 7175
rect 205 7075 240 7175
rect 260 7075 295 7175
rect 455 7075 490 7175
rect 510 7075 545 7175
rect 705 7075 740 7175
rect 760 7075 795 7175
rect 955 7075 990 7175
rect 1010 7075 1045 7175
rect 1205 7075 1240 7175
rect 1260 7075 1295 7175
rect 1455 7075 1490 7175
rect 1510 7075 1545 7175
rect 1705 7075 1740 7175
rect 1760 7075 1795 7175
rect 1955 7075 1990 7175
rect 2010 7075 2045 7175
rect 2205 7075 2240 7175
rect 2260 7075 2295 7175
rect 2455 7075 2490 7175
rect 2510 7075 2545 7175
rect 2705 7075 2740 7175
rect 2760 7075 2795 7175
rect 2955 7075 2990 7175
rect 3010 7075 3045 7175
rect 3205 7075 3240 7175
rect 3260 7075 3295 7175
rect 3455 7075 3490 7175
rect 3510 7075 3545 7175
rect 3705 7075 3740 7175
rect 3760 7075 3795 7175
rect 3955 7075 3990 7175
rect 4010 7075 4045 7175
rect 4205 7075 4240 7175
rect 4260 7075 4295 7175
rect 4455 7075 4490 7175
rect 4510 7075 4545 7175
rect 4705 7075 4740 7175
rect 4760 7075 4795 7175
rect 4955 7075 4990 7175
rect 5010 7075 5045 7175
rect 5205 7075 5240 7175
rect 5260 7075 5295 7175
rect 5455 7075 5490 7175
rect 5510 7075 5545 7175
rect 5705 7075 5740 7175
rect 5760 7075 5795 7175
rect 5955 7075 5990 7175
rect 6010 7075 6045 7175
rect 6205 7075 6240 7175
rect 6260 7075 6295 7175
rect 6455 7075 6490 7175
rect 6510 7075 6545 7175
rect 6705 7075 6740 7175
rect 6760 7075 6795 7175
rect 6955 7075 6990 7175
rect 7010 7075 7045 7175
rect 7205 7075 7240 7175
rect 7260 7075 7295 7175
rect 7455 7075 7490 7175
rect 7510 7075 7545 7175
rect 7705 7075 7740 7175
rect 7760 7075 7795 7175
rect 7955 7075 7990 7175
rect 75 7010 175 7045
rect 325 7010 425 7045
rect 575 7010 675 7045
rect 825 7010 925 7045
rect 1075 7010 1175 7045
rect 1325 7010 1425 7045
rect 1575 7010 1675 7045
rect 1825 7010 1925 7045
rect 2075 7010 2175 7045
rect 2325 7010 2425 7045
rect 2575 7010 2675 7045
rect 2825 7010 2925 7045
rect 3075 7010 3175 7045
rect 3325 7010 3425 7045
rect 3575 7010 3675 7045
rect 3825 7010 3925 7045
rect 4075 7010 4175 7045
rect 4325 7010 4425 7045
rect 4575 7010 4675 7045
rect 4825 7010 4925 7045
rect 5075 7010 5175 7045
rect 5325 7010 5425 7045
rect 5575 7010 5675 7045
rect 5825 7010 5925 7045
rect 6075 7010 6175 7045
rect 6325 7010 6425 7045
rect 6575 7010 6675 7045
rect 6825 7010 6925 7045
rect 7075 7010 7175 7045
rect 7325 7010 7425 7045
rect 7575 7010 7675 7045
rect 7825 7010 7925 7045
rect 75 6955 175 6990
rect 325 6955 425 6990
rect 575 6955 675 6990
rect 825 6955 925 6990
rect 1075 6955 1175 6990
rect 1325 6955 1425 6990
rect 1575 6955 1675 6990
rect 1825 6955 1925 6990
rect 2075 6955 2175 6990
rect 2325 6955 2425 6990
rect 2575 6955 2675 6990
rect 2825 6955 2925 6990
rect 3075 6955 3175 6990
rect 3325 6955 3425 6990
rect 3575 6955 3675 6990
rect 3825 6955 3925 6990
rect 4075 6955 4175 6990
rect 4325 6955 4425 6990
rect 4575 6955 4675 6990
rect 4825 6955 4925 6990
rect 5075 6955 5175 6990
rect 5325 6955 5425 6990
rect 5575 6955 5675 6990
rect 5825 6955 5925 6990
rect 6075 6955 6175 6990
rect 6325 6955 6425 6990
rect 6575 6955 6675 6990
rect 6825 6955 6925 6990
rect 7075 6955 7175 6990
rect 7325 6955 7425 6990
rect 7575 6955 7675 6990
rect 7825 6955 7925 6990
rect 10 6825 45 6925
rect 205 6825 240 6925
rect 260 6825 295 6925
rect 455 6825 490 6925
rect 510 6825 545 6925
rect 705 6825 740 6925
rect 760 6825 795 6925
rect 955 6825 990 6925
rect 1010 6825 1045 6925
rect 1205 6825 1240 6925
rect 1260 6825 1295 6925
rect 1455 6825 1490 6925
rect 1510 6825 1545 6925
rect 1705 6825 1740 6925
rect 1760 6825 1795 6925
rect 1955 6825 1990 6925
rect 2010 6825 2045 6925
rect 2205 6825 2240 6925
rect 2260 6825 2295 6925
rect 2455 6825 2490 6925
rect 2510 6825 2545 6925
rect 2705 6825 2740 6925
rect 2760 6825 2795 6925
rect 2955 6825 2990 6925
rect 3010 6825 3045 6925
rect 3205 6825 3240 6925
rect 3260 6825 3295 6925
rect 3455 6825 3490 6925
rect 3510 6825 3545 6925
rect 3705 6825 3740 6925
rect 3760 6825 3795 6925
rect 3955 6825 3990 6925
rect 4010 6825 4045 6925
rect 4205 6825 4240 6925
rect 4260 6825 4295 6925
rect 4455 6825 4490 6925
rect 4510 6825 4545 6925
rect 4705 6825 4740 6925
rect 4760 6825 4795 6925
rect 4955 6825 4990 6925
rect 5010 6825 5045 6925
rect 5205 6825 5240 6925
rect 5260 6825 5295 6925
rect 5455 6825 5490 6925
rect 5510 6825 5545 6925
rect 5705 6825 5740 6925
rect 5760 6825 5795 6925
rect 5955 6825 5990 6925
rect 6010 6825 6045 6925
rect 6205 6825 6240 6925
rect 6260 6825 6295 6925
rect 6455 6825 6490 6925
rect 6510 6825 6545 6925
rect 6705 6825 6740 6925
rect 6760 6825 6795 6925
rect 6955 6825 6990 6925
rect 7010 6825 7045 6925
rect 7205 6825 7240 6925
rect 7260 6825 7295 6925
rect 7455 6825 7490 6925
rect 7510 6825 7545 6925
rect 7705 6825 7740 6925
rect 7760 6825 7795 6925
rect 7955 6825 7990 6925
rect 75 6760 175 6795
rect 325 6760 425 6795
rect 575 6760 675 6795
rect 825 6760 925 6795
rect 1075 6760 1175 6795
rect 1325 6760 1425 6795
rect 1575 6760 1675 6795
rect 1825 6760 1925 6795
rect 2075 6760 2175 6795
rect 2325 6760 2425 6795
rect 2575 6760 2675 6795
rect 2825 6760 2925 6795
rect 3075 6760 3175 6795
rect 3325 6760 3425 6795
rect 3575 6760 3675 6795
rect 3825 6760 3925 6795
rect 4075 6760 4175 6795
rect 4325 6760 4425 6795
rect 4575 6760 4675 6795
rect 4825 6760 4925 6795
rect 5075 6760 5175 6795
rect 5325 6760 5425 6795
rect 5575 6760 5675 6795
rect 5825 6760 5925 6795
rect 6075 6760 6175 6795
rect 6325 6760 6425 6795
rect 6575 6760 6675 6795
rect 6825 6760 6925 6795
rect 7075 6760 7175 6795
rect 7325 6760 7425 6795
rect 7575 6760 7675 6795
rect 7825 6760 7925 6795
rect 75 6705 175 6740
rect 325 6705 425 6740
rect 575 6705 675 6740
rect 825 6705 925 6740
rect 1075 6705 1175 6740
rect 1325 6705 1425 6740
rect 1575 6705 1675 6740
rect 1825 6705 1925 6740
rect 2075 6705 2175 6740
rect 2325 6705 2425 6740
rect 2575 6705 2675 6740
rect 2825 6705 2925 6740
rect 3075 6705 3175 6740
rect 3325 6705 3425 6740
rect 3575 6705 3675 6740
rect 3825 6705 3925 6740
rect 4075 6705 4175 6740
rect 4325 6705 4425 6740
rect 4575 6705 4675 6740
rect 4825 6705 4925 6740
rect 5075 6705 5175 6740
rect 5325 6705 5425 6740
rect 5575 6705 5675 6740
rect 5825 6705 5925 6740
rect 6075 6705 6175 6740
rect 6325 6705 6425 6740
rect 6575 6705 6675 6740
rect 6825 6705 6925 6740
rect 7075 6705 7175 6740
rect 7325 6705 7425 6740
rect 7575 6705 7675 6740
rect 7825 6705 7925 6740
rect 10 6575 45 6675
rect 205 6575 240 6675
rect 260 6575 295 6675
rect 455 6575 490 6675
rect 510 6575 545 6675
rect 705 6575 740 6675
rect 760 6575 795 6675
rect 955 6575 990 6675
rect 1010 6575 1045 6675
rect 1205 6575 1240 6675
rect 1260 6575 1295 6675
rect 1455 6575 1490 6675
rect 1510 6575 1545 6675
rect 1705 6575 1740 6675
rect 1760 6575 1795 6675
rect 1955 6575 1990 6675
rect 2010 6575 2045 6675
rect 2205 6575 2240 6675
rect 2260 6575 2295 6675
rect 2455 6575 2490 6675
rect 2510 6575 2545 6675
rect 2705 6575 2740 6675
rect 2760 6575 2795 6675
rect 2955 6575 2990 6675
rect 3010 6575 3045 6675
rect 3205 6575 3240 6675
rect 3260 6575 3295 6675
rect 3455 6575 3490 6675
rect 3510 6575 3545 6675
rect 3705 6575 3740 6675
rect 3760 6575 3795 6675
rect 3955 6575 3990 6675
rect 4010 6575 4045 6675
rect 4205 6575 4240 6675
rect 4260 6575 4295 6675
rect 4455 6575 4490 6675
rect 4510 6575 4545 6675
rect 4705 6575 4740 6675
rect 4760 6575 4795 6675
rect 4955 6575 4990 6675
rect 5010 6575 5045 6675
rect 5205 6575 5240 6675
rect 5260 6575 5295 6675
rect 5455 6575 5490 6675
rect 5510 6575 5545 6675
rect 5705 6575 5740 6675
rect 5760 6575 5795 6675
rect 5955 6575 5990 6675
rect 6010 6575 6045 6675
rect 6205 6575 6240 6675
rect 6260 6575 6295 6675
rect 6455 6575 6490 6675
rect 6510 6575 6545 6675
rect 6705 6575 6740 6675
rect 6760 6575 6795 6675
rect 6955 6575 6990 6675
rect 7010 6575 7045 6675
rect 7205 6575 7240 6675
rect 7260 6575 7295 6675
rect 7455 6575 7490 6675
rect 7510 6575 7545 6675
rect 7705 6575 7740 6675
rect 7760 6575 7795 6675
rect 7955 6575 7990 6675
rect 75 6510 175 6545
rect 325 6510 425 6545
rect 575 6510 675 6545
rect 825 6510 925 6545
rect 1075 6510 1175 6545
rect 1325 6510 1425 6545
rect 1575 6510 1675 6545
rect 1825 6510 1925 6545
rect 2075 6510 2175 6545
rect 2325 6510 2425 6545
rect 2575 6510 2675 6545
rect 2825 6510 2925 6545
rect 3075 6510 3175 6545
rect 3325 6510 3425 6545
rect 3575 6510 3675 6545
rect 3825 6510 3925 6545
rect 4075 6510 4175 6545
rect 4325 6510 4425 6545
rect 4575 6510 4675 6545
rect 4825 6510 4925 6545
rect 5075 6510 5175 6545
rect 5325 6510 5425 6545
rect 5575 6510 5675 6545
rect 5825 6510 5925 6545
rect 6075 6510 6175 6545
rect 6325 6510 6425 6545
rect 6575 6510 6675 6545
rect 6825 6510 6925 6545
rect 7075 6510 7175 6545
rect 7325 6510 7425 6545
rect 7575 6510 7675 6545
rect 7825 6510 7925 6545
rect 75 6455 175 6490
rect 325 6455 425 6490
rect 575 6455 675 6490
rect 825 6455 925 6490
rect 1075 6455 1175 6490
rect 1325 6455 1425 6490
rect 1575 6455 1675 6490
rect 1825 6455 1925 6490
rect 2075 6455 2175 6490
rect 2325 6455 2425 6490
rect 2575 6455 2675 6490
rect 2825 6455 2925 6490
rect 3075 6455 3175 6490
rect 3325 6455 3425 6490
rect 3575 6455 3675 6490
rect 3825 6455 3925 6490
rect 4075 6455 4175 6490
rect 4325 6455 4425 6490
rect 4575 6455 4675 6490
rect 4825 6455 4925 6490
rect 5075 6455 5175 6490
rect 5325 6455 5425 6490
rect 5575 6455 5675 6490
rect 5825 6455 5925 6490
rect 6075 6455 6175 6490
rect 6325 6455 6425 6490
rect 6575 6455 6675 6490
rect 6825 6455 6925 6490
rect 7075 6455 7175 6490
rect 7325 6455 7425 6490
rect 7575 6455 7675 6490
rect 7825 6455 7925 6490
rect 10 6325 45 6425
rect 205 6325 240 6425
rect 260 6325 295 6425
rect 455 6325 490 6425
rect 510 6325 545 6425
rect 705 6325 740 6425
rect 760 6325 795 6425
rect 955 6325 990 6425
rect 1010 6325 1045 6425
rect 1205 6325 1240 6425
rect 1260 6325 1295 6425
rect 1455 6325 1490 6425
rect 1510 6325 1545 6425
rect 1705 6325 1740 6425
rect 1760 6325 1795 6425
rect 1955 6325 1990 6425
rect 2010 6325 2045 6425
rect 2205 6325 2240 6425
rect 2260 6325 2295 6425
rect 2455 6325 2490 6425
rect 2510 6325 2545 6425
rect 2705 6325 2740 6425
rect 2760 6325 2795 6425
rect 2955 6325 2990 6425
rect 3010 6325 3045 6425
rect 3205 6325 3240 6425
rect 3260 6325 3295 6425
rect 3455 6325 3490 6425
rect 3510 6325 3545 6425
rect 3705 6325 3740 6425
rect 3760 6325 3795 6425
rect 3955 6325 3990 6425
rect 4010 6325 4045 6425
rect 4205 6325 4240 6425
rect 4260 6325 4295 6425
rect 4455 6325 4490 6425
rect 4510 6325 4545 6425
rect 4705 6325 4740 6425
rect 4760 6325 4795 6425
rect 4955 6325 4990 6425
rect 5010 6325 5045 6425
rect 5205 6325 5240 6425
rect 5260 6325 5295 6425
rect 5455 6325 5490 6425
rect 5510 6325 5545 6425
rect 5705 6325 5740 6425
rect 5760 6325 5795 6425
rect 5955 6325 5990 6425
rect 6010 6325 6045 6425
rect 6205 6325 6240 6425
rect 6260 6325 6295 6425
rect 6455 6325 6490 6425
rect 6510 6325 6545 6425
rect 6705 6325 6740 6425
rect 6760 6325 6795 6425
rect 6955 6325 6990 6425
rect 7010 6325 7045 6425
rect 7205 6325 7240 6425
rect 7260 6325 7295 6425
rect 7455 6325 7490 6425
rect 7510 6325 7545 6425
rect 7705 6325 7740 6425
rect 7760 6325 7795 6425
rect 7955 6325 7990 6425
rect 75 6260 175 6295
rect 325 6260 425 6295
rect 575 6260 675 6295
rect 825 6260 925 6295
rect 1075 6260 1175 6295
rect 1325 6260 1425 6295
rect 1575 6260 1675 6295
rect 1825 6260 1925 6295
rect 2075 6260 2175 6295
rect 2325 6260 2425 6295
rect 2575 6260 2675 6295
rect 2825 6260 2925 6295
rect 3075 6260 3175 6295
rect 3325 6260 3425 6295
rect 3575 6260 3675 6295
rect 3825 6260 3925 6295
rect 4075 6260 4175 6295
rect 4325 6260 4425 6295
rect 4575 6260 4675 6295
rect 4825 6260 4925 6295
rect 5075 6260 5175 6295
rect 5325 6260 5425 6295
rect 5575 6260 5675 6295
rect 5825 6260 5925 6295
rect 6075 6260 6175 6295
rect 6325 6260 6425 6295
rect 6575 6260 6675 6295
rect 6825 6260 6925 6295
rect 7075 6260 7175 6295
rect 7325 6260 7425 6295
rect 7575 6260 7675 6295
rect 7825 6260 7925 6295
rect 75 6205 175 6240
rect 325 6205 425 6240
rect 575 6205 675 6240
rect 825 6205 925 6240
rect 1075 6205 1175 6240
rect 1325 6205 1425 6240
rect 1575 6205 1675 6240
rect 1825 6205 1925 6240
rect 2075 6205 2175 6240
rect 2325 6205 2425 6240
rect 2575 6205 2675 6240
rect 2825 6205 2925 6240
rect 3075 6205 3175 6240
rect 3325 6205 3425 6240
rect 3575 6205 3675 6240
rect 3825 6205 3925 6240
rect 4075 6205 4175 6240
rect 4325 6205 4425 6240
rect 4575 6205 4675 6240
rect 4825 6205 4925 6240
rect 5075 6205 5175 6240
rect 5325 6205 5425 6240
rect 5575 6205 5675 6240
rect 5825 6205 5925 6240
rect 6075 6205 6175 6240
rect 6325 6205 6425 6240
rect 6575 6205 6675 6240
rect 6825 6205 6925 6240
rect 7075 6205 7175 6240
rect 7325 6205 7425 6240
rect 7575 6205 7675 6240
rect 7825 6205 7925 6240
rect 10 6075 45 6175
rect 205 6075 240 6175
rect 260 6075 295 6175
rect 455 6075 490 6175
rect 510 6075 545 6175
rect 705 6075 740 6175
rect 760 6075 795 6175
rect 955 6075 990 6175
rect 1010 6075 1045 6175
rect 1205 6075 1240 6175
rect 1260 6075 1295 6175
rect 1455 6075 1490 6175
rect 1510 6075 1545 6175
rect 1705 6075 1740 6175
rect 1760 6075 1795 6175
rect 1955 6075 1990 6175
rect 2010 6075 2045 6175
rect 2205 6075 2240 6175
rect 2260 6075 2295 6175
rect 2455 6075 2490 6175
rect 2510 6075 2545 6175
rect 2705 6075 2740 6175
rect 2760 6075 2795 6175
rect 2955 6075 2990 6175
rect 3010 6075 3045 6175
rect 3205 6075 3240 6175
rect 3260 6075 3295 6175
rect 3455 6075 3490 6175
rect 3510 6075 3545 6175
rect 3705 6075 3740 6175
rect 3760 6075 3795 6175
rect 3955 6075 3990 6175
rect 4010 6075 4045 6175
rect 4205 6075 4240 6175
rect 4260 6075 4295 6175
rect 4455 6075 4490 6175
rect 4510 6075 4545 6175
rect 4705 6075 4740 6175
rect 4760 6075 4795 6175
rect 4955 6075 4990 6175
rect 5010 6075 5045 6175
rect 5205 6075 5240 6175
rect 5260 6075 5295 6175
rect 5455 6075 5490 6175
rect 5510 6075 5545 6175
rect 5705 6075 5740 6175
rect 5760 6075 5795 6175
rect 5955 6075 5990 6175
rect 6010 6075 6045 6175
rect 6205 6075 6240 6175
rect 6260 6075 6295 6175
rect 6455 6075 6490 6175
rect 6510 6075 6545 6175
rect 6705 6075 6740 6175
rect 6760 6075 6795 6175
rect 6955 6075 6990 6175
rect 7010 6075 7045 6175
rect 7205 6075 7240 6175
rect 7260 6075 7295 6175
rect 7455 6075 7490 6175
rect 7510 6075 7545 6175
rect 7705 6075 7740 6175
rect 7760 6075 7795 6175
rect 7955 6075 7990 6175
rect 75 6010 175 6045
rect 325 6010 425 6045
rect 575 6010 675 6045
rect 825 6010 925 6045
rect 1075 6010 1175 6045
rect 1325 6010 1425 6045
rect 1575 6010 1675 6045
rect 1825 6010 1925 6045
rect 2075 6010 2175 6045
rect 2325 6010 2425 6045
rect 2575 6010 2675 6045
rect 2825 6010 2925 6045
rect 3075 6010 3175 6045
rect 3325 6010 3425 6045
rect 3575 6010 3675 6045
rect 3825 6010 3925 6045
rect 4075 6010 4175 6045
rect 4325 6010 4425 6045
rect 4575 6010 4675 6045
rect 4825 6010 4925 6045
rect 5075 6010 5175 6045
rect 5325 6010 5425 6045
rect 5575 6010 5675 6045
rect 5825 6010 5925 6045
rect 6075 6010 6175 6045
rect 6325 6010 6425 6045
rect 6575 6010 6675 6045
rect 6825 6010 6925 6045
rect 7075 6010 7175 6045
rect 7325 6010 7425 6045
rect 7575 6010 7675 6045
rect 7825 6010 7925 6045
rect 75 5955 175 5990
rect 325 5955 425 5990
rect 575 5955 675 5990
rect 825 5955 925 5990
rect 1075 5955 1175 5990
rect 1325 5955 1425 5990
rect 1575 5955 1675 5990
rect 1825 5955 1925 5990
rect 2075 5955 2175 5990
rect 2325 5955 2425 5990
rect 2575 5955 2675 5990
rect 2825 5955 2925 5990
rect 3075 5955 3175 5990
rect 3325 5955 3425 5990
rect 3575 5955 3675 5990
rect 3825 5955 3925 5990
rect 4075 5955 4175 5990
rect 4325 5955 4425 5990
rect 4575 5955 4675 5990
rect 4825 5955 4925 5990
rect 5075 5955 5175 5990
rect 5325 5955 5425 5990
rect 5575 5955 5675 5990
rect 5825 5955 5925 5990
rect 6075 5955 6175 5990
rect 6325 5955 6425 5990
rect 6575 5955 6675 5990
rect 6825 5955 6925 5990
rect 7075 5955 7175 5990
rect 7325 5955 7425 5990
rect 7575 5955 7675 5990
rect 7825 5955 7925 5990
rect 10 5825 45 5925
rect 205 5825 240 5925
rect 260 5825 295 5925
rect 455 5825 490 5925
rect 510 5825 545 5925
rect 705 5825 740 5925
rect 760 5825 795 5925
rect 955 5825 990 5925
rect 1010 5825 1045 5925
rect 1205 5825 1240 5925
rect 1260 5825 1295 5925
rect 1455 5825 1490 5925
rect 1510 5825 1545 5925
rect 1705 5825 1740 5925
rect 1760 5825 1795 5925
rect 1955 5825 1990 5925
rect 2010 5825 2045 5925
rect 2205 5825 2240 5925
rect 2260 5825 2295 5925
rect 2455 5825 2490 5925
rect 2510 5825 2545 5925
rect 2705 5825 2740 5925
rect 2760 5825 2795 5925
rect 2955 5825 2990 5925
rect 3010 5825 3045 5925
rect 3205 5825 3240 5925
rect 3260 5825 3295 5925
rect 3455 5825 3490 5925
rect 3510 5825 3545 5925
rect 3705 5825 3740 5925
rect 3760 5825 3795 5925
rect 3955 5825 3990 5925
rect 4010 5825 4045 5925
rect 4205 5825 4240 5925
rect 4260 5825 4295 5925
rect 4455 5825 4490 5925
rect 4510 5825 4545 5925
rect 4705 5825 4740 5925
rect 4760 5825 4795 5925
rect 4955 5825 4990 5925
rect 5010 5825 5045 5925
rect 5205 5825 5240 5925
rect 5260 5825 5295 5925
rect 5455 5825 5490 5925
rect 5510 5825 5545 5925
rect 5705 5825 5740 5925
rect 5760 5825 5795 5925
rect 5955 5825 5990 5925
rect 6010 5825 6045 5925
rect 6205 5825 6240 5925
rect 6260 5825 6295 5925
rect 6455 5825 6490 5925
rect 6510 5825 6545 5925
rect 6705 5825 6740 5925
rect 6760 5825 6795 5925
rect 6955 5825 6990 5925
rect 7010 5825 7045 5925
rect 7205 5825 7240 5925
rect 7260 5825 7295 5925
rect 7455 5825 7490 5925
rect 7510 5825 7545 5925
rect 7705 5825 7740 5925
rect 7760 5825 7795 5925
rect 7955 5825 7990 5925
rect 75 5760 175 5795
rect 325 5760 425 5795
rect 575 5760 675 5795
rect 825 5760 925 5795
rect 1075 5760 1175 5795
rect 1325 5760 1425 5795
rect 1575 5760 1675 5795
rect 1825 5760 1925 5795
rect 2075 5760 2175 5795
rect 2325 5760 2425 5795
rect 2575 5760 2675 5795
rect 2825 5760 2925 5795
rect 3075 5760 3175 5795
rect 3325 5760 3425 5795
rect 3575 5760 3675 5795
rect 3825 5760 3925 5795
rect 4075 5760 4175 5795
rect 4325 5760 4425 5795
rect 4575 5760 4675 5795
rect 4825 5760 4925 5795
rect 5075 5760 5175 5795
rect 5325 5760 5425 5795
rect 5575 5760 5675 5795
rect 5825 5760 5925 5795
rect 6075 5760 6175 5795
rect 6325 5760 6425 5795
rect 6575 5760 6675 5795
rect 6825 5760 6925 5795
rect 7075 5760 7175 5795
rect 7325 5760 7425 5795
rect 7575 5760 7675 5795
rect 7825 5760 7925 5795
rect 75 5705 175 5740
rect 325 5705 425 5740
rect 575 5705 675 5740
rect 825 5705 925 5740
rect 1075 5705 1175 5740
rect 1325 5705 1425 5740
rect 1575 5705 1675 5740
rect 1825 5705 1925 5740
rect 2075 5705 2175 5740
rect 2325 5705 2425 5740
rect 2575 5705 2675 5740
rect 2825 5705 2925 5740
rect 3075 5705 3175 5740
rect 3325 5705 3425 5740
rect 3575 5705 3675 5740
rect 3825 5705 3925 5740
rect 4075 5705 4175 5740
rect 4325 5705 4425 5740
rect 4575 5705 4675 5740
rect 4825 5705 4925 5740
rect 5075 5705 5175 5740
rect 5325 5705 5425 5740
rect 5575 5705 5675 5740
rect 5825 5705 5925 5740
rect 6075 5705 6175 5740
rect 6325 5705 6425 5740
rect 6575 5705 6675 5740
rect 6825 5705 6925 5740
rect 7075 5705 7175 5740
rect 7325 5705 7425 5740
rect 7575 5705 7675 5740
rect 7825 5705 7925 5740
rect 10 5575 45 5675
rect 205 5575 240 5675
rect 260 5575 295 5675
rect 455 5575 490 5675
rect 510 5575 545 5675
rect 705 5575 740 5675
rect 760 5575 795 5675
rect 955 5575 990 5675
rect 1010 5575 1045 5675
rect 1205 5575 1240 5675
rect 1260 5575 1295 5675
rect 1455 5575 1490 5675
rect 1510 5575 1545 5675
rect 1705 5575 1740 5675
rect 1760 5575 1795 5675
rect 1955 5575 1990 5675
rect 2010 5575 2045 5675
rect 2205 5575 2240 5675
rect 2260 5575 2295 5675
rect 2455 5575 2490 5675
rect 2510 5575 2545 5675
rect 2705 5575 2740 5675
rect 2760 5575 2795 5675
rect 2955 5575 2990 5675
rect 3010 5575 3045 5675
rect 3205 5575 3240 5675
rect 3260 5575 3295 5675
rect 3455 5575 3490 5675
rect 3510 5575 3545 5675
rect 3705 5575 3740 5675
rect 3760 5575 3795 5675
rect 3955 5575 3990 5675
rect 4010 5575 4045 5675
rect 4205 5575 4240 5675
rect 4260 5575 4295 5675
rect 4455 5575 4490 5675
rect 4510 5575 4545 5675
rect 4705 5575 4740 5675
rect 4760 5575 4795 5675
rect 4955 5575 4990 5675
rect 5010 5575 5045 5675
rect 5205 5575 5240 5675
rect 5260 5575 5295 5675
rect 5455 5575 5490 5675
rect 5510 5575 5545 5675
rect 5705 5575 5740 5675
rect 5760 5575 5795 5675
rect 5955 5575 5990 5675
rect 6010 5575 6045 5675
rect 6205 5575 6240 5675
rect 6260 5575 6295 5675
rect 6455 5575 6490 5675
rect 6510 5575 6545 5675
rect 6705 5575 6740 5675
rect 6760 5575 6795 5675
rect 6955 5575 6990 5675
rect 7010 5575 7045 5675
rect 7205 5575 7240 5675
rect 7260 5575 7295 5675
rect 7455 5575 7490 5675
rect 7510 5575 7545 5675
rect 7705 5575 7740 5675
rect 7760 5575 7795 5675
rect 7955 5575 7990 5675
rect 75 5510 175 5545
rect 325 5510 425 5545
rect 575 5510 675 5545
rect 825 5510 925 5545
rect 1075 5510 1175 5545
rect 1325 5510 1425 5545
rect 1575 5510 1675 5545
rect 1825 5510 1925 5545
rect 2075 5510 2175 5545
rect 2325 5510 2425 5545
rect 2575 5510 2675 5545
rect 2825 5510 2925 5545
rect 3075 5510 3175 5545
rect 3325 5510 3425 5545
rect 3575 5510 3675 5545
rect 3825 5510 3925 5545
rect 4075 5510 4175 5545
rect 4325 5510 4425 5545
rect 4575 5510 4675 5545
rect 4825 5510 4925 5545
rect 5075 5510 5175 5545
rect 5325 5510 5425 5545
rect 5575 5510 5675 5545
rect 5825 5510 5925 5545
rect 6075 5510 6175 5545
rect 6325 5510 6425 5545
rect 6575 5510 6675 5545
rect 6825 5510 6925 5545
rect 7075 5510 7175 5545
rect 7325 5510 7425 5545
rect 7575 5510 7675 5545
rect 7825 5510 7925 5545
rect 75 5455 175 5490
rect 325 5455 425 5490
rect 575 5455 675 5490
rect 825 5455 925 5490
rect 1075 5455 1175 5490
rect 1325 5455 1425 5490
rect 1575 5455 1675 5490
rect 1825 5455 1925 5490
rect 2075 5455 2175 5490
rect 2325 5455 2425 5490
rect 2575 5455 2675 5490
rect 2825 5455 2925 5490
rect 3075 5455 3175 5490
rect 3325 5455 3425 5490
rect 3575 5455 3675 5490
rect 3825 5455 3925 5490
rect 4075 5455 4175 5490
rect 4325 5455 4425 5490
rect 4575 5455 4675 5490
rect 4825 5455 4925 5490
rect 5075 5455 5175 5490
rect 5325 5455 5425 5490
rect 5575 5455 5675 5490
rect 5825 5455 5925 5490
rect 6075 5455 6175 5490
rect 6325 5455 6425 5490
rect 6575 5455 6675 5490
rect 6825 5455 6925 5490
rect 7075 5455 7175 5490
rect 7325 5455 7425 5490
rect 7575 5455 7675 5490
rect 7825 5455 7925 5490
rect 10 5325 45 5425
rect 205 5325 240 5425
rect 260 5325 295 5425
rect 455 5325 490 5425
rect 510 5325 545 5425
rect 705 5325 740 5425
rect 760 5325 795 5425
rect 955 5325 990 5425
rect 1010 5325 1045 5425
rect 1205 5325 1240 5425
rect 1260 5325 1295 5425
rect 1455 5325 1490 5425
rect 1510 5325 1545 5425
rect 1705 5325 1740 5425
rect 1760 5325 1795 5425
rect 1955 5325 1990 5425
rect 2010 5325 2045 5425
rect 2205 5325 2240 5425
rect 2260 5325 2295 5425
rect 2455 5325 2490 5425
rect 2510 5325 2545 5425
rect 2705 5325 2740 5425
rect 2760 5325 2795 5425
rect 2955 5325 2990 5425
rect 3010 5325 3045 5425
rect 3205 5325 3240 5425
rect 3260 5325 3295 5425
rect 3455 5325 3490 5425
rect 3510 5325 3545 5425
rect 3705 5325 3740 5425
rect 3760 5325 3795 5425
rect 3955 5325 3990 5425
rect 4010 5325 4045 5425
rect 4205 5325 4240 5425
rect 4260 5325 4295 5425
rect 4455 5325 4490 5425
rect 4510 5325 4545 5425
rect 4705 5325 4740 5425
rect 4760 5325 4795 5425
rect 4955 5325 4990 5425
rect 5010 5325 5045 5425
rect 5205 5325 5240 5425
rect 5260 5325 5295 5425
rect 5455 5325 5490 5425
rect 5510 5325 5545 5425
rect 5705 5325 5740 5425
rect 5760 5325 5795 5425
rect 5955 5325 5990 5425
rect 6010 5325 6045 5425
rect 6205 5325 6240 5425
rect 6260 5325 6295 5425
rect 6455 5325 6490 5425
rect 6510 5325 6545 5425
rect 6705 5325 6740 5425
rect 6760 5325 6795 5425
rect 6955 5325 6990 5425
rect 7010 5325 7045 5425
rect 7205 5325 7240 5425
rect 7260 5325 7295 5425
rect 7455 5325 7490 5425
rect 7510 5325 7545 5425
rect 7705 5325 7740 5425
rect 7760 5325 7795 5425
rect 7955 5325 7990 5425
rect 75 5260 175 5295
rect 325 5260 425 5295
rect 575 5260 675 5295
rect 825 5260 925 5295
rect 1075 5260 1175 5295
rect 1325 5260 1425 5295
rect 1575 5260 1675 5295
rect 1825 5260 1925 5295
rect 2075 5260 2175 5295
rect 2325 5260 2425 5295
rect 2575 5260 2675 5295
rect 2825 5260 2925 5295
rect 3075 5260 3175 5295
rect 3325 5260 3425 5295
rect 3575 5260 3675 5295
rect 3825 5260 3925 5295
rect 4075 5260 4175 5295
rect 4325 5260 4425 5295
rect 4575 5260 4675 5295
rect 4825 5260 4925 5295
rect 5075 5260 5175 5295
rect 5325 5260 5425 5295
rect 5575 5260 5675 5295
rect 5825 5260 5925 5295
rect 6075 5260 6175 5295
rect 6325 5260 6425 5295
rect 6575 5260 6675 5295
rect 6825 5260 6925 5295
rect 7075 5260 7175 5295
rect 7325 5260 7425 5295
rect 7575 5260 7675 5295
rect 7825 5260 7925 5295
rect 75 5205 175 5240
rect 325 5205 425 5240
rect 575 5205 675 5240
rect 825 5205 925 5240
rect 1075 5205 1175 5240
rect 1325 5205 1425 5240
rect 1575 5205 1675 5240
rect 1825 5205 1925 5240
rect 2075 5205 2175 5240
rect 2325 5205 2425 5240
rect 2575 5205 2675 5240
rect 2825 5205 2925 5240
rect 3075 5205 3175 5240
rect 3325 5205 3425 5240
rect 3575 5205 3675 5240
rect 3825 5205 3925 5240
rect 4075 5205 4175 5240
rect 4325 5205 4425 5240
rect 4575 5205 4675 5240
rect 4825 5205 4925 5240
rect 5075 5205 5175 5240
rect 5325 5205 5425 5240
rect 5575 5205 5675 5240
rect 5825 5205 5925 5240
rect 6075 5205 6175 5240
rect 6325 5205 6425 5240
rect 6575 5205 6675 5240
rect 6825 5205 6925 5240
rect 7075 5205 7175 5240
rect 7325 5205 7425 5240
rect 7575 5205 7675 5240
rect 7825 5205 7925 5240
rect 10 5075 45 5175
rect 205 5075 240 5175
rect 260 5075 295 5175
rect 455 5075 490 5175
rect 510 5075 545 5175
rect 705 5075 740 5175
rect 760 5075 795 5175
rect 955 5075 990 5175
rect 1010 5075 1045 5175
rect 1205 5075 1240 5175
rect 1260 5075 1295 5175
rect 1455 5075 1490 5175
rect 1510 5075 1545 5175
rect 1705 5075 1740 5175
rect 1760 5075 1795 5175
rect 1955 5075 1990 5175
rect 2010 5075 2045 5175
rect 2205 5075 2240 5175
rect 2260 5075 2295 5175
rect 2455 5075 2490 5175
rect 2510 5075 2545 5175
rect 2705 5075 2740 5175
rect 2760 5075 2795 5175
rect 2955 5075 2990 5175
rect 3010 5075 3045 5175
rect 3205 5075 3240 5175
rect 3260 5075 3295 5175
rect 3455 5075 3490 5175
rect 3510 5075 3545 5175
rect 3705 5075 3740 5175
rect 3760 5075 3795 5175
rect 3955 5075 3990 5175
rect 4010 5075 4045 5175
rect 4205 5075 4240 5175
rect 4260 5075 4295 5175
rect 4455 5075 4490 5175
rect 4510 5075 4545 5175
rect 4705 5075 4740 5175
rect 4760 5075 4795 5175
rect 4955 5075 4990 5175
rect 5010 5075 5045 5175
rect 5205 5075 5240 5175
rect 5260 5075 5295 5175
rect 5455 5075 5490 5175
rect 5510 5075 5545 5175
rect 5705 5075 5740 5175
rect 5760 5075 5795 5175
rect 5955 5075 5990 5175
rect 6010 5075 6045 5175
rect 6205 5075 6240 5175
rect 6260 5075 6295 5175
rect 6455 5075 6490 5175
rect 6510 5075 6545 5175
rect 6705 5075 6740 5175
rect 6760 5075 6795 5175
rect 6955 5075 6990 5175
rect 7010 5075 7045 5175
rect 7205 5075 7240 5175
rect 7260 5075 7295 5175
rect 7455 5075 7490 5175
rect 7510 5075 7545 5175
rect 7705 5075 7740 5175
rect 7760 5075 7795 5175
rect 7955 5075 7990 5175
rect 75 5010 175 5045
rect 325 5010 425 5045
rect 575 5010 675 5045
rect 825 5010 925 5045
rect 1075 5010 1175 5045
rect 1325 5010 1425 5045
rect 1575 5010 1675 5045
rect 1825 5010 1925 5045
rect 2075 5010 2175 5045
rect 2325 5010 2425 5045
rect 2575 5010 2675 5045
rect 2825 5010 2925 5045
rect 3075 5010 3175 5045
rect 3325 5010 3425 5045
rect 3575 5010 3675 5045
rect 3825 5010 3925 5045
rect 4075 5010 4175 5045
rect 4325 5010 4425 5045
rect 4575 5010 4675 5045
rect 4825 5010 4925 5045
rect 5075 5010 5175 5045
rect 5325 5010 5425 5045
rect 5575 5010 5675 5045
rect 5825 5010 5925 5045
rect 6075 5010 6175 5045
rect 6325 5010 6425 5045
rect 6575 5010 6675 5045
rect 6825 5010 6925 5045
rect 7075 5010 7175 5045
rect 7325 5010 7425 5045
rect 7575 5010 7675 5045
rect 7825 5010 7925 5045
rect 75 4955 175 4990
rect 325 4955 425 4990
rect 575 4955 675 4990
rect 825 4955 925 4990
rect 1075 4955 1175 4990
rect 1325 4955 1425 4990
rect 1575 4955 1675 4990
rect 1825 4955 1925 4990
rect 2075 4955 2175 4990
rect 2325 4955 2425 4990
rect 2575 4955 2675 4990
rect 2825 4955 2925 4990
rect 3075 4955 3175 4990
rect 3325 4955 3425 4990
rect 3575 4955 3675 4990
rect 3825 4955 3925 4990
rect 4075 4955 4175 4990
rect 4325 4955 4425 4990
rect 4575 4955 4675 4990
rect 4825 4955 4925 4990
rect 5075 4955 5175 4990
rect 5325 4955 5425 4990
rect 5575 4955 5675 4990
rect 5825 4955 5925 4990
rect 6075 4955 6175 4990
rect 6325 4955 6425 4990
rect 6575 4955 6675 4990
rect 6825 4955 6925 4990
rect 7075 4955 7175 4990
rect 7325 4955 7425 4990
rect 7575 4955 7675 4990
rect 7825 4955 7925 4990
rect 10 4825 45 4925
rect 205 4825 240 4925
rect 260 4825 295 4925
rect 455 4825 490 4925
rect 510 4825 545 4925
rect 705 4825 740 4925
rect 760 4825 795 4925
rect 955 4825 990 4925
rect 1010 4825 1045 4925
rect 1205 4825 1240 4925
rect 1260 4825 1295 4925
rect 1455 4825 1490 4925
rect 1510 4825 1545 4925
rect 1705 4825 1740 4925
rect 1760 4825 1795 4925
rect 1955 4825 1990 4925
rect 2010 4825 2045 4925
rect 2205 4825 2240 4925
rect 2260 4825 2295 4925
rect 2455 4825 2490 4925
rect 2510 4825 2545 4925
rect 2705 4825 2740 4925
rect 2760 4825 2795 4925
rect 2955 4825 2990 4925
rect 3010 4825 3045 4925
rect 3205 4825 3240 4925
rect 3260 4825 3295 4925
rect 3455 4825 3490 4925
rect 3510 4825 3545 4925
rect 3705 4825 3740 4925
rect 3760 4825 3795 4925
rect 3955 4825 3990 4925
rect 4010 4825 4045 4925
rect 4205 4825 4240 4925
rect 4260 4825 4295 4925
rect 4455 4825 4490 4925
rect 4510 4825 4545 4925
rect 4705 4825 4740 4925
rect 4760 4825 4795 4925
rect 4955 4825 4990 4925
rect 5010 4825 5045 4925
rect 5205 4825 5240 4925
rect 5260 4825 5295 4925
rect 5455 4825 5490 4925
rect 5510 4825 5545 4925
rect 5705 4825 5740 4925
rect 5760 4825 5795 4925
rect 5955 4825 5990 4925
rect 6010 4825 6045 4925
rect 6205 4825 6240 4925
rect 6260 4825 6295 4925
rect 6455 4825 6490 4925
rect 6510 4825 6545 4925
rect 6705 4825 6740 4925
rect 6760 4825 6795 4925
rect 6955 4825 6990 4925
rect 7010 4825 7045 4925
rect 7205 4825 7240 4925
rect 7260 4825 7295 4925
rect 7455 4825 7490 4925
rect 7510 4825 7545 4925
rect 7705 4825 7740 4925
rect 7760 4825 7795 4925
rect 7955 4825 7990 4925
rect 75 4760 175 4795
rect 325 4760 425 4795
rect 575 4760 675 4795
rect 825 4760 925 4795
rect 1075 4760 1175 4795
rect 1325 4760 1425 4795
rect 1575 4760 1675 4795
rect 1825 4760 1925 4795
rect 2075 4760 2175 4795
rect 2325 4760 2425 4795
rect 2575 4760 2675 4795
rect 2825 4760 2925 4795
rect 3075 4760 3175 4795
rect 3325 4760 3425 4795
rect 3575 4760 3675 4795
rect 3825 4760 3925 4795
rect 4075 4760 4175 4795
rect 4325 4760 4425 4795
rect 4575 4760 4675 4795
rect 4825 4760 4925 4795
rect 5075 4760 5175 4795
rect 5325 4760 5425 4795
rect 5575 4760 5675 4795
rect 5825 4760 5925 4795
rect 6075 4760 6175 4795
rect 6325 4760 6425 4795
rect 6575 4760 6675 4795
rect 6825 4760 6925 4795
rect 7075 4760 7175 4795
rect 7325 4760 7425 4795
rect 7575 4760 7675 4795
rect 7825 4760 7925 4795
rect 75 4705 175 4740
rect 325 4705 425 4740
rect 575 4705 675 4740
rect 825 4705 925 4740
rect 1075 4705 1175 4740
rect 1325 4705 1425 4740
rect 1575 4705 1675 4740
rect 1825 4705 1925 4740
rect 2075 4705 2175 4740
rect 2325 4705 2425 4740
rect 2575 4705 2675 4740
rect 2825 4705 2925 4740
rect 3075 4705 3175 4740
rect 3325 4705 3425 4740
rect 3575 4705 3675 4740
rect 3825 4705 3925 4740
rect 4075 4705 4175 4740
rect 4325 4705 4425 4740
rect 4575 4705 4675 4740
rect 4825 4705 4925 4740
rect 5075 4705 5175 4740
rect 5325 4705 5425 4740
rect 5575 4705 5675 4740
rect 5825 4705 5925 4740
rect 6075 4705 6175 4740
rect 6325 4705 6425 4740
rect 6575 4705 6675 4740
rect 6825 4705 6925 4740
rect 7075 4705 7175 4740
rect 7325 4705 7425 4740
rect 7575 4705 7675 4740
rect 7825 4705 7925 4740
rect 10 4575 45 4675
rect 205 4575 240 4675
rect 260 4575 295 4675
rect 455 4575 490 4675
rect 510 4575 545 4675
rect 705 4575 740 4675
rect 760 4575 795 4675
rect 955 4575 990 4675
rect 1010 4575 1045 4675
rect 1205 4575 1240 4675
rect 1260 4575 1295 4675
rect 1455 4575 1490 4675
rect 1510 4575 1545 4675
rect 1705 4575 1740 4675
rect 1760 4575 1795 4675
rect 1955 4575 1990 4675
rect 2010 4575 2045 4675
rect 2205 4575 2240 4675
rect 2260 4575 2295 4675
rect 2455 4575 2490 4675
rect 2510 4575 2545 4675
rect 2705 4575 2740 4675
rect 2760 4575 2795 4675
rect 2955 4575 2990 4675
rect 3010 4575 3045 4675
rect 3205 4575 3240 4675
rect 3260 4575 3295 4675
rect 3455 4575 3490 4675
rect 3510 4575 3545 4675
rect 3705 4575 3740 4675
rect 3760 4575 3795 4675
rect 3955 4575 3990 4675
rect 4010 4575 4045 4675
rect 4205 4575 4240 4675
rect 4260 4575 4295 4675
rect 4455 4575 4490 4675
rect 4510 4575 4545 4675
rect 4705 4575 4740 4675
rect 4760 4575 4795 4675
rect 4955 4575 4990 4675
rect 5010 4575 5045 4675
rect 5205 4575 5240 4675
rect 5260 4575 5295 4675
rect 5455 4575 5490 4675
rect 5510 4575 5545 4675
rect 5705 4575 5740 4675
rect 5760 4575 5795 4675
rect 5955 4575 5990 4675
rect 6010 4575 6045 4675
rect 6205 4575 6240 4675
rect 6260 4575 6295 4675
rect 6455 4575 6490 4675
rect 6510 4575 6545 4675
rect 6705 4575 6740 4675
rect 6760 4575 6795 4675
rect 6955 4575 6990 4675
rect 7010 4575 7045 4675
rect 7205 4575 7240 4675
rect 7260 4575 7295 4675
rect 7455 4575 7490 4675
rect 7510 4575 7545 4675
rect 7705 4575 7740 4675
rect 7760 4575 7795 4675
rect 7955 4575 7990 4675
rect 75 4510 175 4545
rect 325 4510 425 4545
rect 575 4510 675 4545
rect 825 4510 925 4545
rect 1075 4510 1175 4545
rect 1325 4510 1425 4545
rect 1575 4510 1675 4545
rect 1825 4510 1925 4545
rect 2075 4510 2175 4545
rect 2325 4510 2425 4545
rect 2575 4510 2675 4545
rect 2825 4510 2925 4545
rect 3075 4510 3175 4545
rect 3325 4510 3425 4545
rect 3575 4510 3675 4545
rect 3825 4510 3925 4545
rect 4075 4510 4175 4545
rect 4325 4510 4425 4545
rect 4575 4510 4675 4545
rect 4825 4510 4925 4545
rect 5075 4510 5175 4545
rect 5325 4510 5425 4545
rect 5575 4510 5675 4545
rect 5825 4510 5925 4545
rect 6075 4510 6175 4545
rect 6325 4510 6425 4545
rect 6575 4510 6675 4545
rect 6825 4510 6925 4545
rect 7075 4510 7175 4545
rect 7325 4510 7425 4545
rect 7575 4510 7675 4545
rect 7825 4510 7925 4545
rect 75 4455 175 4490
rect 325 4455 425 4490
rect 575 4455 675 4490
rect 825 4455 925 4490
rect 1075 4455 1175 4490
rect 1325 4455 1425 4490
rect 1575 4455 1675 4490
rect 1825 4455 1925 4490
rect 2075 4455 2175 4490
rect 2325 4455 2425 4490
rect 2575 4455 2675 4490
rect 2825 4455 2925 4490
rect 3075 4455 3175 4490
rect 3325 4455 3425 4490
rect 3575 4455 3675 4490
rect 3825 4455 3925 4490
rect 4075 4455 4175 4490
rect 4325 4455 4425 4490
rect 4575 4455 4675 4490
rect 4825 4455 4925 4490
rect 5075 4455 5175 4490
rect 5325 4455 5425 4490
rect 5575 4455 5675 4490
rect 5825 4455 5925 4490
rect 6075 4455 6175 4490
rect 6325 4455 6425 4490
rect 6575 4455 6675 4490
rect 6825 4455 6925 4490
rect 7075 4455 7175 4490
rect 7325 4455 7425 4490
rect 7575 4455 7675 4490
rect 7825 4455 7925 4490
rect 10 4325 45 4425
rect 205 4325 240 4425
rect 260 4325 295 4425
rect 455 4325 490 4425
rect 510 4325 545 4425
rect 705 4325 740 4425
rect 760 4325 795 4425
rect 955 4325 990 4425
rect 1010 4325 1045 4425
rect 1205 4325 1240 4425
rect 1260 4325 1295 4425
rect 1455 4325 1490 4425
rect 1510 4325 1545 4425
rect 1705 4325 1740 4425
rect 1760 4325 1795 4425
rect 1955 4325 1990 4425
rect 2010 4325 2045 4425
rect 2205 4325 2240 4425
rect 2260 4325 2295 4425
rect 2455 4325 2490 4425
rect 2510 4325 2545 4425
rect 2705 4325 2740 4425
rect 2760 4325 2795 4425
rect 2955 4325 2990 4425
rect 3010 4325 3045 4425
rect 3205 4325 3240 4425
rect 3260 4325 3295 4425
rect 3455 4325 3490 4425
rect 3510 4325 3545 4425
rect 3705 4325 3740 4425
rect 3760 4325 3795 4425
rect 3955 4325 3990 4425
rect 4010 4325 4045 4425
rect 4205 4325 4240 4425
rect 4260 4325 4295 4425
rect 4455 4325 4490 4425
rect 4510 4325 4545 4425
rect 4705 4325 4740 4425
rect 4760 4325 4795 4425
rect 4955 4325 4990 4425
rect 5010 4325 5045 4425
rect 5205 4325 5240 4425
rect 5260 4325 5295 4425
rect 5455 4325 5490 4425
rect 5510 4325 5545 4425
rect 5705 4325 5740 4425
rect 5760 4325 5795 4425
rect 5955 4325 5990 4425
rect 6010 4325 6045 4425
rect 6205 4325 6240 4425
rect 6260 4325 6295 4425
rect 6455 4325 6490 4425
rect 6510 4325 6545 4425
rect 6705 4325 6740 4425
rect 6760 4325 6795 4425
rect 6955 4325 6990 4425
rect 7010 4325 7045 4425
rect 7205 4325 7240 4425
rect 7260 4325 7295 4425
rect 7455 4325 7490 4425
rect 7510 4325 7545 4425
rect 7705 4325 7740 4425
rect 7760 4325 7795 4425
rect 7955 4325 7990 4425
rect 75 4260 175 4295
rect 325 4260 425 4295
rect 575 4260 675 4295
rect 825 4260 925 4295
rect 1075 4260 1175 4295
rect 1325 4260 1425 4295
rect 1575 4260 1675 4295
rect 1825 4260 1925 4295
rect 2075 4260 2175 4295
rect 2325 4260 2425 4295
rect 2575 4260 2675 4295
rect 2825 4260 2925 4295
rect 3075 4260 3175 4295
rect 3325 4260 3425 4295
rect 3575 4260 3675 4295
rect 3825 4260 3925 4295
rect 4075 4260 4175 4295
rect 4325 4260 4425 4295
rect 4575 4260 4675 4295
rect 4825 4260 4925 4295
rect 5075 4260 5175 4295
rect 5325 4260 5425 4295
rect 5575 4260 5675 4295
rect 5825 4260 5925 4295
rect 6075 4260 6175 4295
rect 6325 4260 6425 4295
rect 6575 4260 6675 4295
rect 6825 4260 6925 4295
rect 7075 4260 7175 4295
rect 7325 4260 7425 4295
rect 7575 4260 7675 4295
rect 7825 4260 7925 4295
rect 75 4205 175 4240
rect 325 4205 425 4240
rect 575 4205 675 4240
rect 825 4205 925 4240
rect 1075 4205 1175 4240
rect 1325 4205 1425 4240
rect 1575 4205 1675 4240
rect 1825 4205 1925 4240
rect 2075 4205 2175 4240
rect 2325 4205 2425 4240
rect 2575 4205 2675 4240
rect 2825 4205 2925 4240
rect 3075 4205 3175 4240
rect 3325 4205 3425 4240
rect 3575 4205 3675 4240
rect 3825 4205 3925 4240
rect 4075 4205 4175 4240
rect 4325 4205 4425 4240
rect 4575 4205 4675 4240
rect 4825 4205 4925 4240
rect 5075 4205 5175 4240
rect 5325 4205 5425 4240
rect 5575 4205 5675 4240
rect 5825 4205 5925 4240
rect 6075 4205 6175 4240
rect 6325 4205 6425 4240
rect 6575 4205 6675 4240
rect 6825 4205 6925 4240
rect 7075 4205 7175 4240
rect 7325 4205 7425 4240
rect 7575 4205 7675 4240
rect 7825 4205 7925 4240
rect 10 4075 45 4175
rect 205 4075 240 4175
rect 260 4075 295 4175
rect 455 4075 490 4175
rect 510 4075 545 4175
rect 705 4075 740 4175
rect 760 4075 795 4175
rect 955 4075 990 4175
rect 1010 4075 1045 4175
rect 1205 4075 1240 4175
rect 1260 4075 1295 4175
rect 1455 4075 1490 4175
rect 1510 4075 1545 4175
rect 1705 4075 1740 4175
rect 1760 4075 1795 4175
rect 1955 4075 1990 4175
rect 2010 4075 2045 4175
rect 2205 4075 2240 4175
rect 2260 4075 2295 4175
rect 2455 4075 2490 4175
rect 2510 4075 2545 4175
rect 2705 4075 2740 4175
rect 2760 4075 2795 4175
rect 2955 4075 2990 4175
rect 3010 4075 3045 4175
rect 3205 4075 3240 4175
rect 3260 4075 3295 4175
rect 3455 4075 3490 4175
rect 3510 4075 3545 4175
rect 3705 4075 3740 4175
rect 3760 4075 3795 4175
rect 3955 4075 3990 4175
rect 4010 4075 4045 4175
rect 4205 4075 4240 4175
rect 4260 4075 4295 4175
rect 4455 4075 4490 4175
rect 4510 4075 4545 4175
rect 4705 4075 4740 4175
rect 4760 4075 4795 4175
rect 4955 4075 4990 4175
rect 5010 4075 5045 4175
rect 5205 4075 5240 4175
rect 5260 4075 5295 4175
rect 5455 4075 5490 4175
rect 5510 4075 5545 4175
rect 5705 4075 5740 4175
rect 5760 4075 5795 4175
rect 5955 4075 5990 4175
rect 6010 4075 6045 4175
rect 6205 4075 6240 4175
rect 6260 4075 6295 4175
rect 6455 4075 6490 4175
rect 6510 4075 6545 4175
rect 6705 4075 6740 4175
rect 6760 4075 6795 4175
rect 6955 4075 6990 4175
rect 7010 4075 7045 4175
rect 7205 4075 7240 4175
rect 7260 4075 7295 4175
rect 7455 4075 7490 4175
rect 7510 4075 7545 4175
rect 7705 4075 7740 4175
rect 7760 4075 7795 4175
rect 7955 4075 7990 4175
rect 75 4010 175 4045
rect 325 4010 425 4045
rect 575 4010 675 4045
rect 825 4010 925 4045
rect 1075 4010 1175 4045
rect 1325 4010 1425 4045
rect 1575 4010 1675 4045
rect 1825 4010 1925 4045
rect 2075 4010 2175 4045
rect 2325 4010 2425 4045
rect 2575 4010 2675 4045
rect 2825 4010 2925 4045
rect 3075 4010 3175 4045
rect 3325 4010 3425 4045
rect 3575 4010 3675 4045
rect 3825 4010 3925 4045
rect 4075 4010 4175 4045
rect 4325 4010 4425 4045
rect 4575 4010 4675 4045
rect 4825 4010 4925 4045
rect 5075 4010 5175 4045
rect 5325 4010 5425 4045
rect 5575 4010 5675 4045
rect 5825 4010 5925 4045
rect 6075 4010 6175 4045
rect 6325 4010 6425 4045
rect 6575 4010 6675 4045
rect 6825 4010 6925 4045
rect 7075 4010 7175 4045
rect 7325 4010 7425 4045
rect 7575 4010 7675 4045
rect 7825 4010 7925 4045
rect 75 3955 175 3990
rect 325 3955 425 3990
rect 575 3955 675 3990
rect 825 3955 925 3990
rect 1075 3955 1175 3990
rect 1325 3955 1425 3990
rect 1575 3955 1675 3990
rect 1825 3955 1925 3990
rect 2075 3955 2175 3990
rect 2325 3955 2425 3990
rect 2575 3955 2675 3990
rect 2825 3955 2925 3990
rect 3075 3955 3175 3990
rect 3325 3955 3425 3990
rect 3575 3955 3675 3990
rect 3825 3955 3925 3990
rect 4075 3955 4175 3990
rect 4325 3955 4425 3990
rect 4575 3955 4675 3990
rect 4825 3955 4925 3990
rect 5075 3955 5175 3990
rect 5325 3955 5425 3990
rect 5575 3955 5675 3990
rect 5825 3955 5925 3990
rect 6075 3955 6175 3990
rect 6325 3955 6425 3990
rect 6575 3955 6675 3990
rect 6825 3955 6925 3990
rect 7075 3955 7175 3990
rect 7325 3955 7425 3990
rect 7575 3955 7675 3990
rect 7825 3955 7925 3990
rect 10 3825 45 3925
rect 205 3825 240 3925
rect 260 3825 295 3925
rect 455 3825 490 3925
rect 510 3825 545 3925
rect 705 3825 740 3925
rect 760 3825 795 3925
rect 955 3825 990 3925
rect 1010 3825 1045 3925
rect 1205 3825 1240 3925
rect 1260 3825 1295 3925
rect 1455 3825 1490 3925
rect 1510 3825 1545 3925
rect 1705 3825 1740 3925
rect 1760 3825 1795 3925
rect 1955 3825 1990 3925
rect 2010 3825 2045 3925
rect 2205 3825 2240 3925
rect 2260 3825 2295 3925
rect 2455 3825 2490 3925
rect 2510 3825 2545 3925
rect 2705 3825 2740 3925
rect 2760 3825 2795 3925
rect 2955 3825 2990 3925
rect 3010 3825 3045 3925
rect 3205 3825 3240 3925
rect 3260 3825 3295 3925
rect 3455 3825 3490 3925
rect 3510 3825 3545 3925
rect 3705 3825 3740 3925
rect 3760 3825 3795 3925
rect 3955 3825 3990 3925
rect 4010 3825 4045 3925
rect 4205 3825 4240 3925
rect 4260 3825 4295 3925
rect 4455 3825 4490 3925
rect 4510 3825 4545 3925
rect 4705 3825 4740 3925
rect 4760 3825 4795 3925
rect 4955 3825 4990 3925
rect 5010 3825 5045 3925
rect 5205 3825 5240 3925
rect 5260 3825 5295 3925
rect 5455 3825 5490 3925
rect 5510 3825 5545 3925
rect 5705 3825 5740 3925
rect 5760 3825 5795 3925
rect 5955 3825 5990 3925
rect 6010 3825 6045 3925
rect 6205 3825 6240 3925
rect 6260 3825 6295 3925
rect 6455 3825 6490 3925
rect 6510 3825 6545 3925
rect 6705 3825 6740 3925
rect 6760 3825 6795 3925
rect 6955 3825 6990 3925
rect 7010 3825 7045 3925
rect 7205 3825 7240 3925
rect 7260 3825 7295 3925
rect 7455 3825 7490 3925
rect 7510 3825 7545 3925
rect 7705 3825 7740 3925
rect 7760 3825 7795 3925
rect 7955 3825 7990 3925
rect 75 3760 175 3795
rect 325 3760 425 3795
rect 575 3760 675 3795
rect 825 3760 925 3795
rect 1075 3760 1175 3795
rect 1325 3760 1425 3795
rect 1575 3760 1675 3795
rect 1825 3760 1925 3795
rect 2075 3760 2175 3795
rect 2325 3760 2425 3795
rect 2575 3760 2675 3795
rect 2825 3760 2925 3795
rect 3075 3760 3175 3795
rect 3325 3760 3425 3795
rect 3575 3760 3675 3795
rect 3825 3760 3925 3795
rect 4075 3760 4175 3795
rect 4325 3760 4425 3795
rect 4575 3760 4675 3795
rect 4825 3760 4925 3795
rect 5075 3760 5175 3795
rect 5325 3760 5425 3795
rect 5575 3760 5675 3795
rect 5825 3760 5925 3795
rect 6075 3760 6175 3795
rect 6325 3760 6425 3795
rect 6575 3760 6675 3795
rect 6825 3760 6925 3795
rect 7075 3760 7175 3795
rect 7325 3760 7425 3795
rect 7575 3760 7675 3795
rect 7825 3760 7925 3795
rect 75 3705 175 3740
rect 325 3705 425 3740
rect 575 3705 675 3740
rect 825 3705 925 3740
rect 1075 3705 1175 3740
rect 1325 3705 1425 3740
rect 1575 3705 1675 3740
rect 1825 3705 1925 3740
rect 2075 3705 2175 3740
rect 2325 3705 2425 3740
rect 2575 3705 2675 3740
rect 2825 3705 2925 3740
rect 3075 3705 3175 3740
rect 3325 3705 3425 3740
rect 3575 3705 3675 3740
rect 3825 3705 3925 3740
rect 4075 3705 4175 3740
rect 4325 3705 4425 3740
rect 4575 3705 4675 3740
rect 4825 3705 4925 3740
rect 5075 3705 5175 3740
rect 5325 3705 5425 3740
rect 5575 3705 5675 3740
rect 5825 3705 5925 3740
rect 6075 3705 6175 3740
rect 6325 3705 6425 3740
rect 6575 3705 6675 3740
rect 6825 3705 6925 3740
rect 7075 3705 7175 3740
rect 7325 3705 7425 3740
rect 7575 3705 7675 3740
rect 7825 3705 7925 3740
rect 10 3575 45 3675
rect 205 3575 240 3675
rect 260 3575 295 3675
rect 455 3575 490 3675
rect 510 3575 545 3675
rect 705 3575 740 3675
rect 760 3575 795 3675
rect 955 3575 990 3675
rect 1010 3575 1045 3675
rect 1205 3575 1240 3675
rect 1260 3575 1295 3675
rect 1455 3575 1490 3675
rect 1510 3575 1545 3675
rect 1705 3575 1740 3675
rect 1760 3575 1795 3675
rect 1955 3575 1990 3675
rect 2010 3575 2045 3675
rect 2205 3575 2240 3675
rect 2260 3575 2295 3675
rect 2455 3575 2490 3675
rect 2510 3575 2545 3675
rect 2705 3575 2740 3675
rect 2760 3575 2795 3675
rect 2955 3575 2990 3675
rect 3010 3575 3045 3675
rect 3205 3575 3240 3675
rect 3260 3575 3295 3675
rect 3455 3575 3490 3675
rect 3510 3575 3545 3675
rect 3705 3575 3740 3675
rect 3760 3575 3795 3675
rect 3955 3575 3990 3675
rect 4010 3575 4045 3675
rect 4205 3575 4240 3675
rect 4260 3575 4295 3675
rect 4455 3575 4490 3675
rect 4510 3575 4545 3675
rect 4705 3575 4740 3675
rect 4760 3575 4795 3675
rect 4955 3575 4990 3675
rect 5010 3575 5045 3675
rect 5205 3575 5240 3675
rect 5260 3575 5295 3675
rect 5455 3575 5490 3675
rect 5510 3575 5545 3675
rect 5705 3575 5740 3675
rect 5760 3575 5795 3675
rect 5955 3575 5990 3675
rect 6010 3575 6045 3675
rect 6205 3575 6240 3675
rect 6260 3575 6295 3675
rect 6455 3575 6490 3675
rect 6510 3575 6545 3675
rect 6705 3575 6740 3675
rect 6760 3575 6795 3675
rect 6955 3575 6990 3675
rect 7010 3575 7045 3675
rect 7205 3575 7240 3675
rect 7260 3575 7295 3675
rect 7455 3575 7490 3675
rect 7510 3575 7545 3675
rect 7705 3575 7740 3675
rect 7760 3575 7795 3675
rect 7955 3575 7990 3675
rect 75 3510 175 3545
rect 325 3510 425 3545
rect 575 3510 675 3545
rect 825 3510 925 3545
rect 1075 3510 1175 3545
rect 1325 3510 1425 3545
rect 1575 3510 1675 3545
rect 1825 3510 1925 3545
rect 2075 3510 2175 3545
rect 2325 3510 2425 3545
rect 2575 3510 2675 3545
rect 2825 3510 2925 3545
rect 3075 3510 3175 3545
rect 3325 3510 3425 3545
rect 3575 3510 3675 3545
rect 3825 3510 3925 3545
rect 4075 3510 4175 3545
rect 4325 3510 4425 3545
rect 4575 3510 4675 3545
rect 4825 3510 4925 3545
rect 5075 3510 5175 3545
rect 5325 3510 5425 3545
rect 5575 3510 5675 3545
rect 5825 3510 5925 3545
rect 6075 3510 6175 3545
rect 6325 3510 6425 3545
rect 6575 3510 6675 3545
rect 6825 3510 6925 3545
rect 7075 3510 7175 3545
rect 7325 3510 7425 3545
rect 7575 3510 7675 3545
rect 7825 3510 7925 3545
rect 75 3455 175 3490
rect 325 3455 425 3490
rect 575 3455 675 3490
rect 825 3455 925 3490
rect 1075 3455 1175 3490
rect 1325 3455 1425 3490
rect 1575 3455 1675 3490
rect 1825 3455 1925 3490
rect 2075 3455 2175 3490
rect 2325 3455 2425 3490
rect 2575 3455 2675 3490
rect 2825 3455 2925 3490
rect 3075 3455 3175 3490
rect 3325 3455 3425 3490
rect 3575 3455 3675 3490
rect 3825 3455 3925 3490
rect 4075 3455 4175 3490
rect 4325 3455 4425 3490
rect 4575 3455 4675 3490
rect 4825 3455 4925 3490
rect 5075 3455 5175 3490
rect 5325 3455 5425 3490
rect 5575 3455 5675 3490
rect 5825 3455 5925 3490
rect 6075 3455 6175 3490
rect 6325 3455 6425 3490
rect 6575 3455 6675 3490
rect 6825 3455 6925 3490
rect 7075 3455 7175 3490
rect 7325 3455 7425 3490
rect 7575 3455 7675 3490
rect 7825 3455 7925 3490
rect 10 3325 45 3425
rect 205 3325 240 3425
rect 260 3325 295 3425
rect 455 3325 490 3425
rect 510 3325 545 3425
rect 705 3325 740 3425
rect 760 3325 795 3425
rect 955 3325 990 3425
rect 1010 3325 1045 3425
rect 1205 3325 1240 3425
rect 1260 3325 1295 3425
rect 1455 3325 1490 3425
rect 1510 3325 1545 3425
rect 1705 3325 1740 3425
rect 1760 3325 1795 3425
rect 1955 3325 1990 3425
rect 2010 3325 2045 3425
rect 2205 3325 2240 3425
rect 2260 3325 2295 3425
rect 2455 3325 2490 3425
rect 2510 3325 2545 3425
rect 2705 3325 2740 3425
rect 2760 3325 2795 3425
rect 2955 3325 2990 3425
rect 3010 3325 3045 3425
rect 3205 3325 3240 3425
rect 3260 3325 3295 3425
rect 3455 3325 3490 3425
rect 3510 3325 3545 3425
rect 3705 3325 3740 3425
rect 3760 3325 3795 3425
rect 3955 3325 3990 3425
rect 4010 3325 4045 3425
rect 4205 3325 4240 3425
rect 4260 3325 4295 3425
rect 4455 3325 4490 3425
rect 4510 3325 4545 3425
rect 4705 3325 4740 3425
rect 4760 3325 4795 3425
rect 4955 3325 4990 3425
rect 5010 3325 5045 3425
rect 5205 3325 5240 3425
rect 5260 3325 5295 3425
rect 5455 3325 5490 3425
rect 5510 3325 5545 3425
rect 5705 3325 5740 3425
rect 5760 3325 5795 3425
rect 5955 3325 5990 3425
rect 6010 3325 6045 3425
rect 6205 3325 6240 3425
rect 6260 3325 6295 3425
rect 6455 3325 6490 3425
rect 6510 3325 6545 3425
rect 6705 3325 6740 3425
rect 6760 3325 6795 3425
rect 6955 3325 6990 3425
rect 7010 3325 7045 3425
rect 7205 3325 7240 3425
rect 7260 3325 7295 3425
rect 7455 3325 7490 3425
rect 7510 3325 7545 3425
rect 7705 3325 7740 3425
rect 7760 3325 7795 3425
rect 7955 3325 7990 3425
rect 75 3260 175 3295
rect 325 3260 425 3295
rect 575 3260 675 3295
rect 825 3260 925 3295
rect 1075 3260 1175 3295
rect 1325 3260 1425 3295
rect 1575 3260 1675 3295
rect 1825 3260 1925 3295
rect 2075 3260 2175 3295
rect 2325 3260 2425 3295
rect 2575 3260 2675 3295
rect 2825 3260 2925 3295
rect 3075 3260 3175 3295
rect 3325 3260 3425 3295
rect 3575 3260 3675 3295
rect 3825 3260 3925 3295
rect 4075 3260 4175 3295
rect 4325 3260 4425 3295
rect 4575 3260 4675 3295
rect 4825 3260 4925 3295
rect 5075 3260 5175 3295
rect 5325 3260 5425 3295
rect 5575 3260 5675 3295
rect 5825 3260 5925 3295
rect 6075 3260 6175 3295
rect 6325 3260 6425 3295
rect 6575 3260 6675 3295
rect 6825 3260 6925 3295
rect 7075 3260 7175 3295
rect 7325 3260 7425 3295
rect 7575 3260 7675 3295
rect 7825 3260 7925 3295
rect 75 3205 175 3240
rect 325 3205 425 3240
rect 575 3205 675 3240
rect 825 3205 925 3240
rect 1075 3205 1175 3240
rect 1325 3205 1425 3240
rect 1575 3205 1675 3240
rect 1825 3205 1925 3240
rect 2075 3205 2175 3240
rect 2325 3205 2425 3240
rect 2575 3205 2675 3240
rect 2825 3205 2925 3240
rect 3075 3205 3175 3240
rect 3325 3205 3425 3240
rect 3575 3205 3675 3240
rect 3825 3205 3925 3240
rect 4075 3205 4175 3240
rect 4325 3205 4425 3240
rect 4575 3205 4675 3240
rect 4825 3205 4925 3240
rect 5075 3205 5175 3240
rect 5325 3205 5425 3240
rect 5575 3205 5675 3240
rect 5825 3205 5925 3240
rect 6075 3205 6175 3240
rect 6325 3205 6425 3240
rect 6575 3205 6675 3240
rect 6825 3205 6925 3240
rect 7075 3205 7175 3240
rect 7325 3205 7425 3240
rect 7575 3205 7675 3240
rect 7825 3205 7925 3240
rect 10 3075 45 3175
rect 205 3075 240 3175
rect 260 3075 295 3175
rect 455 3075 490 3175
rect 510 3075 545 3175
rect 705 3075 740 3175
rect 760 3075 795 3175
rect 955 3075 990 3175
rect 1010 3075 1045 3175
rect 1205 3075 1240 3175
rect 1260 3075 1295 3175
rect 1455 3075 1490 3175
rect 1510 3075 1545 3175
rect 1705 3075 1740 3175
rect 1760 3075 1795 3175
rect 1955 3075 1990 3175
rect 2010 3075 2045 3175
rect 2205 3075 2240 3175
rect 2260 3075 2295 3175
rect 2455 3075 2490 3175
rect 2510 3075 2545 3175
rect 2705 3075 2740 3175
rect 2760 3075 2795 3175
rect 2955 3075 2990 3175
rect 3010 3075 3045 3175
rect 3205 3075 3240 3175
rect 3260 3075 3295 3175
rect 3455 3075 3490 3175
rect 3510 3075 3545 3175
rect 3705 3075 3740 3175
rect 3760 3075 3795 3175
rect 3955 3075 3990 3175
rect 4010 3075 4045 3175
rect 4205 3075 4240 3175
rect 4260 3075 4295 3175
rect 4455 3075 4490 3175
rect 4510 3075 4545 3175
rect 4705 3075 4740 3175
rect 4760 3075 4795 3175
rect 4955 3075 4990 3175
rect 5010 3075 5045 3175
rect 5205 3075 5240 3175
rect 5260 3075 5295 3175
rect 5455 3075 5490 3175
rect 5510 3075 5545 3175
rect 5705 3075 5740 3175
rect 5760 3075 5795 3175
rect 5955 3075 5990 3175
rect 6010 3075 6045 3175
rect 6205 3075 6240 3175
rect 6260 3075 6295 3175
rect 6455 3075 6490 3175
rect 6510 3075 6545 3175
rect 6705 3075 6740 3175
rect 6760 3075 6795 3175
rect 6955 3075 6990 3175
rect 7010 3075 7045 3175
rect 7205 3075 7240 3175
rect 7260 3075 7295 3175
rect 7455 3075 7490 3175
rect 7510 3075 7545 3175
rect 7705 3075 7740 3175
rect 7760 3075 7795 3175
rect 7955 3075 7990 3175
rect 75 3010 175 3045
rect 325 3010 425 3045
rect 575 3010 675 3045
rect 825 3010 925 3045
rect 1075 3010 1175 3045
rect 1325 3010 1425 3045
rect 1575 3010 1675 3045
rect 1825 3010 1925 3045
rect 2075 3010 2175 3045
rect 2325 3010 2425 3045
rect 2575 3010 2675 3045
rect 2825 3010 2925 3045
rect 3075 3010 3175 3045
rect 3325 3010 3425 3045
rect 3575 3010 3675 3045
rect 3825 3010 3925 3045
rect 4075 3010 4175 3045
rect 4325 3010 4425 3045
rect 4575 3010 4675 3045
rect 4825 3010 4925 3045
rect 5075 3010 5175 3045
rect 5325 3010 5425 3045
rect 5575 3010 5675 3045
rect 5825 3010 5925 3045
rect 6075 3010 6175 3045
rect 6325 3010 6425 3045
rect 6575 3010 6675 3045
rect 6825 3010 6925 3045
rect 7075 3010 7175 3045
rect 7325 3010 7425 3045
rect 7575 3010 7675 3045
rect 7825 3010 7925 3045
rect 75 2955 175 2990
rect 325 2955 425 2990
rect 575 2955 675 2990
rect 825 2955 925 2990
rect 1075 2955 1175 2990
rect 1325 2955 1425 2990
rect 1575 2955 1675 2990
rect 1825 2955 1925 2990
rect 2075 2955 2175 2990
rect 2325 2955 2425 2990
rect 2575 2955 2675 2990
rect 2825 2955 2925 2990
rect 3075 2955 3175 2990
rect 3325 2955 3425 2990
rect 3575 2955 3675 2990
rect 3825 2955 3925 2990
rect 4075 2955 4175 2990
rect 4325 2955 4425 2990
rect 4575 2955 4675 2990
rect 4825 2955 4925 2990
rect 5075 2955 5175 2990
rect 5325 2955 5425 2990
rect 5575 2955 5675 2990
rect 5825 2955 5925 2990
rect 6075 2955 6175 2990
rect 6325 2955 6425 2990
rect 6575 2955 6675 2990
rect 6825 2955 6925 2990
rect 7075 2955 7175 2990
rect 7325 2955 7425 2990
rect 7575 2955 7675 2990
rect 7825 2955 7925 2990
rect 10 2825 45 2925
rect 205 2825 240 2925
rect 260 2825 295 2925
rect 455 2825 490 2925
rect 510 2825 545 2925
rect 705 2825 740 2925
rect 760 2825 795 2925
rect 955 2825 990 2925
rect 1010 2825 1045 2925
rect 1205 2825 1240 2925
rect 1260 2825 1295 2925
rect 1455 2825 1490 2925
rect 1510 2825 1545 2925
rect 1705 2825 1740 2925
rect 1760 2825 1795 2925
rect 1955 2825 1990 2925
rect 2010 2825 2045 2925
rect 2205 2825 2240 2925
rect 2260 2825 2295 2925
rect 2455 2825 2490 2925
rect 2510 2825 2545 2925
rect 2705 2825 2740 2925
rect 2760 2825 2795 2925
rect 2955 2825 2990 2925
rect 3010 2825 3045 2925
rect 3205 2825 3240 2925
rect 3260 2825 3295 2925
rect 3455 2825 3490 2925
rect 3510 2825 3545 2925
rect 3705 2825 3740 2925
rect 3760 2825 3795 2925
rect 3955 2825 3990 2925
rect 4010 2825 4045 2925
rect 4205 2825 4240 2925
rect 4260 2825 4295 2925
rect 4455 2825 4490 2925
rect 4510 2825 4545 2925
rect 4705 2825 4740 2925
rect 4760 2825 4795 2925
rect 4955 2825 4990 2925
rect 5010 2825 5045 2925
rect 5205 2825 5240 2925
rect 5260 2825 5295 2925
rect 5455 2825 5490 2925
rect 5510 2825 5545 2925
rect 5705 2825 5740 2925
rect 5760 2825 5795 2925
rect 5955 2825 5990 2925
rect 6010 2825 6045 2925
rect 6205 2825 6240 2925
rect 6260 2825 6295 2925
rect 6455 2825 6490 2925
rect 6510 2825 6545 2925
rect 6705 2825 6740 2925
rect 6760 2825 6795 2925
rect 6955 2825 6990 2925
rect 7010 2825 7045 2925
rect 7205 2825 7240 2925
rect 7260 2825 7295 2925
rect 7455 2825 7490 2925
rect 7510 2825 7545 2925
rect 7705 2825 7740 2925
rect 7760 2825 7795 2925
rect 7955 2825 7990 2925
rect 75 2760 175 2795
rect 325 2760 425 2795
rect 575 2760 675 2795
rect 825 2760 925 2795
rect 1075 2760 1175 2795
rect 1325 2760 1425 2795
rect 1575 2760 1675 2795
rect 1825 2760 1925 2795
rect 2075 2760 2175 2795
rect 2325 2760 2425 2795
rect 2575 2760 2675 2795
rect 2825 2760 2925 2795
rect 3075 2760 3175 2795
rect 3325 2760 3425 2795
rect 3575 2760 3675 2795
rect 3825 2760 3925 2795
rect 4075 2760 4175 2795
rect 4325 2760 4425 2795
rect 4575 2760 4675 2795
rect 4825 2760 4925 2795
rect 5075 2760 5175 2795
rect 5325 2760 5425 2795
rect 5575 2760 5675 2795
rect 5825 2760 5925 2795
rect 6075 2760 6175 2795
rect 6325 2760 6425 2795
rect 6575 2760 6675 2795
rect 6825 2760 6925 2795
rect 7075 2760 7175 2795
rect 7325 2760 7425 2795
rect 7575 2760 7675 2795
rect 7825 2760 7925 2795
rect 75 2705 175 2740
rect 325 2705 425 2740
rect 575 2705 675 2740
rect 825 2705 925 2740
rect 1075 2705 1175 2740
rect 1325 2705 1425 2740
rect 1575 2705 1675 2740
rect 1825 2705 1925 2740
rect 2075 2705 2175 2740
rect 2325 2705 2425 2740
rect 2575 2705 2675 2740
rect 2825 2705 2925 2740
rect 3075 2705 3175 2740
rect 3325 2705 3425 2740
rect 3575 2705 3675 2740
rect 3825 2705 3925 2740
rect 4075 2705 4175 2740
rect 4325 2705 4425 2740
rect 4575 2705 4675 2740
rect 4825 2705 4925 2740
rect 5075 2705 5175 2740
rect 5325 2705 5425 2740
rect 5575 2705 5675 2740
rect 5825 2705 5925 2740
rect 6075 2705 6175 2740
rect 6325 2705 6425 2740
rect 6575 2705 6675 2740
rect 6825 2705 6925 2740
rect 7075 2705 7175 2740
rect 7325 2705 7425 2740
rect 7575 2705 7675 2740
rect 7825 2705 7925 2740
rect 10 2575 45 2675
rect 205 2575 240 2675
rect 260 2575 295 2675
rect 455 2575 490 2675
rect 510 2575 545 2675
rect 705 2575 740 2675
rect 760 2575 795 2675
rect 955 2575 990 2675
rect 1010 2575 1045 2675
rect 1205 2575 1240 2675
rect 1260 2575 1295 2675
rect 1455 2575 1490 2675
rect 1510 2575 1545 2675
rect 1705 2575 1740 2675
rect 1760 2575 1795 2675
rect 1955 2575 1990 2675
rect 2010 2575 2045 2675
rect 2205 2575 2240 2675
rect 2260 2575 2295 2675
rect 2455 2575 2490 2675
rect 2510 2575 2545 2675
rect 2705 2575 2740 2675
rect 2760 2575 2795 2675
rect 2955 2575 2990 2675
rect 3010 2575 3045 2675
rect 3205 2575 3240 2675
rect 3260 2575 3295 2675
rect 3455 2575 3490 2675
rect 3510 2575 3545 2675
rect 3705 2575 3740 2675
rect 3760 2575 3795 2675
rect 3955 2575 3990 2675
rect 4010 2575 4045 2675
rect 4205 2575 4240 2675
rect 4260 2575 4295 2675
rect 4455 2575 4490 2675
rect 4510 2575 4545 2675
rect 4705 2575 4740 2675
rect 4760 2575 4795 2675
rect 4955 2575 4990 2675
rect 5010 2575 5045 2675
rect 5205 2575 5240 2675
rect 5260 2575 5295 2675
rect 5455 2575 5490 2675
rect 5510 2575 5545 2675
rect 5705 2575 5740 2675
rect 5760 2575 5795 2675
rect 5955 2575 5990 2675
rect 6010 2575 6045 2675
rect 6205 2575 6240 2675
rect 6260 2575 6295 2675
rect 6455 2575 6490 2675
rect 6510 2575 6545 2675
rect 6705 2575 6740 2675
rect 6760 2575 6795 2675
rect 6955 2575 6990 2675
rect 7010 2575 7045 2675
rect 7205 2575 7240 2675
rect 7260 2575 7295 2675
rect 7455 2575 7490 2675
rect 7510 2575 7545 2675
rect 7705 2575 7740 2675
rect 7760 2575 7795 2675
rect 7955 2575 7990 2675
rect 75 2510 175 2545
rect 325 2510 425 2545
rect 575 2510 675 2545
rect 825 2510 925 2545
rect 1075 2510 1175 2545
rect 1325 2510 1425 2545
rect 1575 2510 1675 2545
rect 1825 2510 1925 2545
rect 2075 2510 2175 2545
rect 2325 2510 2425 2545
rect 2575 2510 2675 2545
rect 2825 2510 2925 2545
rect 3075 2510 3175 2545
rect 3325 2510 3425 2545
rect 3575 2510 3675 2545
rect 3825 2510 3925 2545
rect 4075 2510 4175 2545
rect 4325 2510 4425 2545
rect 4575 2510 4675 2545
rect 4825 2510 4925 2545
rect 5075 2510 5175 2545
rect 5325 2510 5425 2545
rect 5575 2510 5675 2545
rect 5825 2510 5925 2545
rect 6075 2510 6175 2545
rect 6325 2510 6425 2545
rect 6575 2510 6675 2545
rect 6825 2510 6925 2545
rect 7075 2510 7175 2545
rect 7325 2510 7425 2545
rect 7575 2510 7675 2545
rect 7825 2510 7925 2545
rect 75 2455 175 2490
rect 325 2455 425 2490
rect 575 2455 675 2490
rect 825 2455 925 2490
rect 1075 2455 1175 2490
rect 1325 2455 1425 2490
rect 1575 2455 1675 2490
rect 1825 2455 1925 2490
rect 2075 2455 2175 2490
rect 2325 2455 2425 2490
rect 2575 2455 2675 2490
rect 2825 2455 2925 2490
rect 3075 2455 3175 2490
rect 3325 2455 3425 2490
rect 3575 2455 3675 2490
rect 3825 2455 3925 2490
rect 4075 2455 4175 2490
rect 4325 2455 4425 2490
rect 4575 2455 4675 2490
rect 4825 2455 4925 2490
rect 5075 2455 5175 2490
rect 5325 2455 5425 2490
rect 5575 2455 5675 2490
rect 5825 2455 5925 2490
rect 6075 2455 6175 2490
rect 6325 2455 6425 2490
rect 6575 2455 6675 2490
rect 6825 2455 6925 2490
rect 7075 2455 7175 2490
rect 7325 2455 7425 2490
rect 7575 2455 7675 2490
rect 7825 2455 7925 2490
rect 10 2325 45 2425
rect 205 2325 240 2425
rect 260 2325 295 2425
rect 455 2325 490 2425
rect 510 2325 545 2425
rect 705 2325 740 2425
rect 760 2325 795 2425
rect 955 2325 990 2425
rect 1010 2325 1045 2425
rect 1205 2325 1240 2425
rect 1260 2325 1295 2425
rect 1455 2325 1490 2425
rect 1510 2325 1545 2425
rect 1705 2325 1740 2425
rect 1760 2325 1795 2425
rect 1955 2325 1990 2425
rect 2010 2325 2045 2425
rect 2205 2325 2240 2425
rect 2260 2325 2295 2425
rect 2455 2325 2490 2425
rect 2510 2325 2545 2425
rect 2705 2325 2740 2425
rect 2760 2325 2795 2425
rect 2955 2325 2990 2425
rect 3010 2325 3045 2425
rect 3205 2325 3240 2425
rect 3260 2325 3295 2425
rect 3455 2325 3490 2425
rect 3510 2325 3545 2425
rect 3705 2325 3740 2425
rect 3760 2325 3795 2425
rect 3955 2325 3990 2425
rect 4010 2325 4045 2425
rect 4205 2325 4240 2425
rect 4260 2325 4295 2425
rect 4455 2325 4490 2425
rect 4510 2325 4545 2425
rect 4705 2325 4740 2425
rect 4760 2325 4795 2425
rect 4955 2325 4990 2425
rect 5010 2325 5045 2425
rect 5205 2325 5240 2425
rect 5260 2325 5295 2425
rect 5455 2325 5490 2425
rect 5510 2325 5545 2425
rect 5705 2325 5740 2425
rect 5760 2325 5795 2425
rect 5955 2325 5990 2425
rect 6010 2325 6045 2425
rect 6205 2325 6240 2425
rect 6260 2325 6295 2425
rect 6455 2325 6490 2425
rect 6510 2325 6545 2425
rect 6705 2325 6740 2425
rect 6760 2325 6795 2425
rect 6955 2325 6990 2425
rect 7010 2325 7045 2425
rect 7205 2325 7240 2425
rect 7260 2325 7295 2425
rect 7455 2325 7490 2425
rect 7510 2325 7545 2425
rect 7705 2325 7740 2425
rect 7760 2325 7795 2425
rect 7955 2325 7990 2425
rect 75 2260 175 2295
rect 325 2260 425 2295
rect 575 2260 675 2295
rect 825 2260 925 2295
rect 1075 2260 1175 2295
rect 1325 2260 1425 2295
rect 1575 2260 1675 2295
rect 1825 2260 1925 2295
rect 2075 2260 2175 2295
rect 2325 2260 2425 2295
rect 2575 2260 2675 2295
rect 2825 2260 2925 2295
rect 3075 2260 3175 2295
rect 3325 2260 3425 2295
rect 3575 2260 3675 2295
rect 3825 2260 3925 2295
rect 4075 2260 4175 2295
rect 4325 2260 4425 2295
rect 4575 2260 4675 2295
rect 4825 2260 4925 2295
rect 5075 2260 5175 2295
rect 5325 2260 5425 2295
rect 5575 2260 5675 2295
rect 5825 2260 5925 2295
rect 6075 2260 6175 2295
rect 6325 2260 6425 2295
rect 6575 2260 6675 2295
rect 6825 2260 6925 2295
rect 7075 2260 7175 2295
rect 7325 2260 7425 2295
rect 7575 2260 7675 2295
rect 7825 2260 7925 2295
rect 75 2205 175 2240
rect 325 2205 425 2240
rect 575 2205 675 2240
rect 825 2205 925 2240
rect 1075 2205 1175 2240
rect 1325 2205 1425 2240
rect 1575 2205 1675 2240
rect 1825 2205 1925 2240
rect 2075 2205 2175 2240
rect 2325 2205 2425 2240
rect 2575 2205 2675 2240
rect 2825 2205 2925 2240
rect 3075 2205 3175 2240
rect 3325 2205 3425 2240
rect 3575 2205 3675 2240
rect 3825 2205 3925 2240
rect 4075 2205 4175 2240
rect 4325 2205 4425 2240
rect 4575 2205 4675 2240
rect 4825 2205 4925 2240
rect 5075 2205 5175 2240
rect 5325 2205 5425 2240
rect 5575 2205 5675 2240
rect 5825 2205 5925 2240
rect 6075 2205 6175 2240
rect 6325 2205 6425 2240
rect 6575 2205 6675 2240
rect 6825 2205 6925 2240
rect 7075 2205 7175 2240
rect 7325 2205 7425 2240
rect 7575 2205 7675 2240
rect 7825 2205 7925 2240
rect 10 2075 45 2175
rect 205 2075 240 2175
rect 260 2075 295 2175
rect 455 2075 490 2175
rect 510 2075 545 2175
rect 705 2075 740 2175
rect 760 2075 795 2175
rect 955 2075 990 2175
rect 1010 2075 1045 2175
rect 1205 2075 1240 2175
rect 1260 2075 1295 2175
rect 1455 2075 1490 2175
rect 1510 2075 1545 2175
rect 1705 2075 1740 2175
rect 1760 2075 1795 2175
rect 1955 2075 1990 2175
rect 2010 2075 2045 2175
rect 2205 2075 2240 2175
rect 2260 2075 2295 2175
rect 2455 2075 2490 2175
rect 2510 2075 2545 2175
rect 2705 2075 2740 2175
rect 2760 2075 2795 2175
rect 2955 2075 2990 2175
rect 3010 2075 3045 2175
rect 3205 2075 3240 2175
rect 3260 2075 3295 2175
rect 3455 2075 3490 2175
rect 3510 2075 3545 2175
rect 3705 2075 3740 2175
rect 3760 2075 3795 2175
rect 3955 2075 3990 2175
rect 4010 2075 4045 2175
rect 4205 2075 4240 2175
rect 4260 2075 4295 2175
rect 4455 2075 4490 2175
rect 4510 2075 4545 2175
rect 4705 2075 4740 2175
rect 4760 2075 4795 2175
rect 4955 2075 4990 2175
rect 5010 2075 5045 2175
rect 5205 2075 5240 2175
rect 5260 2075 5295 2175
rect 5455 2075 5490 2175
rect 5510 2075 5545 2175
rect 5705 2075 5740 2175
rect 5760 2075 5795 2175
rect 5955 2075 5990 2175
rect 6010 2075 6045 2175
rect 6205 2075 6240 2175
rect 6260 2075 6295 2175
rect 6455 2075 6490 2175
rect 6510 2075 6545 2175
rect 6705 2075 6740 2175
rect 6760 2075 6795 2175
rect 6955 2075 6990 2175
rect 7010 2075 7045 2175
rect 7205 2075 7240 2175
rect 7260 2075 7295 2175
rect 7455 2075 7490 2175
rect 7510 2075 7545 2175
rect 7705 2075 7740 2175
rect 7760 2075 7795 2175
rect 7955 2075 7990 2175
rect 75 2010 175 2045
rect 325 2010 425 2045
rect 575 2010 675 2045
rect 825 2010 925 2045
rect 1075 2010 1175 2045
rect 1325 2010 1425 2045
rect 1575 2010 1675 2045
rect 1825 2010 1925 2045
rect 2075 2010 2175 2045
rect 2325 2010 2425 2045
rect 2575 2010 2675 2045
rect 2825 2010 2925 2045
rect 3075 2010 3175 2045
rect 3325 2010 3425 2045
rect 3575 2010 3675 2045
rect 3825 2010 3925 2045
rect 4075 2010 4175 2045
rect 4325 2010 4425 2045
rect 4575 2010 4675 2045
rect 4825 2010 4925 2045
rect 5075 2010 5175 2045
rect 5325 2010 5425 2045
rect 5575 2010 5675 2045
rect 5825 2010 5925 2045
rect 6075 2010 6175 2045
rect 6325 2010 6425 2045
rect 6575 2010 6675 2045
rect 6825 2010 6925 2045
rect 7075 2010 7175 2045
rect 7325 2010 7425 2045
rect 7575 2010 7675 2045
rect 7825 2010 7925 2045
rect 75 1955 175 1990
rect 325 1955 425 1990
rect 575 1955 675 1990
rect 825 1955 925 1990
rect 1075 1955 1175 1990
rect 1325 1955 1425 1990
rect 1575 1955 1675 1990
rect 1825 1955 1925 1990
rect 2075 1955 2175 1990
rect 2325 1955 2425 1990
rect 2575 1955 2675 1990
rect 2825 1955 2925 1990
rect 3075 1955 3175 1990
rect 3325 1955 3425 1990
rect 3575 1955 3675 1990
rect 3825 1955 3925 1990
rect 4075 1955 4175 1990
rect 4325 1955 4425 1990
rect 4575 1955 4675 1990
rect 4825 1955 4925 1990
rect 5075 1955 5175 1990
rect 5325 1955 5425 1990
rect 5575 1955 5675 1990
rect 5825 1955 5925 1990
rect 6075 1955 6175 1990
rect 6325 1955 6425 1990
rect 6575 1955 6675 1990
rect 6825 1955 6925 1990
rect 7075 1955 7175 1990
rect 7325 1955 7425 1990
rect 7575 1955 7675 1990
rect 7825 1955 7925 1990
rect 10 1825 45 1925
rect 205 1825 240 1925
rect 260 1825 295 1925
rect 455 1825 490 1925
rect 510 1825 545 1925
rect 705 1825 740 1925
rect 760 1825 795 1925
rect 955 1825 990 1925
rect 1010 1825 1045 1925
rect 1205 1825 1240 1925
rect 1260 1825 1295 1925
rect 1455 1825 1490 1925
rect 1510 1825 1545 1925
rect 1705 1825 1740 1925
rect 1760 1825 1795 1925
rect 1955 1825 1990 1925
rect 2010 1825 2045 1925
rect 2205 1825 2240 1925
rect 2260 1825 2295 1925
rect 2455 1825 2490 1925
rect 2510 1825 2545 1925
rect 2705 1825 2740 1925
rect 2760 1825 2795 1925
rect 2955 1825 2990 1925
rect 3010 1825 3045 1925
rect 3205 1825 3240 1925
rect 3260 1825 3295 1925
rect 3455 1825 3490 1925
rect 3510 1825 3545 1925
rect 3705 1825 3740 1925
rect 3760 1825 3795 1925
rect 3955 1825 3990 1925
rect 4010 1825 4045 1925
rect 4205 1825 4240 1925
rect 4260 1825 4295 1925
rect 4455 1825 4490 1925
rect 4510 1825 4545 1925
rect 4705 1825 4740 1925
rect 4760 1825 4795 1925
rect 4955 1825 4990 1925
rect 5010 1825 5045 1925
rect 5205 1825 5240 1925
rect 5260 1825 5295 1925
rect 5455 1825 5490 1925
rect 5510 1825 5545 1925
rect 5705 1825 5740 1925
rect 5760 1825 5795 1925
rect 5955 1825 5990 1925
rect 6010 1825 6045 1925
rect 6205 1825 6240 1925
rect 6260 1825 6295 1925
rect 6455 1825 6490 1925
rect 6510 1825 6545 1925
rect 6705 1825 6740 1925
rect 6760 1825 6795 1925
rect 6955 1825 6990 1925
rect 7010 1825 7045 1925
rect 7205 1825 7240 1925
rect 7260 1825 7295 1925
rect 7455 1825 7490 1925
rect 7510 1825 7545 1925
rect 7705 1825 7740 1925
rect 7760 1825 7795 1925
rect 7955 1825 7990 1925
rect 75 1760 175 1795
rect 325 1760 425 1795
rect 575 1760 675 1795
rect 825 1760 925 1795
rect 1075 1760 1175 1795
rect 1325 1760 1425 1795
rect 1575 1760 1675 1795
rect 1825 1760 1925 1795
rect 2075 1760 2175 1795
rect 2325 1760 2425 1795
rect 2575 1760 2675 1795
rect 2825 1760 2925 1795
rect 3075 1760 3175 1795
rect 3325 1760 3425 1795
rect 3575 1760 3675 1795
rect 3825 1760 3925 1795
rect 4075 1760 4175 1795
rect 4325 1760 4425 1795
rect 4575 1760 4675 1795
rect 4825 1760 4925 1795
rect 5075 1760 5175 1795
rect 5325 1760 5425 1795
rect 5575 1760 5675 1795
rect 5825 1760 5925 1795
rect 6075 1760 6175 1795
rect 6325 1760 6425 1795
rect 6575 1760 6675 1795
rect 6825 1760 6925 1795
rect 7075 1760 7175 1795
rect 7325 1760 7425 1795
rect 7575 1760 7675 1795
rect 7825 1760 7925 1795
rect 75 1705 175 1740
rect 325 1705 425 1740
rect 575 1705 675 1740
rect 825 1705 925 1740
rect 1075 1705 1175 1740
rect 1325 1705 1425 1740
rect 1575 1705 1675 1740
rect 1825 1705 1925 1740
rect 2075 1705 2175 1740
rect 2325 1705 2425 1740
rect 2575 1705 2675 1740
rect 2825 1705 2925 1740
rect 3075 1705 3175 1740
rect 3325 1705 3425 1740
rect 3575 1705 3675 1740
rect 3825 1705 3925 1740
rect 4075 1705 4175 1740
rect 4325 1705 4425 1740
rect 4575 1705 4675 1740
rect 4825 1705 4925 1740
rect 5075 1705 5175 1740
rect 5325 1705 5425 1740
rect 5575 1705 5675 1740
rect 5825 1705 5925 1740
rect 6075 1705 6175 1740
rect 6325 1705 6425 1740
rect 6575 1705 6675 1740
rect 6825 1705 6925 1740
rect 7075 1705 7175 1740
rect 7325 1705 7425 1740
rect 7575 1705 7675 1740
rect 7825 1705 7925 1740
rect 10 1575 45 1675
rect 205 1575 240 1675
rect 260 1575 295 1675
rect 455 1575 490 1675
rect 510 1575 545 1675
rect 705 1575 740 1675
rect 760 1575 795 1675
rect 955 1575 990 1675
rect 1010 1575 1045 1675
rect 1205 1575 1240 1675
rect 1260 1575 1295 1675
rect 1455 1575 1490 1675
rect 1510 1575 1545 1675
rect 1705 1575 1740 1675
rect 1760 1575 1795 1675
rect 1955 1575 1990 1675
rect 2010 1575 2045 1675
rect 2205 1575 2240 1675
rect 2260 1575 2295 1675
rect 2455 1575 2490 1675
rect 2510 1575 2545 1675
rect 2705 1575 2740 1675
rect 2760 1575 2795 1675
rect 2955 1575 2990 1675
rect 3010 1575 3045 1675
rect 3205 1575 3240 1675
rect 3260 1575 3295 1675
rect 3455 1575 3490 1675
rect 3510 1575 3545 1675
rect 3705 1575 3740 1675
rect 3760 1575 3795 1675
rect 3955 1575 3990 1675
rect 4010 1575 4045 1675
rect 4205 1575 4240 1675
rect 4260 1575 4295 1675
rect 4455 1575 4490 1675
rect 4510 1575 4545 1675
rect 4705 1575 4740 1675
rect 4760 1575 4795 1675
rect 4955 1575 4990 1675
rect 5010 1575 5045 1675
rect 5205 1575 5240 1675
rect 5260 1575 5295 1675
rect 5455 1575 5490 1675
rect 5510 1575 5545 1675
rect 5705 1575 5740 1675
rect 5760 1575 5795 1675
rect 5955 1575 5990 1675
rect 6010 1575 6045 1675
rect 6205 1575 6240 1675
rect 6260 1575 6295 1675
rect 6455 1575 6490 1675
rect 6510 1575 6545 1675
rect 6705 1575 6740 1675
rect 6760 1575 6795 1675
rect 6955 1575 6990 1675
rect 7010 1575 7045 1675
rect 7205 1575 7240 1675
rect 7260 1575 7295 1675
rect 7455 1575 7490 1675
rect 7510 1575 7545 1675
rect 7705 1575 7740 1675
rect 7760 1575 7795 1675
rect 7955 1575 7990 1675
rect 75 1510 175 1545
rect 325 1510 425 1545
rect 575 1510 675 1545
rect 825 1510 925 1545
rect 1075 1510 1175 1545
rect 1325 1510 1425 1545
rect 1575 1510 1675 1545
rect 1825 1510 1925 1545
rect 2075 1510 2175 1545
rect 2325 1510 2425 1545
rect 2575 1510 2675 1545
rect 2825 1510 2925 1545
rect 3075 1510 3175 1545
rect 3325 1510 3425 1545
rect 3575 1510 3675 1545
rect 3825 1510 3925 1545
rect 4075 1510 4175 1545
rect 4325 1510 4425 1545
rect 4575 1510 4675 1545
rect 4825 1510 4925 1545
rect 5075 1510 5175 1545
rect 5325 1510 5425 1545
rect 5575 1510 5675 1545
rect 5825 1510 5925 1545
rect 6075 1510 6175 1545
rect 6325 1510 6425 1545
rect 6575 1510 6675 1545
rect 6825 1510 6925 1545
rect 7075 1510 7175 1545
rect 7325 1510 7425 1545
rect 7575 1510 7675 1545
rect 7825 1510 7925 1545
rect 75 1455 175 1490
rect 325 1455 425 1490
rect 575 1455 675 1490
rect 825 1455 925 1490
rect 1075 1455 1175 1490
rect 1325 1455 1425 1490
rect 1575 1455 1675 1490
rect 1825 1455 1925 1490
rect 2075 1455 2175 1490
rect 2325 1455 2425 1490
rect 2575 1455 2675 1490
rect 2825 1455 2925 1490
rect 3075 1455 3175 1490
rect 3325 1455 3425 1490
rect 3575 1455 3675 1490
rect 3825 1455 3925 1490
rect 4075 1455 4175 1490
rect 4325 1455 4425 1490
rect 4575 1455 4675 1490
rect 4825 1455 4925 1490
rect 5075 1455 5175 1490
rect 5325 1455 5425 1490
rect 5575 1455 5675 1490
rect 5825 1455 5925 1490
rect 6075 1455 6175 1490
rect 6325 1455 6425 1490
rect 6575 1455 6675 1490
rect 6825 1455 6925 1490
rect 7075 1455 7175 1490
rect 7325 1455 7425 1490
rect 7575 1455 7675 1490
rect 7825 1455 7925 1490
rect 10 1325 45 1425
rect 205 1325 240 1425
rect 260 1325 295 1425
rect 455 1325 490 1425
rect 510 1325 545 1425
rect 705 1325 740 1425
rect 760 1325 795 1425
rect 955 1325 990 1425
rect 1010 1325 1045 1425
rect 1205 1325 1240 1425
rect 1260 1325 1295 1425
rect 1455 1325 1490 1425
rect 1510 1325 1545 1425
rect 1705 1325 1740 1425
rect 1760 1325 1795 1425
rect 1955 1325 1990 1425
rect 2010 1325 2045 1425
rect 2205 1325 2240 1425
rect 2260 1325 2295 1425
rect 2455 1325 2490 1425
rect 2510 1325 2545 1425
rect 2705 1325 2740 1425
rect 2760 1325 2795 1425
rect 2955 1325 2990 1425
rect 3010 1325 3045 1425
rect 3205 1325 3240 1425
rect 3260 1325 3295 1425
rect 3455 1325 3490 1425
rect 3510 1325 3545 1425
rect 3705 1325 3740 1425
rect 3760 1325 3795 1425
rect 3955 1325 3990 1425
rect 4010 1325 4045 1425
rect 4205 1325 4240 1425
rect 4260 1325 4295 1425
rect 4455 1325 4490 1425
rect 4510 1325 4545 1425
rect 4705 1325 4740 1425
rect 4760 1325 4795 1425
rect 4955 1325 4990 1425
rect 5010 1325 5045 1425
rect 5205 1325 5240 1425
rect 5260 1325 5295 1425
rect 5455 1325 5490 1425
rect 5510 1325 5545 1425
rect 5705 1325 5740 1425
rect 5760 1325 5795 1425
rect 5955 1325 5990 1425
rect 6010 1325 6045 1425
rect 6205 1325 6240 1425
rect 6260 1325 6295 1425
rect 6455 1325 6490 1425
rect 6510 1325 6545 1425
rect 6705 1325 6740 1425
rect 6760 1325 6795 1425
rect 6955 1325 6990 1425
rect 7010 1325 7045 1425
rect 7205 1325 7240 1425
rect 7260 1325 7295 1425
rect 7455 1325 7490 1425
rect 7510 1325 7545 1425
rect 7705 1325 7740 1425
rect 7760 1325 7795 1425
rect 7955 1325 7990 1425
rect 75 1260 175 1295
rect 325 1260 425 1295
rect 575 1260 675 1295
rect 825 1260 925 1295
rect 1075 1260 1175 1295
rect 1325 1260 1425 1295
rect 1575 1260 1675 1295
rect 1825 1260 1925 1295
rect 2075 1260 2175 1295
rect 2325 1260 2425 1295
rect 2575 1260 2675 1295
rect 2825 1260 2925 1295
rect 3075 1260 3175 1295
rect 3325 1260 3425 1295
rect 3575 1260 3675 1295
rect 3825 1260 3925 1295
rect 4075 1260 4175 1295
rect 4325 1260 4425 1295
rect 4575 1260 4675 1295
rect 4825 1260 4925 1295
rect 5075 1260 5175 1295
rect 5325 1260 5425 1295
rect 5575 1260 5675 1295
rect 5825 1260 5925 1295
rect 6075 1260 6175 1295
rect 6325 1260 6425 1295
rect 6575 1260 6675 1295
rect 6825 1260 6925 1295
rect 7075 1260 7175 1295
rect 7325 1260 7425 1295
rect 7575 1260 7675 1295
rect 7825 1260 7925 1295
rect 75 1205 175 1240
rect 325 1205 425 1240
rect 575 1205 675 1240
rect 825 1205 925 1240
rect 1075 1205 1175 1240
rect 1325 1205 1425 1240
rect 1575 1205 1675 1240
rect 1825 1205 1925 1240
rect 2075 1205 2175 1240
rect 2325 1205 2425 1240
rect 2575 1205 2675 1240
rect 2825 1205 2925 1240
rect 3075 1205 3175 1240
rect 3325 1205 3425 1240
rect 3575 1205 3675 1240
rect 3825 1205 3925 1240
rect 4075 1205 4175 1240
rect 4325 1205 4425 1240
rect 4575 1205 4675 1240
rect 4825 1205 4925 1240
rect 5075 1205 5175 1240
rect 5325 1205 5425 1240
rect 5575 1205 5675 1240
rect 5825 1205 5925 1240
rect 6075 1205 6175 1240
rect 6325 1205 6425 1240
rect 6575 1205 6675 1240
rect 6825 1205 6925 1240
rect 7075 1205 7175 1240
rect 7325 1205 7425 1240
rect 7575 1205 7675 1240
rect 7825 1205 7925 1240
rect 10 1075 45 1175
rect 205 1075 240 1175
rect 260 1075 295 1175
rect 455 1075 490 1175
rect 510 1075 545 1175
rect 705 1075 740 1175
rect 760 1075 795 1175
rect 955 1075 990 1175
rect 1010 1075 1045 1175
rect 1205 1075 1240 1175
rect 1260 1075 1295 1175
rect 1455 1075 1490 1175
rect 1510 1075 1545 1175
rect 1705 1075 1740 1175
rect 1760 1075 1795 1175
rect 1955 1075 1990 1175
rect 2010 1075 2045 1175
rect 2205 1075 2240 1175
rect 2260 1075 2295 1175
rect 2455 1075 2490 1175
rect 2510 1075 2545 1175
rect 2705 1075 2740 1175
rect 2760 1075 2795 1175
rect 2955 1075 2990 1175
rect 3010 1075 3045 1175
rect 3205 1075 3240 1175
rect 3260 1075 3295 1175
rect 3455 1075 3490 1175
rect 3510 1075 3545 1175
rect 3705 1075 3740 1175
rect 3760 1075 3795 1175
rect 3955 1075 3990 1175
rect 4010 1075 4045 1175
rect 4205 1075 4240 1175
rect 4260 1075 4295 1175
rect 4455 1075 4490 1175
rect 4510 1075 4545 1175
rect 4705 1075 4740 1175
rect 4760 1075 4795 1175
rect 4955 1075 4990 1175
rect 5010 1075 5045 1175
rect 5205 1075 5240 1175
rect 5260 1075 5295 1175
rect 5455 1075 5490 1175
rect 5510 1075 5545 1175
rect 5705 1075 5740 1175
rect 5760 1075 5795 1175
rect 5955 1075 5990 1175
rect 6010 1075 6045 1175
rect 6205 1075 6240 1175
rect 6260 1075 6295 1175
rect 6455 1075 6490 1175
rect 6510 1075 6545 1175
rect 6705 1075 6740 1175
rect 6760 1075 6795 1175
rect 6955 1075 6990 1175
rect 7010 1075 7045 1175
rect 7205 1075 7240 1175
rect 7260 1075 7295 1175
rect 7455 1075 7490 1175
rect 7510 1075 7545 1175
rect 7705 1075 7740 1175
rect 7760 1075 7795 1175
rect 7955 1075 7990 1175
rect 75 1010 175 1045
rect 325 1010 425 1045
rect 575 1010 675 1045
rect 825 1010 925 1045
rect 1075 1010 1175 1045
rect 1325 1010 1425 1045
rect 1575 1010 1675 1045
rect 1825 1010 1925 1045
rect 2075 1010 2175 1045
rect 2325 1010 2425 1045
rect 2575 1010 2675 1045
rect 2825 1010 2925 1045
rect 3075 1010 3175 1045
rect 3325 1010 3425 1045
rect 3575 1010 3675 1045
rect 3825 1010 3925 1045
rect 4075 1010 4175 1045
rect 4325 1010 4425 1045
rect 4575 1010 4675 1045
rect 4825 1010 4925 1045
rect 5075 1010 5175 1045
rect 5325 1010 5425 1045
rect 5575 1010 5675 1045
rect 5825 1010 5925 1045
rect 6075 1010 6175 1045
rect 6325 1010 6425 1045
rect 6575 1010 6675 1045
rect 6825 1010 6925 1045
rect 7075 1010 7175 1045
rect 7325 1010 7425 1045
rect 7575 1010 7675 1045
rect 7825 1010 7925 1045
rect 75 955 175 990
rect 325 955 425 990
rect 575 955 675 990
rect 825 955 925 990
rect 1075 955 1175 990
rect 1325 955 1425 990
rect 1575 955 1675 990
rect 1825 955 1925 990
rect 2075 955 2175 990
rect 2325 955 2425 990
rect 2575 955 2675 990
rect 2825 955 2925 990
rect 3075 955 3175 990
rect 3325 955 3425 990
rect 3575 955 3675 990
rect 3825 955 3925 990
rect 4075 955 4175 990
rect 4325 955 4425 990
rect 4575 955 4675 990
rect 4825 955 4925 990
rect 5075 955 5175 990
rect 5325 955 5425 990
rect 5575 955 5675 990
rect 5825 955 5925 990
rect 6075 955 6175 990
rect 6325 955 6425 990
rect 6575 955 6675 990
rect 6825 955 6925 990
rect 7075 955 7175 990
rect 7325 955 7425 990
rect 7575 955 7675 990
rect 7825 955 7925 990
rect 10 825 45 925
rect 205 825 240 925
rect 260 825 295 925
rect 455 825 490 925
rect 510 825 545 925
rect 705 825 740 925
rect 760 825 795 925
rect 955 825 990 925
rect 1010 825 1045 925
rect 1205 825 1240 925
rect 1260 825 1295 925
rect 1455 825 1490 925
rect 1510 825 1545 925
rect 1705 825 1740 925
rect 1760 825 1795 925
rect 1955 825 1990 925
rect 2010 825 2045 925
rect 2205 825 2240 925
rect 2260 825 2295 925
rect 2455 825 2490 925
rect 2510 825 2545 925
rect 2705 825 2740 925
rect 2760 825 2795 925
rect 2955 825 2990 925
rect 3010 825 3045 925
rect 3205 825 3240 925
rect 3260 825 3295 925
rect 3455 825 3490 925
rect 3510 825 3545 925
rect 3705 825 3740 925
rect 3760 825 3795 925
rect 3955 825 3990 925
rect 4010 825 4045 925
rect 4205 825 4240 925
rect 4260 825 4295 925
rect 4455 825 4490 925
rect 4510 825 4545 925
rect 4705 825 4740 925
rect 4760 825 4795 925
rect 4955 825 4990 925
rect 5010 825 5045 925
rect 5205 825 5240 925
rect 5260 825 5295 925
rect 5455 825 5490 925
rect 5510 825 5545 925
rect 5705 825 5740 925
rect 5760 825 5795 925
rect 5955 825 5990 925
rect 6010 825 6045 925
rect 6205 825 6240 925
rect 6260 825 6295 925
rect 6455 825 6490 925
rect 6510 825 6545 925
rect 6705 825 6740 925
rect 6760 825 6795 925
rect 6955 825 6990 925
rect 7010 825 7045 925
rect 7205 825 7240 925
rect 7260 825 7295 925
rect 7455 825 7490 925
rect 7510 825 7545 925
rect 7705 825 7740 925
rect 7760 825 7795 925
rect 7955 825 7990 925
rect 75 760 175 795
rect 325 760 425 795
rect 575 760 675 795
rect 825 760 925 795
rect 1075 760 1175 795
rect 1325 760 1425 795
rect 1575 760 1675 795
rect 1825 760 1925 795
rect 2075 760 2175 795
rect 2325 760 2425 795
rect 2575 760 2675 795
rect 2825 760 2925 795
rect 3075 760 3175 795
rect 3325 760 3425 795
rect 3575 760 3675 795
rect 3825 760 3925 795
rect 4075 760 4175 795
rect 4325 760 4425 795
rect 4575 760 4675 795
rect 4825 760 4925 795
rect 5075 760 5175 795
rect 5325 760 5425 795
rect 5575 760 5675 795
rect 5825 760 5925 795
rect 6075 760 6175 795
rect 6325 760 6425 795
rect 6575 760 6675 795
rect 6825 760 6925 795
rect 7075 760 7175 795
rect 7325 760 7425 795
rect 7575 760 7675 795
rect 7825 760 7925 795
rect 75 705 175 740
rect 325 705 425 740
rect 575 705 675 740
rect 825 705 925 740
rect 1075 705 1175 740
rect 1325 705 1425 740
rect 1575 705 1675 740
rect 1825 705 1925 740
rect 2075 705 2175 740
rect 2325 705 2425 740
rect 2575 705 2675 740
rect 2825 705 2925 740
rect 3075 705 3175 740
rect 3325 705 3425 740
rect 3575 705 3675 740
rect 3825 705 3925 740
rect 4075 705 4175 740
rect 4325 705 4425 740
rect 4575 705 4675 740
rect 4825 705 4925 740
rect 5075 705 5175 740
rect 5325 705 5425 740
rect 5575 705 5675 740
rect 5825 705 5925 740
rect 6075 705 6175 740
rect 6325 705 6425 740
rect 6575 705 6675 740
rect 6825 705 6925 740
rect 7075 705 7175 740
rect 7325 705 7425 740
rect 7575 705 7675 740
rect 7825 705 7925 740
rect 10 575 45 675
rect 205 575 240 675
rect 260 575 295 675
rect 455 575 490 675
rect 510 575 545 675
rect 705 575 740 675
rect 760 575 795 675
rect 955 575 990 675
rect 1010 575 1045 675
rect 1205 575 1240 675
rect 1260 575 1295 675
rect 1455 575 1490 675
rect 1510 575 1545 675
rect 1705 575 1740 675
rect 1760 575 1795 675
rect 1955 575 1990 675
rect 2010 575 2045 675
rect 2205 575 2240 675
rect 2260 575 2295 675
rect 2455 575 2490 675
rect 2510 575 2545 675
rect 2705 575 2740 675
rect 2760 575 2795 675
rect 2955 575 2990 675
rect 3010 575 3045 675
rect 3205 575 3240 675
rect 3260 575 3295 675
rect 3455 575 3490 675
rect 3510 575 3545 675
rect 3705 575 3740 675
rect 3760 575 3795 675
rect 3955 575 3990 675
rect 4010 575 4045 675
rect 4205 575 4240 675
rect 4260 575 4295 675
rect 4455 575 4490 675
rect 4510 575 4545 675
rect 4705 575 4740 675
rect 4760 575 4795 675
rect 4955 575 4990 675
rect 5010 575 5045 675
rect 5205 575 5240 675
rect 5260 575 5295 675
rect 5455 575 5490 675
rect 5510 575 5545 675
rect 5705 575 5740 675
rect 5760 575 5795 675
rect 5955 575 5990 675
rect 6010 575 6045 675
rect 6205 575 6240 675
rect 6260 575 6295 675
rect 6455 575 6490 675
rect 6510 575 6545 675
rect 6705 575 6740 675
rect 6760 575 6795 675
rect 6955 575 6990 675
rect 7010 575 7045 675
rect 7205 575 7240 675
rect 7260 575 7295 675
rect 7455 575 7490 675
rect 7510 575 7545 675
rect 7705 575 7740 675
rect 7760 575 7795 675
rect 7955 575 7990 675
rect 75 510 175 545
rect 325 510 425 545
rect 575 510 675 545
rect 825 510 925 545
rect 1075 510 1175 545
rect 1325 510 1425 545
rect 1575 510 1675 545
rect 1825 510 1925 545
rect 2075 510 2175 545
rect 2325 510 2425 545
rect 2575 510 2675 545
rect 2825 510 2925 545
rect 3075 510 3175 545
rect 3325 510 3425 545
rect 3575 510 3675 545
rect 3825 510 3925 545
rect 4075 510 4175 545
rect 4325 510 4425 545
rect 4575 510 4675 545
rect 4825 510 4925 545
rect 5075 510 5175 545
rect 5325 510 5425 545
rect 5575 510 5675 545
rect 5825 510 5925 545
rect 6075 510 6175 545
rect 6325 510 6425 545
rect 6575 510 6675 545
rect 6825 510 6925 545
rect 7075 510 7175 545
rect 7325 510 7425 545
rect 7575 510 7675 545
rect 7825 510 7925 545
rect 75 455 175 490
rect 325 455 425 490
rect 575 455 675 490
rect 825 455 925 490
rect 1075 455 1175 490
rect 1325 455 1425 490
rect 1575 455 1675 490
rect 1825 455 1925 490
rect 2075 455 2175 490
rect 2325 455 2425 490
rect 2575 455 2675 490
rect 2825 455 2925 490
rect 3075 455 3175 490
rect 3325 455 3425 490
rect 3575 455 3675 490
rect 3825 455 3925 490
rect 4075 455 4175 490
rect 4325 455 4425 490
rect 4575 455 4675 490
rect 4825 455 4925 490
rect 5075 455 5175 490
rect 5325 455 5425 490
rect 5575 455 5675 490
rect 5825 455 5925 490
rect 6075 455 6175 490
rect 6325 455 6425 490
rect 6575 455 6675 490
rect 6825 455 6925 490
rect 7075 455 7175 490
rect 7325 455 7425 490
rect 7575 455 7675 490
rect 7825 455 7925 490
rect 10 325 45 425
rect 205 325 240 425
rect 260 325 295 425
rect 455 325 490 425
rect 510 325 545 425
rect 705 325 740 425
rect 760 325 795 425
rect 955 325 990 425
rect 1010 325 1045 425
rect 1205 325 1240 425
rect 1260 325 1295 425
rect 1455 325 1490 425
rect 1510 325 1545 425
rect 1705 325 1740 425
rect 1760 325 1795 425
rect 1955 325 1990 425
rect 2010 325 2045 425
rect 2205 325 2240 425
rect 2260 325 2295 425
rect 2455 325 2490 425
rect 2510 325 2545 425
rect 2705 325 2740 425
rect 2760 325 2795 425
rect 2955 325 2990 425
rect 3010 325 3045 425
rect 3205 325 3240 425
rect 3260 325 3295 425
rect 3455 325 3490 425
rect 3510 325 3545 425
rect 3705 325 3740 425
rect 3760 325 3795 425
rect 3955 325 3990 425
rect 4010 325 4045 425
rect 4205 325 4240 425
rect 4260 325 4295 425
rect 4455 325 4490 425
rect 4510 325 4545 425
rect 4705 325 4740 425
rect 4760 325 4795 425
rect 4955 325 4990 425
rect 5010 325 5045 425
rect 5205 325 5240 425
rect 5260 325 5295 425
rect 5455 325 5490 425
rect 5510 325 5545 425
rect 5705 325 5740 425
rect 5760 325 5795 425
rect 5955 325 5990 425
rect 6010 325 6045 425
rect 6205 325 6240 425
rect 6260 325 6295 425
rect 6455 325 6490 425
rect 6510 325 6545 425
rect 6705 325 6740 425
rect 6760 325 6795 425
rect 6955 325 6990 425
rect 7010 325 7045 425
rect 7205 325 7240 425
rect 7260 325 7295 425
rect 7455 325 7490 425
rect 7510 325 7545 425
rect 7705 325 7740 425
rect 7760 325 7795 425
rect 7955 325 7990 425
rect 75 260 175 295
rect 325 260 425 295
rect 575 260 675 295
rect 825 260 925 295
rect 1075 260 1175 295
rect 1325 260 1425 295
rect 1575 260 1675 295
rect 1825 260 1925 295
rect 2075 260 2175 295
rect 2325 260 2425 295
rect 2575 260 2675 295
rect 2825 260 2925 295
rect 3075 260 3175 295
rect 3325 260 3425 295
rect 3575 260 3675 295
rect 3825 260 3925 295
rect 4075 260 4175 295
rect 4325 260 4425 295
rect 4575 260 4675 295
rect 4825 260 4925 295
rect 5075 260 5175 295
rect 5325 260 5425 295
rect 5575 260 5675 295
rect 5825 260 5925 295
rect 6075 260 6175 295
rect 6325 260 6425 295
rect 6575 260 6675 295
rect 6825 260 6925 295
rect 7075 260 7175 295
rect 7325 260 7425 295
rect 7575 260 7675 295
rect 7825 260 7925 295
rect 75 205 175 240
rect 325 205 425 240
rect 575 205 675 240
rect 825 205 925 240
rect 1075 205 1175 240
rect 1325 205 1425 240
rect 1575 205 1675 240
rect 1825 205 1925 240
rect 2075 205 2175 240
rect 2325 205 2425 240
rect 2575 205 2675 240
rect 2825 205 2925 240
rect 3075 205 3175 240
rect 3325 205 3425 240
rect 3575 205 3675 240
rect 3825 205 3925 240
rect 4075 205 4175 240
rect 4325 205 4425 240
rect 4575 205 4675 240
rect 4825 205 4925 240
rect 5075 205 5175 240
rect 5325 205 5425 240
rect 5575 205 5675 240
rect 5825 205 5925 240
rect 6075 205 6175 240
rect 6325 205 6425 240
rect 6575 205 6675 240
rect 6825 205 6925 240
rect 7075 205 7175 240
rect 7325 205 7425 240
rect 7575 205 7675 240
rect 7825 205 7925 240
rect 10 75 45 175
rect 205 75 240 175
rect 260 75 295 175
rect 455 75 490 175
rect 510 75 545 175
rect 705 75 740 175
rect 760 75 795 175
rect 955 75 990 175
rect 1010 75 1045 175
rect 1205 75 1240 175
rect 1260 75 1295 175
rect 1455 75 1490 175
rect 1510 75 1545 175
rect 1705 75 1740 175
rect 1760 75 1795 175
rect 1955 75 1990 175
rect 2010 75 2045 175
rect 2205 75 2240 175
rect 2260 75 2295 175
rect 2455 75 2490 175
rect 2510 75 2545 175
rect 2705 75 2740 175
rect 2760 75 2795 175
rect 2955 75 2990 175
rect 3010 75 3045 175
rect 3205 75 3240 175
rect 3260 75 3295 175
rect 3455 75 3490 175
rect 3510 75 3545 175
rect 3705 75 3740 175
rect 3760 75 3795 175
rect 3955 75 3990 175
rect 4010 75 4045 175
rect 4205 75 4240 175
rect 4260 75 4295 175
rect 4455 75 4490 175
rect 4510 75 4545 175
rect 4705 75 4740 175
rect 4760 75 4795 175
rect 4955 75 4990 175
rect 5010 75 5045 175
rect 5205 75 5240 175
rect 5260 75 5295 175
rect 5455 75 5490 175
rect 5510 75 5545 175
rect 5705 75 5740 175
rect 5760 75 5795 175
rect 5955 75 5990 175
rect 6010 75 6045 175
rect 6205 75 6240 175
rect 6260 75 6295 175
rect 6455 75 6490 175
rect 6510 75 6545 175
rect 6705 75 6740 175
rect 6760 75 6795 175
rect 6955 75 6990 175
rect 7010 75 7045 175
rect 7205 75 7240 175
rect 7260 75 7295 175
rect 7455 75 7490 175
rect 7510 75 7545 175
rect 7705 75 7740 175
rect 7760 75 7795 175
rect 7955 75 7990 175
rect 75 10 175 45
rect 325 10 425 45
rect 575 10 675 45
rect 825 10 925 45
rect 1075 10 1175 45
rect 1325 10 1425 45
rect 1575 10 1675 45
rect 1825 10 1925 45
rect 2075 10 2175 45
rect 2325 10 2425 45
rect 2575 10 2675 45
rect 2825 10 2925 45
rect 3075 10 3175 45
rect 3325 10 3425 45
rect 3575 10 3675 45
rect 3825 10 3925 45
rect 4075 10 4175 45
rect 4325 10 4425 45
rect 4575 10 4675 45
rect 4825 10 4925 45
rect 5075 10 5175 45
rect 5325 10 5425 45
rect 5575 10 5675 45
rect 5825 10 5925 45
rect 6075 10 6175 45
rect 6325 10 6425 45
rect 6575 10 6675 45
rect 6825 10 6925 45
rect 7075 10 7175 45
rect 7325 10 7425 45
rect 7575 10 7675 45
rect 7825 10 7925 45
<< metal2 >>
rect 70 7990 180 8000
rect 70 7955 75 7990
rect 175 7955 180 7990
rect 70 7930 180 7955
rect 320 7990 430 8000
rect 320 7955 325 7990
rect 425 7955 430 7990
rect 320 7930 430 7955
rect 570 7990 680 8000
rect 570 7955 575 7990
rect 675 7955 680 7990
rect 570 7930 680 7955
rect 820 7990 930 8000
rect 820 7955 825 7990
rect 925 7955 930 7990
rect 820 7930 930 7955
rect 1070 7990 1180 8000
rect 1070 7955 1075 7990
rect 1175 7955 1180 7990
rect 1070 7930 1180 7955
rect 1320 7990 1430 8000
rect 1320 7955 1325 7990
rect 1425 7955 1430 7990
rect 1320 7930 1430 7955
rect 1570 7990 1680 8000
rect 1570 7955 1575 7990
rect 1675 7955 1680 7990
rect 1570 7930 1680 7955
rect 1820 7990 1930 8000
rect 1820 7955 1825 7990
rect 1925 7955 1930 7990
rect 1820 7930 1930 7955
rect 2070 7990 2180 8000
rect 2070 7955 2075 7990
rect 2175 7955 2180 7990
rect 2070 7930 2180 7955
rect 2320 7990 2430 8000
rect 2320 7955 2325 7990
rect 2425 7955 2430 7990
rect 2320 7930 2430 7955
rect 2570 7990 2680 8000
rect 2570 7955 2575 7990
rect 2675 7955 2680 7990
rect 2570 7930 2680 7955
rect 2820 7990 2930 8000
rect 2820 7955 2825 7990
rect 2925 7955 2930 7990
rect 2820 7930 2930 7955
rect 3070 7990 3180 8000
rect 3070 7955 3075 7990
rect 3175 7955 3180 7990
rect 3070 7930 3180 7955
rect 3320 7990 3430 8000
rect 3320 7955 3325 7990
rect 3425 7955 3430 7990
rect 3320 7930 3430 7955
rect 3570 7990 3680 8000
rect 3570 7955 3575 7990
rect 3675 7955 3680 7990
rect 3570 7930 3680 7955
rect 3820 7990 3930 8000
rect 3820 7955 3825 7990
rect 3925 7955 3930 7990
rect 3820 7930 3930 7955
rect 4070 7990 4180 8000
rect 4070 7955 4075 7990
rect 4175 7955 4180 7990
rect 4070 7930 4180 7955
rect 4320 7990 4430 8000
rect 4320 7955 4325 7990
rect 4425 7955 4430 7990
rect 4320 7930 4430 7955
rect 4570 7990 4680 8000
rect 4570 7955 4575 7990
rect 4675 7955 4680 7990
rect 4570 7930 4680 7955
rect 4820 7990 4930 8000
rect 4820 7955 4825 7990
rect 4925 7955 4930 7990
rect 4820 7930 4930 7955
rect 5070 7990 5180 8000
rect 5070 7955 5075 7990
rect 5175 7955 5180 7990
rect 5070 7930 5180 7955
rect 5320 7990 5430 8000
rect 5320 7955 5325 7990
rect 5425 7955 5430 7990
rect 5320 7930 5430 7955
rect 5570 7990 5680 8000
rect 5570 7955 5575 7990
rect 5675 7955 5680 7990
rect 5570 7930 5680 7955
rect 5820 7990 5930 8000
rect 5820 7955 5825 7990
rect 5925 7955 5930 7990
rect 5820 7930 5930 7955
rect 6070 7990 6180 8000
rect 6070 7955 6075 7990
rect 6175 7955 6180 7990
rect 6070 7930 6180 7955
rect 6320 7990 6430 8000
rect 6320 7955 6325 7990
rect 6425 7955 6430 7990
rect 6320 7930 6430 7955
rect 6570 7990 6680 8000
rect 6570 7955 6575 7990
rect 6675 7955 6680 7990
rect 6570 7930 6680 7955
rect 6820 7990 6930 8000
rect 6820 7955 6825 7990
rect 6925 7955 6930 7990
rect 6820 7930 6930 7955
rect 7070 7990 7180 8000
rect 7070 7955 7075 7990
rect 7175 7955 7180 7990
rect 7070 7930 7180 7955
rect 7320 7990 7430 8000
rect 7320 7955 7325 7990
rect 7425 7955 7430 7990
rect 7320 7930 7430 7955
rect 7570 7990 7680 8000
rect 7570 7955 7575 7990
rect 7675 7955 7680 7990
rect 7570 7930 7680 7955
rect 7820 7990 7930 8000
rect 7820 7955 7825 7990
rect 7925 7955 7930 7990
rect 7820 7930 7930 7955
rect 0 7925 8000 7930
rect 0 7825 10 7925
rect 45 7825 205 7925
rect 240 7825 260 7925
rect 295 7825 455 7925
rect 490 7825 510 7925
rect 545 7825 705 7925
rect 740 7825 760 7925
rect 795 7825 955 7925
rect 990 7825 1010 7925
rect 1045 7825 1205 7925
rect 1240 7825 1260 7925
rect 1295 7825 1455 7925
rect 1490 7825 1510 7925
rect 1545 7825 1705 7925
rect 1740 7825 1760 7925
rect 1795 7825 1955 7925
rect 1990 7825 2010 7925
rect 2045 7825 2205 7925
rect 2240 7825 2260 7925
rect 2295 7825 2455 7925
rect 2490 7825 2510 7925
rect 2545 7825 2705 7925
rect 2740 7825 2760 7925
rect 2795 7825 2955 7925
rect 2990 7825 3010 7925
rect 3045 7825 3205 7925
rect 3240 7825 3260 7925
rect 3295 7825 3455 7925
rect 3490 7825 3510 7925
rect 3545 7825 3705 7925
rect 3740 7825 3760 7925
rect 3795 7825 3955 7925
rect 3990 7825 4010 7925
rect 4045 7825 4205 7925
rect 4240 7825 4260 7925
rect 4295 7825 4455 7925
rect 4490 7825 4510 7925
rect 4545 7825 4705 7925
rect 4740 7825 4760 7925
rect 4795 7825 4955 7925
rect 4990 7825 5010 7925
rect 5045 7825 5205 7925
rect 5240 7825 5260 7925
rect 5295 7825 5455 7925
rect 5490 7825 5510 7925
rect 5545 7825 5705 7925
rect 5740 7825 5760 7925
rect 5795 7825 5955 7925
rect 5990 7825 6010 7925
rect 6045 7825 6205 7925
rect 6240 7825 6260 7925
rect 6295 7825 6455 7925
rect 6490 7825 6510 7925
rect 6545 7825 6705 7925
rect 6740 7825 6760 7925
rect 6795 7825 6955 7925
rect 6990 7825 7010 7925
rect 7045 7825 7205 7925
rect 7240 7825 7260 7925
rect 7295 7825 7455 7925
rect 7490 7825 7510 7925
rect 7545 7825 7705 7925
rect 7740 7825 7760 7925
rect 7795 7825 7955 7925
rect 7990 7825 8000 7925
rect 0 7820 8000 7825
rect 70 7795 180 7820
rect 70 7760 75 7795
rect 175 7760 180 7795
rect 70 7740 180 7760
rect 70 7705 75 7740
rect 175 7705 180 7740
rect 70 7680 180 7705
rect 320 7795 430 7820
rect 320 7760 325 7795
rect 425 7760 430 7795
rect 320 7740 430 7760
rect 320 7705 325 7740
rect 425 7705 430 7740
rect 320 7680 430 7705
rect 570 7795 680 7820
rect 570 7760 575 7795
rect 675 7760 680 7795
rect 570 7740 680 7760
rect 570 7705 575 7740
rect 675 7705 680 7740
rect 570 7680 680 7705
rect 820 7795 930 7820
rect 820 7760 825 7795
rect 925 7760 930 7795
rect 820 7740 930 7760
rect 820 7705 825 7740
rect 925 7705 930 7740
rect 820 7680 930 7705
rect 1070 7795 1180 7820
rect 1070 7760 1075 7795
rect 1175 7760 1180 7795
rect 1070 7740 1180 7760
rect 1070 7705 1075 7740
rect 1175 7705 1180 7740
rect 1070 7680 1180 7705
rect 1320 7795 1430 7820
rect 1320 7760 1325 7795
rect 1425 7760 1430 7795
rect 1320 7740 1430 7760
rect 1320 7705 1325 7740
rect 1425 7705 1430 7740
rect 1320 7680 1430 7705
rect 1570 7795 1680 7820
rect 1570 7760 1575 7795
rect 1675 7760 1680 7795
rect 1570 7740 1680 7760
rect 1570 7705 1575 7740
rect 1675 7705 1680 7740
rect 1570 7680 1680 7705
rect 1820 7795 1930 7820
rect 1820 7760 1825 7795
rect 1925 7760 1930 7795
rect 1820 7740 1930 7760
rect 1820 7705 1825 7740
rect 1925 7705 1930 7740
rect 1820 7680 1930 7705
rect 2070 7795 2180 7820
rect 2070 7760 2075 7795
rect 2175 7760 2180 7795
rect 2070 7740 2180 7760
rect 2070 7705 2075 7740
rect 2175 7705 2180 7740
rect 2070 7680 2180 7705
rect 2320 7795 2430 7820
rect 2320 7760 2325 7795
rect 2425 7760 2430 7795
rect 2320 7740 2430 7760
rect 2320 7705 2325 7740
rect 2425 7705 2430 7740
rect 2320 7680 2430 7705
rect 2570 7795 2680 7820
rect 2570 7760 2575 7795
rect 2675 7760 2680 7795
rect 2570 7740 2680 7760
rect 2570 7705 2575 7740
rect 2675 7705 2680 7740
rect 2570 7680 2680 7705
rect 2820 7795 2930 7820
rect 2820 7760 2825 7795
rect 2925 7760 2930 7795
rect 2820 7740 2930 7760
rect 2820 7705 2825 7740
rect 2925 7705 2930 7740
rect 2820 7680 2930 7705
rect 3070 7795 3180 7820
rect 3070 7760 3075 7795
rect 3175 7760 3180 7795
rect 3070 7740 3180 7760
rect 3070 7705 3075 7740
rect 3175 7705 3180 7740
rect 3070 7680 3180 7705
rect 3320 7795 3430 7820
rect 3320 7760 3325 7795
rect 3425 7760 3430 7795
rect 3320 7740 3430 7760
rect 3320 7705 3325 7740
rect 3425 7705 3430 7740
rect 3320 7680 3430 7705
rect 3570 7795 3680 7820
rect 3570 7760 3575 7795
rect 3675 7760 3680 7795
rect 3570 7740 3680 7760
rect 3570 7705 3575 7740
rect 3675 7705 3680 7740
rect 3570 7680 3680 7705
rect 3820 7795 3930 7820
rect 3820 7760 3825 7795
rect 3925 7760 3930 7795
rect 3820 7740 3930 7760
rect 3820 7705 3825 7740
rect 3925 7705 3930 7740
rect 3820 7680 3930 7705
rect 4070 7795 4180 7820
rect 4070 7760 4075 7795
rect 4175 7760 4180 7795
rect 4070 7740 4180 7760
rect 4070 7705 4075 7740
rect 4175 7705 4180 7740
rect 4070 7680 4180 7705
rect 4320 7795 4430 7820
rect 4320 7760 4325 7795
rect 4425 7760 4430 7795
rect 4320 7740 4430 7760
rect 4320 7705 4325 7740
rect 4425 7705 4430 7740
rect 4320 7680 4430 7705
rect 4570 7795 4680 7820
rect 4570 7760 4575 7795
rect 4675 7760 4680 7795
rect 4570 7740 4680 7760
rect 4570 7705 4575 7740
rect 4675 7705 4680 7740
rect 4570 7680 4680 7705
rect 4820 7795 4930 7820
rect 4820 7760 4825 7795
rect 4925 7760 4930 7795
rect 4820 7740 4930 7760
rect 4820 7705 4825 7740
rect 4925 7705 4930 7740
rect 4820 7680 4930 7705
rect 5070 7795 5180 7820
rect 5070 7760 5075 7795
rect 5175 7760 5180 7795
rect 5070 7740 5180 7760
rect 5070 7705 5075 7740
rect 5175 7705 5180 7740
rect 5070 7680 5180 7705
rect 5320 7795 5430 7820
rect 5320 7760 5325 7795
rect 5425 7760 5430 7795
rect 5320 7740 5430 7760
rect 5320 7705 5325 7740
rect 5425 7705 5430 7740
rect 5320 7680 5430 7705
rect 5570 7795 5680 7820
rect 5570 7760 5575 7795
rect 5675 7760 5680 7795
rect 5570 7740 5680 7760
rect 5570 7705 5575 7740
rect 5675 7705 5680 7740
rect 5570 7680 5680 7705
rect 5820 7795 5930 7820
rect 5820 7760 5825 7795
rect 5925 7760 5930 7795
rect 5820 7740 5930 7760
rect 5820 7705 5825 7740
rect 5925 7705 5930 7740
rect 5820 7680 5930 7705
rect 6070 7795 6180 7820
rect 6070 7760 6075 7795
rect 6175 7760 6180 7795
rect 6070 7740 6180 7760
rect 6070 7705 6075 7740
rect 6175 7705 6180 7740
rect 6070 7680 6180 7705
rect 6320 7795 6430 7820
rect 6320 7760 6325 7795
rect 6425 7760 6430 7795
rect 6320 7740 6430 7760
rect 6320 7705 6325 7740
rect 6425 7705 6430 7740
rect 6320 7680 6430 7705
rect 6570 7795 6680 7820
rect 6570 7760 6575 7795
rect 6675 7760 6680 7795
rect 6570 7740 6680 7760
rect 6570 7705 6575 7740
rect 6675 7705 6680 7740
rect 6570 7680 6680 7705
rect 6820 7795 6930 7820
rect 6820 7760 6825 7795
rect 6925 7760 6930 7795
rect 6820 7740 6930 7760
rect 6820 7705 6825 7740
rect 6925 7705 6930 7740
rect 6820 7680 6930 7705
rect 7070 7795 7180 7820
rect 7070 7760 7075 7795
rect 7175 7760 7180 7795
rect 7070 7740 7180 7760
rect 7070 7705 7075 7740
rect 7175 7705 7180 7740
rect 7070 7680 7180 7705
rect 7320 7795 7430 7820
rect 7320 7760 7325 7795
rect 7425 7760 7430 7795
rect 7320 7740 7430 7760
rect 7320 7705 7325 7740
rect 7425 7705 7430 7740
rect 7320 7680 7430 7705
rect 7570 7795 7680 7820
rect 7570 7760 7575 7795
rect 7675 7760 7680 7795
rect 7570 7740 7680 7760
rect 7570 7705 7575 7740
rect 7675 7705 7680 7740
rect 7570 7680 7680 7705
rect 7820 7795 7930 7820
rect 7820 7760 7825 7795
rect 7925 7760 7930 7795
rect 7820 7740 7930 7760
rect 7820 7705 7825 7740
rect 7925 7705 7930 7740
rect 7820 7680 7930 7705
rect 0 7675 8000 7680
rect 0 7575 10 7675
rect 45 7575 205 7675
rect 240 7575 260 7675
rect 295 7575 455 7675
rect 490 7575 510 7675
rect 545 7575 705 7675
rect 740 7575 760 7675
rect 795 7575 955 7675
rect 990 7575 1010 7675
rect 1045 7575 1205 7675
rect 1240 7575 1260 7675
rect 1295 7575 1455 7675
rect 1490 7575 1510 7675
rect 1545 7575 1705 7675
rect 1740 7575 1760 7675
rect 1795 7575 1955 7675
rect 1990 7575 2010 7675
rect 2045 7575 2205 7675
rect 2240 7575 2260 7675
rect 2295 7575 2455 7675
rect 2490 7575 2510 7675
rect 2545 7575 2705 7675
rect 2740 7575 2760 7675
rect 2795 7575 2955 7675
rect 2990 7575 3010 7675
rect 3045 7575 3205 7675
rect 3240 7575 3260 7675
rect 3295 7575 3455 7675
rect 3490 7575 3510 7675
rect 3545 7575 3705 7675
rect 3740 7575 3760 7675
rect 3795 7575 3955 7675
rect 3990 7575 4010 7675
rect 4045 7575 4205 7675
rect 4240 7575 4260 7675
rect 4295 7575 4455 7675
rect 4490 7575 4510 7675
rect 4545 7575 4705 7675
rect 4740 7575 4760 7675
rect 4795 7575 4955 7675
rect 4990 7575 5010 7675
rect 5045 7575 5205 7675
rect 5240 7575 5260 7675
rect 5295 7575 5455 7675
rect 5490 7575 5510 7675
rect 5545 7575 5705 7675
rect 5740 7575 5760 7675
rect 5795 7575 5955 7675
rect 5990 7575 6010 7675
rect 6045 7575 6205 7675
rect 6240 7575 6260 7675
rect 6295 7575 6455 7675
rect 6490 7575 6510 7675
rect 6545 7575 6705 7675
rect 6740 7575 6760 7675
rect 6795 7575 6955 7675
rect 6990 7575 7010 7675
rect 7045 7575 7205 7675
rect 7240 7575 7260 7675
rect 7295 7575 7455 7675
rect 7490 7575 7510 7675
rect 7545 7575 7705 7675
rect 7740 7575 7760 7675
rect 7795 7575 7955 7675
rect 7990 7575 8000 7675
rect 0 7570 8000 7575
rect 70 7545 180 7570
rect 70 7510 75 7545
rect 175 7510 180 7545
rect 70 7490 180 7510
rect 70 7455 75 7490
rect 175 7455 180 7490
rect 70 7430 180 7455
rect 320 7545 430 7570
rect 320 7510 325 7545
rect 425 7510 430 7545
rect 320 7490 430 7510
rect 320 7455 325 7490
rect 425 7455 430 7490
rect 320 7430 430 7455
rect 570 7545 680 7570
rect 570 7510 575 7545
rect 675 7510 680 7545
rect 570 7490 680 7510
rect 570 7455 575 7490
rect 675 7455 680 7490
rect 570 7430 680 7455
rect 820 7545 930 7570
rect 820 7510 825 7545
rect 925 7510 930 7545
rect 820 7490 930 7510
rect 820 7455 825 7490
rect 925 7455 930 7490
rect 820 7430 930 7455
rect 1070 7545 1180 7570
rect 1070 7510 1075 7545
rect 1175 7510 1180 7545
rect 1070 7490 1180 7510
rect 1070 7455 1075 7490
rect 1175 7455 1180 7490
rect 1070 7430 1180 7455
rect 1320 7545 1430 7570
rect 1320 7510 1325 7545
rect 1425 7510 1430 7545
rect 1320 7490 1430 7510
rect 1320 7455 1325 7490
rect 1425 7455 1430 7490
rect 1320 7430 1430 7455
rect 1570 7545 1680 7570
rect 1570 7510 1575 7545
rect 1675 7510 1680 7545
rect 1570 7490 1680 7510
rect 1570 7455 1575 7490
rect 1675 7455 1680 7490
rect 1570 7430 1680 7455
rect 1820 7545 1930 7570
rect 1820 7510 1825 7545
rect 1925 7510 1930 7545
rect 1820 7490 1930 7510
rect 1820 7455 1825 7490
rect 1925 7455 1930 7490
rect 1820 7430 1930 7455
rect 2070 7545 2180 7570
rect 2070 7510 2075 7545
rect 2175 7510 2180 7545
rect 2070 7490 2180 7510
rect 2070 7455 2075 7490
rect 2175 7455 2180 7490
rect 2070 7430 2180 7455
rect 2320 7545 2430 7570
rect 2320 7510 2325 7545
rect 2425 7510 2430 7545
rect 2320 7490 2430 7510
rect 2320 7455 2325 7490
rect 2425 7455 2430 7490
rect 2320 7430 2430 7455
rect 2570 7545 2680 7570
rect 2570 7510 2575 7545
rect 2675 7510 2680 7545
rect 2570 7490 2680 7510
rect 2570 7455 2575 7490
rect 2675 7455 2680 7490
rect 2570 7430 2680 7455
rect 2820 7545 2930 7570
rect 2820 7510 2825 7545
rect 2925 7510 2930 7545
rect 2820 7490 2930 7510
rect 2820 7455 2825 7490
rect 2925 7455 2930 7490
rect 2820 7430 2930 7455
rect 3070 7545 3180 7570
rect 3070 7510 3075 7545
rect 3175 7510 3180 7545
rect 3070 7490 3180 7510
rect 3070 7455 3075 7490
rect 3175 7455 3180 7490
rect 3070 7430 3180 7455
rect 3320 7545 3430 7570
rect 3320 7510 3325 7545
rect 3425 7510 3430 7545
rect 3320 7490 3430 7510
rect 3320 7455 3325 7490
rect 3425 7455 3430 7490
rect 3320 7430 3430 7455
rect 3570 7545 3680 7570
rect 3570 7510 3575 7545
rect 3675 7510 3680 7545
rect 3570 7490 3680 7510
rect 3570 7455 3575 7490
rect 3675 7455 3680 7490
rect 3570 7430 3680 7455
rect 3820 7545 3930 7570
rect 3820 7510 3825 7545
rect 3925 7510 3930 7545
rect 3820 7490 3930 7510
rect 3820 7455 3825 7490
rect 3925 7455 3930 7490
rect 3820 7430 3930 7455
rect 4070 7545 4180 7570
rect 4070 7510 4075 7545
rect 4175 7510 4180 7545
rect 4070 7490 4180 7510
rect 4070 7455 4075 7490
rect 4175 7455 4180 7490
rect 4070 7430 4180 7455
rect 4320 7545 4430 7570
rect 4320 7510 4325 7545
rect 4425 7510 4430 7545
rect 4320 7490 4430 7510
rect 4320 7455 4325 7490
rect 4425 7455 4430 7490
rect 4320 7430 4430 7455
rect 4570 7545 4680 7570
rect 4570 7510 4575 7545
rect 4675 7510 4680 7545
rect 4570 7490 4680 7510
rect 4570 7455 4575 7490
rect 4675 7455 4680 7490
rect 4570 7430 4680 7455
rect 4820 7545 4930 7570
rect 4820 7510 4825 7545
rect 4925 7510 4930 7545
rect 4820 7490 4930 7510
rect 4820 7455 4825 7490
rect 4925 7455 4930 7490
rect 4820 7430 4930 7455
rect 5070 7545 5180 7570
rect 5070 7510 5075 7545
rect 5175 7510 5180 7545
rect 5070 7490 5180 7510
rect 5070 7455 5075 7490
rect 5175 7455 5180 7490
rect 5070 7430 5180 7455
rect 5320 7545 5430 7570
rect 5320 7510 5325 7545
rect 5425 7510 5430 7545
rect 5320 7490 5430 7510
rect 5320 7455 5325 7490
rect 5425 7455 5430 7490
rect 5320 7430 5430 7455
rect 5570 7545 5680 7570
rect 5570 7510 5575 7545
rect 5675 7510 5680 7545
rect 5570 7490 5680 7510
rect 5570 7455 5575 7490
rect 5675 7455 5680 7490
rect 5570 7430 5680 7455
rect 5820 7545 5930 7570
rect 5820 7510 5825 7545
rect 5925 7510 5930 7545
rect 5820 7490 5930 7510
rect 5820 7455 5825 7490
rect 5925 7455 5930 7490
rect 5820 7430 5930 7455
rect 6070 7545 6180 7570
rect 6070 7510 6075 7545
rect 6175 7510 6180 7545
rect 6070 7490 6180 7510
rect 6070 7455 6075 7490
rect 6175 7455 6180 7490
rect 6070 7430 6180 7455
rect 6320 7545 6430 7570
rect 6320 7510 6325 7545
rect 6425 7510 6430 7545
rect 6320 7490 6430 7510
rect 6320 7455 6325 7490
rect 6425 7455 6430 7490
rect 6320 7430 6430 7455
rect 6570 7545 6680 7570
rect 6570 7510 6575 7545
rect 6675 7510 6680 7545
rect 6570 7490 6680 7510
rect 6570 7455 6575 7490
rect 6675 7455 6680 7490
rect 6570 7430 6680 7455
rect 6820 7545 6930 7570
rect 6820 7510 6825 7545
rect 6925 7510 6930 7545
rect 6820 7490 6930 7510
rect 6820 7455 6825 7490
rect 6925 7455 6930 7490
rect 6820 7430 6930 7455
rect 7070 7545 7180 7570
rect 7070 7510 7075 7545
rect 7175 7510 7180 7545
rect 7070 7490 7180 7510
rect 7070 7455 7075 7490
rect 7175 7455 7180 7490
rect 7070 7430 7180 7455
rect 7320 7545 7430 7570
rect 7320 7510 7325 7545
rect 7425 7510 7430 7545
rect 7320 7490 7430 7510
rect 7320 7455 7325 7490
rect 7425 7455 7430 7490
rect 7320 7430 7430 7455
rect 7570 7545 7680 7570
rect 7570 7510 7575 7545
rect 7675 7510 7680 7545
rect 7570 7490 7680 7510
rect 7570 7455 7575 7490
rect 7675 7455 7680 7490
rect 7570 7430 7680 7455
rect 7820 7545 7930 7570
rect 7820 7510 7825 7545
rect 7925 7510 7930 7545
rect 7820 7490 7930 7510
rect 7820 7455 7825 7490
rect 7925 7455 7930 7490
rect 7820 7430 7930 7455
rect 0 7425 8000 7430
rect 0 7325 10 7425
rect 45 7325 205 7425
rect 240 7325 260 7425
rect 295 7325 455 7425
rect 490 7325 510 7425
rect 545 7325 705 7425
rect 740 7325 760 7425
rect 795 7325 955 7425
rect 990 7325 1010 7425
rect 1045 7325 1205 7425
rect 1240 7325 1260 7425
rect 1295 7325 1455 7425
rect 1490 7325 1510 7425
rect 1545 7325 1705 7425
rect 1740 7325 1760 7425
rect 1795 7325 1955 7425
rect 1990 7325 2010 7425
rect 2045 7325 2205 7425
rect 2240 7325 2260 7425
rect 2295 7325 2455 7425
rect 2490 7325 2510 7425
rect 2545 7325 2705 7425
rect 2740 7325 2760 7425
rect 2795 7325 2955 7425
rect 2990 7325 3010 7425
rect 3045 7325 3205 7425
rect 3240 7325 3260 7425
rect 3295 7325 3455 7425
rect 3490 7325 3510 7425
rect 3545 7325 3705 7425
rect 3740 7325 3760 7425
rect 3795 7325 3955 7425
rect 3990 7325 4010 7425
rect 4045 7325 4205 7425
rect 4240 7325 4260 7425
rect 4295 7325 4455 7425
rect 4490 7325 4510 7425
rect 4545 7325 4705 7425
rect 4740 7325 4760 7425
rect 4795 7325 4955 7425
rect 4990 7325 5010 7425
rect 5045 7325 5205 7425
rect 5240 7325 5260 7425
rect 5295 7325 5455 7425
rect 5490 7325 5510 7425
rect 5545 7325 5705 7425
rect 5740 7325 5760 7425
rect 5795 7325 5955 7425
rect 5990 7325 6010 7425
rect 6045 7325 6205 7425
rect 6240 7325 6260 7425
rect 6295 7325 6455 7425
rect 6490 7325 6510 7425
rect 6545 7325 6705 7425
rect 6740 7325 6760 7425
rect 6795 7325 6955 7425
rect 6990 7325 7010 7425
rect 7045 7325 7205 7425
rect 7240 7325 7260 7425
rect 7295 7325 7455 7425
rect 7490 7325 7510 7425
rect 7545 7325 7705 7425
rect 7740 7325 7760 7425
rect 7795 7325 7955 7425
rect 7990 7325 8000 7425
rect 0 7320 8000 7325
rect 70 7295 180 7320
rect 70 7260 75 7295
rect 175 7260 180 7295
rect 70 7240 180 7260
rect 70 7205 75 7240
rect 175 7205 180 7240
rect 70 7180 180 7205
rect 320 7295 430 7320
rect 320 7260 325 7295
rect 425 7260 430 7295
rect 320 7240 430 7260
rect 320 7205 325 7240
rect 425 7205 430 7240
rect 320 7180 430 7205
rect 570 7295 680 7320
rect 570 7260 575 7295
rect 675 7260 680 7295
rect 570 7240 680 7260
rect 570 7205 575 7240
rect 675 7205 680 7240
rect 570 7180 680 7205
rect 820 7295 930 7320
rect 820 7260 825 7295
rect 925 7260 930 7295
rect 820 7240 930 7260
rect 820 7205 825 7240
rect 925 7205 930 7240
rect 820 7180 930 7205
rect 1070 7295 1180 7320
rect 1070 7260 1075 7295
rect 1175 7260 1180 7295
rect 1070 7240 1180 7260
rect 1070 7205 1075 7240
rect 1175 7205 1180 7240
rect 1070 7180 1180 7205
rect 1320 7295 1430 7320
rect 1320 7260 1325 7295
rect 1425 7260 1430 7295
rect 1320 7240 1430 7260
rect 1320 7205 1325 7240
rect 1425 7205 1430 7240
rect 1320 7180 1430 7205
rect 1570 7295 1680 7320
rect 1570 7260 1575 7295
rect 1675 7260 1680 7295
rect 1570 7240 1680 7260
rect 1570 7205 1575 7240
rect 1675 7205 1680 7240
rect 1570 7180 1680 7205
rect 1820 7295 1930 7320
rect 1820 7260 1825 7295
rect 1925 7260 1930 7295
rect 1820 7240 1930 7260
rect 1820 7205 1825 7240
rect 1925 7205 1930 7240
rect 1820 7180 1930 7205
rect 2070 7295 2180 7320
rect 2070 7260 2075 7295
rect 2175 7260 2180 7295
rect 2070 7240 2180 7260
rect 2070 7205 2075 7240
rect 2175 7205 2180 7240
rect 2070 7180 2180 7205
rect 2320 7295 2430 7320
rect 2320 7260 2325 7295
rect 2425 7260 2430 7295
rect 2320 7240 2430 7260
rect 2320 7205 2325 7240
rect 2425 7205 2430 7240
rect 2320 7180 2430 7205
rect 2570 7295 2680 7320
rect 2570 7260 2575 7295
rect 2675 7260 2680 7295
rect 2570 7240 2680 7260
rect 2570 7205 2575 7240
rect 2675 7205 2680 7240
rect 2570 7180 2680 7205
rect 2820 7295 2930 7320
rect 2820 7260 2825 7295
rect 2925 7260 2930 7295
rect 2820 7240 2930 7260
rect 2820 7205 2825 7240
rect 2925 7205 2930 7240
rect 2820 7180 2930 7205
rect 3070 7295 3180 7320
rect 3070 7260 3075 7295
rect 3175 7260 3180 7295
rect 3070 7240 3180 7260
rect 3070 7205 3075 7240
rect 3175 7205 3180 7240
rect 3070 7180 3180 7205
rect 3320 7295 3430 7320
rect 3320 7260 3325 7295
rect 3425 7260 3430 7295
rect 3320 7240 3430 7260
rect 3320 7205 3325 7240
rect 3425 7205 3430 7240
rect 3320 7180 3430 7205
rect 3570 7295 3680 7320
rect 3570 7260 3575 7295
rect 3675 7260 3680 7295
rect 3570 7240 3680 7260
rect 3570 7205 3575 7240
rect 3675 7205 3680 7240
rect 3570 7180 3680 7205
rect 3820 7295 3930 7320
rect 3820 7260 3825 7295
rect 3925 7260 3930 7295
rect 3820 7240 3930 7260
rect 3820 7205 3825 7240
rect 3925 7205 3930 7240
rect 3820 7180 3930 7205
rect 4070 7295 4180 7320
rect 4070 7260 4075 7295
rect 4175 7260 4180 7295
rect 4070 7240 4180 7260
rect 4070 7205 4075 7240
rect 4175 7205 4180 7240
rect 4070 7180 4180 7205
rect 4320 7295 4430 7320
rect 4320 7260 4325 7295
rect 4425 7260 4430 7295
rect 4320 7240 4430 7260
rect 4320 7205 4325 7240
rect 4425 7205 4430 7240
rect 4320 7180 4430 7205
rect 4570 7295 4680 7320
rect 4570 7260 4575 7295
rect 4675 7260 4680 7295
rect 4570 7240 4680 7260
rect 4570 7205 4575 7240
rect 4675 7205 4680 7240
rect 4570 7180 4680 7205
rect 4820 7295 4930 7320
rect 4820 7260 4825 7295
rect 4925 7260 4930 7295
rect 4820 7240 4930 7260
rect 4820 7205 4825 7240
rect 4925 7205 4930 7240
rect 4820 7180 4930 7205
rect 5070 7295 5180 7320
rect 5070 7260 5075 7295
rect 5175 7260 5180 7295
rect 5070 7240 5180 7260
rect 5070 7205 5075 7240
rect 5175 7205 5180 7240
rect 5070 7180 5180 7205
rect 5320 7295 5430 7320
rect 5320 7260 5325 7295
rect 5425 7260 5430 7295
rect 5320 7240 5430 7260
rect 5320 7205 5325 7240
rect 5425 7205 5430 7240
rect 5320 7180 5430 7205
rect 5570 7295 5680 7320
rect 5570 7260 5575 7295
rect 5675 7260 5680 7295
rect 5570 7240 5680 7260
rect 5570 7205 5575 7240
rect 5675 7205 5680 7240
rect 5570 7180 5680 7205
rect 5820 7295 5930 7320
rect 5820 7260 5825 7295
rect 5925 7260 5930 7295
rect 5820 7240 5930 7260
rect 5820 7205 5825 7240
rect 5925 7205 5930 7240
rect 5820 7180 5930 7205
rect 6070 7295 6180 7320
rect 6070 7260 6075 7295
rect 6175 7260 6180 7295
rect 6070 7240 6180 7260
rect 6070 7205 6075 7240
rect 6175 7205 6180 7240
rect 6070 7180 6180 7205
rect 6320 7295 6430 7320
rect 6320 7260 6325 7295
rect 6425 7260 6430 7295
rect 6320 7240 6430 7260
rect 6320 7205 6325 7240
rect 6425 7205 6430 7240
rect 6320 7180 6430 7205
rect 6570 7295 6680 7320
rect 6570 7260 6575 7295
rect 6675 7260 6680 7295
rect 6570 7240 6680 7260
rect 6570 7205 6575 7240
rect 6675 7205 6680 7240
rect 6570 7180 6680 7205
rect 6820 7295 6930 7320
rect 6820 7260 6825 7295
rect 6925 7260 6930 7295
rect 6820 7240 6930 7260
rect 6820 7205 6825 7240
rect 6925 7205 6930 7240
rect 6820 7180 6930 7205
rect 7070 7295 7180 7320
rect 7070 7260 7075 7295
rect 7175 7260 7180 7295
rect 7070 7240 7180 7260
rect 7070 7205 7075 7240
rect 7175 7205 7180 7240
rect 7070 7180 7180 7205
rect 7320 7295 7430 7320
rect 7320 7260 7325 7295
rect 7425 7260 7430 7295
rect 7320 7240 7430 7260
rect 7320 7205 7325 7240
rect 7425 7205 7430 7240
rect 7320 7180 7430 7205
rect 7570 7295 7680 7320
rect 7570 7260 7575 7295
rect 7675 7260 7680 7295
rect 7570 7240 7680 7260
rect 7570 7205 7575 7240
rect 7675 7205 7680 7240
rect 7570 7180 7680 7205
rect 7820 7295 7930 7320
rect 7820 7260 7825 7295
rect 7925 7260 7930 7295
rect 7820 7240 7930 7260
rect 7820 7205 7825 7240
rect 7925 7205 7930 7240
rect 7820 7180 7930 7205
rect 0 7175 8000 7180
rect 0 7075 10 7175
rect 45 7075 205 7175
rect 240 7075 260 7175
rect 295 7075 455 7175
rect 490 7075 510 7175
rect 545 7075 705 7175
rect 740 7075 760 7175
rect 795 7075 955 7175
rect 990 7075 1010 7175
rect 1045 7075 1205 7175
rect 1240 7075 1260 7175
rect 1295 7075 1455 7175
rect 1490 7075 1510 7175
rect 1545 7075 1705 7175
rect 1740 7075 1760 7175
rect 1795 7075 1955 7175
rect 1990 7075 2010 7175
rect 2045 7075 2205 7175
rect 2240 7075 2260 7175
rect 2295 7075 2455 7175
rect 2490 7075 2510 7175
rect 2545 7075 2705 7175
rect 2740 7075 2760 7175
rect 2795 7075 2955 7175
rect 2990 7075 3010 7175
rect 3045 7075 3205 7175
rect 3240 7075 3260 7175
rect 3295 7075 3455 7175
rect 3490 7075 3510 7175
rect 3545 7075 3705 7175
rect 3740 7075 3760 7175
rect 3795 7075 3955 7175
rect 3990 7075 4010 7175
rect 4045 7075 4205 7175
rect 4240 7075 4260 7175
rect 4295 7075 4455 7175
rect 4490 7075 4510 7175
rect 4545 7075 4705 7175
rect 4740 7075 4760 7175
rect 4795 7075 4955 7175
rect 4990 7075 5010 7175
rect 5045 7075 5205 7175
rect 5240 7075 5260 7175
rect 5295 7075 5455 7175
rect 5490 7075 5510 7175
rect 5545 7075 5705 7175
rect 5740 7075 5760 7175
rect 5795 7075 5955 7175
rect 5990 7075 6010 7175
rect 6045 7075 6205 7175
rect 6240 7075 6260 7175
rect 6295 7075 6455 7175
rect 6490 7075 6510 7175
rect 6545 7075 6705 7175
rect 6740 7075 6760 7175
rect 6795 7075 6955 7175
rect 6990 7075 7010 7175
rect 7045 7075 7205 7175
rect 7240 7075 7260 7175
rect 7295 7075 7455 7175
rect 7490 7075 7510 7175
rect 7545 7075 7705 7175
rect 7740 7075 7760 7175
rect 7795 7075 7955 7175
rect 7990 7075 8000 7175
rect 0 7070 8000 7075
rect 70 7045 180 7070
rect 70 7010 75 7045
rect 175 7010 180 7045
rect 70 6990 180 7010
rect 70 6955 75 6990
rect 175 6955 180 6990
rect 70 6930 180 6955
rect 320 7045 430 7070
rect 320 7010 325 7045
rect 425 7010 430 7045
rect 320 6990 430 7010
rect 320 6955 325 6990
rect 425 6955 430 6990
rect 320 6930 430 6955
rect 570 7045 680 7070
rect 570 7010 575 7045
rect 675 7010 680 7045
rect 570 6990 680 7010
rect 570 6955 575 6990
rect 675 6955 680 6990
rect 570 6930 680 6955
rect 820 7045 930 7070
rect 820 7010 825 7045
rect 925 7010 930 7045
rect 820 6990 930 7010
rect 820 6955 825 6990
rect 925 6955 930 6990
rect 820 6930 930 6955
rect 1070 7045 1180 7070
rect 1070 7010 1075 7045
rect 1175 7010 1180 7045
rect 1070 6990 1180 7010
rect 1070 6955 1075 6990
rect 1175 6955 1180 6990
rect 1070 6930 1180 6955
rect 1320 7045 1430 7070
rect 1320 7010 1325 7045
rect 1425 7010 1430 7045
rect 1320 6990 1430 7010
rect 1320 6955 1325 6990
rect 1425 6955 1430 6990
rect 1320 6930 1430 6955
rect 1570 7045 1680 7070
rect 1570 7010 1575 7045
rect 1675 7010 1680 7045
rect 1570 6990 1680 7010
rect 1570 6955 1575 6990
rect 1675 6955 1680 6990
rect 1570 6930 1680 6955
rect 1820 7045 1930 7070
rect 1820 7010 1825 7045
rect 1925 7010 1930 7045
rect 1820 6990 1930 7010
rect 1820 6955 1825 6990
rect 1925 6955 1930 6990
rect 1820 6930 1930 6955
rect 2070 7045 2180 7070
rect 2070 7010 2075 7045
rect 2175 7010 2180 7045
rect 2070 6990 2180 7010
rect 2070 6955 2075 6990
rect 2175 6955 2180 6990
rect 2070 6930 2180 6955
rect 2320 7045 2430 7070
rect 2320 7010 2325 7045
rect 2425 7010 2430 7045
rect 2320 6990 2430 7010
rect 2320 6955 2325 6990
rect 2425 6955 2430 6990
rect 2320 6930 2430 6955
rect 2570 7045 2680 7070
rect 2570 7010 2575 7045
rect 2675 7010 2680 7045
rect 2570 6990 2680 7010
rect 2570 6955 2575 6990
rect 2675 6955 2680 6990
rect 2570 6930 2680 6955
rect 2820 7045 2930 7070
rect 2820 7010 2825 7045
rect 2925 7010 2930 7045
rect 2820 6990 2930 7010
rect 2820 6955 2825 6990
rect 2925 6955 2930 6990
rect 2820 6930 2930 6955
rect 3070 7045 3180 7070
rect 3070 7010 3075 7045
rect 3175 7010 3180 7045
rect 3070 6990 3180 7010
rect 3070 6955 3075 6990
rect 3175 6955 3180 6990
rect 3070 6930 3180 6955
rect 3320 7045 3430 7070
rect 3320 7010 3325 7045
rect 3425 7010 3430 7045
rect 3320 6990 3430 7010
rect 3320 6955 3325 6990
rect 3425 6955 3430 6990
rect 3320 6930 3430 6955
rect 3570 7045 3680 7070
rect 3570 7010 3575 7045
rect 3675 7010 3680 7045
rect 3570 6990 3680 7010
rect 3570 6955 3575 6990
rect 3675 6955 3680 6990
rect 3570 6930 3680 6955
rect 3820 7045 3930 7070
rect 3820 7010 3825 7045
rect 3925 7010 3930 7045
rect 3820 6990 3930 7010
rect 3820 6955 3825 6990
rect 3925 6955 3930 6990
rect 3820 6930 3930 6955
rect 4070 7045 4180 7070
rect 4070 7010 4075 7045
rect 4175 7010 4180 7045
rect 4070 6990 4180 7010
rect 4070 6955 4075 6990
rect 4175 6955 4180 6990
rect 4070 6930 4180 6955
rect 4320 7045 4430 7070
rect 4320 7010 4325 7045
rect 4425 7010 4430 7045
rect 4320 6990 4430 7010
rect 4320 6955 4325 6990
rect 4425 6955 4430 6990
rect 4320 6930 4430 6955
rect 4570 7045 4680 7070
rect 4570 7010 4575 7045
rect 4675 7010 4680 7045
rect 4570 6990 4680 7010
rect 4570 6955 4575 6990
rect 4675 6955 4680 6990
rect 4570 6930 4680 6955
rect 4820 7045 4930 7070
rect 4820 7010 4825 7045
rect 4925 7010 4930 7045
rect 4820 6990 4930 7010
rect 4820 6955 4825 6990
rect 4925 6955 4930 6990
rect 4820 6930 4930 6955
rect 5070 7045 5180 7070
rect 5070 7010 5075 7045
rect 5175 7010 5180 7045
rect 5070 6990 5180 7010
rect 5070 6955 5075 6990
rect 5175 6955 5180 6990
rect 5070 6930 5180 6955
rect 5320 7045 5430 7070
rect 5320 7010 5325 7045
rect 5425 7010 5430 7045
rect 5320 6990 5430 7010
rect 5320 6955 5325 6990
rect 5425 6955 5430 6990
rect 5320 6930 5430 6955
rect 5570 7045 5680 7070
rect 5570 7010 5575 7045
rect 5675 7010 5680 7045
rect 5570 6990 5680 7010
rect 5570 6955 5575 6990
rect 5675 6955 5680 6990
rect 5570 6930 5680 6955
rect 5820 7045 5930 7070
rect 5820 7010 5825 7045
rect 5925 7010 5930 7045
rect 5820 6990 5930 7010
rect 5820 6955 5825 6990
rect 5925 6955 5930 6990
rect 5820 6930 5930 6955
rect 6070 7045 6180 7070
rect 6070 7010 6075 7045
rect 6175 7010 6180 7045
rect 6070 6990 6180 7010
rect 6070 6955 6075 6990
rect 6175 6955 6180 6990
rect 6070 6930 6180 6955
rect 6320 7045 6430 7070
rect 6320 7010 6325 7045
rect 6425 7010 6430 7045
rect 6320 6990 6430 7010
rect 6320 6955 6325 6990
rect 6425 6955 6430 6990
rect 6320 6930 6430 6955
rect 6570 7045 6680 7070
rect 6570 7010 6575 7045
rect 6675 7010 6680 7045
rect 6570 6990 6680 7010
rect 6570 6955 6575 6990
rect 6675 6955 6680 6990
rect 6570 6930 6680 6955
rect 6820 7045 6930 7070
rect 6820 7010 6825 7045
rect 6925 7010 6930 7045
rect 6820 6990 6930 7010
rect 6820 6955 6825 6990
rect 6925 6955 6930 6990
rect 6820 6930 6930 6955
rect 7070 7045 7180 7070
rect 7070 7010 7075 7045
rect 7175 7010 7180 7045
rect 7070 6990 7180 7010
rect 7070 6955 7075 6990
rect 7175 6955 7180 6990
rect 7070 6930 7180 6955
rect 7320 7045 7430 7070
rect 7320 7010 7325 7045
rect 7425 7010 7430 7045
rect 7320 6990 7430 7010
rect 7320 6955 7325 6990
rect 7425 6955 7430 6990
rect 7320 6930 7430 6955
rect 7570 7045 7680 7070
rect 7570 7010 7575 7045
rect 7675 7010 7680 7045
rect 7570 6990 7680 7010
rect 7570 6955 7575 6990
rect 7675 6955 7680 6990
rect 7570 6930 7680 6955
rect 7820 7045 7930 7070
rect 7820 7010 7825 7045
rect 7925 7010 7930 7045
rect 7820 6990 7930 7010
rect 7820 6955 7825 6990
rect 7925 6955 7930 6990
rect 7820 6930 7930 6955
rect 0 6925 8000 6930
rect 0 6825 10 6925
rect 45 6825 205 6925
rect 240 6825 260 6925
rect 295 6825 455 6925
rect 490 6825 510 6925
rect 545 6825 705 6925
rect 740 6825 760 6925
rect 795 6825 955 6925
rect 990 6825 1010 6925
rect 1045 6825 1205 6925
rect 1240 6825 1260 6925
rect 1295 6825 1455 6925
rect 1490 6825 1510 6925
rect 1545 6825 1705 6925
rect 1740 6825 1760 6925
rect 1795 6825 1955 6925
rect 1990 6825 2010 6925
rect 2045 6825 2205 6925
rect 2240 6825 2260 6925
rect 2295 6825 2455 6925
rect 2490 6825 2510 6925
rect 2545 6825 2705 6925
rect 2740 6825 2760 6925
rect 2795 6825 2955 6925
rect 2990 6825 3010 6925
rect 3045 6825 3205 6925
rect 3240 6825 3260 6925
rect 3295 6825 3455 6925
rect 3490 6825 3510 6925
rect 3545 6825 3705 6925
rect 3740 6825 3760 6925
rect 3795 6825 3955 6925
rect 3990 6825 4010 6925
rect 4045 6825 4205 6925
rect 4240 6825 4260 6925
rect 4295 6825 4455 6925
rect 4490 6825 4510 6925
rect 4545 6825 4705 6925
rect 4740 6825 4760 6925
rect 4795 6825 4955 6925
rect 4990 6825 5010 6925
rect 5045 6825 5205 6925
rect 5240 6825 5260 6925
rect 5295 6825 5455 6925
rect 5490 6825 5510 6925
rect 5545 6825 5705 6925
rect 5740 6825 5760 6925
rect 5795 6825 5955 6925
rect 5990 6825 6010 6925
rect 6045 6825 6205 6925
rect 6240 6825 6260 6925
rect 6295 6825 6455 6925
rect 6490 6825 6510 6925
rect 6545 6825 6705 6925
rect 6740 6825 6760 6925
rect 6795 6825 6955 6925
rect 6990 6825 7010 6925
rect 7045 6825 7205 6925
rect 7240 6825 7260 6925
rect 7295 6825 7455 6925
rect 7490 6825 7510 6925
rect 7545 6825 7705 6925
rect 7740 6825 7760 6925
rect 7795 6825 7955 6925
rect 7990 6825 8000 6925
rect 0 6820 8000 6825
rect 70 6795 180 6820
rect 70 6760 75 6795
rect 175 6760 180 6795
rect 70 6740 180 6760
rect 70 6705 75 6740
rect 175 6705 180 6740
rect 70 6680 180 6705
rect 320 6795 430 6820
rect 320 6760 325 6795
rect 425 6760 430 6795
rect 320 6740 430 6760
rect 320 6705 325 6740
rect 425 6705 430 6740
rect 320 6680 430 6705
rect 570 6795 680 6820
rect 570 6760 575 6795
rect 675 6760 680 6795
rect 570 6740 680 6760
rect 570 6705 575 6740
rect 675 6705 680 6740
rect 570 6680 680 6705
rect 820 6795 930 6820
rect 820 6760 825 6795
rect 925 6760 930 6795
rect 820 6740 930 6760
rect 820 6705 825 6740
rect 925 6705 930 6740
rect 820 6680 930 6705
rect 1070 6795 1180 6820
rect 1070 6760 1075 6795
rect 1175 6760 1180 6795
rect 1070 6740 1180 6760
rect 1070 6705 1075 6740
rect 1175 6705 1180 6740
rect 1070 6680 1180 6705
rect 1320 6795 1430 6820
rect 1320 6760 1325 6795
rect 1425 6760 1430 6795
rect 1320 6740 1430 6760
rect 1320 6705 1325 6740
rect 1425 6705 1430 6740
rect 1320 6680 1430 6705
rect 1570 6795 1680 6820
rect 1570 6760 1575 6795
rect 1675 6760 1680 6795
rect 1570 6740 1680 6760
rect 1570 6705 1575 6740
rect 1675 6705 1680 6740
rect 1570 6680 1680 6705
rect 1820 6795 1930 6820
rect 1820 6760 1825 6795
rect 1925 6760 1930 6795
rect 1820 6740 1930 6760
rect 1820 6705 1825 6740
rect 1925 6705 1930 6740
rect 1820 6680 1930 6705
rect 2070 6795 2180 6820
rect 2070 6760 2075 6795
rect 2175 6760 2180 6795
rect 2070 6740 2180 6760
rect 2070 6705 2075 6740
rect 2175 6705 2180 6740
rect 2070 6680 2180 6705
rect 2320 6795 2430 6820
rect 2320 6760 2325 6795
rect 2425 6760 2430 6795
rect 2320 6740 2430 6760
rect 2320 6705 2325 6740
rect 2425 6705 2430 6740
rect 2320 6680 2430 6705
rect 2570 6795 2680 6820
rect 2570 6760 2575 6795
rect 2675 6760 2680 6795
rect 2570 6740 2680 6760
rect 2570 6705 2575 6740
rect 2675 6705 2680 6740
rect 2570 6680 2680 6705
rect 2820 6795 2930 6820
rect 2820 6760 2825 6795
rect 2925 6760 2930 6795
rect 2820 6740 2930 6760
rect 2820 6705 2825 6740
rect 2925 6705 2930 6740
rect 2820 6680 2930 6705
rect 3070 6795 3180 6820
rect 3070 6760 3075 6795
rect 3175 6760 3180 6795
rect 3070 6740 3180 6760
rect 3070 6705 3075 6740
rect 3175 6705 3180 6740
rect 3070 6680 3180 6705
rect 3320 6795 3430 6820
rect 3320 6760 3325 6795
rect 3425 6760 3430 6795
rect 3320 6740 3430 6760
rect 3320 6705 3325 6740
rect 3425 6705 3430 6740
rect 3320 6680 3430 6705
rect 3570 6795 3680 6820
rect 3570 6760 3575 6795
rect 3675 6760 3680 6795
rect 3570 6740 3680 6760
rect 3570 6705 3575 6740
rect 3675 6705 3680 6740
rect 3570 6680 3680 6705
rect 3820 6795 3930 6820
rect 3820 6760 3825 6795
rect 3925 6760 3930 6795
rect 3820 6740 3930 6760
rect 3820 6705 3825 6740
rect 3925 6705 3930 6740
rect 3820 6680 3930 6705
rect 4070 6795 4180 6820
rect 4070 6760 4075 6795
rect 4175 6760 4180 6795
rect 4070 6740 4180 6760
rect 4070 6705 4075 6740
rect 4175 6705 4180 6740
rect 4070 6680 4180 6705
rect 4320 6795 4430 6820
rect 4320 6760 4325 6795
rect 4425 6760 4430 6795
rect 4320 6740 4430 6760
rect 4320 6705 4325 6740
rect 4425 6705 4430 6740
rect 4320 6680 4430 6705
rect 4570 6795 4680 6820
rect 4570 6760 4575 6795
rect 4675 6760 4680 6795
rect 4570 6740 4680 6760
rect 4570 6705 4575 6740
rect 4675 6705 4680 6740
rect 4570 6680 4680 6705
rect 4820 6795 4930 6820
rect 4820 6760 4825 6795
rect 4925 6760 4930 6795
rect 4820 6740 4930 6760
rect 4820 6705 4825 6740
rect 4925 6705 4930 6740
rect 4820 6680 4930 6705
rect 5070 6795 5180 6820
rect 5070 6760 5075 6795
rect 5175 6760 5180 6795
rect 5070 6740 5180 6760
rect 5070 6705 5075 6740
rect 5175 6705 5180 6740
rect 5070 6680 5180 6705
rect 5320 6795 5430 6820
rect 5320 6760 5325 6795
rect 5425 6760 5430 6795
rect 5320 6740 5430 6760
rect 5320 6705 5325 6740
rect 5425 6705 5430 6740
rect 5320 6680 5430 6705
rect 5570 6795 5680 6820
rect 5570 6760 5575 6795
rect 5675 6760 5680 6795
rect 5570 6740 5680 6760
rect 5570 6705 5575 6740
rect 5675 6705 5680 6740
rect 5570 6680 5680 6705
rect 5820 6795 5930 6820
rect 5820 6760 5825 6795
rect 5925 6760 5930 6795
rect 5820 6740 5930 6760
rect 5820 6705 5825 6740
rect 5925 6705 5930 6740
rect 5820 6680 5930 6705
rect 6070 6795 6180 6820
rect 6070 6760 6075 6795
rect 6175 6760 6180 6795
rect 6070 6740 6180 6760
rect 6070 6705 6075 6740
rect 6175 6705 6180 6740
rect 6070 6680 6180 6705
rect 6320 6795 6430 6820
rect 6320 6760 6325 6795
rect 6425 6760 6430 6795
rect 6320 6740 6430 6760
rect 6320 6705 6325 6740
rect 6425 6705 6430 6740
rect 6320 6680 6430 6705
rect 6570 6795 6680 6820
rect 6570 6760 6575 6795
rect 6675 6760 6680 6795
rect 6570 6740 6680 6760
rect 6570 6705 6575 6740
rect 6675 6705 6680 6740
rect 6570 6680 6680 6705
rect 6820 6795 6930 6820
rect 6820 6760 6825 6795
rect 6925 6760 6930 6795
rect 6820 6740 6930 6760
rect 6820 6705 6825 6740
rect 6925 6705 6930 6740
rect 6820 6680 6930 6705
rect 7070 6795 7180 6820
rect 7070 6760 7075 6795
rect 7175 6760 7180 6795
rect 7070 6740 7180 6760
rect 7070 6705 7075 6740
rect 7175 6705 7180 6740
rect 7070 6680 7180 6705
rect 7320 6795 7430 6820
rect 7320 6760 7325 6795
rect 7425 6760 7430 6795
rect 7320 6740 7430 6760
rect 7320 6705 7325 6740
rect 7425 6705 7430 6740
rect 7320 6680 7430 6705
rect 7570 6795 7680 6820
rect 7570 6760 7575 6795
rect 7675 6760 7680 6795
rect 7570 6740 7680 6760
rect 7570 6705 7575 6740
rect 7675 6705 7680 6740
rect 7570 6680 7680 6705
rect 7820 6795 7930 6820
rect 7820 6760 7825 6795
rect 7925 6760 7930 6795
rect 7820 6740 7930 6760
rect 7820 6705 7825 6740
rect 7925 6705 7930 6740
rect 7820 6680 7930 6705
rect 0 6675 8000 6680
rect 0 6575 10 6675
rect 45 6575 205 6675
rect 240 6575 260 6675
rect 295 6575 455 6675
rect 490 6575 510 6675
rect 545 6575 705 6675
rect 740 6575 760 6675
rect 795 6575 955 6675
rect 990 6575 1010 6675
rect 1045 6575 1205 6675
rect 1240 6575 1260 6675
rect 1295 6575 1455 6675
rect 1490 6575 1510 6675
rect 1545 6575 1705 6675
rect 1740 6575 1760 6675
rect 1795 6575 1955 6675
rect 1990 6575 2010 6675
rect 2045 6575 2205 6675
rect 2240 6575 2260 6675
rect 2295 6575 2455 6675
rect 2490 6575 2510 6675
rect 2545 6575 2705 6675
rect 2740 6575 2760 6675
rect 2795 6575 2955 6675
rect 2990 6575 3010 6675
rect 3045 6575 3205 6675
rect 3240 6575 3260 6675
rect 3295 6575 3455 6675
rect 3490 6575 3510 6675
rect 3545 6575 3705 6675
rect 3740 6575 3760 6675
rect 3795 6575 3955 6675
rect 3990 6575 4010 6675
rect 4045 6575 4205 6675
rect 4240 6575 4260 6675
rect 4295 6575 4455 6675
rect 4490 6575 4510 6675
rect 4545 6575 4705 6675
rect 4740 6575 4760 6675
rect 4795 6575 4955 6675
rect 4990 6575 5010 6675
rect 5045 6575 5205 6675
rect 5240 6575 5260 6675
rect 5295 6575 5455 6675
rect 5490 6575 5510 6675
rect 5545 6575 5705 6675
rect 5740 6575 5760 6675
rect 5795 6575 5955 6675
rect 5990 6575 6010 6675
rect 6045 6575 6205 6675
rect 6240 6575 6260 6675
rect 6295 6575 6455 6675
rect 6490 6575 6510 6675
rect 6545 6575 6705 6675
rect 6740 6575 6760 6675
rect 6795 6575 6955 6675
rect 6990 6575 7010 6675
rect 7045 6575 7205 6675
rect 7240 6575 7260 6675
rect 7295 6575 7455 6675
rect 7490 6575 7510 6675
rect 7545 6575 7705 6675
rect 7740 6575 7760 6675
rect 7795 6575 7955 6675
rect 7990 6575 8000 6675
rect 0 6570 8000 6575
rect 70 6545 180 6570
rect 70 6510 75 6545
rect 175 6510 180 6545
rect 70 6490 180 6510
rect 70 6455 75 6490
rect 175 6455 180 6490
rect 70 6430 180 6455
rect 320 6545 430 6570
rect 320 6510 325 6545
rect 425 6510 430 6545
rect 320 6490 430 6510
rect 320 6455 325 6490
rect 425 6455 430 6490
rect 320 6430 430 6455
rect 570 6545 680 6570
rect 570 6510 575 6545
rect 675 6510 680 6545
rect 570 6490 680 6510
rect 570 6455 575 6490
rect 675 6455 680 6490
rect 570 6430 680 6455
rect 820 6545 930 6570
rect 820 6510 825 6545
rect 925 6510 930 6545
rect 820 6490 930 6510
rect 820 6455 825 6490
rect 925 6455 930 6490
rect 820 6430 930 6455
rect 1070 6545 1180 6570
rect 1070 6510 1075 6545
rect 1175 6510 1180 6545
rect 1070 6490 1180 6510
rect 1070 6455 1075 6490
rect 1175 6455 1180 6490
rect 1070 6430 1180 6455
rect 1320 6545 1430 6570
rect 1320 6510 1325 6545
rect 1425 6510 1430 6545
rect 1320 6490 1430 6510
rect 1320 6455 1325 6490
rect 1425 6455 1430 6490
rect 1320 6430 1430 6455
rect 1570 6545 1680 6570
rect 1570 6510 1575 6545
rect 1675 6510 1680 6545
rect 1570 6490 1680 6510
rect 1570 6455 1575 6490
rect 1675 6455 1680 6490
rect 1570 6430 1680 6455
rect 1820 6545 1930 6570
rect 1820 6510 1825 6545
rect 1925 6510 1930 6545
rect 1820 6490 1930 6510
rect 1820 6455 1825 6490
rect 1925 6455 1930 6490
rect 1820 6430 1930 6455
rect 2070 6545 2180 6570
rect 2070 6510 2075 6545
rect 2175 6510 2180 6545
rect 2070 6490 2180 6510
rect 2070 6455 2075 6490
rect 2175 6455 2180 6490
rect 2070 6430 2180 6455
rect 2320 6545 2430 6570
rect 2320 6510 2325 6545
rect 2425 6510 2430 6545
rect 2320 6490 2430 6510
rect 2320 6455 2325 6490
rect 2425 6455 2430 6490
rect 2320 6430 2430 6455
rect 2570 6545 2680 6570
rect 2570 6510 2575 6545
rect 2675 6510 2680 6545
rect 2570 6490 2680 6510
rect 2570 6455 2575 6490
rect 2675 6455 2680 6490
rect 2570 6430 2680 6455
rect 2820 6545 2930 6570
rect 2820 6510 2825 6545
rect 2925 6510 2930 6545
rect 2820 6490 2930 6510
rect 2820 6455 2825 6490
rect 2925 6455 2930 6490
rect 2820 6430 2930 6455
rect 3070 6545 3180 6570
rect 3070 6510 3075 6545
rect 3175 6510 3180 6545
rect 3070 6490 3180 6510
rect 3070 6455 3075 6490
rect 3175 6455 3180 6490
rect 3070 6430 3180 6455
rect 3320 6545 3430 6570
rect 3320 6510 3325 6545
rect 3425 6510 3430 6545
rect 3320 6490 3430 6510
rect 3320 6455 3325 6490
rect 3425 6455 3430 6490
rect 3320 6430 3430 6455
rect 3570 6545 3680 6570
rect 3570 6510 3575 6545
rect 3675 6510 3680 6545
rect 3570 6490 3680 6510
rect 3570 6455 3575 6490
rect 3675 6455 3680 6490
rect 3570 6430 3680 6455
rect 3820 6545 3930 6570
rect 3820 6510 3825 6545
rect 3925 6510 3930 6545
rect 3820 6490 3930 6510
rect 3820 6455 3825 6490
rect 3925 6455 3930 6490
rect 3820 6430 3930 6455
rect 4070 6545 4180 6570
rect 4070 6510 4075 6545
rect 4175 6510 4180 6545
rect 4070 6490 4180 6510
rect 4070 6455 4075 6490
rect 4175 6455 4180 6490
rect 4070 6430 4180 6455
rect 4320 6545 4430 6570
rect 4320 6510 4325 6545
rect 4425 6510 4430 6545
rect 4320 6490 4430 6510
rect 4320 6455 4325 6490
rect 4425 6455 4430 6490
rect 4320 6430 4430 6455
rect 4570 6545 4680 6570
rect 4570 6510 4575 6545
rect 4675 6510 4680 6545
rect 4570 6490 4680 6510
rect 4570 6455 4575 6490
rect 4675 6455 4680 6490
rect 4570 6430 4680 6455
rect 4820 6545 4930 6570
rect 4820 6510 4825 6545
rect 4925 6510 4930 6545
rect 4820 6490 4930 6510
rect 4820 6455 4825 6490
rect 4925 6455 4930 6490
rect 4820 6430 4930 6455
rect 5070 6545 5180 6570
rect 5070 6510 5075 6545
rect 5175 6510 5180 6545
rect 5070 6490 5180 6510
rect 5070 6455 5075 6490
rect 5175 6455 5180 6490
rect 5070 6430 5180 6455
rect 5320 6545 5430 6570
rect 5320 6510 5325 6545
rect 5425 6510 5430 6545
rect 5320 6490 5430 6510
rect 5320 6455 5325 6490
rect 5425 6455 5430 6490
rect 5320 6430 5430 6455
rect 5570 6545 5680 6570
rect 5570 6510 5575 6545
rect 5675 6510 5680 6545
rect 5570 6490 5680 6510
rect 5570 6455 5575 6490
rect 5675 6455 5680 6490
rect 5570 6430 5680 6455
rect 5820 6545 5930 6570
rect 5820 6510 5825 6545
rect 5925 6510 5930 6545
rect 5820 6490 5930 6510
rect 5820 6455 5825 6490
rect 5925 6455 5930 6490
rect 5820 6430 5930 6455
rect 6070 6545 6180 6570
rect 6070 6510 6075 6545
rect 6175 6510 6180 6545
rect 6070 6490 6180 6510
rect 6070 6455 6075 6490
rect 6175 6455 6180 6490
rect 6070 6430 6180 6455
rect 6320 6545 6430 6570
rect 6320 6510 6325 6545
rect 6425 6510 6430 6545
rect 6320 6490 6430 6510
rect 6320 6455 6325 6490
rect 6425 6455 6430 6490
rect 6320 6430 6430 6455
rect 6570 6545 6680 6570
rect 6570 6510 6575 6545
rect 6675 6510 6680 6545
rect 6570 6490 6680 6510
rect 6570 6455 6575 6490
rect 6675 6455 6680 6490
rect 6570 6430 6680 6455
rect 6820 6545 6930 6570
rect 6820 6510 6825 6545
rect 6925 6510 6930 6545
rect 6820 6490 6930 6510
rect 6820 6455 6825 6490
rect 6925 6455 6930 6490
rect 6820 6430 6930 6455
rect 7070 6545 7180 6570
rect 7070 6510 7075 6545
rect 7175 6510 7180 6545
rect 7070 6490 7180 6510
rect 7070 6455 7075 6490
rect 7175 6455 7180 6490
rect 7070 6430 7180 6455
rect 7320 6545 7430 6570
rect 7320 6510 7325 6545
rect 7425 6510 7430 6545
rect 7320 6490 7430 6510
rect 7320 6455 7325 6490
rect 7425 6455 7430 6490
rect 7320 6430 7430 6455
rect 7570 6545 7680 6570
rect 7570 6510 7575 6545
rect 7675 6510 7680 6545
rect 7570 6490 7680 6510
rect 7570 6455 7575 6490
rect 7675 6455 7680 6490
rect 7570 6430 7680 6455
rect 7820 6545 7930 6570
rect 7820 6510 7825 6545
rect 7925 6510 7930 6545
rect 7820 6490 7930 6510
rect 7820 6455 7825 6490
rect 7925 6455 7930 6490
rect 7820 6430 7930 6455
rect 0 6425 8000 6430
rect 0 6325 10 6425
rect 45 6325 205 6425
rect 240 6325 260 6425
rect 295 6325 455 6425
rect 490 6325 510 6425
rect 545 6325 705 6425
rect 740 6325 760 6425
rect 795 6325 955 6425
rect 990 6325 1010 6425
rect 1045 6325 1205 6425
rect 1240 6325 1260 6425
rect 1295 6325 1455 6425
rect 1490 6325 1510 6425
rect 1545 6325 1705 6425
rect 1740 6325 1760 6425
rect 1795 6325 1955 6425
rect 1990 6325 2010 6425
rect 2045 6325 2205 6425
rect 2240 6325 2260 6425
rect 2295 6325 2455 6425
rect 2490 6325 2510 6425
rect 2545 6325 2705 6425
rect 2740 6325 2760 6425
rect 2795 6325 2955 6425
rect 2990 6325 3010 6425
rect 3045 6325 3205 6425
rect 3240 6325 3260 6425
rect 3295 6325 3455 6425
rect 3490 6325 3510 6425
rect 3545 6325 3705 6425
rect 3740 6325 3760 6425
rect 3795 6325 3955 6425
rect 3990 6325 4010 6425
rect 4045 6325 4205 6425
rect 4240 6325 4260 6425
rect 4295 6325 4455 6425
rect 4490 6325 4510 6425
rect 4545 6325 4705 6425
rect 4740 6325 4760 6425
rect 4795 6325 4955 6425
rect 4990 6325 5010 6425
rect 5045 6325 5205 6425
rect 5240 6325 5260 6425
rect 5295 6325 5455 6425
rect 5490 6325 5510 6425
rect 5545 6325 5705 6425
rect 5740 6325 5760 6425
rect 5795 6325 5955 6425
rect 5990 6325 6010 6425
rect 6045 6325 6205 6425
rect 6240 6325 6260 6425
rect 6295 6325 6455 6425
rect 6490 6325 6510 6425
rect 6545 6325 6705 6425
rect 6740 6325 6760 6425
rect 6795 6325 6955 6425
rect 6990 6325 7010 6425
rect 7045 6325 7205 6425
rect 7240 6325 7260 6425
rect 7295 6325 7455 6425
rect 7490 6325 7510 6425
rect 7545 6325 7705 6425
rect 7740 6325 7760 6425
rect 7795 6325 7955 6425
rect 7990 6325 8000 6425
rect 0 6320 8000 6325
rect 70 6295 180 6320
rect 70 6260 75 6295
rect 175 6260 180 6295
rect 70 6240 180 6260
rect 70 6205 75 6240
rect 175 6205 180 6240
rect 70 6180 180 6205
rect 320 6295 430 6320
rect 320 6260 325 6295
rect 425 6260 430 6295
rect 320 6240 430 6260
rect 320 6205 325 6240
rect 425 6205 430 6240
rect 320 6180 430 6205
rect 570 6295 680 6320
rect 570 6260 575 6295
rect 675 6260 680 6295
rect 570 6240 680 6260
rect 570 6205 575 6240
rect 675 6205 680 6240
rect 570 6180 680 6205
rect 820 6295 930 6320
rect 820 6260 825 6295
rect 925 6260 930 6295
rect 820 6240 930 6260
rect 820 6205 825 6240
rect 925 6205 930 6240
rect 820 6180 930 6205
rect 1070 6295 1180 6320
rect 1070 6260 1075 6295
rect 1175 6260 1180 6295
rect 1070 6240 1180 6260
rect 1070 6205 1075 6240
rect 1175 6205 1180 6240
rect 1070 6180 1180 6205
rect 1320 6295 1430 6320
rect 1320 6260 1325 6295
rect 1425 6260 1430 6295
rect 1320 6240 1430 6260
rect 1320 6205 1325 6240
rect 1425 6205 1430 6240
rect 1320 6180 1430 6205
rect 1570 6295 1680 6320
rect 1570 6260 1575 6295
rect 1675 6260 1680 6295
rect 1570 6240 1680 6260
rect 1570 6205 1575 6240
rect 1675 6205 1680 6240
rect 1570 6180 1680 6205
rect 1820 6295 1930 6320
rect 1820 6260 1825 6295
rect 1925 6260 1930 6295
rect 1820 6240 1930 6260
rect 1820 6205 1825 6240
rect 1925 6205 1930 6240
rect 1820 6180 1930 6205
rect 2070 6295 2180 6320
rect 2070 6260 2075 6295
rect 2175 6260 2180 6295
rect 2070 6240 2180 6260
rect 2070 6205 2075 6240
rect 2175 6205 2180 6240
rect 2070 6180 2180 6205
rect 2320 6295 2430 6320
rect 2320 6260 2325 6295
rect 2425 6260 2430 6295
rect 2320 6240 2430 6260
rect 2320 6205 2325 6240
rect 2425 6205 2430 6240
rect 2320 6180 2430 6205
rect 2570 6295 2680 6320
rect 2570 6260 2575 6295
rect 2675 6260 2680 6295
rect 2570 6240 2680 6260
rect 2570 6205 2575 6240
rect 2675 6205 2680 6240
rect 2570 6180 2680 6205
rect 2820 6295 2930 6320
rect 2820 6260 2825 6295
rect 2925 6260 2930 6295
rect 2820 6240 2930 6260
rect 2820 6205 2825 6240
rect 2925 6205 2930 6240
rect 2820 6180 2930 6205
rect 3070 6295 3180 6320
rect 3070 6260 3075 6295
rect 3175 6260 3180 6295
rect 3070 6240 3180 6260
rect 3070 6205 3075 6240
rect 3175 6205 3180 6240
rect 3070 6180 3180 6205
rect 3320 6295 3430 6320
rect 3320 6260 3325 6295
rect 3425 6260 3430 6295
rect 3320 6240 3430 6260
rect 3320 6205 3325 6240
rect 3425 6205 3430 6240
rect 3320 6180 3430 6205
rect 3570 6295 3680 6320
rect 3570 6260 3575 6295
rect 3675 6260 3680 6295
rect 3570 6240 3680 6260
rect 3570 6205 3575 6240
rect 3675 6205 3680 6240
rect 3570 6180 3680 6205
rect 3820 6295 3930 6320
rect 3820 6260 3825 6295
rect 3925 6260 3930 6295
rect 3820 6240 3930 6260
rect 3820 6205 3825 6240
rect 3925 6205 3930 6240
rect 3820 6180 3930 6205
rect 4070 6295 4180 6320
rect 4070 6260 4075 6295
rect 4175 6260 4180 6295
rect 4070 6240 4180 6260
rect 4070 6205 4075 6240
rect 4175 6205 4180 6240
rect 4070 6180 4180 6205
rect 4320 6295 4430 6320
rect 4320 6260 4325 6295
rect 4425 6260 4430 6295
rect 4320 6240 4430 6260
rect 4320 6205 4325 6240
rect 4425 6205 4430 6240
rect 4320 6180 4430 6205
rect 4570 6295 4680 6320
rect 4570 6260 4575 6295
rect 4675 6260 4680 6295
rect 4570 6240 4680 6260
rect 4570 6205 4575 6240
rect 4675 6205 4680 6240
rect 4570 6180 4680 6205
rect 4820 6295 4930 6320
rect 4820 6260 4825 6295
rect 4925 6260 4930 6295
rect 4820 6240 4930 6260
rect 4820 6205 4825 6240
rect 4925 6205 4930 6240
rect 4820 6180 4930 6205
rect 5070 6295 5180 6320
rect 5070 6260 5075 6295
rect 5175 6260 5180 6295
rect 5070 6240 5180 6260
rect 5070 6205 5075 6240
rect 5175 6205 5180 6240
rect 5070 6180 5180 6205
rect 5320 6295 5430 6320
rect 5320 6260 5325 6295
rect 5425 6260 5430 6295
rect 5320 6240 5430 6260
rect 5320 6205 5325 6240
rect 5425 6205 5430 6240
rect 5320 6180 5430 6205
rect 5570 6295 5680 6320
rect 5570 6260 5575 6295
rect 5675 6260 5680 6295
rect 5570 6240 5680 6260
rect 5570 6205 5575 6240
rect 5675 6205 5680 6240
rect 5570 6180 5680 6205
rect 5820 6295 5930 6320
rect 5820 6260 5825 6295
rect 5925 6260 5930 6295
rect 5820 6240 5930 6260
rect 5820 6205 5825 6240
rect 5925 6205 5930 6240
rect 5820 6180 5930 6205
rect 6070 6295 6180 6320
rect 6070 6260 6075 6295
rect 6175 6260 6180 6295
rect 6070 6240 6180 6260
rect 6070 6205 6075 6240
rect 6175 6205 6180 6240
rect 6070 6180 6180 6205
rect 6320 6295 6430 6320
rect 6320 6260 6325 6295
rect 6425 6260 6430 6295
rect 6320 6240 6430 6260
rect 6320 6205 6325 6240
rect 6425 6205 6430 6240
rect 6320 6180 6430 6205
rect 6570 6295 6680 6320
rect 6570 6260 6575 6295
rect 6675 6260 6680 6295
rect 6570 6240 6680 6260
rect 6570 6205 6575 6240
rect 6675 6205 6680 6240
rect 6570 6180 6680 6205
rect 6820 6295 6930 6320
rect 6820 6260 6825 6295
rect 6925 6260 6930 6295
rect 6820 6240 6930 6260
rect 6820 6205 6825 6240
rect 6925 6205 6930 6240
rect 6820 6180 6930 6205
rect 7070 6295 7180 6320
rect 7070 6260 7075 6295
rect 7175 6260 7180 6295
rect 7070 6240 7180 6260
rect 7070 6205 7075 6240
rect 7175 6205 7180 6240
rect 7070 6180 7180 6205
rect 7320 6295 7430 6320
rect 7320 6260 7325 6295
rect 7425 6260 7430 6295
rect 7320 6240 7430 6260
rect 7320 6205 7325 6240
rect 7425 6205 7430 6240
rect 7320 6180 7430 6205
rect 7570 6295 7680 6320
rect 7570 6260 7575 6295
rect 7675 6260 7680 6295
rect 7570 6240 7680 6260
rect 7570 6205 7575 6240
rect 7675 6205 7680 6240
rect 7570 6180 7680 6205
rect 7820 6295 7930 6320
rect 7820 6260 7825 6295
rect 7925 6260 7930 6295
rect 7820 6240 7930 6260
rect 7820 6205 7825 6240
rect 7925 6205 7930 6240
rect 7820 6180 7930 6205
rect 0 6175 8000 6180
rect 0 6075 10 6175
rect 45 6075 205 6175
rect 240 6075 260 6175
rect 295 6075 455 6175
rect 490 6075 510 6175
rect 545 6075 705 6175
rect 740 6075 760 6175
rect 795 6075 955 6175
rect 990 6075 1010 6175
rect 1045 6075 1205 6175
rect 1240 6075 1260 6175
rect 1295 6075 1455 6175
rect 1490 6075 1510 6175
rect 1545 6075 1705 6175
rect 1740 6075 1760 6175
rect 1795 6075 1955 6175
rect 1990 6075 2010 6175
rect 2045 6075 2205 6175
rect 2240 6075 2260 6175
rect 2295 6075 2455 6175
rect 2490 6075 2510 6175
rect 2545 6075 2705 6175
rect 2740 6075 2760 6175
rect 2795 6075 2955 6175
rect 2990 6075 3010 6175
rect 3045 6075 3205 6175
rect 3240 6075 3260 6175
rect 3295 6075 3455 6175
rect 3490 6075 3510 6175
rect 3545 6075 3705 6175
rect 3740 6075 3760 6175
rect 3795 6075 3955 6175
rect 3990 6075 4010 6175
rect 4045 6075 4205 6175
rect 4240 6075 4260 6175
rect 4295 6075 4455 6175
rect 4490 6075 4510 6175
rect 4545 6075 4705 6175
rect 4740 6075 4760 6175
rect 4795 6075 4955 6175
rect 4990 6075 5010 6175
rect 5045 6075 5205 6175
rect 5240 6075 5260 6175
rect 5295 6075 5455 6175
rect 5490 6075 5510 6175
rect 5545 6075 5705 6175
rect 5740 6075 5760 6175
rect 5795 6075 5955 6175
rect 5990 6075 6010 6175
rect 6045 6075 6205 6175
rect 6240 6075 6260 6175
rect 6295 6075 6455 6175
rect 6490 6075 6510 6175
rect 6545 6075 6705 6175
rect 6740 6075 6760 6175
rect 6795 6075 6955 6175
rect 6990 6075 7010 6175
rect 7045 6075 7205 6175
rect 7240 6075 7260 6175
rect 7295 6075 7455 6175
rect 7490 6075 7510 6175
rect 7545 6075 7705 6175
rect 7740 6075 7760 6175
rect 7795 6075 7955 6175
rect 7990 6075 8000 6175
rect 0 6070 8000 6075
rect 70 6045 180 6070
rect 70 6010 75 6045
rect 175 6010 180 6045
rect 70 5990 180 6010
rect 70 5955 75 5990
rect 175 5955 180 5990
rect 70 5930 180 5955
rect 320 6045 430 6070
rect 320 6010 325 6045
rect 425 6010 430 6045
rect 320 5990 430 6010
rect 320 5955 325 5990
rect 425 5955 430 5990
rect 320 5930 430 5955
rect 570 6045 680 6070
rect 570 6010 575 6045
rect 675 6010 680 6045
rect 570 5990 680 6010
rect 570 5955 575 5990
rect 675 5955 680 5990
rect 570 5930 680 5955
rect 820 6045 930 6070
rect 820 6010 825 6045
rect 925 6010 930 6045
rect 820 5990 930 6010
rect 820 5955 825 5990
rect 925 5955 930 5990
rect 820 5930 930 5955
rect 1070 6045 1180 6070
rect 1070 6010 1075 6045
rect 1175 6010 1180 6045
rect 1070 5990 1180 6010
rect 1070 5955 1075 5990
rect 1175 5955 1180 5990
rect 1070 5930 1180 5955
rect 1320 6045 1430 6070
rect 1320 6010 1325 6045
rect 1425 6010 1430 6045
rect 1320 5990 1430 6010
rect 1320 5955 1325 5990
rect 1425 5955 1430 5990
rect 1320 5930 1430 5955
rect 1570 6045 1680 6070
rect 1570 6010 1575 6045
rect 1675 6010 1680 6045
rect 1570 5990 1680 6010
rect 1570 5955 1575 5990
rect 1675 5955 1680 5990
rect 1570 5930 1680 5955
rect 1820 6045 1930 6070
rect 1820 6010 1825 6045
rect 1925 6010 1930 6045
rect 1820 5990 1930 6010
rect 1820 5955 1825 5990
rect 1925 5955 1930 5990
rect 1820 5930 1930 5955
rect 2070 6045 2180 6070
rect 2070 6010 2075 6045
rect 2175 6010 2180 6045
rect 2070 5990 2180 6010
rect 2070 5955 2075 5990
rect 2175 5955 2180 5990
rect 2070 5930 2180 5955
rect 2320 6045 2430 6070
rect 2320 6010 2325 6045
rect 2425 6010 2430 6045
rect 2320 5990 2430 6010
rect 2320 5955 2325 5990
rect 2425 5955 2430 5990
rect 2320 5930 2430 5955
rect 2570 6045 2680 6070
rect 2570 6010 2575 6045
rect 2675 6010 2680 6045
rect 2570 5990 2680 6010
rect 2570 5955 2575 5990
rect 2675 5955 2680 5990
rect 2570 5930 2680 5955
rect 2820 6045 2930 6070
rect 2820 6010 2825 6045
rect 2925 6010 2930 6045
rect 2820 5990 2930 6010
rect 2820 5955 2825 5990
rect 2925 5955 2930 5990
rect 2820 5930 2930 5955
rect 3070 6045 3180 6070
rect 3070 6010 3075 6045
rect 3175 6010 3180 6045
rect 3070 5990 3180 6010
rect 3070 5955 3075 5990
rect 3175 5955 3180 5990
rect 3070 5930 3180 5955
rect 3320 6045 3430 6070
rect 3320 6010 3325 6045
rect 3425 6010 3430 6045
rect 3320 5990 3430 6010
rect 3320 5955 3325 5990
rect 3425 5955 3430 5990
rect 3320 5930 3430 5955
rect 3570 6045 3680 6070
rect 3570 6010 3575 6045
rect 3675 6010 3680 6045
rect 3570 5990 3680 6010
rect 3570 5955 3575 5990
rect 3675 5955 3680 5990
rect 3570 5930 3680 5955
rect 3820 6045 3930 6070
rect 3820 6010 3825 6045
rect 3925 6010 3930 6045
rect 3820 5990 3930 6010
rect 3820 5955 3825 5990
rect 3925 5955 3930 5990
rect 3820 5930 3930 5955
rect 4070 6045 4180 6070
rect 4070 6010 4075 6045
rect 4175 6010 4180 6045
rect 4070 5990 4180 6010
rect 4070 5955 4075 5990
rect 4175 5955 4180 5990
rect 4070 5930 4180 5955
rect 4320 6045 4430 6070
rect 4320 6010 4325 6045
rect 4425 6010 4430 6045
rect 4320 5990 4430 6010
rect 4320 5955 4325 5990
rect 4425 5955 4430 5990
rect 4320 5930 4430 5955
rect 4570 6045 4680 6070
rect 4570 6010 4575 6045
rect 4675 6010 4680 6045
rect 4570 5990 4680 6010
rect 4570 5955 4575 5990
rect 4675 5955 4680 5990
rect 4570 5930 4680 5955
rect 4820 6045 4930 6070
rect 4820 6010 4825 6045
rect 4925 6010 4930 6045
rect 4820 5990 4930 6010
rect 4820 5955 4825 5990
rect 4925 5955 4930 5990
rect 4820 5930 4930 5955
rect 5070 6045 5180 6070
rect 5070 6010 5075 6045
rect 5175 6010 5180 6045
rect 5070 5990 5180 6010
rect 5070 5955 5075 5990
rect 5175 5955 5180 5990
rect 5070 5930 5180 5955
rect 5320 6045 5430 6070
rect 5320 6010 5325 6045
rect 5425 6010 5430 6045
rect 5320 5990 5430 6010
rect 5320 5955 5325 5990
rect 5425 5955 5430 5990
rect 5320 5930 5430 5955
rect 5570 6045 5680 6070
rect 5570 6010 5575 6045
rect 5675 6010 5680 6045
rect 5570 5990 5680 6010
rect 5570 5955 5575 5990
rect 5675 5955 5680 5990
rect 5570 5930 5680 5955
rect 5820 6045 5930 6070
rect 5820 6010 5825 6045
rect 5925 6010 5930 6045
rect 5820 5990 5930 6010
rect 5820 5955 5825 5990
rect 5925 5955 5930 5990
rect 5820 5930 5930 5955
rect 6070 6045 6180 6070
rect 6070 6010 6075 6045
rect 6175 6010 6180 6045
rect 6070 5990 6180 6010
rect 6070 5955 6075 5990
rect 6175 5955 6180 5990
rect 6070 5930 6180 5955
rect 6320 6045 6430 6070
rect 6320 6010 6325 6045
rect 6425 6010 6430 6045
rect 6320 5990 6430 6010
rect 6320 5955 6325 5990
rect 6425 5955 6430 5990
rect 6320 5930 6430 5955
rect 6570 6045 6680 6070
rect 6570 6010 6575 6045
rect 6675 6010 6680 6045
rect 6570 5990 6680 6010
rect 6570 5955 6575 5990
rect 6675 5955 6680 5990
rect 6570 5930 6680 5955
rect 6820 6045 6930 6070
rect 6820 6010 6825 6045
rect 6925 6010 6930 6045
rect 6820 5990 6930 6010
rect 6820 5955 6825 5990
rect 6925 5955 6930 5990
rect 6820 5930 6930 5955
rect 7070 6045 7180 6070
rect 7070 6010 7075 6045
rect 7175 6010 7180 6045
rect 7070 5990 7180 6010
rect 7070 5955 7075 5990
rect 7175 5955 7180 5990
rect 7070 5930 7180 5955
rect 7320 6045 7430 6070
rect 7320 6010 7325 6045
rect 7425 6010 7430 6045
rect 7320 5990 7430 6010
rect 7320 5955 7325 5990
rect 7425 5955 7430 5990
rect 7320 5930 7430 5955
rect 7570 6045 7680 6070
rect 7570 6010 7575 6045
rect 7675 6010 7680 6045
rect 7570 5990 7680 6010
rect 7570 5955 7575 5990
rect 7675 5955 7680 5990
rect 7570 5930 7680 5955
rect 7820 6045 7930 6070
rect 7820 6010 7825 6045
rect 7925 6010 7930 6045
rect 7820 5990 7930 6010
rect 7820 5955 7825 5990
rect 7925 5955 7930 5990
rect 7820 5930 7930 5955
rect 0 5925 8000 5930
rect 0 5825 10 5925
rect 45 5825 205 5925
rect 240 5825 260 5925
rect 295 5825 455 5925
rect 490 5825 510 5925
rect 545 5825 705 5925
rect 740 5825 760 5925
rect 795 5825 955 5925
rect 990 5825 1010 5925
rect 1045 5825 1205 5925
rect 1240 5825 1260 5925
rect 1295 5825 1455 5925
rect 1490 5825 1510 5925
rect 1545 5825 1705 5925
rect 1740 5825 1760 5925
rect 1795 5825 1955 5925
rect 1990 5825 2010 5925
rect 2045 5825 2205 5925
rect 2240 5825 2260 5925
rect 2295 5825 2455 5925
rect 2490 5825 2510 5925
rect 2545 5825 2705 5925
rect 2740 5825 2760 5925
rect 2795 5825 2955 5925
rect 2990 5825 3010 5925
rect 3045 5825 3205 5925
rect 3240 5825 3260 5925
rect 3295 5825 3455 5925
rect 3490 5825 3510 5925
rect 3545 5825 3705 5925
rect 3740 5825 3760 5925
rect 3795 5825 3955 5925
rect 3990 5825 4010 5925
rect 4045 5825 4205 5925
rect 4240 5825 4260 5925
rect 4295 5825 4455 5925
rect 4490 5825 4510 5925
rect 4545 5825 4705 5925
rect 4740 5825 4760 5925
rect 4795 5825 4955 5925
rect 4990 5825 5010 5925
rect 5045 5825 5205 5925
rect 5240 5825 5260 5925
rect 5295 5825 5455 5925
rect 5490 5825 5510 5925
rect 5545 5825 5705 5925
rect 5740 5825 5760 5925
rect 5795 5825 5955 5925
rect 5990 5825 6010 5925
rect 6045 5825 6205 5925
rect 6240 5825 6260 5925
rect 6295 5825 6455 5925
rect 6490 5825 6510 5925
rect 6545 5825 6705 5925
rect 6740 5825 6760 5925
rect 6795 5825 6955 5925
rect 6990 5825 7010 5925
rect 7045 5825 7205 5925
rect 7240 5825 7260 5925
rect 7295 5825 7455 5925
rect 7490 5825 7510 5925
rect 7545 5825 7705 5925
rect 7740 5825 7760 5925
rect 7795 5825 7955 5925
rect 7990 5825 8000 5925
rect 0 5820 8000 5825
rect 70 5795 180 5820
rect 70 5760 75 5795
rect 175 5760 180 5795
rect 70 5740 180 5760
rect 70 5705 75 5740
rect 175 5705 180 5740
rect 70 5680 180 5705
rect 320 5795 430 5820
rect 320 5760 325 5795
rect 425 5760 430 5795
rect 320 5740 430 5760
rect 320 5705 325 5740
rect 425 5705 430 5740
rect 320 5680 430 5705
rect 570 5795 680 5820
rect 570 5760 575 5795
rect 675 5760 680 5795
rect 570 5740 680 5760
rect 570 5705 575 5740
rect 675 5705 680 5740
rect 570 5680 680 5705
rect 820 5795 930 5820
rect 820 5760 825 5795
rect 925 5760 930 5795
rect 820 5740 930 5760
rect 820 5705 825 5740
rect 925 5705 930 5740
rect 820 5680 930 5705
rect 1070 5795 1180 5820
rect 1070 5760 1075 5795
rect 1175 5760 1180 5795
rect 1070 5740 1180 5760
rect 1070 5705 1075 5740
rect 1175 5705 1180 5740
rect 1070 5680 1180 5705
rect 1320 5795 1430 5820
rect 1320 5760 1325 5795
rect 1425 5760 1430 5795
rect 1320 5740 1430 5760
rect 1320 5705 1325 5740
rect 1425 5705 1430 5740
rect 1320 5680 1430 5705
rect 1570 5795 1680 5820
rect 1570 5760 1575 5795
rect 1675 5760 1680 5795
rect 1570 5740 1680 5760
rect 1570 5705 1575 5740
rect 1675 5705 1680 5740
rect 1570 5680 1680 5705
rect 1820 5795 1930 5820
rect 1820 5760 1825 5795
rect 1925 5760 1930 5795
rect 1820 5740 1930 5760
rect 1820 5705 1825 5740
rect 1925 5705 1930 5740
rect 1820 5680 1930 5705
rect 2070 5795 2180 5820
rect 2070 5760 2075 5795
rect 2175 5760 2180 5795
rect 2070 5740 2180 5760
rect 2070 5705 2075 5740
rect 2175 5705 2180 5740
rect 2070 5680 2180 5705
rect 2320 5795 2430 5820
rect 2320 5760 2325 5795
rect 2425 5760 2430 5795
rect 2320 5740 2430 5760
rect 2320 5705 2325 5740
rect 2425 5705 2430 5740
rect 2320 5680 2430 5705
rect 2570 5795 2680 5820
rect 2570 5760 2575 5795
rect 2675 5760 2680 5795
rect 2570 5740 2680 5760
rect 2570 5705 2575 5740
rect 2675 5705 2680 5740
rect 2570 5680 2680 5705
rect 2820 5795 2930 5820
rect 2820 5760 2825 5795
rect 2925 5760 2930 5795
rect 2820 5740 2930 5760
rect 2820 5705 2825 5740
rect 2925 5705 2930 5740
rect 2820 5680 2930 5705
rect 3070 5795 3180 5820
rect 3070 5760 3075 5795
rect 3175 5760 3180 5795
rect 3070 5740 3180 5760
rect 3070 5705 3075 5740
rect 3175 5705 3180 5740
rect 3070 5680 3180 5705
rect 3320 5795 3430 5820
rect 3320 5760 3325 5795
rect 3425 5760 3430 5795
rect 3320 5740 3430 5760
rect 3320 5705 3325 5740
rect 3425 5705 3430 5740
rect 3320 5680 3430 5705
rect 3570 5795 3680 5820
rect 3570 5760 3575 5795
rect 3675 5760 3680 5795
rect 3570 5740 3680 5760
rect 3570 5705 3575 5740
rect 3675 5705 3680 5740
rect 3570 5680 3680 5705
rect 3820 5795 3930 5820
rect 3820 5760 3825 5795
rect 3925 5760 3930 5795
rect 3820 5740 3930 5760
rect 3820 5705 3825 5740
rect 3925 5705 3930 5740
rect 3820 5680 3930 5705
rect 4070 5795 4180 5820
rect 4070 5760 4075 5795
rect 4175 5760 4180 5795
rect 4070 5740 4180 5760
rect 4070 5705 4075 5740
rect 4175 5705 4180 5740
rect 4070 5680 4180 5705
rect 4320 5795 4430 5820
rect 4320 5760 4325 5795
rect 4425 5760 4430 5795
rect 4320 5740 4430 5760
rect 4320 5705 4325 5740
rect 4425 5705 4430 5740
rect 4320 5680 4430 5705
rect 4570 5795 4680 5820
rect 4570 5760 4575 5795
rect 4675 5760 4680 5795
rect 4570 5740 4680 5760
rect 4570 5705 4575 5740
rect 4675 5705 4680 5740
rect 4570 5680 4680 5705
rect 4820 5795 4930 5820
rect 4820 5760 4825 5795
rect 4925 5760 4930 5795
rect 4820 5740 4930 5760
rect 4820 5705 4825 5740
rect 4925 5705 4930 5740
rect 4820 5680 4930 5705
rect 5070 5795 5180 5820
rect 5070 5760 5075 5795
rect 5175 5760 5180 5795
rect 5070 5740 5180 5760
rect 5070 5705 5075 5740
rect 5175 5705 5180 5740
rect 5070 5680 5180 5705
rect 5320 5795 5430 5820
rect 5320 5760 5325 5795
rect 5425 5760 5430 5795
rect 5320 5740 5430 5760
rect 5320 5705 5325 5740
rect 5425 5705 5430 5740
rect 5320 5680 5430 5705
rect 5570 5795 5680 5820
rect 5570 5760 5575 5795
rect 5675 5760 5680 5795
rect 5570 5740 5680 5760
rect 5570 5705 5575 5740
rect 5675 5705 5680 5740
rect 5570 5680 5680 5705
rect 5820 5795 5930 5820
rect 5820 5760 5825 5795
rect 5925 5760 5930 5795
rect 5820 5740 5930 5760
rect 5820 5705 5825 5740
rect 5925 5705 5930 5740
rect 5820 5680 5930 5705
rect 6070 5795 6180 5820
rect 6070 5760 6075 5795
rect 6175 5760 6180 5795
rect 6070 5740 6180 5760
rect 6070 5705 6075 5740
rect 6175 5705 6180 5740
rect 6070 5680 6180 5705
rect 6320 5795 6430 5820
rect 6320 5760 6325 5795
rect 6425 5760 6430 5795
rect 6320 5740 6430 5760
rect 6320 5705 6325 5740
rect 6425 5705 6430 5740
rect 6320 5680 6430 5705
rect 6570 5795 6680 5820
rect 6570 5760 6575 5795
rect 6675 5760 6680 5795
rect 6570 5740 6680 5760
rect 6570 5705 6575 5740
rect 6675 5705 6680 5740
rect 6570 5680 6680 5705
rect 6820 5795 6930 5820
rect 6820 5760 6825 5795
rect 6925 5760 6930 5795
rect 6820 5740 6930 5760
rect 6820 5705 6825 5740
rect 6925 5705 6930 5740
rect 6820 5680 6930 5705
rect 7070 5795 7180 5820
rect 7070 5760 7075 5795
rect 7175 5760 7180 5795
rect 7070 5740 7180 5760
rect 7070 5705 7075 5740
rect 7175 5705 7180 5740
rect 7070 5680 7180 5705
rect 7320 5795 7430 5820
rect 7320 5760 7325 5795
rect 7425 5760 7430 5795
rect 7320 5740 7430 5760
rect 7320 5705 7325 5740
rect 7425 5705 7430 5740
rect 7320 5680 7430 5705
rect 7570 5795 7680 5820
rect 7570 5760 7575 5795
rect 7675 5760 7680 5795
rect 7570 5740 7680 5760
rect 7570 5705 7575 5740
rect 7675 5705 7680 5740
rect 7570 5680 7680 5705
rect 7820 5795 7930 5820
rect 7820 5760 7825 5795
rect 7925 5760 7930 5795
rect 7820 5740 7930 5760
rect 7820 5705 7825 5740
rect 7925 5705 7930 5740
rect 7820 5680 7930 5705
rect 0 5675 8000 5680
rect 0 5575 10 5675
rect 45 5575 205 5675
rect 240 5575 260 5675
rect 295 5575 455 5675
rect 490 5575 510 5675
rect 545 5575 705 5675
rect 740 5575 760 5675
rect 795 5575 955 5675
rect 990 5575 1010 5675
rect 1045 5575 1205 5675
rect 1240 5575 1260 5675
rect 1295 5575 1455 5675
rect 1490 5575 1510 5675
rect 1545 5575 1705 5675
rect 1740 5575 1760 5675
rect 1795 5575 1955 5675
rect 1990 5575 2010 5675
rect 2045 5575 2205 5675
rect 2240 5575 2260 5675
rect 2295 5575 2455 5675
rect 2490 5575 2510 5675
rect 2545 5575 2705 5675
rect 2740 5575 2760 5675
rect 2795 5575 2955 5675
rect 2990 5575 3010 5675
rect 3045 5575 3205 5675
rect 3240 5575 3260 5675
rect 3295 5575 3455 5675
rect 3490 5575 3510 5675
rect 3545 5575 3705 5675
rect 3740 5575 3760 5675
rect 3795 5575 3955 5675
rect 3990 5575 4010 5675
rect 4045 5575 4205 5675
rect 4240 5575 4260 5675
rect 4295 5575 4455 5675
rect 4490 5575 4510 5675
rect 4545 5575 4705 5675
rect 4740 5575 4760 5675
rect 4795 5575 4955 5675
rect 4990 5575 5010 5675
rect 5045 5575 5205 5675
rect 5240 5575 5260 5675
rect 5295 5575 5455 5675
rect 5490 5575 5510 5675
rect 5545 5575 5705 5675
rect 5740 5575 5760 5675
rect 5795 5575 5955 5675
rect 5990 5575 6010 5675
rect 6045 5575 6205 5675
rect 6240 5575 6260 5675
rect 6295 5575 6455 5675
rect 6490 5575 6510 5675
rect 6545 5575 6705 5675
rect 6740 5575 6760 5675
rect 6795 5575 6955 5675
rect 6990 5575 7010 5675
rect 7045 5575 7205 5675
rect 7240 5575 7260 5675
rect 7295 5575 7455 5675
rect 7490 5575 7510 5675
rect 7545 5575 7705 5675
rect 7740 5575 7760 5675
rect 7795 5575 7955 5675
rect 7990 5575 8000 5675
rect 0 5570 8000 5575
rect 70 5545 180 5570
rect 70 5510 75 5545
rect 175 5510 180 5545
rect 70 5490 180 5510
rect 70 5455 75 5490
rect 175 5455 180 5490
rect 70 5430 180 5455
rect 320 5545 430 5570
rect 320 5510 325 5545
rect 425 5510 430 5545
rect 320 5490 430 5510
rect 320 5455 325 5490
rect 425 5455 430 5490
rect 320 5430 430 5455
rect 570 5545 680 5570
rect 570 5510 575 5545
rect 675 5510 680 5545
rect 570 5490 680 5510
rect 570 5455 575 5490
rect 675 5455 680 5490
rect 570 5430 680 5455
rect 820 5545 930 5570
rect 820 5510 825 5545
rect 925 5510 930 5545
rect 820 5490 930 5510
rect 820 5455 825 5490
rect 925 5455 930 5490
rect 820 5430 930 5455
rect 1070 5545 1180 5570
rect 1070 5510 1075 5545
rect 1175 5510 1180 5545
rect 1070 5490 1180 5510
rect 1070 5455 1075 5490
rect 1175 5455 1180 5490
rect 1070 5430 1180 5455
rect 1320 5545 1430 5570
rect 1320 5510 1325 5545
rect 1425 5510 1430 5545
rect 1320 5490 1430 5510
rect 1320 5455 1325 5490
rect 1425 5455 1430 5490
rect 1320 5430 1430 5455
rect 1570 5545 1680 5570
rect 1570 5510 1575 5545
rect 1675 5510 1680 5545
rect 1570 5490 1680 5510
rect 1570 5455 1575 5490
rect 1675 5455 1680 5490
rect 1570 5430 1680 5455
rect 1820 5545 1930 5570
rect 1820 5510 1825 5545
rect 1925 5510 1930 5545
rect 1820 5490 1930 5510
rect 1820 5455 1825 5490
rect 1925 5455 1930 5490
rect 1820 5430 1930 5455
rect 2070 5545 2180 5570
rect 2070 5510 2075 5545
rect 2175 5510 2180 5545
rect 2070 5490 2180 5510
rect 2070 5455 2075 5490
rect 2175 5455 2180 5490
rect 2070 5430 2180 5455
rect 2320 5545 2430 5570
rect 2320 5510 2325 5545
rect 2425 5510 2430 5545
rect 2320 5490 2430 5510
rect 2320 5455 2325 5490
rect 2425 5455 2430 5490
rect 2320 5430 2430 5455
rect 2570 5545 2680 5570
rect 2570 5510 2575 5545
rect 2675 5510 2680 5545
rect 2570 5490 2680 5510
rect 2570 5455 2575 5490
rect 2675 5455 2680 5490
rect 2570 5430 2680 5455
rect 2820 5545 2930 5570
rect 2820 5510 2825 5545
rect 2925 5510 2930 5545
rect 2820 5490 2930 5510
rect 2820 5455 2825 5490
rect 2925 5455 2930 5490
rect 2820 5430 2930 5455
rect 3070 5545 3180 5570
rect 3070 5510 3075 5545
rect 3175 5510 3180 5545
rect 3070 5490 3180 5510
rect 3070 5455 3075 5490
rect 3175 5455 3180 5490
rect 3070 5430 3180 5455
rect 3320 5545 3430 5570
rect 3320 5510 3325 5545
rect 3425 5510 3430 5545
rect 3320 5490 3430 5510
rect 3320 5455 3325 5490
rect 3425 5455 3430 5490
rect 3320 5430 3430 5455
rect 3570 5545 3680 5570
rect 3570 5510 3575 5545
rect 3675 5510 3680 5545
rect 3570 5490 3680 5510
rect 3570 5455 3575 5490
rect 3675 5455 3680 5490
rect 3570 5430 3680 5455
rect 3820 5545 3930 5570
rect 3820 5510 3825 5545
rect 3925 5510 3930 5545
rect 3820 5490 3930 5510
rect 3820 5455 3825 5490
rect 3925 5455 3930 5490
rect 3820 5430 3930 5455
rect 4070 5545 4180 5570
rect 4070 5510 4075 5545
rect 4175 5510 4180 5545
rect 4070 5490 4180 5510
rect 4070 5455 4075 5490
rect 4175 5455 4180 5490
rect 4070 5430 4180 5455
rect 4320 5545 4430 5570
rect 4320 5510 4325 5545
rect 4425 5510 4430 5545
rect 4320 5490 4430 5510
rect 4320 5455 4325 5490
rect 4425 5455 4430 5490
rect 4320 5430 4430 5455
rect 4570 5545 4680 5570
rect 4570 5510 4575 5545
rect 4675 5510 4680 5545
rect 4570 5490 4680 5510
rect 4570 5455 4575 5490
rect 4675 5455 4680 5490
rect 4570 5430 4680 5455
rect 4820 5545 4930 5570
rect 4820 5510 4825 5545
rect 4925 5510 4930 5545
rect 4820 5490 4930 5510
rect 4820 5455 4825 5490
rect 4925 5455 4930 5490
rect 4820 5430 4930 5455
rect 5070 5545 5180 5570
rect 5070 5510 5075 5545
rect 5175 5510 5180 5545
rect 5070 5490 5180 5510
rect 5070 5455 5075 5490
rect 5175 5455 5180 5490
rect 5070 5430 5180 5455
rect 5320 5545 5430 5570
rect 5320 5510 5325 5545
rect 5425 5510 5430 5545
rect 5320 5490 5430 5510
rect 5320 5455 5325 5490
rect 5425 5455 5430 5490
rect 5320 5430 5430 5455
rect 5570 5545 5680 5570
rect 5570 5510 5575 5545
rect 5675 5510 5680 5545
rect 5570 5490 5680 5510
rect 5570 5455 5575 5490
rect 5675 5455 5680 5490
rect 5570 5430 5680 5455
rect 5820 5545 5930 5570
rect 5820 5510 5825 5545
rect 5925 5510 5930 5545
rect 5820 5490 5930 5510
rect 5820 5455 5825 5490
rect 5925 5455 5930 5490
rect 5820 5430 5930 5455
rect 6070 5545 6180 5570
rect 6070 5510 6075 5545
rect 6175 5510 6180 5545
rect 6070 5490 6180 5510
rect 6070 5455 6075 5490
rect 6175 5455 6180 5490
rect 6070 5430 6180 5455
rect 6320 5545 6430 5570
rect 6320 5510 6325 5545
rect 6425 5510 6430 5545
rect 6320 5490 6430 5510
rect 6320 5455 6325 5490
rect 6425 5455 6430 5490
rect 6320 5430 6430 5455
rect 6570 5545 6680 5570
rect 6570 5510 6575 5545
rect 6675 5510 6680 5545
rect 6570 5490 6680 5510
rect 6570 5455 6575 5490
rect 6675 5455 6680 5490
rect 6570 5430 6680 5455
rect 6820 5545 6930 5570
rect 6820 5510 6825 5545
rect 6925 5510 6930 5545
rect 6820 5490 6930 5510
rect 6820 5455 6825 5490
rect 6925 5455 6930 5490
rect 6820 5430 6930 5455
rect 7070 5545 7180 5570
rect 7070 5510 7075 5545
rect 7175 5510 7180 5545
rect 7070 5490 7180 5510
rect 7070 5455 7075 5490
rect 7175 5455 7180 5490
rect 7070 5430 7180 5455
rect 7320 5545 7430 5570
rect 7320 5510 7325 5545
rect 7425 5510 7430 5545
rect 7320 5490 7430 5510
rect 7320 5455 7325 5490
rect 7425 5455 7430 5490
rect 7320 5430 7430 5455
rect 7570 5545 7680 5570
rect 7570 5510 7575 5545
rect 7675 5510 7680 5545
rect 7570 5490 7680 5510
rect 7570 5455 7575 5490
rect 7675 5455 7680 5490
rect 7570 5430 7680 5455
rect 7820 5545 7930 5570
rect 7820 5510 7825 5545
rect 7925 5510 7930 5545
rect 7820 5490 7930 5510
rect 7820 5455 7825 5490
rect 7925 5455 7930 5490
rect 7820 5430 7930 5455
rect 0 5425 8000 5430
rect 0 5325 10 5425
rect 45 5325 205 5425
rect 240 5325 260 5425
rect 295 5325 455 5425
rect 490 5325 510 5425
rect 545 5325 705 5425
rect 740 5325 760 5425
rect 795 5325 955 5425
rect 990 5325 1010 5425
rect 1045 5325 1205 5425
rect 1240 5325 1260 5425
rect 1295 5325 1455 5425
rect 1490 5325 1510 5425
rect 1545 5325 1705 5425
rect 1740 5325 1760 5425
rect 1795 5325 1955 5425
rect 1990 5325 2010 5425
rect 2045 5325 2205 5425
rect 2240 5325 2260 5425
rect 2295 5325 2455 5425
rect 2490 5325 2510 5425
rect 2545 5325 2705 5425
rect 2740 5325 2760 5425
rect 2795 5325 2955 5425
rect 2990 5325 3010 5425
rect 3045 5325 3205 5425
rect 3240 5325 3260 5425
rect 3295 5325 3455 5425
rect 3490 5325 3510 5425
rect 3545 5325 3705 5425
rect 3740 5325 3760 5425
rect 3795 5325 3955 5425
rect 3990 5325 4010 5425
rect 4045 5325 4205 5425
rect 4240 5325 4260 5425
rect 4295 5325 4455 5425
rect 4490 5325 4510 5425
rect 4545 5325 4705 5425
rect 4740 5325 4760 5425
rect 4795 5325 4955 5425
rect 4990 5325 5010 5425
rect 5045 5325 5205 5425
rect 5240 5325 5260 5425
rect 5295 5325 5455 5425
rect 5490 5325 5510 5425
rect 5545 5325 5705 5425
rect 5740 5325 5760 5425
rect 5795 5325 5955 5425
rect 5990 5325 6010 5425
rect 6045 5325 6205 5425
rect 6240 5325 6260 5425
rect 6295 5325 6455 5425
rect 6490 5325 6510 5425
rect 6545 5325 6705 5425
rect 6740 5325 6760 5425
rect 6795 5325 6955 5425
rect 6990 5325 7010 5425
rect 7045 5325 7205 5425
rect 7240 5325 7260 5425
rect 7295 5325 7455 5425
rect 7490 5325 7510 5425
rect 7545 5325 7705 5425
rect 7740 5325 7760 5425
rect 7795 5325 7955 5425
rect 7990 5325 8000 5425
rect 0 5320 8000 5325
rect 70 5295 180 5320
rect 70 5260 75 5295
rect 175 5260 180 5295
rect 70 5240 180 5260
rect 70 5205 75 5240
rect 175 5205 180 5240
rect 70 5180 180 5205
rect 320 5295 430 5320
rect 320 5260 325 5295
rect 425 5260 430 5295
rect 320 5240 430 5260
rect 320 5205 325 5240
rect 425 5205 430 5240
rect 320 5180 430 5205
rect 570 5295 680 5320
rect 570 5260 575 5295
rect 675 5260 680 5295
rect 570 5240 680 5260
rect 570 5205 575 5240
rect 675 5205 680 5240
rect 570 5180 680 5205
rect 820 5295 930 5320
rect 820 5260 825 5295
rect 925 5260 930 5295
rect 820 5240 930 5260
rect 820 5205 825 5240
rect 925 5205 930 5240
rect 820 5180 930 5205
rect 1070 5295 1180 5320
rect 1070 5260 1075 5295
rect 1175 5260 1180 5295
rect 1070 5240 1180 5260
rect 1070 5205 1075 5240
rect 1175 5205 1180 5240
rect 1070 5180 1180 5205
rect 1320 5295 1430 5320
rect 1320 5260 1325 5295
rect 1425 5260 1430 5295
rect 1320 5240 1430 5260
rect 1320 5205 1325 5240
rect 1425 5205 1430 5240
rect 1320 5180 1430 5205
rect 1570 5295 1680 5320
rect 1570 5260 1575 5295
rect 1675 5260 1680 5295
rect 1570 5240 1680 5260
rect 1570 5205 1575 5240
rect 1675 5205 1680 5240
rect 1570 5180 1680 5205
rect 1820 5295 1930 5320
rect 1820 5260 1825 5295
rect 1925 5260 1930 5295
rect 1820 5240 1930 5260
rect 1820 5205 1825 5240
rect 1925 5205 1930 5240
rect 1820 5180 1930 5205
rect 2070 5295 2180 5320
rect 2070 5260 2075 5295
rect 2175 5260 2180 5295
rect 2070 5240 2180 5260
rect 2070 5205 2075 5240
rect 2175 5205 2180 5240
rect 2070 5180 2180 5205
rect 2320 5295 2430 5320
rect 2320 5260 2325 5295
rect 2425 5260 2430 5295
rect 2320 5240 2430 5260
rect 2320 5205 2325 5240
rect 2425 5205 2430 5240
rect 2320 5180 2430 5205
rect 2570 5295 2680 5320
rect 2570 5260 2575 5295
rect 2675 5260 2680 5295
rect 2570 5240 2680 5260
rect 2570 5205 2575 5240
rect 2675 5205 2680 5240
rect 2570 5180 2680 5205
rect 2820 5295 2930 5320
rect 2820 5260 2825 5295
rect 2925 5260 2930 5295
rect 2820 5240 2930 5260
rect 2820 5205 2825 5240
rect 2925 5205 2930 5240
rect 2820 5180 2930 5205
rect 3070 5295 3180 5320
rect 3070 5260 3075 5295
rect 3175 5260 3180 5295
rect 3070 5240 3180 5260
rect 3070 5205 3075 5240
rect 3175 5205 3180 5240
rect 3070 5180 3180 5205
rect 3320 5295 3430 5320
rect 3320 5260 3325 5295
rect 3425 5260 3430 5295
rect 3320 5240 3430 5260
rect 3320 5205 3325 5240
rect 3425 5205 3430 5240
rect 3320 5180 3430 5205
rect 3570 5295 3680 5320
rect 3570 5260 3575 5295
rect 3675 5260 3680 5295
rect 3570 5240 3680 5260
rect 3570 5205 3575 5240
rect 3675 5205 3680 5240
rect 3570 5180 3680 5205
rect 3820 5295 3930 5320
rect 3820 5260 3825 5295
rect 3925 5260 3930 5295
rect 3820 5240 3930 5260
rect 3820 5205 3825 5240
rect 3925 5205 3930 5240
rect 3820 5180 3930 5205
rect 4070 5295 4180 5320
rect 4070 5260 4075 5295
rect 4175 5260 4180 5295
rect 4070 5240 4180 5260
rect 4070 5205 4075 5240
rect 4175 5205 4180 5240
rect 4070 5180 4180 5205
rect 4320 5295 4430 5320
rect 4320 5260 4325 5295
rect 4425 5260 4430 5295
rect 4320 5240 4430 5260
rect 4320 5205 4325 5240
rect 4425 5205 4430 5240
rect 4320 5180 4430 5205
rect 4570 5295 4680 5320
rect 4570 5260 4575 5295
rect 4675 5260 4680 5295
rect 4570 5240 4680 5260
rect 4570 5205 4575 5240
rect 4675 5205 4680 5240
rect 4570 5180 4680 5205
rect 4820 5295 4930 5320
rect 4820 5260 4825 5295
rect 4925 5260 4930 5295
rect 4820 5240 4930 5260
rect 4820 5205 4825 5240
rect 4925 5205 4930 5240
rect 4820 5180 4930 5205
rect 5070 5295 5180 5320
rect 5070 5260 5075 5295
rect 5175 5260 5180 5295
rect 5070 5240 5180 5260
rect 5070 5205 5075 5240
rect 5175 5205 5180 5240
rect 5070 5180 5180 5205
rect 5320 5295 5430 5320
rect 5320 5260 5325 5295
rect 5425 5260 5430 5295
rect 5320 5240 5430 5260
rect 5320 5205 5325 5240
rect 5425 5205 5430 5240
rect 5320 5180 5430 5205
rect 5570 5295 5680 5320
rect 5570 5260 5575 5295
rect 5675 5260 5680 5295
rect 5570 5240 5680 5260
rect 5570 5205 5575 5240
rect 5675 5205 5680 5240
rect 5570 5180 5680 5205
rect 5820 5295 5930 5320
rect 5820 5260 5825 5295
rect 5925 5260 5930 5295
rect 5820 5240 5930 5260
rect 5820 5205 5825 5240
rect 5925 5205 5930 5240
rect 5820 5180 5930 5205
rect 6070 5295 6180 5320
rect 6070 5260 6075 5295
rect 6175 5260 6180 5295
rect 6070 5240 6180 5260
rect 6070 5205 6075 5240
rect 6175 5205 6180 5240
rect 6070 5180 6180 5205
rect 6320 5295 6430 5320
rect 6320 5260 6325 5295
rect 6425 5260 6430 5295
rect 6320 5240 6430 5260
rect 6320 5205 6325 5240
rect 6425 5205 6430 5240
rect 6320 5180 6430 5205
rect 6570 5295 6680 5320
rect 6570 5260 6575 5295
rect 6675 5260 6680 5295
rect 6570 5240 6680 5260
rect 6570 5205 6575 5240
rect 6675 5205 6680 5240
rect 6570 5180 6680 5205
rect 6820 5295 6930 5320
rect 6820 5260 6825 5295
rect 6925 5260 6930 5295
rect 6820 5240 6930 5260
rect 6820 5205 6825 5240
rect 6925 5205 6930 5240
rect 6820 5180 6930 5205
rect 7070 5295 7180 5320
rect 7070 5260 7075 5295
rect 7175 5260 7180 5295
rect 7070 5240 7180 5260
rect 7070 5205 7075 5240
rect 7175 5205 7180 5240
rect 7070 5180 7180 5205
rect 7320 5295 7430 5320
rect 7320 5260 7325 5295
rect 7425 5260 7430 5295
rect 7320 5240 7430 5260
rect 7320 5205 7325 5240
rect 7425 5205 7430 5240
rect 7320 5180 7430 5205
rect 7570 5295 7680 5320
rect 7570 5260 7575 5295
rect 7675 5260 7680 5295
rect 7570 5240 7680 5260
rect 7570 5205 7575 5240
rect 7675 5205 7680 5240
rect 7570 5180 7680 5205
rect 7820 5295 7930 5320
rect 7820 5260 7825 5295
rect 7925 5260 7930 5295
rect 7820 5240 7930 5260
rect 7820 5205 7825 5240
rect 7925 5205 7930 5240
rect 7820 5180 7930 5205
rect 0 5175 8000 5180
rect 0 5075 10 5175
rect 45 5075 205 5175
rect 240 5075 260 5175
rect 295 5075 455 5175
rect 490 5075 510 5175
rect 545 5075 705 5175
rect 740 5075 760 5175
rect 795 5075 955 5175
rect 990 5075 1010 5175
rect 1045 5075 1205 5175
rect 1240 5075 1260 5175
rect 1295 5075 1455 5175
rect 1490 5075 1510 5175
rect 1545 5075 1705 5175
rect 1740 5075 1760 5175
rect 1795 5075 1955 5175
rect 1990 5075 2010 5175
rect 2045 5075 2205 5175
rect 2240 5075 2260 5175
rect 2295 5075 2455 5175
rect 2490 5075 2510 5175
rect 2545 5075 2705 5175
rect 2740 5075 2760 5175
rect 2795 5075 2955 5175
rect 2990 5075 3010 5175
rect 3045 5075 3205 5175
rect 3240 5075 3260 5175
rect 3295 5075 3455 5175
rect 3490 5075 3510 5175
rect 3545 5075 3705 5175
rect 3740 5075 3760 5175
rect 3795 5075 3955 5175
rect 3990 5075 4010 5175
rect 4045 5075 4205 5175
rect 4240 5075 4260 5175
rect 4295 5075 4455 5175
rect 4490 5075 4510 5175
rect 4545 5075 4705 5175
rect 4740 5075 4760 5175
rect 4795 5075 4955 5175
rect 4990 5075 5010 5175
rect 5045 5075 5205 5175
rect 5240 5075 5260 5175
rect 5295 5075 5455 5175
rect 5490 5075 5510 5175
rect 5545 5075 5705 5175
rect 5740 5075 5760 5175
rect 5795 5075 5955 5175
rect 5990 5075 6010 5175
rect 6045 5075 6205 5175
rect 6240 5075 6260 5175
rect 6295 5075 6455 5175
rect 6490 5075 6510 5175
rect 6545 5075 6705 5175
rect 6740 5075 6760 5175
rect 6795 5075 6955 5175
rect 6990 5075 7010 5175
rect 7045 5075 7205 5175
rect 7240 5075 7260 5175
rect 7295 5075 7455 5175
rect 7490 5075 7510 5175
rect 7545 5075 7705 5175
rect 7740 5075 7760 5175
rect 7795 5075 7955 5175
rect 7990 5075 8000 5175
rect 0 5070 8000 5075
rect 70 5045 180 5070
rect 70 5010 75 5045
rect 175 5010 180 5045
rect 70 4990 180 5010
rect 70 4955 75 4990
rect 175 4955 180 4990
rect 70 4930 180 4955
rect 320 5045 430 5070
rect 320 5010 325 5045
rect 425 5010 430 5045
rect 320 4990 430 5010
rect 320 4955 325 4990
rect 425 4955 430 4990
rect 320 4930 430 4955
rect 570 5045 680 5070
rect 570 5010 575 5045
rect 675 5010 680 5045
rect 570 4990 680 5010
rect 570 4955 575 4990
rect 675 4955 680 4990
rect 570 4930 680 4955
rect 820 5045 930 5070
rect 820 5010 825 5045
rect 925 5010 930 5045
rect 820 4990 930 5010
rect 820 4955 825 4990
rect 925 4955 930 4990
rect 820 4930 930 4955
rect 1070 5045 1180 5070
rect 1070 5010 1075 5045
rect 1175 5010 1180 5045
rect 1070 4990 1180 5010
rect 1070 4955 1075 4990
rect 1175 4955 1180 4990
rect 1070 4930 1180 4955
rect 1320 5045 1430 5070
rect 1320 5010 1325 5045
rect 1425 5010 1430 5045
rect 1320 4990 1430 5010
rect 1320 4955 1325 4990
rect 1425 4955 1430 4990
rect 1320 4930 1430 4955
rect 1570 5045 1680 5070
rect 1570 5010 1575 5045
rect 1675 5010 1680 5045
rect 1570 4990 1680 5010
rect 1570 4955 1575 4990
rect 1675 4955 1680 4990
rect 1570 4930 1680 4955
rect 1820 5045 1930 5070
rect 1820 5010 1825 5045
rect 1925 5010 1930 5045
rect 1820 4990 1930 5010
rect 1820 4955 1825 4990
rect 1925 4955 1930 4990
rect 1820 4930 1930 4955
rect 2070 5045 2180 5070
rect 2070 5010 2075 5045
rect 2175 5010 2180 5045
rect 2070 4990 2180 5010
rect 2070 4955 2075 4990
rect 2175 4955 2180 4990
rect 2070 4930 2180 4955
rect 2320 5045 2430 5070
rect 2320 5010 2325 5045
rect 2425 5010 2430 5045
rect 2320 4990 2430 5010
rect 2320 4955 2325 4990
rect 2425 4955 2430 4990
rect 2320 4930 2430 4955
rect 2570 5045 2680 5070
rect 2570 5010 2575 5045
rect 2675 5010 2680 5045
rect 2570 4990 2680 5010
rect 2570 4955 2575 4990
rect 2675 4955 2680 4990
rect 2570 4930 2680 4955
rect 2820 5045 2930 5070
rect 2820 5010 2825 5045
rect 2925 5010 2930 5045
rect 2820 4990 2930 5010
rect 2820 4955 2825 4990
rect 2925 4955 2930 4990
rect 2820 4930 2930 4955
rect 3070 5045 3180 5070
rect 3070 5010 3075 5045
rect 3175 5010 3180 5045
rect 3070 4990 3180 5010
rect 3070 4955 3075 4990
rect 3175 4955 3180 4990
rect 3070 4930 3180 4955
rect 3320 5045 3430 5070
rect 3320 5010 3325 5045
rect 3425 5010 3430 5045
rect 3320 4990 3430 5010
rect 3320 4955 3325 4990
rect 3425 4955 3430 4990
rect 3320 4930 3430 4955
rect 3570 5045 3680 5070
rect 3570 5010 3575 5045
rect 3675 5010 3680 5045
rect 3570 4990 3680 5010
rect 3570 4955 3575 4990
rect 3675 4955 3680 4990
rect 3570 4930 3680 4955
rect 3820 5045 3930 5070
rect 3820 5010 3825 5045
rect 3925 5010 3930 5045
rect 3820 4990 3930 5010
rect 3820 4955 3825 4990
rect 3925 4955 3930 4990
rect 3820 4930 3930 4955
rect 4070 5045 4180 5070
rect 4070 5010 4075 5045
rect 4175 5010 4180 5045
rect 4070 4990 4180 5010
rect 4070 4955 4075 4990
rect 4175 4955 4180 4990
rect 4070 4930 4180 4955
rect 4320 5045 4430 5070
rect 4320 5010 4325 5045
rect 4425 5010 4430 5045
rect 4320 4990 4430 5010
rect 4320 4955 4325 4990
rect 4425 4955 4430 4990
rect 4320 4930 4430 4955
rect 4570 5045 4680 5070
rect 4570 5010 4575 5045
rect 4675 5010 4680 5045
rect 4570 4990 4680 5010
rect 4570 4955 4575 4990
rect 4675 4955 4680 4990
rect 4570 4930 4680 4955
rect 4820 5045 4930 5070
rect 4820 5010 4825 5045
rect 4925 5010 4930 5045
rect 4820 4990 4930 5010
rect 4820 4955 4825 4990
rect 4925 4955 4930 4990
rect 4820 4930 4930 4955
rect 5070 5045 5180 5070
rect 5070 5010 5075 5045
rect 5175 5010 5180 5045
rect 5070 4990 5180 5010
rect 5070 4955 5075 4990
rect 5175 4955 5180 4990
rect 5070 4930 5180 4955
rect 5320 5045 5430 5070
rect 5320 5010 5325 5045
rect 5425 5010 5430 5045
rect 5320 4990 5430 5010
rect 5320 4955 5325 4990
rect 5425 4955 5430 4990
rect 5320 4930 5430 4955
rect 5570 5045 5680 5070
rect 5570 5010 5575 5045
rect 5675 5010 5680 5045
rect 5570 4990 5680 5010
rect 5570 4955 5575 4990
rect 5675 4955 5680 4990
rect 5570 4930 5680 4955
rect 5820 5045 5930 5070
rect 5820 5010 5825 5045
rect 5925 5010 5930 5045
rect 5820 4990 5930 5010
rect 5820 4955 5825 4990
rect 5925 4955 5930 4990
rect 5820 4930 5930 4955
rect 6070 5045 6180 5070
rect 6070 5010 6075 5045
rect 6175 5010 6180 5045
rect 6070 4990 6180 5010
rect 6070 4955 6075 4990
rect 6175 4955 6180 4990
rect 6070 4930 6180 4955
rect 6320 5045 6430 5070
rect 6320 5010 6325 5045
rect 6425 5010 6430 5045
rect 6320 4990 6430 5010
rect 6320 4955 6325 4990
rect 6425 4955 6430 4990
rect 6320 4930 6430 4955
rect 6570 5045 6680 5070
rect 6570 5010 6575 5045
rect 6675 5010 6680 5045
rect 6570 4990 6680 5010
rect 6570 4955 6575 4990
rect 6675 4955 6680 4990
rect 6570 4930 6680 4955
rect 6820 5045 6930 5070
rect 6820 5010 6825 5045
rect 6925 5010 6930 5045
rect 6820 4990 6930 5010
rect 6820 4955 6825 4990
rect 6925 4955 6930 4990
rect 6820 4930 6930 4955
rect 7070 5045 7180 5070
rect 7070 5010 7075 5045
rect 7175 5010 7180 5045
rect 7070 4990 7180 5010
rect 7070 4955 7075 4990
rect 7175 4955 7180 4990
rect 7070 4930 7180 4955
rect 7320 5045 7430 5070
rect 7320 5010 7325 5045
rect 7425 5010 7430 5045
rect 7320 4990 7430 5010
rect 7320 4955 7325 4990
rect 7425 4955 7430 4990
rect 7320 4930 7430 4955
rect 7570 5045 7680 5070
rect 7570 5010 7575 5045
rect 7675 5010 7680 5045
rect 7570 4990 7680 5010
rect 7570 4955 7575 4990
rect 7675 4955 7680 4990
rect 7570 4930 7680 4955
rect 7820 5045 7930 5070
rect 7820 5010 7825 5045
rect 7925 5010 7930 5045
rect 7820 4990 7930 5010
rect 7820 4955 7825 4990
rect 7925 4955 7930 4990
rect 7820 4930 7930 4955
rect 0 4925 8000 4930
rect 0 4825 10 4925
rect 45 4825 205 4925
rect 240 4825 260 4925
rect 295 4825 455 4925
rect 490 4825 510 4925
rect 545 4825 705 4925
rect 740 4825 760 4925
rect 795 4825 955 4925
rect 990 4825 1010 4925
rect 1045 4825 1205 4925
rect 1240 4825 1260 4925
rect 1295 4825 1455 4925
rect 1490 4825 1510 4925
rect 1545 4825 1705 4925
rect 1740 4825 1760 4925
rect 1795 4825 1955 4925
rect 1990 4825 2010 4925
rect 2045 4825 2205 4925
rect 2240 4825 2260 4925
rect 2295 4825 2455 4925
rect 2490 4825 2510 4925
rect 2545 4825 2705 4925
rect 2740 4825 2760 4925
rect 2795 4825 2955 4925
rect 2990 4825 3010 4925
rect 3045 4825 3205 4925
rect 3240 4825 3260 4925
rect 3295 4825 3455 4925
rect 3490 4825 3510 4925
rect 3545 4825 3705 4925
rect 3740 4825 3760 4925
rect 3795 4825 3955 4925
rect 3990 4825 4010 4925
rect 4045 4825 4205 4925
rect 4240 4825 4260 4925
rect 4295 4825 4455 4925
rect 4490 4825 4510 4925
rect 4545 4825 4705 4925
rect 4740 4825 4760 4925
rect 4795 4825 4955 4925
rect 4990 4825 5010 4925
rect 5045 4825 5205 4925
rect 5240 4825 5260 4925
rect 5295 4825 5455 4925
rect 5490 4825 5510 4925
rect 5545 4825 5705 4925
rect 5740 4825 5760 4925
rect 5795 4825 5955 4925
rect 5990 4825 6010 4925
rect 6045 4825 6205 4925
rect 6240 4825 6260 4925
rect 6295 4825 6455 4925
rect 6490 4825 6510 4925
rect 6545 4825 6705 4925
rect 6740 4825 6760 4925
rect 6795 4825 6955 4925
rect 6990 4825 7010 4925
rect 7045 4825 7205 4925
rect 7240 4825 7260 4925
rect 7295 4825 7455 4925
rect 7490 4825 7510 4925
rect 7545 4825 7705 4925
rect 7740 4825 7760 4925
rect 7795 4825 7955 4925
rect 7990 4825 8000 4925
rect 0 4820 8000 4825
rect 70 4795 180 4820
rect 70 4760 75 4795
rect 175 4760 180 4795
rect 70 4740 180 4760
rect 70 4705 75 4740
rect 175 4705 180 4740
rect 70 4680 180 4705
rect 320 4795 430 4820
rect 320 4760 325 4795
rect 425 4760 430 4795
rect 320 4740 430 4760
rect 320 4705 325 4740
rect 425 4705 430 4740
rect 320 4680 430 4705
rect 570 4795 680 4820
rect 570 4760 575 4795
rect 675 4760 680 4795
rect 570 4740 680 4760
rect 570 4705 575 4740
rect 675 4705 680 4740
rect 570 4680 680 4705
rect 820 4795 930 4820
rect 820 4760 825 4795
rect 925 4760 930 4795
rect 820 4740 930 4760
rect 820 4705 825 4740
rect 925 4705 930 4740
rect 820 4680 930 4705
rect 1070 4795 1180 4820
rect 1070 4760 1075 4795
rect 1175 4760 1180 4795
rect 1070 4740 1180 4760
rect 1070 4705 1075 4740
rect 1175 4705 1180 4740
rect 1070 4680 1180 4705
rect 1320 4795 1430 4820
rect 1320 4760 1325 4795
rect 1425 4760 1430 4795
rect 1320 4740 1430 4760
rect 1320 4705 1325 4740
rect 1425 4705 1430 4740
rect 1320 4680 1430 4705
rect 1570 4795 1680 4820
rect 1570 4760 1575 4795
rect 1675 4760 1680 4795
rect 1570 4740 1680 4760
rect 1570 4705 1575 4740
rect 1675 4705 1680 4740
rect 1570 4680 1680 4705
rect 1820 4795 1930 4820
rect 1820 4760 1825 4795
rect 1925 4760 1930 4795
rect 1820 4740 1930 4760
rect 1820 4705 1825 4740
rect 1925 4705 1930 4740
rect 1820 4680 1930 4705
rect 2070 4795 2180 4820
rect 2070 4760 2075 4795
rect 2175 4760 2180 4795
rect 2070 4740 2180 4760
rect 2070 4705 2075 4740
rect 2175 4705 2180 4740
rect 2070 4680 2180 4705
rect 2320 4795 2430 4820
rect 2320 4760 2325 4795
rect 2425 4760 2430 4795
rect 2320 4740 2430 4760
rect 2320 4705 2325 4740
rect 2425 4705 2430 4740
rect 2320 4680 2430 4705
rect 2570 4795 2680 4820
rect 2570 4760 2575 4795
rect 2675 4760 2680 4795
rect 2570 4740 2680 4760
rect 2570 4705 2575 4740
rect 2675 4705 2680 4740
rect 2570 4680 2680 4705
rect 2820 4795 2930 4820
rect 2820 4760 2825 4795
rect 2925 4760 2930 4795
rect 2820 4740 2930 4760
rect 2820 4705 2825 4740
rect 2925 4705 2930 4740
rect 2820 4680 2930 4705
rect 3070 4795 3180 4820
rect 3070 4760 3075 4795
rect 3175 4760 3180 4795
rect 3070 4740 3180 4760
rect 3070 4705 3075 4740
rect 3175 4705 3180 4740
rect 3070 4680 3180 4705
rect 3320 4795 3430 4820
rect 3320 4760 3325 4795
rect 3425 4760 3430 4795
rect 3320 4740 3430 4760
rect 3320 4705 3325 4740
rect 3425 4705 3430 4740
rect 3320 4680 3430 4705
rect 3570 4795 3680 4820
rect 3570 4760 3575 4795
rect 3675 4760 3680 4795
rect 3570 4740 3680 4760
rect 3570 4705 3575 4740
rect 3675 4705 3680 4740
rect 3570 4680 3680 4705
rect 3820 4795 3930 4820
rect 3820 4760 3825 4795
rect 3925 4760 3930 4795
rect 3820 4740 3930 4760
rect 3820 4705 3825 4740
rect 3925 4705 3930 4740
rect 3820 4680 3930 4705
rect 4070 4795 4180 4820
rect 4070 4760 4075 4795
rect 4175 4760 4180 4795
rect 4070 4740 4180 4760
rect 4070 4705 4075 4740
rect 4175 4705 4180 4740
rect 4070 4680 4180 4705
rect 4320 4795 4430 4820
rect 4320 4760 4325 4795
rect 4425 4760 4430 4795
rect 4320 4740 4430 4760
rect 4320 4705 4325 4740
rect 4425 4705 4430 4740
rect 4320 4680 4430 4705
rect 4570 4795 4680 4820
rect 4570 4760 4575 4795
rect 4675 4760 4680 4795
rect 4570 4740 4680 4760
rect 4570 4705 4575 4740
rect 4675 4705 4680 4740
rect 4570 4680 4680 4705
rect 4820 4795 4930 4820
rect 4820 4760 4825 4795
rect 4925 4760 4930 4795
rect 4820 4740 4930 4760
rect 4820 4705 4825 4740
rect 4925 4705 4930 4740
rect 4820 4680 4930 4705
rect 5070 4795 5180 4820
rect 5070 4760 5075 4795
rect 5175 4760 5180 4795
rect 5070 4740 5180 4760
rect 5070 4705 5075 4740
rect 5175 4705 5180 4740
rect 5070 4680 5180 4705
rect 5320 4795 5430 4820
rect 5320 4760 5325 4795
rect 5425 4760 5430 4795
rect 5320 4740 5430 4760
rect 5320 4705 5325 4740
rect 5425 4705 5430 4740
rect 5320 4680 5430 4705
rect 5570 4795 5680 4820
rect 5570 4760 5575 4795
rect 5675 4760 5680 4795
rect 5570 4740 5680 4760
rect 5570 4705 5575 4740
rect 5675 4705 5680 4740
rect 5570 4680 5680 4705
rect 5820 4795 5930 4820
rect 5820 4760 5825 4795
rect 5925 4760 5930 4795
rect 5820 4740 5930 4760
rect 5820 4705 5825 4740
rect 5925 4705 5930 4740
rect 5820 4680 5930 4705
rect 6070 4795 6180 4820
rect 6070 4760 6075 4795
rect 6175 4760 6180 4795
rect 6070 4740 6180 4760
rect 6070 4705 6075 4740
rect 6175 4705 6180 4740
rect 6070 4680 6180 4705
rect 6320 4795 6430 4820
rect 6320 4760 6325 4795
rect 6425 4760 6430 4795
rect 6320 4740 6430 4760
rect 6320 4705 6325 4740
rect 6425 4705 6430 4740
rect 6320 4680 6430 4705
rect 6570 4795 6680 4820
rect 6570 4760 6575 4795
rect 6675 4760 6680 4795
rect 6570 4740 6680 4760
rect 6570 4705 6575 4740
rect 6675 4705 6680 4740
rect 6570 4680 6680 4705
rect 6820 4795 6930 4820
rect 6820 4760 6825 4795
rect 6925 4760 6930 4795
rect 6820 4740 6930 4760
rect 6820 4705 6825 4740
rect 6925 4705 6930 4740
rect 6820 4680 6930 4705
rect 7070 4795 7180 4820
rect 7070 4760 7075 4795
rect 7175 4760 7180 4795
rect 7070 4740 7180 4760
rect 7070 4705 7075 4740
rect 7175 4705 7180 4740
rect 7070 4680 7180 4705
rect 7320 4795 7430 4820
rect 7320 4760 7325 4795
rect 7425 4760 7430 4795
rect 7320 4740 7430 4760
rect 7320 4705 7325 4740
rect 7425 4705 7430 4740
rect 7320 4680 7430 4705
rect 7570 4795 7680 4820
rect 7570 4760 7575 4795
rect 7675 4760 7680 4795
rect 7570 4740 7680 4760
rect 7570 4705 7575 4740
rect 7675 4705 7680 4740
rect 7570 4680 7680 4705
rect 7820 4795 7930 4820
rect 7820 4760 7825 4795
rect 7925 4760 7930 4795
rect 7820 4740 7930 4760
rect 7820 4705 7825 4740
rect 7925 4705 7930 4740
rect 7820 4680 7930 4705
rect 0 4675 8000 4680
rect 0 4575 10 4675
rect 45 4575 205 4675
rect 240 4575 260 4675
rect 295 4575 455 4675
rect 490 4575 510 4675
rect 545 4575 705 4675
rect 740 4575 760 4675
rect 795 4575 955 4675
rect 990 4575 1010 4675
rect 1045 4575 1205 4675
rect 1240 4575 1260 4675
rect 1295 4575 1455 4675
rect 1490 4575 1510 4675
rect 1545 4575 1705 4675
rect 1740 4575 1760 4675
rect 1795 4575 1955 4675
rect 1990 4575 2010 4675
rect 2045 4575 2205 4675
rect 2240 4575 2260 4675
rect 2295 4575 2455 4675
rect 2490 4575 2510 4675
rect 2545 4575 2705 4675
rect 2740 4575 2760 4675
rect 2795 4575 2955 4675
rect 2990 4575 3010 4675
rect 3045 4575 3205 4675
rect 3240 4575 3260 4675
rect 3295 4575 3455 4675
rect 3490 4575 3510 4675
rect 3545 4575 3705 4675
rect 3740 4575 3760 4675
rect 3795 4575 3955 4675
rect 3990 4575 4010 4675
rect 4045 4575 4205 4675
rect 4240 4575 4260 4675
rect 4295 4575 4455 4675
rect 4490 4575 4510 4675
rect 4545 4575 4705 4675
rect 4740 4575 4760 4675
rect 4795 4575 4955 4675
rect 4990 4575 5010 4675
rect 5045 4575 5205 4675
rect 5240 4575 5260 4675
rect 5295 4575 5455 4675
rect 5490 4575 5510 4675
rect 5545 4575 5705 4675
rect 5740 4575 5760 4675
rect 5795 4575 5955 4675
rect 5990 4575 6010 4675
rect 6045 4575 6205 4675
rect 6240 4575 6260 4675
rect 6295 4575 6455 4675
rect 6490 4575 6510 4675
rect 6545 4575 6705 4675
rect 6740 4575 6760 4675
rect 6795 4575 6955 4675
rect 6990 4575 7010 4675
rect 7045 4575 7205 4675
rect 7240 4575 7260 4675
rect 7295 4575 7455 4675
rect 7490 4575 7510 4675
rect 7545 4575 7705 4675
rect 7740 4575 7760 4675
rect 7795 4575 7955 4675
rect 7990 4575 8000 4675
rect 0 4570 8000 4575
rect 70 4545 180 4570
rect 70 4510 75 4545
rect 175 4510 180 4545
rect 70 4490 180 4510
rect 70 4455 75 4490
rect 175 4455 180 4490
rect 70 4430 180 4455
rect 320 4545 430 4570
rect 320 4510 325 4545
rect 425 4510 430 4545
rect 320 4490 430 4510
rect 320 4455 325 4490
rect 425 4455 430 4490
rect 320 4430 430 4455
rect 570 4545 680 4570
rect 570 4510 575 4545
rect 675 4510 680 4545
rect 570 4490 680 4510
rect 570 4455 575 4490
rect 675 4455 680 4490
rect 570 4430 680 4455
rect 820 4545 930 4570
rect 820 4510 825 4545
rect 925 4510 930 4545
rect 820 4490 930 4510
rect 820 4455 825 4490
rect 925 4455 930 4490
rect 820 4430 930 4455
rect 1070 4545 1180 4570
rect 1070 4510 1075 4545
rect 1175 4510 1180 4545
rect 1070 4490 1180 4510
rect 1070 4455 1075 4490
rect 1175 4455 1180 4490
rect 1070 4430 1180 4455
rect 1320 4545 1430 4570
rect 1320 4510 1325 4545
rect 1425 4510 1430 4545
rect 1320 4490 1430 4510
rect 1320 4455 1325 4490
rect 1425 4455 1430 4490
rect 1320 4430 1430 4455
rect 1570 4545 1680 4570
rect 1570 4510 1575 4545
rect 1675 4510 1680 4545
rect 1570 4490 1680 4510
rect 1570 4455 1575 4490
rect 1675 4455 1680 4490
rect 1570 4430 1680 4455
rect 1820 4545 1930 4570
rect 1820 4510 1825 4545
rect 1925 4510 1930 4545
rect 1820 4490 1930 4510
rect 1820 4455 1825 4490
rect 1925 4455 1930 4490
rect 1820 4430 1930 4455
rect 2070 4545 2180 4570
rect 2070 4510 2075 4545
rect 2175 4510 2180 4545
rect 2070 4490 2180 4510
rect 2070 4455 2075 4490
rect 2175 4455 2180 4490
rect 2070 4430 2180 4455
rect 2320 4545 2430 4570
rect 2320 4510 2325 4545
rect 2425 4510 2430 4545
rect 2320 4490 2430 4510
rect 2320 4455 2325 4490
rect 2425 4455 2430 4490
rect 2320 4430 2430 4455
rect 2570 4545 2680 4570
rect 2570 4510 2575 4545
rect 2675 4510 2680 4545
rect 2570 4490 2680 4510
rect 2570 4455 2575 4490
rect 2675 4455 2680 4490
rect 2570 4430 2680 4455
rect 2820 4545 2930 4570
rect 2820 4510 2825 4545
rect 2925 4510 2930 4545
rect 2820 4490 2930 4510
rect 2820 4455 2825 4490
rect 2925 4455 2930 4490
rect 2820 4430 2930 4455
rect 3070 4545 3180 4570
rect 3070 4510 3075 4545
rect 3175 4510 3180 4545
rect 3070 4490 3180 4510
rect 3070 4455 3075 4490
rect 3175 4455 3180 4490
rect 3070 4430 3180 4455
rect 3320 4545 3430 4570
rect 3320 4510 3325 4545
rect 3425 4510 3430 4545
rect 3320 4490 3430 4510
rect 3320 4455 3325 4490
rect 3425 4455 3430 4490
rect 3320 4430 3430 4455
rect 3570 4545 3680 4570
rect 3570 4510 3575 4545
rect 3675 4510 3680 4545
rect 3570 4490 3680 4510
rect 3570 4455 3575 4490
rect 3675 4455 3680 4490
rect 3570 4430 3680 4455
rect 3820 4545 3930 4570
rect 3820 4510 3825 4545
rect 3925 4510 3930 4545
rect 3820 4490 3930 4510
rect 3820 4455 3825 4490
rect 3925 4455 3930 4490
rect 3820 4430 3930 4455
rect 4070 4545 4180 4570
rect 4070 4510 4075 4545
rect 4175 4510 4180 4545
rect 4070 4490 4180 4510
rect 4070 4455 4075 4490
rect 4175 4455 4180 4490
rect 4070 4430 4180 4455
rect 4320 4545 4430 4570
rect 4320 4510 4325 4545
rect 4425 4510 4430 4545
rect 4320 4490 4430 4510
rect 4320 4455 4325 4490
rect 4425 4455 4430 4490
rect 4320 4430 4430 4455
rect 4570 4545 4680 4570
rect 4570 4510 4575 4545
rect 4675 4510 4680 4545
rect 4570 4490 4680 4510
rect 4570 4455 4575 4490
rect 4675 4455 4680 4490
rect 4570 4430 4680 4455
rect 4820 4545 4930 4570
rect 4820 4510 4825 4545
rect 4925 4510 4930 4545
rect 4820 4490 4930 4510
rect 4820 4455 4825 4490
rect 4925 4455 4930 4490
rect 4820 4430 4930 4455
rect 5070 4545 5180 4570
rect 5070 4510 5075 4545
rect 5175 4510 5180 4545
rect 5070 4490 5180 4510
rect 5070 4455 5075 4490
rect 5175 4455 5180 4490
rect 5070 4430 5180 4455
rect 5320 4545 5430 4570
rect 5320 4510 5325 4545
rect 5425 4510 5430 4545
rect 5320 4490 5430 4510
rect 5320 4455 5325 4490
rect 5425 4455 5430 4490
rect 5320 4430 5430 4455
rect 5570 4545 5680 4570
rect 5570 4510 5575 4545
rect 5675 4510 5680 4545
rect 5570 4490 5680 4510
rect 5570 4455 5575 4490
rect 5675 4455 5680 4490
rect 5570 4430 5680 4455
rect 5820 4545 5930 4570
rect 5820 4510 5825 4545
rect 5925 4510 5930 4545
rect 5820 4490 5930 4510
rect 5820 4455 5825 4490
rect 5925 4455 5930 4490
rect 5820 4430 5930 4455
rect 6070 4545 6180 4570
rect 6070 4510 6075 4545
rect 6175 4510 6180 4545
rect 6070 4490 6180 4510
rect 6070 4455 6075 4490
rect 6175 4455 6180 4490
rect 6070 4430 6180 4455
rect 6320 4545 6430 4570
rect 6320 4510 6325 4545
rect 6425 4510 6430 4545
rect 6320 4490 6430 4510
rect 6320 4455 6325 4490
rect 6425 4455 6430 4490
rect 6320 4430 6430 4455
rect 6570 4545 6680 4570
rect 6570 4510 6575 4545
rect 6675 4510 6680 4545
rect 6570 4490 6680 4510
rect 6570 4455 6575 4490
rect 6675 4455 6680 4490
rect 6570 4430 6680 4455
rect 6820 4545 6930 4570
rect 6820 4510 6825 4545
rect 6925 4510 6930 4545
rect 6820 4490 6930 4510
rect 6820 4455 6825 4490
rect 6925 4455 6930 4490
rect 6820 4430 6930 4455
rect 7070 4545 7180 4570
rect 7070 4510 7075 4545
rect 7175 4510 7180 4545
rect 7070 4490 7180 4510
rect 7070 4455 7075 4490
rect 7175 4455 7180 4490
rect 7070 4430 7180 4455
rect 7320 4545 7430 4570
rect 7320 4510 7325 4545
rect 7425 4510 7430 4545
rect 7320 4490 7430 4510
rect 7320 4455 7325 4490
rect 7425 4455 7430 4490
rect 7320 4430 7430 4455
rect 7570 4545 7680 4570
rect 7570 4510 7575 4545
rect 7675 4510 7680 4545
rect 7570 4490 7680 4510
rect 7570 4455 7575 4490
rect 7675 4455 7680 4490
rect 7570 4430 7680 4455
rect 7820 4545 7930 4570
rect 7820 4510 7825 4545
rect 7925 4510 7930 4545
rect 7820 4490 7930 4510
rect 7820 4455 7825 4490
rect 7925 4455 7930 4490
rect 7820 4430 7930 4455
rect 0 4425 8000 4430
rect 0 4325 10 4425
rect 45 4325 205 4425
rect 240 4325 260 4425
rect 295 4325 455 4425
rect 490 4325 510 4425
rect 545 4325 705 4425
rect 740 4325 760 4425
rect 795 4325 955 4425
rect 990 4325 1010 4425
rect 1045 4325 1205 4425
rect 1240 4325 1260 4425
rect 1295 4325 1455 4425
rect 1490 4325 1510 4425
rect 1545 4325 1705 4425
rect 1740 4325 1760 4425
rect 1795 4325 1955 4425
rect 1990 4325 2010 4425
rect 2045 4325 2205 4425
rect 2240 4325 2260 4425
rect 2295 4325 2455 4425
rect 2490 4325 2510 4425
rect 2545 4325 2705 4425
rect 2740 4325 2760 4425
rect 2795 4325 2955 4425
rect 2990 4325 3010 4425
rect 3045 4325 3205 4425
rect 3240 4325 3260 4425
rect 3295 4325 3455 4425
rect 3490 4325 3510 4425
rect 3545 4325 3705 4425
rect 3740 4325 3760 4425
rect 3795 4325 3955 4425
rect 3990 4325 4010 4425
rect 4045 4325 4205 4425
rect 4240 4325 4260 4425
rect 4295 4325 4455 4425
rect 4490 4325 4510 4425
rect 4545 4325 4705 4425
rect 4740 4325 4760 4425
rect 4795 4325 4955 4425
rect 4990 4325 5010 4425
rect 5045 4325 5205 4425
rect 5240 4325 5260 4425
rect 5295 4325 5455 4425
rect 5490 4325 5510 4425
rect 5545 4325 5705 4425
rect 5740 4325 5760 4425
rect 5795 4325 5955 4425
rect 5990 4325 6010 4425
rect 6045 4325 6205 4425
rect 6240 4325 6260 4425
rect 6295 4325 6455 4425
rect 6490 4325 6510 4425
rect 6545 4325 6705 4425
rect 6740 4325 6760 4425
rect 6795 4325 6955 4425
rect 6990 4325 7010 4425
rect 7045 4325 7205 4425
rect 7240 4325 7260 4425
rect 7295 4325 7455 4425
rect 7490 4325 7510 4425
rect 7545 4325 7705 4425
rect 7740 4325 7760 4425
rect 7795 4325 7955 4425
rect 7990 4325 8000 4425
rect 0 4320 8000 4325
rect 70 4295 180 4320
rect 70 4260 75 4295
rect 175 4260 180 4295
rect 70 4240 180 4260
rect 70 4205 75 4240
rect 175 4205 180 4240
rect 70 4180 180 4205
rect 320 4295 430 4320
rect 320 4260 325 4295
rect 425 4260 430 4295
rect 320 4240 430 4260
rect 320 4205 325 4240
rect 425 4205 430 4240
rect 320 4180 430 4205
rect 570 4295 680 4320
rect 570 4260 575 4295
rect 675 4260 680 4295
rect 570 4240 680 4260
rect 570 4205 575 4240
rect 675 4205 680 4240
rect 570 4180 680 4205
rect 820 4295 930 4320
rect 820 4260 825 4295
rect 925 4260 930 4295
rect 820 4240 930 4260
rect 820 4205 825 4240
rect 925 4205 930 4240
rect 820 4180 930 4205
rect 1070 4295 1180 4320
rect 1070 4260 1075 4295
rect 1175 4260 1180 4295
rect 1070 4240 1180 4260
rect 1070 4205 1075 4240
rect 1175 4205 1180 4240
rect 1070 4180 1180 4205
rect 1320 4295 1430 4320
rect 1320 4260 1325 4295
rect 1425 4260 1430 4295
rect 1320 4240 1430 4260
rect 1320 4205 1325 4240
rect 1425 4205 1430 4240
rect 1320 4180 1430 4205
rect 1570 4295 1680 4320
rect 1570 4260 1575 4295
rect 1675 4260 1680 4295
rect 1570 4240 1680 4260
rect 1570 4205 1575 4240
rect 1675 4205 1680 4240
rect 1570 4180 1680 4205
rect 1820 4295 1930 4320
rect 1820 4260 1825 4295
rect 1925 4260 1930 4295
rect 1820 4240 1930 4260
rect 1820 4205 1825 4240
rect 1925 4205 1930 4240
rect 1820 4180 1930 4205
rect 2070 4295 2180 4320
rect 2070 4260 2075 4295
rect 2175 4260 2180 4295
rect 2070 4240 2180 4260
rect 2070 4205 2075 4240
rect 2175 4205 2180 4240
rect 2070 4180 2180 4205
rect 2320 4295 2430 4320
rect 2320 4260 2325 4295
rect 2425 4260 2430 4295
rect 2320 4240 2430 4260
rect 2320 4205 2325 4240
rect 2425 4205 2430 4240
rect 2320 4180 2430 4205
rect 2570 4295 2680 4320
rect 2570 4260 2575 4295
rect 2675 4260 2680 4295
rect 2570 4240 2680 4260
rect 2570 4205 2575 4240
rect 2675 4205 2680 4240
rect 2570 4180 2680 4205
rect 2820 4295 2930 4320
rect 2820 4260 2825 4295
rect 2925 4260 2930 4295
rect 2820 4240 2930 4260
rect 2820 4205 2825 4240
rect 2925 4205 2930 4240
rect 2820 4180 2930 4205
rect 3070 4295 3180 4320
rect 3070 4260 3075 4295
rect 3175 4260 3180 4295
rect 3070 4240 3180 4260
rect 3070 4205 3075 4240
rect 3175 4205 3180 4240
rect 3070 4180 3180 4205
rect 3320 4295 3430 4320
rect 3320 4260 3325 4295
rect 3425 4260 3430 4295
rect 3320 4240 3430 4260
rect 3320 4205 3325 4240
rect 3425 4205 3430 4240
rect 3320 4180 3430 4205
rect 3570 4295 3680 4320
rect 3570 4260 3575 4295
rect 3675 4260 3680 4295
rect 3570 4240 3680 4260
rect 3570 4205 3575 4240
rect 3675 4205 3680 4240
rect 3570 4180 3680 4205
rect 3820 4295 3930 4320
rect 3820 4260 3825 4295
rect 3925 4260 3930 4295
rect 3820 4240 3930 4260
rect 3820 4205 3825 4240
rect 3925 4205 3930 4240
rect 3820 4180 3930 4205
rect 4070 4295 4180 4320
rect 4070 4260 4075 4295
rect 4175 4260 4180 4295
rect 4070 4240 4180 4260
rect 4070 4205 4075 4240
rect 4175 4205 4180 4240
rect 4070 4180 4180 4205
rect 4320 4295 4430 4320
rect 4320 4260 4325 4295
rect 4425 4260 4430 4295
rect 4320 4240 4430 4260
rect 4320 4205 4325 4240
rect 4425 4205 4430 4240
rect 4320 4180 4430 4205
rect 4570 4295 4680 4320
rect 4570 4260 4575 4295
rect 4675 4260 4680 4295
rect 4570 4240 4680 4260
rect 4570 4205 4575 4240
rect 4675 4205 4680 4240
rect 4570 4180 4680 4205
rect 4820 4295 4930 4320
rect 4820 4260 4825 4295
rect 4925 4260 4930 4295
rect 4820 4240 4930 4260
rect 4820 4205 4825 4240
rect 4925 4205 4930 4240
rect 4820 4180 4930 4205
rect 5070 4295 5180 4320
rect 5070 4260 5075 4295
rect 5175 4260 5180 4295
rect 5070 4240 5180 4260
rect 5070 4205 5075 4240
rect 5175 4205 5180 4240
rect 5070 4180 5180 4205
rect 5320 4295 5430 4320
rect 5320 4260 5325 4295
rect 5425 4260 5430 4295
rect 5320 4240 5430 4260
rect 5320 4205 5325 4240
rect 5425 4205 5430 4240
rect 5320 4180 5430 4205
rect 5570 4295 5680 4320
rect 5570 4260 5575 4295
rect 5675 4260 5680 4295
rect 5570 4240 5680 4260
rect 5570 4205 5575 4240
rect 5675 4205 5680 4240
rect 5570 4180 5680 4205
rect 5820 4295 5930 4320
rect 5820 4260 5825 4295
rect 5925 4260 5930 4295
rect 5820 4240 5930 4260
rect 5820 4205 5825 4240
rect 5925 4205 5930 4240
rect 5820 4180 5930 4205
rect 6070 4295 6180 4320
rect 6070 4260 6075 4295
rect 6175 4260 6180 4295
rect 6070 4240 6180 4260
rect 6070 4205 6075 4240
rect 6175 4205 6180 4240
rect 6070 4180 6180 4205
rect 6320 4295 6430 4320
rect 6320 4260 6325 4295
rect 6425 4260 6430 4295
rect 6320 4240 6430 4260
rect 6320 4205 6325 4240
rect 6425 4205 6430 4240
rect 6320 4180 6430 4205
rect 6570 4295 6680 4320
rect 6570 4260 6575 4295
rect 6675 4260 6680 4295
rect 6570 4240 6680 4260
rect 6570 4205 6575 4240
rect 6675 4205 6680 4240
rect 6570 4180 6680 4205
rect 6820 4295 6930 4320
rect 6820 4260 6825 4295
rect 6925 4260 6930 4295
rect 6820 4240 6930 4260
rect 6820 4205 6825 4240
rect 6925 4205 6930 4240
rect 6820 4180 6930 4205
rect 7070 4295 7180 4320
rect 7070 4260 7075 4295
rect 7175 4260 7180 4295
rect 7070 4240 7180 4260
rect 7070 4205 7075 4240
rect 7175 4205 7180 4240
rect 7070 4180 7180 4205
rect 7320 4295 7430 4320
rect 7320 4260 7325 4295
rect 7425 4260 7430 4295
rect 7320 4240 7430 4260
rect 7320 4205 7325 4240
rect 7425 4205 7430 4240
rect 7320 4180 7430 4205
rect 7570 4295 7680 4320
rect 7570 4260 7575 4295
rect 7675 4260 7680 4295
rect 7570 4240 7680 4260
rect 7570 4205 7575 4240
rect 7675 4205 7680 4240
rect 7570 4180 7680 4205
rect 7820 4295 7930 4320
rect 7820 4260 7825 4295
rect 7925 4260 7930 4295
rect 7820 4240 7930 4260
rect 7820 4205 7825 4240
rect 7925 4205 7930 4240
rect 7820 4180 7930 4205
rect 0 4175 8000 4180
rect 0 4075 10 4175
rect 45 4075 205 4175
rect 240 4075 260 4175
rect 295 4075 455 4175
rect 490 4075 510 4175
rect 545 4075 705 4175
rect 740 4075 760 4175
rect 795 4075 955 4175
rect 990 4075 1010 4175
rect 1045 4075 1205 4175
rect 1240 4075 1260 4175
rect 1295 4075 1455 4175
rect 1490 4075 1510 4175
rect 1545 4075 1705 4175
rect 1740 4075 1760 4175
rect 1795 4075 1955 4175
rect 1990 4075 2010 4175
rect 2045 4075 2205 4175
rect 2240 4075 2260 4175
rect 2295 4075 2455 4175
rect 2490 4075 2510 4175
rect 2545 4075 2705 4175
rect 2740 4075 2760 4175
rect 2795 4075 2955 4175
rect 2990 4075 3010 4175
rect 3045 4075 3205 4175
rect 3240 4075 3260 4175
rect 3295 4075 3455 4175
rect 3490 4075 3510 4175
rect 3545 4075 3705 4175
rect 3740 4075 3760 4175
rect 3795 4075 3955 4175
rect 3990 4075 4010 4175
rect 4045 4075 4205 4175
rect 4240 4075 4260 4175
rect 4295 4075 4455 4175
rect 4490 4075 4510 4175
rect 4545 4075 4705 4175
rect 4740 4075 4760 4175
rect 4795 4075 4955 4175
rect 4990 4075 5010 4175
rect 5045 4075 5205 4175
rect 5240 4075 5260 4175
rect 5295 4075 5455 4175
rect 5490 4075 5510 4175
rect 5545 4075 5705 4175
rect 5740 4075 5760 4175
rect 5795 4075 5955 4175
rect 5990 4075 6010 4175
rect 6045 4075 6205 4175
rect 6240 4075 6260 4175
rect 6295 4075 6455 4175
rect 6490 4075 6510 4175
rect 6545 4075 6705 4175
rect 6740 4075 6760 4175
rect 6795 4075 6955 4175
rect 6990 4075 7010 4175
rect 7045 4075 7205 4175
rect 7240 4075 7260 4175
rect 7295 4075 7455 4175
rect 7490 4075 7510 4175
rect 7545 4075 7705 4175
rect 7740 4075 7760 4175
rect 7795 4075 7955 4175
rect 7990 4075 8000 4175
rect 0 4070 8000 4075
rect 70 4045 180 4070
rect 70 4010 75 4045
rect 175 4010 180 4045
rect 70 3990 180 4010
rect 70 3955 75 3990
rect 175 3955 180 3990
rect 70 3930 180 3955
rect 320 4045 430 4070
rect 320 4010 325 4045
rect 425 4010 430 4045
rect 320 3990 430 4010
rect 320 3955 325 3990
rect 425 3955 430 3990
rect 320 3930 430 3955
rect 570 4045 680 4070
rect 570 4010 575 4045
rect 675 4010 680 4045
rect 570 3990 680 4010
rect 570 3955 575 3990
rect 675 3955 680 3990
rect 570 3930 680 3955
rect 820 4045 930 4070
rect 820 4010 825 4045
rect 925 4010 930 4045
rect 820 3990 930 4010
rect 820 3955 825 3990
rect 925 3955 930 3990
rect 820 3930 930 3955
rect 1070 4045 1180 4070
rect 1070 4010 1075 4045
rect 1175 4010 1180 4045
rect 1070 3990 1180 4010
rect 1070 3955 1075 3990
rect 1175 3955 1180 3990
rect 1070 3930 1180 3955
rect 1320 4045 1430 4070
rect 1320 4010 1325 4045
rect 1425 4010 1430 4045
rect 1320 3990 1430 4010
rect 1320 3955 1325 3990
rect 1425 3955 1430 3990
rect 1320 3930 1430 3955
rect 1570 4045 1680 4070
rect 1570 4010 1575 4045
rect 1675 4010 1680 4045
rect 1570 3990 1680 4010
rect 1570 3955 1575 3990
rect 1675 3955 1680 3990
rect 1570 3930 1680 3955
rect 1820 4045 1930 4070
rect 1820 4010 1825 4045
rect 1925 4010 1930 4045
rect 1820 3990 1930 4010
rect 1820 3955 1825 3990
rect 1925 3955 1930 3990
rect 1820 3930 1930 3955
rect 2070 4045 2180 4070
rect 2070 4010 2075 4045
rect 2175 4010 2180 4045
rect 2070 3990 2180 4010
rect 2070 3955 2075 3990
rect 2175 3955 2180 3990
rect 2070 3930 2180 3955
rect 2320 4045 2430 4070
rect 2320 4010 2325 4045
rect 2425 4010 2430 4045
rect 2320 3990 2430 4010
rect 2320 3955 2325 3990
rect 2425 3955 2430 3990
rect 2320 3930 2430 3955
rect 2570 4045 2680 4070
rect 2570 4010 2575 4045
rect 2675 4010 2680 4045
rect 2570 3990 2680 4010
rect 2570 3955 2575 3990
rect 2675 3955 2680 3990
rect 2570 3930 2680 3955
rect 2820 4045 2930 4070
rect 2820 4010 2825 4045
rect 2925 4010 2930 4045
rect 2820 3990 2930 4010
rect 2820 3955 2825 3990
rect 2925 3955 2930 3990
rect 2820 3930 2930 3955
rect 3070 4045 3180 4070
rect 3070 4010 3075 4045
rect 3175 4010 3180 4045
rect 3070 3990 3180 4010
rect 3070 3955 3075 3990
rect 3175 3955 3180 3990
rect 3070 3930 3180 3955
rect 3320 4045 3430 4070
rect 3320 4010 3325 4045
rect 3425 4010 3430 4045
rect 3320 3990 3430 4010
rect 3320 3955 3325 3990
rect 3425 3955 3430 3990
rect 3320 3930 3430 3955
rect 3570 4045 3680 4070
rect 3570 4010 3575 4045
rect 3675 4010 3680 4045
rect 3570 3990 3680 4010
rect 3570 3955 3575 3990
rect 3675 3955 3680 3990
rect 3570 3930 3680 3955
rect 3820 4045 3930 4070
rect 3820 4010 3825 4045
rect 3925 4010 3930 4045
rect 3820 3990 3930 4010
rect 3820 3955 3825 3990
rect 3925 3955 3930 3990
rect 3820 3930 3930 3955
rect 4070 4045 4180 4070
rect 4070 4010 4075 4045
rect 4175 4010 4180 4045
rect 4070 3990 4180 4010
rect 4070 3955 4075 3990
rect 4175 3955 4180 3990
rect 4070 3930 4180 3955
rect 4320 4045 4430 4070
rect 4320 4010 4325 4045
rect 4425 4010 4430 4045
rect 4320 3990 4430 4010
rect 4320 3955 4325 3990
rect 4425 3955 4430 3990
rect 4320 3930 4430 3955
rect 4570 4045 4680 4070
rect 4570 4010 4575 4045
rect 4675 4010 4680 4045
rect 4570 3990 4680 4010
rect 4570 3955 4575 3990
rect 4675 3955 4680 3990
rect 4570 3930 4680 3955
rect 4820 4045 4930 4070
rect 4820 4010 4825 4045
rect 4925 4010 4930 4045
rect 4820 3990 4930 4010
rect 4820 3955 4825 3990
rect 4925 3955 4930 3990
rect 4820 3930 4930 3955
rect 5070 4045 5180 4070
rect 5070 4010 5075 4045
rect 5175 4010 5180 4045
rect 5070 3990 5180 4010
rect 5070 3955 5075 3990
rect 5175 3955 5180 3990
rect 5070 3930 5180 3955
rect 5320 4045 5430 4070
rect 5320 4010 5325 4045
rect 5425 4010 5430 4045
rect 5320 3990 5430 4010
rect 5320 3955 5325 3990
rect 5425 3955 5430 3990
rect 5320 3930 5430 3955
rect 5570 4045 5680 4070
rect 5570 4010 5575 4045
rect 5675 4010 5680 4045
rect 5570 3990 5680 4010
rect 5570 3955 5575 3990
rect 5675 3955 5680 3990
rect 5570 3930 5680 3955
rect 5820 4045 5930 4070
rect 5820 4010 5825 4045
rect 5925 4010 5930 4045
rect 5820 3990 5930 4010
rect 5820 3955 5825 3990
rect 5925 3955 5930 3990
rect 5820 3930 5930 3955
rect 6070 4045 6180 4070
rect 6070 4010 6075 4045
rect 6175 4010 6180 4045
rect 6070 3990 6180 4010
rect 6070 3955 6075 3990
rect 6175 3955 6180 3990
rect 6070 3930 6180 3955
rect 6320 4045 6430 4070
rect 6320 4010 6325 4045
rect 6425 4010 6430 4045
rect 6320 3990 6430 4010
rect 6320 3955 6325 3990
rect 6425 3955 6430 3990
rect 6320 3930 6430 3955
rect 6570 4045 6680 4070
rect 6570 4010 6575 4045
rect 6675 4010 6680 4045
rect 6570 3990 6680 4010
rect 6570 3955 6575 3990
rect 6675 3955 6680 3990
rect 6570 3930 6680 3955
rect 6820 4045 6930 4070
rect 6820 4010 6825 4045
rect 6925 4010 6930 4045
rect 6820 3990 6930 4010
rect 6820 3955 6825 3990
rect 6925 3955 6930 3990
rect 6820 3930 6930 3955
rect 7070 4045 7180 4070
rect 7070 4010 7075 4045
rect 7175 4010 7180 4045
rect 7070 3990 7180 4010
rect 7070 3955 7075 3990
rect 7175 3955 7180 3990
rect 7070 3930 7180 3955
rect 7320 4045 7430 4070
rect 7320 4010 7325 4045
rect 7425 4010 7430 4045
rect 7320 3990 7430 4010
rect 7320 3955 7325 3990
rect 7425 3955 7430 3990
rect 7320 3930 7430 3955
rect 7570 4045 7680 4070
rect 7570 4010 7575 4045
rect 7675 4010 7680 4045
rect 7570 3990 7680 4010
rect 7570 3955 7575 3990
rect 7675 3955 7680 3990
rect 7570 3930 7680 3955
rect 7820 4045 7930 4070
rect 7820 4010 7825 4045
rect 7925 4010 7930 4045
rect 7820 3990 7930 4010
rect 7820 3955 7825 3990
rect 7925 3955 7930 3990
rect 7820 3930 7930 3955
rect 0 3925 8000 3930
rect 0 3825 10 3925
rect 45 3825 205 3925
rect 240 3825 260 3925
rect 295 3825 455 3925
rect 490 3825 510 3925
rect 545 3825 705 3925
rect 740 3825 760 3925
rect 795 3825 955 3925
rect 990 3825 1010 3925
rect 1045 3825 1205 3925
rect 1240 3825 1260 3925
rect 1295 3825 1455 3925
rect 1490 3825 1510 3925
rect 1545 3825 1705 3925
rect 1740 3825 1760 3925
rect 1795 3825 1955 3925
rect 1990 3825 2010 3925
rect 2045 3825 2205 3925
rect 2240 3825 2260 3925
rect 2295 3825 2455 3925
rect 2490 3825 2510 3925
rect 2545 3825 2705 3925
rect 2740 3825 2760 3925
rect 2795 3825 2955 3925
rect 2990 3825 3010 3925
rect 3045 3825 3205 3925
rect 3240 3825 3260 3925
rect 3295 3825 3455 3925
rect 3490 3825 3510 3925
rect 3545 3825 3705 3925
rect 3740 3825 3760 3925
rect 3795 3825 3955 3925
rect 3990 3825 4010 3925
rect 4045 3825 4205 3925
rect 4240 3825 4260 3925
rect 4295 3825 4455 3925
rect 4490 3825 4510 3925
rect 4545 3825 4705 3925
rect 4740 3825 4760 3925
rect 4795 3825 4955 3925
rect 4990 3825 5010 3925
rect 5045 3825 5205 3925
rect 5240 3825 5260 3925
rect 5295 3825 5455 3925
rect 5490 3825 5510 3925
rect 5545 3825 5705 3925
rect 5740 3825 5760 3925
rect 5795 3825 5955 3925
rect 5990 3825 6010 3925
rect 6045 3825 6205 3925
rect 6240 3825 6260 3925
rect 6295 3825 6455 3925
rect 6490 3825 6510 3925
rect 6545 3825 6705 3925
rect 6740 3825 6760 3925
rect 6795 3825 6955 3925
rect 6990 3825 7010 3925
rect 7045 3825 7205 3925
rect 7240 3825 7260 3925
rect 7295 3825 7455 3925
rect 7490 3825 7510 3925
rect 7545 3825 7705 3925
rect 7740 3825 7760 3925
rect 7795 3825 7955 3925
rect 7990 3825 8000 3925
rect 0 3820 8000 3825
rect 70 3795 180 3820
rect 70 3760 75 3795
rect 175 3760 180 3795
rect 70 3740 180 3760
rect 70 3705 75 3740
rect 175 3705 180 3740
rect 70 3680 180 3705
rect 320 3795 430 3820
rect 320 3760 325 3795
rect 425 3760 430 3795
rect 320 3740 430 3760
rect 320 3705 325 3740
rect 425 3705 430 3740
rect 320 3680 430 3705
rect 570 3795 680 3820
rect 570 3760 575 3795
rect 675 3760 680 3795
rect 570 3740 680 3760
rect 570 3705 575 3740
rect 675 3705 680 3740
rect 570 3680 680 3705
rect 820 3795 930 3820
rect 820 3760 825 3795
rect 925 3760 930 3795
rect 820 3740 930 3760
rect 820 3705 825 3740
rect 925 3705 930 3740
rect 820 3680 930 3705
rect 1070 3795 1180 3820
rect 1070 3760 1075 3795
rect 1175 3760 1180 3795
rect 1070 3740 1180 3760
rect 1070 3705 1075 3740
rect 1175 3705 1180 3740
rect 1070 3680 1180 3705
rect 1320 3795 1430 3820
rect 1320 3760 1325 3795
rect 1425 3760 1430 3795
rect 1320 3740 1430 3760
rect 1320 3705 1325 3740
rect 1425 3705 1430 3740
rect 1320 3680 1430 3705
rect 1570 3795 1680 3820
rect 1570 3760 1575 3795
rect 1675 3760 1680 3795
rect 1570 3740 1680 3760
rect 1570 3705 1575 3740
rect 1675 3705 1680 3740
rect 1570 3680 1680 3705
rect 1820 3795 1930 3820
rect 1820 3760 1825 3795
rect 1925 3760 1930 3795
rect 1820 3740 1930 3760
rect 1820 3705 1825 3740
rect 1925 3705 1930 3740
rect 1820 3680 1930 3705
rect 2070 3795 2180 3820
rect 2070 3760 2075 3795
rect 2175 3760 2180 3795
rect 2070 3740 2180 3760
rect 2070 3705 2075 3740
rect 2175 3705 2180 3740
rect 2070 3680 2180 3705
rect 2320 3795 2430 3820
rect 2320 3760 2325 3795
rect 2425 3760 2430 3795
rect 2320 3740 2430 3760
rect 2320 3705 2325 3740
rect 2425 3705 2430 3740
rect 2320 3680 2430 3705
rect 2570 3795 2680 3820
rect 2570 3760 2575 3795
rect 2675 3760 2680 3795
rect 2570 3740 2680 3760
rect 2570 3705 2575 3740
rect 2675 3705 2680 3740
rect 2570 3680 2680 3705
rect 2820 3795 2930 3820
rect 2820 3760 2825 3795
rect 2925 3760 2930 3795
rect 2820 3740 2930 3760
rect 2820 3705 2825 3740
rect 2925 3705 2930 3740
rect 2820 3680 2930 3705
rect 3070 3795 3180 3820
rect 3070 3760 3075 3795
rect 3175 3760 3180 3795
rect 3070 3740 3180 3760
rect 3070 3705 3075 3740
rect 3175 3705 3180 3740
rect 3070 3680 3180 3705
rect 3320 3795 3430 3820
rect 3320 3760 3325 3795
rect 3425 3760 3430 3795
rect 3320 3740 3430 3760
rect 3320 3705 3325 3740
rect 3425 3705 3430 3740
rect 3320 3680 3430 3705
rect 3570 3795 3680 3820
rect 3570 3760 3575 3795
rect 3675 3760 3680 3795
rect 3570 3740 3680 3760
rect 3570 3705 3575 3740
rect 3675 3705 3680 3740
rect 3570 3680 3680 3705
rect 3820 3795 3930 3820
rect 3820 3760 3825 3795
rect 3925 3760 3930 3795
rect 3820 3740 3930 3760
rect 3820 3705 3825 3740
rect 3925 3705 3930 3740
rect 3820 3680 3930 3705
rect 4070 3795 4180 3820
rect 4070 3760 4075 3795
rect 4175 3760 4180 3795
rect 4070 3740 4180 3760
rect 4070 3705 4075 3740
rect 4175 3705 4180 3740
rect 4070 3680 4180 3705
rect 4320 3795 4430 3820
rect 4320 3760 4325 3795
rect 4425 3760 4430 3795
rect 4320 3740 4430 3760
rect 4320 3705 4325 3740
rect 4425 3705 4430 3740
rect 4320 3680 4430 3705
rect 4570 3795 4680 3820
rect 4570 3760 4575 3795
rect 4675 3760 4680 3795
rect 4570 3740 4680 3760
rect 4570 3705 4575 3740
rect 4675 3705 4680 3740
rect 4570 3680 4680 3705
rect 4820 3795 4930 3820
rect 4820 3760 4825 3795
rect 4925 3760 4930 3795
rect 4820 3740 4930 3760
rect 4820 3705 4825 3740
rect 4925 3705 4930 3740
rect 4820 3680 4930 3705
rect 5070 3795 5180 3820
rect 5070 3760 5075 3795
rect 5175 3760 5180 3795
rect 5070 3740 5180 3760
rect 5070 3705 5075 3740
rect 5175 3705 5180 3740
rect 5070 3680 5180 3705
rect 5320 3795 5430 3820
rect 5320 3760 5325 3795
rect 5425 3760 5430 3795
rect 5320 3740 5430 3760
rect 5320 3705 5325 3740
rect 5425 3705 5430 3740
rect 5320 3680 5430 3705
rect 5570 3795 5680 3820
rect 5570 3760 5575 3795
rect 5675 3760 5680 3795
rect 5570 3740 5680 3760
rect 5570 3705 5575 3740
rect 5675 3705 5680 3740
rect 5570 3680 5680 3705
rect 5820 3795 5930 3820
rect 5820 3760 5825 3795
rect 5925 3760 5930 3795
rect 5820 3740 5930 3760
rect 5820 3705 5825 3740
rect 5925 3705 5930 3740
rect 5820 3680 5930 3705
rect 6070 3795 6180 3820
rect 6070 3760 6075 3795
rect 6175 3760 6180 3795
rect 6070 3740 6180 3760
rect 6070 3705 6075 3740
rect 6175 3705 6180 3740
rect 6070 3680 6180 3705
rect 6320 3795 6430 3820
rect 6320 3760 6325 3795
rect 6425 3760 6430 3795
rect 6320 3740 6430 3760
rect 6320 3705 6325 3740
rect 6425 3705 6430 3740
rect 6320 3680 6430 3705
rect 6570 3795 6680 3820
rect 6570 3760 6575 3795
rect 6675 3760 6680 3795
rect 6570 3740 6680 3760
rect 6570 3705 6575 3740
rect 6675 3705 6680 3740
rect 6570 3680 6680 3705
rect 6820 3795 6930 3820
rect 6820 3760 6825 3795
rect 6925 3760 6930 3795
rect 6820 3740 6930 3760
rect 6820 3705 6825 3740
rect 6925 3705 6930 3740
rect 6820 3680 6930 3705
rect 7070 3795 7180 3820
rect 7070 3760 7075 3795
rect 7175 3760 7180 3795
rect 7070 3740 7180 3760
rect 7070 3705 7075 3740
rect 7175 3705 7180 3740
rect 7070 3680 7180 3705
rect 7320 3795 7430 3820
rect 7320 3760 7325 3795
rect 7425 3760 7430 3795
rect 7320 3740 7430 3760
rect 7320 3705 7325 3740
rect 7425 3705 7430 3740
rect 7320 3680 7430 3705
rect 7570 3795 7680 3820
rect 7570 3760 7575 3795
rect 7675 3760 7680 3795
rect 7570 3740 7680 3760
rect 7570 3705 7575 3740
rect 7675 3705 7680 3740
rect 7570 3680 7680 3705
rect 7820 3795 7930 3820
rect 7820 3760 7825 3795
rect 7925 3760 7930 3795
rect 7820 3740 7930 3760
rect 7820 3705 7825 3740
rect 7925 3705 7930 3740
rect 7820 3680 7930 3705
rect 0 3675 8000 3680
rect 0 3575 10 3675
rect 45 3575 205 3675
rect 240 3575 260 3675
rect 295 3575 455 3675
rect 490 3575 510 3675
rect 545 3575 705 3675
rect 740 3575 760 3675
rect 795 3575 955 3675
rect 990 3575 1010 3675
rect 1045 3575 1205 3675
rect 1240 3575 1260 3675
rect 1295 3575 1455 3675
rect 1490 3575 1510 3675
rect 1545 3575 1705 3675
rect 1740 3575 1760 3675
rect 1795 3575 1955 3675
rect 1990 3575 2010 3675
rect 2045 3575 2205 3675
rect 2240 3575 2260 3675
rect 2295 3575 2455 3675
rect 2490 3575 2510 3675
rect 2545 3575 2705 3675
rect 2740 3575 2760 3675
rect 2795 3575 2955 3675
rect 2990 3575 3010 3675
rect 3045 3575 3205 3675
rect 3240 3575 3260 3675
rect 3295 3575 3455 3675
rect 3490 3575 3510 3675
rect 3545 3575 3705 3675
rect 3740 3575 3760 3675
rect 3795 3575 3955 3675
rect 3990 3575 4010 3675
rect 4045 3575 4205 3675
rect 4240 3575 4260 3675
rect 4295 3575 4455 3675
rect 4490 3575 4510 3675
rect 4545 3575 4705 3675
rect 4740 3575 4760 3675
rect 4795 3575 4955 3675
rect 4990 3575 5010 3675
rect 5045 3575 5205 3675
rect 5240 3575 5260 3675
rect 5295 3575 5455 3675
rect 5490 3575 5510 3675
rect 5545 3575 5705 3675
rect 5740 3575 5760 3675
rect 5795 3575 5955 3675
rect 5990 3575 6010 3675
rect 6045 3575 6205 3675
rect 6240 3575 6260 3675
rect 6295 3575 6455 3675
rect 6490 3575 6510 3675
rect 6545 3575 6705 3675
rect 6740 3575 6760 3675
rect 6795 3575 6955 3675
rect 6990 3575 7010 3675
rect 7045 3575 7205 3675
rect 7240 3575 7260 3675
rect 7295 3575 7455 3675
rect 7490 3575 7510 3675
rect 7545 3575 7705 3675
rect 7740 3575 7760 3675
rect 7795 3575 7955 3675
rect 7990 3575 8000 3675
rect 0 3570 8000 3575
rect 70 3545 180 3570
rect 70 3510 75 3545
rect 175 3510 180 3545
rect 70 3490 180 3510
rect 70 3455 75 3490
rect 175 3455 180 3490
rect 70 3430 180 3455
rect 320 3545 430 3570
rect 320 3510 325 3545
rect 425 3510 430 3545
rect 320 3490 430 3510
rect 320 3455 325 3490
rect 425 3455 430 3490
rect 320 3430 430 3455
rect 570 3545 680 3570
rect 570 3510 575 3545
rect 675 3510 680 3545
rect 570 3490 680 3510
rect 570 3455 575 3490
rect 675 3455 680 3490
rect 570 3430 680 3455
rect 820 3545 930 3570
rect 820 3510 825 3545
rect 925 3510 930 3545
rect 820 3490 930 3510
rect 820 3455 825 3490
rect 925 3455 930 3490
rect 820 3430 930 3455
rect 1070 3545 1180 3570
rect 1070 3510 1075 3545
rect 1175 3510 1180 3545
rect 1070 3490 1180 3510
rect 1070 3455 1075 3490
rect 1175 3455 1180 3490
rect 1070 3430 1180 3455
rect 1320 3545 1430 3570
rect 1320 3510 1325 3545
rect 1425 3510 1430 3545
rect 1320 3490 1430 3510
rect 1320 3455 1325 3490
rect 1425 3455 1430 3490
rect 1320 3430 1430 3455
rect 1570 3545 1680 3570
rect 1570 3510 1575 3545
rect 1675 3510 1680 3545
rect 1570 3490 1680 3510
rect 1570 3455 1575 3490
rect 1675 3455 1680 3490
rect 1570 3430 1680 3455
rect 1820 3545 1930 3570
rect 1820 3510 1825 3545
rect 1925 3510 1930 3545
rect 1820 3490 1930 3510
rect 1820 3455 1825 3490
rect 1925 3455 1930 3490
rect 1820 3430 1930 3455
rect 2070 3545 2180 3570
rect 2070 3510 2075 3545
rect 2175 3510 2180 3545
rect 2070 3490 2180 3510
rect 2070 3455 2075 3490
rect 2175 3455 2180 3490
rect 2070 3430 2180 3455
rect 2320 3545 2430 3570
rect 2320 3510 2325 3545
rect 2425 3510 2430 3545
rect 2320 3490 2430 3510
rect 2320 3455 2325 3490
rect 2425 3455 2430 3490
rect 2320 3430 2430 3455
rect 2570 3545 2680 3570
rect 2570 3510 2575 3545
rect 2675 3510 2680 3545
rect 2570 3490 2680 3510
rect 2570 3455 2575 3490
rect 2675 3455 2680 3490
rect 2570 3430 2680 3455
rect 2820 3545 2930 3570
rect 2820 3510 2825 3545
rect 2925 3510 2930 3545
rect 2820 3490 2930 3510
rect 2820 3455 2825 3490
rect 2925 3455 2930 3490
rect 2820 3430 2930 3455
rect 3070 3545 3180 3570
rect 3070 3510 3075 3545
rect 3175 3510 3180 3545
rect 3070 3490 3180 3510
rect 3070 3455 3075 3490
rect 3175 3455 3180 3490
rect 3070 3430 3180 3455
rect 3320 3545 3430 3570
rect 3320 3510 3325 3545
rect 3425 3510 3430 3545
rect 3320 3490 3430 3510
rect 3320 3455 3325 3490
rect 3425 3455 3430 3490
rect 3320 3430 3430 3455
rect 3570 3545 3680 3570
rect 3570 3510 3575 3545
rect 3675 3510 3680 3545
rect 3570 3490 3680 3510
rect 3570 3455 3575 3490
rect 3675 3455 3680 3490
rect 3570 3430 3680 3455
rect 3820 3545 3930 3570
rect 3820 3510 3825 3545
rect 3925 3510 3930 3545
rect 3820 3490 3930 3510
rect 3820 3455 3825 3490
rect 3925 3455 3930 3490
rect 3820 3430 3930 3455
rect 4070 3545 4180 3570
rect 4070 3510 4075 3545
rect 4175 3510 4180 3545
rect 4070 3490 4180 3510
rect 4070 3455 4075 3490
rect 4175 3455 4180 3490
rect 4070 3430 4180 3455
rect 4320 3545 4430 3570
rect 4320 3510 4325 3545
rect 4425 3510 4430 3545
rect 4320 3490 4430 3510
rect 4320 3455 4325 3490
rect 4425 3455 4430 3490
rect 4320 3430 4430 3455
rect 4570 3545 4680 3570
rect 4570 3510 4575 3545
rect 4675 3510 4680 3545
rect 4570 3490 4680 3510
rect 4570 3455 4575 3490
rect 4675 3455 4680 3490
rect 4570 3430 4680 3455
rect 4820 3545 4930 3570
rect 4820 3510 4825 3545
rect 4925 3510 4930 3545
rect 4820 3490 4930 3510
rect 4820 3455 4825 3490
rect 4925 3455 4930 3490
rect 4820 3430 4930 3455
rect 5070 3545 5180 3570
rect 5070 3510 5075 3545
rect 5175 3510 5180 3545
rect 5070 3490 5180 3510
rect 5070 3455 5075 3490
rect 5175 3455 5180 3490
rect 5070 3430 5180 3455
rect 5320 3545 5430 3570
rect 5320 3510 5325 3545
rect 5425 3510 5430 3545
rect 5320 3490 5430 3510
rect 5320 3455 5325 3490
rect 5425 3455 5430 3490
rect 5320 3430 5430 3455
rect 5570 3545 5680 3570
rect 5570 3510 5575 3545
rect 5675 3510 5680 3545
rect 5570 3490 5680 3510
rect 5570 3455 5575 3490
rect 5675 3455 5680 3490
rect 5570 3430 5680 3455
rect 5820 3545 5930 3570
rect 5820 3510 5825 3545
rect 5925 3510 5930 3545
rect 5820 3490 5930 3510
rect 5820 3455 5825 3490
rect 5925 3455 5930 3490
rect 5820 3430 5930 3455
rect 6070 3545 6180 3570
rect 6070 3510 6075 3545
rect 6175 3510 6180 3545
rect 6070 3490 6180 3510
rect 6070 3455 6075 3490
rect 6175 3455 6180 3490
rect 6070 3430 6180 3455
rect 6320 3545 6430 3570
rect 6320 3510 6325 3545
rect 6425 3510 6430 3545
rect 6320 3490 6430 3510
rect 6320 3455 6325 3490
rect 6425 3455 6430 3490
rect 6320 3430 6430 3455
rect 6570 3545 6680 3570
rect 6570 3510 6575 3545
rect 6675 3510 6680 3545
rect 6570 3490 6680 3510
rect 6570 3455 6575 3490
rect 6675 3455 6680 3490
rect 6570 3430 6680 3455
rect 6820 3545 6930 3570
rect 6820 3510 6825 3545
rect 6925 3510 6930 3545
rect 6820 3490 6930 3510
rect 6820 3455 6825 3490
rect 6925 3455 6930 3490
rect 6820 3430 6930 3455
rect 7070 3545 7180 3570
rect 7070 3510 7075 3545
rect 7175 3510 7180 3545
rect 7070 3490 7180 3510
rect 7070 3455 7075 3490
rect 7175 3455 7180 3490
rect 7070 3430 7180 3455
rect 7320 3545 7430 3570
rect 7320 3510 7325 3545
rect 7425 3510 7430 3545
rect 7320 3490 7430 3510
rect 7320 3455 7325 3490
rect 7425 3455 7430 3490
rect 7320 3430 7430 3455
rect 7570 3545 7680 3570
rect 7570 3510 7575 3545
rect 7675 3510 7680 3545
rect 7570 3490 7680 3510
rect 7570 3455 7575 3490
rect 7675 3455 7680 3490
rect 7570 3430 7680 3455
rect 7820 3545 7930 3570
rect 7820 3510 7825 3545
rect 7925 3510 7930 3545
rect 7820 3490 7930 3510
rect 7820 3455 7825 3490
rect 7925 3455 7930 3490
rect 7820 3430 7930 3455
rect 0 3425 8000 3430
rect 0 3325 10 3425
rect 45 3325 205 3425
rect 240 3325 260 3425
rect 295 3325 455 3425
rect 490 3325 510 3425
rect 545 3325 705 3425
rect 740 3325 760 3425
rect 795 3325 955 3425
rect 990 3325 1010 3425
rect 1045 3325 1205 3425
rect 1240 3325 1260 3425
rect 1295 3325 1455 3425
rect 1490 3325 1510 3425
rect 1545 3325 1705 3425
rect 1740 3325 1760 3425
rect 1795 3325 1955 3425
rect 1990 3325 2010 3425
rect 2045 3325 2205 3425
rect 2240 3325 2260 3425
rect 2295 3325 2455 3425
rect 2490 3325 2510 3425
rect 2545 3325 2705 3425
rect 2740 3325 2760 3425
rect 2795 3325 2955 3425
rect 2990 3325 3010 3425
rect 3045 3325 3205 3425
rect 3240 3325 3260 3425
rect 3295 3325 3455 3425
rect 3490 3325 3510 3425
rect 3545 3325 3705 3425
rect 3740 3325 3760 3425
rect 3795 3325 3955 3425
rect 3990 3325 4010 3425
rect 4045 3325 4205 3425
rect 4240 3325 4260 3425
rect 4295 3325 4455 3425
rect 4490 3325 4510 3425
rect 4545 3325 4705 3425
rect 4740 3325 4760 3425
rect 4795 3325 4955 3425
rect 4990 3325 5010 3425
rect 5045 3325 5205 3425
rect 5240 3325 5260 3425
rect 5295 3325 5455 3425
rect 5490 3325 5510 3425
rect 5545 3325 5705 3425
rect 5740 3325 5760 3425
rect 5795 3325 5955 3425
rect 5990 3325 6010 3425
rect 6045 3325 6205 3425
rect 6240 3325 6260 3425
rect 6295 3325 6455 3425
rect 6490 3325 6510 3425
rect 6545 3325 6705 3425
rect 6740 3325 6760 3425
rect 6795 3325 6955 3425
rect 6990 3325 7010 3425
rect 7045 3325 7205 3425
rect 7240 3325 7260 3425
rect 7295 3325 7455 3425
rect 7490 3325 7510 3425
rect 7545 3325 7705 3425
rect 7740 3325 7760 3425
rect 7795 3325 7955 3425
rect 7990 3325 8000 3425
rect 0 3320 8000 3325
rect 70 3295 180 3320
rect 70 3260 75 3295
rect 175 3260 180 3295
rect 70 3240 180 3260
rect 70 3205 75 3240
rect 175 3205 180 3240
rect 70 3180 180 3205
rect 320 3295 430 3320
rect 320 3260 325 3295
rect 425 3260 430 3295
rect 320 3240 430 3260
rect 320 3205 325 3240
rect 425 3205 430 3240
rect 320 3180 430 3205
rect 570 3295 680 3320
rect 570 3260 575 3295
rect 675 3260 680 3295
rect 570 3240 680 3260
rect 570 3205 575 3240
rect 675 3205 680 3240
rect 570 3180 680 3205
rect 820 3295 930 3320
rect 820 3260 825 3295
rect 925 3260 930 3295
rect 820 3240 930 3260
rect 820 3205 825 3240
rect 925 3205 930 3240
rect 820 3180 930 3205
rect 1070 3295 1180 3320
rect 1070 3260 1075 3295
rect 1175 3260 1180 3295
rect 1070 3240 1180 3260
rect 1070 3205 1075 3240
rect 1175 3205 1180 3240
rect 1070 3180 1180 3205
rect 1320 3295 1430 3320
rect 1320 3260 1325 3295
rect 1425 3260 1430 3295
rect 1320 3240 1430 3260
rect 1320 3205 1325 3240
rect 1425 3205 1430 3240
rect 1320 3180 1430 3205
rect 1570 3295 1680 3320
rect 1570 3260 1575 3295
rect 1675 3260 1680 3295
rect 1570 3240 1680 3260
rect 1570 3205 1575 3240
rect 1675 3205 1680 3240
rect 1570 3180 1680 3205
rect 1820 3295 1930 3320
rect 1820 3260 1825 3295
rect 1925 3260 1930 3295
rect 1820 3240 1930 3260
rect 1820 3205 1825 3240
rect 1925 3205 1930 3240
rect 1820 3180 1930 3205
rect 2070 3295 2180 3320
rect 2070 3260 2075 3295
rect 2175 3260 2180 3295
rect 2070 3240 2180 3260
rect 2070 3205 2075 3240
rect 2175 3205 2180 3240
rect 2070 3180 2180 3205
rect 2320 3295 2430 3320
rect 2320 3260 2325 3295
rect 2425 3260 2430 3295
rect 2320 3240 2430 3260
rect 2320 3205 2325 3240
rect 2425 3205 2430 3240
rect 2320 3180 2430 3205
rect 2570 3295 2680 3320
rect 2570 3260 2575 3295
rect 2675 3260 2680 3295
rect 2570 3240 2680 3260
rect 2570 3205 2575 3240
rect 2675 3205 2680 3240
rect 2570 3180 2680 3205
rect 2820 3295 2930 3320
rect 2820 3260 2825 3295
rect 2925 3260 2930 3295
rect 2820 3240 2930 3260
rect 2820 3205 2825 3240
rect 2925 3205 2930 3240
rect 2820 3180 2930 3205
rect 3070 3295 3180 3320
rect 3070 3260 3075 3295
rect 3175 3260 3180 3295
rect 3070 3240 3180 3260
rect 3070 3205 3075 3240
rect 3175 3205 3180 3240
rect 3070 3180 3180 3205
rect 3320 3295 3430 3320
rect 3320 3260 3325 3295
rect 3425 3260 3430 3295
rect 3320 3240 3430 3260
rect 3320 3205 3325 3240
rect 3425 3205 3430 3240
rect 3320 3180 3430 3205
rect 3570 3295 3680 3320
rect 3570 3260 3575 3295
rect 3675 3260 3680 3295
rect 3570 3240 3680 3260
rect 3570 3205 3575 3240
rect 3675 3205 3680 3240
rect 3570 3180 3680 3205
rect 3820 3295 3930 3320
rect 3820 3260 3825 3295
rect 3925 3260 3930 3295
rect 3820 3240 3930 3260
rect 3820 3205 3825 3240
rect 3925 3205 3930 3240
rect 3820 3180 3930 3205
rect 4070 3295 4180 3320
rect 4070 3260 4075 3295
rect 4175 3260 4180 3295
rect 4070 3240 4180 3260
rect 4070 3205 4075 3240
rect 4175 3205 4180 3240
rect 4070 3180 4180 3205
rect 4320 3295 4430 3320
rect 4320 3260 4325 3295
rect 4425 3260 4430 3295
rect 4320 3240 4430 3260
rect 4320 3205 4325 3240
rect 4425 3205 4430 3240
rect 4320 3180 4430 3205
rect 4570 3295 4680 3320
rect 4570 3260 4575 3295
rect 4675 3260 4680 3295
rect 4570 3240 4680 3260
rect 4570 3205 4575 3240
rect 4675 3205 4680 3240
rect 4570 3180 4680 3205
rect 4820 3295 4930 3320
rect 4820 3260 4825 3295
rect 4925 3260 4930 3295
rect 4820 3240 4930 3260
rect 4820 3205 4825 3240
rect 4925 3205 4930 3240
rect 4820 3180 4930 3205
rect 5070 3295 5180 3320
rect 5070 3260 5075 3295
rect 5175 3260 5180 3295
rect 5070 3240 5180 3260
rect 5070 3205 5075 3240
rect 5175 3205 5180 3240
rect 5070 3180 5180 3205
rect 5320 3295 5430 3320
rect 5320 3260 5325 3295
rect 5425 3260 5430 3295
rect 5320 3240 5430 3260
rect 5320 3205 5325 3240
rect 5425 3205 5430 3240
rect 5320 3180 5430 3205
rect 5570 3295 5680 3320
rect 5570 3260 5575 3295
rect 5675 3260 5680 3295
rect 5570 3240 5680 3260
rect 5570 3205 5575 3240
rect 5675 3205 5680 3240
rect 5570 3180 5680 3205
rect 5820 3295 5930 3320
rect 5820 3260 5825 3295
rect 5925 3260 5930 3295
rect 5820 3240 5930 3260
rect 5820 3205 5825 3240
rect 5925 3205 5930 3240
rect 5820 3180 5930 3205
rect 6070 3295 6180 3320
rect 6070 3260 6075 3295
rect 6175 3260 6180 3295
rect 6070 3240 6180 3260
rect 6070 3205 6075 3240
rect 6175 3205 6180 3240
rect 6070 3180 6180 3205
rect 6320 3295 6430 3320
rect 6320 3260 6325 3295
rect 6425 3260 6430 3295
rect 6320 3240 6430 3260
rect 6320 3205 6325 3240
rect 6425 3205 6430 3240
rect 6320 3180 6430 3205
rect 6570 3295 6680 3320
rect 6570 3260 6575 3295
rect 6675 3260 6680 3295
rect 6570 3240 6680 3260
rect 6570 3205 6575 3240
rect 6675 3205 6680 3240
rect 6570 3180 6680 3205
rect 6820 3295 6930 3320
rect 6820 3260 6825 3295
rect 6925 3260 6930 3295
rect 6820 3240 6930 3260
rect 6820 3205 6825 3240
rect 6925 3205 6930 3240
rect 6820 3180 6930 3205
rect 7070 3295 7180 3320
rect 7070 3260 7075 3295
rect 7175 3260 7180 3295
rect 7070 3240 7180 3260
rect 7070 3205 7075 3240
rect 7175 3205 7180 3240
rect 7070 3180 7180 3205
rect 7320 3295 7430 3320
rect 7320 3260 7325 3295
rect 7425 3260 7430 3295
rect 7320 3240 7430 3260
rect 7320 3205 7325 3240
rect 7425 3205 7430 3240
rect 7320 3180 7430 3205
rect 7570 3295 7680 3320
rect 7570 3260 7575 3295
rect 7675 3260 7680 3295
rect 7570 3240 7680 3260
rect 7570 3205 7575 3240
rect 7675 3205 7680 3240
rect 7570 3180 7680 3205
rect 7820 3295 7930 3320
rect 7820 3260 7825 3295
rect 7925 3260 7930 3295
rect 7820 3240 7930 3260
rect 7820 3205 7825 3240
rect 7925 3205 7930 3240
rect 7820 3180 7930 3205
rect 0 3175 8000 3180
rect 0 3075 10 3175
rect 45 3075 205 3175
rect 240 3075 260 3175
rect 295 3075 455 3175
rect 490 3075 510 3175
rect 545 3075 705 3175
rect 740 3075 760 3175
rect 795 3075 955 3175
rect 990 3075 1010 3175
rect 1045 3075 1205 3175
rect 1240 3075 1260 3175
rect 1295 3075 1455 3175
rect 1490 3075 1510 3175
rect 1545 3075 1705 3175
rect 1740 3075 1760 3175
rect 1795 3075 1955 3175
rect 1990 3075 2010 3175
rect 2045 3075 2205 3175
rect 2240 3075 2260 3175
rect 2295 3075 2455 3175
rect 2490 3075 2510 3175
rect 2545 3075 2705 3175
rect 2740 3075 2760 3175
rect 2795 3075 2955 3175
rect 2990 3075 3010 3175
rect 3045 3075 3205 3175
rect 3240 3075 3260 3175
rect 3295 3075 3455 3175
rect 3490 3075 3510 3175
rect 3545 3075 3705 3175
rect 3740 3075 3760 3175
rect 3795 3075 3955 3175
rect 3990 3075 4010 3175
rect 4045 3075 4205 3175
rect 4240 3075 4260 3175
rect 4295 3075 4455 3175
rect 4490 3075 4510 3175
rect 4545 3075 4705 3175
rect 4740 3075 4760 3175
rect 4795 3075 4955 3175
rect 4990 3075 5010 3175
rect 5045 3075 5205 3175
rect 5240 3075 5260 3175
rect 5295 3075 5455 3175
rect 5490 3075 5510 3175
rect 5545 3075 5705 3175
rect 5740 3075 5760 3175
rect 5795 3075 5955 3175
rect 5990 3075 6010 3175
rect 6045 3075 6205 3175
rect 6240 3075 6260 3175
rect 6295 3075 6455 3175
rect 6490 3075 6510 3175
rect 6545 3075 6705 3175
rect 6740 3075 6760 3175
rect 6795 3075 6955 3175
rect 6990 3075 7010 3175
rect 7045 3075 7205 3175
rect 7240 3075 7260 3175
rect 7295 3075 7455 3175
rect 7490 3075 7510 3175
rect 7545 3075 7705 3175
rect 7740 3075 7760 3175
rect 7795 3075 7955 3175
rect 7990 3075 8000 3175
rect 0 3070 8000 3075
rect 70 3045 180 3070
rect 70 3010 75 3045
rect 175 3010 180 3045
rect 70 2990 180 3010
rect 70 2955 75 2990
rect 175 2955 180 2990
rect 70 2930 180 2955
rect 320 3045 430 3070
rect 320 3010 325 3045
rect 425 3010 430 3045
rect 320 2990 430 3010
rect 320 2955 325 2990
rect 425 2955 430 2990
rect 320 2930 430 2955
rect 570 3045 680 3070
rect 570 3010 575 3045
rect 675 3010 680 3045
rect 570 2990 680 3010
rect 570 2955 575 2990
rect 675 2955 680 2990
rect 570 2930 680 2955
rect 820 3045 930 3070
rect 820 3010 825 3045
rect 925 3010 930 3045
rect 820 2990 930 3010
rect 820 2955 825 2990
rect 925 2955 930 2990
rect 820 2930 930 2955
rect 1070 3045 1180 3070
rect 1070 3010 1075 3045
rect 1175 3010 1180 3045
rect 1070 2990 1180 3010
rect 1070 2955 1075 2990
rect 1175 2955 1180 2990
rect 1070 2930 1180 2955
rect 1320 3045 1430 3070
rect 1320 3010 1325 3045
rect 1425 3010 1430 3045
rect 1320 2990 1430 3010
rect 1320 2955 1325 2990
rect 1425 2955 1430 2990
rect 1320 2930 1430 2955
rect 1570 3045 1680 3070
rect 1570 3010 1575 3045
rect 1675 3010 1680 3045
rect 1570 2990 1680 3010
rect 1570 2955 1575 2990
rect 1675 2955 1680 2990
rect 1570 2930 1680 2955
rect 1820 3045 1930 3070
rect 1820 3010 1825 3045
rect 1925 3010 1930 3045
rect 1820 2990 1930 3010
rect 1820 2955 1825 2990
rect 1925 2955 1930 2990
rect 1820 2930 1930 2955
rect 2070 3045 2180 3070
rect 2070 3010 2075 3045
rect 2175 3010 2180 3045
rect 2070 2990 2180 3010
rect 2070 2955 2075 2990
rect 2175 2955 2180 2990
rect 2070 2930 2180 2955
rect 2320 3045 2430 3070
rect 2320 3010 2325 3045
rect 2425 3010 2430 3045
rect 2320 2990 2430 3010
rect 2320 2955 2325 2990
rect 2425 2955 2430 2990
rect 2320 2930 2430 2955
rect 2570 3045 2680 3070
rect 2570 3010 2575 3045
rect 2675 3010 2680 3045
rect 2570 2990 2680 3010
rect 2570 2955 2575 2990
rect 2675 2955 2680 2990
rect 2570 2930 2680 2955
rect 2820 3045 2930 3070
rect 2820 3010 2825 3045
rect 2925 3010 2930 3045
rect 2820 2990 2930 3010
rect 2820 2955 2825 2990
rect 2925 2955 2930 2990
rect 2820 2930 2930 2955
rect 3070 3045 3180 3070
rect 3070 3010 3075 3045
rect 3175 3010 3180 3045
rect 3070 2990 3180 3010
rect 3070 2955 3075 2990
rect 3175 2955 3180 2990
rect 3070 2930 3180 2955
rect 3320 3045 3430 3070
rect 3320 3010 3325 3045
rect 3425 3010 3430 3045
rect 3320 2990 3430 3010
rect 3320 2955 3325 2990
rect 3425 2955 3430 2990
rect 3320 2930 3430 2955
rect 3570 3045 3680 3070
rect 3570 3010 3575 3045
rect 3675 3010 3680 3045
rect 3570 2990 3680 3010
rect 3570 2955 3575 2990
rect 3675 2955 3680 2990
rect 3570 2930 3680 2955
rect 3820 3045 3930 3070
rect 3820 3010 3825 3045
rect 3925 3010 3930 3045
rect 3820 2990 3930 3010
rect 3820 2955 3825 2990
rect 3925 2955 3930 2990
rect 3820 2930 3930 2955
rect 4070 3045 4180 3070
rect 4070 3010 4075 3045
rect 4175 3010 4180 3045
rect 4070 2990 4180 3010
rect 4070 2955 4075 2990
rect 4175 2955 4180 2990
rect 4070 2930 4180 2955
rect 4320 3045 4430 3070
rect 4320 3010 4325 3045
rect 4425 3010 4430 3045
rect 4320 2990 4430 3010
rect 4320 2955 4325 2990
rect 4425 2955 4430 2990
rect 4320 2930 4430 2955
rect 4570 3045 4680 3070
rect 4570 3010 4575 3045
rect 4675 3010 4680 3045
rect 4570 2990 4680 3010
rect 4570 2955 4575 2990
rect 4675 2955 4680 2990
rect 4570 2930 4680 2955
rect 4820 3045 4930 3070
rect 4820 3010 4825 3045
rect 4925 3010 4930 3045
rect 4820 2990 4930 3010
rect 4820 2955 4825 2990
rect 4925 2955 4930 2990
rect 4820 2930 4930 2955
rect 5070 3045 5180 3070
rect 5070 3010 5075 3045
rect 5175 3010 5180 3045
rect 5070 2990 5180 3010
rect 5070 2955 5075 2990
rect 5175 2955 5180 2990
rect 5070 2930 5180 2955
rect 5320 3045 5430 3070
rect 5320 3010 5325 3045
rect 5425 3010 5430 3045
rect 5320 2990 5430 3010
rect 5320 2955 5325 2990
rect 5425 2955 5430 2990
rect 5320 2930 5430 2955
rect 5570 3045 5680 3070
rect 5570 3010 5575 3045
rect 5675 3010 5680 3045
rect 5570 2990 5680 3010
rect 5570 2955 5575 2990
rect 5675 2955 5680 2990
rect 5570 2930 5680 2955
rect 5820 3045 5930 3070
rect 5820 3010 5825 3045
rect 5925 3010 5930 3045
rect 5820 2990 5930 3010
rect 5820 2955 5825 2990
rect 5925 2955 5930 2990
rect 5820 2930 5930 2955
rect 6070 3045 6180 3070
rect 6070 3010 6075 3045
rect 6175 3010 6180 3045
rect 6070 2990 6180 3010
rect 6070 2955 6075 2990
rect 6175 2955 6180 2990
rect 6070 2930 6180 2955
rect 6320 3045 6430 3070
rect 6320 3010 6325 3045
rect 6425 3010 6430 3045
rect 6320 2990 6430 3010
rect 6320 2955 6325 2990
rect 6425 2955 6430 2990
rect 6320 2930 6430 2955
rect 6570 3045 6680 3070
rect 6570 3010 6575 3045
rect 6675 3010 6680 3045
rect 6570 2990 6680 3010
rect 6570 2955 6575 2990
rect 6675 2955 6680 2990
rect 6570 2930 6680 2955
rect 6820 3045 6930 3070
rect 6820 3010 6825 3045
rect 6925 3010 6930 3045
rect 6820 2990 6930 3010
rect 6820 2955 6825 2990
rect 6925 2955 6930 2990
rect 6820 2930 6930 2955
rect 7070 3045 7180 3070
rect 7070 3010 7075 3045
rect 7175 3010 7180 3045
rect 7070 2990 7180 3010
rect 7070 2955 7075 2990
rect 7175 2955 7180 2990
rect 7070 2930 7180 2955
rect 7320 3045 7430 3070
rect 7320 3010 7325 3045
rect 7425 3010 7430 3045
rect 7320 2990 7430 3010
rect 7320 2955 7325 2990
rect 7425 2955 7430 2990
rect 7320 2930 7430 2955
rect 7570 3045 7680 3070
rect 7570 3010 7575 3045
rect 7675 3010 7680 3045
rect 7570 2990 7680 3010
rect 7570 2955 7575 2990
rect 7675 2955 7680 2990
rect 7570 2930 7680 2955
rect 7820 3045 7930 3070
rect 7820 3010 7825 3045
rect 7925 3010 7930 3045
rect 7820 2990 7930 3010
rect 7820 2955 7825 2990
rect 7925 2955 7930 2990
rect 7820 2930 7930 2955
rect 0 2925 8000 2930
rect 0 2825 10 2925
rect 45 2825 205 2925
rect 240 2825 260 2925
rect 295 2825 455 2925
rect 490 2825 510 2925
rect 545 2825 705 2925
rect 740 2825 760 2925
rect 795 2825 955 2925
rect 990 2825 1010 2925
rect 1045 2825 1205 2925
rect 1240 2825 1260 2925
rect 1295 2825 1455 2925
rect 1490 2825 1510 2925
rect 1545 2825 1705 2925
rect 1740 2825 1760 2925
rect 1795 2825 1955 2925
rect 1990 2825 2010 2925
rect 2045 2825 2205 2925
rect 2240 2825 2260 2925
rect 2295 2825 2455 2925
rect 2490 2825 2510 2925
rect 2545 2825 2705 2925
rect 2740 2825 2760 2925
rect 2795 2825 2955 2925
rect 2990 2825 3010 2925
rect 3045 2825 3205 2925
rect 3240 2825 3260 2925
rect 3295 2825 3455 2925
rect 3490 2825 3510 2925
rect 3545 2825 3705 2925
rect 3740 2825 3760 2925
rect 3795 2825 3955 2925
rect 3990 2825 4010 2925
rect 4045 2825 4205 2925
rect 4240 2825 4260 2925
rect 4295 2825 4455 2925
rect 4490 2825 4510 2925
rect 4545 2825 4705 2925
rect 4740 2825 4760 2925
rect 4795 2825 4955 2925
rect 4990 2825 5010 2925
rect 5045 2825 5205 2925
rect 5240 2825 5260 2925
rect 5295 2825 5455 2925
rect 5490 2825 5510 2925
rect 5545 2825 5705 2925
rect 5740 2825 5760 2925
rect 5795 2825 5955 2925
rect 5990 2825 6010 2925
rect 6045 2825 6205 2925
rect 6240 2825 6260 2925
rect 6295 2825 6455 2925
rect 6490 2825 6510 2925
rect 6545 2825 6705 2925
rect 6740 2825 6760 2925
rect 6795 2825 6955 2925
rect 6990 2825 7010 2925
rect 7045 2825 7205 2925
rect 7240 2825 7260 2925
rect 7295 2825 7455 2925
rect 7490 2825 7510 2925
rect 7545 2825 7705 2925
rect 7740 2825 7760 2925
rect 7795 2825 7955 2925
rect 7990 2825 8000 2925
rect 0 2820 8000 2825
rect 70 2795 180 2820
rect 70 2760 75 2795
rect 175 2760 180 2795
rect 70 2740 180 2760
rect 70 2705 75 2740
rect 175 2705 180 2740
rect 70 2680 180 2705
rect 320 2795 430 2820
rect 320 2760 325 2795
rect 425 2760 430 2795
rect 320 2740 430 2760
rect 320 2705 325 2740
rect 425 2705 430 2740
rect 320 2680 430 2705
rect 570 2795 680 2820
rect 570 2760 575 2795
rect 675 2760 680 2795
rect 570 2740 680 2760
rect 570 2705 575 2740
rect 675 2705 680 2740
rect 570 2680 680 2705
rect 820 2795 930 2820
rect 820 2760 825 2795
rect 925 2760 930 2795
rect 820 2740 930 2760
rect 820 2705 825 2740
rect 925 2705 930 2740
rect 820 2680 930 2705
rect 1070 2795 1180 2820
rect 1070 2760 1075 2795
rect 1175 2760 1180 2795
rect 1070 2740 1180 2760
rect 1070 2705 1075 2740
rect 1175 2705 1180 2740
rect 1070 2680 1180 2705
rect 1320 2795 1430 2820
rect 1320 2760 1325 2795
rect 1425 2760 1430 2795
rect 1320 2740 1430 2760
rect 1320 2705 1325 2740
rect 1425 2705 1430 2740
rect 1320 2680 1430 2705
rect 1570 2795 1680 2820
rect 1570 2760 1575 2795
rect 1675 2760 1680 2795
rect 1570 2740 1680 2760
rect 1570 2705 1575 2740
rect 1675 2705 1680 2740
rect 1570 2680 1680 2705
rect 1820 2795 1930 2820
rect 1820 2760 1825 2795
rect 1925 2760 1930 2795
rect 1820 2740 1930 2760
rect 1820 2705 1825 2740
rect 1925 2705 1930 2740
rect 1820 2680 1930 2705
rect 2070 2795 2180 2820
rect 2070 2760 2075 2795
rect 2175 2760 2180 2795
rect 2070 2740 2180 2760
rect 2070 2705 2075 2740
rect 2175 2705 2180 2740
rect 2070 2680 2180 2705
rect 2320 2795 2430 2820
rect 2320 2760 2325 2795
rect 2425 2760 2430 2795
rect 2320 2740 2430 2760
rect 2320 2705 2325 2740
rect 2425 2705 2430 2740
rect 2320 2680 2430 2705
rect 2570 2795 2680 2820
rect 2570 2760 2575 2795
rect 2675 2760 2680 2795
rect 2570 2740 2680 2760
rect 2570 2705 2575 2740
rect 2675 2705 2680 2740
rect 2570 2680 2680 2705
rect 2820 2795 2930 2820
rect 2820 2760 2825 2795
rect 2925 2760 2930 2795
rect 2820 2740 2930 2760
rect 2820 2705 2825 2740
rect 2925 2705 2930 2740
rect 2820 2680 2930 2705
rect 3070 2795 3180 2820
rect 3070 2760 3075 2795
rect 3175 2760 3180 2795
rect 3070 2740 3180 2760
rect 3070 2705 3075 2740
rect 3175 2705 3180 2740
rect 3070 2680 3180 2705
rect 3320 2795 3430 2820
rect 3320 2760 3325 2795
rect 3425 2760 3430 2795
rect 3320 2740 3430 2760
rect 3320 2705 3325 2740
rect 3425 2705 3430 2740
rect 3320 2680 3430 2705
rect 3570 2795 3680 2820
rect 3570 2760 3575 2795
rect 3675 2760 3680 2795
rect 3570 2740 3680 2760
rect 3570 2705 3575 2740
rect 3675 2705 3680 2740
rect 3570 2680 3680 2705
rect 3820 2795 3930 2820
rect 3820 2760 3825 2795
rect 3925 2760 3930 2795
rect 3820 2740 3930 2760
rect 3820 2705 3825 2740
rect 3925 2705 3930 2740
rect 3820 2680 3930 2705
rect 4070 2795 4180 2820
rect 4070 2760 4075 2795
rect 4175 2760 4180 2795
rect 4070 2740 4180 2760
rect 4070 2705 4075 2740
rect 4175 2705 4180 2740
rect 4070 2680 4180 2705
rect 4320 2795 4430 2820
rect 4320 2760 4325 2795
rect 4425 2760 4430 2795
rect 4320 2740 4430 2760
rect 4320 2705 4325 2740
rect 4425 2705 4430 2740
rect 4320 2680 4430 2705
rect 4570 2795 4680 2820
rect 4570 2760 4575 2795
rect 4675 2760 4680 2795
rect 4570 2740 4680 2760
rect 4570 2705 4575 2740
rect 4675 2705 4680 2740
rect 4570 2680 4680 2705
rect 4820 2795 4930 2820
rect 4820 2760 4825 2795
rect 4925 2760 4930 2795
rect 4820 2740 4930 2760
rect 4820 2705 4825 2740
rect 4925 2705 4930 2740
rect 4820 2680 4930 2705
rect 5070 2795 5180 2820
rect 5070 2760 5075 2795
rect 5175 2760 5180 2795
rect 5070 2740 5180 2760
rect 5070 2705 5075 2740
rect 5175 2705 5180 2740
rect 5070 2680 5180 2705
rect 5320 2795 5430 2820
rect 5320 2760 5325 2795
rect 5425 2760 5430 2795
rect 5320 2740 5430 2760
rect 5320 2705 5325 2740
rect 5425 2705 5430 2740
rect 5320 2680 5430 2705
rect 5570 2795 5680 2820
rect 5570 2760 5575 2795
rect 5675 2760 5680 2795
rect 5570 2740 5680 2760
rect 5570 2705 5575 2740
rect 5675 2705 5680 2740
rect 5570 2680 5680 2705
rect 5820 2795 5930 2820
rect 5820 2760 5825 2795
rect 5925 2760 5930 2795
rect 5820 2740 5930 2760
rect 5820 2705 5825 2740
rect 5925 2705 5930 2740
rect 5820 2680 5930 2705
rect 6070 2795 6180 2820
rect 6070 2760 6075 2795
rect 6175 2760 6180 2795
rect 6070 2740 6180 2760
rect 6070 2705 6075 2740
rect 6175 2705 6180 2740
rect 6070 2680 6180 2705
rect 6320 2795 6430 2820
rect 6320 2760 6325 2795
rect 6425 2760 6430 2795
rect 6320 2740 6430 2760
rect 6320 2705 6325 2740
rect 6425 2705 6430 2740
rect 6320 2680 6430 2705
rect 6570 2795 6680 2820
rect 6570 2760 6575 2795
rect 6675 2760 6680 2795
rect 6570 2740 6680 2760
rect 6570 2705 6575 2740
rect 6675 2705 6680 2740
rect 6570 2680 6680 2705
rect 6820 2795 6930 2820
rect 6820 2760 6825 2795
rect 6925 2760 6930 2795
rect 6820 2740 6930 2760
rect 6820 2705 6825 2740
rect 6925 2705 6930 2740
rect 6820 2680 6930 2705
rect 7070 2795 7180 2820
rect 7070 2760 7075 2795
rect 7175 2760 7180 2795
rect 7070 2740 7180 2760
rect 7070 2705 7075 2740
rect 7175 2705 7180 2740
rect 7070 2680 7180 2705
rect 7320 2795 7430 2820
rect 7320 2760 7325 2795
rect 7425 2760 7430 2795
rect 7320 2740 7430 2760
rect 7320 2705 7325 2740
rect 7425 2705 7430 2740
rect 7320 2680 7430 2705
rect 7570 2795 7680 2820
rect 7570 2760 7575 2795
rect 7675 2760 7680 2795
rect 7570 2740 7680 2760
rect 7570 2705 7575 2740
rect 7675 2705 7680 2740
rect 7570 2680 7680 2705
rect 7820 2795 7930 2820
rect 7820 2760 7825 2795
rect 7925 2760 7930 2795
rect 7820 2740 7930 2760
rect 7820 2705 7825 2740
rect 7925 2705 7930 2740
rect 7820 2680 7930 2705
rect 0 2675 8000 2680
rect 0 2575 10 2675
rect 45 2575 205 2675
rect 240 2575 260 2675
rect 295 2575 455 2675
rect 490 2575 510 2675
rect 545 2575 705 2675
rect 740 2575 760 2675
rect 795 2575 955 2675
rect 990 2575 1010 2675
rect 1045 2575 1205 2675
rect 1240 2575 1260 2675
rect 1295 2575 1455 2675
rect 1490 2575 1510 2675
rect 1545 2575 1705 2675
rect 1740 2575 1760 2675
rect 1795 2575 1955 2675
rect 1990 2575 2010 2675
rect 2045 2575 2205 2675
rect 2240 2575 2260 2675
rect 2295 2575 2455 2675
rect 2490 2575 2510 2675
rect 2545 2575 2705 2675
rect 2740 2575 2760 2675
rect 2795 2575 2955 2675
rect 2990 2575 3010 2675
rect 3045 2575 3205 2675
rect 3240 2575 3260 2675
rect 3295 2575 3455 2675
rect 3490 2575 3510 2675
rect 3545 2575 3705 2675
rect 3740 2575 3760 2675
rect 3795 2575 3955 2675
rect 3990 2575 4010 2675
rect 4045 2575 4205 2675
rect 4240 2575 4260 2675
rect 4295 2575 4455 2675
rect 4490 2575 4510 2675
rect 4545 2575 4705 2675
rect 4740 2575 4760 2675
rect 4795 2575 4955 2675
rect 4990 2575 5010 2675
rect 5045 2575 5205 2675
rect 5240 2575 5260 2675
rect 5295 2575 5455 2675
rect 5490 2575 5510 2675
rect 5545 2575 5705 2675
rect 5740 2575 5760 2675
rect 5795 2575 5955 2675
rect 5990 2575 6010 2675
rect 6045 2575 6205 2675
rect 6240 2575 6260 2675
rect 6295 2575 6455 2675
rect 6490 2575 6510 2675
rect 6545 2575 6705 2675
rect 6740 2575 6760 2675
rect 6795 2575 6955 2675
rect 6990 2575 7010 2675
rect 7045 2575 7205 2675
rect 7240 2575 7260 2675
rect 7295 2575 7455 2675
rect 7490 2575 7510 2675
rect 7545 2575 7705 2675
rect 7740 2575 7760 2675
rect 7795 2575 7955 2675
rect 7990 2575 8000 2675
rect 0 2570 8000 2575
rect 70 2545 180 2570
rect 70 2510 75 2545
rect 175 2510 180 2545
rect 70 2490 180 2510
rect 70 2455 75 2490
rect 175 2455 180 2490
rect 70 2430 180 2455
rect 320 2545 430 2570
rect 320 2510 325 2545
rect 425 2510 430 2545
rect 320 2490 430 2510
rect 320 2455 325 2490
rect 425 2455 430 2490
rect 320 2430 430 2455
rect 570 2545 680 2570
rect 570 2510 575 2545
rect 675 2510 680 2545
rect 570 2490 680 2510
rect 570 2455 575 2490
rect 675 2455 680 2490
rect 570 2430 680 2455
rect 820 2545 930 2570
rect 820 2510 825 2545
rect 925 2510 930 2545
rect 820 2490 930 2510
rect 820 2455 825 2490
rect 925 2455 930 2490
rect 820 2430 930 2455
rect 1070 2545 1180 2570
rect 1070 2510 1075 2545
rect 1175 2510 1180 2545
rect 1070 2490 1180 2510
rect 1070 2455 1075 2490
rect 1175 2455 1180 2490
rect 1070 2430 1180 2455
rect 1320 2545 1430 2570
rect 1320 2510 1325 2545
rect 1425 2510 1430 2545
rect 1320 2490 1430 2510
rect 1320 2455 1325 2490
rect 1425 2455 1430 2490
rect 1320 2430 1430 2455
rect 1570 2545 1680 2570
rect 1570 2510 1575 2545
rect 1675 2510 1680 2545
rect 1570 2490 1680 2510
rect 1570 2455 1575 2490
rect 1675 2455 1680 2490
rect 1570 2430 1680 2455
rect 1820 2545 1930 2570
rect 1820 2510 1825 2545
rect 1925 2510 1930 2545
rect 1820 2490 1930 2510
rect 1820 2455 1825 2490
rect 1925 2455 1930 2490
rect 1820 2430 1930 2455
rect 2070 2545 2180 2570
rect 2070 2510 2075 2545
rect 2175 2510 2180 2545
rect 2070 2490 2180 2510
rect 2070 2455 2075 2490
rect 2175 2455 2180 2490
rect 2070 2430 2180 2455
rect 2320 2545 2430 2570
rect 2320 2510 2325 2545
rect 2425 2510 2430 2545
rect 2320 2490 2430 2510
rect 2320 2455 2325 2490
rect 2425 2455 2430 2490
rect 2320 2430 2430 2455
rect 2570 2545 2680 2570
rect 2570 2510 2575 2545
rect 2675 2510 2680 2545
rect 2570 2490 2680 2510
rect 2570 2455 2575 2490
rect 2675 2455 2680 2490
rect 2570 2430 2680 2455
rect 2820 2545 2930 2570
rect 2820 2510 2825 2545
rect 2925 2510 2930 2545
rect 2820 2490 2930 2510
rect 2820 2455 2825 2490
rect 2925 2455 2930 2490
rect 2820 2430 2930 2455
rect 3070 2545 3180 2570
rect 3070 2510 3075 2545
rect 3175 2510 3180 2545
rect 3070 2490 3180 2510
rect 3070 2455 3075 2490
rect 3175 2455 3180 2490
rect 3070 2430 3180 2455
rect 3320 2545 3430 2570
rect 3320 2510 3325 2545
rect 3425 2510 3430 2545
rect 3320 2490 3430 2510
rect 3320 2455 3325 2490
rect 3425 2455 3430 2490
rect 3320 2430 3430 2455
rect 3570 2545 3680 2570
rect 3570 2510 3575 2545
rect 3675 2510 3680 2545
rect 3570 2490 3680 2510
rect 3570 2455 3575 2490
rect 3675 2455 3680 2490
rect 3570 2430 3680 2455
rect 3820 2545 3930 2570
rect 3820 2510 3825 2545
rect 3925 2510 3930 2545
rect 3820 2490 3930 2510
rect 3820 2455 3825 2490
rect 3925 2455 3930 2490
rect 3820 2430 3930 2455
rect 4070 2545 4180 2570
rect 4070 2510 4075 2545
rect 4175 2510 4180 2545
rect 4070 2490 4180 2510
rect 4070 2455 4075 2490
rect 4175 2455 4180 2490
rect 4070 2430 4180 2455
rect 4320 2545 4430 2570
rect 4320 2510 4325 2545
rect 4425 2510 4430 2545
rect 4320 2490 4430 2510
rect 4320 2455 4325 2490
rect 4425 2455 4430 2490
rect 4320 2430 4430 2455
rect 4570 2545 4680 2570
rect 4570 2510 4575 2545
rect 4675 2510 4680 2545
rect 4570 2490 4680 2510
rect 4570 2455 4575 2490
rect 4675 2455 4680 2490
rect 4570 2430 4680 2455
rect 4820 2545 4930 2570
rect 4820 2510 4825 2545
rect 4925 2510 4930 2545
rect 4820 2490 4930 2510
rect 4820 2455 4825 2490
rect 4925 2455 4930 2490
rect 4820 2430 4930 2455
rect 5070 2545 5180 2570
rect 5070 2510 5075 2545
rect 5175 2510 5180 2545
rect 5070 2490 5180 2510
rect 5070 2455 5075 2490
rect 5175 2455 5180 2490
rect 5070 2430 5180 2455
rect 5320 2545 5430 2570
rect 5320 2510 5325 2545
rect 5425 2510 5430 2545
rect 5320 2490 5430 2510
rect 5320 2455 5325 2490
rect 5425 2455 5430 2490
rect 5320 2430 5430 2455
rect 5570 2545 5680 2570
rect 5570 2510 5575 2545
rect 5675 2510 5680 2545
rect 5570 2490 5680 2510
rect 5570 2455 5575 2490
rect 5675 2455 5680 2490
rect 5570 2430 5680 2455
rect 5820 2545 5930 2570
rect 5820 2510 5825 2545
rect 5925 2510 5930 2545
rect 5820 2490 5930 2510
rect 5820 2455 5825 2490
rect 5925 2455 5930 2490
rect 5820 2430 5930 2455
rect 6070 2545 6180 2570
rect 6070 2510 6075 2545
rect 6175 2510 6180 2545
rect 6070 2490 6180 2510
rect 6070 2455 6075 2490
rect 6175 2455 6180 2490
rect 6070 2430 6180 2455
rect 6320 2545 6430 2570
rect 6320 2510 6325 2545
rect 6425 2510 6430 2545
rect 6320 2490 6430 2510
rect 6320 2455 6325 2490
rect 6425 2455 6430 2490
rect 6320 2430 6430 2455
rect 6570 2545 6680 2570
rect 6570 2510 6575 2545
rect 6675 2510 6680 2545
rect 6570 2490 6680 2510
rect 6570 2455 6575 2490
rect 6675 2455 6680 2490
rect 6570 2430 6680 2455
rect 6820 2545 6930 2570
rect 6820 2510 6825 2545
rect 6925 2510 6930 2545
rect 6820 2490 6930 2510
rect 6820 2455 6825 2490
rect 6925 2455 6930 2490
rect 6820 2430 6930 2455
rect 7070 2545 7180 2570
rect 7070 2510 7075 2545
rect 7175 2510 7180 2545
rect 7070 2490 7180 2510
rect 7070 2455 7075 2490
rect 7175 2455 7180 2490
rect 7070 2430 7180 2455
rect 7320 2545 7430 2570
rect 7320 2510 7325 2545
rect 7425 2510 7430 2545
rect 7320 2490 7430 2510
rect 7320 2455 7325 2490
rect 7425 2455 7430 2490
rect 7320 2430 7430 2455
rect 7570 2545 7680 2570
rect 7570 2510 7575 2545
rect 7675 2510 7680 2545
rect 7570 2490 7680 2510
rect 7570 2455 7575 2490
rect 7675 2455 7680 2490
rect 7570 2430 7680 2455
rect 7820 2545 7930 2570
rect 7820 2510 7825 2545
rect 7925 2510 7930 2545
rect 7820 2490 7930 2510
rect 7820 2455 7825 2490
rect 7925 2455 7930 2490
rect 7820 2430 7930 2455
rect 0 2425 8000 2430
rect 0 2325 10 2425
rect 45 2325 205 2425
rect 240 2325 260 2425
rect 295 2325 455 2425
rect 490 2325 510 2425
rect 545 2325 705 2425
rect 740 2325 760 2425
rect 795 2325 955 2425
rect 990 2325 1010 2425
rect 1045 2325 1205 2425
rect 1240 2325 1260 2425
rect 1295 2325 1455 2425
rect 1490 2325 1510 2425
rect 1545 2325 1705 2425
rect 1740 2325 1760 2425
rect 1795 2325 1955 2425
rect 1990 2325 2010 2425
rect 2045 2325 2205 2425
rect 2240 2325 2260 2425
rect 2295 2325 2455 2425
rect 2490 2325 2510 2425
rect 2545 2325 2705 2425
rect 2740 2325 2760 2425
rect 2795 2325 2955 2425
rect 2990 2325 3010 2425
rect 3045 2325 3205 2425
rect 3240 2325 3260 2425
rect 3295 2325 3455 2425
rect 3490 2325 3510 2425
rect 3545 2325 3705 2425
rect 3740 2325 3760 2425
rect 3795 2325 3955 2425
rect 3990 2325 4010 2425
rect 4045 2325 4205 2425
rect 4240 2325 4260 2425
rect 4295 2325 4455 2425
rect 4490 2325 4510 2425
rect 4545 2325 4705 2425
rect 4740 2325 4760 2425
rect 4795 2325 4955 2425
rect 4990 2325 5010 2425
rect 5045 2325 5205 2425
rect 5240 2325 5260 2425
rect 5295 2325 5455 2425
rect 5490 2325 5510 2425
rect 5545 2325 5705 2425
rect 5740 2325 5760 2425
rect 5795 2325 5955 2425
rect 5990 2325 6010 2425
rect 6045 2325 6205 2425
rect 6240 2325 6260 2425
rect 6295 2325 6455 2425
rect 6490 2325 6510 2425
rect 6545 2325 6705 2425
rect 6740 2325 6760 2425
rect 6795 2325 6955 2425
rect 6990 2325 7010 2425
rect 7045 2325 7205 2425
rect 7240 2325 7260 2425
rect 7295 2325 7455 2425
rect 7490 2325 7510 2425
rect 7545 2325 7705 2425
rect 7740 2325 7760 2425
rect 7795 2325 7955 2425
rect 7990 2325 8000 2425
rect 0 2320 8000 2325
rect 70 2295 180 2320
rect 70 2260 75 2295
rect 175 2260 180 2295
rect 70 2240 180 2260
rect 70 2205 75 2240
rect 175 2205 180 2240
rect 70 2180 180 2205
rect 320 2295 430 2320
rect 320 2260 325 2295
rect 425 2260 430 2295
rect 320 2240 430 2260
rect 320 2205 325 2240
rect 425 2205 430 2240
rect 320 2180 430 2205
rect 570 2295 680 2320
rect 570 2260 575 2295
rect 675 2260 680 2295
rect 570 2240 680 2260
rect 570 2205 575 2240
rect 675 2205 680 2240
rect 570 2180 680 2205
rect 820 2295 930 2320
rect 820 2260 825 2295
rect 925 2260 930 2295
rect 820 2240 930 2260
rect 820 2205 825 2240
rect 925 2205 930 2240
rect 820 2180 930 2205
rect 1070 2295 1180 2320
rect 1070 2260 1075 2295
rect 1175 2260 1180 2295
rect 1070 2240 1180 2260
rect 1070 2205 1075 2240
rect 1175 2205 1180 2240
rect 1070 2180 1180 2205
rect 1320 2295 1430 2320
rect 1320 2260 1325 2295
rect 1425 2260 1430 2295
rect 1320 2240 1430 2260
rect 1320 2205 1325 2240
rect 1425 2205 1430 2240
rect 1320 2180 1430 2205
rect 1570 2295 1680 2320
rect 1570 2260 1575 2295
rect 1675 2260 1680 2295
rect 1570 2240 1680 2260
rect 1570 2205 1575 2240
rect 1675 2205 1680 2240
rect 1570 2180 1680 2205
rect 1820 2295 1930 2320
rect 1820 2260 1825 2295
rect 1925 2260 1930 2295
rect 1820 2240 1930 2260
rect 1820 2205 1825 2240
rect 1925 2205 1930 2240
rect 1820 2180 1930 2205
rect 2070 2295 2180 2320
rect 2070 2260 2075 2295
rect 2175 2260 2180 2295
rect 2070 2240 2180 2260
rect 2070 2205 2075 2240
rect 2175 2205 2180 2240
rect 2070 2180 2180 2205
rect 2320 2295 2430 2320
rect 2320 2260 2325 2295
rect 2425 2260 2430 2295
rect 2320 2240 2430 2260
rect 2320 2205 2325 2240
rect 2425 2205 2430 2240
rect 2320 2180 2430 2205
rect 2570 2295 2680 2320
rect 2570 2260 2575 2295
rect 2675 2260 2680 2295
rect 2570 2240 2680 2260
rect 2570 2205 2575 2240
rect 2675 2205 2680 2240
rect 2570 2180 2680 2205
rect 2820 2295 2930 2320
rect 2820 2260 2825 2295
rect 2925 2260 2930 2295
rect 2820 2240 2930 2260
rect 2820 2205 2825 2240
rect 2925 2205 2930 2240
rect 2820 2180 2930 2205
rect 3070 2295 3180 2320
rect 3070 2260 3075 2295
rect 3175 2260 3180 2295
rect 3070 2240 3180 2260
rect 3070 2205 3075 2240
rect 3175 2205 3180 2240
rect 3070 2180 3180 2205
rect 3320 2295 3430 2320
rect 3320 2260 3325 2295
rect 3425 2260 3430 2295
rect 3320 2240 3430 2260
rect 3320 2205 3325 2240
rect 3425 2205 3430 2240
rect 3320 2180 3430 2205
rect 3570 2295 3680 2320
rect 3570 2260 3575 2295
rect 3675 2260 3680 2295
rect 3570 2240 3680 2260
rect 3570 2205 3575 2240
rect 3675 2205 3680 2240
rect 3570 2180 3680 2205
rect 3820 2295 3930 2320
rect 3820 2260 3825 2295
rect 3925 2260 3930 2295
rect 3820 2240 3930 2260
rect 3820 2205 3825 2240
rect 3925 2205 3930 2240
rect 3820 2180 3930 2205
rect 4070 2295 4180 2320
rect 4070 2260 4075 2295
rect 4175 2260 4180 2295
rect 4070 2240 4180 2260
rect 4070 2205 4075 2240
rect 4175 2205 4180 2240
rect 4070 2180 4180 2205
rect 4320 2295 4430 2320
rect 4320 2260 4325 2295
rect 4425 2260 4430 2295
rect 4320 2240 4430 2260
rect 4320 2205 4325 2240
rect 4425 2205 4430 2240
rect 4320 2180 4430 2205
rect 4570 2295 4680 2320
rect 4570 2260 4575 2295
rect 4675 2260 4680 2295
rect 4570 2240 4680 2260
rect 4570 2205 4575 2240
rect 4675 2205 4680 2240
rect 4570 2180 4680 2205
rect 4820 2295 4930 2320
rect 4820 2260 4825 2295
rect 4925 2260 4930 2295
rect 4820 2240 4930 2260
rect 4820 2205 4825 2240
rect 4925 2205 4930 2240
rect 4820 2180 4930 2205
rect 5070 2295 5180 2320
rect 5070 2260 5075 2295
rect 5175 2260 5180 2295
rect 5070 2240 5180 2260
rect 5070 2205 5075 2240
rect 5175 2205 5180 2240
rect 5070 2180 5180 2205
rect 5320 2295 5430 2320
rect 5320 2260 5325 2295
rect 5425 2260 5430 2295
rect 5320 2240 5430 2260
rect 5320 2205 5325 2240
rect 5425 2205 5430 2240
rect 5320 2180 5430 2205
rect 5570 2295 5680 2320
rect 5570 2260 5575 2295
rect 5675 2260 5680 2295
rect 5570 2240 5680 2260
rect 5570 2205 5575 2240
rect 5675 2205 5680 2240
rect 5570 2180 5680 2205
rect 5820 2295 5930 2320
rect 5820 2260 5825 2295
rect 5925 2260 5930 2295
rect 5820 2240 5930 2260
rect 5820 2205 5825 2240
rect 5925 2205 5930 2240
rect 5820 2180 5930 2205
rect 6070 2295 6180 2320
rect 6070 2260 6075 2295
rect 6175 2260 6180 2295
rect 6070 2240 6180 2260
rect 6070 2205 6075 2240
rect 6175 2205 6180 2240
rect 6070 2180 6180 2205
rect 6320 2295 6430 2320
rect 6320 2260 6325 2295
rect 6425 2260 6430 2295
rect 6320 2240 6430 2260
rect 6320 2205 6325 2240
rect 6425 2205 6430 2240
rect 6320 2180 6430 2205
rect 6570 2295 6680 2320
rect 6570 2260 6575 2295
rect 6675 2260 6680 2295
rect 6570 2240 6680 2260
rect 6570 2205 6575 2240
rect 6675 2205 6680 2240
rect 6570 2180 6680 2205
rect 6820 2295 6930 2320
rect 6820 2260 6825 2295
rect 6925 2260 6930 2295
rect 6820 2240 6930 2260
rect 6820 2205 6825 2240
rect 6925 2205 6930 2240
rect 6820 2180 6930 2205
rect 7070 2295 7180 2320
rect 7070 2260 7075 2295
rect 7175 2260 7180 2295
rect 7070 2240 7180 2260
rect 7070 2205 7075 2240
rect 7175 2205 7180 2240
rect 7070 2180 7180 2205
rect 7320 2295 7430 2320
rect 7320 2260 7325 2295
rect 7425 2260 7430 2295
rect 7320 2240 7430 2260
rect 7320 2205 7325 2240
rect 7425 2205 7430 2240
rect 7320 2180 7430 2205
rect 7570 2295 7680 2320
rect 7570 2260 7575 2295
rect 7675 2260 7680 2295
rect 7570 2240 7680 2260
rect 7570 2205 7575 2240
rect 7675 2205 7680 2240
rect 7570 2180 7680 2205
rect 7820 2295 7930 2320
rect 7820 2260 7825 2295
rect 7925 2260 7930 2295
rect 7820 2240 7930 2260
rect 7820 2205 7825 2240
rect 7925 2205 7930 2240
rect 7820 2180 7930 2205
rect 0 2175 8000 2180
rect 0 2075 10 2175
rect 45 2075 205 2175
rect 240 2075 260 2175
rect 295 2075 455 2175
rect 490 2075 510 2175
rect 545 2075 705 2175
rect 740 2075 760 2175
rect 795 2075 955 2175
rect 990 2075 1010 2175
rect 1045 2075 1205 2175
rect 1240 2075 1260 2175
rect 1295 2075 1455 2175
rect 1490 2075 1510 2175
rect 1545 2075 1705 2175
rect 1740 2075 1760 2175
rect 1795 2075 1955 2175
rect 1990 2075 2010 2175
rect 2045 2075 2205 2175
rect 2240 2075 2260 2175
rect 2295 2075 2455 2175
rect 2490 2075 2510 2175
rect 2545 2075 2705 2175
rect 2740 2075 2760 2175
rect 2795 2075 2955 2175
rect 2990 2075 3010 2175
rect 3045 2075 3205 2175
rect 3240 2075 3260 2175
rect 3295 2075 3455 2175
rect 3490 2075 3510 2175
rect 3545 2075 3705 2175
rect 3740 2075 3760 2175
rect 3795 2075 3955 2175
rect 3990 2075 4010 2175
rect 4045 2075 4205 2175
rect 4240 2075 4260 2175
rect 4295 2075 4455 2175
rect 4490 2075 4510 2175
rect 4545 2075 4705 2175
rect 4740 2075 4760 2175
rect 4795 2075 4955 2175
rect 4990 2075 5010 2175
rect 5045 2075 5205 2175
rect 5240 2075 5260 2175
rect 5295 2075 5455 2175
rect 5490 2075 5510 2175
rect 5545 2075 5705 2175
rect 5740 2075 5760 2175
rect 5795 2075 5955 2175
rect 5990 2075 6010 2175
rect 6045 2075 6205 2175
rect 6240 2075 6260 2175
rect 6295 2075 6455 2175
rect 6490 2075 6510 2175
rect 6545 2075 6705 2175
rect 6740 2075 6760 2175
rect 6795 2075 6955 2175
rect 6990 2075 7010 2175
rect 7045 2075 7205 2175
rect 7240 2075 7260 2175
rect 7295 2075 7455 2175
rect 7490 2075 7510 2175
rect 7545 2075 7705 2175
rect 7740 2075 7760 2175
rect 7795 2075 7955 2175
rect 7990 2075 8000 2175
rect 0 2070 8000 2075
rect 70 2045 180 2070
rect 70 2010 75 2045
rect 175 2010 180 2045
rect 70 1990 180 2010
rect 70 1955 75 1990
rect 175 1955 180 1990
rect 70 1930 180 1955
rect 320 2045 430 2070
rect 320 2010 325 2045
rect 425 2010 430 2045
rect 320 1990 430 2010
rect 320 1955 325 1990
rect 425 1955 430 1990
rect 320 1930 430 1955
rect 570 2045 680 2070
rect 570 2010 575 2045
rect 675 2010 680 2045
rect 570 1990 680 2010
rect 570 1955 575 1990
rect 675 1955 680 1990
rect 570 1930 680 1955
rect 820 2045 930 2070
rect 820 2010 825 2045
rect 925 2010 930 2045
rect 820 1990 930 2010
rect 820 1955 825 1990
rect 925 1955 930 1990
rect 820 1930 930 1955
rect 1070 2045 1180 2070
rect 1070 2010 1075 2045
rect 1175 2010 1180 2045
rect 1070 1990 1180 2010
rect 1070 1955 1075 1990
rect 1175 1955 1180 1990
rect 1070 1930 1180 1955
rect 1320 2045 1430 2070
rect 1320 2010 1325 2045
rect 1425 2010 1430 2045
rect 1320 1990 1430 2010
rect 1320 1955 1325 1990
rect 1425 1955 1430 1990
rect 1320 1930 1430 1955
rect 1570 2045 1680 2070
rect 1570 2010 1575 2045
rect 1675 2010 1680 2045
rect 1570 1990 1680 2010
rect 1570 1955 1575 1990
rect 1675 1955 1680 1990
rect 1570 1930 1680 1955
rect 1820 2045 1930 2070
rect 1820 2010 1825 2045
rect 1925 2010 1930 2045
rect 1820 1990 1930 2010
rect 1820 1955 1825 1990
rect 1925 1955 1930 1990
rect 1820 1930 1930 1955
rect 2070 2045 2180 2070
rect 2070 2010 2075 2045
rect 2175 2010 2180 2045
rect 2070 1990 2180 2010
rect 2070 1955 2075 1990
rect 2175 1955 2180 1990
rect 2070 1930 2180 1955
rect 2320 2045 2430 2070
rect 2320 2010 2325 2045
rect 2425 2010 2430 2045
rect 2320 1990 2430 2010
rect 2320 1955 2325 1990
rect 2425 1955 2430 1990
rect 2320 1930 2430 1955
rect 2570 2045 2680 2070
rect 2570 2010 2575 2045
rect 2675 2010 2680 2045
rect 2570 1990 2680 2010
rect 2570 1955 2575 1990
rect 2675 1955 2680 1990
rect 2570 1930 2680 1955
rect 2820 2045 2930 2070
rect 2820 2010 2825 2045
rect 2925 2010 2930 2045
rect 2820 1990 2930 2010
rect 2820 1955 2825 1990
rect 2925 1955 2930 1990
rect 2820 1930 2930 1955
rect 3070 2045 3180 2070
rect 3070 2010 3075 2045
rect 3175 2010 3180 2045
rect 3070 1990 3180 2010
rect 3070 1955 3075 1990
rect 3175 1955 3180 1990
rect 3070 1930 3180 1955
rect 3320 2045 3430 2070
rect 3320 2010 3325 2045
rect 3425 2010 3430 2045
rect 3320 1990 3430 2010
rect 3320 1955 3325 1990
rect 3425 1955 3430 1990
rect 3320 1930 3430 1955
rect 3570 2045 3680 2070
rect 3570 2010 3575 2045
rect 3675 2010 3680 2045
rect 3570 1990 3680 2010
rect 3570 1955 3575 1990
rect 3675 1955 3680 1990
rect 3570 1930 3680 1955
rect 3820 2045 3930 2070
rect 3820 2010 3825 2045
rect 3925 2010 3930 2045
rect 3820 1990 3930 2010
rect 3820 1955 3825 1990
rect 3925 1955 3930 1990
rect 3820 1930 3930 1955
rect 4070 2045 4180 2070
rect 4070 2010 4075 2045
rect 4175 2010 4180 2045
rect 4070 1990 4180 2010
rect 4070 1955 4075 1990
rect 4175 1955 4180 1990
rect 4070 1930 4180 1955
rect 4320 2045 4430 2070
rect 4320 2010 4325 2045
rect 4425 2010 4430 2045
rect 4320 1990 4430 2010
rect 4320 1955 4325 1990
rect 4425 1955 4430 1990
rect 4320 1930 4430 1955
rect 4570 2045 4680 2070
rect 4570 2010 4575 2045
rect 4675 2010 4680 2045
rect 4570 1990 4680 2010
rect 4570 1955 4575 1990
rect 4675 1955 4680 1990
rect 4570 1930 4680 1955
rect 4820 2045 4930 2070
rect 4820 2010 4825 2045
rect 4925 2010 4930 2045
rect 4820 1990 4930 2010
rect 4820 1955 4825 1990
rect 4925 1955 4930 1990
rect 4820 1930 4930 1955
rect 5070 2045 5180 2070
rect 5070 2010 5075 2045
rect 5175 2010 5180 2045
rect 5070 1990 5180 2010
rect 5070 1955 5075 1990
rect 5175 1955 5180 1990
rect 5070 1930 5180 1955
rect 5320 2045 5430 2070
rect 5320 2010 5325 2045
rect 5425 2010 5430 2045
rect 5320 1990 5430 2010
rect 5320 1955 5325 1990
rect 5425 1955 5430 1990
rect 5320 1930 5430 1955
rect 5570 2045 5680 2070
rect 5570 2010 5575 2045
rect 5675 2010 5680 2045
rect 5570 1990 5680 2010
rect 5570 1955 5575 1990
rect 5675 1955 5680 1990
rect 5570 1930 5680 1955
rect 5820 2045 5930 2070
rect 5820 2010 5825 2045
rect 5925 2010 5930 2045
rect 5820 1990 5930 2010
rect 5820 1955 5825 1990
rect 5925 1955 5930 1990
rect 5820 1930 5930 1955
rect 6070 2045 6180 2070
rect 6070 2010 6075 2045
rect 6175 2010 6180 2045
rect 6070 1990 6180 2010
rect 6070 1955 6075 1990
rect 6175 1955 6180 1990
rect 6070 1930 6180 1955
rect 6320 2045 6430 2070
rect 6320 2010 6325 2045
rect 6425 2010 6430 2045
rect 6320 1990 6430 2010
rect 6320 1955 6325 1990
rect 6425 1955 6430 1990
rect 6320 1930 6430 1955
rect 6570 2045 6680 2070
rect 6570 2010 6575 2045
rect 6675 2010 6680 2045
rect 6570 1990 6680 2010
rect 6570 1955 6575 1990
rect 6675 1955 6680 1990
rect 6570 1930 6680 1955
rect 6820 2045 6930 2070
rect 6820 2010 6825 2045
rect 6925 2010 6930 2045
rect 6820 1990 6930 2010
rect 6820 1955 6825 1990
rect 6925 1955 6930 1990
rect 6820 1930 6930 1955
rect 7070 2045 7180 2070
rect 7070 2010 7075 2045
rect 7175 2010 7180 2045
rect 7070 1990 7180 2010
rect 7070 1955 7075 1990
rect 7175 1955 7180 1990
rect 7070 1930 7180 1955
rect 7320 2045 7430 2070
rect 7320 2010 7325 2045
rect 7425 2010 7430 2045
rect 7320 1990 7430 2010
rect 7320 1955 7325 1990
rect 7425 1955 7430 1990
rect 7320 1930 7430 1955
rect 7570 2045 7680 2070
rect 7570 2010 7575 2045
rect 7675 2010 7680 2045
rect 7570 1990 7680 2010
rect 7570 1955 7575 1990
rect 7675 1955 7680 1990
rect 7570 1930 7680 1955
rect 7820 2045 7930 2070
rect 7820 2010 7825 2045
rect 7925 2010 7930 2045
rect 7820 1990 7930 2010
rect 7820 1955 7825 1990
rect 7925 1955 7930 1990
rect 7820 1930 7930 1955
rect 0 1925 8000 1930
rect 0 1825 10 1925
rect 45 1825 205 1925
rect 240 1825 260 1925
rect 295 1825 455 1925
rect 490 1825 510 1925
rect 545 1825 705 1925
rect 740 1825 760 1925
rect 795 1825 955 1925
rect 990 1825 1010 1925
rect 1045 1825 1205 1925
rect 1240 1825 1260 1925
rect 1295 1825 1455 1925
rect 1490 1825 1510 1925
rect 1545 1825 1705 1925
rect 1740 1825 1760 1925
rect 1795 1825 1955 1925
rect 1990 1825 2010 1925
rect 2045 1825 2205 1925
rect 2240 1825 2260 1925
rect 2295 1825 2455 1925
rect 2490 1825 2510 1925
rect 2545 1825 2705 1925
rect 2740 1825 2760 1925
rect 2795 1825 2955 1925
rect 2990 1825 3010 1925
rect 3045 1825 3205 1925
rect 3240 1825 3260 1925
rect 3295 1825 3455 1925
rect 3490 1825 3510 1925
rect 3545 1825 3705 1925
rect 3740 1825 3760 1925
rect 3795 1825 3955 1925
rect 3990 1825 4010 1925
rect 4045 1825 4205 1925
rect 4240 1825 4260 1925
rect 4295 1825 4455 1925
rect 4490 1825 4510 1925
rect 4545 1825 4705 1925
rect 4740 1825 4760 1925
rect 4795 1825 4955 1925
rect 4990 1825 5010 1925
rect 5045 1825 5205 1925
rect 5240 1825 5260 1925
rect 5295 1825 5455 1925
rect 5490 1825 5510 1925
rect 5545 1825 5705 1925
rect 5740 1825 5760 1925
rect 5795 1825 5955 1925
rect 5990 1825 6010 1925
rect 6045 1825 6205 1925
rect 6240 1825 6260 1925
rect 6295 1825 6455 1925
rect 6490 1825 6510 1925
rect 6545 1825 6705 1925
rect 6740 1825 6760 1925
rect 6795 1825 6955 1925
rect 6990 1825 7010 1925
rect 7045 1825 7205 1925
rect 7240 1825 7260 1925
rect 7295 1825 7455 1925
rect 7490 1825 7510 1925
rect 7545 1825 7705 1925
rect 7740 1825 7760 1925
rect 7795 1825 7955 1925
rect 7990 1825 8000 1925
rect 0 1820 8000 1825
rect 70 1795 180 1820
rect 70 1760 75 1795
rect 175 1760 180 1795
rect 70 1740 180 1760
rect 70 1705 75 1740
rect 175 1705 180 1740
rect 70 1680 180 1705
rect 320 1795 430 1820
rect 320 1760 325 1795
rect 425 1760 430 1795
rect 320 1740 430 1760
rect 320 1705 325 1740
rect 425 1705 430 1740
rect 320 1680 430 1705
rect 570 1795 680 1820
rect 570 1760 575 1795
rect 675 1760 680 1795
rect 570 1740 680 1760
rect 570 1705 575 1740
rect 675 1705 680 1740
rect 570 1680 680 1705
rect 820 1795 930 1820
rect 820 1760 825 1795
rect 925 1760 930 1795
rect 820 1740 930 1760
rect 820 1705 825 1740
rect 925 1705 930 1740
rect 820 1680 930 1705
rect 1070 1795 1180 1820
rect 1070 1760 1075 1795
rect 1175 1760 1180 1795
rect 1070 1740 1180 1760
rect 1070 1705 1075 1740
rect 1175 1705 1180 1740
rect 1070 1680 1180 1705
rect 1320 1795 1430 1820
rect 1320 1760 1325 1795
rect 1425 1760 1430 1795
rect 1320 1740 1430 1760
rect 1320 1705 1325 1740
rect 1425 1705 1430 1740
rect 1320 1680 1430 1705
rect 1570 1795 1680 1820
rect 1570 1760 1575 1795
rect 1675 1760 1680 1795
rect 1570 1740 1680 1760
rect 1570 1705 1575 1740
rect 1675 1705 1680 1740
rect 1570 1680 1680 1705
rect 1820 1795 1930 1820
rect 1820 1760 1825 1795
rect 1925 1760 1930 1795
rect 1820 1740 1930 1760
rect 1820 1705 1825 1740
rect 1925 1705 1930 1740
rect 1820 1680 1930 1705
rect 2070 1795 2180 1820
rect 2070 1760 2075 1795
rect 2175 1760 2180 1795
rect 2070 1740 2180 1760
rect 2070 1705 2075 1740
rect 2175 1705 2180 1740
rect 2070 1680 2180 1705
rect 2320 1795 2430 1820
rect 2320 1760 2325 1795
rect 2425 1760 2430 1795
rect 2320 1740 2430 1760
rect 2320 1705 2325 1740
rect 2425 1705 2430 1740
rect 2320 1680 2430 1705
rect 2570 1795 2680 1820
rect 2570 1760 2575 1795
rect 2675 1760 2680 1795
rect 2570 1740 2680 1760
rect 2570 1705 2575 1740
rect 2675 1705 2680 1740
rect 2570 1680 2680 1705
rect 2820 1795 2930 1820
rect 2820 1760 2825 1795
rect 2925 1760 2930 1795
rect 2820 1740 2930 1760
rect 2820 1705 2825 1740
rect 2925 1705 2930 1740
rect 2820 1680 2930 1705
rect 3070 1795 3180 1820
rect 3070 1760 3075 1795
rect 3175 1760 3180 1795
rect 3070 1740 3180 1760
rect 3070 1705 3075 1740
rect 3175 1705 3180 1740
rect 3070 1680 3180 1705
rect 3320 1795 3430 1820
rect 3320 1760 3325 1795
rect 3425 1760 3430 1795
rect 3320 1740 3430 1760
rect 3320 1705 3325 1740
rect 3425 1705 3430 1740
rect 3320 1680 3430 1705
rect 3570 1795 3680 1820
rect 3570 1760 3575 1795
rect 3675 1760 3680 1795
rect 3570 1740 3680 1760
rect 3570 1705 3575 1740
rect 3675 1705 3680 1740
rect 3570 1680 3680 1705
rect 3820 1795 3930 1820
rect 3820 1760 3825 1795
rect 3925 1760 3930 1795
rect 3820 1740 3930 1760
rect 3820 1705 3825 1740
rect 3925 1705 3930 1740
rect 3820 1680 3930 1705
rect 4070 1795 4180 1820
rect 4070 1760 4075 1795
rect 4175 1760 4180 1795
rect 4070 1740 4180 1760
rect 4070 1705 4075 1740
rect 4175 1705 4180 1740
rect 4070 1680 4180 1705
rect 4320 1795 4430 1820
rect 4320 1760 4325 1795
rect 4425 1760 4430 1795
rect 4320 1740 4430 1760
rect 4320 1705 4325 1740
rect 4425 1705 4430 1740
rect 4320 1680 4430 1705
rect 4570 1795 4680 1820
rect 4570 1760 4575 1795
rect 4675 1760 4680 1795
rect 4570 1740 4680 1760
rect 4570 1705 4575 1740
rect 4675 1705 4680 1740
rect 4570 1680 4680 1705
rect 4820 1795 4930 1820
rect 4820 1760 4825 1795
rect 4925 1760 4930 1795
rect 4820 1740 4930 1760
rect 4820 1705 4825 1740
rect 4925 1705 4930 1740
rect 4820 1680 4930 1705
rect 5070 1795 5180 1820
rect 5070 1760 5075 1795
rect 5175 1760 5180 1795
rect 5070 1740 5180 1760
rect 5070 1705 5075 1740
rect 5175 1705 5180 1740
rect 5070 1680 5180 1705
rect 5320 1795 5430 1820
rect 5320 1760 5325 1795
rect 5425 1760 5430 1795
rect 5320 1740 5430 1760
rect 5320 1705 5325 1740
rect 5425 1705 5430 1740
rect 5320 1680 5430 1705
rect 5570 1795 5680 1820
rect 5570 1760 5575 1795
rect 5675 1760 5680 1795
rect 5570 1740 5680 1760
rect 5570 1705 5575 1740
rect 5675 1705 5680 1740
rect 5570 1680 5680 1705
rect 5820 1795 5930 1820
rect 5820 1760 5825 1795
rect 5925 1760 5930 1795
rect 5820 1740 5930 1760
rect 5820 1705 5825 1740
rect 5925 1705 5930 1740
rect 5820 1680 5930 1705
rect 6070 1795 6180 1820
rect 6070 1760 6075 1795
rect 6175 1760 6180 1795
rect 6070 1740 6180 1760
rect 6070 1705 6075 1740
rect 6175 1705 6180 1740
rect 6070 1680 6180 1705
rect 6320 1795 6430 1820
rect 6320 1760 6325 1795
rect 6425 1760 6430 1795
rect 6320 1740 6430 1760
rect 6320 1705 6325 1740
rect 6425 1705 6430 1740
rect 6320 1680 6430 1705
rect 6570 1795 6680 1820
rect 6570 1760 6575 1795
rect 6675 1760 6680 1795
rect 6570 1740 6680 1760
rect 6570 1705 6575 1740
rect 6675 1705 6680 1740
rect 6570 1680 6680 1705
rect 6820 1795 6930 1820
rect 6820 1760 6825 1795
rect 6925 1760 6930 1795
rect 6820 1740 6930 1760
rect 6820 1705 6825 1740
rect 6925 1705 6930 1740
rect 6820 1680 6930 1705
rect 7070 1795 7180 1820
rect 7070 1760 7075 1795
rect 7175 1760 7180 1795
rect 7070 1740 7180 1760
rect 7070 1705 7075 1740
rect 7175 1705 7180 1740
rect 7070 1680 7180 1705
rect 7320 1795 7430 1820
rect 7320 1760 7325 1795
rect 7425 1760 7430 1795
rect 7320 1740 7430 1760
rect 7320 1705 7325 1740
rect 7425 1705 7430 1740
rect 7320 1680 7430 1705
rect 7570 1795 7680 1820
rect 7570 1760 7575 1795
rect 7675 1760 7680 1795
rect 7570 1740 7680 1760
rect 7570 1705 7575 1740
rect 7675 1705 7680 1740
rect 7570 1680 7680 1705
rect 7820 1795 7930 1820
rect 7820 1760 7825 1795
rect 7925 1760 7930 1795
rect 7820 1740 7930 1760
rect 7820 1705 7825 1740
rect 7925 1705 7930 1740
rect 7820 1680 7930 1705
rect 0 1675 8000 1680
rect 0 1575 10 1675
rect 45 1575 205 1675
rect 240 1575 260 1675
rect 295 1575 455 1675
rect 490 1575 510 1675
rect 545 1575 705 1675
rect 740 1575 760 1675
rect 795 1575 955 1675
rect 990 1575 1010 1675
rect 1045 1575 1205 1675
rect 1240 1575 1260 1675
rect 1295 1575 1455 1675
rect 1490 1575 1510 1675
rect 1545 1575 1705 1675
rect 1740 1575 1760 1675
rect 1795 1575 1955 1675
rect 1990 1575 2010 1675
rect 2045 1575 2205 1675
rect 2240 1575 2260 1675
rect 2295 1575 2455 1675
rect 2490 1575 2510 1675
rect 2545 1575 2705 1675
rect 2740 1575 2760 1675
rect 2795 1575 2955 1675
rect 2990 1575 3010 1675
rect 3045 1575 3205 1675
rect 3240 1575 3260 1675
rect 3295 1575 3455 1675
rect 3490 1575 3510 1675
rect 3545 1575 3705 1675
rect 3740 1575 3760 1675
rect 3795 1575 3955 1675
rect 3990 1575 4010 1675
rect 4045 1575 4205 1675
rect 4240 1575 4260 1675
rect 4295 1575 4455 1675
rect 4490 1575 4510 1675
rect 4545 1575 4705 1675
rect 4740 1575 4760 1675
rect 4795 1575 4955 1675
rect 4990 1575 5010 1675
rect 5045 1575 5205 1675
rect 5240 1575 5260 1675
rect 5295 1575 5455 1675
rect 5490 1575 5510 1675
rect 5545 1575 5705 1675
rect 5740 1575 5760 1675
rect 5795 1575 5955 1675
rect 5990 1575 6010 1675
rect 6045 1575 6205 1675
rect 6240 1575 6260 1675
rect 6295 1575 6455 1675
rect 6490 1575 6510 1675
rect 6545 1575 6705 1675
rect 6740 1575 6760 1675
rect 6795 1575 6955 1675
rect 6990 1575 7010 1675
rect 7045 1575 7205 1675
rect 7240 1575 7260 1675
rect 7295 1575 7455 1675
rect 7490 1575 7510 1675
rect 7545 1575 7705 1675
rect 7740 1575 7760 1675
rect 7795 1575 7955 1675
rect 7990 1575 8000 1675
rect 0 1570 8000 1575
rect 70 1545 180 1570
rect 70 1510 75 1545
rect 175 1510 180 1545
rect 70 1490 180 1510
rect 70 1455 75 1490
rect 175 1455 180 1490
rect 70 1430 180 1455
rect 320 1545 430 1570
rect 320 1510 325 1545
rect 425 1510 430 1545
rect 320 1490 430 1510
rect 320 1455 325 1490
rect 425 1455 430 1490
rect 320 1430 430 1455
rect 570 1545 680 1570
rect 570 1510 575 1545
rect 675 1510 680 1545
rect 570 1490 680 1510
rect 570 1455 575 1490
rect 675 1455 680 1490
rect 570 1430 680 1455
rect 820 1545 930 1570
rect 820 1510 825 1545
rect 925 1510 930 1545
rect 820 1490 930 1510
rect 820 1455 825 1490
rect 925 1455 930 1490
rect 820 1430 930 1455
rect 1070 1545 1180 1570
rect 1070 1510 1075 1545
rect 1175 1510 1180 1545
rect 1070 1490 1180 1510
rect 1070 1455 1075 1490
rect 1175 1455 1180 1490
rect 1070 1430 1180 1455
rect 1320 1545 1430 1570
rect 1320 1510 1325 1545
rect 1425 1510 1430 1545
rect 1320 1490 1430 1510
rect 1320 1455 1325 1490
rect 1425 1455 1430 1490
rect 1320 1430 1430 1455
rect 1570 1545 1680 1570
rect 1570 1510 1575 1545
rect 1675 1510 1680 1545
rect 1570 1490 1680 1510
rect 1570 1455 1575 1490
rect 1675 1455 1680 1490
rect 1570 1430 1680 1455
rect 1820 1545 1930 1570
rect 1820 1510 1825 1545
rect 1925 1510 1930 1545
rect 1820 1490 1930 1510
rect 1820 1455 1825 1490
rect 1925 1455 1930 1490
rect 1820 1430 1930 1455
rect 2070 1545 2180 1570
rect 2070 1510 2075 1545
rect 2175 1510 2180 1545
rect 2070 1490 2180 1510
rect 2070 1455 2075 1490
rect 2175 1455 2180 1490
rect 2070 1430 2180 1455
rect 2320 1545 2430 1570
rect 2320 1510 2325 1545
rect 2425 1510 2430 1545
rect 2320 1490 2430 1510
rect 2320 1455 2325 1490
rect 2425 1455 2430 1490
rect 2320 1430 2430 1455
rect 2570 1545 2680 1570
rect 2570 1510 2575 1545
rect 2675 1510 2680 1545
rect 2570 1490 2680 1510
rect 2570 1455 2575 1490
rect 2675 1455 2680 1490
rect 2570 1430 2680 1455
rect 2820 1545 2930 1570
rect 2820 1510 2825 1545
rect 2925 1510 2930 1545
rect 2820 1490 2930 1510
rect 2820 1455 2825 1490
rect 2925 1455 2930 1490
rect 2820 1430 2930 1455
rect 3070 1545 3180 1570
rect 3070 1510 3075 1545
rect 3175 1510 3180 1545
rect 3070 1490 3180 1510
rect 3070 1455 3075 1490
rect 3175 1455 3180 1490
rect 3070 1430 3180 1455
rect 3320 1545 3430 1570
rect 3320 1510 3325 1545
rect 3425 1510 3430 1545
rect 3320 1490 3430 1510
rect 3320 1455 3325 1490
rect 3425 1455 3430 1490
rect 3320 1430 3430 1455
rect 3570 1545 3680 1570
rect 3570 1510 3575 1545
rect 3675 1510 3680 1545
rect 3570 1490 3680 1510
rect 3570 1455 3575 1490
rect 3675 1455 3680 1490
rect 3570 1430 3680 1455
rect 3820 1545 3930 1570
rect 3820 1510 3825 1545
rect 3925 1510 3930 1545
rect 3820 1490 3930 1510
rect 3820 1455 3825 1490
rect 3925 1455 3930 1490
rect 3820 1430 3930 1455
rect 4070 1545 4180 1570
rect 4070 1510 4075 1545
rect 4175 1510 4180 1545
rect 4070 1490 4180 1510
rect 4070 1455 4075 1490
rect 4175 1455 4180 1490
rect 4070 1430 4180 1455
rect 4320 1545 4430 1570
rect 4320 1510 4325 1545
rect 4425 1510 4430 1545
rect 4320 1490 4430 1510
rect 4320 1455 4325 1490
rect 4425 1455 4430 1490
rect 4320 1430 4430 1455
rect 4570 1545 4680 1570
rect 4570 1510 4575 1545
rect 4675 1510 4680 1545
rect 4570 1490 4680 1510
rect 4570 1455 4575 1490
rect 4675 1455 4680 1490
rect 4570 1430 4680 1455
rect 4820 1545 4930 1570
rect 4820 1510 4825 1545
rect 4925 1510 4930 1545
rect 4820 1490 4930 1510
rect 4820 1455 4825 1490
rect 4925 1455 4930 1490
rect 4820 1430 4930 1455
rect 5070 1545 5180 1570
rect 5070 1510 5075 1545
rect 5175 1510 5180 1545
rect 5070 1490 5180 1510
rect 5070 1455 5075 1490
rect 5175 1455 5180 1490
rect 5070 1430 5180 1455
rect 5320 1545 5430 1570
rect 5320 1510 5325 1545
rect 5425 1510 5430 1545
rect 5320 1490 5430 1510
rect 5320 1455 5325 1490
rect 5425 1455 5430 1490
rect 5320 1430 5430 1455
rect 5570 1545 5680 1570
rect 5570 1510 5575 1545
rect 5675 1510 5680 1545
rect 5570 1490 5680 1510
rect 5570 1455 5575 1490
rect 5675 1455 5680 1490
rect 5570 1430 5680 1455
rect 5820 1545 5930 1570
rect 5820 1510 5825 1545
rect 5925 1510 5930 1545
rect 5820 1490 5930 1510
rect 5820 1455 5825 1490
rect 5925 1455 5930 1490
rect 5820 1430 5930 1455
rect 6070 1545 6180 1570
rect 6070 1510 6075 1545
rect 6175 1510 6180 1545
rect 6070 1490 6180 1510
rect 6070 1455 6075 1490
rect 6175 1455 6180 1490
rect 6070 1430 6180 1455
rect 6320 1545 6430 1570
rect 6320 1510 6325 1545
rect 6425 1510 6430 1545
rect 6320 1490 6430 1510
rect 6320 1455 6325 1490
rect 6425 1455 6430 1490
rect 6320 1430 6430 1455
rect 6570 1545 6680 1570
rect 6570 1510 6575 1545
rect 6675 1510 6680 1545
rect 6570 1490 6680 1510
rect 6570 1455 6575 1490
rect 6675 1455 6680 1490
rect 6570 1430 6680 1455
rect 6820 1545 6930 1570
rect 6820 1510 6825 1545
rect 6925 1510 6930 1545
rect 6820 1490 6930 1510
rect 6820 1455 6825 1490
rect 6925 1455 6930 1490
rect 6820 1430 6930 1455
rect 7070 1545 7180 1570
rect 7070 1510 7075 1545
rect 7175 1510 7180 1545
rect 7070 1490 7180 1510
rect 7070 1455 7075 1490
rect 7175 1455 7180 1490
rect 7070 1430 7180 1455
rect 7320 1545 7430 1570
rect 7320 1510 7325 1545
rect 7425 1510 7430 1545
rect 7320 1490 7430 1510
rect 7320 1455 7325 1490
rect 7425 1455 7430 1490
rect 7320 1430 7430 1455
rect 7570 1545 7680 1570
rect 7570 1510 7575 1545
rect 7675 1510 7680 1545
rect 7570 1490 7680 1510
rect 7570 1455 7575 1490
rect 7675 1455 7680 1490
rect 7570 1430 7680 1455
rect 7820 1545 7930 1570
rect 7820 1510 7825 1545
rect 7925 1510 7930 1545
rect 7820 1490 7930 1510
rect 7820 1455 7825 1490
rect 7925 1455 7930 1490
rect 7820 1430 7930 1455
rect 0 1425 8000 1430
rect 0 1325 10 1425
rect 45 1325 205 1425
rect 240 1325 260 1425
rect 295 1325 455 1425
rect 490 1325 510 1425
rect 545 1325 705 1425
rect 740 1325 760 1425
rect 795 1325 955 1425
rect 990 1325 1010 1425
rect 1045 1325 1205 1425
rect 1240 1325 1260 1425
rect 1295 1325 1455 1425
rect 1490 1325 1510 1425
rect 1545 1325 1705 1425
rect 1740 1325 1760 1425
rect 1795 1325 1955 1425
rect 1990 1325 2010 1425
rect 2045 1325 2205 1425
rect 2240 1325 2260 1425
rect 2295 1325 2455 1425
rect 2490 1325 2510 1425
rect 2545 1325 2705 1425
rect 2740 1325 2760 1425
rect 2795 1325 2955 1425
rect 2990 1325 3010 1425
rect 3045 1325 3205 1425
rect 3240 1325 3260 1425
rect 3295 1325 3455 1425
rect 3490 1325 3510 1425
rect 3545 1325 3705 1425
rect 3740 1325 3760 1425
rect 3795 1325 3955 1425
rect 3990 1325 4010 1425
rect 4045 1325 4205 1425
rect 4240 1325 4260 1425
rect 4295 1325 4455 1425
rect 4490 1325 4510 1425
rect 4545 1325 4705 1425
rect 4740 1325 4760 1425
rect 4795 1325 4955 1425
rect 4990 1325 5010 1425
rect 5045 1325 5205 1425
rect 5240 1325 5260 1425
rect 5295 1325 5455 1425
rect 5490 1325 5510 1425
rect 5545 1325 5705 1425
rect 5740 1325 5760 1425
rect 5795 1325 5955 1425
rect 5990 1325 6010 1425
rect 6045 1325 6205 1425
rect 6240 1325 6260 1425
rect 6295 1325 6455 1425
rect 6490 1325 6510 1425
rect 6545 1325 6705 1425
rect 6740 1325 6760 1425
rect 6795 1325 6955 1425
rect 6990 1325 7010 1425
rect 7045 1325 7205 1425
rect 7240 1325 7260 1425
rect 7295 1325 7455 1425
rect 7490 1325 7510 1425
rect 7545 1325 7705 1425
rect 7740 1325 7760 1425
rect 7795 1325 7955 1425
rect 7990 1325 8000 1425
rect 0 1320 8000 1325
rect 70 1295 180 1320
rect 70 1260 75 1295
rect 175 1260 180 1295
rect 70 1240 180 1260
rect 70 1205 75 1240
rect 175 1205 180 1240
rect 70 1180 180 1205
rect 320 1295 430 1320
rect 320 1260 325 1295
rect 425 1260 430 1295
rect 320 1240 430 1260
rect 320 1205 325 1240
rect 425 1205 430 1240
rect 320 1180 430 1205
rect 570 1295 680 1320
rect 570 1260 575 1295
rect 675 1260 680 1295
rect 570 1240 680 1260
rect 570 1205 575 1240
rect 675 1205 680 1240
rect 570 1180 680 1205
rect 820 1295 930 1320
rect 820 1260 825 1295
rect 925 1260 930 1295
rect 820 1240 930 1260
rect 820 1205 825 1240
rect 925 1205 930 1240
rect 820 1180 930 1205
rect 1070 1295 1180 1320
rect 1070 1260 1075 1295
rect 1175 1260 1180 1295
rect 1070 1240 1180 1260
rect 1070 1205 1075 1240
rect 1175 1205 1180 1240
rect 1070 1180 1180 1205
rect 1320 1295 1430 1320
rect 1320 1260 1325 1295
rect 1425 1260 1430 1295
rect 1320 1240 1430 1260
rect 1320 1205 1325 1240
rect 1425 1205 1430 1240
rect 1320 1180 1430 1205
rect 1570 1295 1680 1320
rect 1570 1260 1575 1295
rect 1675 1260 1680 1295
rect 1570 1240 1680 1260
rect 1570 1205 1575 1240
rect 1675 1205 1680 1240
rect 1570 1180 1680 1205
rect 1820 1295 1930 1320
rect 1820 1260 1825 1295
rect 1925 1260 1930 1295
rect 1820 1240 1930 1260
rect 1820 1205 1825 1240
rect 1925 1205 1930 1240
rect 1820 1180 1930 1205
rect 2070 1295 2180 1320
rect 2070 1260 2075 1295
rect 2175 1260 2180 1295
rect 2070 1240 2180 1260
rect 2070 1205 2075 1240
rect 2175 1205 2180 1240
rect 2070 1180 2180 1205
rect 2320 1295 2430 1320
rect 2320 1260 2325 1295
rect 2425 1260 2430 1295
rect 2320 1240 2430 1260
rect 2320 1205 2325 1240
rect 2425 1205 2430 1240
rect 2320 1180 2430 1205
rect 2570 1295 2680 1320
rect 2570 1260 2575 1295
rect 2675 1260 2680 1295
rect 2570 1240 2680 1260
rect 2570 1205 2575 1240
rect 2675 1205 2680 1240
rect 2570 1180 2680 1205
rect 2820 1295 2930 1320
rect 2820 1260 2825 1295
rect 2925 1260 2930 1295
rect 2820 1240 2930 1260
rect 2820 1205 2825 1240
rect 2925 1205 2930 1240
rect 2820 1180 2930 1205
rect 3070 1295 3180 1320
rect 3070 1260 3075 1295
rect 3175 1260 3180 1295
rect 3070 1240 3180 1260
rect 3070 1205 3075 1240
rect 3175 1205 3180 1240
rect 3070 1180 3180 1205
rect 3320 1295 3430 1320
rect 3320 1260 3325 1295
rect 3425 1260 3430 1295
rect 3320 1240 3430 1260
rect 3320 1205 3325 1240
rect 3425 1205 3430 1240
rect 3320 1180 3430 1205
rect 3570 1295 3680 1320
rect 3570 1260 3575 1295
rect 3675 1260 3680 1295
rect 3570 1240 3680 1260
rect 3570 1205 3575 1240
rect 3675 1205 3680 1240
rect 3570 1180 3680 1205
rect 3820 1295 3930 1320
rect 3820 1260 3825 1295
rect 3925 1260 3930 1295
rect 3820 1240 3930 1260
rect 3820 1205 3825 1240
rect 3925 1205 3930 1240
rect 3820 1180 3930 1205
rect 4070 1295 4180 1320
rect 4070 1260 4075 1295
rect 4175 1260 4180 1295
rect 4070 1240 4180 1260
rect 4070 1205 4075 1240
rect 4175 1205 4180 1240
rect 4070 1180 4180 1205
rect 4320 1295 4430 1320
rect 4320 1260 4325 1295
rect 4425 1260 4430 1295
rect 4320 1240 4430 1260
rect 4320 1205 4325 1240
rect 4425 1205 4430 1240
rect 4320 1180 4430 1205
rect 4570 1295 4680 1320
rect 4570 1260 4575 1295
rect 4675 1260 4680 1295
rect 4570 1240 4680 1260
rect 4570 1205 4575 1240
rect 4675 1205 4680 1240
rect 4570 1180 4680 1205
rect 4820 1295 4930 1320
rect 4820 1260 4825 1295
rect 4925 1260 4930 1295
rect 4820 1240 4930 1260
rect 4820 1205 4825 1240
rect 4925 1205 4930 1240
rect 4820 1180 4930 1205
rect 5070 1295 5180 1320
rect 5070 1260 5075 1295
rect 5175 1260 5180 1295
rect 5070 1240 5180 1260
rect 5070 1205 5075 1240
rect 5175 1205 5180 1240
rect 5070 1180 5180 1205
rect 5320 1295 5430 1320
rect 5320 1260 5325 1295
rect 5425 1260 5430 1295
rect 5320 1240 5430 1260
rect 5320 1205 5325 1240
rect 5425 1205 5430 1240
rect 5320 1180 5430 1205
rect 5570 1295 5680 1320
rect 5570 1260 5575 1295
rect 5675 1260 5680 1295
rect 5570 1240 5680 1260
rect 5570 1205 5575 1240
rect 5675 1205 5680 1240
rect 5570 1180 5680 1205
rect 5820 1295 5930 1320
rect 5820 1260 5825 1295
rect 5925 1260 5930 1295
rect 5820 1240 5930 1260
rect 5820 1205 5825 1240
rect 5925 1205 5930 1240
rect 5820 1180 5930 1205
rect 6070 1295 6180 1320
rect 6070 1260 6075 1295
rect 6175 1260 6180 1295
rect 6070 1240 6180 1260
rect 6070 1205 6075 1240
rect 6175 1205 6180 1240
rect 6070 1180 6180 1205
rect 6320 1295 6430 1320
rect 6320 1260 6325 1295
rect 6425 1260 6430 1295
rect 6320 1240 6430 1260
rect 6320 1205 6325 1240
rect 6425 1205 6430 1240
rect 6320 1180 6430 1205
rect 6570 1295 6680 1320
rect 6570 1260 6575 1295
rect 6675 1260 6680 1295
rect 6570 1240 6680 1260
rect 6570 1205 6575 1240
rect 6675 1205 6680 1240
rect 6570 1180 6680 1205
rect 6820 1295 6930 1320
rect 6820 1260 6825 1295
rect 6925 1260 6930 1295
rect 6820 1240 6930 1260
rect 6820 1205 6825 1240
rect 6925 1205 6930 1240
rect 6820 1180 6930 1205
rect 7070 1295 7180 1320
rect 7070 1260 7075 1295
rect 7175 1260 7180 1295
rect 7070 1240 7180 1260
rect 7070 1205 7075 1240
rect 7175 1205 7180 1240
rect 7070 1180 7180 1205
rect 7320 1295 7430 1320
rect 7320 1260 7325 1295
rect 7425 1260 7430 1295
rect 7320 1240 7430 1260
rect 7320 1205 7325 1240
rect 7425 1205 7430 1240
rect 7320 1180 7430 1205
rect 7570 1295 7680 1320
rect 7570 1260 7575 1295
rect 7675 1260 7680 1295
rect 7570 1240 7680 1260
rect 7570 1205 7575 1240
rect 7675 1205 7680 1240
rect 7570 1180 7680 1205
rect 7820 1295 7930 1320
rect 7820 1260 7825 1295
rect 7925 1260 7930 1295
rect 7820 1240 7930 1260
rect 7820 1205 7825 1240
rect 7925 1205 7930 1240
rect 7820 1180 7930 1205
rect 0 1175 8000 1180
rect 0 1075 10 1175
rect 45 1075 205 1175
rect 240 1075 260 1175
rect 295 1075 455 1175
rect 490 1075 510 1175
rect 545 1075 705 1175
rect 740 1075 760 1175
rect 795 1075 955 1175
rect 990 1075 1010 1175
rect 1045 1075 1205 1175
rect 1240 1075 1260 1175
rect 1295 1075 1455 1175
rect 1490 1075 1510 1175
rect 1545 1075 1705 1175
rect 1740 1075 1760 1175
rect 1795 1075 1955 1175
rect 1990 1075 2010 1175
rect 2045 1075 2205 1175
rect 2240 1075 2260 1175
rect 2295 1075 2455 1175
rect 2490 1075 2510 1175
rect 2545 1075 2705 1175
rect 2740 1075 2760 1175
rect 2795 1075 2955 1175
rect 2990 1075 3010 1175
rect 3045 1075 3205 1175
rect 3240 1075 3260 1175
rect 3295 1075 3455 1175
rect 3490 1075 3510 1175
rect 3545 1075 3705 1175
rect 3740 1075 3760 1175
rect 3795 1075 3955 1175
rect 3990 1075 4010 1175
rect 4045 1075 4205 1175
rect 4240 1075 4260 1175
rect 4295 1075 4455 1175
rect 4490 1075 4510 1175
rect 4545 1075 4705 1175
rect 4740 1075 4760 1175
rect 4795 1075 4955 1175
rect 4990 1075 5010 1175
rect 5045 1075 5205 1175
rect 5240 1075 5260 1175
rect 5295 1075 5455 1175
rect 5490 1075 5510 1175
rect 5545 1075 5705 1175
rect 5740 1075 5760 1175
rect 5795 1075 5955 1175
rect 5990 1075 6010 1175
rect 6045 1075 6205 1175
rect 6240 1075 6260 1175
rect 6295 1075 6455 1175
rect 6490 1075 6510 1175
rect 6545 1075 6705 1175
rect 6740 1075 6760 1175
rect 6795 1075 6955 1175
rect 6990 1075 7010 1175
rect 7045 1075 7205 1175
rect 7240 1075 7260 1175
rect 7295 1075 7455 1175
rect 7490 1075 7510 1175
rect 7545 1075 7705 1175
rect 7740 1075 7760 1175
rect 7795 1075 7955 1175
rect 7990 1075 8000 1175
rect 0 1070 8000 1075
rect 70 1045 180 1070
rect 70 1010 75 1045
rect 175 1010 180 1045
rect 70 990 180 1010
rect 70 955 75 990
rect 175 955 180 990
rect 70 930 180 955
rect 320 1045 430 1070
rect 320 1010 325 1045
rect 425 1010 430 1045
rect 320 990 430 1010
rect 320 955 325 990
rect 425 955 430 990
rect 320 930 430 955
rect 570 1045 680 1070
rect 570 1010 575 1045
rect 675 1010 680 1045
rect 570 990 680 1010
rect 570 955 575 990
rect 675 955 680 990
rect 570 930 680 955
rect 820 1045 930 1070
rect 820 1010 825 1045
rect 925 1010 930 1045
rect 820 990 930 1010
rect 820 955 825 990
rect 925 955 930 990
rect 820 930 930 955
rect 1070 1045 1180 1070
rect 1070 1010 1075 1045
rect 1175 1010 1180 1045
rect 1070 990 1180 1010
rect 1070 955 1075 990
rect 1175 955 1180 990
rect 1070 930 1180 955
rect 1320 1045 1430 1070
rect 1320 1010 1325 1045
rect 1425 1010 1430 1045
rect 1320 990 1430 1010
rect 1320 955 1325 990
rect 1425 955 1430 990
rect 1320 930 1430 955
rect 1570 1045 1680 1070
rect 1570 1010 1575 1045
rect 1675 1010 1680 1045
rect 1570 990 1680 1010
rect 1570 955 1575 990
rect 1675 955 1680 990
rect 1570 930 1680 955
rect 1820 1045 1930 1070
rect 1820 1010 1825 1045
rect 1925 1010 1930 1045
rect 1820 990 1930 1010
rect 1820 955 1825 990
rect 1925 955 1930 990
rect 1820 930 1930 955
rect 2070 1045 2180 1070
rect 2070 1010 2075 1045
rect 2175 1010 2180 1045
rect 2070 990 2180 1010
rect 2070 955 2075 990
rect 2175 955 2180 990
rect 2070 930 2180 955
rect 2320 1045 2430 1070
rect 2320 1010 2325 1045
rect 2425 1010 2430 1045
rect 2320 990 2430 1010
rect 2320 955 2325 990
rect 2425 955 2430 990
rect 2320 930 2430 955
rect 2570 1045 2680 1070
rect 2570 1010 2575 1045
rect 2675 1010 2680 1045
rect 2570 990 2680 1010
rect 2570 955 2575 990
rect 2675 955 2680 990
rect 2570 930 2680 955
rect 2820 1045 2930 1070
rect 2820 1010 2825 1045
rect 2925 1010 2930 1045
rect 2820 990 2930 1010
rect 2820 955 2825 990
rect 2925 955 2930 990
rect 2820 930 2930 955
rect 3070 1045 3180 1070
rect 3070 1010 3075 1045
rect 3175 1010 3180 1045
rect 3070 990 3180 1010
rect 3070 955 3075 990
rect 3175 955 3180 990
rect 3070 930 3180 955
rect 3320 1045 3430 1070
rect 3320 1010 3325 1045
rect 3425 1010 3430 1045
rect 3320 990 3430 1010
rect 3320 955 3325 990
rect 3425 955 3430 990
rect 3320 930 3430 955
rect 3570 1045 3680 1070
rect 3570 1010 3575 1045
rect 3675 1010 3680 1045
rect 3570 990 3680 1010
rect 3570 955 3575 990
rect 3675 955 3680 990
rect 3570 930 3680 955
rect 3820 1045 3930 1070
rect 3820 1010 3825 1045
rect 3925 1010 3930 1045
rect 3820 990 3930 1010
rect 3820 955 3825 990
rect 3925 955 3930 990
rect 3820 930 3930 955
rect 4070 1045 4180 1070
rect 4070 1010 4075 1045
rect 4175 1010 4180 1045
rect 4070 990 4180 1010
rect 4070 955 4075 990
rect 4175 955 4180 990
rect 4070 930 4180 955
rect 4320 1045 4430 1070
rect 4320 1010 4325 1045
rect 4425 1010 4430 1045
rect 4320 990 4430 1010
rect 4320 955 4325 990
rect 4425 955 4430 990
rect 4320 930 4430 955
rect 4570 1045 4680 1070
rect 4570 1010 4575 1045
rect 4675 1010 4680 1045
rect 4570 990 4680 1010
rect 4570 955 4575 990
rect 4675 955 4680 990
rect 4570 930 4680 955
rect 4820 1045 4930 1070
rect 4820 1010 4825 1045
rect 4925 1010 4930 1045
rect 4820 990 4930 1010
rect 4820 955 4825 990
rect 4925 955 4930 990
rect 4820 930 4930 955
rect 5070 1045 5180 1070
rect 5070 1010 5075 1045
rect 5175 1010 5180 1045
rect 5070 990 5180 1010
rect 5070 955 5075 990
rect 5175 955 5180 990
rect 5070 930 5180 955
rect 5320 1045 5430 1070
rect 5320 1010 5325 1045
rect 5425 1010 5430 1045
rect 5320 990 5430 1010
rect 5320 955 5325 990
rect 5425 955 5430 990
rect 5320 930 5430 955
rect 5570 1045 5680 1070
rect 5570 1010 5575 1045
rect 5675 1010 5680 1045
rect 5570 990 5680 1010
rect 5570 955 5575 990
rect 5675 955 5680 990
rect 5570 930 5680 955
rect 5820 1045 5930 1070
rect 5820 1010 5825 1045
rect 5925 1010 5930 1045
rect 5820 990 5930 1010
rect 5820 955 5825 990
rect 5925 955 5930 990
rect 5820 930 5930 955
rect 6070 1045 6180 1070
rect 6070 1010 6075 1045
rect 6175 1010 6180 1045
rect 6070 990 6180 1010
rect 6070 955 6075 990
rect 6175 955 6180 990
rect 6070 930 6180 955
rect 6320 1045 6430 1070
rect 6320 1010 6325 1045
rect 6425 1010 6430 1045
rect 6320 990 6430 1010
rect 6320 955 6325 990
rect 6425 955 6430 990
rect 6320 930 6430 955
rect 6570 1045 6680 1070
rect 6570 1010 6575 1045
rect 6675 1010 6680 1045
rect 6570 990 6680 1010
rect 6570 955 6575 990
rect 6675 955 6680 990
rect 6570 930 6680 955
rect 6820 1045 6930 1070
rect 6820 1010 6825 1045
rect 6925 1010 6930 1045
rect 6820 990 6930 1010
rect 6820 955 6825 990
rect 6925 955 6930 990
rect 6820 930 6930 955
rect 7070 1045 7180 1070
rect 7070 1010 7075 1045
rect 7175 1010 7180 1045
rect 7070 990 7180 1010
rect 7070 955 7075 990
rect 7175 955 7180 990
rect 7070 930 7180 955
rect 7320 1045 7430 1070
rect 7320 1010 7325 1045
rect 7425 1010 7430 1045
rect 7320 990 7430 1010
rect 7320 955 7325 990
rect 7425 955 7430 990
rect 7320 930 7430 955
rect 7570 1045 7680 1070
rect 7570 1010 7575 1045
rect 7675 1010 7680 1045
rect 7570 990 7680 1010
rect 7570 955 7575 990
rect 7675 955 7680 990
rect 7570 930 7680 955
rect 7820 1045 7930 1070
rect 7820 1010 7825 1045
rect 7925 1010 7930 1045
rect 7820 990 7930 1010
rect 7820 955 7825 990
rect 7925 955 7930 990
rect 7820 930 7930 955
rect 0 925 8000 930
rect 0 825 10 925
rect 45 825 205 925
rect 240 825 260 925
rect 295 825 455 925
rect 490 825 510 925
rect 545 825 705 925
rect 740 825 760 925
rect 795 825 955 925
rect 990 825 1010 925
rect 1045 825 1205 925
rect 1240 825 1260 925
rect 1295 825 1455 925
rect 1490 825 1510 925
rect 1545 825 1705 925
rect 1740 825 1760 925
rect 1795 825 1955 925
rect 1990 825 2010 925
rect 2045 825 2205 925
rect 2240 825 2260 925
rect 2295 825 2455 925
rect 2490 825 2510 925
rect 2545 825 2705 925
rect 2740 825 2760 925
rect 2795 825 2955 925
rect 2990 825 3010 925
rect 3045 825 3205 925
rect 3240 825 3260 925
rect 3295 825 3455 925
rect 3490 825 3510 925
rect 3545 825 3705 925
rect 3740 825 3760 925
rect 3795 825 3955 925
rect 3990 825 4010 925
rect 4045 825 4205 925
rect 4240 825 4260 925
rect 4295 825 4455 925
rect 4490 825 4510 925
rect 4545 825 4705 925
rect 4740 825 4760 925
rect 4795 825 4955 925
rect 4990 825 5010 925
rect 5045 825 5205 925
rect 5240 825 5260 925
rect 5295 825 5455 925
rect 5490 825 5510 925
rect 5545 825 5705 925
rect 5740 825 5760 925
rect 5795 825 5955 925
rect 5990 825 6010 925
rect 6045 825 6205 925
rect 6240 825 6260 925
rect 6295 825 6455 925
rect 6490 825 6510 925
rect 6545 825 6705 925
rect 6740 825 6760 925
rect 6795 825 6955 925
rect 6990 825 7010 925
rect 7045 825 7205 925
rect 7240 825 7260 925
rect 7295 825 7455 925
rect 7490 825 7510 925
rect 7545 825 7705 925
rect 7740 825 7760 925
rect 7795 825 7955 925
rect 7990 825 8000 925
rect 0 820 8000 825
rect 70 795 180 820
rect 70 760 75 795
rect 175 760 180 795
rect 70 740 180 760
rect 70 705 75 740
rect 175 705 180 740
rect 70 680 180 705
rect 320 795 430 820
rect 320 760 325 795
rect 425 760 430 795
rect 320 740 430 760
rect 320 705 325 740
rect 425 705 430 740
rect 320 680 430 705
rect 570 795 680 820
rect 570 760 575 795
rect 675 760 680 795
rect 570 740 680 760
rect 570 705 575 740
rect 675 705 680 740
rect 570 680 680 705
rect 820 795 930 820
rect 820 760 825 795
rect 925 760 930 795
rect 820 740 930 760
rect 820 705 825 740
rect 925 705 930 740
rect 820 680 930 705
rect 1070 795 1180 820
rect 1070 760 1075 795
rect 1175 760 1180 795
rect 1070 740 1180 760
rect 1070 705 1075 740
rect 1175 705 1180 740
rect 1070 680 1180 705
rect 1320 795 1430 820
rect 1320 760 1325 795
rect 1425 760 1430 795
rect 1320 740 1430 760
rect 1320 705 1325 740
rect 1425 705 1430 740
rect 1320 680 1430 705
rect 1570 795 1680 820
rect 1570 760 1575 795
rect 1675 760 1680 795
rect 1570 740 1680 760
rect 1570 705 1575 740
rect 1675 705 1680 740
rect 1570 680 1680 705
rect 1820 795 1930 820
rect 1820 760 1825 795
rect 1925 760 1930 795
rect 1820 740 1930 760
rect 1820 705 1825 740
rect 1925 705 1930 740
rect 1820 680 1930 705
rect 2070 795 2180 820
rect 2070 760 2075 795
rect 2175 760 2180 795
rect 2070 740 2180 760
rect 2070 705 2075 740
rect 2175 705 2180 740
rect 2070 680 2180 705
rect 2320 795 2430 820
rect 2320 760 2325 795
rect 2425 760 2430 795
rect 2320 740 2430 760
rect 2320 705 2325 740
rect 2425 705 2430 740
rect 2320 680 2430 705
rect 2570 795 2680 820
rect 2570 760 2575 795
rect 2675 760 2680 795
rect 2570 740 2680 760
rect 2570 705 2575 740
rect 2675 705 2680 740
rect 2570 680 2680 705
rect 2820 795 2930 820
rect 2820 760 2825 795
rect 2925 760 2930 795
rect 2820 740 2930 760
rect 2820 705 2825 740
rect 2925 705 2930 740
rect 2820 680 2930 705
rect 3070 795 3180 820
rect 3070 760 3075 795
rect 3175 760 3180 795
rect 3070 740 3180 760
rect 3070 705 3075 740
rect 3175 705 3180 740
rect 3070 680 3180 705
rect 3320 795 3430 820
rect 3320 760 3325 795
rect 3425 760 3430 795
rect 3320 740 3430 760
rect 3320 705 3325 740
rect 3425 705 3430 740
rect 3320 680 3430 705
rect 3570 795 3680 820
rect 3570 760 3575 795
rect 3675 760 3680 795
rect 3570 740 3680 760
rect 3570 705 3575 740
rect 3675 705 3680 740
rect 3570 680 3680 705
rect 3820 795 3930 820
rect 3820 760 3825 795
rect 3925 760 3930 795
rect 3820 740 3930 760
rect 3820 705 3825 740
rect 3925 705 3930 740
rect 3820 680 3930 705
rect 4070 795 4180 820
rect 4070 760 4075 795
rect 4175 760 4180 795
rect 4070 740 4180 760
rect 4070 705 4075 740
rect 4175 705 4180 740
rect 4070 680 4180 705
rect 4320 795 4430 820
rect 4320 760 4325 795
rect 4425 760 4430 795
rect 4320 740 4430 760
rect 4320 705 4325 740
rect 4425 705 4430 740
rect 4320 680 4430 705
rect 4570 795 4680 820
rect 4570 760 4575 795
rect 4675 760 4680 795
rect 4570 740 4680 760
rect 4570 705 4575 740
rect 4675 705 4680 740
rect 4570 680 4680 705
rect 4820 795 4930 820
rect 4820 760 4825 795
rect 4925 760 4930 795
rect 4820 740 4930 760
rect 4820 705 4825 740
rect 4925 705 4930 740
rect 4820 680 4930 705
rect 5070 795 5180 820
rect 5070 760 5075 795
rect 5175 760 5180 795
rect 5070 740 5180 760
rect 5070 705 5075 740
rect 5175 705 5180 740
rect 5070 680 5180 705
rect 5320 795 5430 820
rect 5320 760 5325 795
rect 5425 760 5430 795
rect 5320 740 5430 760
rect 5320 705 5325 740
rect 5425 705 5430 740
rect 5320 680 5430 705
rect 5570 795 5680 820
rect 5570 760 5575 795
rect 5675 760 5680 795
rect 5570 740 5680 760
rect 5570 705 5575 740
rect 5675 705 5680 740
rect 5570 680 5680 705
rect 5820 795 5930 820
rect 5820 760 5825 795
rect 5925 760 5930 795
rect 5820 740 5930 760
rect 5820 705 5825 740
rect 5925 705 5930 740
rect 5820 680 5930 705
rect 6070 795 6180 820
rect 6070 760 6075 795
rect 6175 760 6180 795
rect 6070 740 6180 760
rect 6070 705 6075 740
rect 6175 705 6180 740
rect 6070 680 6180 705
rect 6320 795 6430 820
rect 6320 760 6325 795
rect 6425 760 6430 795
rect 6320 740 6430 760
rect 6320 705 6325 740
rect 6425 705 6430 740
rect 6320 680 6430 705
rect 6570 795 6680 820
rect 6570 760 6575 795
rect 6675 760 6680 795
rect 6570 740 6680 760
rect 6570 705 6575 740
rect 6675 705 6680 740
rect 6570 680 6680 705
rect 6820 795 6930 820
rect 6820 760 6825 795
rect 6925 760 6930 795
rect 6820 740 6930 760
rect 6820 705 6825 740
rect 6925 705 6930 740
rect 6820 680 6930 705
rect 7070 795 7180 820
rect 7070 760 7075 795
rect 7175 760 7180 795
rect 7070 740 7180 760
rect 7070 705 7075 740
rect 7175 705 7180 740
rect 7070 680 7180 705
rect 7320 795 7430 820
rect 7320 760 7325 795
rect 7425 760 7430 795
rect 7320 740 7430 760
rect 7320 705 7325 740
rect 7425 705 7430 740
rect 7320 680 7430 705
rect 7570 795 7680 820
rect 7570 760 7575 795
rect 7675 760 7680 795
rect 7570 740 7680 760
rect 7570 705 7575 740
rect 7675 705 7680 740
rect 7570 680 7680 705
rect 7820 795 7930 820
rect 7820 760 7825 795
rect 7925 760 7930 795
rect 7820 740 7930 760
rect 7820 705 7825 740
rect 7925 705 7930 740
rect 7820 680 7930 705
rect 0 675 8000 680
rect 0 575 10 675
rect 45 575 205 675
rect 240 575 260 675
rect 295 575 455 675
rect 490 575 510 675
rect 545 575 705 675
rect 740 575 760 675
rect 795 575 955 675
rect 990 575 1010 675
rect 1045 575 1205 675
rect 1240 575 1260 675
rect 1295 575 1455 675
rect 1490 575 1510 675
rect 1545 575 1705 675
rect 1740 575 1760 675
rect 1795 575 1955 675
rect 1990 575 2010 675
rect 2045 575 2205 675
rect 2240 575 2260 675
rect 2295 575 2455 675
rect 2490 575 2510 675
rect 2545 575 2705 675
rect 2740 575 2760 675
rect 2795 575 2955 675
rect 2990 575 3010 675
rect 3045 575 3205 675
rect 3240 575 3260 675
rect 3295 575 3455 675
rect 3490 575 3510 675
rect 3545 575 3705 675
rect 3740 575 3760 675
rect 3795 575 3955 675
rect 3990 575 4010 675
rect 4045 575 4205 675
rect 4240 575 4260 675
rect 4295 575 4455 675
rect 4490 575 4510 675
rect 4545 575 4705 675
rect 4740 575 4760 675
rect 4795 575 4955 675
rect 4990 575 5010 675
rect 5045 575 5205 675
rect 5240 575 5260 675
rect 5295 575 5455 675
rect 5490 575 5510 675
rect 5545 575 5705 675
rect 5740 575 5760 675
rect 5795 575 5955 675
rect 5990 575 6010 675
rect 6045 575 6205 675
rect 6240 575 6260 675
rect 6295 575 6455 675
rect 6490 575 6510 675
rect 6545 575 6705 675
rect 6740 575 6760 675
rect 6795 575 6955 675
rect 6990 575 7010 675
rect 7045 575 7205 675
rect 7240 575 7260 675
rect 7295 575 7455 675
rect 7490 575 7510 675
rect 7545 575 7705 675
rect 7740 575 7760 675
rect 7795 575 7955 675
rect 7990 575 8000 675
rect 0 570 8000 575
rect 70 545 180 570
rect 70 510 75 545
rect 175 510 180 545
rect 70 490 180 510
rect 70 455 75 490
rect 175 455 180 490
rect 70 430 180 455
rect 320 545 430 570
rect 320 510 325 545
rect 425 510 430 545
rect 320 490 430 510
rect 320 455 325 490
rect 425 455 430 490
rect 320 430 430 455
rect 570 545 680 570
rect 570 510 575 545
rect 675 510 680 545
rect 570 490 680 510
rect 570 455 575 490
rect 675 455 680 490
rect 570 430 680 455
rect 820 545 930 570
rect 820 510 825 545
rect 925 510 930 545
rect 820 490 930 510
rect 820 455 825 490
rect 925 455 930 490
rect 820 430 930 455
rect 1070 545 1180 570
rect 1070 510 1075 545
rect 1175 510 1180 545
rect 1070 490 1180 510
rect 1070 455 1075 490
rect 1175 455 1180 490
rect 1070 430 1180 455
rect 1320 545 1430 570
rect 1320 510 1325 545
rect 1425 510 1430 545
rect 1320 490 1430 510
rect 1320 455 1325 490
rect 1425 455 1430 490
rect 1320 430 1430 455
rect 1570 545 1680 570
rect 1570 510 1575 545
rect 1675 510 1680 545
rect 1570 490 1680 510
rect 1570 455 1575 490
rect 1675 455 1680 490
rect 1570 430 1680 455
rect 1820 545 1930 570
rect 1820 510 1825 545
rect 1925 510 1930 545
rect 1820 490 1930 510
rect 1820 455 1825 490
rect 1925 455 1930 490
rect 1820 430 1930 455
rect 2070 545 2180 570
rect 2070 510 2075 545
rect 2175 510 2180 545
rect 2070 490 2180 510
rect 2070 455 2075 490
rect 2175 455 2180 490
rect 2070 430 2180 455
rect 2320 545 2430 570
rect 2320 510 2325 545
rect 2425 510 2430 545
rect 2320 490 2430 510
rect 2320 455 2325 490
rect 2425 455 2430 490
rect 2320 430 2430 455
rect 2570 545 2680 570
rect 2570 510 2575 545
rect 2675 510 2680 545
rect 2570 490 2680 510
rect 2570 455 2575 490
rect 2675 455 2680 490
rect 2570 430 2680 455
rect 2820 545 2930 570
rect 2820 510 2825 545
rect 2925 510 2930 545
rect 2820 490 2930 510
rect 2820 455 2825 490
rect 2925 455 2930 490
rect 2820 430 2930 455
rect 3070 545 3180 570
rect 3070 510 3075 545
rect 3175 510 3180 545
rect 3070 490 3180 510
rect 3070 455 3075 490
rect 3175 455 3180 490
rect 3070 430 3180 455
rect 3320 545 3430 570
rect 3320 510 3325 545
rect 3425 510 3430 545
rect 3320 490 3430 510
rect 3320 455 3325 490
rect 3425 455 3430 490
rect 3320 430 3430 455
rect 3570 545 3680 570
rect 3570 510 3575 545
rect 3675 510 3680 545
rect 3570 490 3680 510
rect 3570 455 3575 490
rect 3675 455 3680 490
rect 3570 430 3680 455
rect 3820 545 3930 570
rect 3820 510 3825 545
rect 3925 510 3930 545
rect 3820 490 3930 510
rect 3820 455 3825 490
rect 3925 455 3930 490
rect 3820 430 3930 455
rect 4070 545 4180 570
rect 4070 510 4075 545
rect 4175 510 4180 545
rect 4070 490 4180 510
rect 4070 455 4075 490
rect 4175 455 4180 490
rect 4070 430 4180 455
rect 4320 545 4430 570
rect 4320 510 4325 545
rect 4425 510 4430 545
rect 4320 490 4430 510
rect 4320 455 4325 490
rect 4425 455 4430 490
rect 4320 430 4430 455
rect 4570 545 4680 570
rect 4570 510 4575 545
rect 4675 510 4680 545
rect 4570 490 4680 510
rect 4570 455 4575 490
rect 4675 455 4680 490
rect 4570 430 4680 455
rect 4820 545 4930 570
rect 4820 510 4825 545
rect 4925 510 4930 545
rect 4820 490 4930 510
rect 4820 455 4825 490
rect 4925 455 4930 490
rect 4820 430 4930 455
rect 5070 545 5180 570
rect 5070 510 5075 545
rect 5175 510 5180 545
rect 5070 490 5180 510
rect 5070 455 5075 490
rect 5175 455 5180 490
rect 5070 430 5180 455
rect 5320 545 5430 570
rect 5320 510 5325 545
rect 5425 510 5430 545
rect 5320 490 5430 510
rect 5320 455 5325 490
rect 5425 455 5430 490
rect 5320 430 5430 455
rect 5570 545 5680 570
rect 5570 510 5575 545
rect 5675 510 5680 545
rect 5570 490 5680 510
rect 5570 455 5575 490
rect 5675 455 5680 490
rect 5570 430 5680 455
rect 5820 545 5930 570
rect 5820 510 5825 545
rect 5925 510 5930 545
rect 5820 490 5930 510
rect 5820 455 5825 490
rect 5925 455 5930 490
rect 5820 430 5930 455
rect 6070 545 6180 570
rect 6070 510 6075 545
rect 6175 510 6180 545
rect 6070 490 6180 510
rect 6070 455 6075 490
rect 6175 455 6180 490
rect 6070 430 6180 455
rect 6320 545 6430 570
rect 6320 510 6325 545
rect 6425 510 6430 545
rect 6320 490 6430 510
rect 6320 455 6325 490
rect 6425 455 6430 490
rect 6320 430 6430 455
rect 6570 545 6680 570
rect 6570 510 6575 545
rect 6675 510 6680 545
rect 6570 490 6680 510
rect 6570 455 6575 490
rect 6675 455 6680 490
rect 6570 430 6680 455
rect 6820 545 6930 570
rect 6820 510 6825 545
rect 6925 510 6930 545
rect 6820 490 6930 510
rect 6820 455 6825 490
rect 6925 455 6930 490
rect 6820 430 6930 455
rect 7070 545 7180 570
rect 7070 510 7075 545
rect 7175 510 7180 545
rect 7070 490 7180 510
rect 7070 455 7075 490
rect 7175 455 7180 490
rect 7070 430 7180 455
rect 7320 545 7430 570
rect 7320 510 7325 545
rect 7425 510 7430 545
rect 7320 490 7430 510
rect 7320 455 7325 490
rect 7425 455 7430 490
rect 7320 430 7430 455
rect 7570 545 7680 570
rect 7570 510 7575 545
rect 7675 510 7680 545
rect 7570 490 7680 510
rect 7570 455 7575 490
rect 7675 455 7680 490
rect 7570 430 7680 455
rect 7820 545 7930 570
rect 7820 510 7825 545
rect 7925 510 7930 545
rect 7820 490 7930 510
rect 7820 455 7825 490
rect 7925 455 7930 490
rect 7820 430 7930 455
rect 0 425 8000 430
rect 0 325 10 425
rect 45 325 205 425
rect 240 325 260 425
rect 295 325 455 425
rect 490 325 510 425
rect 545 325 705 425
rect 740 325 760 425
rect 795 325 955 425
rect 990 325 1010 425
rect 1045 325 1205 425
rect 1240 325 1260 425
rect 1295 325 1455 425
rect 1490 325 1510 425
rect 1545 325 1705 425
rect 1740 325 1760 425
rect 1795 325 1955 425
rect 1990 325 2010 425
rect 2045 325 2205 425
rect 2240 325 2260 425
rect 2295 325 2455 425
rect 2490 325 2510 425
rect 2545 325 2705 425
rect 2740 325 2760 425
rect 2795 325 2955 425
rect 2990 325 3010 425
rect 3045 325 3205 425
rect 3240 325 3260 425
rect 3295 325 3455 425
rect 3490 325 3510 425
rect 3545 325 3705 425
rect 3740 325 3760 425
rect 3795 325 3955 425
rect 3990 325 4010 425
rect 4045 325 4205 425
rect 4240 325 4260 425
rect 4295 325 4455 425
rect 4490 325 4510 425
rect 4545 325 4705 425
rect 4740 325 4760 425
rect 4795 325 4955 425
rect 4990 325 5010 425
rect 5045 325 5205 425
rect 5240 325 5260 425
rect 5295 325 5455 425
rect 5490 325 5510 425
rect 5545 325 5705 425
rect 5740 325 5760 425
rect 5795 325 5955 425
rect 5990 325 6010 425
rect 6045 325 6205 425
rect 6240 325 6260 425
rect 6295 325 6455 425
rect 6490 325 6510 425
rect 6545 325 6705 425
rect 6740 325 6760 425
rect 6795 325 6955 425
rect 6990 325 7010 425
rect 7045 325 7205 425
rect 7240 325 7260 425
rect 7295 325 7455 425
rect 7490 325 7510 425
rect 7545 325 7705 425
rect 7740 325 7760 425
rect 7795 325 7955 425
rect 7990 325 8000 425
rect 0 320 8000 325
rect 70 295 180 320
rect 70 260 75 295
rect 175 260 180 295
rect 70 240 180 260
rect 70 205 75 240
rect 175 205 180 240
rect 70 180 180 205
rect 320 295 430 320
rect 320 260 325 295
rect 425 260 430 295
rect 320 240 430 260
rect 320 205 325 240
rect 425 205 430 240
rect 320 180 430 205
rect 570 295 680 320
rect 570 260 575 295
rect 675 260 680 295
rect 570 240 680 260
rect 570 205 575 240
rect 675 205 680 240
rect 570 180 680 205
rect 820 295 930 320
rect 820 260 825 295
rect 925 260 930 295
rect 820 240 930 260
rect 820 205 825 240
rect 925 205 930 240
rect 820 180 930 205
rect 1070 295 1180 320
rect 1070 260 1075 295
rect 1175 260 1180 295
rect 1070 240 1180 260
rect 1070 205 1075 240
rect 1175 205 1180 240
rect 1070 180 1180 205
rect 1320 295 1430 320
rect 1320 260 1325 295
rect 1425 260 1430 295
rect 1320 240 1430 260
rect 1320 205 1325 240
rect 1425 205 1430 240
rect 1320 180 1430 205
rect 1570 295 1680 320
rect 1570 260 1575 295
rect 1675 260 1680 295
rect 1570 240 1680 260
rect 1570 205 1575 240
rect 1675 205 1680 240
rect 1570 180 1680 205
rect 1820 295 1930 320
rect 1820 260 1825 295
rect 1925 260 1930 295
rect 1820 240 1930 260
rect 1820 205 1825 240
rect 1925 205 1930 240
rect 1820 180 1930 205
rect 2070 295 2180 320
rect 2070 260 2075 295
rect 2175 260 2180 295
rect 2070 240 2180 260
rect 2070 205 2075 240
rect 2175 205 2180 240
rect 2070 180 2180 205
rect 2320 295 2430 320
rect 2320 260 2325 295
rect 2425 260 2430 295
rect 2320 240 2430 260
rect 2320 205 2325 240
rect 2425 205 2430 240
rect 2320 180 2430 205
rect 2570 295 2680 320
rect 2570 260 2575 295
rect 2675 260 2680 295
rect 2570 240 2680 260
rect 2570 205 2575 240
rect 2675 205 2680 240
rect 2570 180 2680 205
rect 2820 295 2930 320
rect 2820 260 2825 295
rect 2925 260 2930 295
rect 2820 240 2930 260
rect 2820 205 2825 240
rect 2925 205 2930 240
rect 2820 180 2930 205
rect 3070 295 3180 320
rect 3070 260 3075 295
rect 3175 260 3180 295
rect 3070 240 3180 260
rect 3070 205 3075 240
rect 3175 205 3180 240
rect 3070 180 3180 205
rect 3320 295 3430 320
rect 3320 260 3325 295
rect 3425 260 3430 295
rect 3320 240 3430 260
rect 3320 205 3325 240
rect 3425 205 3430 240
rect 3320 180 3430 205
rect 3570 295 3680 320
rect 3570 260 3575 295
rect 3675 260 3680 295
rect 3570 240 3680 260
rect 3570 205 3575 240
rect 3675 205 3680 240
rect 3570 180 3680 205
rect 3820 295 3930 320
rect 3820 260 3825 295
rect 3925 260 3930 295
rect 3820 240 3930 260
rect 3820 205 3825 240
rect 3925 205 3930 240
rect 3820 180 3930 205
rect 4070 295 4180 320
rect 4070 260 4075 295
rect 4175 260 4180 295
rect 4070 240 4180 260
rect 4070 205 4075 240
rect 4175 205 4180 240
rect 4070 180 4180 205
rect 4320 295 4430 320
rect 4320 260 4325 295
rect 4425 260 4430 295
rect 4320 240 4430 260
rect 4320 205 4325 240
rect 4425 205 4430 240
rect 4320 180 4430 205
rect 4570 295 4680 320
rect 4570 260 4575 295
rect 4675 260 4680 295
rect 4570 240 4680 260
rect 4570 205 4575 240
rect 4675 205 4680 240
rect 4570 180 4680 205
rect 4820 295 4930 320
rect 4820 260 4825 295
rect 4925 260 4930 295
rect 4820 240 4930 260
rect 4820 205 4825 240
rect 4925 205 4930 240
rect 4820 180 4930 205
rect 5070 295 5180 320
rect 5070 260 5075 295
rect 5175 260 5180 295
rect 5070 240 5180 260
rect 5070 205 5075 240
rect 5175 205 5180 240
rect 5070 180 5180 205
rect 5320 295 5430 320
rect 5320 260 5325 295
rect 5425 260 5430 295
rect 5320 240 5430 260
rect 5320 205 5325 240
rect 5425 205 5430 240
rect 5320 180 5430 205
rect 5570 295 5680 320
rect 5570 260 5575 295
rect 5675 260 5680 295
rect 5570 240 5680 260
rect 5570 205 5575 240
rect 5675 205 5680 240
rect 5570 180 5680 205
rect 5820 295 5930 320
rect 5820 260 5825 295
rect 5925 260 5930 295
rect 5820 240 5930 260
rect 5820 205 5825 240
rect 5925 205 5930 240
rect 5820 180 5930 205
rect 6070 295 6180 320
rect 6070 260 6075 295
rect 6175 260 6180 295
rect 6070 240 6180 260
rect 6070 205 6075 240
rect 6175 205 6180 240
rect 6070 180 6180 205
rect 6320 295 6430 320
rect 6320 260 6325 295
rect 6425 260 6430 295
rect 6320 240 6430 260
rect 6320 205 6325 240
rect 6425 205 6430 240
rect 6320 180 6430 205
rect 6570 295 6680 320
rect 6570 260 6575 295
rect 6675 260 6680 295
rect 6570 240 6680 260
rect 6570 205 6575 240
rect 6675 205 6680 240
rect 6570 180 6680 205
rect 6820 295 6930 320
rect 6820 260 6825 295
rect 6925 260 6930 295
rect 6820 240 6930 260
rect 6820 205 6825 240
rect 6925 205 6930 240
rect 6820 180 6930 205
rect 7070 295 7180 320
rect 7070 260 7075 295
rect 7175 260 7180 295
rect 7070 240 7180 260
rect 7070 205 7075 240
rect 7175 205 7180 240
rect 7070 180 7180 205
rect 7320 295 7430 320
rect 7320 260 7325 295
rect 7425 260 7430 295
rect 7320 240 7430 260
rect 7320 205 7325 240
rect 7425 205 7430 240
rect 7320 180 7430 205
rect 7570 295 7680 320
rect 7570 260 7575 295
rect 7675 260 7680 295
rect 7570 240 7680 260
rect 7570 205 7575 240
rect 7675 205 7680 240
rect 7570 180 7680 205
rect 7820 295 7930 320
rect 7820 260 7825 295
rect 7925 260 7930 295
rect 7820 240 7930 260
rect 7820 205 7825 240
rect 7925 205 7930 240
rect 7820 180 7930 205
rect 0 175 8000 180
rect 0 75 10 175
rect 45 75 205 175
rect 240 75 260 175
rect 295 75 455 175
rect 490 75 510 175
rect 545 75 705 175
rect 740 75 760 175
rect 795 75 955 175
rect 990 75 1010 175
rect 1045 75 1205 175
rect 1240 75 1260 175
rect 1295 75 1455 175
rect 1490 75 1510 175
rect 1545 75 1705 175
rect 1740 75 1760 175
rect 1795 75 1955 175
rect 1990 75 2010 175
rect 2045 75 2205 175
rect 2240 75 2260 175
rect 2295 75 2455 175
rect 2490 75 2510 175
rect 2545 75 2705 175
rect 2740 75 2760 175
rect 2795 75 2955 175
rect 2990 75 3010 175
rect 3045 75 3205 175
rect 3240 75 3260 175
rect 3295 75 3455 175
rect 3490 75 3510 175
rect 3545 75 3705 175
rect 3740 75 3760 175
rect 3795 75 3955 175
rect 3990 75 4010 175
rect 4045 75 4205 175
rect 4240 75 4260 175
rect 4295 75 4455 175
rect 4490 75 4510 175
rect 4545 75 4705 175
rect 4740 75 4760 175
rect 4795 75 4955 175
rect 4990 75 5010 175
rect 5045 75 5205 175
rect 5240 75 5260 175
rect 5295 75 5455 175
rect 5490 75 5510 175
rect 5545 75 5705 175
rect 5740 75 5760 175
rect 5795 75 5955 175
rect 5990 75 6010 175
rect 6045 75 6205 175
rect 6240 75 6260 175
rect 6295 75 6455 175
rect 6490 75 6510 175
rect 6545 75 6705 175
rect 6740 75 6760 175
rect 6795 75 6955 175
rect 6990 75 7010 175
rect 7045 75 7205 175
rect 7240 75 7260 175
rect 7295 75 7455 175
rect 7490 75 7510 175
rect 7545 75 7705 175
rect 7740 75 7760 175
rect 7795 75 7955 175
rect 7990 75 8000 175
rect 0 70 8000 75
rect 70 45 180 70
rect 70 10 75 45
rect 175 10 180 45
rect 70 0 180 10
rect 320 45 430 70
rect 320 10 325 45
rect 425 10 430 45
rect 320 0 430 10
rect 570 45 680 70
rect 570 10 575 45
rect 675 10 680 45
rect 570 0 680 10
rect 820 45 930 70
rect 820 10 825 45
rect 925 10 930 45
rect 820 0 930 10
rect 1070 45 1180 70
rect 1070 10 1075 45
rect 1175 10 1180 45
rect 1070 0 1180 10
rect 1320 45 1430 70
rect 1320 10 1325 45
rect 1425 10 1430 45
rect 1320 0 1430 10
rect 1570 45 1680 70
rect 1570 10 1575 45
rect 1675 10 1680 45
rect 1570 0 1680 10
rect 1820 45 1930 70
rect 1820 10 1825 45
rect 1925 10 1930 45
rect 1820 0 1930 10
rect 2070 45 2180 70
rect 2070 10 2075 45
rect 2175 10 2180 45
rect 2070 0 2180 10
rect 2320 45 2430 70
rect 2320 10 2325 45
rect 2425 10 2430 45
rect 2320 0 2430 10
rect 2570 45 2680 70
rect 2570 10 2575 45
rect 2675 10 2680 45
rect 2570 0 2680 10
rect 2820 45 2930 70
rect 2820 10 2825 45
rect 2925 10 2930 45
rect 2820 0 2930 10
rect 3070 45 3180 70
rect 3070 10 3075 45
rect 3175 10 3180 45
rect 3070 0 3180 10
rect 3320 45 3430 70
rect 3320 10 3325 45
rect 3425 10 3430 45
rect 3320 0 3430 10
rect 3570 45 3680 70
rect 3570 10 3575 45
rect 3675 10 3680 45
rect 3570 0 3680 10
rect 3820 45 3930 70
rect 3820 10 3825 45
rect 3925 10 3930 45
rect 3820 0 3930 10
rect 4070 45 4180 70
rect 4070 10 4075 45
rect 4175 10 4180 45
rect 4070 0 4180 10
rect 4320 45 4430 70
rect 4320 10 4325 45
rect 4425 10 4430 45
rect 4320 0 4430 10
rect 4570 45 4680 70
rect 4570 10 4575 45
rect 4675 10 4680 45
rect 4570 0 4680 10
rect 4820 45 4930 70
rect 4820 10 4825 45
rect 4925 10 4930 45
rect 4820 0 4930 10
rect 5070 45 5180 70
rect 5070 10 5075 45
rect 5175 10 5180 45
rect 5070 0 5180 10
rect 5320 45 5430 70
rect 5320 10 5325 45
rect 5425 10 5430 45
rect 5320 0 5430 10
rect 5570 45 5680 70
rect 5570 10 5575 45
rect 5675 10 5680 45
rect 5570 0 5680 10
rect 5820 45 5930 70
rect 5820 10 5825 45
rect 5925 10 5930 45
rect 5820 0 5930 10
rect 6070 45 6180 70
rect 6070 10 6075 45
rect 6175 10 6180 45
rect 6070 0 6180 10
rect 6320 45 6430 70
rect 6320 10 6325 45
rect 6425 10 6430 45
rect 6320 0 6430 10
rect 6570 45 6680 70
rect 6570 10 6575 45
rect 6675 10 6680 45
rect 6570 0 6680 10
rect 6820 45 6930 70
rect 6820 10 6825 45
rect 6925 10 6930 45
rect 6820 0 6930 10
rect 7070 45 7180 70
rect 7070 10 7075 45
rect 7175 10 7180 45
rect 7070 0 7180 10
rect 7320 45 7430 70
rect 7320 10 7325 45
rect 7425 10 7430 45
rect 7320 0 7430 10
rect 7570 45 7680 70
rect 7570 10 7575 45
rect 7675 10 7680 45
rect 7570 0 7680 10
rect 7820 45 7930 70
rect 7820 10 7825 45
rect 7925 10 7930 45
rect 7820 0 7930 10
<< via2 >>
rect 75 7955 175 7990
rect 325 7955 425 7990
rect 575 7955 675 7990
rect 825 7955 925 7990
rect 1075 7955 1175 7990
rect 1325 7955 1425 7990
rect 1575 7955 1675 7990
rect 1825 7955 1925 7990
rect 2075 7955 2175 7990
rect 2325 7955 2425 7990
rect 2575 7955 2675 7990
rect 2825 7955 2925 7990
rect 3075 7955 3175 7990
rect 3325 7955 3425 7990
rect 3575 7955 3675 7990
rect 3825 7955 3925 7990
rect 4075 7955 4175 7990
rect 4325 7955 4425 7990
rect 4575 7955 4675 7990
rect 4825 7955 4925 7990
rect 5075 7955 5175 7990
rect 5325 7955 5425 7990
rect 5575 7955 5675 7990
rect 5825 7955 5925 7990
rect 6075 7955 6175 7990
rect 6325 7955 6425 7990
rect 6575 7955 6675 7990
rect 6825 7955 6925 7990
rect 7075 7955 7175 7990
rect 7325 7955 7425 7990
rect 7575 7955 7675 7990
rect 7825 7955 7925 7990
rect 10 7825 45 7925
rect 205 7825 240 7925
rect 260 7825 295 7925
rect 455 7825 490 7925
rect 510 7825 545 7925
rect 705 7825 740 7925
rect 760 7825 795 7925
rect 955 7825 990 7925
rect 1010 7825 1045 7925
rect 1205 7825 1240 7925
rect 1260 7825 1295 7925
rect 1455 7825 1490 7925
rect 1510 7825 1545 7925
rect 1705 7825 1740 7925
rect 1760 7825 1795 7925
rect 1955 7825 1990 7925
rect 2010 7825 2045 7925
rect 2205 7825 2240 7925
rect 2260 7825 2295 7925
rect 2455 7825 2490 7925
rect 2510 7825 2545 7925
rect 2705 7825 2740 7925
rect 2760 7825 2795 7925
rect 2955 7825 2990 7925
rect 3010 7825 3045 7925
rect 3205 7825 3240 7925
rect 3260 7825 3295 7925
rect 3455 7825 3490 7925
rect 3510 7825 3545 7925
rect 3705 7825 3740 7925
rect 3760 7825 3795 7925
rect 3955 7825 3990 7925
rect 4010 7825 4045 7925
rect 4205 7825 4240 7925
rect 4260 7825 4295 7925
rect 4455 7825 4490 7925
rect 4510 7825 4545 7925
rect 4705 7825 4740 7925
rect 4760 7825 4795 7925
rect 4955 7825 4990 7925
rect 5010 7825 5045 7925
rect 5205 7825 5240 7925
rect 5260 7825 5295 7925
rect 5455 7825 5490 7925
rect 5510 7825 5545 7925
rect 5705 7825 5740 7925
rect 5760 7825 5795 7925
rect 5955 7825 5990 7925
rect 6010 7825 6045 7925
rect 6205 7825 6240 7925
rect 6260 7825 6295 7925
rect 6455 7825 6490 7925
rect 6510 7825 6545 7925
rect 6705 7825 6740 7925
rect 6760 7825 6795 7925
rect 6955 7825 6990 7925
rect 7010 7825 7045 7925
rect 7205 7825 7240 7925
rect 7260 7825 7295 7925
rect 7455 7825 7490 7925
rect 7510 7825 7545 7925
rect 7705 7825 7740 7925
rect 7760 7825 7795 7925
rect 7955 7825 7990 7925
rect 75 7760 175 7795
rect 75 7705 175 7740
rect 325 7760 425 7795
rect 325 7705 425 7740
rect 575 7760 675 7795
rect 575 7705 675 7740
rect 825 7760 925 7795
rect 825 7705 925 7740
rect 1075 7760 1175 7795
rect 1075 7705 1175 7740
rect 1325 7760 1425 7795
rect 1325 7705 1425 7740
rect 1575 7760 1675 7795
rect 1575 7705 1675 7740
rect 1825 7760 1925 7795
rect 1825 7705 1925 7740
rect 2075 7760 2175 7795
rect 2075 7705 2175 7740
rect 2325 7760 2425 7795
rect 2325 7705 2425 7740
rect 2575 7760 2675 7795
rect 2575 7705 2675 7740
rect 2825 7760 2925 7795
rect 2825 7705 2925 7740
rect 3075 7760 3175 7795
rect 3075 7705 3175 7740
rect 3325 7760 3425 7795
rect 3325 7705 3425 7740
rect 3575 7760 3675 7795
rect 3575 7705 3675 7740
rect 3825 7760 3925 7795
rect 3825 7705 3925 7740
rect 4075 7760 4175 7795
rect 4075 7705 4175 7740
rect 4325 7760 4425 7795
rect 4325 7705 4425 7740
rect 4575 7760 4675 7795
rect 4575 7705 4675 7740
rect 4825 7760 4925 7795
rect 4825 7705 4925 7740
rect 5075 7760 5175 7795
rect 5075 7705 5175 7740
rect 5325 7760 5425 7795
rect 5325 7705 5425 7740
rect 5575 7760 5675 7795
rect 5575 7705 5675 7740
rect 5825 7760 5925 7795
rect 5825 7705 5925 7740
rect 6075 7760 6175 7795
rect 6075 7705 6175 7740
rect 6325 7760 6425 7795
rect 6325 7705 6425 7740
rect 6575 7760 6675 7795
rect 6575 7705 6675 7740
rect 6825 7760 6925 7795
rect 6825 7705 6925 7740
rect 7075 7760 7175 7795
rect 7075 7705 7175 7740
rect 7325 7760 7425 7795
rect 7325 7705 7425 7740
rect 7575 7760 7675 7795
rect 7575 7705 7675 7740
rect 7825 7760 7925 7795
rect 7825 7705 7925 7740
rect 10 7575 45 7675
rect 205 7575 240 7675
rect 260 7575 295 7675
rect 455 7575 490 7675
rect 510 7575 545 7675
rect 705 7575 740 7675
rect 760 7575 795 7675
rect 955 7575 990 7675
rect 1010 7575 1045 7675
rect 1205 7575 1240 7675
rect 1260 7575 1295 7675
rect 1455 7575 1490 7675
rect 1510 7575 1545 7675
rect 1705 7575 1740 7675
rect 1760 7575 1795 7675
rect 1955 7575 1990 7675
rect 2010 7575 2045 7675
rect 2205 7575 2240 7675
rect 2260 7575 2295 7675
rect 2455 7575 2490 7675
rect 2510 7575 2545 7675
rect 2705 7575 2740 7675
rect 2760 7575 2795 7675
rect 2955 7575 2990 7675
rect 3010 7575 3045 7675
rect 3205 7575 3240 7675
rect 3260 7575 3295 7675
rect 3455 7575 3490 7675
rect 3510 7575 3545 7675
rect 3705 7575 3740 7675
rect 3760 7575 3795 7675
rect 3955 7575 3990 7675
rect 4010 7575 4045 7675
rect 4205 7575 4240 7675
rect 4260 7575 4295 7675
rect 4455 7575 4490 7675
rect 4510 7575 4545 7675
rect 4705 7575 4740 7675
rect 4760 7575 4795 7675
rect 4955 7575 4990 7675
rect 5010 7575 5045 7675
rect 5205 7575 5240 7675
rect 5260 7575 5295 7675
rect 5455 7575 5490 7675
rect 5510 7575 5545 7675
rect 5705 7575 5740 7675
rect 5760 7575 5795 7675
rect 5955 7575 5990 7675
rect 6010 7575 6045 7675
rect 6205 7575 6240 7675
rect 6260 7575 6295 7675
rect 6455 7575 6490 7675
rect 6510 7575 6545 7675
rect 6705 7575 6740 7675
rect 6760 7575 6795 7675
rect 6955 7575 6990 7675
rect 7010 7575 7045 7675
rect 7205 7575 7240 7675
rect 7260 7575 7295 7675
rect 7455 7575 7490 7675
rect 7510 7575 7545 7675
rect 7705 7575 7740 7675
rect 7760 7575 7795 7675
rect 7955 7575 7990 7675
rect 75 7510 175 7545
rect 75 7455 175 7490
rect 325 7510 425 7545
rect 325 7455 425 7490
rect 575 7510 675 7545
rect 575 7455 675 7490
rect 825 7510 925 7545
rect 825 7455 925 7490
rect 1075 7510 1175 7545
rect 1075 7455 1175 7490
rect 1325 7510 1425 7545
rect 1325 7455 1425 7490
rect 1575 7510 1675 7545
rect 1575 7455 1675 7490
rect 1825 7510 1925 7545
rect 1825 7455 1925 7490
rect 2075 7510 2175 7545
rect 2075 7455 2175 7490
rect 2325 7510 2425 7545
rect 2325 7455 2425 7490
rect 2575 7510 2675 7545
rect 2575 7455 2675 7490
rect 2825 7510 2925 7545
rect 2825 7455 2925 7490
rect 3075 7510 3175 7545
rect 3075 7455 3175 7490
rect 3325 7510 3425 7545
rect 3325 7455 3425 7490
rect 3575 7510 3675 7545
rect 3575 7455 3675 7490
rect 3825 7510 3925 7545
rect 3825 7455 3925 7490
rect 4075 7510 4175 7545
rect 4075 7455 4175 7490
rect 4325 7510 4425 7545
rect 4325 7455 4425 7490
rect 4575 7510 4675 7545
rect 4575 7455 4675 7490
rect 4825 7510 4925 7545
rect 4825 7455 4925 7490
rect 5075 7510 5175 7545
rect 5075 7455 5175 7490
rect 5325 7510 5425 7545
rect 5325 7455 5425 7490
rect 5575 7510 5675 7545
rect 5575 7455 5675 7490
rect 5825 7510 5925 7545
rect 5825 7455 5925 7490
rect 6075 7510 6175 7545
rect 6075 7455 6175 7490
rect 6325 7510 6425 7545
rect 6325 7455 6425 7490
rect 6575 7510 6675 7545
rect 6575 7455 6675 7490
rect 6825 7510 6925 7545
rect 6825 7455 6925 7490
rect 7075 7510 7175 7545
rect 7075 7455 7175 7490
rect 7325 7510 7425 7545
rect 7325 7455 7425 7490
rect 7575 7510 7675 7545
rect 7575 7455 7675 7490
rect 7825 7510 7925 7545
rect 7825 7455 7925 7490
rect 10 7325 45 7425
rect 205 7325 240 7425
rect 260 7325 295 7425
rect 455 7325 490 7425
rect 510 7325 545 7425
rect 705 7325 740 7425
rect 760 7325 795 7425
rect 955 7325 990 7425
rect 1010 7325 1045 7425
rect 1205 7325 1240 7425
rect 1260 7325 1295 7425
rect 1455 7325 1490 7425
rect 1510 7325 1545 7425
rect 1705 7325 1740 7425
rect 1760 7325 1795 7425
rect 1955 7325 1990 7425
rect 2010 7325 2045 7425
rect 2205 7325 2240 7425
rect 2260 7325 2295 7425
rect 2455 7325 2490 7425
rect 2510 7325 2545 7425
rect 2705 7325 2740 7425
rect 2760 7325 2795 7425
rect 2955 7325 2990 7425
rect 3010 7325 3045 7425
rect 3205 7325 3240 7425
rect 3260 7325 3295 7425
rect 3455 7325 3490 7425
rect 3510 7325 3545 7425
rect 3705 7325 3740 7425
rect 3760 7325 3795 7425
rect 3955 7325 3990 7425
rect 4010 7325 4045 7425
rect 4205 7325 4240 7425
rect 4260 7325 4295 7425
rect 4455 7325 4490 7425
rect 4510 7325 4545 7425
rect 4705 7325 4740 7425
rect 4760 7325 4795 7425
rect 4955 7325 4990 7425
rect 5010 7325 5045 7425
rect 5205 7325 5240 7425
rect 5260 7325 5295 7425
rect 5455 7325 5490 7425
rect 5510 7325 5545 7425
rect 5705 7325 5740 7425
rect 5760 7325 5795 7425
rect 5955 7325 5990 7425
rect 6010 7325 6045 7425
rect 6205 7325 6240 7425
rect 6260 7325 6295 7425
rect 6455 7325 6490 7425
rect 6510 7325 6545 7425
rect 6705 7325 6740 7425
rect 6760 7325 6795 7425
rect 6955 7325 6990 7425
rect 7010 7325 7045 7425
rect 7205 7325 7240 7425
rect 7260 7325 7295 7425
rect 7455 7325 7490 7425
rect 7510 7325 7545 7425
rect 7705 7325 7740 7425
rect 7760 7325 7795 7425
rect 7955 7325 7990 7425
rect 75 7260 175 7295
rect 75 7205 175 7240
rect 325 7260 425 7295
rect 325 7205 425 7240
rect 575 7260 675 7295
rect 575 7205 675 7240
rect 825 7260 925 7295
rect 825 7205 925 7240
rect 1075 7260 1175 7295
rect 1075 7205 1175 7240
rect 1325 7260 1425 7295
rect 1325 7205 1425 7240
rect 1575 7260 1675 7295
rect 1575 7205 1675 7240
rect 1825 7260 1925 7295
rect 1825 7205 1925 7240
rect 2075 7260 2175 7295
rect 2075 7205 2175 7240
rect 2325 7260 2425 7295
rect 2325 7205 2425 7240
rect 2575 7260 2675 7295
rect 2575 7205 2675 7240
rect 2825 7260 2925 7295
rect 2825 7205 2925 7240
rect 3075 7260 3175 7295
rect 3075 7205 3175 7240
rect 3325 7260 3425 7295
rect 3325 7205 3425 7240
rect 3575 7260 3675 7295
rect 3575 7205 3675 7240
rect 3825 7260 3925 7295
rect 3825 7205 3925 7240
rect 4075 7260 4175 7295
rect 4075 7205 4175 7240
rect 4325 7260 4425 7295
rect 4325 7205 4425 7240
rect 4575 7260 4675 7295
rect 4575 7205 4675 7240
rect 4825 7260 4925 7295
rect 4825 7205 4925 7240
rect 5075 7260 5175 7295
rect 5075 7205 5175 7240
rect 5325 7260 5425 7295
rect 5325 7205 5425 7240
rect 5575 7260 5675 7295
rect 5575 7205 5675 7240
rect 5825 7260 5925 7295
rect 5825 7205 5925 7240
rect 6075 7260 6175 7295
rect 6075 7205 6175 7240
rect 6325 7260 6425 7295
rect 6325 7205 6425 7240
rect 6575 7260 6675 7295
rect 6575 7205 6675 7240
rect 6825 7260 6925 7295
rect 6825 7205 6925 7240
rect 7075 7260 7175 7295
rect 7075 7205 7175 7240
rect 7325 7260 7425 7295
rect 7325 7205 7425 7240
rect 7575 7260 7675 7295
rect 7575 7205 7675 7240
rect 7825 7260 7925 7295
rect 7825 7205 7925 7240
rect 10 7075 45 7175
rect 205 7075 240 7175
rect 260 7075 295 7175
rect 455 7075 490 7175
rect 510 7075 545 7175
rect 705 7075 740 7175
rect 760 7075 795 7175
rect 955 7075 990 7175
rect 1010 7075 1045 7175
rect 1205 7075 1240 7175
rect 1260 7075 1295 7175
rect 1455 7075 1490 7175
rect 1510 7075 1545 7175
rect 1705 7075 1740 7175
rect 1760 7075 1795 7175
rect 1955 7075 1990 7175
rect 2010 7075 2045 7175
rect 2205 7075 2240 7175
rect 2260 7075 2295 7175
rect 2455 7075 2490 7175
rect 2510 7075 2545 7175
rect 2705 7075 2740 7175
rect 2760 7075 2795 7175
rect 2955 7075 2990 7175
rect 3010 7075 3045 7175
rect 3205 7075 3240 7175
rect 3260 7075 3295 7175
rect 3455 7075 3490 7175
rect 3510 7075 3545 7175
rect 3705 7075 3740 7175
rect 3760 7075 3795 7175
rect 3955 7075 3990 7175
rect 4010 7075 4045 7175
rect 4205 7075 4240 7175
rect 4260 7075 4295 7175
rect 4455 7075 4490 7175
rect 4510 7075 4545 7175
rect 4705 7075 4740 7175
rect 4760 7075 4795 7175
rect 4955 7075 4990 7175
rect 5010 7075 5045 7175
rect 5205 7075 5240 7175
rect 5260 7075 5295 7175
rect 5455 7075 5490 7175
rect 5510 7075 5545 7175
rect 5705 7075 5740 7175
rect 5760 7075 5795 7175
rect 5955 7075 5990 7175
rect 6010 7075 6045 7175
rect 6205 7075 6240 7175
rect 6260 7075 6295 7175
rect 6455 7075 6490 7175
rect 6510 7075 6545 7175
rect 6705 7075 6740 7175
rect 6760 7075 6795 7175
rect 6955 7075 6990 7175
rect 7010 7075 7045 7175
rect 7205 7075 7240 7175
rect 7260 7075 7295 7175
rect 7455 7075 7490 7175
rect 7510 7075 7545 7175
rect 7705 7075 7740 7175
rect 7760 7075 7795 7175
rect 7955 7075 7990 7175
rect 75 7010 175 7045
rect 75 6955 175 6990
rect 325 7010 425 7045
rect 325 6955 425 6990
rect 575 7010 675 7045
rect 575 6955 675 6990
rect 825 7010 925 7045
rect 825 6955 925 6990
rect 1075 7010 1175 7045
rect 1075 6955 1175 6990
rect 1325 7010 1425 7045
rect 1325 6955 1425 6990
rect 1575 7010 1675 7045
rect 1575 6955 1675 6990
rect 1825 7010 1925 7045
rect 1825 6955 1925 6990
rect 2075 7010 2175 7045
rect 2075 6955 2175 6990
rect 2325 7010 2425 7045
rect 2325 6955 2425 6990
rect 2575 7010 2675 7045
rect 2575 6955 2675 6990
rect 2825 7010 2925 7045
rect 2825 6955 2925 6990
rect 3075 7010 3175 7045
rect 3075 6955 3175 6990
rect 3325 7010 3425 7045
rect 3325 6955 3425 6990
rect 3575 7010 3675 7045
rect 3575 6955 3675 6990
rect 3825 7010 3925 7045
rect 3825 6955 3925 6990
rect 4075 7010 4175 7045
rect 4075 6955 4175 6990
rect 4325 7010 4425 7045
rect 4325 6955 4425 6990
rect 4575 7010 4675 7045
rect 4575 6955 4675 6990
rect 4825 7010 4925 7045
rect 4825 6955 4925 6990
rect 5075 7010 5175 7045
rect 5075 6955 5175 6990
rect 5325 7010 5425 7045
rect 5325 6955 5425 6990
rect 5575 7010 5675 7045
rect 5575 6955 5675 6990
rect 5825 7010 5925 7045
rect 5825 6955 5925 6990
rect 6075 7010 6175 7045
rect 6075 6955 6175 6990
rect 6325 7010 6425 7045
rect 6325 6955 6425 6990
rect 6575 7010 6675 7045
rect 6575 6955 6675 6990
rect 6825 7010 6925 7045
rect 6825 6955 6925 6990
rect 7075 7010 7175 7045
rect 7075 6955 7175 6990
rect 7325 7010 7425 7045
rect 7325 6955 7425 6990
rect 7575 7010 7675 7045
rect 7575 6955 7675 6990
rect 7825 7010 7925 7045
rect 7825 6955 7925 6990
rect 10 6825 45 6925
rect 205 6825 240 6925
rect 260 6825 295 6925
rect 455 6825 490 6925
rect 510 6825 545 6925
rect 705 6825 740 6925
rect 760 6825 795 6925
rect 955 6825 990 6925
rect 1010 6825 1045 6925
rect 1205 6825 1240 6925
rect 1260 6825 1295 6925
rect 1455 6825 1490 6925
rect 1510 6825 1545 6925
rect 1705 6825 1740 6925
rect 1760 6825 1795 6925
rect 1955 6825 1990 6925
rect 2010 6825 2045 6925
rect 2205 6825 2240 6925
rect 2260 6825 2295 6925
rect 2455 6825 2490 6925
rect 2510 6825 2545 6925
rect 2705 6825 2740 6925
rect 2760 6825 2795 6925
rect 2955 6825 2990 6925
rect 3010 6825 3045 6925
rect 3205 6825 3240 6925
rect 3260 6825 3295 6925
rect 3455 6825 3490 6925
rect 3510 6825 3545 6925
rect 3705 6825 3740 6925
rect 3760 6825 3795 6925
rect 3955 6825 3990 6925
rect 4010 6825 4045 6925
rect 4205 6825 4240 6925
rect 4260 6825 4295 6925
rect 4455 6825 4490 6925
rect 4510 6825 4545 6925
rect 4705 6825 4740 6925
rect 4760 6825 4795 6925
rect 4955 6825 4990 6925
rect 5010 6825 5045 6925
rect 5205 6825 5240 6925
rect 5260 6825 5295 6925
rect 5455 6825 5490 6925
rect 5510 6825 5545 6925
rect 5705 6825 5740 6925
rect 5760 6825 5795 6925
rect 5955 6825 5990 6925
rect 6010 6825 6045 6925
rect 6205 6825 6240 6925
rect 6260 6825 6295 6925
rect 6455 6825 6490 6925
rect 6510 6825 6545 6925
rect 6705 6825 6740 6925
rect 6760 6825 6795 6925
rect 6955 6825 6990 6925
rect 7010 6825 7045 6925
rect 7205 6825 7240 6925
rect 7260 6825 7295 6925
rect 7455 6825 7490 6925
rect 7510 6825 7545 6925
rect 7705 6825 7740 6925
rect 7760 6825 7795 6925
rect 7955 6825 7990 6925
rect 75 6760 175 6795
rect 75 6705 175 6740
rect 325 6760 425 6795
rect 325 6705 425 6740
rect 575 6760 675 6795
rect 575 6705 675 6740
rect 825 6760 925 6795
rect 825 6705 925 6740
rect 1075 6760 1175 6795
rect 1075 6705 1175 6740
rect 1325 6760 1425 6795
rect 1325 6705 1425 6740
rect 1575 6760 1675 6795
rect 1575 6705 1675 6740
rect 1825 6760 1925 6795
rect 1825 6705 1925 6740
rect 2075 6760 2175 6795
rect 2075 6705 2175 6740
rect 2325 6760 2425 6795
rect 2325 6705 2425 6740
rect 2575 6760 2675 6795
rect 2575 6705 2675 6740
rect 2825 6760 2925 6795
rect 2825 6705 2925 6740
rect 3075 6760 3175 6795
rect 3075 6705 3175 6740
rect 3325 6760 3425 6795
rect 3325 6705 3425 6740
rect 3575 6760 3675 6795
rect 3575 6705 3675 6740
rect 3825 6760 3925 6795
rect 3825 6705 3925 6740
rect 4075 6760 4175 6795
rect 4075 6705 4175 6740
rect 4325 6760 4425 6795
rect 4325 6705 4425 6740
rect 4575 6760 4675 6795
rect 4575 6705 4675 6740
rect 4825 6760 4925 6795
rect 4825 6705 4925 6740
rect 5075 6760 5175 6795
rect 5075 6705 5175 6740
rect 5325 6760 5425 6795
rect 5325 6705 5425 6740
rect 5575 6760 5675 6795
rect 5575 6705 5675 6740
rect 5825 6760 5925 6795
rect 5825 6705 5925 6740
rect 6075 6760 6175 6795
rect 6075 6705 6175 6740
rect 6325 6760 6425 6795
rect 6325 6705 6425 6740
rect 6575 6760 6675 6795
rect 6575 6705 6675 6740
rect 6825 6760 6925 6795
rect 6825 6705 6925 6740
rect 7075 6760 7175 6795
rect 7075 6705 7175 6740
rect 7325 6760 7425 6795
rect 7325 6705 7425 6740
rect 7575 6760 7675 6795
rect 7575 6705 7675 6740
rect 7825 6760 7925 6795
rect 7825 6705 7925 6740
rect 10 6575 45 6675
rect 205 6575 240 6675
rect 260 6575 295 6675
rect 455 6575 490 6675
rect 510 6575 545 6675
rect 705 6575 740 6675
rect 760 6575 795 6675
rect 955 6575 990 6675
rect 1010 6575 1045 6675
rect 1205 6575 1240 6675
rect 1260 6575 1295 6675
rect 1455 6575 1490 6675
rect 1510 6575 1545 6675
rect 1705 6575 1740 6675
rect 1760 6575 1795 6675
rect 1955 6575 1990 6675
rect 2010 6575 2045 6675
rect 2205 6575 2240 6675
rect 2260 6575 2295 6675
rect 2455 6575 2490 6675
rect 2510 6575 2545 6675
rect 2705 6575 2740 6675
rect 2760 6575 2795 6675
rect 2955 6575 2990 6675
rect 3010 6575 3045 6675
rect 3205 6575 3240 6675
rect 3260 6575 3295 6675
rect 3455 6575 3490 6675
rect 3510 6575 3545 6675
rect 3705 6575 3740 6675
rect 3760 6575 3795 6675
rect 3955 6575 3990 6675
rect 4010 6575 4045 6675
rect 4205 6575 4240 6675
rect 4260 6575 4295 6675
rect 4455 6575 4490 6675
rect 4510 6575 4545 6675
rect 4705 6575 4740 6675
rect 4760 6575 4795 6675
rect 4955 6575 4990 6675
rect 5010 6575 5045 6675
rect 5205 6575 5240 6675
rect 5260 6575 5295 6675
rect 5455 6575 5490 6675
rect 5510 6575 5545 6675
rect 5705 6575 5740 6675
rect 5760 6575 5795 6675
rect 5955 6575 5990 6675
rect 6010 6575 6045 6675
rect 6205 6575 6240 6675
rect 6260 6575 6295 6675
rect 6455 6575 6490 6675
rect 6510 6575 6545 6675
rect 6705 6575 6740 6675
rect 6760 6575 6795 6675
rect 6955 6575 6990 6675
rect 7010 6575 7045 6675
rect 7205 6575 7240 6675
rect 7260 6575 7295 6675
rect 7455 6575 7490 6675
rect 7510 6575 7545 6675
rect 7705 6575 7740 6675
rect 7760 6575 7795 6675
rect 7955 6575 7990 6675
rect 75 6510 175 6545
rect 75 6455 175 6490
rect 325 6510 425 6545
rect 325 6455 425 6490
rect 575 6510 675 6545
rect 575 6455 675 6490
rect 825 6510 925 6545
rect 825 6455 925 6490
rect 1075 6510 1175 6545
rect 1075 6455 1175 6490
rect 1325 6510 1425 6545
rect 1325 6455 1425 6490
rect 1575 6510 1675 6545
rect 1575 6455 1675 6490
rect 1825 6510 1925 6545
rect 1825 6455 1925 6490
rect 2075 6510 2175 6545
rect 2075 6455 2175 6490
rect 2325 6510 2425 6545
rect 2325 6455 2425 6490
rect 2575 6510 2675 6545
rect 2575 6455 2675 6490
rect 2825 6510 2925 6545
rect 2825 6455 2925 6490
rect 3075 6510 3175 6545
rect 3075 6455 3175 6490
rect 3325 6510 3425 6545
rect 3325 6455 3425 6490
rect 3575 6510 3675 6545
rect 3575 6455 3675 6490
rect 3825 6510 3925 6545
rect 3825 6455 3925 6490
rect 4075 6510 4175 6545
rect 4075 6455 4175 6490
rect 4325 6510 4425 6545
rect 4325 6455 4425 6490
rect 4575 6510 4675 6545
rect 4575 6455 4675 6490
rect 4825 6510 4925 6545
rect 4825 6455 4925 6490
rect 5075 6510 5175 6545
rect 5075 6455 5175 6490
rect 5325 6510 5425 6545
rect 5325 6455 5425 6490
rect 5575 6510 5675 6545
rect 5575 6455 5675 6490
rect 5825 6510 5925 6545
rect 5825 6455 5925 6490
rect 6075 6510 6175 6545
rect 6075 6455 6175 6490
rect 6325 6510 6425 6545
rect 6325 6455 6425 6490
rect 6575 6510 6675 6545
rect 6575 6455 6675 6490
rect 6825 6510 6925 6545
rect 6825 6455 6925 6490
rect 7075 6510 7175 6545
rect 7075 6455 7175 6490
rect 7325 6510 7425 6545
rect 7325 6455 7425 6490
rect 7575 6510 7675 6545
rect 7575 6455 7675 6490
rect 7825 6510 7925 6545
rect 7825 6455 7925 6490
rect 10 6325 45 6425
rect 205 6325 240 6425
rect 260 6325 295 6425
rect 455 6325 490 6425
rect 510 6325 545 6425
rect 705 6325 740 6425
rect 760 6325 795 6425
rect 955 6325 990 6425
rect 1010 6325 1045 6425
rect 1205 6325 1240 6425
rect 1260 6325 1295 6425
rect 1455 6325 1490 6425
rect 1510 6325 1545 6425
rect 1705 6325 1740 6425
rect 1760 6325 1795 6425
rect 1955 6325 1990 6425
rect 2010 6325 2045 6425
rect 2205 6325 2240 6425
rect 2260 6325 2295 6425
rect 2455 6325 2490 6425
rect 2510 6325 2545 6425
rect 2705 6325 2740 6425
rect 2760 6325 2795 6425
rect 2955 6325 2990 6425
rect 3010 6325 3045 6425
rect 3205 6325 3240 6425
rect 3260 6325 3295 6425
rect 3455 6325 3490 6425
rect 3510 6325 3545 6425
rect 3705 6325 3740 6425
rect 3760 6325 3795 6425
rect 3955 6325 3990 6425
rect 4010 6325 4045 6425
rect 4205 6325 4240 6425
rect 4260 6325 4295 6425
rect 4455 6325 4490 6425
rect 4510 6325 4545 6425
rect 4705 6325 4740 6425
rect 4760 6325 4795 6425
rect 4955 6325 4990 6425
rect 5010 6325 5045 6425
rect 5205 6325 5240 6425
rect 5260 6325 5295 6425
rect 5455 6325 5490 6425
rect 5510 6325 5545 6425
rect 5705 6325 5740 6425
rect 5760 6325 5795 6425
rect 5955 6325 5990 6425
rect 6010 6325 6045 6425
rect 6205 6325 6240 6425
rect 6260 6325 6295 6425
rect 6455 6325 6490 6425
rect 6510 6325 6545 6425
rect 6705 6325 6740 6425
rect 6760 6325 6795 6425
rect 6955 6325 6990 6425
rect 7010 6325 7045 6425
rect 7205 6325 7240 6425
rect 7260 6325 7295 6425
rect 7455 6325 7490 6425
rect 7510 6325 7545 6425
rect 7705 6325 7740 6425
rect 7760 6325 7795 6425
rect 7955 6325 7990 6425
rect 75 6260 175 6295
rect 75 6205 175 6240
rect 325 6260 425 6295
rect 325 6205 425 6240
rect 575 6260 675 6295
rect 575 6205 675 6240
rect 825 6260 925 6295
rect 825 6205 925 6240
rect 1075 6260 1175 6295
rect 1075 6205 1175 6240
rect 1325 6260 1425 6295
rect 1325 6205 1425 6240
rect 1575 6260 1675 6295
rect 1575 6205 1675 6240
rect 1825 6260 1925 6295
rect 1825 6205 1925 6240
rect 2075 6260 2175 6295
rect 2075 6205 2175 6240
rect 2325 6260 2425 6295
rect 2325 6205 2425 6240
rect 2575 6260 2675 6295
rect 2575 6205 2675 6240
rect 2825 6260 2925 6295
rect 2825 6205 2925 6240
rect 3075 6260 3175 6295
rect 3075 6205 3175 6240
rect 3325 6260 3425 6295
rect 3325 6205 3425 6240
rect 3575 6260 3675 6295
rect 3575 6205 3675 6240
rect 3825 6260 3925 6295
rect 3825 6205 3925 6240
rect 4075 6260 4175 6295
rect 4075 6205 4175 6240
rect 4325 6260 4425 6295
rect 4325 6205 4425 6240
rect 4575 6260 4675 6295
rect 4575 6205 4675 6240
rect 4825 6260 4925 6295
rect 4825 6205 4925 6240
rect 5075 6260 5175 6295
rect 5075 6205 5175 6240
rect 5325 6260 5425 6295
rect 5325 6205 5425 6240
rect 5575 6260 5675 6295
rect 5575 6205 5675 6240
rect 5825 6260 5925 6295
rect 5825 6205 5925 6240
rect 6075 6260 6175 6295
rect 6075 6205 6175 6240
rect 6325 6260 6425 6295
rect 6325 6205 6425 6240
rect 6575 6260 6675 6295
rect 6575 6205 6675 6240
rect 6825 6260 6925 6295
rect 6825 6205 6925 6240
rect 7075 6260 7175 6295
rect 7075 6205 7175 6240
rect 7325 6260 7425 6295
rect 7325 6205 7425 6240
rect 7575 6260 7675 6295
rect 7575 6205 7675 6240
rect 7825 6260 7925 6295
rect 7825 6205 7925 6240
rect 10 6075 45 6175
rect 205 6075 240 6175
rect 260 6075 295 6175
rect 455 6075 490 6175
rect 510 6075 545 6175
rect 705 6075 740 6175
rect 760 6075 795 6175
rect 955 6075 990 6175
rect 1010 6075 1045 6175
rect 1205 6075 1240 6175
rect 1260 6075 1295 6175
rect 1455 6075 1490 6175
rect 1510 6075 1545 6175
rect 1705 6075 1740 6175
rect 1760 6075 1795 6175
rect 1955 6075 1990 6175
rect 2010 6075 2045 6175
rect 2205 6075 2240 6175
rect 2260 6075 2295 6175
rect 2455 6075 2490 6175
rect 2510 6075 2545 6175
rect 2705 6075 2740 6175
rect 2760 6075 2795 6175
rect 2955 6075 2990 6175
rect 3010 6075 3045 6175
rect 3205 6075 3240 6175
rect 3260 6075 3295 6175
rect 3455 6075 3490 6175
rect 3510 6075 3545 6175
rect 3705 6075 3740 6175
rect 3760 6075 3795 6175
rect 3955 6075 3990 6175
rect 4010 6075 4045 6175
rect 4205 6075 4240 6175
rect 4260 6075 4295 6175
rect 4455 6075 4490 6175
rect 4510 6075 4545 6175
rect 4705 6075 4740 6175
rect 4760 6075 4795 6175
rect 4955 6075 4990 6175
rect 5010 6075 5045 6175
rect 5205 6075 5240 6175
rect 5260 6075 5295 6175
rect 5455 6075 5490 6175
rect 5510 6075 5545 6175
rect 5705 6075 5740 6175
rect 5760 6075 5795 6175
rect 5955 6075 5990 6175
rect 6010 6075 6045 6175
rect 6205 6075 6240 6175
rect 6260 6075 6295 6175
rect 6455 6075 6490 6175
rect 6510 6075 6545 6175
rect 6705 6075 6740 6175
rect 6760 6075 6795 6175
rect 6955 6075 6990 6175
rect 7010 6075 7045 6175
rect 7205 6075 7240 6175
rect 7260 6075 7295 6175
rect 7455 6075 7490 6175
rect 7510 6075 7545 6175
rect 7705 6075 7740 6175
rect 7760 6075 7795 6175
rect 7955 6075 7990 6175
rect 75 6010 175 6045
rect 75 5955 175 5990
rect 325 6010 425 6045
rect 325 5955 425 5990
rect 575 6010 675 6045
rect 575 5955 675 5990
rect 825 6010 925 6045
rect 825 5955 925 5990
rect 1075 6010 1175 6045
rect 1075 5955 1175 5990
rect 1325 6010 1425 6045
rect 1325 5955 1425 5990
rect 1575 6010 1675 6045
rect 1575 5955 1675 5990
rect 1825 6010 1925 6045
rect 1825 5955 1925 5990
rect 2075 6010 2175 6045
rect 2075 5955 2175 5990
rect 2325 6010 2425 6045
rect 2325 5955 2425 5990
rect 2575 6010 2675 6045
rect 2575 5955 2675 5990
rect 2825 6010 2925 6045
rect 2825 5955 2925 5990
rect 3075 6010 3175 6045
rect 3075 5955 3175 5990
rect 3325 6010 3425 6045
rect 3325 5955 3425 5990
rect 3575 6010 3675 6045
rect 3575 5955 3675 5990
rect 3825 6010 3925 6045
rect 3825 5955 3925 5990
rect 4075 6010 4175 6045
rect 4075 5955 4175 5990
rect 4325 6010 4425 6045
rect 4325 5955 4425 5990
rect 4575 6010 4675 6045
rect 4575 5955 4675 5990
rect 4825 6010 4925 6045
rect 4825 5955 4925 5990
rect 5075 6010 5175 6045
rect 5075 5955 5175 5990
rect 5325 6010 5425 6045
rect 5325 5955 5425 5990
rect 5575 6010 5675 6045
rect 5575 5955 5675 5990
rect 5825 6010 5925 6045
rect 5825 5955 5925 5990
rect 6075 6010 6175 6045
rect 6075 5955 6175 5990
rect 6325 6010 6425 6045
rect 6325 5955 6425 5990
rect 6575 6010 6675 6045
rect 6575 5955 6675 5990
rect 6825 6010 6925 6045
rect 6825 5955 6925 5990
rect 7075 6010 7175 6045
rect 7075 5955 7175 5990
rect 7325 6010 7425 6045
rect 7325 5955 7425 5990
rect 7575 6010 7675 6045
rect 7575 5955 7675 5990
rect 7825 6010 7925 6045
rect 7825 5955 7925 5990
rect 10 5825 45 5925
rect 205 5825 240 5925
rect 260 5825 295 5925
rect 455 5825 490 5925
rect 510 5825 545 5925
rect 705 5825 740 5925
rect 760 5825 795 5925
rect 955 5825 990 5925
rect 1010 5825 1045 5925
rect 1205 5825 1240 5925
rect 1260 5825 1295 5925
rect 1455 5825 1490 5925
rect 1510 5825 1545 5925
rect 1705 5825 1740 5925
rect 1760 5825 1795 5925
rect 1955 5825 1990 5925
rect 2010 5825 2045 5925
rect 2205 5825 2240 5925
rect 2260 5825 2295 5925
rect 2455 5825 2490 5925
rect 2510 5825 2545 5925
rect 2705 5825 2740 5925
rect 2760 5825 2795 5925
rect 2955 5825 2990 5925
rect 3010 5825 3045 5925
rect 3205 5825 3240 5925
rect 3260 5825 3295 5925
rect 3455 5825 3490 5925
rect 3510 5825 3545 5925
rect 3705 5825 3740 5925
rect 3760 5825 3795 5925
rect 3955 5825 3990 5925
rect 4010 5825 4045 5925
rect 4205 5825 4240 5925
rect 4260 5825 4295 5925
rect 4455 5825 4490 5925
rect 4510 5825 4545 5925
rect 4705 5825 4740 5925
rect 4760 5825 4795 5925
rect 4955 5825 4990 5925
rect 5010 5825 5045 5925
rect 5205 5825 5240 5925
rect 5260 5825 5295 5925
rect 5455 5825 5490 5925
rect 5510 5825 5545 5925
rect 5705 5825 5740 5925
rect 5760 5825 5795 5925
rect 5955 5825 5990 5925
rect 6010 5825 6045 5925
rect 6205 5825 6240 5925
rect 6260 5825 6295 5925
rect 6455 5825 6490 5925
rect 6510 5825 6545 5925
rect 6705 5825 6740 5925
rect 6760 5825 6795 5925
rect 6955 5825 6990 5925
rect 7010 5825 7045 5925
rect 7205 5825 7240 5925
rect 7260 5825 7295 5925
rect 7455 5825 7490 5925
rect 7510 5825 7545 5925
rect 7705 5825 7740 5925
rect 7760 5825 7795 5925
rect 7955 5825 7990 5925
rect 75 5760 175 5795
rect 75 5705 175 5740
rect 325 5760 425 5795
rect 325 5705 425 5740
rect 575 5760 675 5795
rect 575 5705 675 5740
rect 825 5760 925 5795
rect 825 5705 925 5740
rect 1075 5760 1175 5795
rect 1075 5705 1175 5740
rect 1325 5760 1425 5795
rect 1325 5705 1425 5740
rect 1575 5760 1675 5795
rect 1575 5705 1675 5740
rect 1825 5760 1925 5795
rect 1825 5705 1925 5740
rect 2075 5760 2175 5795
rect 2075 5705 2175 5740
rect 2325 5760 2425 5795
rect 2325 5705 2425 5740
rect 2575 5760 2675 5795
rect 2575 5705 2675 5740
rect 2825 5760 2925 5795
rect 2825 5705 2925 5740
rect 3075 5760 3175 5795
rect 3075 5705 3175 5740
rect 3325 5760 3425 5795
rect 3325 5705 3425 5740
rect 3575 5760 3675 5795
rect 3575 5705 3675 5740
rect 3825 5760 3925 5795
rect 3825 5705 3925 5740
rect 4075 5760 4175 5795
rect 4075 5705 4175 5740
rect 4325 5760 4425 5795
rect 4325 5705 4425 5740
rect 4575 5760 4675 5795
rect 4575 5705 4675 5740
rect 4825 5760 4925 5795
rect 4825 5705 4925 5740
rect 5075 5760 5175 5795
rect 5075 5705 5175 5740
rect 5325 5760 5425 5795
rect 5325 5705 5425 5740
rect 5575 5760 5675 5795
rect 5575 5705 5675 5740
rect 5825 5760 5925 5795
rect 5825 5705 5925 5740
rect 6075 5760 6175 5795
rect 6075 5705 6175 5740
rect 6325 5760 6425 5795
rect 6325 5705 6425 5740
rect 6575 5760 6675 5795
rect 6575 5705 6675 5740
rect 6825 5760 6925 5795
rect 6825 5705 6925 5740
rect 7075 5760 7175 5795
rect 7075 5705 7175 5740
rect 7325 5760 7425 5795
rect 7325 5705 7425 5740
rect 7575 5760 7675 5795
rect 7575 5705 7675 5740
rect 7825 5760 7925 5795
rect 7825 5705 7925 5740
rect 10 5575 45 5675
rect 205 5575 240 5675
rect 260 5575 295 5675
rect 455 5575 490 5675
rect 510 5575 545 5675
rect 705 5575 740 5675
rect 760 5575 795 5675
rect 955 5575 990 5675
rect 1010 5575 1045 5675
rect 1205 5575 1240 5675
rect 1260 5575 1295 5675
rect 1455 5575 1490 5675
rect 1510 5575 1545 5675
rect 1705 5575 1740 5675
rect 1760 5575 1795 5675
rect 1955 5575 1990 5675
rect 2010 5575 2045 5675
rect 2205 5575 2240 5675
rect 2260 5575 2295 5675
rect 2455 5575 2490 5675
rect 2510 5575 2545 5675
rect 2705 5575 2740 5675
rect 2760 5575 2795 5675
rect 2955 5575 2990 5675
rect 3010 5575 3045 5675
rect 3205 5575 3240 5675
rect 3260 5575 3295 5675
rect 3455 5575 3490 5675
rect 3510 5575 3545 5675
rect 3705 5575 3740 5675
rect 3760 5575 3795 5675
rect 3955 5575 3990 5675
rect 4010 5575 4045 5675
rect 4205 5575 4240 5675
rect 4260 5575 4295 5675
rect 4455 5575 4490 5675
rect 4510 5575 4545 5675
rect 4705 5575 4740 5675
rect 4760 5575 4795 5675
rect 4955 5575 4990 5675
rect 5010 5575 5045 5675
rect 5205 5575 5240 5675
rect 5260 5575 5295 5675
rect 5455 5575 5490 5675
rect 5510 5575 5545 5675
rect 5705 5575 5740 5675
rect 5760 5575 5795 5675
rect 5955 5575 5990 5675
rect 6010 5575 6045 5675
rect 6205 5575 6240 5675
rect 6260 5575 6295 5675
rect 6455 5575 6490 5675
rect 6510 5575 6545 5675
rect 6705 5575 6740 5675
rect 6760 5575 6795 5675
rect 6955 5575 6990 5675
rect 7010 5575 7045 5675
rect 7205 5575 7240 5675
rect 7260 5575 7295 5675
rect 7455 5575 7490 5675
rect 7510 5575 7545 5675
rect 7705 5575 7740 5675
rect 7760 5575 7795 5675
rect 7955 5575 7990 5675
rect 75 5510 175 5545
rect 75 5455 175 5490
rect 325 5510 425 5545
rect 325 5455 425 5490
rect 575 5510 675 5545
rect 575 5455 675 5490
rect 825 5510 925 5545
rect 825 5455 925 5490
rect 1075 5510 1175 5545
rect 1075 5455 1175 5490
rect 1325 5510 1425 5545
rect 1325 5455 1425 5490
rect 1575 5510 1675 5545
rect 1575 5455 1675 5490
rect 1825 5510 1925 5545
rect 1825 5455 1925 5490
rect 2075 5510 2175 5545
rect 2075 5455 2175 5490
rect 2325 5510 2425 5545
rect 2325 5455 2425 5490
rect 2575 5510 2675 5545
rect 2575 5455 2675 5490
rect 2825 5510 2925 5545
rect 2825 5455 2925 5490
rect 3075 5510 3175 5545
rect 3075 5455 3175 5490
rect 3325 5510 3425 5545
rect 3325 5455 3425 5490
rect 3575 5510 3675 5545
rect 3575 5455 3675 5490
rect 3825 5510 3925 5545
rect 3825 5455 3925 5490
rect 4075 5510 4175 5545
rect 4075 5455 4175 5490
rect 4325 5510 4425 5545
rect 4325 5455 4425 5490
rect 4575 5510 4675 5545
rect 4575 5455 4675 5490
rect 4825 5510 4925 5545
rect 4825 5455 4925 5490
rect 5075 5510 5175 5545
rect 5075 5455 5175 5490
rect 5325 5510 5425 5545
rect 5325 5455 5425 5490
rect 5575 5510 5675 5545
rect 5575 5455 5675 5490
rect 5825 5510 5925 5545
rect 5825 5455 5925 5490
rect 6075 5510 6175 5545
rect 6075 5455 6175 5490
rect 6325 5510 6425 5545
rect 6325 5455 6425 5490
rect 6575 5510 6675 5545
rect 6575 5455 6675 5490
rect 6825 5510 6925 5545
rect 6825 5455 6925 5490
rect 7075 5510 7175 5545
rect 7075 5455 7175 5490
rect 7325 5510 7425 5545
rect 7325 5455 7425 5490
rect 7575 5510 7675 5545
rect 7575 5455 7675 5490
rect 7825 5510 7925 5545
rect 7825 5455 7925 5490
rect 10 5325 45 5425
rect 205 5325 240 5425
rect 260 5325 295 5425
rect 455 5325 490 5425
rect 510 5325 545 5425
rect 705 5325 740 5425
rect 760 5325 795 5425
rect 955 5325 990 5425
rect 1010 5325 1045 5425
rect 1205 5325 1240 5425
rect 1260 5325 1295 5425
rect 1455 5325 1490 5425
rect 1510 5325 1545 5425
rect 1705 5325 1740 5425
rect 1760 5325 1795 5425
rect 1955 5325 1990 5425
rect 2010 5325 2045 5425
rect 2205 5325 2240 5425
rect 2260 5325 2295 5425
rect 2455 5325 2490 5425
rect 2510 5325 2545 5425
rect 2705 5325 2740 5425
rect 2760 5325 2795 5425
rect 2955 5325 2990 5425
rect 3010 5325 3045 5425
rect 3205 5325 3240 5425
rect 3260 5325 3295 5425
rect 3455 5325 3490 5425
rect 3510 5325 3545 5425
rect 3705 5325 3740 5425
rect 3760 5325 3795 5425
rect 3955 5325 3990 5425
rect 4010 5325 4045 5425
rect 4205 5325 4240 5425
rect 4260 5325 4295 5425
rect 4455 5325 4490 5425
rect 4510 5325 4545 5425
rect 4705 5325 4740 5425
rect 4760 5325 4795 5425
rect 4955 5325 4990 5425
rect 5010 5325 5045 5425
rect 5205 5325 5240 5425
rect 5260 5325 5295 5425
rect 5455 5325 5490 5425
rect 5510 5325 5545 5425
rect 5705 5325 5740 5425
rect 5760 5325 5795 5425
rect 5955 5325 5990 5425
rect 6010 5325 6045 5425
rect 6205 5325 6240 5425
rect 6260 5325 6295 5425
rect 6455 5325 6490 5425
rect 6510 5325 6545 5425
rect 6705 5325 6740 5425
rect 6760 5325 6795 5425
rect 6955 5325 6990 5425
rect 7010 5325 7045 5425
rect 7205 5325 7240 5425
rect 7260 5325 7295 5425
rect 7455 5325 7490 5425
rect 7510 5325 7545 5425
rect 7705 5325 7740 5425
rect 7760 5325 7795 5425
rect 7955 5325 7990 5425
rect 75 5260 175 5295
rect 75 5205 175 5240
rect 325 5260 425 5295
rect 325 5205 425 5240
rect 575 5260 675 5295
rect 575 5205 675 5240
rect 825 5260 925 5295
rect 825 5205 925 5240
rect 1075 5260 1175 5295
rect 1075 5205 1175 5240
rect 1325 5260 1425 5295
rect 1325 5205 1425 5240
rect 1575 5260 1675 5295
rect 1575 5205 1675 5240
rect 1825 5260 1925 5295
rect 1825 5205 1925 5240
rect 2075 5260 2175 5295
rect 2075 5205 2175 5240
rect 2325 5260 2425 5295
rect 2325 5205 2425 5240
rect 2575 5260 2675 5295
rect 2575 5205 2675 5240
rect 2825 5260 2925 5295
rect 2825 5205 2925 5240
rect 3075 5260 3175 5295
rect 3075 5205 3175 5240
rect 3325 5260 3425 5295
rect 3325 5205 3425 5240
rect 3575 5260 3675 5295
rect 3575 5205 3675 5240
rect 3825 5260 3925 5295
rect 3825 5205 3925 5240
rect 4075 5260 4175 5295
rect 4075 5205 4175 5240
rect 4325 5260 4425 5295
rect 4325 5205 4425 5240
rect 4575 5260 4675 5295
rect 4575 5205 4675 5240
rect 4825 5260 4925 5295
rect 4825 5205 4925 5240
rect 5075 5260 5175 5295
rect 5075 5205 5175 5240
rect 5325 5260 5425 5295
rect 5325 5205 5425 5240
rect 5575 5260 5675 5295
rect 5575 5205 5675 5240
rect 5825 5260 5925 5295
rect 5825 5205 5925 5240
rect 6075 5260 6175 5295
rect 6075 5205 6175 5240
rect 6325 5260 6425 5295
rect 6325 5205 6425 5240
rect 6575 5260 6675 5295
rect 6575 5205 6675 5240
rect 6825 5260 6925 5295
rect 6825 5205 6925 5240
rect 7075 5260 7175 5295
rect 7075 5205 7175 5240
rect 7325 5260 7425 5295
rect 7325 5205 7425 5240
rect 7575 5260 7675 5295
rect 7575 5205 7675 5240
rect 7825 5260 7925 5295
rect 7825 5205 7925 5240
rect 10 5075 45 5175
rect 205 5075 240 5175
rect 260 5075 295 5175
rect 455 5075 490 5175
rect 510 5075 545 5175
rect 705 5075 740 5175
rect 760 5075 795 5175
rect 955 5075 990 5175
rect 1010 5075 1045 5175
rect 1205 5075 1240 5175
rect 1260 5075 1295 5175
rect 1455 5075 1490 5175
rect 1510 5075 1545 5175
rect 1705 5075 1740 5175
rect 1760 5075 1795 5175
rect 1955 5075 1990 5175
rect 2010 5075 2045 5175
rect 2205 5075 2240 5175
rect 2260 5075 2295 5175
rect 2455 5075 2490 5175
rect 2510 5075 2545 5175
rect 2705 5075 2740 5175
rect 2760 5075 2795 5175
rect 2955 5075 2990 5175
rect 3010 5075 3045 5175
rect 3205 5075 3240 5175
rect 3260 5075 3295 5175
rect 3455 5075 3490 5175
rect 3510 5075 3545 5175
rect 3705 5075 3740 5175
rect 3760 5075 3795 5175
rect 3955 5075 3990 5175
rect 4010 5075 4045 5175
rect 4205 5075 4240 5175
rect 4260 5075 4295 5175
rect 4455 5075 4490 5175
rect 4510 5075 4545 5175
rect 4705 5075 4740 5175
rect 4760 5075 4795 5175
rect 4955 5075 4990 5175
rect 5010 5075 5045 5175
rect 5205 5075 5240 5175
rect 5260 5075 5295 5175
rect 5455 5075 5490 5175
rect 5510 5075 5545 5175
rect 5705 5075 5740 5175
rect 5760 5075 5795 5175
rect 5955 5075 5990 5175
rect 6010 5075 6045 5175
rect 6205 5075 6240 5175
rect 6260 5075 6295 5175
rect 6455 5075 6490 5175
rect 6510 5075 6545 5175
rect 6705 5075 6740 5175
rect 6760 5075 6795 5175
rect 6955 5075 6990 5175
rect 7010 5075 7045 5175
rect 7205 5075 7240 5175
rect 7260 5075 7295 5175
rect 7455 5075 7490 5175
rect 7510 5075 7545 5175
rect 7705 5075 7740 5175
rect 7760 5075 7795 5175
rect 7955 5075 7990 5175
rect 75 5010 175 5045
rect 75 4955 175 4990
rect 325 5010 425 5045
rect 325 4955 425 4990
rect 575 5010 675 5045
rect 575 4955 675 4990
rect 825 5010 925 5045
rect 825 4955 925 4990
rect 1075 5010 1175 5045
rect 1075 4955 1175 4990
rect 1325 5010 1425 5045
rect 1325 4955 1425 4990
rect 1575 5010 1675 5045
rect 1575 4955 1675 4990
rect 1825 5010 1925 5045
rect 1825 4955 1925 4990
rect 2075 5010 2175 5045
rect 2075 4955 2175 4990
rect 2325 5010 2425 5045
rect 2325 4955 2425 4990
rect 2575 5010 2675 5045
rect 2575 4955 2675 4990
rect 2825 5010 2925 5045
rect 2825 4955 2925 4990
rect 3075 5010 3175 5045
rect 3075 4955 3175 4990
rect 3325 5010 3425 5045
rect 3325 4955 3425 4990
rect 3575 5010 3675 5045
rect 3575 4955 3675 4990
rect 3825 5010 3925 5045
rect 3825 4955 3925 4990
rect 4075 5010 4175 5045
rect 4075 4955 4175 4990
rect 4325 5010 4425 5045
rect 4325 4955 4425 4990
rect 4575 5010 4675 5045
rect 4575 4955 4675 4990
rect 4825 5010 4925 5045
rect 4825 4955 4925 4990
rect 5075 5010 5175 5045
rect 5075 4955 5175 4990
rect 5325 5010 5425 5045
rect 5325 4955 5425 4990
rect 5575 5010 5675 5045
rect 5575 4955 5675 4990
rect 5825 5010 5925 5045
rect 5825 4955 5925 4990
rect 6075 5010 6175 5045
rect 6075 4955 6175 4990
rect 6325 5010 6425 5045
rect 6325 4955 6425 4990
rect 6575 5010 6675 5045
rect 6575 4955 6675 4990
rect 6825 5010 6925 5045
rect 6825 4955 6925 4990
rect 7075 5010 7175 5045
rect 7075 4955 7175 4990
rect 7325 5010 7425 5045
rect 7325 4955 7425 4990
rect 7575 5010 7675 5045
rect 7575 4955 7675 4990
rect 7825 5010 7925 5045
rect 7825 4955 7925 4990
rect 10 4825 45 4925
rect 205 4825 240 4925
rect 260 4825 295 4925
rect 455 4825 490 4925
rect 510 4825 545 4925
rect 705 4825 740 4925
rect 760 4825 795 4925
rect 955 4825 990 4925
rect 1010 4825 1045 4925
rect 1205 4825 1240 4925
rect 1260 4825 1295 4925
rect 1455 4825 1490 4925
rect 1510 4825 1545 4925
rect 1705 4825 1740 4925
rect 1760 4825 1795 4925
rect 1955 4825 1990 4925
rect 2010 4825 2045 4925
rect 2205 4825 2240 4925
rect 2260 4825 2295 4925
rect 2455 4825 2490 4925
rect 2510 4825 2545 4925
rect 2705 4825 2740 4925
rect 2760 4825 2795 4925
rect 2955 4825 2990 4925
rect 3010 4825 3045 4925
rect 3205 4825 3240 4925
rect 3260 4825 3295 4925
rect 3455 4825 3490 4925
rect 3510 4825 3545 4925
rect 3705 4825 3740 4925
rect 3760 4825 3795 4925
rect 3955 4825 3990 4925
rect 4010 4825 4045 4925
rect 4205 4825 4240 4925
rect 4260 4825 4295 4925
rect 4455 4825 4490 4925
rect 4510 4825 4545 4925
rect 4705 4825 4740 4925
rect 4760 4825 4795 4925
rect 4955 4825 4990 4925
rect 5010 4825 5045 4925
rect 5205 4825 5240 4925
rect 5260 4825 5295 4925
rect 5455 4825 5490 4925
rect 5510 4825 5545 4925
rect 5705 4825 5740 4925
rect 5760 4825 5795 4925
rect 5955 4825 5990 4925
rect 6010 4825 6045 4925
rect 6205 4825 6240 4925
rect 6260 4825 6295 4925
rect 6455 4825 6490 4925
rect 6510 4825 6545 4925
rect 6705 4825 6740 4925
rect 6760 4825 6795 4925
rect 6955 4825 6990 4925
rect 7010 4825 7045 4925
rect 7205 4825 7240 4925
rect 7260 4825 7295 4925
rect 7455 4825 7490 4925
rect 7510 4825 7545 4925
rect 7705 4825 7740 4925
rect 7760 4825 7795 4925
rect 7955 4825 7990 4925
rect 75 4760 175 4795
rect 75 4705 175 4740
rect 325 4760 425 4795
rect 325 4705 425 4740
rect 575 4760 675 4795
rect 575 4705 675 4740
rect 825 4760 925 4795
rect 825 4705 925 4740
rect 1075 4760 1175 4795
rect 1075 4705 1175 4740
rect 1325 4760 1425 4795
rect 1325 4705 1425 4740
rect 1575 4760 1675 4795
rect 1575 4705 1675 4740
rect 1825 4760 1925 4795
rect 1825 4705 1925 4740
rect 2075 4760 2175 4795
rect 2075 4705 2175 4740
rect 2325 4760 2425 4795
rect 2325 4705 2425 4740
rect 2575 4760 2675 4795
rect 2575 4705 2675 4740
rect 2825 4760 2925 4795
rect 2825 4705 2925 4740
rect 3075 4760 3175 4795
rect 3075 4705 3175 4740
rect 3325 4760 3425 4795
rect 3325 4705 3425 4740
rect 3575 4760 3675 4795
rect 3575 4705 3675 4740
rect 3825 4760 3925 4795
rect 3825 4705 3925 4740
rect 4075 4760 4175 4795
rect 4075 4705 4175 4740
rect 4325 4760 4425 4795
rect 4325 4705 4425 4740
rect 4575 4760 4675 4795
rect 4575 4705 4675 4740
rect 4825 4760 4925 4795
rect 4825 4705 4925 4740
rect 5075 4760 5175 4795
rect 5075 4705 5175 4740
rect 5325 4760 5425 4795
rect 5325 4705 5425 4740
rect 5575 4760 5675 4795
rect 5575 4705 5675 4740
rect 5825 4760 5925 4795
rect 5825 4705 5925 4740
rect 6075 4760 6175 4795
rect 6075 4705 6175 4740
rect 6325 4760 6425 4795
rect 6325 4705 6425 4740
rect 6575 4760 6675 4795
rect 6575 4705 6675 4740
rect 6825 4760 6925 4795
rect 6825 4705 6925 4740
rect 7075 4760 7175 4795
rect 7075 4705 7175 4740
rect 7325 4760 7425 4795
rect 7325 4705 7425 4740
rect 7575 4760 7675 4795
rect 7575 4705 7675 4740
rect 7825 4760 7925 4795
rect 7825 4705 7925 4740
rect 10 4575 45 4675
rect 205 4575 240 4675
rect 260 4575 295 4675
rect 455 4575 490 4675
rect 510 4575 545 4675
rect 705 4575 740 4675
rect 760 4575 795 4675
rect 955 4575 990 4675
rect 1010 4575 1045 4675
rect 1205 4575 1240 4675
rect 1260 4575 1295 4675
rect 1455 4575 1490 4675
rect 1510 4575 1545 4675
rect 1705 4575 1740 4675
rect 1760 4575 1795 4675
rect 1955 4575 1990 4675
rect 2010 4575 2045 4675
rect 2205 4575 2240 4675
rect 2260 4575 2295 4675
rect 2455 4575 2490 4675
rect 2510 4575 2545 4675
rect 2705 4575 2740 4675
rect 2760 4575 2795 4675
rect 2955 4575 2990 4675
rect 3010 4575 3045 4675
rect 3205 4575 3240 4675
rect 3260 4575 3295 4675
rect 3455 4575 3490 4675
rect 3510 4575 3545 4675
rect 3705 4575 3740 4675
rect 3760 4575 3795 4675
rect 3955 4575 3990 4675
rect 4010 4575 4045 4675
rect 4205 4575 4240 4675
rect 4260 4575 4295 4675
rect 4455 4575 4490 4675
rect 4510 4575 4545 4675
rect 4705 4575 4740 4675
rect 4760 4575 4795 4675
rect 4955 4575 4990 4675
rect 5010 4575 5045 4675
rect 5205 4575 5240 4675
rect 5260 4575 5295 4675
rect 5455 4575 5490 4675
rect 5510 4575 5545 4675
rect 5705 4575 5740 4675
rect 5760 4575 5795 4675
rect 5955 4575 5990 4675
rect 6010 4575 6045 4675
rect 6205 4575 6240 4675
rect 6260 4575 6295 4675
rect 6455 4575 6490 4675
rect 6510 4575 6545 4675
rect 6705 4575 6740 4675
rect 6760 4575 6795 4675
rect 6955 4575 6990 4675
rect 7010 4575 7045 4675
rect 7205 4575 7240 4675
rect 7260 4575 7295 4675
rect 7455 4575 7490 4675
rect 7510 4575 7545 4675
rect 7705 4575 7740 4675
rect 7760 4575 7795 4675
rect 7955 4575 7990 4675
rect 75 4510 175 4545
rect 75 4455 175 4490
rect 325 4510 425 4545
rect 325 4455 425 4490
rect 575 4510 675 4545
rect 575 4455 675 4490
rect 825 4510 925 4545
rect 825 4455 925 4490
rect 1075 4510 1175 4545
rect 1075 4455 1175 4490
rect 1325 4510 1425 4545
rect 1325 4455 1425 4490
rect 1575 4510 1675 4545
rect 1575 4455 1675 4490
rect 1825 4510 1925 4545
rect 1825 4455 1925 4490
rect 2075 4510 2175 4545
rect 2075 4455 2175 4490
rect 2325 4510 2425 4545
rect 2325 4455 2425 4490
rect 2575 4510 2675 4545
rect 2575 4455 2675 4490
rect 2825 4510 2925 4545
rect 2825 4455 2925 4490
rect 3075 4510 3175 4545
rect 3075 4455 3175 4490
rect 3325 4510 3425 4545
rect 3325 4455 3425 4490
rect 3575 4510 3675 4545
rect 3575 4455 3675 4490
rect 3825 4510 3925 4545
rect 3825 4455 3925 4490
rect 4075 4510 4175 4545
rect 4075 4455 4175 4490
rect 4325 4510 4425 4545
rect 4325 4455 4425 4490
rect 4575 4510 4675 4545
rect 4575 4455 4675 4490
rect 4825 4510 4925 4545
rect 4825 4455 4925 4490
rect 5075 4510 5175 4545
rect 5075 4455 5175 4490
rect 5325 4510 5425 4545
rect 5325 4455 5425 4490
rect 5575 4510 5675 4545
rect 5575 4455 5675 4490
rect 5825 4510 5925 4545
rect 5825 4455 5925 4490
rect 6075 4510 6175 4545
rect 6075 4455 6175 4490
rect 6325 4510 6425 4545
rect 6325 4455 6425 4490
rect 6575 4510 6675 4545
rect 6575 4455 6675 4490
rect 6825 4510 6925 4545
rect 6825 4455 6925 4490
rect 7075 4510 7175 4545
rect 7075 4455 7175 4490
rect 7325 4510 7425 4545
rect 7325 4455 7425 4490
rect 7575 4510 7675 4545
rect 7575 4455 7675 4490
rect 7825 4510 7925 4545
rect 7825 4455 7925 4490
rect 10 4325 45 4425
rect 205 4325 240 4425
rect 260 4325 295 4425
rect 455 4325 490 4425
rect 510 4325 545 4425
rect 705 4325 740 4425
rect 760 4325 795 4425
rect 955 4325 990 4425
rect 1010 4325 1045 4425
rect 1205 4325 1240 4425
rect 1260 4325 1295 4425
rect 1455 4325 1490 4425
rect 1510 4325 1545 4425
rect 1705 4325 1740 4425
rect 1760 4325 1795 4425
rect 1955 4325 1990 4425
rect 2010 4325 2045 4425
rect 2205 4325 2240 4425
rect 2260 4325 2295 4425
rect 2455 4325 2490 4425
rect 2510 4325 2545 4425
rect 2705 4325 2740 4425
rect 2760 4325 2795 4425
rect 2955 4325 2990 4425
rect 3010 4325 3045 4425
rect 3205 4325 3240 4425
rect 3260 4325 3295 4425
rect 3455 4325 3490 4425
rect 3510 4325 3545 4425
rect 3705 4325 3740 4425
rect 3760 4325 3795 4425
rect 3955 4325 3990 4425
rect 4010 4325 4045 4425
rect 4205 4325 4240 4425
rect 4260 4325 4295 4425
rect 4455 4325 4490 4425
rect 4510 4325 4545 4425
rect 4705 4325 4740 4425
rect 4760 4325 4795 4425
rect 4955 4325 4990 4425
rect 5010 4325 5045 4425
rect 5205 4325 5240 4425
rect 5260 4325 5295 4425
rect 5455 4325 5490 4425
rect 5510 4325 5545 4425
rect 5705 4325 5740 4425
rect 5760 4325 5795 4425
rect 5955 4325 5990 4425
rect 6010 4325 6045 4425
rect 6205 4325 6240 4425
rect 6260 4325 6295 4425
rect 6455 4325 6490 4425
rect 6510 4325 6545 4425
rect 6705 4325 6740 4425
rect 6760 4325 6795 4425
rect 6955 4325 6990 4425
rect 7010 4325 7045 4425
rect 7205 4325 7240 4425
rect 7260 4325 7295 4425
rect 7455 4325 7490 4425
rect 7510 4325 7545 4425
rect 7705 4325 7740 4425
rect 7760 4325 7795 4425
rect 7955 4325 7990 4425
rect 75 4260 175 4295
rect 75 4205 175 4240
rect 325 4260 425 4295
rect 325 4205 425 4240
rect 575 4260 675 4295
rect 575 4205 675 4240
rect 825 4260 925 4295
rect 825 4205 925 4240
rect 1075 4260 1175 4295
rect 1075 4205 1175 4240
rect 1325 4260 1425 4295
rect 1325 4205 1425 4240
rect 1575 4260 1675 4295
rect 1575 4205 1675 4240
rect 1825 4260 1925 4295
rect 1825 4205 1925 4240
rect 2075 4260 2175 4295
rect 2075 4205 2175 4240
rect 2325 4260 2425 4295
rect 2325 4205 2425 4240
rect 2575 4260 2675 4295
rect 2575 4205 2675 4240
rect 2825 4260 2925 4295
rect 2825 4205 2925 4240
rect 3075 4260 3175 4295
rect 3075 4205 3175 4240
rect 3325 4260 3425 4295
rect 3325 4205 3425 4240
rect 3575 4260 3675 4295
rect 3575 4205 3675 4240
rect 3825 4260 3925 4295
rect 3825 4205 3925 4240
rect 4075 4260 4175 4295
rect 4075 4205 4175 4240
rect 4325 4260 4425 4295
rect 4325 4205 4425 4240
rect 4575 4260 4675 4295
rect 4575 4205 4675 4240
rect 4825 4260 4925 4295
rect 4825 4205 4925 4240
rect 5075 4260 5175 4295
rect 5075 4205 5175 4240
rect 5325 4260 5425 4295
rect 5325 4205 5425 4240
rect 5575 4260 5675 4295
rect 5575 4205 5675 4240
rect 5825 4260 5925 4295
rect 5825 4205 5925 4240
rect 6075 4260 6175 4295
rect 6075 4205 6175 4240
rect 6325 4260 6425 4295
rect 6325 4205 6425 4240
rect 6575 4260 6675 4295
rect 6575 4205 6675 4240
rect 6825 4260 6925 4295
rect 6825 4205 6925 4240
rect 7075 4260 7175 4295
rect 7075 4205 7175 4240
rect 7325 4260 7425 4295
rect 7325 4205 7425 4240
rect 7575 4260 7675 4295
rect 7575 4205 7675 4240
rect 7825 4260 7925 4295
rect 7825 4205 7925 4240
rect 10 4075 45 4175
rect 205 4075 240 4175
rect 260 4075 295 4175
rect 455 4075 490 4175
rect 510 4075 545 4175
rect 705 4075 740 4175
rect 760 4075 795 4175
rect 955 4075 990 4175
rect 1010 4075 1045 4175
rect 1205 4075 1240 4175
rect 1260 4075 1295 4175
rect 1455 4075 1490 4175
rect 1510 4075 1545 4175
rect 1705 4075 1740 4175
rect 1760 4075 1795 4175
rect 1955 4075 1990 4175
rect 2010 4075 2045 4175
rect 2205 4075 2240 4175
rect 2260 4075 2295 4175
rect 2455 4075 2490 4175
rect 2510 4075 2545 4175
rect 2705 4075 2740 4175
rect 2760 4075 2795 4175
rect 2955 4075 2990 4175
rect 3010 4075 3045 4175
rect 3205 4075 3240 4175
rect 3260 4075 3295 4175
rect 3455 4075 3490 4175
rect 3510 4075 3545 4175
rect 3705 4075 3740 4175
rect 3760 4075 3795 4175
rect 3955 4075 3990 4175
rect 4010 4075 4045 4175
rect 4205 4075 4240 4175
rect 4260 4075 4295 4175
rect 4455 4075 4490 4175
rect 4510 4075 4545 4175
rect 4705 4075 4740 4175
rect 4760 4075 4795 4175
rect 4955 4075 4990 4175
rect 5010 4075 5045 4175
rect 5205 4075 5240 4175
rect 5260 4075 5295 4175
rect 5455 4075 5490 4175
rect 5510 4075 5545 4175
rect 5705 4075 5740 4175
rect 5760 4075 5795 4175
rect 5955 4075 5990 4175
rect 6010 4075 6045 4175
rect 6205 4075 6240 4175
rect 6260 4075 6295 4175
rect 6455 4075 6490 4175
rect 6510 4075 6545 4175
rect 6705 4075 6740 4175
rect 6760 4075 6795 4175
rect 6955 4075 6990 4175
rect 7010 4075 7045 4175
rect 7205 4075 7240 4175
rect 7260 4075 7295 4175
rect 7455 4075 7490 4175
rect 7510 4075 7545 4175
rect 7705 4075 7740 4175
rect 7760 4075 7795 4175
rect 7955 4075 7990 4175
rect 75 4010 175 4045
rect 75 3955 175 3990
rect 325 4010 425 4045
rect 325 3955 425 3990
rect 575 4010 675 4045
rect 575 3955 675 3990
rect 825 4010 925 4045
rect 825 3955 925 3990
rect 1075 4010 1175 4045
rect 1075 3955 1175 3990
rect 1325 4010 1425 4045
rect 1325 3955 1425 3990
rect 1575 4010 1675 4045
rect 1575 3955 1675 3990
rect 1825 4010 1925 4045
rect 1825 3955 1925 3990
rect 2075 4010 2175 4045
rect 2075 3955 2175 3990
rect 2325 4010 2425 4045
rect 2325 3955 2425 3990
rect 2575 4010 2675 4045
rect 2575 3955 2675 3990
rect 2825 4010 2925 4045
rect 2825 3955 2925 3990
rect 3075 4010 3175 4045
rect 3075 3955 3175 3990
rect 3325 4010 3425 4045
rect 3325 3955 3425 3990
rect 3575 4010 3675 4045
rect 3575 3955 3675 3990
rect 3825 4010 3925 4045
rect 3825 3955 3925 3990
rect 4075 4010 4175 4045
rect 4075 3955 4175 3990
rect 4325 4010 4425 4045
rect 4325 3955 4425 3990
rect 4575 4010 4675 4045
rect 4575 3955 4675 3990
rect 4825 4010 4925 4045
rect 4825 3955 4925 3990
rect 5075 4010 5175 4045
rect 5075 3955 5175 3990
rect 5325 4010 5425 4045
rect 5325 3955 5425 3990
rect 5575 4010 5675 4045
rect 5575 3955 5675 3990
rect 5825 4010 5925 4045
rect 5825 3955 5925 3990
rect 6075 4010 6175 4045
rect 6075 3955 6175 3990
rect 6325 4010 6425 4045
rect 6325 3955 6425 3990
rect 6575 4010 6675 4045
rect 6575 3955 6675 3990
rect 6825 4010 6925 4045
rect 6825 3955 6925 3990
rect 7075 4010 7175 4045
rect 7075 3955 7175 3990
rect 7325 4010 7425 4045
rect 7325 3955 7425 3990
rect 7575 4010 7675 4045
rect 7575 3955 7675 3990
rect 7825 4010 7925 4045
rect 7825 3955 7925 3990
rect 10 3825 45 3925
rect 205 3825 240 3925
rect 260 3825 295 3925
rect 455 3825 490 3925
rect 510 3825 545 3925
rect 705 3825 740 3925
rect 760 3825 795 3925
rect 955 3825 990 3925
rect 1010 3825 1045 3925
rect 1205 3825 1240 3925
rect 1260 3825 1295 3925
rect 1455 3825 1490 3925
rect 1510 3825 1545 3925
rect 1705 3825 1740 3925
rect 1760 3825 1795 3925
rect 1955 3825 1990 3925
rect 2010 3825 2045 3925
rect 2205 3825 2240 3925
rect 2260 3825 2295 3925
rect 2455 3825 2490 3925
rect 2510 3825 2545 3925
rect 2705 3825 2740 3925
rect 2760 3825 2795 3925
rect 2955 3825 2990 3925
rect 3010 3825 3045 3925
rect 3205 3825 3240 3925
rect 3260 3825 3295 3925
rect 3455 3825 3490 3925
rect 3510 3825 3545 3925
rect 3705 3825 3740 3925
rect 3760 3825 3795 3925
rect 3955 3825 3990 3925
rect 4010 3825 4045 3925
rect 4205 3825 4240 3925
rect 4260 3825 4295 3925
rect 4455 3825 4490 3925
rect 4510 3825 4545 3925
rect 4705 3825 4740 3925
rect 4760 3825 4795 3925
rect 4955 3825 4990 3925
rect 5010 3825 5045 3925
rect 5205 3825 5240 3925
rect 5260 3825 5295 3925
rect 5455 3825 5490 3925
rect 5510 3825 5545 3925
rect 5705 3825 5740 3925
rect 5760 3825 5795 3925
rect 5955 3825 5990 3925
rect 6010 3825 6045 3925
rect 6205 3825 6240 3925
rect 6260 3825 6295 3925
rect 6455 3825 6490 3925
rect 6510 3825 6545 3925
rect 6705 3825 6740 3925
rect 6760 3825 6795 3925
rect 6955 3825 6990 3925
rect 7010 3825 7045 3925
rect 7205 3825 7240 3925
rect 7260 3825 7295 3925
rect 7455 3825 7490 3925
rect 7510 3825 7545 3925
rect 7705 3825 7740 3925
rect 7760 3825 7795 3925
rect 7955 3825 7990 3925
rect 75 3760 175 3795
rect 75 3705 175 3740
rect 325 3760 425 3795
rect 325 3705 425 3740
rect 575 3760 675 3795
rect 575 3705 675 3740
rect 825 3760 925 3795
rect 825 3705 925 3740
rect 1075 3760 1175 3795
rect 1075 3705 1175 3740
rect 1325 3760 1425 3795
rect 1325 3705 1425 3740
rect 1575 3760 1675 3795
rect 1575 3705 1675 3740
rect 1825 3760 1925 3795
rect 1825 3705 1925 3740
rect 2075 3760 2175 3795
rect 2075 3705 2175 3740
rect 2325 3760 2425 3795
rect 2325 3705 2425 3740
rect 2575 3760 2675 3795
rect 2575 3705 2675 3740
rect 2825 3760 2925 3795
rect 2825 3705 2925 3740
rect 3075 3760 3175 3795
rect 3075 3705 3175 3740
rect 3325 3760 3425 3795
rect 3325 3705 3425 3740
rect 3575 3760 3675 3795
rect 3575 3705 3675 3740
rect 3825 3760 3925 3795
rect 3825 3705 3925 3740
rect 4075 3760 4175 3795
rect 4075 3705 4175 3740
rect 4325 3760 4425 3795
rect 4325 3705 4425 3740
rect 4575 3760 4675 3795
rect 4575 3705 4675 3740
rect 4825 3760 4925 3795
rect 4825 3705 4925 3740
rect 5075 3760 5175 3795
rect 5075 3705 5175 3740
rect 5325 3760 5425 3795
rect 5325 3705 5425 3740
rect 5575 3760 5675 3795
rect 5575 3705 5675 3740
rect 5825 3760 5925 3795
rect 5825 3705 5925 3740
rect 6075 3760 6175 3795
rect 6075 3705 6175 3740
rect 6325 3760 6425 3795
rect 6325 3705 6425 3740
rect 6575 3760 6675 3795
rect 6575 3705 6675 3740
rect 6825 3760 6925 3795
rect 6825 3705 6925 3740
rect 7075 3760 7175 3795
rect 7075 3705 7175 3740
rect 7325 3760 7425 3795
rect 7325 3705 7425 3740
rect 7575 3760 7675 3795
rect 7575 3705 7675 3740
rect 7825 3760 7925 3795
rect 7825 3705 7925 3740
rect 10 3575 45 3675
rect 205 3575 240 3675
rect 260 3575 295 3675
rect 455 3575 490 3675
rect 510 3575 545 3675
rect 705 3575 740 3675
rect 760 3575 795 3675
rect 955 3575 990 3675
rect 1010 3575 1045 3675
rect 1205 3575 1240 3675
rect 1260 3575 1295 3675
rect 1455 3575 1490 3675
rect 1510 3575 1545 3675
rect 1705 3575 1740 3675
rect 1760 3575 1795 3675
rect 1955 3575 1990 3675
rect 2010 3575 2045 3675
rect 2205 3575 2240 3675
rect 2260 3575 2295 3675
rect 2455 3575 2490 3675
rect 2510 3575 2545 3675
rect 2705 3575 2740 3675
rect 2760 3575 2795 3675
rect 2955 3575 2990 3675
rect 3010 3575 3045 3675
rect 3205 3575 3240 3675
rect 3260 3575 3295 3675
rect 3455 3575 3490 3675
rect 3510 3575 3545 3675
rect 3705 3575 3740 3675
rect 3760 3575 3795 3675
rect 3955 3575 3990 3675
rect 4010 3575 4045 3675
rect 4205 3575 4240 3675
rect 4260 3575 4295 3675
rect 4455 3575 4490 3675
rect 4510 3575 4545 3675
rect 4705 3575 4740 3675
rect 4760 3575 4795 3675
rect 4955 3575 4990 3675
rect 5010 3575 5045 3675
rect 5205 3575 5240 3675
rect 5260 3575 5295 3675
rect 5455 3575 5490 3675
rect 5510 3575 5545 3675
rect 5705 3575 5740 3675
rect 5760 3575 5795 3675
rect 5955 3575 5990 3675
rect 6010 3575 6045 3675
rect 6205 3575 6240 3675
rect 6260 3575 6295 3675
rect 6455 3575 6490 3675
rect 6510 3575 6545 3675
rect 6705 3575 6740 3675
rect 6760 3575 6795 3675
rect 6955 3575 6990 3675
rect 7010 3575 7045 3675
rect 7205 3575 7240 3675
rect 7260 3575 7295 3675
rect 7455 3575 7490 3675
rect 7510 3575 7545 3675
rect 7705 3575 7740 3675
rect 7760 3575 7795 3675
rect 7955 3575 7990 3675
rect 75 3510 175 3545
rect 75 3455 175 3490
rect 325 3510 425 3545
rect 325 3455 425 3490
rect 575 3510 675 3545
rect 575 3455 675 3490
rect 825 3510 925 3545
rect 825 3455 925 3490
rect 1075 3510 1175 3545
rect 1075 3455 1175 3490
rect 1325 3510 1425 3545
rect 1325 3455 1425 3490
rect 1575 3510 1675 3545
rect 1575 3455 1675 3490
rect 1825 3510 1925 3545
rect 1825 3455 1925 3490
rect 2075 3510 2175 3545
rect 2075 3455 2175 3490
rect 2325 3510 2425 3545
rect 2325 3455 2425 3490
rect 2575 3510 2675 3545
rect 2575 3455 2675 3490
rect 2825 3510 2925 3545
rect 2825 3455 2925 3490
rect 3075 3510 3175 3545
rect 3075 3455 3175 3490
rect 3325 3510 3425 3545
rect 3325 3455 3425 3490
rect 3575 3510 3675 3545
rect 3575 3455 3675 3490
rect 3825 3510 3925 3545
rect 3825 3455 3925 3490
rect 4075 3510 4175 3545
rect 4075 3455 4175 3490
rect 4325 3510 4425 3545
rect 4325 3455 4425 3490
rect 4575 3510 4675 3545
rect 4575 3455 4675 3490
rect 4825 3510 4925 3545
rect 4825 3455 4925 3490
rect 5075 3510 5175 3545
rect 5075 3455 5175 3490
rect 5325 3510 5425 3545
rect 5325 3455 5425 3490
rect 5575 3510 5675 3545
rect 5575 3455 5675 3490
rect 5825 3510 5925 3545
rect 5825 3455 5925 3490
rect 6075 3510 6175 3545
rect 6075 3455 6175 3490
rect 6325 3510 6425 3545
rect 6325 3455 6425 3490
rect 6575 3510 6675 3545
rect 6575 3455 6675 3490
rect 6825 3510 6925 3545
rect 6825 3455 6925 3490
rect 7075 3510 7175 3545
rect 7075 3455 7175 3490
rect 7325 3510 7425 3545
rect 7325 3455 7425 3490
rect 7575 3510 7675 3545
rect 7575 3455 7675 3490
rect 7825 3510 7925 3545
rect 7825 3455 7925 3490
rect 10 3325 45 3425
rect 205 3325 240 3425
rect 260 3325 295 3425
rect 455 3325 490 3425
rect 510 3325 545 3425
rect 705 3325 740 3425
rect 760 3325 795 3425
rect 955 3325 990 3425
rect 1010 3325 1045 3425
rect 1205 3325 1240 3425
rect 1260 3325 1295 3425
rect 1455 3325 1490 3425
rect 1510 3325 1545 3425
rect 1705 3325 1740 3425
rect 1760 3325 1795 3425
rect 1955 3325 1990 3425
rect 2010 3325 2045 3425
rect 2205 3325 2240 3425
rect 2260 3325 2295 3425
rect 2455 3325 2490 3425
rect 2510 3325 2545 3425
rect 2705 3325 2740 3425
rect 2760 3325 2795 3425
rect 2955 3325 2990 3425
rect 3010 3325 3045 3425
rect 3205 3325 3240 3425
rect 3260 3325 3295 3425
rect 3455 3325 3490 3425
rect 3510 3325 3545 3425
rect 3705 3325 3740 3425
rect 3760 3325 3795 3425
rect 3955 3325 3990 3425
rect 4010 3325 4045 3425
rect 4205 3325 4240 3425
rect 4260 3325 4295 3425
rect 4455 3325 4490 3425
rect 4510 3325 4545 3425
rect 4705 3325 4740 3425
rect 4760 3325 4795 3425
rect 4955 3325 4990 3425
rect 5010 3325 5045 3425
rect 5205 3325 5240 3425
rect 5260 3325 5295 3425
rect 5455 3325 5490 3425
rect 5510 3325 5545 3425
rect 5705 3325 5740 3425
rect 5760 3325 5795 3425
rect 5955 3325 5990 3425
rect 6010 3325 6045 3425
rect 6205 3325 6240 3425
rect 6260 3325 6295 3425
rect 6455 3325 6490 3425
rect 6510 3325 6545 3425
rect 6705 3325 6740 3425
rect 6760 3325 6795 3425
rect 6955 3325 6990 3425
rect 7010 3325 7045 3425
rect 7205 3325 7240 3425
rect 7260 3325 7295 3425
rect 7455 3325 7490 3425
rect 7510 3325 7545 3425
rect 7705 3325 7740 3425
rect 7760 3325 7795 3425
rect 7955 3325 7990 3425
rect 75 3260 175 3295
rect 75 3205 175 3240
rect 325 3260 425 3295
rect 325 3205 425 3240
rect 575 3260 675 3295
rect 575 3205 675 3240
rect 825 3260 925 3295
rect 825 3205 925 3240
rect 1075 3260 1175 3295
rect 1075 3205 1175 3240
rect 1325 3260 1425 3295
rect 1325 3205 1425 3240
rect 1575 3260 1675 3295
rect 1575 3205 1675 3240
rect 1825 3260 1925 3295
rect 1825 3205 1925 3240
rect 2075 3260 2175 3295
rect 2075 3205 2175 3240
rect 2325 3260 2425 3295
rect 2325 3205 2425 3240
rect 2575 3260 2675 3295
rect 2575 3205 2675 3240
rect 2825 3260 2925 3295
rect 2825 3205 2925 3240
rect 3075 3260 3175 3295
rect 3075 3205 3175 3240
rect 3325 3260 3425 3295
rect 3325 3205 3425 3240
rect 3575 3260 3675 3295
rect 3575 3205 3675 3240
rect 3825 3260 3925 3295
rect 3825 3205 3925 3240
rect 4075 3260 4175 3295
rect 4075 3205 4175 3240
rect 4325 3260 4425 3295
rect 4325 3205 4425 3240
rect 4575 3260 4675 3295
rect 4575 3205 4675 3240
rect 4825 3260 4925 3295
rect 4825 3205 4925 3240
rect 5075 3260 5175 3295
rect 5075 3205 5175 3240
rect 5325 3260 5425 3295
rect 5325 3205 5425 3240
rect 5575 3260 5675 3295
rect 5575 3205 5675 3240
rect 5825 3260 5925 3295
rect 5825 3205 5925 3240
rect 6075 3260 6175 3295
rect 6075 3205 6175 3240
rect 6325 3260 6425 3295
rect 6325 3205 6425 3240
rect 6575 3260 6675 3295
rect 6575 3205 6675 3240
rect 6825 3260 6925 3295
rect 6825 3205 6925 3240
rect 7075 3260 7175 3295
rect 7075 3205 7175 3240
rect 7325 3260 7425 3295
rect 7325 3205 7425 3240
rect 7575 3260 7675 3295
rect 7575 3205 7675 3240
rect 7825 3260 7925 3295
rect 7825 3205 7925 3240
rect 10 3075 45 3175
rect 205 3075 240 3175
rect 260 3075 295 3175
rect 455 3075 490 3175
rect 510 3075 545 3175
rect 705 3075 740 3175
rect 760 3075 795 3175
rect 955 3075 990 3175
rect 1010 3075 1045 3175
rect 1205 3075 1240 3175
rect 1260 3075 1295 3175
rect 1455 3075 1490 3175
rect 1510 3075 1545 3175
rect 1705 3075 1740 3175
rect 1760 3075 1795 3175
rect 1955 3075 1990 3175
rect 2010 3075 2045 3175
rect 2205 3075 2240 3175
rect 2260 3075 2295 3175
rect 2455 3075 2490 3175
rect 2510 3075 2545 3175
rect 2705 3075 2740 3175
rect 2760 3075 2795 3175
rect 2955 3075 2990 3175
rect 3010 3075 3045 3175
rect 3205 3075 3240 3175
rect 3260 3075 3295 3175
rect 3455 3075 3490 3175
rect 3510 3075 3545 3175
rect 3705 3075 3740 3175
rect 3760 3075 3795 3175
rect 3955 3075 3990 3175
rect 4010 3075 4045 3175
rect 4205 3075 4240 3175
rect 4260 3075 4295 3175
rect 4455 3075 4490 3175
rect 4510 3075 4545 3175
rect 4705 3075 4740 3175
rect 4760 3075 4795 3175
rect 4955 3075 4990 3175
rect 5010 3075 5045 3175
rect 5205 3075 5240 3175
rect 5260 3075 5295 3175
rect 5455 3075 5490 3175
rect 5510 3075 5545 3175
rect 5705 3075 5740 3175
rect 5760 3075 5795 3175
rect 5955 3075 5990 3175
rect 6010 3075 6045 3175
rect 6205 3075 6240 3175
rect 6260 3075 6295 3175
rect 6455 3075 6490 3175
rect 6510 3075 6545 3175
rect 6705 3075 6740 3175
rect 6760 3075 6795 3175
rect 6955 3075 6990 3175
rect 7010 3075 7045 3175
rect 7205 3075 7240 3175
rect 7260 3075 7295 3175
rect 7455 3075 7490 3175
rect 7510 3075 7545 3175
rect 7705 3075 7740 3175
rect 7760 3075 7795 3175
rect 7955 3075 7990 3175
rect 75 3010 175 3045
rect 75 2955 175 2990
rect 325 3010 425 3045
rect 325 2955 425 2990
rect 575 3010 675 3045
rect 575 2955 675 2990
rect 825 3010 925 3045
rect 825 2955 925 2990
rect 1075 3010 1175 3045
rect 1075 2955 1175 2990
rect 1325 3010 1425 3045
rect 1325 2955 1425 2990
rect 1575 3010 1675 3045
rect 1575 2955 1675 2990
rect 1825 3010 1925 3045
rect 1825 2955 1925 2990
rect 2075 3010 2175 3045
rect 2075 2955 2175 2990
rect 2325 3010 2425 3045
rect 2325 2955 2425 2990
rect 2575 3010 2675 3045
rect 2575 2955 2675 2990
rect 2825 3010 2925 3045
rect 2825 2955 2925 2990
rect 3075 3010 3175 3045
rect 3075 2955 3175 2990
rect 3325 3010 3425 3045
rect 3325 2955 3425 2990
rect 3575 3010 3675 3045
rect 3575 2955 3675 2990
rect 3825 3010 3925 3045
rect 3825 2955 3925 2990
rect 4075 3010 4175 3045
rect 4075 2955 4175 2990
rect 4325 3010 4425 3045
rect 4325 2955 4425 2990
rect 4575 3010 4675 3045
rect 4575 2955 4675 2990
rect 4825 3010 4925 3045
rect 4825 2955 4925 2990
rect 5075 3010 5175 3045
rect 5075 2955 5175 2990
rect 5325 3010 5425 3045
rect 5325 2955 5425 2990
rect 5575 3010 5675 3045
rect 5575 2955 5675 2990
rect 5825 3010 5925 3045
rect 5825 2955 5925 2990
rect 6075 3010 6175 3045
rect 6075 2955 6175 2990
rect 6325 3010 6425 3045
rect 6325 2955 6425 2990
rect 6575 3010 6675 3045
rect 6575 2955 6675 2990
rect 6825 3010 6925 3045
rect 6825 2955 6925 2990
rect 7075 3010 7175 3045
rect 7075 2955 7175 2990
rect 7325 3010 7425 3045
rect 7325 2955 7425 2990
rect 7575 3010 7675 3045
rect 7575 2955 7675 2990
rect 7825 3010 7925 3045
rect 7825 2955 7925 2990
rect 10 2825 45 2925
rect 205 2825 240 2925
rect 260 2825 295 2925
rect 455 2825 490 2925
rect 510 2825 545 2925
rect 705 2825 740 2925
rect 760 2825 795 2925
rect 955 2825 990 2925
rect 1010 2825 1045 2925
rect 1205 2825 1240 2925
rect 1260 2825 1295 2925
rect 1455 2825 1490 2925
rect 1510 2825 1545 2925
rect 1705 2825 1740 2925
rect 1760 2825 1795 2925
rect 1955 2825 1990 2925
rect 2010 2825 2045 2925
rect 2205 2825 2240 2925
rect 2260 2825 2295 2925
rect 2455 2825 2490 2925
rect 2510 2825 2545 2925
rect 2705 2825 2740 2925
rect 2760 2825 2795 2925
rect 2955 2825 2990 2925
rect 3010 2825 3045 2925
rect 3205 2825 3240 2925
rect 3260 2825 3295 2925
rect 3455 2825 3490 2925
rect 3510 2825 3545 2925
rect 3705 2825 3740 2925
rect 3760 2825 3795 2925
rect 3955 2825 3990 2925
rect 4010 2825 4045 2925
rect 4205 2825 4240 2925
rect 4260 2825 4295 2925
rect 4455 2825 4490 2925
rect 4510 2825 4545 2925
rect 4705 2825 4740 2925
rect 4760 2825 4795 2925
rect 4955 2825 4990 2925
rect 5010 2825 5045 2925
rect 5205 2825 5240 2925
rect 5260 2825 5295 2925
rect 5455 2825 5490 2925
rect 5510 2825 5545 2925
rect 5705 2825 5740 2925
rect 5760 2825 5795 2925
rect 5955 2825 5990 2925
rect 6010 2825 6045 2925
rect 6205 2825 6240 2925
rect 6260 2825 6295 2925
rect 6455 2825 6490 2925
rect 6510 2825 6545 2925
rect 6705 2825 6740 2925
rect 6760 2825 6795 2925
rect 6955 2825 6990 2925
rect 7010 2825 7045 2925
rect 7205 2825 7240 2925
rect 7260 2825 7295 2925
rect 7455 2825 7490 2925
rect 7510 2825 7545 2925
rect 7705 2825 7740 2925
rect 7760 2825 7795 2925
rect 7955 2825 7990 2925
rect 75 2760 175 2795
rect 75 2705 175 2740
rect 325 2760 425 2795
rect 325 2705 425 2740
rect 575 2760 675 2795
rect 575 2705 675 2740
rect 825 2760 925 2795
rect 825 2705 925 2740
rect 1075 2760 1175 2795
rect 1075 2705 1175 2740
rect 1325 2760 1425 2795
rect 1325 2705 1425 2740
rect 1575 2760 1675 2795
rect 1575 2705 1675 2740
rect 1825 2760 1925 2795
rect 1825 2705 1925 2740
rect 2075 2760 2175 2795
rect 2075 2705 2175 2740
rect 2325 2760 2425 2795
rect 2325 2705 2425 2740
rect 2575 2760 2675 2795
rect 2575 2705 2675 2740
rect 2825 2760 2925 2795
rect 2825 2705 2925 2740
rect 3075 2760 3175 2795
rect 3075 2705 3175 2740
rect 3325 2760 3425 2795
rect 3325 2705 3425 2740
rect 3575 2760 3675 2795
rect 3575 2705 3675 2740
rect 3825 2760 3925 2795
rect 3825 2705 3925 2740
rect 4075 2760 4175 2795
rect 4075 2705 4175 2740
rect 4325 2760 4425 2795
rect 4325 2705 4425 2740
rect 4575 2760 4675 2795
rect 4575 2705 4675 2740
rect 4825 2760 4925 2795
rect 4825 2705 4925 2740
rect 5075 2760 5175 2795
rect 5075 2705 5175 2740
rect 5325 2760 5425 2795
rect 5325 2705 5425 2740
rect 5575 2760 5675 2795
rect 5575 2705 5675 2740
rect 5825 2760 5925 2795
rect 5825 2705 5925 2740
rect 6075 2760 6175 2795
rect 6075 2705 6175 2740
rect 6325 2760 6425 2795
rect 6325 2705 6425 2740
rect 6575 2760 6675 2795
rect 6575 2705 6675 2740
rect 6825 2760 6925 2795
rect 6825 2705 6925 2740
rect 7075 2760 7175 2795
rect 7075 2705 7175 2740
rect 7325 2760 7425 2795
rect 7325 2705 7425 2740
rect 7575 2760 7675 2795
rect 7575 2705 7675 2740
rect 7825 2760 7925 2795
rect 7825 2705 7925 2740
rect 10 2575 45 2675
rect 205 2575 240 2675
rect 260 2575 295 2675
rect 455 2575 490 2675
rect 510 2575 545 2675
rect 705 2575 740 2675
rect 760 2575 795 2675
rect 955 2575 990 2675
rect 1010 2575 1045 2675
rect 1205 2575 1240 2675
rect 1260 2575 1295 2675
rect 1455 2575 1490 2675
rect 1510 2575 1545 2675
rect 1705 2575 1740 2675
rect 1760 2575 1795 2675
rect 1955 2575 1990 2675
rect 2010 2575 2045 2675
rect 2205 2575 2240 2675
rect 2260 2575 2295 2675
rect 2455 2575 2490 2675
rect 2510 2575 2545 2675
rect 2705 2575 2740 2675
rect 2760 2575 2795 2675
rect 2955 2575 2990 2675
rect 3010 2575 3045 2675
rect 3205 2575 3240 2675
rect 3260 2575 3295 2675
rect 3455 2575 3490 2675
rect 3510 2575 3545 2675
rect 3705 2575 3740 2675
rect 3760 2575 3795 2675
rect 3955 2575 3990 2675
rect 4010 2575 4045 2675
rect 4205 2575 4240 2675
rect 4260 2575 4295 2675
rect 4455 2575 4490 2675
rect 4510 2575 4545 2675
rect 4705 2575 4740 2675
rect 4760 2575 4795 2675
rect 4955 2575 4990 2675
rect 5010 2575 5045 2675
rect 5205 2575 5240 2675
rect 5260 2575 5295 2675
rect 5455 2575 5490 2675
rect 5510 2575 5545 2675
rect 5705 2575 5740 2675
rect 5760 2575 5795 2675
rect 5955 2575 5990 2675
rect 6010 2575 6045 2675
rect 6205 2575 6240 2675
rect 6260 2575 6295 2675
rect 6455 2575 6490 2675
rect 6510 2575 6545 2675
rect 6705 2575 6740 2675
rect 6760 2575 6795 2675
rect 6955 2575 6990 2675
rect 7010 2575 7045 2675
rect 7205 2575 7240 2675
rect 7260 2575 7295 2675
rect 7455 2575 7490 2675
rect 7510 2575 7545 2675
rect 7705 2575 7740 2675
rect 7760 2575 7795 2675
rect 7955 2575 7990 2675
rect 75 2510 175 2545
rect 75 2455 175 2490
rect 325 2510 425 2545
rect 325 2455 425 2490
rect 575 2510 675 2545
rect 575 2455 675 2490
rect 825 2510 925 2545
rect 825 2455 925 2490
rect 1075 2510 1175 2545
rect 1075 2455 1175 2490
rect 1325 2510 1425 2545
rect 1325 2455 1425 2490
rect 1575 2510 1675 2545
rect 1575 2455 1675 2490
rect 1825 2510 1925 2545
rect 1825 2455 1925 2490
rect 2075 2510 2175 2545
rect 2075 2455 2175 2490
rect 2325 2510 2425 2545
rect 2325 2455 2425 2490
rect 2575 2510 2675 2545
rect 2575 2455 2675 2490
rect 2825 2510 2925 2545
rect 2825 2455 2925 2490
rect 3075 2510 3175 2545
rect 3075 2455 3175 2490
rect 3325 2510 3425 2545
rect 3325 2455 3425 2490
rect 3575 2510 3675 2545
rect 3575 2455 3675 2490
rect 3825 2510 3925 2545
rect 3825 2455 3925 2490
rect 4075 2510 4175 2545
rect 4075 2455 4175 2490
rect 4325 2510 4425 2545
rect 4325 2455 4425 2490
rect 4575 2510 4675 2545
rect 4575 2455 4675 2490
rect 4825 2510 4925 2545
rect 4825 2455 4925 2490
rect 5075 2510 5175 2545
rect 5075 2455 5175 2490
rect 5325 2510 5425 2545
rect 5325 2455 5425 2490
rect 5575 2510 5675 2545
rect 5575 2455 5675 2490
rect 5825 2510 5925 2545
rect 5825 2455 5925 2490
rect 6075 2510 6175 2545
rect 6075 2455 6175 2490
rect 6325 2510 6425 2545
rect 6325 2455 6425 2490
rect 6575 2510 6675 2545
rect 6575 2455 6675 2490
rect 6825 2510 6925 2545
rect 6825 2455 6925 2490
rect 7075 2510 7175 2545
rect 7075 2455 7175 2490
rect 7325 2510 7425 2545
rect 7325 2455 7425 2490
rect 7575 2510 7675 2545
rect 7575 2455 7675 2490
rect 7825 2510 7925 2545
rect 7825 2455 7925 2490
rect 10 2325 45 2425
rect 205 2325 240 2425
rect 260 2325 295 2425
rect 455 2325 490 2425
rect 510 2325 545 2425
rect 705 2325 740 2425
rect 760 2325 795 2425
rect 955 2325 990 2425
rect 1010 2325 1045 2425
rect 1205 2325 1240 2425
rect 1260 2325 1295 2425
rect 1455 2325 1490 2425
rect 1510 2325 1545 2425
rect 1705 2325 1740 2425
rect 1760 2325 1795 2425
rect 1955 2325 1990 2425
rect 2010 2325 2045 2425
rect 2205 2325 2240 2425
rect 2260 2325 2295 2425
rect 2455 2325 2490 2425
rect 2510 2325 2545 2425
rect 2705 2325 2740 2425
rect 2760 2325 2795 2425
rect 2955 2325 2990 2425
rect 3010 2325 3045 2425
rect 3205 2325 3240 2425
rect 3260 2325 3295 2425
rect 3455 2325 3490 2425
rect 3510 2325 3545 2425
rect 3705 2325 3740 2425
rect 3760 2325 3795 2425
rect 3955 2325 3990 2425
rect 4010 2325 4045 2425
rect 4205 2325 4240 2425
rect 4260 2325 4295 2425
rect 4455 2325 4490 2425
rect 4510 2325 4545 2425
rect 4705 2325 4740 2425
rect 4760 2325 4795 2425
rect 4955 2325 4990 2425
rect 5010 2325 5045 2425
rect 5205 2325 5240 2425
rect 5260 2325 5295 2425
rect 5455 2325 5490 2425
rect 5510 2325 5545 2425
rect 5705 2325 5740 2425
rect 5760 2325 5795 2425
rect 5955 2325 5990 2425
rect 6010 2325 6045 2425
rect 6205 2325 6240 2425
rect 6260 2325 6295 2425
rect 6455 2325 6490 2425
rect 6510 2325 6545 2425
rect 6705 2325 6740 2425
rect 6760 2325 6795 2425
rect 6955 2325 6990 2425
rect 7010 2325 7045 2425
rect 7205 2325 7240 2425
rect 7260 2325 7295 2425
rect 7455 2325 7490 2425
rect 7510 2325 7545 2425
rect 7705 2325 7740 2425
rect 7760 2325 7795 2425
rect 7955 2325 7990 2425
rect 75 2260 175 2295
rect 75 2205 175 2240
rect 325 2260 425 2295
rect 325 2205 425 2240
rect 575 2260 675 2295
rect 575 2205 675 2240
rect 825 2260 925 2295
rect 825 2205 925 2240
rect 1075 2260 1175 2295
rect 1075 2205 1175 2240
rect 1325 2260 1425 2295
rect 1325 2205 1425 2240
rect 1575 2260 1675 2295
rect 1575 2205 1675 2240
rect 1825 2260 1925 2295
rect 1825 2205 1925 2240
rect 2075 2260 2175 2295
rect 2075 2205 2175 2240
rect 2325 2260 2425 2295
rect 2325 2205 2425 2240
rect 2575 2260 2675 2295
rect 2575 2205 2675 2240
rect 2825 2260 2925 2295
rect 2825 2205 2925 2240
rect 3075 2260 3175 2295
rect 3075 2205 3175 2240
rect 3325 2260 3425 2295
rect 3325 2205 3425 2240
rect 3575 2260 3675 2295
rect 3575 2205 3675 2240
rect 3825 2260 3925 2295
rect 3825 2205 3925 2240
rect 4075 2260 4175 2295
rect 4075 2205 4175 2240
rect 4325 2260 4425 2295
rect 4325 2205 4425 2240
rect 4575 2260 4675 2295
rect 4575 2205 4675 2240
rect 4825 2260 4925 2295
rect 4825 2205 4925 2240
rect 5075 2260 5175 2295
rect 5075 2205 5175 2240
rect 5325 2260 5425 2295
rect 5325 2205 5425 2240
rect 5575 2260 5675 2295
rect 5575 2205 5675 2240
rect 5825 2260 5925 2295
rect 5825 2205 5925 2240
rect 6075 2260 6175 2295
rect 6075 2205 6175 2240
rect 6325 2260 6425 2295
rect 6325 2205 6425 2240
rect 6575 2260 6675 2295
rect 6575 2205 6675 2240
rect 6825 2260 6925 2295
rect 6825 2205 6925 2240
rect 7075 2260 7175 2295
rect 7075 2205 7175 2240
rect 7325 2260 7425 2295
rect 7325 2205 7425 2240
rect 7575 2260 7675 2295
rect 7575 2205 7675 2240
rect 7825 2260 7925 2295
rect 7825 2205 7925 2240
rect 10 2075 45 2175
rect 205 2075 240 2175
rect 260 2075 295 2175
rect 455 2075 490 2175
rect 510 2075 545 2175
rect 705 2075 740 2175
rect 760 2075 795 2175
rect 955 2075 990 2175
rect 1010 2075 1045 2175
rect 1205 2075 1240 2175
rect 1260 2075 1295 2175
rect 1455 2075 1490 2175
rect 1510 2075 1545 2175
rect 1705 2075 1740 2175
rect 1760 2075 1795 2175
rect 1955 2075 1990 2175
rect 2010 2075 2045 2175
rect 2205 2075 2240 2175
rect 2260 2075 2295 2175
rect 2455 2075 2490 2175
rect 2510 2075 2545 2175
rect 2705 2075 2740 2175
rect 2760 2075 2795 2175
rect 2955 2075 2990 2175
rect 3010 2075 3045 2175
rect 3205 2075 3240 2175
rect 3260 2075 3295 2175
rect 3455 2075 3490 2175
rect 3510 2075 3545 2175
rect 3705 2075 3740 2175
rect 3760 2075 3795 2175
rect 3955 2075 3990 2175
rect 4010 2075 4045 2175
rect 4205 2075 4240 2175
rect 4260 2075 4295 2175
rect 4455 2075 4490 2175
rect 4510 2075 4545 2175
rect 4705 2075 4740 2175
rect 4760 2075 4795 2175
rect 4955 2075 4990 2175
rect 5010 2075 5045 2175
rect 5205 2075 5240 2175
rect 5260 2075 5295 2175
rect 5455 2075 5490 2175
rect 5510 2075 5545 2175
rect 5705 2075 5740 2175
rect 5760 2075 5795 2175
rect 5955 2075 5990 2175
rect 6010 2075 6045 2175
rect 6205 2075 6240 2175
rect 6260 2075 6295 2175
rect 6455 2075 6490 2175
rect 6510 2075 6545 2175
rect 6705 2075 6740 2175
rect 6760 2075 6795 2175
rect 6955 2075 6990 2175
rect 7010 2075 7045 2175
rect 7205 2075 7240 2175
rect 7260 2075 7295 2175
rect 7455 2075 7490 2175
rect 7510 2075 7545 2175
rect 7705 2075 7740 2175
rect 7760 2075 7795 2175
rect 7955 2075 7990 2175
rect 75 2010 175 2045
rect 75 1955 175 1990
rect 325 2010 425 2045
rect 325 1955 425 1990
rect 575 2010 675 2045
rect 575 1955 675 1990
rect 825 2010 925 2045
rect 825 1955 925 1990
rect 1075 2010 1175 2045
rect 1075 1955 1175 1990
rect 1325 2010 1425 2045
rect 1325 1955 1425 1990
rect 1575 2010 1675 2045
rect 1575 1955 1675 1990
rect 1825 2010 1925 2045
rect 1825 1955 1925 1990
rect 2075 2010 2175 2045
rect 2075 1955 2175 1990
rect 2325 2010 2425 2045
rect 2325 1955 2425 1990
rect 2575 2010 2675 2045
rect 2575 1955 2675 1990
rect 2825 2010 2925 2045
rect 2825 1955 2925 1990
rect 3075 2010 3175 2045
rect 3075 1955 3175 1990
rect 3325 2010 3425 2045
rect 3325 1955 3425 1990
rect 3575 2010 3675 2045
rect 3575 1955 3675 1990
rect 3825 2010 3925 2045
rect 3825 1955 3925 1990
rect 4075 2010 4175 2045
rect 4075 1955 4175 1990
rect 4325 2010 4425 2045
rect 4325 1955 4425 1990
rect 4575 2010 4675 2045
rect 4575 1955 4675 1990
rect 4825 2010 4925 2045
rect 4825 1955 4925 1990
rect 5075 2010 5175 2045
rect 5075 1955 5175 1990
rect 5325 2010 5425 2045
rect 5325 1955 5425 1990
rect 5575 2010 5675 2045
rect 5575 1955 5675 1990
rect 5825 2010 5925 2045
rect 5825 1955 5925 1990
rect 6075 2010 6175 2045
rect 6075 1955 6175 1990
rect 6325 2010 6425 2045
rect 6325 1955 6425 1990
rect 6575 2010 6675 2045
rect 6575 1955 6675 1990
rect 6825 2010 6925 2045
rect 6825 1955 6925 1990
rect 7075 2010 7175 2045
rect 7075 1955 7175 1990
rect 7325 2010 7425 2045
rect 7325 1955 7425 1990
rect 7575 2010 7675 2045
rect 7575 1955 7675 1990
rect 7825 2010 7925 2045
rect 7825 1955 7925 1990
rect 10 1825 45 1925
rect 205 1825 240 1925
rect 260 1825 295 1925
rect 455 1825 490 1925
rect 510 1825 545 1925
rect 705 1825 740 1925
rect 760 1825 795 1925
rect 955 1825 990 1925
rect 1010 1825 1045 1925
rect 1205 1825 1240 1925
rect 1260 1825 1295 1925
rect 1455 1825 1490 1925
rect 1510 1825 1545 1925
rect 1705 1825 1740 1925
rect 1760 1825 1795 1925
rect 1955 1825 1990 1925
rect 2010 1825 2045 1925
rect 2205 1825 2240 1925
rect 2260 1825 2295 1925
rect 2455 1825 2490 1925
rect 2510 1825 2545 1925
rect 2705 1825 2740 1925
rect 2760 1825 2795 1925
rect 2955 1825 2990 1925
rect 3010 1825 3045 1925
rect 3205 1825 3240 1925
rect 3260 1825 3295 1925
rect 3455 1825 3490 1925
rect 3510 1825 3545 1925
rect 3705 1825 3740 1925
rect 3760 1825 3795 1925
rect 3955 1825 3990 1925
rect 4010 1825 4045 1925
rect 4205 1825 4240 1925
rect 4260 1825 4295 1925
rect 4455 1825 4490 1925
rect 4510 1825 4545 1925
rect 4705 1825 4740 1925
rect 4760 1825 4795 1925
rect 4955 1825 4990 1925
rect 5010 1825 5045 1925
rect 5205 1825 5240 1925
rect 5260 1825 5295 1925
rect 5455 1825 5490 1925
rect 5510 1825 5545 1925
rect 5705 1825 5740 1925
rect 5760 1825 5795 1925
rect 5955 1825 5990 1925
rect 6010 1825 6045 1925
rect 6205 1825 6240 1925
rect 6260 1825 6295 1925
rect 6455 1825 6490 1925
rect 6510 1825 6545 1925
rect 6705 1825 6740 1925
rect 6760 1825 6795 1925
rect 6955 1825 6990 1925
rect 7010 1825 7045 1925
rect 7205 1825 7240 1925
rect 7260 1825 7295 1925
rect 7455 1825 7490 1925
rect 7510 1825 7545 1925
rect 7705 1825 7740 1925
rect 7760 1825 7795 1925
rect 7955 1825 7990 1925
rect 75 1760 175 1795
rect 75 1705 175 1740
rect 325 1760 425 1795
rect 325 1705 425 1740
rect 575 1760 675 1795
rect 575 1705 675 1740
rect 825 1760 925 1795
rect 825 1705 925 1740
rect 1075 1760 1175 1795
rect 1075 1705 1175 1740
rect 1325 1760 1425 1795
rect 1325 1705 1425 1740
rect 1575 1760 1675 1795
rect 1575 1705 1675 1740
rect 1825 1760 1925 1795
rect 1825 1705 1925 1740
rect 2075 1760 2175 1795
rect 2075 1705 2175 1740
rect 2325 1760 2425 1795
rect 2325 1705 2425 1740
rect 2575 1760 2675 1795
rect 2575 1705 2675 1740
rect 2825 1760 2925 1795
rect 2825 1705 2925 1740
rect 3075 1760 3175 1795
rect 3075 1705 3175 1740
rect 3325 1760 3425 1795
rect 3325 1705 3425 1740
rect 3575 1760 3675 1795
rect 3575 1705 3675 1740
rect 3825 1760 3925 1795
rect 3825 1705 3925 1740
rect 4075 1760 4175 1795
rect 4075 1705 4175 1740
rect 4325 1760 4425 1795
rect 4325 1705 4425 1740
rect 4575 1760 4675 1795
rect 4575 1705 4675 1740
rect 4825 1760 4925 1795
rect 4825 1705 4925 1740
rect 5075 1760 5175 1795
rect 5075 1705 5175 1740
rect 5325 1760 5425 1795
rect 5325 1705 5425 1740
rect 5575 1760 5675 1795
rect 5575 1705 5675 1740
rect 5825 1760 5925 1795
rect 5825 1705 5925 1740
rect 6075 1760 6175 1795
rect 6075 1705 6175 1740
rect 6325 1760 6425 1795
rect 6325 1705 6425 1740
rect 6575 1760 6675 1795
rect 6575 1705 6675 1740
rect 6825 1760 6925 1795
rect 6825 1705 6925 1740
rect 7075 1760 7175 1795
rect 7075 1705 7175 1740
rect 7325 1760 7425 1795
rect 7325 1705 7425 1740
rect 7575 1760 7675 1795
rect 7575 1705 7675 1740
rect 7825 1760 7925 1795
rect 7825 1705 7925 1740
rect 10 1575 45 1675
rect 205 1575 240 1675
rect 260 1575 295 1675
rect 455 1575 490 1675
rect 510 1575 545 1675
rect 705 1575 740 1675
rect 760 1575 795 1675
rect 955 1575 990 1675
rect 1010 1575 1045 1675
rect 1205 1575 1240 1675
rect 1260 1575 1295 1675
rect 1455 1575 1490 1675
rect 1510 1575 1545 1675
rect 1705 1575 1740 1675
rect 1760 1575 1795 1675
rect 1955 1575 1990 1675
rect 2010 1575 2045 1675
rect 2205 1575 2240 1675
rect 2260 1575 2295 1675
rect 2455 1575 2490 1675
rect 2510 1575 2545 1675
rect 2705 1575 2740 1675
rect 2760 1575 2795 1675
rect 2955 1575 2990 1675
rect 3010 1575 3045 1675
rect 3205 1575 3240 1675
rect 3260 1575 3295 1675
rect 3455 1575 3490 1675
rect 3510 1575 3545 1675
rect 3705 1575 3740 1675
rect 3760 1575 3795 1675
rect 3955 1575 3990 1675
rect 4010 1575 4045 1675
rect 4205 1575 4240 1675
rect 4260 1575 4295 1675
rect 4455 1575 4490 1675
rect 4510 1575 4545 1675
rect 4705 1575 4740 1675
rect 4760 1575 4795 1675
rect 4955 1575 4990 1675
rect 5010 1575 5045 1675
rect 5205 1575 5240 1675
rect 5260 1575 5295 1675
rect 5455 1575 5490 1675
rect 5510 1575 5545 1675
rect 5705 1575 5740 1675
rect 5760 1575 5795 1675
rect 5955 1575 5990 1675
rect 6010 1575 6045 1675
rect 6205 1575 6240 1675
rect 6260 1575 6295 1675
rect 6455 1575 6490 1675
rect 6510 1575 6545 1675
rect 6705 1575 6740 1675
rect 6760 1575 6795 1675
rect 6955 1575 6990 1675
rect 7010 1575 7045 1675
rect 7205 1575 7240 1675
rect 7260 1575 7295 1675
rect 7455 1575 7490 1675
rect 7510 1575 7545 1675
rect 7705 1575 7740 1675
rect 7760 1575 7795 1675
rect 7955 1575 7990 1675
rect 75 1510 175 1545
rect 75 1455 175 1490
rect 325 1510 425 1545
rect 325 1455 425 1490
rect 575 1510 675 1545
rect 575 1455 675 1490
rect 825 1510 925 1545
rect 825 1455 925 1490
rect 1075 1510 1175 1545
rect 1075 1455 1175 1490
rect 1325 1510 1425 1545
rect 1325 1455 1425 1490
rect 1575 1510 1675 1545
rect 1575 1455 1675 1490
rect 1825 1510 1925 1545
rect 1825 1455 1925 1490
rect 2075 1510 2175 1545
rect 2075 1455 2175 1490
rect 2325 1510 2425 1545
rect 2325 1455 2425 1490
rect 2575 1510 2675 1545
rect 2575 1455 2675 1490
rect 2825 1510 2925 1545
rect 2825 1455 2925 1490
rect 3075 1510 3175 1545
rect 3075 1455 3175 1490
rect 3325 1510 3425 1545
rect 3325 1455 3425 1490
rect 3575 1510 3675 1545
rect 3575 1455 3675 1490
rect 3825 1510 3925 1545
rect 3825 1455 3925 1490
rect 4075 1510 4175 1545
rect 4075 1455 4175 1490
rect 4325 1510 4425 1545
rect 4325 1455 4425 1490
rect 4575 1510 4675 1545
rect 4575 1455 4675 1490
rect 4825 1510 4925 1545
rect 4825 1455 4925 1490
rect 5075 1510 5175 1545
rect 5075 1455 5175 1490
rect 5325 1510 5425 1545
rect 5325 1455 5425 1490
rect 5575 1510 5675 1545
rect 5575 1455 5675 1490
rect 5825 1510 5925 1545
rect 5825 1455 5925 1490
rect 6075 1510 6175 1545
rect 6075 1455 6175 1490
rect 6325 1510 6425 1545
rect 6325 1455 6425 1490
rect 6575 1510 6675 1545
rect 6575 1455 6675 1490
rect 6825 1510 6925 1545
rect 6825 1455 6925 1490
rect 7075 1510 7175 1545
rect 7075 1455 7175 1490
rect 7325 1510 7425 1545
rect 7325 1455 7425 1490
rect 7575 1510 7675 1545
rect 7575 1455 7675 1490
rect 7825 1510 7925 1545
rect 7825 1455 7925 1490
rect 10 1325 45 1425
rect 205 1325 240 1425
rect 260 1325 295 1425
rect 455 1325 490 1425
rect 510 1325 545 1425
rect 705 1325 740 1425
rect 760 1325 795 1425
rect 955 1325 990 1425
rect 1010 1325 1045 1425
rect 1205 1325 1240 1425
rect 1260 1325 1295 1425
rect 1455 1325 1490 1425
rect 1510 1325 1545 1425
rect 1705 1325 1740 1425
rect 1760 1325 1795 1425
rect 1955 1325 1990 1425
rect 2010 1325 2045 1425
rect 2205 1325 2240 1425
rect 2260 1325 2295 1425
rect 2455 1325 2490 1425
rect 2510 1325 2545 1425
rect 2705 1325 2740 1425
rect 2760 1325 2795 1425
rect 2955 1325 2990 1425
rect 3010 1325 3045 1425
rect 3205 1325 3240 1425
rect 3260 1325 3295 1425
rect 3455 1325 3490 1425
rect 3510 1325 3545 1425
rect 3705 1325 3740 1425
rect 3760 1325 3795 1425
rect 3955 1325 3990 1425
rect 4010 1325 4045 1425
rect 4205 1325 4240 1425
rect 4260 1325 4295 1425
rect 4455 1325 4490 1425
rect 4510 1325 4545 1425
rect 4705 1325 4740 1425
rect 4760 1325 4795 1425
rect 4955 1325 4990 1425
rect 5010 1325 5045 1425
rect 5205 1325 5240 1425
rect 5260 1325 5295 1425
rect 5455 1325 5490 1425
rect 5510 1325 5545 1425
rect 5705 1325 5740 1425
rect 5760 1325 5795 1425
rect 5955 1325 5990 1425
rect 6010 1325 6045 1425
rect 6205 1325 6240 1425
rect 6260 1325 6295 1425
rect 6455 1325 6490 1425
rect 6510 1325 6545 1425
rect 6705 1325 6740 1425
rect 6760 1325 6795 1425
rect 6955 1325 6990 1425
rect 7010 1325 7045 1425
rect 7205 1325 7240 1425
rect 7260 1325 7295 1425
rect 7455 1325 7490 1425
rect 7510 1325 7545 1425
rect 7705 1325 7740 1425
rect 7760 1325 7795 1425
rect 7955 1325 7990 1425
rect 75 1260 175 1295
rect 75 1205 175 1240
rect 325 1260 425 1295
rect 325 1205 425 1240
rect 575 1260 675 1295
rect 575 1205 675 1240
rect 825 1260 925 1295
rect 825 1205 925 1240
rect 1075 1260 1175 1295
rect 1075 1205 1175 1240
rect 1325 1260 1425 1295
rect 1325 1205 1425 1240
rect 1575 1260 1675 1295
rect 1575 1205 1675 1240
rect 1825 1260 1925 1295
rect 1825 1205 1925 1240
rect 2075 1260 2175 1295
rect 2075 1205 2175 1240
rect 2325 1260 2425 1295
rect 2325 1205 2425 1240
rect 2575 1260 2675 1295
rect 2575 1205 2675 1240
rect 2825 1260 2925 1295
rect 2825 1205 2925 1240
rect 3075 1260 3175 1295
rect 3075 1205 3175 1240
rect 3325 1260 3425 1295
rect 3325 1205 3425 1240
rect 3575 1260 3675 1295
rect 3575 1205 3675 1240
rect 3825 1260 3925 1295
rect 3825 1205 3925 1240
rect 4075 1260 4175 1295
rect 4075 1205 4175 1240
rect 4325 1260 4425 1295
rect 4325 1205 4425 1240
rect 4575 1260 4675 1295
rect 4575 1205 4675 1240
rect 4825 1260 4925 1295
rect 4825 1205 4925 1240
rect 5075 1260 5175 1295
rect 5075 1205 5175 1240
rect 5325 1260 5425 1295
rect 5325 1205 5425 1240
rect 5575 1260 5675 1295
rect 5575 1205 5675 1240
rect 5825 1260 5925 1295
rect 5825 1205 5925 1240
rect 6075 1260 6175 1295
rect 6075 1205 6175 1240
rect 6325 1260 6425 1295
rect 6325 1205 6425 1240
rect 6575 1260 6675 1295
rect 6575 1205 6675 1240
rect 6825 1260 6925 1295
rect 6825 1205 6925 1240
rect 7075 1260 7175 1295
rect 7075 1205 7175 1240
rect 7325 1260 7425 1295
rect 7325 1205 7425 1240
rect 7575 1260 7675 1295
rect 7575 1205 7675 1240
rect 7825 1260 7925 1295
rect 7825 1205 7925 1240
rect 10 1075 45 1175
rect 205 1075 240 1175
rect 260 1075 295 1175
rect 455 1075 490 1175
rect 510 1075 545 1175
rect 705 1075 740 1175
rect 760 1075 795 1175
rect 955 1075 990 1175
rect 1010 1075 1045 1175
rect 1205 1075 1240 1175
rect 1260 1075 1295 1175
rect 1455 1075 1490 1175
rect 1510 1075 1545 1175
rect 1705 1075 1740 1175
rect 1760 1075 1795 1175
rect 1955 1075 1990 1175
rect 2010 1075 2045 1175
rect 2205 1075 2240 1175
rect 2260 1075 2295 1175
rect 2455 1075 2490 1175
rect 2510 1075 2545 1175
rect 2705 1075 2740 1175
rect 2760 1075 2795 1175
rect 2955 1075 2990 1175
rect 3010 1075 3045 1175
rect 3205 1075 3240 1175
rect 3260 1075 3295 1175
rect 3455 1075 3490 1175
rect 3510 1075 3545 1175
rect 3705 1075 3740 1175
rect 3760 1075 3795 1175
rect 3955 1075 3990 1175
rect 4010 1075 4045 1175
rect 4205 1075 4240 1175
rect 4260 1075 4295 1175
rect 4455 1075 4490 1175
rect 4510 1075 4545 1175
rect 4705 1075 4740 1175
rect 4760 1075 4795 1175
rect 4955 1075 4990 1175
rect 5010 1075 5045 1175
rect 5205 1075 5240 1175
rect 5260 1075 5295 1175
rect 5455 1075 5490 1175
rect 5510 1075 5545 1175
rect 5705 1075 5740 1175
rect 5760 1075 5795 1175
rect 5955 1075 5990 1175
rect 6010 1075 6045 1175
rect 6205 1075 6240 1175
rect 6260 1075 6295 1175
rect 6455 1075 6490 1175
rect 6510 1075 6545 1175
rect 6705 1075 6740 1175
rect 6760 1075 6795 1175
rect 6955 1075 6990 1175
rect 7010 1075 7045 1175
rect 7205 1075 7240 1175
rect 7260 1075 7295 1175
rect 7455 1075 7490 1175
rect 7510 1075 7545 1175
rect 7705 1075 7740 1175
rect 7760 1075 7795 1175
rect 7955 1075 7990 1175
rect 75 1010 175 1045
rect 75 955 175 990
rect 325 1010 425 1045
rect 325 955 425 990
rect 575 1010 675 1045
rect 575 955 675 990
rect 825 1010 925 1045
rect 825 955 925 990
rect 1075 1010 1175 1045
rect 1075 955 1175 990
rect 1325 1010 1425 1045
rect 1325 955 1425 990
rect 1575 1010 1675 1045
rect 1575 955 1675 990
rect 1825 1010 1925 1045
rect 1825 955 1925 990
rect 2075 1010 2175 1045
rect 2075 955 2175 990
rect 2325 1010 2425 1045
rect 2325 955 2425 990
rect 2575 1010 2675 1045
rect 2575 955 2675 990
rect 2825 1010 2925 1045
rect 2825 955 2925 990
rect 3075 1010 3175 1045
rect 3075 955 3175 990
rect 3325 1010 3425 1045
rect 3325 955 3425 990
rect 3575 1010 3675 1045
rect 3575 955 3675 990
rect 3825 1010 3925 1045
rect 3825 955 3925 990
rect 4075 1010 4175 1045
rect 4075 955 4175 990
rect 4325 1010 4425 1045
rect 4325 955 4425 990
rect 4575 1010 4675 1045
rect 4575 955 4675 990
rect 4825 1010 4925 1045
rect 4825 955 4925 990
rect 5075 1010 5175 1045
rect 5075 955 5175 990
rect 5325 1010 5425 1045
rect 5325 955 5425 990
rect 5575 1010 5675 1045
rect 5575 955 5675 990
rect 5825 1010 5925 1045
rect 5825 955 5925 990
rect 6075 1010 6175 1045
rect 6075 955 6175 990
rect 6325 1010 6425 1045
rect 6325 955 6425 990
rect 6575 1010 6675 1045
rect 6575 955 6675 990
rect 6825 1010 6925 1045
rect 6825 955 6925 990
rect 7075 1010 7175 1045
rect 7075 955 7175 990
rect 7325 1010 7425 1045
rect 7325 955 7425 990
rect 7575 1010 7675 1045
rect 7575 955 7675 990
rect 7825 1010 7925 1045
rect 7825 955 7925 990
rect 10 825 45 925
rect 205 825 240 925
rect 260 825 295 925
rect 455 825 490 925
rect 510 825 545 925
rect 705 825 740 925
rect 760 825 795 925
rect 955 825 990 925
rect 1010 825 1045 925
rect 1205 825 1240 925
rect 1260 825 1295 925
rect 1455 825 1490 925
rect 1510 825 1545 925
rect 1705 825 1740 925
rect 1760 825 1795 925
rect 1955 825 1990 925
rect 2010 825 2045 925
rect 2205 825 2240 925
rect 2260 825 2295 925
rect 2455 825 2490 925
rect 2510 825 2545 925
rect 2705 825 2740 925
rect 2760 825 2795 925
rect 2955 825 2990 925
rect 3010 825 3045 925
rect 3205 825 3240 925
rect 3260 825 3295 925
rect 3455 825 3490 925
rect 3510 825 3545 925
rect 3705 825 3740 925
rect 3760 825 3795 925
rect 3955 825 3990 925
rect 4010 825 4045 925
rect 4205 825 4240 925
rect 4260 825 4295 925
rect 4455 825 4490 925
rect 4510 825 4545 925
rect 4705 825 4740 925
rect 4760 825 4795 925
rect 4955 825 4990 925
rect 5010 825 5045 925
rect 5205 825 5240 925
rect 5260 825 5295 925
rect 5455 825 5490 925
rect 5510 825 5545 925
rect 5705 825 5740 925
rect 5760 825 5795 925
rect 5955 825 5990 925
rect 6010 825 6045 925
rect 6205 825 6240 925
rect 6260 825 6295 925
rect 6455 825 6490 925
rect 6510 825 6545 925
rect 6705 825 6740 925
rect 6760 825 6795 925
rect 6955 825 6990 925
rect 7010 825 7045 925
rect 7205 825 7240 925
rect 7260 825 7295 925
rect 7455 825 7490 925
rect 7510 825 7545 925
rect 7705 825 7740 925
rect 7760 825 7795 925
rect 7955 825 7990 925
rect 75 760 175 795
rect 75 705 175 740
rect 325 760 425 795
rect 325 705 425 740
rect 575 760 675 795
rect 575 705 675 740
rect 825 760 925 795
rect 825 705 925 740
rect 1075 760 1175 795
rect 1075 705 1175 740
rect 1325 760 1425 795
rect 1325 705 1425 740
rect 1575 760 1675 795
rect 1575 705 1675 740
rect 1825 760 1925 795
rect 1825 705 1925 740
rect 2075 760 2175 795
rect 2075 705 2175 740
rect 2325 760 2425 795
rect 2325 705 2425 740
rect 2575 760 2675 795
rect 2575 705 2675 740
rect 2825 760 2925 795
rect 2825 705 2925 740
rect 3075 760 3175 795
rect 3075 705 3175 740
rect 3325 760 3425 795
rect 3325 705 3425 740
rect 3575 760 3675 795
rect 3575 705 3675 740
rect 3825 760 3925 795
rect 3825 705 3925 740
rect 4075 760 4175 795
rect 4075 705 4175 740
rect 4325 760 4425 795
rect 4325 705 4425 740
rect 4575 760 4675 795
rect 4575 705 4675 740
rect 4825 760 4925 795
rect 4825 705 4925 740
rect 5075 760 5175 795
rect 5075 705 5175 740
rect 5325 760 5425 795
rect 5325 705 5425 740
rect 5575 760 5675 795
rect 5575 705 5675 740
rect 5825 760 5925 795
rect 5825 705 5925 740
rect 6075 760 6175 795
rect 6075 705 6175 740
rect 6325 760 6425 795
rect 6325 705 6425 740
rect 6575 760 6675 795
rect 6575 705 6675 740
rect 6825 760 6925 795
rect 6825 705 6925 740
rect 7075 760 7175 795
rect 7075 705 7175 740
rect 7325 760 7425 795
rect 7325 705 7425 740
rect 7575 760 7675 795
rect 7575 705 7675 740
rect 7825 760 7925 795
rect 7825 705 7925 740
rect 10 575 45 675
rect 205 575 240 675
rect 260 575 295 675
rect 455 575 490 675
rect 510 575 545 675
rect 705 575 740 675
rect 760 575 795 675
rect 955 575 990 675
rect 1010 575 1045 675
rect 1205 575 1240 675
rect 1260 575 1295 675
rect 1455 575 1490 675
rect 1510 575 1545 675
rect 1705 575 1740 675
rect 1760 575 1795 675
rect 1955 575 1990 675
rect 2010 575 2045 675
rect 2205 575 2240 675
rect 2260 575 2295 675
rect 2455 575 2490 675
rect 2510 575 2545 675
rect 2705 575 2740 675
rect 2760 575 2795 675
rect 2955 575 2990 675
rect 3010 575 3045 675
rect 3205 575 3240 675
rect 3260 575 3295 675
rect 3455 575 3490 675
rect 3510 575 3545 675
rect 3705 575 3740 675
rect 3760 575 3795 675
rect 3955 575 3990 675
rect 4010 575 4045 675
rect 4205 575 4240 675
rect 4260 575 4295 675
rect 4455 575 4490 675
rect 4510 575 4545 675
rect 4705 575 4740 675
rect 4760 575 4795 675
rect 4955 575 4990 675
rect 5010 575 5045 675
rect 5205 575 5240 675
rect 5260 575 5295 675
rect 5455 575 5490 675
rect 5510 575 5545 675
rect 5705 575 5740 675
rect 5760 575 5795 675
rect 5955 575 5990 675
rect 6010 575 6045 675
rect 6205 575 6240 675
rect 6260 575 6295 675
rect 6455 575 6490 675
rect 6510 575 6545 675
rect 6705 575 6740 675
rect 6760 575 6795 675
rect 6955 575 6990 675
rect 7010 575 7045 675
rect 7205 575 7240 675
rect 7260 575 7295 675
rect 7455 575 7490 675
rect 7510 575 7545 675
rect 7705 575 7740 675
rect 7760 575 7795 675
rect 7955 575 7990 675
rect 75 510 175 545
rect 75 455 175 490
rect 325 510 425 545
rect 325 455 425 490
rect 575 510 675 545
rect 575 455 675 490
rect 825 510 925 545
rect 825 455 925 490
rect 1075 510 1175 545
rect 1075 455 1175 490
rect 1325 510 1425 545
rect 1325 455 1425 490
rect 1575 510 1675 545
rect 1575 455 1675 490
rect 1825 510 1925 545
rect 1825 455 1925 490
rect 2075 510 2175 545
rect 2075 455 2175 490
rect 2325 510 2425 545
rect 2325 455 2425 490
rect 2575 510 2675 545
rect 2575 455 2675 490
rect 2825 510 2925 545
rect 2825 455 2925 490
rect 3075 510 3175 545
rect 3075 455 3175 490
rect 3325 510 3425 545
rect 3325 455 3425 490
rect 3575 510 3675 545
rect 3575 455 3675 490
rect 3825 510 3925 545
rect 3825 455 3925 490
rect 4075 510 4175 545
rect 4075 455 4175 490
rect 4325 510 4425 545
rect 4325 455 4425 490
rect 4575 510 4675 545
rect 4575 455 4675 490
rect 4825 510 4925 545
rect 4825 455 4925 490
rect 5075 510 5175 545
rect 5075 455 5175 490
rect 5325 510 5425 545
rect 5325 455 5425 490
rect 5575 510 5675 545
rect 5575 455 5675 490
rect 5825 510 5925 545
rect 5825 455 5925 490
rect 6075 510 6175 545
rect 6075 455 6175 490
rect 6325 510 6425 545
rect 6325 455 6425 490
rect 6575 510 6675 545
rect 6575 455 6675 490
rect 6825 510 6925 545
rect 6825 455 6925 490
rect 7075 510 7175 545
rect 7075 455 7175 490
rect 7325 510 7425 545
rect 7325 455 7425 490
rect 7575 510 7675 545
rect 7575 455 7675 490
rect 7825 510 7925 545
rect 7825 455 7925 490
rect 10 325 45 425
rect 205 325 240 425
rect 260 325 295 425
rect 455 325 490 425
rect 510 325 545 425
rect 705 325 740 425
rect 760 325 795 425
rect 955 325 990 425
rect 1010 325 1045 425
rect 1205 325 1240 425
rect 1260 325 1295 425
rect 1455 325 1490 425
rect 1510 325 1545 425
rect 1705 325 1740 425
rect 1760 325 1795 425
rect 1955 325 1990 425
rect 2010 325 2045 425
rect 2205 325 2240 425
rect 2260 325 2295 425
rect 2455 325 2490 425
rect 2510 325 2545 425
rect 2705 325 2740 425
rect 2760 325 2795 425
rect 2955 325 2990 425
rect 3010 325 3045 425
rect 3205 325 3240 425
rect 3260 325 3295 425
rect 3455 325 3490 425
rect 3510 325 3545 425
rect 3705 325 3740 425
rect 3760 325 3795 425
rect 3955 325 3990 425
rect 4010 325 4045 425
rect 4205 325 4240 425
rect 4260 325 4295 425
rect 4455 325 4490 425
rect 4510 325 4545 425
rect 4705 325 4740 425
rect 4760 325 4795 425
rect 4955 325 4990 425
rect 5010 325 5045 425
rect 5205 325 5240 425
rect 5260 325 5295 425
rect 5455 325 5490 425
rect 5510 325 5545 425
rect 5705 325 5740 425
rect 5760 325 5795 425
rect 5955 325 5990 425
rect 6010 325 6045 425
rect 6205 325 6240 425
rect 6260 325 6295 425
rect 6455 325 6490 425
rect 6510 325 6545 425
rect 6705 325 6740 425
rect 6760 325 6795 425
rect 6955 325 6990 425
rect 7010 325 7045 425
rect 7205 325 7240 425
rect 7260 325 7295 425
rect 7455 325 7490 425
rect 7510 325 7545 425
rect 7705 325 7740 425
rect 7760 325 7795 425
rect 7955 325 7990 425
rect 75 260 175 295
rect 75 205 175 240
rect 325 260 425 295
rect 325 205 425 240
rect 575 260 675 295
rect 575 205 675 240
rect 825 260 925 295
rect 825 205 925 240
rect 1075 260 1175 295
rect 1075 205 1175 240
rect 1325 260 1425 295
rect 1325 205 1425 240
rect 1575 260 1675 295
rect 1575 205 1675 240
rect 1825 260 1925 295
rect 1825 205 1925 240
rect 2075 260 2175 295
rect 2075 205 2175 240
rect 2325 260 2425 295
rect 2325 205 2425 240
rect 2575 260 2675 295
rect 2575 205 2675 240
rect 2825 260 2925 295
rect 2825 205 2925 240
rect 3075 260 3175 295
rect 3075 205 3175 240
rect 3325 260 3425 295
rect 3325 205 3425 240
rect 3575 260 3675 295
rect 3575 205 3675 240
rect 3825 260 3925 295
rect 3825 205 3925 240
rect 4075 260 4175 295
rect 4075 205 4175 240
rect 4325 260 4425 295
rect 4325 205 4425 240
rect 4575 260 4675 295
rect 4575 205 4675 240
rect 4825 260 4925 295
rect 4825 205 4925 240
rect 5075 260 5175 295
rect 5075 205 5175 240
rect 5325 260 5425 295
rect 5325 205 5425 240
rect 5575 260 5675 295
rect 5575 205 5675 240
rect 5825 260 5925 295
rect 5825 205 5925 240
rect 6075 260 6175 295
rect 6075 205 6175 240
rect 6325 260 6425 295
rect 6325 205 6425 240
rect 6575 260 6675 295
rect 6575 205 6675 240
rect 6825 260 6925 295
rect 6825 205 6925 240
rect 7075 260 7175 295
rect 7075 205 7175 240
rect 7325 260 7425 295
rect 7325 205 7425 240
rect 7575 260 7675 295
rect 7575 205 7675 240
rect 7825 260 7925 295
rect 7825 205 7925 240
rect 10 75 45 175
rect 205 75 240 175
rect 260 75 295 175
rect 455 75 490 175
rect 510 75 545 175
rect 705 75 740 175
rect 760 75 795 175
rect 955 75 990 175
rect 1010 75 1045 175
rect 1205 75 1240 175
rect 1260 75 1295 175
rect 1455 75 1490 175
rect 1510 75 1545 175
rect 1705 75 1740 175
rect 1760 75 1795 175
rect 1955 75 1990 175
rect 2010 75 2045 175
rect 2205 75 2240 175
rect 2260 75 2295 175
rect 2455 75 2490 175
rect 2510 75 2545 175
rect 2705 75 2740 175
rect 2760 75 2795 175
rect 2955 75 2990 175
rect 3010 75 3045 175
rect 3205 75 3240 175
rect 3260 75 3295 175
rect 3455 75 3490 175
rect 3510 75 3545 175
rect 3705 75 3740 175
rect 3760 75 3795 175
rect 3955 75 3990 175
rect 4010 75 4045 175
rect 4205 75 4240 175
rect 4260 75 4295 175
rect 4455 75 4490 175
rect 4510 75 4545 175
rect 4705 75 4740 175
rect 4760 75 4795 175
rect 4955 75 4990 175
rect 5010 75 5045 175
rect 5205 75 5240 175
rect 5260 75 5295 175
rect 5455 75 5490 175
rect 5510 75 5545 175
rect 5705 75 5740 175
rect 5760 75 5795 175
rect 5955 75 5990 175
rect 6010 75 6045 175
rect 6205 75 6240 175
rect 6260 75 6295 175
rect 6455 75 6490 175
rect 6510 75 6545 175
rect 6705 75 6740 175
rect 6760 75 6795 175
rect 6955 75 6990 175
rect 7010 75 7045 175
rect 7205 75 7240 175
rect 7260 75 7295 175
rect 7455 75 7490 175
rect 7510 75 7545 175
rect 7705 75 7740 175
rect 7760 75 7795 175
rect 7955 75 7990 175
rect 75 10 175 45
rect 325 10 425 45
rect 575 10 675 45
rect 825 10 925 45
rect 1075 10 1175 45
rect 1325 10 1425 45
rect 1575 10 1675 45
rect 1825 10 1925 45
rect 2075 10 2175 45
rect 2325 10 2425 45
rect 2575 10 2675 45
rect 2825 10 2925 45
rect 3075 10 3175 45
rect 3325 10 3425 45
rect 3575 10 3675 45
rect 3825 10 3925 45
rect 4075 10 4175 45
rect 4325 10 4425 45
rect 4575 10 4675 45
rect 4825 10 4925 45
rect 5075 10 5175 45
rect 5325 10 5425 45
rect 5575 10 5675 45
rect 5825 10 5925 45
rect 6075 10 6175 45
rect 6325 10 6425 45
rect 6575 10 6675 45
rect 6825 10 6925 45
rect 7075 10 7175 45
rect 7325 10 7425 45
rect 7575 10 7675 45
rect 7825 10 7925 45
<< metal3 >>
rect 0 7990 8000 8000
rect 0 7955 75 7990
rect 175 7955 325 7990
rect 425 7955 575 7990
rect 675 7955 825 7990
rect 925 7955 1075 7990
rect 1175 7955 1325 7990
rect 1425 7955 1575 7990
rect 1675 7955 1825 7990
rect 1925 7955 2075 7990
rect 2175 7955 2325 7990
rect 2425 7955 2575 7990
rect 2675 7955 2825 7990
rect 2925 7955 3075 7990
rect 3175 7955 3325 7990
rect 3425 7955 3575 7990
rect 3675 7955 3825 7990
rect 3925 7955 4075 7990
rect 4175 7955 4325 7990
rect 4425 7955 4575 7990
rect 4675 7955 4825 7990
rect 4925 7955 5075 7990
rect 5175 7955 5325 7990
rect 5425 7955 5575 7990
rect 5675 7955 5825 7990
rect 5925 7955 6075 7990
rect 6175 7955 6325 7990
rect 6425 7955 6575 7990
rect 6675 7955 6825 7990
rect 6925 7955 7075 7990
rect 7175 7955 7325 7990
rect 7425 7955 7575 7990
rect 7675 7955 7825 7990
rect 7925 7955 8000 7990
rect 0 7950 8000 7955
rect 0 7940 60 7950
rect 190 7940 310 7950
rect 440 7940 560 7950
rect 690 7940 810 7950
rect 940 7940 1060 7950
rect 1190 7940 1310 7950
rect 1440 7940 1560 7950
rect 1690 7940 1810 7950
rect 1940 7940 2060 7950
rect 2190 7940 2310 7950
rect 2440 7940 2560 7950
rect 2690 7940 2810 7950
rect 2940 7940 3060 7950
rect 3190 7940 3310 7950
rect 3440 7940 3560 7950
rect 3690 7940 3810 7950
rect 3940 7940 4060 7950
rect 4190 7940 4310 7950
rect 4440 7940 4560 7950
rect 4690 7940 4810 7950
rect 4940 7940 5060 7950
rect 5190 7940 5310 7950
rect 5440 7940 5560 7950
rect 5690 7940 5810 7950
rect 5940 7940 6060 7950
rect 6190 7940 6310 7950
rect 6440 7940 6560 7950
rect 6690 7940 6810 7950
rect 6940 7940 7060 7950
rect 7190 7940 7310 7950
rect 7440 7940 7560 7950
rect 7690 7940 7810 7950
rect 7940 7940 8000 7950
rect 0 7925 50 7940
rect 0 7825 10 7925
rect 45 7825 50 7925
rect 0 7810 50 7825
rect 200 7925 300 7940
rect 200 7825 205 7925
rect 240 7825 260 7925
rect 295 7825 300 7925
rect 200 7810 300 7825
rect 450 7925 550 7940
rect 450 7825 455 7925
rect 490 7825 510 7925
rect 545 7825 550 7925
rect 450 7810 550 7825
rect 700 7925 800 7940
rect 700 7825 705 7925
rect 740 7825 760 7925
rect 795 7825 800 7925
rect 700 7810 800 7825
rect 950 7925 1050 7940
rect 950 7825 955 7925
rect 990 7825 1010 7925
rect 1045 7825 1050 7925
rect 950 7810 1050 7825
rect 1200 7925 1300 7940
rect 1200 7825 1205 7925
rect 1240 7825 1260 7925
rect 1295 7825 1300 7925
rect 1200 7810 1300 7825
rect 1450 7925 1550 7940
rect 1450 7825 1455 7925
rect 1490 7825 1510 7925
rect 1545 7825 1550 7925
rect 1450 7810 1550 7825
rect 1700 7925 1800 7940
rect 1700 7825 1705 7925
rect 1740 7825 1760 7925
rect 1795 7825 1800 7925
rect 1700 7810 1800 7825
rect 1950 7925 2050 7940
rect 1950 7825 1955 7925
rect 1990 7825 2010 7925
rect 2045 7825 2050 7925
rect 1950 7810 2050 7825
rect 2200 7925 2300 7940
rect 2200 7825 2205 7925
rect 2240 7825 2260 7925
rect 2295 7825 2300 7925
rect 2200 7810 2300 7825
rect 2450 7925 2550 7940
rect 2450 7825 2455 7925
rect 2490 7825 2510 7925
rect 2545 7825 2550 7925
rect 2450 7810 2550 7825
rect 2700 7925 2800 7940
rect 2700 7825 2705 7925
rect 2740 7825 2760 7925
rect 2795 7825 2800 7925
rect 2700 7810 2800 7825
rect 2950 7925 3050 7940
rect 2950 7825 2955 7925
rect 2990 7825 3010 7925
rect 3045 7825 3050 7925
rect 2950 7810 3050 7825
rect 3200 7925 3300 7940
rect 3200 7825 3205 7925
rect 3240 7825 3260 7925
rect 3295 7825 3300 7925
rect 3200 7810 3300 7825
rect 3450 7925 3550 7940
rect 3450 7825 3455 7925
rect 3490 7825 3510 7925
rect 3545 7825 3550 7925
rect 3450 7810 3550 7825
rect 3700 7925 3800 7940
rect 3700 7825 3705 7925
rect 3740 7825 3760 7925
rect 3795 7825 3800 7925
rect 3700 7810 3800 7825
rect 3950 7925 4050 7940
rect 3950 7825 3955 7925
rect 3990 7825 4010 7925
rect 4045 7825 4050 7925
rect 3950 7810 4050 7825
rect 4200 7925 4300 7940
rect 4200 7825 4205 7925
rect 4240 7825 4260 7925
rect 4295 7825 4300 7925
rect 4200 7810 4300 7825
rect 4450 7925 4550 7940
rect 4450 7825 4455 7925
rect 4490 7825 4510 7925
rect 4545 7825 4550 7925
rect 4450 7810 4550 7825
rect 4700 7925 4800 7940
rect 4700 7825 4705 7925
rect 4740 7825 4760 7925
rect 4795 7825 4800 7925
rect 4700 7810 4800 7825
rect 4950 7925 5050 7940
rect 4950 7825 4955 7925
rect 4990 7825 5010 7925
rect 5045 7825 5050 7925
rect 4950 7810 5050 7825
rect 5200 7925 5300 7940
rect 5200 7825 5205 7925
rect 5240 7825 5260 7925
rect 5295 7825 5300 7925
rect 5200 7810 5300 7825
rect 5450 7925 5550 7940
rect 5450 7825 5455 7925
rect 5490 7825 5510 7925
rect 5545 7825 5550 7925
rect 5450 7810 5550 7825
rect 5700 7925 5800 7940
rect 5700 7825 5705 7925
rect 5740 7825 5760 7925
rect 5795 7825 5800 7925
rect 5700 7810 5800 7825
rect 5950 7925 6050 7940
rect 5950 7825 5955 7925
rect 5990 7825 6010 7925
rect 6045 7825 6050 7925
rect 5950 7810 6050 7825
rect 6200 7925 6300 7940
rect 6200 7825 6205 7925
rect 6240 7825 6260 7925
rect 6295 7825 6300 7925
rect 6200 7810 6300 7825
rect 6450 7925 6550 7940
rect 6450 7825 6455 7925
rect 6490 7825 6510 7925
rect 6545 7825 6550 7925
rect 6450 7810 6550 7825
rect 6700 7925 6800 7940
rect 6700 7825 6705 7925
rect 6740 7825 6760 7925
rect 6795 7825 6800 7925
rect 6700 7810 6800 7825
rect 6950 7925 7050 7940
rect 6950 7825 6955 7925
rect 6990 7825 7010 7925
rect 7045 7825 7050 7925
rect 6950 7810 7050 7825
rect 7200 7925 7300 7940
rect 7200 7825 7205 7925
rect 7240 7825 7260 7925
rect 7295 7825 7300 7925
rect 7200 7810 7300 7825
rect 7450 7925 7550 7940
rect 7450 7825 7455 7925
rect 7490 7825 7510 7925
rect 7545 7825 7550 7925
rect 7450 7810 7550 7825
rect 7700 7925 7800 7940
rect 7700 7825 7705 7925
rect 7740 7825 7760 7925
rect 7795 7825 7800 7925
rect 7700 7810 7800 7825
rect 7950 7925 8000 7940
rect 7950 7825 7955 7925
rect 7990 7825 8000 7925
rect 7950 7810 8000 7825
rect 0 7800 60 7810
rect 190 7800 310 7810
rect 440 7800 560 7810
rect 690 7800 810 7810
rect 940 7800 1060 7810
rect 1190 7800 1310 7810
rect 1440 7800 1560 7810
rect 1690 7800 1810 7810
rect 1940 7800 2060 7810
rect 2190 7800 2310 7810
rect 2440 7800 2560 7810
rect 2690 7800 2810 7810
rect 2940 7800 3060 7810
rect 3190 7800 3310 7810
rect 3440 7800 3560 7810
rect 3690 7800 3810 7810
rect 3940 7800 4060 7810
rect 4190 7800 4310 7810
rect 4440 7800 4560 7810
rect 4690 7800 4810 7810
rect 4940 7800 5060 7810
rect 5190 7800 5310 7810
rect 5440 7800 5560 7810
rect 5690 7800 5810 7810
rect 5940 7800 6060 7810
rect 6190 7800 6310 7810
rect 6440 7800 6560 7810
rect 6690 7800 6810 7810
rect 6940 7800 7060 7810
rect 7190 7800 7310 7810
rect 7440 7800 7560 7810
rect 7690 7800 7810 7810
rect 7940 7800 8000 7810
rect 0 7795 200 7800
rect 0 7760 75 7795
rect 175 7760 200 7795
rect 0 7740 200 7760
rect 0 7705 75 7740
rect 175 7705 200 7740
rect 0 7700 200 7705
rect 300 7795 450 7800
rect 300 7760 325 7795
rect 425 7760 450 7795
rect 300 7740 450 7760
rect 300 7705 325 7740
rect 425 7705 450 7740
rect 300 7700 450 7705
rect 550 7795 700 7800
rect 550 7760 575 7795
rect 675 7760 700 7795
rect 550 7740 700 7760
rect 550 7705 575 7740
rect 675 7705 700 7740
rect 550 7700 700 7705
rect 800 7795 1200 7800
rect 800 7760 825 7795
rect 925 7760 1075 7795
rect 1175 7760 1200 7795
rect 800 7740 1200 7760
rect 800 7705 825 7740
rect 925 7705 1075 7740
rect 1175 7705 1200 7740
rect 800 7700 1200 7705
rect 1300 7795 1450 7800
rect 1300 7760 1325 7795
rect 1425 7760 1450 7795
rect 1300 7740 1450 7760
rect 1300 7705 1325 7740
rect 1425 7705 1450 7740
rect 1300 7700 1450 7705
rect 1550 7795 1700 7800
rect 1550 7760 1575 7795
rect 1675 7760 1700 7795
rect 1550 7740 1700 7760
rect 1550 7705 1575 7740
rect 1675 7705 1700 7740
rect 1550 7700 1700 7705
rect 1800 7795 2200 7800
rect 1800 7760 1825 7795
rect 1925 7760 2075 7795
rect 2175 7760 2200 7795
rect 1800 7740 2200 7760
rect 1800 7705 1825 7740
rect 1925 7705 2075 7740
rect 2175 7705 2200 7740
rect 1800 7700 2200 7705
rect 2300 7795 2450 7800
rect 2300 7760 2325 7795
rect 2425 7760 2450 7795
rect 2300 7740 2450 7760
rect 2300 7705 2325 7740
rect 2425 7705 2450 7740
rect 2300 7700 2450 7705
rect 2550 7795 2700 7800
rect 2550 7760 2575 7795
rect 2675 7760 2700 7795
rect 2550 7740 2700 7760
rect 2550 7705 2575 7740
rect 2675 7705 2700 7740
rect 2550 7700 2700 7705
rect 2800 7795 3200 7800
rect 2800 7760 2825 7795
rect 2925 7760 3075 7795
rect 3175 7760 3200 7795
rect 2800 7740 3200 7760
rect 2800 7705 2825 7740
rect 2925 7705 3075 7740
rect 3175 7705 3200 7740
rect 2800 7700 3200 7705
rect 3300 7795 3450 7800
rect 3300 7760 3325 7795
rect 3425 7760 3450 7795
rect 3300 7740 3450 7760
rect 3300 7705 3325 7740
rect 3425 7705 3450 7740
rect 3300 7700 3450 7705
rect 3550 7795 3700 7800
rect 3550 7760 3575 7795
rect 3675 7760 3700 7795
rect 3550 7740 3700 7760
rect 3550 7705 3575 7740
rect 3675 7705 3700 7740
rect 3550 7700 3700 7705
rect 3800 7795 4200 7800
rect 3800 7760 3825 7795
rect 3925 7760 4075 7795
rect 4175 7760 4200 7795
rect 3800 7740 4200 7760
rect 3800 7705 3825 7740
rect 3925 7705 4075 7740
rect 4175 7705 4200 7740
rect 3800 7700 4200 7705
rect 4300 7795 4450 7800
rect 4300 7760 4325 7795
rect 4425 7760 4450 7795
rect 4300 7740 4450 7760
rect 4300 7705 4325 7740
rect 4425 7705 4450 7740
rect 4300 7700 4450 7705
rect 4550 7795 4700 7800
rect 4550 7760 4575 7795
rect 4675 7760 4700 7795
rect 4550 7740 4700 7760
rect 4550 7705 4575 7740
rect 4675 7705 4700 7740
rect 4550 7700 4700 7705
rect 4800 7795 5200 7800
rect 4800 7760 4825 7795
rect 4925 7760 5075 7795
rect 5175 7760 5200 7795
rect 4800 7740 5200 7760
rect 4800 7705 4825 7740
rect 4925 7705 5075 7740
rect 5175 7705 5200 7740
rect 4800 7700 5200 7705
rect 5300 7795 5450 7800
rect 5300 7760 5325 7795
rect 5425 7760 5450 7795
rect 5300 7740 5450 7760
rect 5300 7705 5325 7740
rect 5425 7705 5450 7740
rect 5300 7700 5450 7705
rect 5550 7795 5700 7800
rect 5550 7760 5575 7795
rect 5675 7760 5700 7795
rect 5550 7740 5700 7760
rect 5550 7705 5575 7740
rect 5675 7705 5700 7740
rect 5550 7700 5700 7705
rect 5800 7795 6200 7800
rect 5800 7760 5825 7795
rect 5925 7760 6075 7795
rect 6175 7760 6200 7795
rect 5800 7740 6200 7760
rect 5800 7705 5825 7740
rect 5925 7705 6075 7740
rect 6175 7705 6200 7740
rect 5800 7700 6200 7705
rect 6300 7795 6450 7800
rect 6300 7760 6325 7795
rect 6425 7760 6450 7795
rect 6300 7740 6450 7760
rect 6300 7705 6325 7740
rect 6425 7705 6450 7740
rect 6300 7700 6450 7705
rect 6550 7795 6700 7800
rect 6550 7760 6575 7795
rect 6675 7760 6700 7795
rect 6550 7740 6700 7760
rect 6550 7705 6575 7740
rect 6675 7705 6700 7740
rect 6550 7700 6700 7705
rect 6800 7795 7200 7800
rect 6800 7760 6825 7795
rect 6925 7760 7075 7795
rect 7175 7760 7200 7795
rect 6800 7740 7200 7760
rect 6800 7705 6825 7740
rect 6925 7705 7075 7740
rect 7175 7705 7200 7740
rect 6800 7700 7200 7705
rect 7300 7795 7450 7800
rect 7300 7760 7325 7795
rect 7425 7760 7450 7795
rect 7300 7740 7450 7760
rect 7300 7705 7325 7740
rect 7425 7705 7450 7740
rect 7300 7700 7450 7705
rect 7550 7795 7700 7800
rect 7550 7760 7575 7795
rect 7675 7760 7700 7795
rect 7550 7740 7700 7760
rect 7550 7705 7575 7740
rect 7675 7705 7700 7740
rect 7550 7700 7700 7705
rect 7800 7795 8000 7800
rect 7800 7760 7825 7795
rect 7925 7760 8000 7795
rect 7800 7740 8000 7760
rect 7800 7705 7825 7740
rect 7925 7705 8000 7740
rect 7800 7700 8000 7705
rect 0 7690 60 7700
rect 190 7690 310 7700
rect 440 7690 560 7700
rect 690 7690 810 7700
rect 940 7690 1060 7700
rect 1190 7690 1310 7700
rect 1440 7690 1560 7700
rect 1690 7690 1810 7700
rect 1940 7690 2060 7700
rect 2190 7690 2310 7700
rect 2440 7690 2560 7700
rect 2690 7690 2810 7700
rect 2940 7690 3060 7700
rect 3190 7690 3310 7700
rect 3440 7690 3560 7700
rect 3690 7690 3810 7700
rect 3940 7690 4060 7700
rect 4190 7690 4310 7700
rect 4440 7690 4560 7700
rect 4690 7690 4810 7700
rect 4940 7690 5060 7700
rect 5190 7690 5310 7700
rect 5440 7690 5560 7700
rect 5690 7690 5810 7700
rect 5940 7690 6060 7700
rect 6190 7690 6310 7700
rect 6440 7690 6560 7700
rect 6690 7690 6810 7700
rect 6940 7690 7060 7700
rect 7190 7690 7310 7700
rect 7440 7690 7560 7700
rect 7690 7690 7810 7700
rect 7940 7690 8000 7700
rect 0 7675 50 7690
rect 0 7575 10 7675
rect 45 7575 50 7675
rect 0 7560 50 7575
rect 200 7675 300 7690
rect 200 7575 205 7675
rect 240 7575 260 7675
rect 295 7575 300 7675
rect 200 7560 300 7575
rect 450 7675 550 7690
rect 450 7575 455 7675
rect 490 7575 510 7675
rect 545 7575 550 7675
rect 450 7560 550 7575
rect 700 7675 800 7690
rect 700 7575 705 7675
rect 740 7575 760 7675
rect 795 7575 800 7675
rect 700 7560 800 7575
rect 950 7675 1050 7690
rect 950 7575 955 7675
rect 990 7575 1010 7675
rect 1045 7575 1050 7675
rect 950 7560 1050 7575
rect 1200 7675 1300 7690
rect 1200 7575 1205 7675
rect 1240 7575 1260 7675
rect 1295 7575 1300 7675
rect 1200 7560 1300 7575
rect 1450 7675 1550 7690
rect 1450 7575 1455 7675
rect 1490 7575 1510 7675
rect 1545 7575 1550 7675
rect 1450 7560 1550 7575
rect 1700 7675 1800 7690
rect 1700 7575 1705 7675
rect 1740 7575 1760 7675
rect 1795 7575 1800 7675
rect 1700 7560 1800 7575
rect 1950 7675 2050 7690
rect 1950 7575 1955 7675
rect 1990 7575 2010 7675
rect 2045 7575 2050 7675
rect 1950 7560 2050 7575
rect 2200 7675 2300 7690
rect 2200 7575 2205 7675
rect 2240 7575 2260 7675
rect 2295 7575 2300 7675
rect 2200 7560 2300 7575
rect 2450 7675 2550 7690
rect 2450 7575 2455 7675
rect 2490 7575 2510 7675
rect 2545 7575 2550 7675
rect 2450 7560 2550 7575
rect 2700 7675 2800 7690
rect 2700 7575 2705 7675
rect 2740 7575 2760 7675
rect 2795 7575 2800 7675
rect 2700 7560 2800 7575
rect 2950 7675 3050 7690
rect 2950 7575 2955 7675
rect 2990 7575 3010 7675
rect 3045 7575 3050 7675
rect 2950 7560 3050 7575
rect 3200 7675 3300 7690
rect 3200 7575 3205 7675
rect 3240 7575 3260 7675
rect 3295 7575 3300 7675
rect 3200 7560 3300 7575
rect 3450 7675 3550 7690
rect 3450 7575 3455 7675
rect 3490 7575 3510 7675
rect 3545 7575 3550 7675
rect 3450 7560 3550 7575
rect 3700 7675 3800 7690
rect 3700 7575 3705 7675
rect 3740 7575 3760 7675
rect 3795 7575 3800 7675
rect 3700 7560 3800 7575
rect 3950 7675 4050 7690
rect 3950 7575 3955 7675
rect 3990 7575 4010 7675
rect 4045 7575 4050 7675
rect 3950 7560 4050 7575
rect 4200 7675 4300 7690
rect 4200 7575 4205 7675
rect 4240 7575 4260 7675
rect 4295 7575 4300 7675
rect 4200 7560 4300 7575
rect 4450 7675 4550 7690
rect 4450 7575 4455 7675
rect 4490 7575 4510 7675
rect 4545 7575 4550 7675
rect 4450 7560 4550 7575
rect 4700 7675 4800 7690
rect 4700 7575 4705 7675
rect 4740 7575 4760 7675
rect 4795 7575 4800 7675
rect 4700 7560 4800 7575
rect 4950 7675 5050 7690
rect 4950 7575 4955 7675
rect 4990 7575 5010 7675
rect 5045 7575 5050 7675
rect 4950 7560 5050 7575
rect 5200 7675 5300 7690
rect 5200 7575 5205 7675
rect 5240 7575 5260 7675
rect 5295 7575 5300 7675
rect 5200 7560 5300 7575
rect 5450 7675 5550 7690
rect 5450 7575 5455 7675
rect 5490 7575 5510 7675
rect 5545 7575 5550 7675
rect 5450 7560 5550 7575
rect 5700 7675 5800 7690
rect 5700 7575 5705 7675
rect 5740 7575 5760 7675
rect 5795 7575 5800 7675
rect 5700 7560 5800 7575
rect 5950 7675 6050 7690
rect 5950 7575 5955 7675
rect 5990 7575 6010 7675
rect 6045 7575 6050 7675
rect 5950 7560 6050 7575
rect 6200 7675 6300 7690
rect 6200 7575 6205 7675
rect 6240 7575 6260 7675
rect 6295 7575 6300 7675
rect 6200 7560 6300 7575
rect 6450 7675 6550 7690
rect 6450 7575 6455 7675
rect 6490 7575 6510 7675
rect 6545 7575 6550 7675
rect 6450 7560 6550 7575
rect 6700 7675 6800 7690
rect 6700 7575 6705 7675
rect 6740 7575 6760 7675
rect 6795 7575 6800 7675
rect 6700 7560 6800 7575
rect 6950 7675 7050 7690
rect 6950 7575 6955 7675
rect 6990 7575 7010 7675
rect 7045 7575 7050 7675
rect 6950 7560 7050 7575
rect 7200 7675 7300 7690
rect 7200 7575 7205 7675
rect 7240 7575 7260 7675
rect 7295 7575 7300 7675
rect 7200 7560 7300 7575
rect 7450 7675 7550 7690
rect 7450 7575 7455 7675
rect 7490 7575 7510 7675
rect 7545 7575 7550 7675
rect 7450 7560 7550 7575
rect 7700 7675 7800 7690
rect 7700 7575 7705 7675
rect 7740 7575 7760 7675
rect 7795 7575 7800 7675
rect 7700 7560 7800 7575
rect 7950 7675 8000 7690
rect 7950 7575 7955 7675
rect 7990 7575 8000 7675
rect 7950 7560 8000 7575
rect 0 7550 60 7560
rect 190 7550 310 7560
rect 440 7550 560 7560
rect 690 7550 810 7560
rect 940 7550 1060 7560
rect 1190 7550 1310 7560
rect 1440 7550 1560 7560
rect 1690 7550 1810 7560
rect 1940 7550 2060 7560
rect 2190 7550 2310 7560
rect 2440 7550 2560 7560
rect 2690 7550 2810 7560
rect 2940 7550 3060 7560
rect 3190 7550 3310 7560
rect 3440 7550 3560 7560
rect 3690 7550 3810 7560
rect 3940 7550 4060 7560
rect 4190 7550 4310 7560
rect 4440 7550 4560 7560
rect 4690 7550 4810 7560
rect 4940 7550 5060 7560
rect 5190 7550 5310 7560
rect 5440 7550 5560 7560
rect 5690 7550 5810 7560
rect 5940 7550 6060 7560
rect 6190 7550 6310 7560
rect 6440 7550 6560 7560
rect 6690 7550 6810 7560
rect 6940 7550 7060 7560
rect 7190 7550 7310 7560
rect 7440 7550 7560 7560
rect 7690 7550 7810 7560
rect 7940 7550 8000 7560
rect 0 7545 200 7550
rect 0 7510 75 7545
rect 175 7510 200 7545
rect 0 7490 200 7510
rect 0 7455 75 7490
rect 175 7455 200 7490
rect 0 7450 200 7455
rect 300 7545 450 7550
rect 300 7510 325 7545
rect 425 7510 450 7545
rect 300 7490 450 7510
rect 300 7455 325 7490
rect 425 7455 450 7490
rect 300 7450 450 7455
rect 550 7545 700 7550
rect 550 7510 575 7545
rect 675 7510 700 7545
rect 550 7490 700 7510
rect 550 7455 575 7490
rect 675 7455 700 7490
rect 550 7450 700 7455
rect 800 7545 950 7550
rect 800 7510 825 7545
rect 925 7510 950 7545
rect 800 7490 950 7510
rect 800 7455 825 7490
rect 925 7455 950 7490
rect 800 7450 950 7455
rect 1050 7545 1200 7550
rect 1050 7510 1075 7545
rect 1175 7510 1200 7545
rect 1050 7490 1200 7510
rect 1050 7455 1075 7490
rect 1175 7455 1200 7490
rect 1050 7450 1200 7455
rect 1300 7545 1450 7550
rect 1300 7510 1325 7545
rect 1425 7510 1450 7545
rect 1300 7490 1450 7510
rect 1300 7455 1325 7490
rect 1425 7455 1450 7490
rect 1300 7450 1450 7455
rect 1550 7545 1700 7550
rect 1550 7510 1575 7545
rect 1675 7510 1700 7545
rect 1550 7490 1700 7510
rect 1550 7455 1575 7490
rect 1675 7455 1700 7490
rect 1550 7450 1700 7455
rect 1800 7545 2200 7550
rect 1800 7510 1825 7545
rect 1925 7510 2075 7545
rect 2175 7510 2200 7545
rect 1800 7490 2200 7510
rect 1800 7455 1825 7490
rect 1925 7455 2075 7490
rect 2175 7455 2200 7490
rect 1800 7450 2200 7455
rect 2300 7545 2450 7550
rect 2300 7510 2325 7545
rect 2425 7510 2450 7545
rect 2300 7490 2450 7510
rect 2300 7455 2325 7490
rect 2425 7455 2450 7490
rect 2300 7450 2450 7455
rect 2550 7545 2700 7550
rect 2550 7510 2575 7545
rect 2675 7510 2700 7545
rect 2550 7490 2700 7510
rect 2550 7455 2575 7490
rect 2675 7455 2700 7490
rect 2550 7450 2700 7455
rect 2800 7545 2950 7550
rect 2800 7510 2825 7545
rect 2925 7510 2950 7545
rect 2800 7490 2950 7510
rect 2800 7455 2825 7490
rect 2925 7455 2950 7490
rect 2800 7450 2950 7455
rect 3050 7545 3200 7550
rect 3050 7510 3075 7545
rect 3175 7510 3200 7545
rect 3050 7490 3200 7510
rect 3050 7455 3075 7490
rect 3175 7455 3200 7490
rect 3050 7450 3200 7455
rect 3300 7545 3450 7550
rect 3300 7510 3325 7545
rect 3425 7510 3450 7545
rect 3300 7490 3450 7510
rect 3300 7455 3325 7490
rect 3425 7455 3450 7490
rect 3300 7450 3450 7455
rect 3550 7545 3700 7550
rect 3550 7510 3575 7545
rect 3675 7510 3700 7545
rect 3550 7490 3700 7510
rect 3550 7455 3575 7490
rect 3675 7455 3700 7490
rect 3550 7450 3700 7455
rect 3800 7545 4200 7550
rect 3800 7510 3825 7545
rect 3925 7510 4075 7545
rect 4175 7510 4200 7545
rect 3800 7490 4200 7510
rect 3800 7455 3825 7490
rect 3925 7455 4075 7490
rect 4175 7455 4200 7490
rect 3800 7450 4200 7455
rect 4300 7545 4450 7550
rect 4300 7510 4325 7545
rect 4425 7510 4450 7545
rect 4300 7490 4450 7510
rect 4300 7455 4325 7490
rect 4425 7455 4450 7490
rect 4300 7450 4450 7455
rect 4550 7545 4700 7550
rect 4550 7510 4575 7545
rect 4675 7510 4700 7545
rect 4550 7490 4700 7510
rect 4550 7455 4575 7490
rect 4675 7455 4700 7490
rect 4550 7450 4700 7455
rect 4800 7545 4950 7550
rect 4800 7510 4825 7545
rect 4925 7510 4950 7545
rect 4800 7490 4950 7510
rect 4800 7455 4825 7490
rect 4925 7455 4950 7490
rect 4800 7450 4950 7455
rect 5050 7545 5200 7550
rect 5050 7510 5075 7545
rect 5175 7510 5200 7545
rect 5050 7490 5200 7510
rect 5050 7455 5075 7490
rect 5175 7455 5200 7490
rect 5050 7450 5200 7455
rect 5300 7545 5450 7550
rect 5300 7510 5325 7545
rect 5425 7510 5450 7545
rect 5300 7490 5450 7510
rect 5300 7455 5325 7490
rect 5425 7455 5450 7490
rect 5300 7450 5450 7455
rect 5550 7545 5700 7550
rect 5550 7510 5575 7545
rect 5675 7510 5700 7545
rect 5550 7490 5700 7510
rect 5550 7455 5575 7490
rect 5675 7455 5700 7490
rect 5550 7450 5700 7455
rect 5800 7545 6200 7550
rect 5800 7510 5825 7545
rect 5925 7510 6075 7545
rect 6175 7510 6200 7545
rect 5800 7490 6200 7510
rect 5800 7455 5825 7490
rect 5925 7455 6075 7490
rect 6175 7455 6200 7490
rect 5800 7450 6200 7455
rect 6300 7545 6450 7550
rect 6300 7510 6325 7545
rect 6425 7510 6450 7545
rect 6300 7490 6450 7510
rect 6300 7455 6325 7490
rect 6425 7455 6450 7490
rect 6300 7450 6450 7455
rect 6550 7545 6700 7550
rect 6550 7510 6575 7545
rect 6675 7510 6700 7545
rect 6550 7490 6700 7510
rect 6550 7455 6575 7490
rect 6675 7455 6700 7490
rect 6550 7450 6700 7455
rect 6800 7545 6950 7550
rect 6800 7510 6825 7545
rect 6925 7510 6950 7545
rect 6800 7490 6950 7510
rect 6800 7455 6825 7490
rect 6925 7455 6950 7490
rect 6800 7450 6950 7455
rect 7050 7545 7200 7550
rect 7050 7510 7075 7545
rect 7175 7510 7200 7545
rect 7050 7490 7200 7510
rect 7050 7455 7075 7490
rect 7175 7455 7200 7490
rect 7050 7450 7200 7455
rect 7300 7545 7450 7550
rect 7300 7510 7325 7545
rect 7425 7510 7450 7545
rect 7300 7490 7450 7510
rect 7300 7455 7325 7490
rect 7425 7455 7450 7490
rect 7300 7450 7450 7455
rect 7550 7545 7700 7550
rect 7550 7510 7575 7545
rect 7675 7510 7700 7545
rect 7550 7490 7700 7510
rect 7550 7455 7575 7490
rect 7675 7455 7700 7490
rect 7550 7450 7700 7455
rect 7800 7545 8000 7550
rect 7800 7510 7825 7545
rect 7925 7510 8000 7545
rect 7800 7490 8000 7510
rect 7800 7455 7825 7490
rect 7925 7455 8000 7490
rect 7800 7450 8000 7455
rect 0 7440 60 7450
rect 190 7440 310 7450
rect 440 7440 560 7450
rect 690 7440 810 7450
rect 940 7440 1060 7450
rect 1190 7440 1310 7450
rect 1440 7440 1560 7450
rect 1690 7440 1810 7450
rect 1940 7440 2060 7450
rect 2190 7440 2310 7450
rect 2440 7440 2560 7450
rect 2690 7440 2810 7450
rect 2940 7440 3060 7450
rect 3190 7440 3310 7450
rect 3440 7440 3560 7450
rect 3690 7440 3810 7450
rect 3940 7440 4060 7450
rect 4190 7440 4310 7450
rect 4440 7440 4560 7450
rect 4690 7440 4810 7450
rect 4940 7440 5060 7450
rect 5190 7440 5310 7450
rect 5440 7440 5560 7450
rect 5690 7440 5810 7450
rect 5940 7440 6060 7450
rect 6190 7440 6310 7450
rect 6440 7440 6560 7450
rect 6690 7440 6810 7450
rect 6940 7440 7060 7450
rect 7190 7440 7310 7450
rect 7440 7440 7560 7450
rect 7690 7440 7810 7450
rect 7940 7440 8000 7450
rect 0 7425 50 7440
rect 0 7325 10 7425
rect 45 7325 50 7425
rect 0 7310 50 7325
rect 200 7425 300 7440
rect 200 7325 205 7425
rect 240 7325 260 7425
rect 295 7325 300 7425
rect 200 7310 300 7325
rect 450 7425 550 7440
rect 450 7325 455 7425
rect 490 7325 510 7425
rect 545 7325 550 7425
rect 450 7310 550 7325
rect 700 7425 800 7440
rect 700 7325 705 7425
rect 740 7325 760 7425
rect 795 7325 800 7425
rect 700 7310 800 7325
rect 950 7425 1050 7440
rect 950 7325 955 7425
rect 990 7325 1010 7425
rect 1045 7325 1050 7425
rect 950 7310 1050 7325
rect 1200 7425 1300 7440
rect 1200 7325 1205 7425
rect 1240 7325 1260 7425
rect 1295 7325 1300 7425
rect 1200 7310 1300 7325
rect 1450 7425 1550 7440
rect 1450 7325 1455 7425
rect 1490 7325 1510 7425
rect 1545 7325 1550 7425
rect 1450 7310 1550 7325
rect 1700 7425 1800 7440
rect 1700 7325 1705 7425
rect 1740 7325 1760 7425
rect 1795 7325 1800 7425
rect 1700 7310 1800 7325
rect 1950 7425 2050 7440
rect 1950 7325 1955 7425
rect 1990 7325 2010 7425
rect 2045 7325 2050 7425
rect 1950 7310 2050 7325
rect 2200 7425 2300 7440
rect 2200 7325 2205 7425
rect 2240 7325 2260 7425
rect 2295 7325 2300 7425
rect 2200 7310 2300 7325
rect 2450 7425 2550 7440
rect 2450 7325 2455 7425
rect 2490 7325 2510 7425
rect 2545 7325 2550 7425
rect 2450 7310 2550 7325
rect 2700 7425 2800 7440
rect 2700 7325 2705 7425
rect 2740 7325 2760 7425
rect 2795 7325 2800 7425
rect 2700 7310 2800 7325
rect 2950 7425 3050 7440
rect 2950 7325 2955 7425
rect 2990 7325 3010 7425
rect 3045 7325 3050 7425
rect 2950 7310 3050 7325
rect 3200 7425 3300 7440
rect 3200 7325 3205 7425
rect 3240 7325 3260 7425
rect 3295 7325 3300 7425
rect 3200 7310 3300 7325
rect 3450 7425 3550 7440
rect 3450 7325 3455 7425
rect 3490 7325 3510 7425
rect 3545 7325 3550 7425
rect 3450 7310 3550 7325
rect 3700 7425 3800 7440
rect 3700 7325 3705 7425
rect 3740 7325 3760 7425
rect 3795 7325 3800 7425
rect 3700 7310 3800 7325
rect 3950 7425 4050 7440
rect 3950 7325 3955 7425
rect 3990 7325 4010 7425
rect 4045 7325 4050 7425
rect 3950 7310 4050 7325
rect 4200 7425 4300 7440
rect 4200 7325 4205 7425
rect 4240 7325 4260 7425
rect 4295 7325 4300 7425
rect 4200 7310 4300 7325
rect 4450 7425 4550 7440
rect 4450 7325 4455 7425
rect 4490 7325 4510 7425
rect 4545 7325 4550 7425
rect 4450 7310 4550 7325
rect 4700 7425 4800 7440
rect 4700 7325 4705 7425
rect 4740 7325 4760 7425
rect 4795 7325 4800 7425
rect 4700 7310 4800 7325
rect 4950 7425 5050 7440
rect 4950 7325 4955 7425
rect 4990 7325 5010 7425
rect 5045 7325 5050 7425
rect 4950 7310 5050 7325
rect 5200 7425 5300 7440
rect 5200 7325 5205 7425
rect 5240 7325 5260 7425
rect 5295 7325 5300 7425
rect 5200 7310 5300 7325
rect 5450 7425 5550 7440
rect 5450 7325 5455 7425
rect 5490 7325 5510 7425
rect 5545 7325 5550 7425
rect 5450 7310 5550 7325
rect 5700 7425 5800 7440
rect 5700 7325 5705 7425
rect 5740 7325 5760 7425
rect 5795 7325 5800 7425
rect 5700 7310 5800 7325
rect 5950 7425 6050 7440
rect 5950 7325 5955 7425
rect 5990 7325 6010 7425
rect 6045 7325 6050 7425
rect 5950 7310 6050 7325
rect 6200 7425 6300 7440
rect 6200 7325 6205 7425
rect 6240 7325 6260 7425
rect 6295 7325 6300 7425
rect 6200 7310 6300 7325
rect 6450 7425 6550 7440
rect 6450 7325 6455 7425
rect 6490 7325 6510 7425
rect 6545 7325 6550 7425
rect 6450 7310 6550 7325
rect 6700 7425 6800 7440
rect 6700 7325 6705 7425
rect 6740 7325 6760 7425
rect 6795 7325 6800 7425
rect 6700 7310 6800 7325
rect 6950 7425 7050 7440
rect 6950 7325 6955 7425
rect 6990 7325 7010 7425
rect 7045 7325 7050 7425
rect 6950 7310 7050 7325
rect 7200 7425 7300 7440
rect 7200 7325 7205 7425
rect 7240 7325 7260 7425
rect 7295 7325 7300 7425
rect 7200 7310 7300 7325
rect 7450 7425 7550 7440
rect 7450 7325 7455 7425
rect 7490 7325 7510 7425
rect 7545 7325 7550 7425
rect 7450 7310 7550 7325
rect 7700 7425 7800 7440
rect 7700 7325 7705 7425
rect 7740 7325 7760 7425
rect 7795 7325 7800 7425
rect 7700 7310 7800 7325
rect 7950 7425 8000 7440
rect 7950 7325 7955 7425
rect 7990 7325 8000 7425
rect 7950 7310 8000 7325
rect 0 7300 60 7310
rect 190 7300 310 7310
rect 440 7300 560 7310
rect 690 7300 810 7310
rect 940 7300 1060 7310
rect 1190 7300 1310 7310
rect 1440 7300 1560 7310
rect 1690 7300 1810 7310
rect 1940 7300 2060 7310
rect 2190 7300 2310 7310
rect 2440 7300 2560 7310
rect 2690 7300 2810 7310
rect 2940 7300 3060 7310
rect 3190 7300 3310 7310
rect 3440 7300 3560 7310
rect 3690 7300 3810 7310
rect 3940 7300 4060 7310
rect 4190 7300 4310 7310
rect 4440 7300 4560 7310
rect 4690 7300 4810 7310
rect 4940 7300 5060 7310
rect 5190 7300 5310 7310
rect 5440 7300 5560 7310
rect 5690 7300 5810 7310
rect 5940 7300 6060 7310
rect 6190 7300 6310 7310
rect 6440 7300 6560 7310
rect 6690 7300 6810 7310
rect 6940 7300 7060 7310
rect 7190 7300 7310 7310
rect 7440 7300 7560 7310
rect 7690 7300 7810 7310
rect 7940 7300 8000 7310
rect 0 7295 200 7300
rect 0 7260 75 7295
rect 175 7260 200 7295
rect 0 7240 200 7260
rect 0 7205 75 7240
rect 175 7205 200 7240
rect 0 7200 200 7205
rect 300 7295 450 7300
rect 300 7260 325 7295
rect 425 7260 450 7295
rect 300 7240 450 7260
rect 300 7205 325 7240
rect 425 7205 450 7240
rect 300 7200 450 7205
rect 550 7295 700 7300
rect 550 7260 575 7295
rect 675 7260 700 7295
rect 550 7240 700 7260
rect 550 7205 575 7240
rect 675 7205 700 7240
rect 550 7200 700 7205
rect 800 7295 1200 7300
rect 800 7260 825 7295
rect 925 7260 1075 7295
rect 1175 7260 1200 7295
rect 800 7240 1200 7260
rect 800 7205 825 7240
rect 925 7205 1075 7240
rect 1175 7205 1200 7240
rect 800 7200 1200 7205
rect 1300 7295 1450 7300
rect 1300 7260 1325 7295
rect 1425 7260 1450 7295
rect 1300 7240 1450 7260
rect 1300 7205 1325 7240
rect 1425 7205 1450 7240
rect 1300 7200 1450 7205
rect 1550 7295 1700 7300
rect 1550 7260 1575 7295
rect 1675 7260 1700 7295
rect 1550 7240 1700 7260
rect 1550 7205 1575 7240
rect 1675 7205 1700 7240
rect 1550 7200 1700 7205
rect 1800 7295 2200 7300
rect 1800 7260 1825 7295
rect 1925 7260 2075 7295
rect 2175 7260 2200 7295
rect 1800 7240 2200 7260
rect 1800 7205 1825 7240
rect 1925 7205 2075 7240
rect 2175 7205 2200 7240
rect 1800 7200 2200 7205
rect 2300 7295 2450 7300
rect 2300 7260 2325 7295
rect 2425 7260 2450 7295
rect 2300 7240 2450 7260
rect 2300 7205 2325 7240
rect 2425 7205 2450 7240
rect 2300 7200 2450 7205
rect 2550 7295 2700 7300
rect 2550 7260 2575 7295
rect 2675 7260 2700 7295
rect 2550 7240 2700 7260
rect 2550 7205 2575 7240
rect 2675 7205 2700 7240
rect 2550 7200 2700 7205
rect 2800 7295 3200 7300
rect 2800 7260 2825 7295
rect 2925 7260 3075 7295
rect 3175 7260 3200 7295
rect 2800 7240 3200 7260
rect 2800 7205 2825 7240
rect 2925 7205 3075 7240
rect 3175 7205 3200 7240
rect 2800 7200 3200 7205
rect 3300 7295 3450 7300
rect 3300 7260 3325 7295
rect 3425 7260 3450 7295
rect 3300 7240 3450 7260
rect 3300 7205 3325 7240
rect 3425 7205 3450 7240
rect 3300 7200 3450 7205
rect 3550 7295 3700 7300
rect 3550 7260 3575 7295
rect 3675 7260 3700 7295
rect 3550 7240 3700 7260
rect 3550 7205 3575 7240
rect 3675 7205 3700 7240
rect 3550 7200 3700 7205
rect 3800 7295 4200 7300
rect 3800 7260 3825 7295
rect 3925 7260 4075 7295
rect 4175 7260 4200 7295
rect 3800 7240 4200 7260
rect 3800 7205 3825 7240
rect 3925 7205 4075 7240
rect 4175 7205 4200 7240
rect 3800 7200 4200 7205
rect 4300 7295 4450 7300
rect 4300 7260 4325 7295
rect 4425 7260 4450 7295
rect 4300 7240 4450 7260
rect 4300 7205 4325 7240
rect 4425 7205 4450 7240
rect 4300 7200 4450 7205
rect 4550 7295 4700 7300
rect 4550 7260 4575 7295
rect 4675 7260 4700 7295
rect 4550 7240 4700 7260
rect 4550 7205 4575 7240
rect 4675 7205 4700 7240
rect 4550 7200 4700 7205
rect 4800 7295 5200 7300
rect 4800 7260 4825 7295
rect 4925 7260 5075 7295
rect 5175 7260 5200 7295
rect 4800 7240 5200 7260
rect 4800 7205 4825 7240
rect 4925 7205 5075 7240
rect 5175 7205 5200 7240
rect 4800 7200 5200 7205
rect 5300 7295 5450 7300
rect 5300 7260 5325 7295
rect 5425 7260 5450 7295
rect 5300 7240 5450 7260
rect 5300 7205 5325 7240
rect 5425 7205 5450 7240
rect 5300 7200 5450 7205
rect 5550 7295 5700 7300
rect 5550 7260 5575 7295
rect 5675 7260 5700 7295
rect 5550 7240 5700 7260
rect 5550 7205 5575 7240
rect 5675 7205 5700 7240
rect 5550 7200 5700 7205
rect 5800 7295 6200 7300
rect 5800 7260 5825 7295
rect 5925 7260 6075 7295
rect 6175 7260 6200 7295
rect 5800 7240 6200 7260
rect 5800 7205 5825 7240
rect 5925 7205 6075 7240
rect 6175 7205 6200 7240
rect 5800 7200 6200 7205
rect 6300 7295 6450 7300
rect 6300 7260 6325 7295
rect 6425 7260 6450 7295
rect 6300 7240 6450 7260
rect 6300 7205 6325 7240
rect 6425 7205 6450 7240
rect 6300 7200 6450 7205
rect 6550 7295 6700 7300
rect 6550 7260 6575 7295
rect 6675 7260 6700 7295
rect 6550 7240 6700 7260
rect 6550 7205 6575 7240
rect 6675 7205 6700 7240
rect 6550 7200 6700 7205
rect 6800 7295 7200 7300
rect 6800 7260 6825 7295
rect 6925 7260 7075 7295
rect 7175 7260 7200 7295
rect 6800 7240 7200 7260
rect 6800 7205 6825 7240
rect 6925 7205 7075 7240
rect 7175 7205 7200 7240
rect 6800 7200 7200 7205
rect 7300 7295 7450 7300
rect 7300 7260 7325 7295
rect 7425 7260 7450 7295
rect 7300 7240 7450 7260
rect 7300 7205 7325 7240
rect 7425 7205 7450 7240
rect 7300 7200 7450 7205
rect 7550 7295 7700 7300
rect 7550 7260 7575 7295
rect 7675 7260 7700 7295
rect 7550 7240 7700 7260
rect 7550 7205 7575 7240
rect 7675 7205 7700 7240
rect 7550 7200 7700 7205
rect 7800 7295 8000 7300
rect 7800 7260 7825 7295
rect 7925 7260 8000 7295
rect 7800 7240 8000 7260
rect 7800 7205 7825 7240
rect 7925 7205 8000 7240
rect 7800 7200 8000 7205
rect 0 7190 60 7200
rect 190 7190 310 7200
rect 440 7190 560 7200
rect 690 7190 810 7200
rect 940 7190 1060 7200
rect 1190 7190 1310 7200
rect 1440 7190 1560 7200
rect 1690 7190 1810 7200
rect 1940 7190 2060 7200
rect 2190 7190 2310 7200
rect 2440 7190 2560 7200
rect 2690 7190 2810 7200
rect 2940 7190 3060 7200
rect 3190 7190 3310 7200
rect 3440 7190 3560 7200
rect 3690 7190 3810 7200
rect 3940 7190 4060 7200
rect 4190 7190 4310 7200
rect 4440 7190 4560 7200
rect 4690 7190 4810 7200
rect 4940 7190 5060 7200
rect 5190 7190 5310 7200
rect 5440 7190 5560 7200
rect 5690 7190 5810 7200
rect 5940 7190 6060 7200
rect 6190 7190 6310 7200
rect 6440 7190 6560 7200
rect 6690 7190 6810 7200
rect 6940 7190 7060 7200
rect 7190 7190 7310 7200
rect 7440 7190 7560 7200
rect 7690 7190 7810 7200
rect 7940 7190 8000 7200
rect 0 7175 50 7190
rect 0 7075 10 7175
rect 45 7075 50 7175
rect 0 7060 50 7075
rect 200 7175 300 7190
rect 200 7075 205 7175
rect 240 7075 260 7175
rect 295 7075 300 7175
rect 200 7060 300 7075
rect 450 7175 550 7190
rect 450 7075 455 7175
rect 490 7075 510 7175
rect 545 7075 550 7175
rect 450 7060 550 7075
rect 700 7175 800 7190
rect 700 7075 705 7175
rect 740 7075 760 7175
rect 795 7075 800 7175
rect 700 7060 800 7075
rect 950 7175 1050 7190
rect 950 7075 955 7175
rect 990 7075 1010 7175
rect 1045 7075 1050 7175
rect 950 7060 1050 7075
rect 1200 7175 1300 7190
rect 1200 7075 1205 7175
rect 1240 7075 1260 7175
rect 1295 7075 1300 7175
rect 1200 7060 1300 7075
rect 1450 7175 1550 7190
rect 1450 7075 1455 7175
rect 1490 7075 1510 7175
rect 1545 7075 1550 7175
rect 1450 7060 1550 7075
rect 1700 7175 1800 7190
rect 1700 7075 1705 7175
rect 1740 7075 1760 7175
rect 1795 7075 1800 7175
rect 1700 7060 1800 7075
rect 1950 7175 2050 7190
rect 1950 7075 1955 7175
rect 1990 7075 2010 7175
rect 2045 7075 2050 7175
rect 1950 7060 2050 7075
rect 2200 7175 2300 7190
rect 2200 7075 2205 7175
rect 2240 7075 2260 7175
rect 2295 7075 2300 7175
rect 2200 7060 2300 7075
rect 2450 7175 2550 7190
rect 2450 7075 2455 7175
rect 2490 7075 2510 7175
rect 2545 7075 2550 7175
rect 2450 7060 2550 7075
rect 2700 7175 2800 7190
rect 2700 7075 2705 7175
rect 2740 7075 2760 7175
rect 2795 7075 2800 7175
rect 2700 7060 2800 7075
rect 2950 7175 3050 7190
rect 2950 7075 2955 7175
rect 2990 7075 3010 7175
rect 3045 7075 3050 7175
rect 2950 7060 3050 7075
rect 3200 7175 3300 7190
rect 3200 7075 3205 7175
rect 3240 7075 3260 7175
rect 3295 7075 3300 7175
rect 3200 7060 3300 7075
rect 3450 7175 3550 7190
rect 3450 7075 3455 7175
rect 3490 7075 3510 7175
rect 3545 7075 3550 7175
rect 3450 7060 3550 7075
rect 3700 7175 3800 7190
rect 3700 7075 3705 7175
rect 3740 7075 3760 7175
rect 3795 7075 3800 7175
rect 3700 7060 3800 7075
rect 3950 7175 4050 7190
rect 3950 7075 3955 7175
rect 3990 7075 4010 7175
rect 4045 7075 4050 7175
rect 3950 7060 4050 7075
rect 4200 7175 4300 7190
rect 4200 7075 4205 7175
rect 4240 7075 4260 7175
rect 4295 7075 4300 7175
rect 4200 7060 4300 7075
rect 4450 7175 4550 7190
rect 4450 7075 4455 7175
rect 4490 7075 4510 7175
rect 4545 7075 4550 7175
rect 4450 7060 4550 7075
rect 4700 7175 4800 7190
rect 4700 7075 4705 7175
rect 4740 7075 4760 7175
rect 4795 7075 4800 7175
rect 4700 7060 4800 7075
rect 4950 7175 5050 7190
rect 4950 7075 4955 7175
rect 4990 7075 5010 7175
rect 5045 7075 5050 7175
rect 4950 7060 5050 7075
rect 5200 7175 5300 7190
rect 5200 7075 5205 7175
rect 5240 7075 5260 7175
rect 5295 7075 5300 7175
rect 5200 7060 5300 7075
rect 5450 7175 5550 7190
rect 5450 7075 5455 7175
rect 5490 7075 5510 7175
rect 5545 7075 5550 7175
rect 5450 7060 5550 7075
rect 5700 7175 5800 7190
rect 5700 7075 5705 7175
rect 5740 7075 5760 7175
rect 5795 7075 5800 7175
rect 5700 7060 5800 7075
rect 5950 7175 6050 7190
rect 5950 7075 5955 7175
rect 5990 7075 6010 7175
rect 6045 7075 6050 7175
rect 5950 7060 6050 7075
rect 6200 7175 6300 7190
rect 6200 7075 6205 7175
rect 6240 7075 6260 7175
rect 6295 7075 6300 7175
rect 6200 7060 6300 7075
rect 6450 7175 6550 7190
rect 6450 7075 6455 7175
rect 6490 7075 6510 7175
rect 6545 7075 6550 7175
rect 6450 7060 6550 7075
rect 6700 7175 6800 7190
rect 6700 7075 6705 7175
rect 6740 7075 6760 7175
rect 6795 7075 6800 7175
rect 6700 7060 6800 7075
rect 6950 7175 7050 7190
rect 6950 7075 6955 7175
rect 6990 7075 7010 7175
rect 7045 7075 7050 7175
rect 6950 7060 7050 7075
rect 7200 7175 7300 7190
rect 7200 7075 7205 7175
rect 7240 7075 7260 7175
rect 7295 7075 7300 7175
rect 7200 7060 7300 7075
rect 7450 7175 7550 7190
rect 7450 7075 7455 7175
rect 7490 7075 7510 7175
rect 7545 7075 7550 7175
rect 7450 7060 7550 7075
rect 7700 7175 7800 7190
rect 7700 7075 7705 7175
rect 7740 7075 7760 7175
rect 7795 7075 7800 7175
rect 7700 7060 7800 7075
rect 7950 7175 8000 7190
rect 7950 7075 7955 7175
rect 7990 7075 8000 7175
rect 7950 7060 8000 7075
rect 0 7050 60 7060
rect 190 7050 310 7060
rect 440 7050 560 7060
rect 690 7050 810 7060
rect 940 7050 1060 7060
rect 1190 7050 1310 7060
rect 1440 7050 1560 7060
rect 1690 7050 1810 7060
rect 1940 7050 2060 7060
rect 2190 7050 2310 7060
rect 2440 7050 2560 7060
rect 2690 7050 2810 7060
rect 2940 7050 3060 7060
rect 3190 7050 3310 7060
rect 3440 7050 3560 7060
rect 3690 7050 3810 7060
rect 3940 7050 4060 7060
rect 4190 7050 4310 7060
rect 4440 7050 4560 7060
rect 4690 7050 4810 7060
rect 4940 7050 5060 7060
rect 5190 7050 5310 7060
rect 5440 7050 5560 7060
rect 5690 7050 5810 7060
rect 5940 7050 6060 7060
rect 6190 7050 6310 7060
rect 6440 7050 6560 7060
rect 6690 7050 6810 7060
rect 6940 7050 7060 7060
rect 7190 7050 7310 7060
rect 7440 7050 7560 7060
rect 7690 7050 7810 7060
rect 7940 7050 8000 7060
rect 0 7045 450 7050
rect 0 7010 75 7045
rect 175 7010 325 7045
rect 425 7010 450 7045
rect 0 6990 450 7010
rect 0 6955 75 6990
rect 175 6955 325 6990
rect 425 6955 450 6990
rect 0 6950 450 6955
rect 550 7045 1450 7050
rect 550 7010 575 7045
rect 675 7010 825 7045
rect 925 7010 1075 7045
rect 1175 7010 1325 7045
rect 1425 7010 1450 7045
rect 550 6990 1450 7010
rect 550 6955 575 6990
rect 675 6955 825 6990
rect 925 6955 1075 6990
rect 1175 6955 1325 6990
rect 1425 6955 1450 6990
rect 550 6950 1450 6955
rect 1550 7045 2450 7050
rect 1550 7010 1575 7045
rect 1675 7010 1825 7045
rect 1925 7010 2075 7045
rect 2175 7010 2325 7045
rect 2425 7010 2450 7045
rect 1550 6990 2450 7010
rect 1550 6955 1575 6990
rect 1675 6955 1825 6990
rect 1925 6955 2075 6990
rect 2175 6955 2325 6990
rect 2425 6955 2450 6990
rect 1550 6950 2450 6955
rect 2550 7045 3450 7050
rect 2550 7010 2575 7045
rect 2675 7010 2825 7045
rect 2925 7010 3075 7045
rect 3175 7010 3325 7045
rect 3425 7010 3450 7045
rect 2550 6990 3450 7010
rect 2550 6955 2575 6990
rect 2675 6955 2825 6990
rect 2925 6955 3075 6990
rect 3175 6955 3325 6990
rect 3425 6955 3450 6990
rect 2550 6950 3450 6955
rect 3550 7045 4450 7050
rect 3550 7010 3575 7045
rect 3675 7010 3825 7045
rect 3925 7010 4075 7045
rect 4175 7010 4325 7045
rect 4425 7010 4450 7045
rect 3550 6990 4450 7010
rect 3550 6955 3575 6990
rect 3675 6955 3825 6990
rect 3925 6955 4075 6990
rect 4175 6955 4325 6990
rect 4425 6955 4450 6990
rect 3550 6950 4450 6955
rect 4550 7045 5450 7050
rect 4550 7010 4575 7045
rect 4675 7010 4825 7045
rect 4925 7010 5075 7045
rect 5175 7010 5325 7045
rect 5425 7010 5450 7045
rect 4550 6990 5450 7010
rect 4550 6955 4575 6990
rect 4675 6955 4825 6990
rect 4925 6955 5075 6990
rect 5175 6955 5325 6990
rect 5425 6955 5450 6990
rect 4550 6950 5450 6955
rect 5550 7045 6450 7050
rect 5550 7010 5575 7045
rect 5675 7010 5825 7045
rect 5925 7010 6075 7045
rect 6175 7010 6325 7045
rect 6425 7010 6450 7045
rect 5550 6990 6450 7010
rect 5550 6955 5575 6990
rect 5675 6955 5825 6990
rect 5925 6955 6075 6990
rect 6175 6955 6325 6990
rect 6425 6955 6450 6990
rect 5550 6950 6450 6955
rect 6550 7045 7450 7050
rect 6550 7010 6575 7045
rect 6675 7010 6825 7045
rect 6925 7010 7075 7045
rect 7175 7010 7325 7045
rect 7425 7010 7450 7045
rect 6550 6990 7450 7010
rect 6550 6955 6575 6990
rect 6675 6955 6825 6990
rect 6925 6955 7075 6990
rect 7175 6955 7325 6990
rect 7425 6955 7450 6990
rect 6550 6950 7450 6955
rect 7550 7045 8000 7050
rect 7550 7010 7575 7045
rect 7675 7010 7825 7045
rect 7925 7010 8000 7045
rect 7550 6990 8000 7010
rect 7550 6955 7575 6990
rect 7675 6955 7825 6990
rect 7925 6955 8000 6990
rect 7550 6950 8000 6955
rect 0 6940 60 6950
rect 190 6940 310 6950
rect 440 6940 560 6950
rect 690 6940 810 6950
rect 940 6940 1060 6950
rect 1190 6940 1310 6950
rect 1440 6940 1560 6950
rect 1690 6940 1810 6950
rect 1940 6940 2060 6950
rect 2190 6940 2310 6950
rect 2440 6940 2560 6950
rect 2690 6940 2810 6950
rect 2940 6940 3060 6950
rect 3190 6940 3310 6950
rect 3440 6940 3560 6950
rect 3690 6940 3810 6950
rect 3940 6940 4060 6950
rect 4190 6940 4310 6950
rect 4440 6940 4560 6950
rect 4690 6940 4810 6950
rect 4940 6940 5060 6950
rect 5190 6940 5310 6950
rect 5440 6940 5560 6950
rect 5690 6940 5810 6950
rect 5940 6940 6060 6950
rect 6190 6940 6310 6950
rect 6440 6940 6560 6950
rect 6690 6940 6810 6950
rect 6940 6940 7060 6950
rect 7190 6940 7310 6950
rect 7440 6940 7560 6950
rect 7690 6940 7810 6950
rect 7940 6940 8000 6950
rect 0 6925 50 6940
rect 0 6825 10 6925
rect 45 6825 50 6925
rect 0 6810 50 6825
rect 200 6925 300 6940
rect 200 6825 205 6925
rect 240 6825 260 6925
rect 295 6825 300 6925
rect 200 6810 300 6825
rect 450 6925 550 6940
rect 450 6825 455 6925
rect 490 6825 510 6925
rect 545 6825 550 6925
rect 450 6810 550 6825
rect 700 6925 800 6940
rect 700 6825 705 6925
rect 740 6825 760 6925
rect 795 6825 800 6925
rect 700 6810 800 6825
rect 950 6925 1050 6940
rect 950 6825 955 6925
rect 990 6825 1010 6925
rect 1045 6825 1050 6925
rect 950 6810 1050 6825
rect 1200 6925 1300 6940
rect 1200 6825 1205 6925
rect 1240 6825 1260 6925
rect 1295 6825 1300 6925
rect 1200 6810 1300 6825
rect 1450 6925 1550 6940
rect 1450 6825 1455 6925
rect 1490 6825 1510 6925
rect 1545 6825 1550 6925
rect 1450 6810 1550 6825
rect 1700 6925 1800 6940
rect 1700 6825 1705 6925
rect 1740 6825 1760 6925
rect 1795 6825 1800 6925
rect 1700 6810 1800 6825
rect 1950 6925 2050 6940
rect 1950 6825 1955 6925
rect 1990 6825 2010 6925
rect 2045 6825 2050 6925
rect 1950 6810 2050 6825
rect 2200 6925 2300 6940
rect 2200 6825 2205 6925
rect 2240 6825 2260 6925
rect 2295 6825 2300 6925
rect 2200 6810 2300 6825
rect 2450 6925 2550 6940
rect 2450 6825 2455 6925
rect 2490 6825 2510 6925
rect 2545 6825 2550 6925
rect 2450 6810 2550 6825
rect 2700 6925 2800 6940
rect 2700 6825 2705 6925
rect 2740 6825 2760 6925
rect 2795 6825 2800 6925
rect 2700 6810 2800 6825
rect 2950 6925 3050 6940
rect 2950 6825 2955 6925
rect 2990 6825 3010 6925
rect 3045 6825 3050 6925
rect 2950 6810 3050 6825
rect 3200 6925 3300 6940
rect 3200 6825 3205 6925
rect 3240 6825 3260 6925
rect 3295 6825 3300 6925
rect 3200 6810 3300 6825
rect 3450 6925 3550 6940
rect 3450 6825 3455 6925
rect 3490 6825 3510 6925
rect 3545 6825 3550 6925
rect 3450 6810 3550 6825
rect 3700 6925 3800 6940
rect 3700 6825 3705 6925
rect 3740 6825 3760 6925
rect 3795 6825 3800 6925
rect 3700 6810 3800 6825
rect 3950 6925 4050 6940
rect 3950 6825 3955 6925
rect 3990 6825 4010 6925
rect 4045 6825 4050 6925
rect 3950 6810 4050 6825
rect 4200 6925 4300 6940
rect 4200 6825 4205 6925
rect 4240 6825 4260 6925
rect 4295 6825 4300 6925
rect 4200 6810 4300 6825
rect 4450 6925 4550 6940
rect 4450 6825 4455 6925
rect 4490 6825 4510 6925
rect 4545 6825 4550 6925
rect 4450 6810 4550 6825
rect 4700 6925 4800 6940
rect 4700 6825 4705 6925
rect 4740 6825 4760 6925
rect 4795 6825 4800 6925
rect 4700 6810 4800 6825
rect 4950 6925 5050 6940
rect 4950 6825 4955 6925
rect 4990 6825 5010 6925
rect 5045 6825 5050 6925
rect 4950 6810 5050 6825
rect 5200 6925 5300 6940
rect 5200 6825 5205 6925
rect 5240 6825 5260 6925
rect 5295 6825 5300 6925
rect 5200 6810 5300 6825
rect 5450 6925 5550 6940
rect 5450 6825 5455 6925
rect 5490 6825 5510 6925
rect 5545 6825 5550 6925
rect 5450 6810 5550 6825
rect 5700 6925 5800 6940
rect 5700 6825 5705 6925
rect 5740 6825 5760 6925
rect 5795 6825 5800 6925
rect 5700 6810 5800 6825
rect 5950 6925 6050 6940
rect 5950 6825 5955 6925
rect 5990 6825 6010 6925
rect 6045 6825 6050 6925
rect 5950 6810 6050 6825
rect 6200 6925 6300 6940
rect 6200 6825 6205 6925
rect 6240 6825 6260 6925
rect 6295 6825 6300 6925
rect 6200 6810 6300 6825
rect 6450 6925 6550 6940
rect 6450 6825 6455 6925
rect 6490 6825 6510 6925
rect 6545 6825 6550 6925
rect 6450 6810 6550 6825
rect 6700 6925 6800 6940
rect 6700 6825 6705 6925
rect 6740 6825 6760 6925
rect 6795 6825 6800 6925
rect 6700 6810 6800 6825
rect 6950 6925 7050 6940
rect 6950 6825 6955 6925
rect 6990 6825 7010 6925
rect 7045 6825 7050 6925
rect 6950 6810 7050 6825
rect 7200 6925 7300 6940
rect 7200 6825 7205 6925
rect 7240 6825 7260 6925
rect 7295 6825 7300 6925
rect 7200 6810 7300 6825
rect 7450 6925 7550 6940
rect 7450 6825 7455 6925
rect 7490 6825 7510 6925
rect 7545 6825 7550 6925
rect 7450 6810 7550 6825
rect 7700 6925 7800 6940
rect 7700 6825 7705 6925
rect 7740 6825 7760 6925
rect 7795 6825 7800 6925
rect 7700 6810 7800 6825
rect 7950 6925 8000 6940
rect 7950 6825 7955 6925
rect 7990 6825 8000 6925
rect 7950 6810 8000 6825
rect 0 6800 60 6810
rect 190 6800 310 6810
rect 440 6800 560 6810
rect 690 6800 810 6810
rect 940 6800 1060 6810
rect 1190 6800 1310 6810
rect 1440 6800 1560 6810
rect 1690 6800 1810 6810
rect 1940 6800 2060 6810
rect 2190 6800 2310 6810
rect 2440 6800 2560 6810
rect 2690 6800 2810 6810
rect 2940 6800 3060 6810
rect 3190 6800 3310 6810
rect 3440 6800 3560 6810
rect 3690 6800 3810 6810
rect 3940 6800 4060 6810
rect 4190 6800 4310 6810
rect 4440 6800 4560 6810
rect 4690 6800 4810 6810
rect 4940 6800 5060 6810
rect 5190 6800 5310 6810
rect 5440 6800 5560 6810
rect 5690 6800 5810 6810
rect 5940 6800 6060 6810
rect 6190 6800 6310 6810
rect 6440 6800 6560 6810
rect 6690 6800 6810 6810
rect 6940 6800 7060 6810
rect 7190 6800 7310 6810
rect 7440 6800 7560 6810
rect 7690 6800 7810 6810
rect 7940 6800 8000 6810
rect 0 6795 200 6800
rect 0 6760 75 6795
rect 175 6760 200 6795
rect 0 6740 200 6760
rect 0 6705 75 6740
rect 175 6705 200 6740
rect 0 6700 200 6705
rect 300 6795 450 6800
rect 300 6760 325 6795
rect 425 6760 450 6795
rect 300 6740 450 6760
rect 300 6705 325 6740
rect 425 6705 450 6740
rect 300 6700 450 6705
rect 550 6795 700 6800
rect 550 6760 575 6795
rect 675 6760 700 6795
rect 550 6740 700 6760
rect 550 6705 575 6740
rect 675 6705 700 6740
rect 550 6700 700 6705
rect 800 6795 1200 6800
rect 800 6760 825 6795
rect 925 6760 1075 6795
rect 1175 6760 1200 6795
rect 800 6740 1200 6760
rect 800 6705 825 6740
rect 925 6705 1075 6740
rect 1175 6705 1200 6740
rect 800 6700 1200 6705
rect 1300 6795 1450 6800
rect 1300 6760 1325 6795
rect 1425 6760 1450 6795
rect 1300 6740 1450 6760
rect 1300 6705 1325 6740
rect 1425 6705 1450 6740
rect 1300 6700 1450 6705
rect 1550 6795 1700 6800
rect 1550 6760 1575 6795
rect 1675 6760 1700 6795
rect 1550 6740 1700 6760
rect 1550 6705 1575 6740
rect 1675 6705 1700 6740
rect 1550 6700 1700 6705
rect 1800 6795 2200 6800
rect 1800 6760 1825 6795
rect 1925 6760 2075 6795
rect 2175 6760 2200 6795
rect 1800 6740 2200 6760
rect 1800 6705 1825 6740
rect 1925 6705 2075 6740
rect 2175 6705 2200 6740
rect 1800 6700 2200 6705
rect 2300 6795 2450 6800
rect 2300 6760 2325 6795
rect 2425 6760 2450 6795
rect 2300 6740 2450 6760
rect 2300 6705 2325 6740
rect 2425 6705 2450 6740
rect 2300 6700 2450 6705
rect 2550 6795 2700 6800
rect 2550 6760 2575 6795
rect 2675 6760 2700 6795
rect 2550 6740 2700 6760
rect 2550 6705 2575 6740
rect 2675 6705 2700 6740
rect 2550 6700 2700 6705
rect 2800 6795 3200 6800
rect 2800 6760 2825 6795
rect 2925 6760 3075 6795
rect 3175 6760 3200 6795
rect 2800 6740 3200 6760
rect 2800 6705 2825 6740
rect 2925 6705 3075 6740
rect 3175 6705 3200 6740
rect 2800 6700 3200 6705
rect 3300 6795 3450 6800
rect 3300 6760 3325 6795
rect 3425 6760 3450 6795
rect 3300 6740 3450 6760
rect 3300 6705 3325 6740
rect 3425 6705 3450 6740
rect 3300 6700 3450 6705
rect 3550 6795 3700 6800
rect 3550 6760 3575 6795
rect 3675 6760 3700 6795
rect 3550 6740 3700 6760
rect 3550 6705 3575 6740
rect 3675 6705 3700 6740
rect 3550 6700 3700 6705
rect 3800 6795 4200 6800
rect 3800 6760 3825 6795
rect 3925 6760 4075 6795
rect 4175 6760 4200 6795
rect 3800 6740 4200 6760
rect 3800 6705 3825 6740
rect 3925 6705 4075 6740
rect 4175 6705 4200 6740
rect 3800 6700 4200 6705
rect 4300 6795 4450 6800
rect 4300 6760 4325 6795
rect 4425 6760 4450 6795
rect 4300 6740 4450 6760
rect 4300 6705 4325 6740
rect 4425 6705 4450 6740
rect 4300 6700 4450 6705
rect 4550 6795 4700 6800
rect 4550 6760 4575 6795
rect 4675 6760 4700 6795
rect 4550 6740 4700 6760
rect 4550 6705 4575 6740
rect 4675 6705 4700 6740
rect 4550 6700 4700 6705
rect 4800 6795 5200 6800
rect 4800 6760 4825 6795
rect 4925 6760 5075 6795
rect 5175 6760 5200 6795
rect 4800 6740 5200 6760
rect 4800 6705 4825 6740
rect 4925 6705 5075 6740
rect 5175 6705 5200 6740
rect 4800 6700 5200 6705
rect 5300 6795 5450 6800
rect 5300 6760 5325 6795
rect 5425 6760 5450 6795
rect 5300 6740 5450 6760
rect 5300 6705 5325 6740
rect 5425 6705 5450 6740
rect 5300 6700 5450 6705
rect 5550 6795 5700 6800
rect 5550 6760 5575 6795
rect 5675 6760 5700 6795
rect 5550 6740 5700 6760
rect 5550 6705 5575 6740
rect 5675 6705 5700 6740
rect 5550 6700 5700 6705
rect 5800 6795 6200 6800
rect 5800 6760 5825 6795
rect 5925 6760 6075 6795
rect 6175 6760 6200 6795
rect 5800 6740 6200 6760
rect 5800 6705 5825 6740
rect 5925 6705 6075 6740
rect 6175 6705 6200 6740
rect 5800 6700 6200 6705
rect 6300 6795 6450 6800
rect 6300 6760 6325 6795
rect 6425 6760 6450 6795
rect 6300 6740 6450 6760
rect 6300 6705 6325 6740
rect 6425 6705 6450 6740
rect 6300 6700 6450 6705
rect 6550 6795 6700 6800
rect 6550 6760 6575 6795
rect 6675 6760 6700 6795
rect 6550 6740 6700 6760
rect 6550 6705 6575 6740
rect 6675 6705 6700 6740
rect 6550 6700 6700 6705
rect 6800 6795 7200 6800
rect 6800 6760 6825 6795
rect 6925 6760 7075 6795
rect 7175 6760 7200 6795
rect 6800 6740 7200 6760
rect 6800 6705 6825 6740
rect 6925 6705 7075 6740
rect 7175 6705 7200 6740
rect 6800 6700 7200 6705
rect 7300 6795 7450 6800
rect 7300 6760 7325 6795
rect 7425 6760 7450 6795
rect 7300 6740 7450 6760
rect 7300 6705 7325 6740
rect 7425 6705 7450 6740
rect 7300 6700 7450 6705
rect 7550 6795 7700 6800
rect 7550 6760 7575 6795
rect 7675 6760 7700 6795
rect 7550 6740 7700 6760
rect 7550 6705 7575 6740
rect 7675 6705 7700 6740
rect 7550 6700 7700 6705
rect 7800 6795 8000 6800
rect 7800 6760 7825 6795
rect 7925 6760 8000 6795
rect 7800 6740 8000 6760
rect 7800 6705 7825 6740
rect 7925 6705 8000 6740
rect 7800 6700 8000 6705
rect 0 6690 60 6700
rect 190 6690 310 6700
rect 440 6690 560 6700
rect 690 6690 810 6700
rect 940 6690 1060 6700
rect 1190 6690 1310 6700
rect 1440 6690 1560 6700
rect 1690 6690 1810 6700
rect 1940 6690 2060 6700
rect 2190 6690 2310 6700
rect 2440 6690 2560 6700
rect 2690 6690 2810 6700
rect 2940 6690 3060 6700
rect 3190 6690 3310 6700
rect 3440 6690 3560 6700
rect 3690 6690 3810 6700
rect 3940 6690 4060 6700
rect 4190 6690 4310 6700
rect 4440 6690 4560 6700
rect 4690 6690 4810 6700
rect 4940 6690 5060 6700
rect 5190 6690 5310 6700
rect 5440 6690 5560 6700
rect 5690 6690 5810 6700
rect 5940 6690 6060 6700
rect 6190 6690 6310 6700
rect 6440 6690 6560 6700
rect 6690 6690 6810 6700
rect 6940 6690 7060 6700
rect 7190 6690 7310 6700
rect 7440 6690 7560 6700
rect 7690 6690 7810 6700
rect 7940 6690 8000 6700
rect 0 6675 50 6690
rect 0 6575 10 6675
rect 45 6575 50 6675
rect 0 6560 50 6575
rect 200 6675 300 6690
rect 200 6575 205 6675
rect 240 6575 260 6675
rect 295 6575 300 6675
rect 200 6560 300 6575
rect 450 6675 550 6690
rect 450 6575 455 6675
rect 490 6575 510 6675
rect 545 6575 550 6675
rect 450 6560 550 6575
rect 700 6675 800 6690
rect 700 6575 705 6675
rect 740 6575 760 6675
rect 795 6575 800 6675
rect 700 6560 800 6575
rect 950 6675 1050 6690
rect 950 6575 955 6675
rect 990 6575 1010 6675
rect 1045 6575 1050 6675
rect 950 6560 1050 6575
rect 1200 6675 1300 6690
rect 1200 6575 1205 6675
rect 1240 6575 1260 6675
rect 1295 6575 1300 6675
rect 1200 6560 1300 6575
rect 1450 6675 1550 6690
rect 1450 6575 1455 6675
rect 1490 6575 1510 6675
rect 1545 6575 1550 6675
rect 1450 6560 1550 6575
rect 1700 6675 1800 6690
rect 1700 6575 1705 6675
rect 1740 6575 1760 6675
rect 1795 6575 1800 6675
rect 1700 6560 1800 6575
rect 1950 6675 2050 6690
rect 1950 6575 1955 6675
rect 1990 6575 2010 6675
rect 2045 6575 2050 6675
rect 1950 6560 2050 6575
rect 2200 6675 2300 6690
rect 2200 6575 2205 6675
rect 2240 6575 2260 6675
rect 2295 6575 2300 6675
rect 2200 6560 2300 6575
rect 2450 6675 2550 6690
rect 2450 6575 2455 6675
rect 2490 6575 2510 6675
rect 2545 6575 2550 6675
rect 2450 6560 2550 6575
rect 2700 6675 2800 6690
rect 2700 6575 2705 6675
rect 2740 6575 2760 6675
rect 2795 6575 2800 6675
rect 2700 6560 2800 6575
rect 2950 6675 3050 6690
rect 2950 6575 2955 6675
rect 2990 6575 3010 6675
rect 3045 6575 3050 6675
rect 2950 6560 3050 6575
rect 3200 6675 3300 6690
rect 3200 6575 3205 6675
rect 3240 6575 3260 6675
rect 3295 6575 3300 6675
rect 3200 6560 3300 6575
rect 3450 6675 3550 6690
rect 3450 6575 3455 6675
rect 3490 6575 3510 6675
rect 3545 6575 3550 6675
rect 3450 6560 3550 6575
rect 3700 6675 3800 6690
rect 3700 6575 3705 6675
rect 3740 6575 3760 6675
rect 3795 6575 3800 6675
rect 3700 6560 3800 6575
rect 3950 6675 4050 6690
rect 3950 6575 3955 6675
rect 3990 6575 4010 6675
rect 4045 6575 4050 6675
rect 3950 6560 4050 6575
rect 4200 6675 4300 6690
rect 4200 6575 4205 6675
rect 4240 6575 4260 6675
rect 4295 6575 4300 6675
rect 4200 6560 4300 6575
rect 4450 6675 4550 6690
rect 4450 6575 4455 6675
rect 4490 6575 4510 6675
rect 4545 6575 4550 6675
rect 4450 6560 4550 6575
rect 4700 6675 4800 6690
rect 4700 6575 4705 6675
rect 4740 6575 4760 6675
rect 4795 6575 4800 6675
rect 4700 6560 4800 6575
rect 4950 6675 5050 6690
rect 4950 6575 4955 6675
rect 4990 6575 5010 6675
rect 5045 6575 5050 6675
rect 4950 6560 5050 6575
rect 5200 6675 5300 6690
rect 5200 6575 5205 6675
rect 5240 6575 5260 6675
rect 5295 6575 5300 6675
rect 5200 6560 5300 6575
rect 5450 6675 5550 6690
rect 5450 6575 5455 6675
rect 5490 6575 5510 6675
rect 5545 6575 5550 6675
rect 5450 6560 5550 6575
rect 5700 6675 5800 6690
rect 5700 6575 5705 6675
rect 5740 6575 5760 6675
rect 5795 6575 5800 6675
rect 5700 6560 5800 6575
rect 5950 6675 6050 6690
rect 5950 6575 5955 6675
rect 5990 6575 6010 6675
rect 6045 6575 6050 6675
rect 5950 6560 6050 6575
rect 6200 6675 6300 6690
rect 6200 6575 6205 6675
rect 6240 6575 6260 6675
rect 6295 6575 6300 6675
rect 6200 6560 6300 6575
rect 6450 6675 6550 6690
rect 6450 6575 6455 6675
rect 6490 6575 6510 6675
rect 6545 6575 6550 6675
rect 6450 6560 6550 6575
rect 6700 6675 6800 6690
rect 6700 6575 6705 6675
rect 6740 6575 6760 6675
rect 6795 6575 6800 6675
rect 6700 6560 6800 6575
rect 6950 6675 7050 6690
rect 6950 6575 6955 6675
rect 6990 6575 7010 6675
rect 7045 6575 7050 6675
rect 6950 6560 7050 6575
rect 7200 6675 7300 6690
rect 7200 6575 7205 6675
rect 7240 6575 7260 6675
rect 7295 6575 7300 6675
rect 7200 6560 7300 6575
rect 7450 6675 7550 6690
rect 7450 6575 7455 6675
rect 7490 6575 7510 6675
rect 7545 6575 7550 6675
rect 7450 6560 7550 6575
rect 7700 6675 7800 6690
rect 7700 6575 7705 6675
rect 7740 6575 7760 6675
rect 7795 6575 7800 6675
rect 7700 6560 7800 6575
rect 7950 6675 8000 6690
rect 7950 6575 7955 6675
rect 7990 6575 8000 6675
rect 7950 6560 8000 6575
rect 0 6550 60 6560
rect 190 6550 310 6560
rect 440 6550 560 6560
rect 690 6550 810 6560
rect 940 6550 1060 6560
rect 1190 6550 1310 6560
rect 1440 6550 1560 6560
rect 1690 6550 1810 6560
rect 1940 6550 2060 6560
rect 2190 6550 2310 6560
rect 2440 6550 2560 6560
rect 2690 6550 2810 6560
rect 2940 6550 3060 6560
rect 3190 6550 3310 6560
rect 3440 6550 3560 6560
rect 3690 6550 3810 6560
rect 3940 6550 4060 6560
rect 4190 6550 4310 6560
rect 4440 6550 4560 6560
rect 4690 6550 4810 6560
rect 4940 6550 5060 6560
rect 5190 6550 5310 6560
rect 5440 6550 5560 6560
rect 5690 6550 5810 6560
rect 5940 6550 6060 6560
rect 6190 6550 6310 6560
rect 6440 6550 6560 6560
rect 6690 6550 6810 6560
rect 6940 6550 7060 6560
rect 7190 6550 7310 6560
rect 7440 6550 7560 6560
rect 7690 6550 7810 6560
rect 7940 6550 8000 6560
rect 0 6545 200 6550
rect 0 6510 75 6545
rect 175 6510 200 6545
rect 0 6490 200 6510
rect 0 6455 75 6490
rect 175 6455 200 6490
rect 0 6450 200 6455
rect 300 6545 450 6550
rect 300 6510 325 6545
rect 425 6510 450 6545
rect 300 6490 450 6510
rect 300 6455 325 6490
rect 425 6455 450 6490
rect 300 6450 450 6455
rect 550 6545 700 6550
rect 550 6510 575 6545
rect 675 6510 700 6545
rect 550 6490 700 6510
rect 550 6455 575 6490
rect 675 6455 700 6490
rect 550 6450 700 6455
rect 800 6545 950 6550
rect 800 6510 825 6545
rect 925 6510 950 6545
rect 800 6490 950 6510
rect 800 6455 825 6490
rect 925 6455 950 6490
rect 800 6450 950 6455
rect 1050 6545 1200 6550
rect 1050 6510 1075 6545
rect 1175 6510 1200 6545
rect 1050 6490 1200 6510
rect 1050 6455 1075 6490
rect 1175 6455 1200 6490
rect 1050 6450 1200 6455
rect 1300 6545 1450 6550
rect 1300 6510 1325 6545
rect 1425 6510 1450 6545
rect 1300 6490 1450 6510
rect 1300 6455 1325 6490
rect 1425 6455 1450 6490
rect 1300 6450 1450 6455
rect 1550 6545 1700 6550
rect 1550 6510 1575 6545
rect 1675 6510 1700 6545
rect 1550 6490 1700 6510
rect 1550 6455 1575 6490
rect 1675 6455 1700 6490
rect 1550 6450 1700 6455
rect 1800 6545 2200 6550
rect 1800 6510 1825 6545
rect 1925 6510 2075 6545
rect 2175 6510 2200 6545
rect 1800 6490 2200 6510
rect 1800 6455 1825 6490
rect 1925 6455 2075 6490
rect 2175 6455 2200 6490
rect 1800 6450 2200 6455
rect 2300 6545 2450 6550
rect 2300 6510 2325 6545
rect 2425 6510 2450 6545
rect 2300 6490 2450 6510
rect 2300 6455 2325 6490
rect 2425 6455 2450 6490
rect 2300 6450 2450 6455
rect 2550 6545 2700 6550
rect 2550 6510 2575 6545
rect 2675 6510 2700 6545
rect 2550 6490 2700 6510
rect 2550 6455 2575 6490
rect 2675 6455 2700 6490
rect 2550 6450 2700 6455
rect 2800 6545 2950 6550
rect 2800 6510 2825 6545
rect 2925 6510 2950 6545
rect 2800 6490 2950 6510
rect 2800 6455 2825 6490
rect 2925 6455 2950 6490
rect 2800 6450 2950 6455
rect 3050 6545 3200 6550
rect 3050 6510 3075 6545
rect 3175 6510 3200 6545
rect 3050 6490 3200 6510
rect 3050 6455 3075 6490
rect 3175 6455 3200 6490
rect 3050 6450 3200 6455
rect 3300 6545 3450 6550
rect 3300 6510 3325 6545
rect 3425 6510 3450 6545
rect 3300 6490 3450 6510
rect 3300 6455 3325 6490
rect 3425 6455 3450 6490
rect 3300 6450 3450 6455
rect 3550 6545 3700 6550
rect 3550 6510 3575 6545
rect 3675 6510 3700 6545
rect 3550 6490 3700 6510
rect 3550 6455 3575 6490
rect 3675 6455 3700 6490
rect 3550 6450 3700 6455
rect 3800 6545 4200 6550
rect 3800 6510 3825 6545
rect 3925 6510 4075 6545
rect 4175 6510 4200 6545
rect 3800 6490 4200 6510
rect 3800 6455 3825 6490
rect 3925 6455 4075 6490
rect 4175 6455 4200 6490
rect 3800 6450 4200 6455
rect 4300 6545 4450 6550
rect 4300 6510 4325 6545
rect 4425 6510 4450 6545
rect 4300 6490 4450 6510
rect 4300 6455 4325 6490
rect 4425 6455 4450 6490
rect 4300 6450 4450 6455
rect 4550 6545 4700 6550
rect 4550 6510 4575 6545
rect 4675 6510 4700 6545
rect 4550 6490 4700 6510
rect 4550 6455 4575 6490
rect 4675 6455 4700 6490
rect 4550 6450 4700 6455
rect 4800 6545 4950 6550
rect 4800 6510 4825 6545
rect 4925 6510 4950 6545
rect 4800 6490 4950 6510
rect 4800 6455 4825 6490
rect 4925 6455 4950 6490
rect 4800 6450 4950 6455
rect 5050 6545 5200 6550
rect 5050 6510 5075 6545
rect 5175 6510 5200 6545
rect 5050 6490 5200 6510
rect 5050 6455 5075 6490
rect 5175 6455 5200 6490
rect 5050 6450 5200 6455
rect 5300 6545 5450 6550
rect 5300 6510 5325 6545
rect 5425 6510 5450 6545
rect 5300 6490 5450 6510
rect 5300 6455 5325 6490
rect 5425 6455 5450 6490
rect 5300 6450 5450 6455
rect 5550 6545 5700 6550
rect 5550 6510 5575 6545
rect 5675 6510 5700 6545
rect 5550 6490 5700 6510
rect 5550 6455 5575 6490
rect 5675 6455 5700 6490
rect 5550 6450 5700 6455
rect 5800 6545 6200 6550
rect 5800 6510 5825 6545
rect 5925 6510 6075 6545
rect 6175 6510 6200 6545
rect 5800 6490 6200 6510
rect 5800 6455 5825 6490
rect 5925 6455 6075 6490
rect 6175 6455 6200 6490
rect 5800 6450 6200 6455
rect 6300 6545 6450 6550
rect 6300 6510 6325 6545
rect 6425 6510 6450 6545
rect 6300 6490 6450 6510
rect 6300 6455 6325 6490
rect 6425 6455 6450 6490
rect 6300 6450 6450 6455
rect 6550 6545 6700 6550
rect 6550 6510 6575 6545
rect 6675 6510 6700 6545
rect 6550 6490 6700 6510
rect 6550 6455 6575 6490
rect 6675 6455 6700 6490
rect 6550 6450 6700 6455
rect 6800 6545 6950 6550
rect 6800 6510 6825 6545
rect 6925 6510 6950 6545
rect 6800 6490 6950 6510
rect 6800 6455 6825 6490
rect 6925 6455 6950 6490
rect 6800 6450 6950 6455
rect 7050 6545 7200 6550
rect 7050 6510 7075 6545
rect 7175 6510 7200 6545
rect 7050 6490 7200 6510
rect 7050 6455 7075 6490
rect 7175 6455 7200 6490
rect 7050 6450 7200 6455
rect 7300 6545 7450 6550
rect 7300 6510 7325 6545
rect 7425 6510 7450 6545
rect 7300 6490 7450 6510
rect 7300 6455 7325 6490
rect 7425 6455 7450 6490
rect 7300 6450 7450 6455
rect 7550 6545 7700 6550
rect 7550 6510 7575 6545
rect 7675 6510 7700 6545
rect 7550 6490 7700 6510
rect 7550 6455 7575 6490
rect 7675 6455 7700 6490
rect 7550 6450 7700 6455
rect 7800 6545 8000 6550
rect 7800 6510 7825 6545
rect 7925 6510 8000 6545
rect 7800 6490 8000 6510
rect 7800 6455 7825 6490
rect 7925 6455 8000 6490
rect 7800 6450 8000 6455
rect 0 6440 60 6450
rect 190 6440 310 6450
rect 440 6440 560 6450
rect 690 6440 810 6450
rect 940 6440 1060 6450
rect 1190 6440 1310 6450
rect 1440 6440 1560 6450
rect 1690 6440 1810 6450
rect 1940 6440 2060 6450
rect 2190 6440 2310 6450
rect 2440 6440 2560 6450
rect 2690 6440 2810 6450
rect 2940 6440 3060 6450
rect 3190 6440 3310 6450
rect 3440 6440 3560 6450
rect 3690 6440 3810 6450
rect 3940 6440 4060 6450
rect 4190 6440 4310 6450
rect 4440 6440 4560 6450
rect 4690 6440 4810 6450
rect 4940 6440 5060 6450
rect 5190 6440 5310 6450
rect 5440 6440 5560 6450
rect 5690 6440 5810 6450
rect 5940 6440 6060 6450
rect 6190 6440 6310 6450
rect 6440 6440 6560 6450
rect 6690 6440 6810 6450
rect 6940 6440 7060 6450
rect 7190 6440 7310 6450
rect 7440 6440 7560 6450
rect 7690 6440 7810 6450
rect 7940 6440 8000 6450
rect 0 6425 50 6440
rect 0 6325 10 6425
rect 45 6325 50 6425
rect 0 6310 50 6325
rect 200 6425 300 6440
rect 200 6325 205 6425
rect 240 6325 260 6425
rect 295 6325 300 6425
rect 200 6310 300 6325
rect 450 6425 550 6440
rect 450 6325 455 6425
rect 490 6325 510 6425
rect 545 6325 550 6425
rect 450 6310 550 6325
rect 700 6425 800 6440
rect 700 6325 705 6425
rect 740 6325 760 6425
rect 795 6325 800 6425
rect 700 6310 800 6325
rect 950 6425 1050 6440
rect 950 6325 955 6425
rect 990 6325 1010 6425
rect 1045 6325 1050 6425
rect 950 6310 1050 6325
rect 1200 6425 1300 6440
rect 1200 6325 1205 6425
rect 1240 6325 1260 6425
rect 1295 6325 1300 6425
rect 1200 6310 1300 6325
rect 1450 6425 1550 6440
rect 1450 6325 1455 6425
rect 1490 6325 1510 6425
rect 1545 6325 1550 6425
rect 1450 6310 1550 6325
rect 1700 6425 1800 6440
rect 1700 6325 1705 6425
rect 1740 6325 1760 6425
rect 1795 6325 1800 6425
rect 1700 6310 1800 6325
rect 1950 6425 2050 6440
rect 1950 6325 1955 6425
rect 1990 6325 2010 6425
rect 2045 6325 2050 6425
rect 1950 6310 2050 6325
rect 2200 6425 2300 6440
rect 2200 6325 2205 6425
rect 2240 6325 2260 6425
rect 2295 6325 2300 6425
rect 2200 6310 2300 6325
rect 2450 6425 2550 6440
rect 2450 6325 2455 6425
rect 2490 6325 2510 6425
rect 2545 6325 2550 6425
rect 2450 6310 2550 6325
rect 2700 6425 2800 6440
rect 2700 6325 2705 6425
rect 2740 6325 2760 6425
rect 2795 6325 2800 6425
rect 2700 6310 2800 6325
rect 2950 6425 3050 6440
rect 2950 6325 2955 6425
rect 2990 6325 3010 6425
rect 3045 6325 3050 6425
rect 2950 6310 3050 6325
rect 3200 6425 3300 6440
rect 3200 6325 3205 6425
rect 3240 6325 3260 6425
rect 3295 6325 3300 6425
rect 3200 6310 3300 6325
rect 3450 6425 3550 6440
rect 3450 6325 3455 6425
rect 3490 6325 3510 6425
rect 3545 6325 3550 6425
rect 3450 6310 3550 6325
rect 3700 6425 3800 6440
rect 3700 6325 3705 6425
rect 3740 6325 3760 6425
rect 3795 6325 3800 6425
rect 3700 6310 3800 6325
rect 3950 6425 4050 6440
rect 3950 6325 3955 6425
rect 3990 6325 4010 6425
rect 4045 6325 4050 6425
rect 3950 6310 4050 6325
rect 4200 6425 4300 6440
rect 4200 6325 4205 6425
rect 4240 6325 4260 6425
rect 4295 6325 4300 6425
rect 4200 6310 4300 6325
rect 4450 6425 4550 6440
rect 4450 6325 4455 6425
rect 4490 6325 4510 6425
rect 4545 6325 4550 6425
rect 4450 6310 4550 6325
rect 4700 6425 4800 6440
rect 4700 6325 4705 6425
rect 4740 6325 4760 6425
rect 4795 6325 4800 6425
rect 4700 6310 4800 6325
rect 4950 6425 5050 6440
rect 4950 6325 4955 6425
rect 4990 6325 5010 6425
rect 5045 6325 5050 6425
rect 4950 6310 5050 6325
rect 5200 6425 5300 6440
rect 5200 6325 5205 6425
rect 5240 6325 5260 6425
rect 5295 6325 5300 6425
rect 5200 6310 5300 6325
rect 5450 6425 5550 6440
rect 5450 6325 5455 6425
rect 5490 6325 5510 6425
rect 5545 6325 5550 6425
rect 5450 6310 5550 6325
rect 5700 6425 5800 6440
rect 5700 6325 5705 6425
rect 5740 6325 5760 6425
rect 5795 6325 5800 6425
rect 5700 6310 5800 6325
rect 5950 6425 6050 6440
rect 5950 6325 5955 6425
rect 5990 6325 6010 6425
rect 6045 6325 6050 6425
rect 5950 6310 6050 6325
rect 6200 6425 6300 6440
rect 6200 6325 6205 6425
rect 6240 6325 6260 6425
rect 6295 6325 6300 6425
rect 6200 6310 6300 6325
rect 6450 6425 6550 6440
rect 6450 6325 6455 6425
rect 6490 6325 6510 6425
rect 6545 6325 6550 6425
rect 6450 6310 6550 6325
rect 6700 6425 6800 6440
rect 6700 6325 6705 6425
rect 6740 6325 6760 6425
rect 6795 6325 6800 6425
rect 6700 6310 6800 6325
rect 6950 6425 7050 6440
rect 6950 6325 6955 6425
rect 6990 6325 7010 6425
rect 7045 6325 7050 6425
rect 6950 6310 7050 6325
rect 7200 6425 7300 6440
rect 7200 6325 7205 6425
rect 7240 6325 7260 6425
rect 7295 6325 7300 6425
rect 7200 6310 7300 6325
rect 7450 6425 7550 6440
rect 7450 6325 7455 6425
rect 7490 6325 7510 6425
rect 7545 6325 7550 6425
rect 7450 6310 7550 6325
rect 7700 6425 7800 6440
rect 7700 6325 7705 6425
rect 7740 6325 7760 6425
rect 7795 6325 7800 6425
rect 7700 6310 7800 6325
rect 7950 6425 8000 6440
rect 7950 6325 7955 6425
rect 7990 6325 8000 6425
rect 7950 6310 8000 6325
rect 0 6300 60 6310
rect 190 6300 310 6310
rect 440 6300 560 6310
rect 690 6300 810 6310
rect 940 6300 1060 6310
rect 1190 6300 1310 6310
rect 1440 6300 1560 6310
rect 1690 6300 1810 6310
rect 1940 6300 2060 6310
rect 2190 6300 2310 6310
rect 2440 6300 2560 6310
rect 2690 6300 2810 6310
rect 2940 6300 3060 6310
rect 3190 6300 3310 6310
rect 3440 6300 3560 6310
rect 3690 6300 3810 6310
rect 3940 6300 4060 6310
rect 4190 6300 4310 6310
rect 4440 6300 4560 6310
rect 4690 6300 4810 6310
rect 4940 6300 5060 6310
rect 5190 6300 5310 6310
rect 5440 6300 5560 6310
rect 5690 6300 5810 6310
rect 5940 6300 6060 6310
rect 6190 6300 6310 6310
rect 6440 6300 6560 6310
rect 6690 6300 6810 6310
rect 6940 6300 7060 6310
rect 7190 6300 7310 6310
rect 7440 6300 7560 6310
rect 7690 6300 7810 6310
rect 7940 6300 8000 6310
rect 0 6295 200 6300
rect 0 6260 75 6295
rect 175 6260 200 6295
rect 0 6240 200 6260
rect 0 6205 75 6240
rect 175 6205 200 6240
rect 0 6200 200 6205
rect 300 6295 450 6300
rect 300 6260 325 6295
rect 425 6260 450 6295
rect 300 6240 450 6260
rect 300 6205 325 6240
rect 425 6205 450 6240
rect 300 6200 450 6205
rect 550 6295 700 6300
rect 550 6260 575 6295
rect 675 6260 700 6295
rect 550 6240 700 6260
rect 550 6205 575 6240
rect 675 6205 700 6240
rect 550 6200 700 6205
rect 800 6295 1200 6300
rect 800 6260 825 6295
rect 925 6260 1075 6295
rect 1175 6260 1200 6295
rect 800 6240 1200 6260
rect 800 6205 825 6240
rect 925 6205 1075 6240
rect 1175 6205 1200 6240
rect 800 6200 1200 6205
rect 1300 6295 1450 6300
rect 1300 6260 1325 6295
rect 1425 6260 1450 6295
rect 1300 6240 1450 6260
rect 1300 6205 1325 6240
rect 1425 6205 1450 6240
rect 1300 6200 1450 6205
rect 1550 6295 1700 6300
rect 1550 6260 1575 6295
rect 1675 6260 1700 6295
rect 1550 6240 1700 6260
rect 1550 6205 1575 6240
rect 1675 6205 1700 6240
rect 1550 6200 1700 6205
rect 1800 6295 2200 6300
rect 1800 6260 1825 6295
rect 1925 6260 2075 6295
rect 2175 6260 2200 6295
rect 1800 6240 2200 6260
rect 1800 6205 1825 6240
rect 1925 6205 2075 6240
rect 2175 6205 2200 6240
rect 1800 6200 2200 6205
rect 2300 6295 2450 6300
rect 2300 6260 2325 6295
rect 2425 6260 2450 6295
rect 2300 6240 2450 6260
rect 2300 6205 2325 6240
rect 2425 6205 2450 6240
rect 2300 6200 2450 6205
rect 2550 6295 2700 6300
rect 2550 6260 2575 6295
rect 2675 6260 2700 6295
rect 2550 6240 2700 6260
rect 2550 6205 2575 6240
rect 2675 6205 2700 6240
rect 2550 6200 2700 6205
rect 2800 6295 3200 6300
rect 2800 6260 2825 6295
rect 2925 6260 3075 6295
rect 3175 6260 3200 6295
rect 2800 6240 3200 6260
rect 2800 6205 2825 6240
rect 2925 6205 3075 6240
rect 3175 6205 3200 6240
rect 2800 6200 3200 6205
rect 3300 6295 3450 6300
rect 3300 6260 3325 6295
rect 3425 6260 3450 6295
rect 3300 6240 3450 6260
rect 3300 6205 3325 6240
rect 3425 6205 3450 6240
rect 3300 6200 3450 6205
rect 3550 6295 3700 6300
rect 3550 6260 3575 6295
rect 3675 6260 3700 6295
rect 3550 6240 3700 6260
rect 3550 6205 3575 6240
rect 3675 6205 3700 6240
rect 3550 6200 3700 6205
rect 3800 6295 4200 6300
rect 3800 6260 3825 6295
rect 3925 6260 4075 6295
rect 4175 6260 4200 6295
rect 3800 6240 4200 6260
rect 3800 6205 3825 6240
rect 3925 6205 4075 6240
rect 4175 6205 4200 6240
rect 3800 6200 4200 6205
rect 4300 6295 4450 6300
rect 4300 6260 4325 6295
rect 4425 6260 4450 6295
rect 4300 6240 4450 6260
rect 4300 6205 4325 6240
rect 4425 6205 4450 6240
rect 4300 6200 4450 6205
rect 4550 6295 4700 6300
rect 4550 6260 4575 6295
rect 4675 6260 4700 6295
rect 4550 6240 4700 6260
rect 4550 6205 4575 6240
rect 4675 6205 4700 6240
rect 4550 6200 4700 6205
rect 4800 6295 5200 6300
rect 4800 6260 4825 6295
rect 4925 6260 5075 6295
rect 5175 6260 5200 6295
rect 4800 6240 5200 6260
rect 4800 6205 4825 6240
rect 4925 6205 5075 6240
rect 5175 6205 5200 6240
rect 4800 6200 5200 6205
rect 5300 6295 5450 6300
rect 5300 6260 5325 6295
rect 5425 6260 5450 6295
rect 5300 6240 5450 6260
rect 5300 6205 5325 6240
rect 5425 6205 5450 6240
rect 5300 6200 5450 6205
rect 5550 6295 5700 6300
rect 5550 6260 5575 6295
rect 5675 6260 5700 6295
rect 5550 6240 5700 6260
rect 5550 6205 5575 6240
rect 5675 6205 5700 6240
rect 5550 6200 5700 6205
rect 5800 6295 6200 6300
rect 5800 6260 5825 6295
rect 5925 6260 6075 6295
rect 6175 6260 6200 6295
rect 5800 6240 6200 6260
rect 5800 6205 5825 6240
rect 5925 6205 6075 6240
rect 6175 6205 6200 6240
rect 5800 6200 6200 6205
rect 6300 6295 6450 6300
rect 6300 6260 6325 6295
rect 6425 6260 6450 6295
rect 6300 6240 6450 6260
rect 6300 6205 6325 6240
rect 6425 6205 6450 6240
rect 6300 6200 6450 6205
rect 6550 6295 6700 6300
rect 6550 6260 6575 6295
rect 6675 6260 6700 6295
rect 6550 6240 6700 6260
rect 6550 6205 6575 6240
rect 6675 6205 6700 6240
rect 6550 6200 6700 6205
rect 6800 6295 7200 6300
rect 6800 6260 6825 6295
rect 6925 6260 7075 6295
rect 7175 6260 7200 6295
rect 6800 6240 7200 6260
rect 6800 6205 6825 6240
rect 6925 6205 7075 6240
rect 7175 6205 7200 6240
rect 6800 6200 7200 6205
rect 7300 6295 7450 6300
rect 7300 6260 7325 6295
rect 7425 6260 7450 6295
rect 7300 6240 7450 6260
rect 7300 6205 7325 6240
rect 7425 6205 7450 6240
rect 7300 6200 7450 6205
rect 7550 6295 7700 6300
rect 7550 6260 7575 6295
rect 7675 6260 7700 6295
rect 7550 6240 7700 6260
rect 7550 6205 7575 6240
rect 7675 6205 7700 6240
rect 7550 6200 7700 6205
rect 7800 6295 8000 6300
rect 7800 6260 7825 6295
rect 7925 6260 8000 6295
rect 7800 6240 8000 6260
rect 7800 6205 7825 6240
rect 7925 6205 8000 6240
rect 7800 6200 8000 6205
rect 0 6190 60 6200
rect 190 6190 310 6200
rect 440 6190 560 6200
rect 690 6190 810 6200
rect 940 6190 1060 6200
rect 1190 6190 1310 6200
rect 1440 6190 1560 6200
rect 1690 6190 1810 6200
rect 1940 6190 2060 6200
rect 2190 6190 2310 6200
rect 2440 6190 2560 6200
rect 2690 6190 2810 6200
rect 2940 6190 3060 6200
rect 3190 6190 3310 6200
rect 3440 6190 3560 6200
rect 3690 6190 3810 6200
rect 3940 6190 4060 6200
rect 4190 6190 4310 6200
rect 4440 6190 4560 6200
rect 4690 6190 4810 6200
rect 4940 6190 5060 6200
rect 5190 6190 5310 6200
rect 5440 6190 5560 6200
rect 5690 6190 5810 6200
rect 5940 6190 6060 6200
rect 6190 6190 6310 6200
rect 6440 6190 6560 6200
rect 6690 6190 6810 6200
rect 6940 6190 7060 6200
rect 7190 6190 7310 6200
rect 7440 6190 7560 6200
rect 7690 6190 7810 6200
rect 7940 6190 8000 6200
rect 0 6175 50 6190
rect 0 6075 10 6175
rect 45 6075 50 6175
rect 0 6060 50 6075
rect 200 6175 300 6190
rect 200 6075 205 6175
rect 240 6075 260 6175
rect 295 6075 300 6175
rect 200 6060 300 6075
rect 450 6175 550 6190
rect 450 6075 455 6175
rect 490 6075 510 6175
rect 545 6075 550 6175
rect 450 6060 550 6075
rect 700 6175 800 6190
rect 700 6075 705 6175
rect 740 6075 760 6175
rect 795 6075 800 6175
rect 700 6060 800 6075
rect 950 6175 1050 6190
rect 950 6075 955 6175
rect 990 6075 1010 6175
rect 1045 6075 1050 6175
rect 950 6060 1050 6075
rect 1200 6175 1300 6190
rect 1200 6075 1205 6175
rect 1240 6075 1260 6175
rect 1295 6075 1300 6175
rect 1200 6060 1300 6075
rect 1450 6175 1550 6190
rect 1450 6075 1455 6175
rect 1490 6075 1510 6175
rect 1545 6075 1550 6175
rect 1450 6060 1550 6075
rect 1700 6175 1800 6190
rect 1700 6075 1705 6175
rect 1740 6075 1760 6175
rect 1795 6075 1800 6175
rect 1700 6060 1800 6075
rect 1950 6175 2050 6190
rect 1950 6075 1955 6175
rect 1990 6075 2010 6175
rect 2045 6075 2050 6175
rect 1950 6060 2050 6075
rect 2200 6175 2300 6190
rect 2200 6075 2205 6175
rect 2240 6075 2260 6175
rect 2295 6075 2300 6175
rect 2200 6060 2300 6075
rect 2450 6175 2550 6190
rect 2450 6075 2455 6175
rect 2490 6075 2510 6175
rect 2545 6075 2550 6175
rect 2450 6060 2550 6075
rect 2700 6175 2800 6190
rect 2700 6075 2705 6175
rect 2740 6075 2760 6175
rect 2795 6075 2800 6175
rect 2700 6060 2800 6075
rect 2950 6175 3050 6190
rect 2950 6075 2955 6175
rect 2990 6075 3010 6175
rect 3045 6075 3050 6175
rect 2950 6060 3050 6075
rect 3200 6175 3300 6190
rect 3200 6075 3205 6175
rect 3240 6075 3260 6175
rect 3295 6075 3300 6175
rect 3200 6060 3300 6075
rect 3450 6175 3550 6190
rect 3450 6075 3455 6175
rect 3490 6075 3510 6175
rect 3545 6075 3550 6175
rect 3450 6060 3550 6075
rect 3700 6175 3800 6190
rect 3700 6075 3705 6175
rect 3740 6075 3760 6175
rect 3795 6075 3800 6175
rect 3700 6060 3800 6075
rect 3950 6175 4050 6190
rect 3950 6075 3955 6175
rect 3990 6075 4010 6175
rect 4045 6075 4050 6175
rect 3950 6060 4050 6075
rect 4200 6175 4300 6190
rect 4200 6075 4205 6175
rect 4240 6075 4260 6175
rect 4295 6075 4300 6175
rect 4200 6060 4300 6075
rect 4450 6175 4550 6190
rect 4450 6075 4455 6175
rect 4490 6075 4510 6175
rect 4545 6075 4550 6175
rect 4450 6060 4550 6075
rect 4700 6175 4800 6190
rect 4700 6075 4705 6175
rect 4740 6075 4760 6175
rect 4795 6075 4800 6175
rect 4700 6060 4800 6075
rect 4950 6175 5050 6190
rect 4950 6075 4955 6175
rect 4990 6075 5010 6175
rect 5045 6075 5050 6175
rect 4950 6060 5050 6075
rect 5200 6175 5300 6190
rect 5200 6075 5205 6175
rect 5240 6075 5260 6175
rect 5295 6075 5300 6175
rect 5200 6060 5300 6075
rect 5450 6175 5550 6190
rect 5450 6075 5455 6175
rect 5490 6075 5510 6175
rect 5545 6075 5550 6175
rect 5450 6060 5550 6075
rect 5700 6175 5800 6190
rect 5700 6075 5705 6175
rect 5740 6075 5760 6175
rect 5795 6075 5800 6175
rect 5700 6060 5800 6075
rect 5950 6175 6050 6190
rect 5950 6075 5955 6175
rect 5990 6075 6010 6175
rect 6045 6075 6050 6175
rect 5950 6060 6050 6075
rect 6200 6175 6300 6190
rect 6200 6075 6205 6175
rect 6240 6075 6260 6175
rect 6295 6075 6300 6175
rect 6200 6060 6300 6075
rect 6450 6175 6550 6190
rect 6450 6075 6455 6175
rect 6490 6075 6510 6175
rect 6545 6075 6550 6175
rect 6450 6060 6550 6075
rect 6700 6175 6800 6190
rect 6700 6075 6705 6175
rect 6740 6075 6760 6175
rect 6795 6075 6800 6175
rect 6700 6060 6800 6075
rect 6950 6175 7050 6190
rect 6950 6075 6955 6175
rect 6990 6075 7010 6175
rect 7045 6075 7050 6175
rect 6950 6060 7050 6075
rect 7200 6175 7300 6190
rect 7200 6075 7205 6175
rect 7240 6075 7260 6175
rect 7295 6075 7300 6175
rect 7200 6060 7300 6075
rect 7450 6175 7550 6190
rect 7450 6075 7455 6175
rect 7490 6075 7510 6175
rect 7545 6075 7550 6175
rect 7450 6060 7550 6075
rect 7700 6175 7800 6190
rect 7700 6075 7705 6175
rect 7740 6075 7760 6175
rect 7795 6075 7800 6175
rect 7700 6060 7800 6075
rect 7950 6175 8000 6190
rect 7950 6075 7955 6175
rect 7990 6075 8000 6175
rect 7950 6060 8000 6075
rect 0 6050 60 6060
rect 190 6050 310 6060
rect 440 6050 560 6060
rect 690 6050 810 6060
rect 940 6050 1060 6060
rect 1190 6050 1310 6060
rect 1440 6050 1560 6060
rect 1690 6050 1810 6060
rect 1940 6050 2060 6060
rect 2190 6050 2310 6060
rect 2440 6050 2560 6060
rect 2690 6050 2810 6060
rect 2940 6050 3060 6060
rect 3190 6050 3310 6060
rect 3440 6050 3560 6060
rect 3690 6050 3810 6060
rect 3940 6050 4060 6060
rect 4190 6050 4310 6060
rect 4440 6050 4560 6060
rect 4690 6050 4810 6060
rect 4940 6050 5060 6060
rect 5190 6050 5310 6060
rect 5440 6050 5560 6060
rect 5690 6050 5810 6060
rect 5940 6050 6060 6060
rect 6190 6050 6310 6060
rect 6440 6050 6560 6060
rect 6690 6050 6810 6060
rect 6940 6050 7060 6060
rect 7190 6050 7310 6060
rect 7440 6050 7560 6060
rect 7690 6050 7810 6060
rect 7940 6050 8000 6060
rect 0 6045 8000 6050
rect 0 6010 75 6045
rect 175 6010 325 6045
rect 425 6010 575 6045
rect 675 6010 825 6045
rect 925 6010 1075 6045
rect 1175 6010 1325 6045
rect 1425 6010 1575 6045
rect 1675 6010 1825 6045
rect 1925 6010 2075 6045
rect 2175 6010 2325 6045
rect 2425 6010 2575 6045
rect 2675 6010 2825 6045
rect 2925 6010 3075 6045
rect 3175 6010 3325 6045
rect 3425 6010 3575 6045
rect 3675 6010 3825 6045
rect 3925 6010 4075 6045
rect 4175 6010 4325 6045
rect 4425 6010 4575 6045
rect 4675 6010 4825 6045
rect 4925 6010 5075 6045
rect 5175 6010 5325 6045
rect 5425 6010 5575 6045
rect 5675 6010 5825 6045
rect 5925 6010 6075 6045
rect 6175 6010 6325 6045
rect 6425 6010 6575 6045
rect 6675 6010 6825 6045
rect 6925 6010 7075 6045
rect 7175 6010 7325 6045
rect 7425 6010 7575 6045
rect 7675 6010 7825 6045
rect 7925 6010 8000 6045
rect 0 5990 8000 6010
rect 0 5955 75 5990
rect 175 5955 325 5990
rect 425 5955 575 5990
rect 675 5955 825 5990
rect 925 5955 1075 5990
rect 1175 5955 1325 5990
rect 1425 5955 1575 5990
rect 1675 5955 1825 5990
rect 1925 5955 2075 5990
rect 2175 5955 2325 5990
rect 2425 5955 2575 5990
rect 2675 5955 2825 5990
rect 2925 5955 3075 5990
rect 3175 5955 3325 5990
rect 3425 5955 3575 5990
rect 3675 5955 3825 5990
rect 3925 5955 4075 5990
rect 4175 5955 4325 5990
rect 4425 5955 4575 5990
rect 4675 5955 4825 5990
rect 4925 5955 5075 5990
rect 5175 5955 5325 5990
rect 5425 5955 5575 5990
rect 5675 5955 5825 5990
rect 5925 5955 6075 5990
rect 6175 5955 6325 5990
rect 6425 5955 6575 5990
rect 6675 5955 6825 5990
rect 6925 5955 7075 5990
rect 7175 5955 7325 5990
rect 7425 5955 7575 5990
rect 7675 5955 7825 5990
rect 7925 5955 8000 5990
rect 0 5950 8000 5955
rect 0 5940 60 5950
rect 190 5940 310 5950
rect 440 5940 560 5950
rect 690 5940 810 5950
rect 940 5940 1060 5950
rect 1190 5940 1310 5950
rect 1440 5940 1560 5950
rect 1690 5940 1810 5950
rect 1940 5940 2060 5950
rect 2190 5940 2310 5950
rect 2440 5940 2560 5950
rect 2690 5940 2810 5950
rect 2940 5940 3060 5950
rect 3190 5940 3310 5950
rect 3440 5940 3560 5950
rect 3690 5940 3810 5950
rect 3940 5940 4060 5950
rect 4190 5940 4310 5950
rect 4440 5940 4560 5950
rect 4690 5940 4810 5950
rect 4940 5940 5060 5950
rect 5190 5940 5310 5950
rect 5440 5940 5560 5950
rect 5690 5940 5810 5950
rect 5940 5940 6060 5950
rect 6190 5940 6310 5950
rect 6440 5940 6560 5950
rect 6690 5940 6810 5950
rect 6940 5940 7060 5950
rect 7190 5940 7310 5950
rect 7440 5940 7560 5950
rect 7690 5940 7810 5950
rect 7940 5940 8000 5950
rect 0 5925 50 5940
rect 0 5825 10 5925
rect 45 5825 50 5925
rect 0 5810 50 5825
rect 200 5925 300 5940
rect 200 5825 205 5925
rect 240 5825 260 5925
rect 295 5825 300 5925
rect 200 5810 300 5825
rect 450 5925 550 5940
rect 450 5825 455 5925
rect 490 5825 510 5925
rect 545 5825 550 5925
rect 450 5810 550 5825
rect 700 5925 800 5940
rect 700 5825 705 5925
rect 740 5825 760 5925
rect 795 5825 800 5925
rect 700 5810 800 5825
rect 950 5925 1050 5940
rect 950 5825 955 5925
rect 990 5825 1010 5925
rect 1045 5825 1050 5925
rect 950 5810 1050 5825
rect 1200 5925 1300 5940
rect 1200 5825 1205 5925
rect 1240 5825 1260 5925
rect 1295 5825 1300 5925
rect 1200 5810 1300 5825
rect 1450 5925 1550 5940
rect 1450 5825 1455 5925
rect 1490 5825 1510 5925
rect 1545 5825 1550 5925
rect 1450 5810 1550 5825
rect 1700 5925 1800 5940
rect 1700 5825 1705 5925
rect 1740 5825 1760 5925
rect 1795 5825 1800 5925
rect 1700 5810 1800 5825
rect 1950 5925 2050 5940
rect 1950 5825 1955 5925
rect 1990 5825 2010 5925
rect 2045 5825 2050 5925
rect 1950 5810 2050 5825
rect 2200 5925 2300 5940
rect 2200 5825 2205 5925
rect 2240 5825 2260 5925
rect 2295 5825 2300 5925
rect 2200 5810 2300 5825
rect 2450 5925 2550 5940
rect 2450 5825 2455 5925
rect 2490 5825 2510 5925
rect 2545 5825 2550 5925
rect 2450 5810 2550 5825
rect 2700 5925 2800 5940
rect 2700 5825 2705 5925
rect 2740 5825 2760 5925
rect 2795 5825 2800 5925
rect 2700 5810 2800 5825
rect 2950 5925 3050 5940
rect 2950 5825 2955 5925
rect 2990 5825 3010 5925
rect 3045 5825 3050 5925
rect 2950 5810 3050 5825
rect 3200 5925 3300 5940
rect 3200 5825 3205 5925
rect 3240 5825 3260 5925
rect 3295 5825 3300 5925
rect 3200 5810 3300 5825
rect 3450 5925 3550 5940
rect 3450 5825 3455 5925
rect 3490 5825 3510 5925
rect 3545 5825 3550 5925
rect 3450 5810 3550 5825
rect 3700 5925 3800 5940
rect 3700 5825 3705 5925
rect 3740 5825 3760 5925
rect 3795 5825 3800 5925
rect 3700 5810 3800 5825
rect 3950 5925 4050 5940
rect 3950 5825 3955 5925
rect 3990 5825 4010 5925
rect 4045 5825 4050 5925
rect 3950 5810 4050 5825
rect 4200 5925 4300 5940
rect 4200 5825 4205 5925
rect 4240 5825 4260 5925
rect 4295 5825 4300 5925
rect 4200 5810 4300 5825
rect 4450 5925 4550 5940
rect 4450 5825 4455 5925
rect 4490 5825 4510 5925
rect 4545 5825 4550 5925
rect 4450 5810 4550 5825
rect 4700 5925 4800 5940
rect 4700 5825 4705 5925
rect 4740 5825 4760 5925
rect 4795 5825 4800 5925
rect 4700 5810 4800 5825
rect 4950 5925 5050 5940
rect 4950 5825 4955 5925
rect 4990 5825 5010 5925
rect 5045 5825 5050 5925
rect 4950 5810 5050 5825
rect 5200 5925 5300 5940
rect 5200 5825 5205 5925
rect 5240 5825 5260 5925
rect 5295 5825 5300 5925
rect 5200 5810 5300 5825
rect 5450 5925 5550 5940
rect 5450 5825 5455 5925
rect 5490 5825 5510 5925
rect 5545 5825 5550 5925
rect 5450 5810 5550 5825
rect 5700 5925 5800 5940
rect 5700 5825 5705 5925
rect 5740 5825 5760 5925
rect 5795 5825 5800 5925
rect 5700 5810 5800 5825
rect 5950 5925 6050 5940
rect 5950 5825 5955 5925
rect 5990 5825 6010 5925
rect 6045 5825 6050 5925
rect 5950 5810 6050 5825
rect 6200 5925 6300 5940
rect 6200 5825 6205 5925
rect 6240 5825 6260 5925
rect 6295 5825 6300 5925
rect 6200 5810 6300 5825
rect 6450 5925 6550 5940
rect 6450 5825 6455 5925
rect 6490 5825 6510 5925
rect 6545 5825 6550 5925
rect 6450 5810 6550 5825
rect 6700 5925 6800 5940
rect 6700 5825 6705 5925
rect 6740 5825 6760 5925
rect 6795 5825 6800 5925
rect 6700 5810 6800 5825
rect 6950 5925 7050 5940
rect 6950 5825 6955 5925
rect 6990 5825 7010 5925
rect 7045 5825 7050 5925
rect 6950 5810 7050 5825
rect 7200 5925 7300 5940
rect 7200 5825 7205 5925
rect 7240 5825 7260 5925
rect 7295 5825 7300 5925
rect 7200 5810 7300 5825
rect 7450 5925 7550 5940
rect 7450 5825 7455 5925
rect 7490 5825 7510 5925
rect 7545 5825 7550 5925
rect 7450 5810 7550 5825
rect 7700 5925 7800 5940
rect 7700 5825 7705 5925
rect 7740 5825 7760 5925
rect 7795 5825 7800 5925
rect 7700 5810 7800 5825
rect 7950 5925 8000 5940
rect 7950 5825 7955 5925
rect 7990 5825 8000 5925
rect 7950 5810 8000 5825
rect 0 5800 60 5810
rect 190 5800 310 5810
rect 440 5800 560 5810
rect 690 5800 810 5810
rect 940 5800 1060 5810
rect 1190 5800 1310 5810
rect 1440 5800 1560 5810
rect 1690 5800 1810 5810
rect 1940 5800 2060 5810
rect 2190 5800 2310 5810
rect 2440 5800 2560 5810
rect 2690 5800 2810 5810
rect 2940 5800 3060 5810
rect 3190 5800 3310 5810
rect 3440 5800 3560 5810
rect 3690 5800 3810 5810
rect 3940 5800 4060 5810
rect 4190 5800 4310 5810
rect 4440 5800 4560 5810
rect 4690 5800 4810 5810
rect 4940 5800 5060 5810
rect 5190 5800 5310 5810
rect 5440 5800 5560 5810
rect 5690 5800 5810 5810
rect 5940 5800 6060 5810
rect 6190 5800 6310 5810
rect 6440 5800 6560 5810
rect 6690 5800 6810 5810
rect 6940 5800 7060 5810
rect 7190 5800 7310 5810
rect 7440 5800 7560 5810
rect 7690 5800 7810 5810
rect 7940 5800 8000 5810
rect 0 5795 200 5800
rect 0 5760 75 5795
rect 175 5760 200 5795
rect 0 5740 200 5760
rect 0 5705 75 5740
rect 175 5705 200 5740
rect 0 5700 200 5705
rect 300 5795 450 5800
rect 300 5760 325 5795
rect 425 5760 450 5795
rect 300 5740 450 5760
rect 300 5705 325 5740
rect 425 5705 450 5740
rect 300 5700 450 5705
rect 550 5795 700 5800
rect 550 5760 575 5795
rect 675 5760 700 5795
rect 550 5740 700 5760
rect 550 5705 575 5740
rect 675 5705 700 5740
rect 550 5700 700 5705
rect 800 5795 1200 5800
rect 800 5760 825 5795
rect 925 5760 1075 5795
rect 1175 5760 1200 5795
rect 800 5740 1200 5760
rect 800 5705 825 5740
rect 925 5705 1075 5740
rect 1175 5705 1200 5740
rect 800 5700 1200 5705
rect 1300 5795 1450 5800
rect 1300 5760 1325 5795
rect 1425 5760 1450 5795
rect 1300 5740 1450 5760
rect 1300 5705 1325 5740
rect 1425 5705 1450 5740
rect 1300 5700 1450 5705
rect 1550 5795 1700 5800
rect 1550 5760 1575 5795
rect 1675 5760 1700 5795
rect 1550 5740 1700 5760
rect 1550 5705 1575 5740
rect 1675 5705 1700 5740
rect 1550 5700 1700 5705
rect 1800 5795 2200 5800
rect 1800 5760 1825 5795
rect 1925 5760 2075 5795
rect 2175 5760 2200 5795
rect 1800 5740 2200 5760
rect 1800 5705 1825 5740
rect 1925 5705 2075 5740
rect 2175 5705 2200 5740
rect 1800 5700 2200 5705
rect 2300 5795 2450 5800
rect 2300 5760 2325 5795
rect 2425 5760 2450 5795
rect 2300 5740 2450 5760
rect 2300 5705 2325 5740
rect 2425 5705 2450 5740
rect 2300 5700 2450 5705
rect 2550 5795 2700 5800
rect 2550 5760 2575 5795
rect 2675 5760 2700 5795
rect 2550 5740 2700 5760
rect 2550 5705 2575 5740
rect 2675 5705 2700 5740
rect 2550 5700 2700 5705
rect 2800 5795 3200 5800
rect 2800 5760 2825 5795
rect 2925 5760 3075 5795
rect 3175 5760 3200 5795
rect 2800 5740 3200 5760
rect 2800 5705 2825 5740
rect 2925 5705 3075 5740
rect 3175 5705 3200 5740
rect 2800 5700 3200 5705
rect 3300 5795 3450 5800
rect 3300 5760 3325 5795
rect 3425 5760 3450 5795
rect 3300 5740 3450 5760
rect 3300 5705 3325 5740
rect 3425 5705 3450 5740
rect 3300 5700 3450 5705
rect 3550 5795 3700 5800
rect 3550 5760 3575 5795
rect 3675 5760 3700 5795
rect 3550 5740 3700 5760
rect 3550 5705 3575 5740
rect 3675 5705 3700 5740
rect 3550 5700 3700 5705
rect 3800 5795 4200 5800
rect 3800 5760 3825 5795
rect 3925 5760 4075 5795
rect 4175 5760 4200 5795
rect 3800 5740 4200 5760
rect 3800 5705 3825 5740
rect 3925 5705 4075 5740
rect 4175 5705 4200 5740
rect 3800 5700 4200 5705
rect 4300 5795 4450 5800
rect 4300 5760 4325 5795
rect 4425 5760 4450 5795
rect 4300 5740 4450 5760
rect 4300 5705 4325 5740
rect 4425 5705 4450 5740
rect 4300 5700 4450 5705
rect 4550 5795 4700 5800
rect 4550 5760 4575 5795
rect 4675 5760 4700 5795
rect 4550 5740 4700 5760
rect 4550 5705 4575 5740
rect 4675 5705 4700 5740
rect 4550 5700 4700 5705
rect 4800 5795 5200 5800
rect 4800 5760 4825 5795
rect 4925 5760 5075 5795
rect 5175 5760 5200 5795
rect 4800 5740 5200 5760
rect 4800 5705 4825 5740
rect 4925 5705 5075 5740
rect 5175 5705 5200 5740
rect 4800 5700 5200 5705
rect 5300 5795 5450 5800
rect 5300 5760 5325 5795
rect 5425 5760 5450 5795
rect 5300 5740 5450 5760
rect 5300 5705 5325 5740
rect 5425 5705 5450 5740
rect 5300 5700 5450 5705
rect 5550 5795 5700 5800
rect 5550 5760 5575 5795
rect 5675 5760 5700 5795
rect 5550 5740 5700 5760
rect 5550 5705 5575 5740
rect 5675 5705 5700 5740
rect 5550 5700 5700 5705
rect 5800 5795 6200 5800
rect 5800 5760 5825 5795
rect 5925 5760 6075 5795
rect 6175 5760 6200 5795
rect 5800 5740 6200 5760
rect 5800 5705 5825 5740
rect 5925 5705 6075 5740
rect 6175 5705 6200 5740
rect 5800 5700 6200 5705
rect 6300 5795 6450 5800
rect 6300 5760 6325 5795
rect 6425 5760 6450 5795
rect 6300 5740 6450 5760
rect 6300 5705 6325 5740
rect 6425 5705 6450 5740
rect 6300 5700 6450 5705
rect 6550 5795 6700 5800
rect 6550 5760 6575 5795
rect 6675 5760 6700 5795
rect 6550 5740 6700 5760
rect 6550 5705 6575 5740
rect 6675 5705 6700 5740
rect 6550 5700 6700 5705
rect 6800 5795 7200 5800
rect 6800 5760 6825 5795
rect 6925 5760 7075 5795
rect 7175 5760 7200 5795
rect 6800 5740 7200 5760
rect 6800 5705 6825 5740
rect 6925 5705 7075 5740
rect 7175 5705 7200 5740
rect 6800 5700 7200 5705
rect 7300 5795 7450 5800
rect 7300 5760 7325 5795
rect 7425 5760 7450 5795
rect 7300 5740 7450 5760
rect 7300 5705 7325 5740
rect 7425 5705 7450 5740
rect 7300 5700 7450 5705
rect 7550 5795 7700 5800
rect 7550 5760 7575 5795
rect 7675 5760 7700 5795
rect 7550 5740 7700 5760
rect 7550 5705 7575 5740
rect 7675 5705 7700 5740
rect 7550 5700 7700 5705
rect 7800 5795 8000 5800
rect 7800 5760 7825 5795
rect 7925 5760 8000 5795
rect 7800 5740 8000 5760
rect 7800 5705 7825 5740
rect 7925 5705 8000 5740
rect 7800 5700 8000 5705
rect 0 5690 60 5700
rect 190 5690 310 5700
rect 440 5690 560 5700
rect 690 5690 810 5700
rect 940 5690 1060 5700
rect 1190 5690 1310 5700
rect 1440 5690 1560 5700
rect 1690 5690 1810 5700
rect 1940 5690 2060 5700
rect 2190 5690 2310 5700
rect 2440 5690 2560 5700
rect 2690 5690 2810 5700
rect 2940 5690 3060 5700
rect 3190 5690 3310 5700
rect 3440 5690 3560 5700
rect 3690 5690 3810 5700
rect 3940 5690 4060 5700
rect 4190 5690 4310 5700
rect 4440 5690 4560 5700
rect 4690 5690 4810 5700
rect 4940 5690 5060 5700
rect 5190 5690 5310 5700
rect 5440 5690 5560 5700
rect 5690 5690 5810 5700
rect 5940 5690 6060 5700
rect 6190 5690 6310 5700
rect 6440 5690 6560 5700
rect 6690 5690 6810 5700
rect 6940 5690 7060 5700
rect 7190 5690 7310 5700
rect 7440 5690 7560 5700
rect 7690 5690 7810 5700
rect 7940 5690 8000 5700
rect 0 5675 50 5690
rect 0 5575 10 5675
rect 45 5575 50 5675
rect 0 5560 50 5575
rect 200 5675 300 5690
rect 200 5575 205 5675
rect 240 5575 260 5675
rect 295 5575 300 5675
rect 200 5560 300 5575
rect 450 5675 550 5690
rect 450 5575 455 5675
rect 490 5575 510 5675
rect 545 5575 550 5675
rect 450 5560 550 5575
rect 700 5675 800 5690
rect 700 5575 705 5675
rect 740 5575 760 5675
rect 795 5575 800 5675
rect 700 5560 800 5575
rect 950 5675 1050 5690
rect 950 5575 955 5675
rect 990 5575 1010 5675
rect 1045 5575 1050 5675
rect 950 5560 1050 5575
rect 1200 5675 1300 5690
rect 1200 5575 1205 5675
rect 1240 5575 1260 5675
rect 1295 5575 1300 5675
rect 1200 5560 1300 5575
rect 1450 5675 1550 5690
rect 1450 5575 1455 5675
rect 1490 5575 1510 5675
rect 1545 5575 1550 5675
rect 1450 5560 1550 5575
rect 1700 5675 1800 5690
rect 1700 5575 1705 5675
rect 1740 5575 1760 5675
rect 1795 5575 1800 5675
rect 1700 5560 1800 5575
rect 1950 5675 2050 5690
rect 1950 5575 1955 5675
rect 1990 5575 2010 5675
rect 2045 5575 2050 5675
rect 1950 5560 2050 5575
rect 2200 5675 2300 5690
rect 2200 5575 2205 5675
rect 2240 5575 2260 5675
rect 2295 5575 2300 5675
rect 2200 5560 2300 5575
rect 2450 5675 2550 5690
rect 2450 5575 2455 5675
rect 2490 5575 2510 5675
rect 2545 5575 2550 5675
rect 2450 5560 2550 5575
rect 2700 5675 2800 5690
rect 2700 5575 2705 5675
rect 2740 5575 2760 5675
rect 2795 5575 2800 5675
rect 2700 5560 2800 5575
rect 2950 5675 3050 5690
rect 2950 5575 2955 5675
rect 2990 5575 3010 5675
rect 3045 5575 3050 5675
rect 2950 5560 3050 5575
rect 3200 5675 3300 5690
rect 3200 5575 3205 5675
rect 3240 5575 3260 5675
rect 3295 5575 3300 5675
rect 3200 5560 3300 5575
rect 3450 5675 3550 5690
rect 3450 5575 3455 5675
rect 3490 5575 3510 5675
rect 3545 5575 3550 5675
rect 3450 5560 3550 5575
rect 3700 5675 3800 5690
rect 3700 5575 3705 5675
rect 3740 5575 3760 5675
rect 3795 5575 3800 5675
rect 3700 5560 3800 5575
rect 3950 5675 4050 5690
rect 3950 5575 3955 5675
rect 3990 5575 4010 5675
rect 4045 5575 4050 5675
rect 3950 5560 4050 5575
rect 4200 5675 4300 5690
rect 4200 5575 4205 5675
rect 4240 5575 4260 5675
rect 4295 5575 4300 5675
rect 4200 5560 4300 5575
rect 4450 5675 4550 5690
rect 4450 5575 4455 5675
rect 4490 5575 4510 5675
rect 4545 5575 4550 5675
rect 4450 5560 4550 5575
rect 4700 5675 4800 5690
rect 4700 5575 4705 5675
rect 4740 5575 4760 5675
rect 4795 5575 4800 5675
rect 4700 5560 4800 5575
rect 4950 5675 5050 5690
rect 4950 5575 4955 5675
rect 4990 5575 5010 5675
rect 5045 5575 5050 5675
rect 4950 5560 5050 5575
rect 5200 5675 5300 5690
rect 5200 5575 5205 5675
rect 5240 5575 5260 5675
rect 5295 5575 5300 5675
rect 5200 5560 5300 5575
rect 5450 5675 5550 5690
rect 5450 5575 5455 5675
rect 5490 5575 5510 5675
rect 5545 5575 5550 5675
rect 5450 5560 5550 5575
rect 5700 5675 5800 5690
rect 5700 5575 5705 5675
rect 5740 5575 5760 5675
rect 5795 5575 5800 5675
rect 5700 5560 5800 5575
rect 5950 5675 6050 5690
rect 5950 5575 5955 5675
rect 5990 5575 6010 5675
rect 6045 5575 6050 5675
rect 5950 5560 6050 5575
rect 6200 5675 6300 5690
rect 6200 5575 6205 5675
rect 6240 5575 6260 5675
rect 6295 5575 6300 5675
rect 6200 5560 6300 5575
rect 6450 5675 6550 5690
rect 6450 5575 6455 5675
rect 6490 5575 6510 5675
rect 6545 5575 6550 5675
rect 6450 5560 6550 5575
rect 6700 5675 6800 5690
rect 6700 5575 6705 5675
rect 6740 5575 6760 5675
rect 6795 5575 6800 5675
rect 6700 5560 6800 5575
rect 6950 5675 7050 5690
rect 6950 5575 6955 5675
rect 6990 5575 7010 5675
rect 7045 5575 7050 5675
rect 6950 5560 7050 5575
rect 7200 5675 7300 5690
rect 7200 5575 7205 5675
rect 7240 5575 7260 5675
rect 7295 5575 7300 5675
rect 7200 5560 7300 5575
rect 7450 5675 7550 5690
rect 7450 5575 7455 5675
rect 7490 5575 7510 5675
rect 7545 5575 7550 5675
rect 7450 5560 7550 5575
rect 7700 5675 7800 5690
rect 7700 5575 7705 5675
rect 7740 5575 7760 5675
rect 7795 5575 7800 5675
rect 7700 5560 7800 5575
rect 7950 5675 8000 5690
rect 7950 5575 7955 5675
rect 7990 5575 8000 5675
rect 7950 5560 8000 5575
rect 0 5550 60 5560
rect 190 5550 310 5560
rect 440 5550 560 5560
rect 690 5550 810 5560
rect 940 5550 1060 5560
rect 1190 5550 1310 5560
rect 1440 5550 1560 5560
rect 1690 5550 1810 5560
rect 1940 5550 2060 5560
rect 2190 5550 2310 5560
rect 2440 5550 2560 5560
rect 2690 5550 2810 5560
rect 2940 5550 3060 5560
rect 3190 5550 3310 5560
rect 3440 5550 3560 5560
rect 3690 5550 3810 5560
rect 3940 5550 4060 5560
rect 4190 5550 4310 5560
rect 4440 5550 4560 5560
rect 4690 5550 4810 5560
rect 4940 5550 5060 5560
rect 5190 5550 5310 5560
rect 5440 5550 5560 5560
rect 5690 5550 5810 5560
rect 5940 5550 6060 5560
rect 6190 5550 6310 5560
rect 6440 5550 6560 5560
rect 6690 5550 6810 5560
rect 6940 5550 7060 5560
rect 7190 5550 7310 5560
rect 7440 5550 7560 5560
rect 7690 5550 7810 5560
rect 7940 5550 8000 5560
rect 0 5545 200 5550
rect 0 5510 75 5545
rect 175 5510 200 5545
rect 0 5490 200 5510
rect 0 5455 75 5490
rect 175 5455 200 5490
rect 0 5450 200 5455
rect 300 5545 450 5550
rect 300 5510 325 5545
rect 425 5510 450 5545
rect 300 5490 450 5510
rect 300 5455 325 5490
rect 425 5455 450 5490
rect 300 5450 450 5455
rect 550 5545 700 5550
rect 550 5510 575 5545
rect 675 5510 700 5545
rect 550 5490 700 5510
rect 550 5455 575 5490
rect 675 5455 700 5490
rect 550 5450 700 5455
rect 800 5545 950 5550
rect 800 5510 825 5545
rect 925 5510 950 5545
rect 800 5490 950 5510
rect 800 5455 825 5490
rect 925 5455 950 5490
rect 800 5450 950 5455
rect 1050 5545 1200 5550
rect 1050 5510 1075 5545
rect 1175 5510 1200 5545
rect 1050 5490 1200 5510
rect 1050 5455 1075 5490
rect 1175 5455 1200 5490
rect 1050 5450 1200 5455
rect 1300 5545 1450 5550
rect 1300 5510 1325 5545
rect 1425 5510 1450 5545
rect 1300 5490 1450 5510
rect 1300 5455 1325 5490
rect 1425 5455 1450 5490
rect 1300 5450 1450 5455
rect 1550 5545 1700 5550
rect 1550 5510 1575 5545
rect 1675 5510 1700 5545
rect 1550 5490 1700 5510
rect 1550 5455 1575 5490
rect 1675 5455 1700 5490
rect 1550 5450 1700 5455
rect 1800 5545 2200 5550
rect 1800 5510 1825 5545
rect 1925 5510 2075 5545
rect 2175 5510 2200 5545
rect 1800 5490 2200 5510
rect 1800 5455 1825 5490
rect 1925 5455 2075 5490
rect 2175 5455 2200 5490
rect 1800 5450 2200 5455
rect 2300 5545 2450 5550
rect 2300 5510 2325 5545
rect 2425 5510 2450 5545
rect 2300 5490 2450 5510
rect 2300 5455 2325 5490
rect 2425 5455 2450 5490
rect 2300 5450 2450 5455
rect 2550 5545 2700 5550
rect 2550 5510 2575 5545
rect 2675 5510 2700 5545
rect 2550 5490 2700 5510
rect 2550 5455 2575 5490
rect 2675 5455 2700 5490
rect 2550 5450 2700 5455
rect 2800 5545 2950 5550
rect 2800 5510 2825 5545
rect 2925 5510 2950 5545
rect 2800 5490 2950 5510
rect 2800 5455 2825 5490
rect 2925 5455 2950 5490
rect 2800 5450 2950 5455
rect 3050 5545 3200 5550
rect 3050 5510 3075 5545
rect 3175 5510 3200 5545
rect 3050 5490 3200 5510
rect 3050 5455 3075 5490
rect 3175 5455 3200 5490
rect 3050 5450 3200 5455
rect 3300 5545 3450 5550
rect 3300 5510 3325 5545
rect 3425 5510 3450 5545
rect 3300 5490 3450 5510
rect 3300 5455 3325 5490
rect 3425 5455 3450 5490
rect 3300 5450 3450 5455
rect 3550 5545 3700 5550
rect 3550 5510 3575 5545
rect 3675 5510 3700 5545
rect 3550 5490 3700 5510
rect 3550 5455 3575 5490
rect 3675 5455 3700 5490
rect 3550 5450 3700 5455
rect 3800 5545 4200 5550
rect 3800 5510 3825 5545
rect 3925 5510 4075 5545
rect 4175 5510 4200 5545
rect 3800 5490 4200 5510
rect 3800 5455 3825 5490
rect 3925 5455 4075 5490
rect 4175 5455 4200 5490
rect 3800 5450 4200 5455
rect 4300 5545 4450 5550
rect 4300 5510 4325 5545
rect 4425 5510 4450 5545
rect 4300 5490 4450 5510
rect 4300 5455 4325 5490
rect 4425 5455 4450 5490
rect 4300 5450 4450 5455
rect 4550 5545 4700 5550
rect 4550 5510 4575 5545
rect 4675 5510 4700 5545
rect 4550 5490 4700 5510
rect 4550 5455 4575 5490
rect 4675 5455 4700 5490
rect 4550 5450 4700 5455
rect 4800 5545 4950 5550
rect 4800 5510 4825 5545
rect 4925 5510 4950 5545
rect 4800 5490 4950 5510
rect 4800 5455 4825 5490
rect 4925 5455 4950 5490
rect 4800 5450 4950 5455
rect 5050 5545 5200 5550
rect 5050 5510 5075 5545
rect 5175 5510 5200 5545
rect 5050 5490 5200 5510
rect 5050 5455 5075 5490
rect 5175 5455 5200 5490
rect 5050 5450 5200 5455
rect 5300 5545 5450 5550
rect 5300 5510 5325 5545
rect 5425 5510 5450 5545
rect 5300 5490 5450 5510
rect 5300 5455 5325 5490
rect 5425 5455 5450 5490
rect 5300 5450 5450 5455
rect 5550 5545 5700 5550
rect 5550 5510 5575 5545
rect 5675 5510 5700 5545
rect 5550 5490 5700 5510
rect 5550 5455 5575 5490
rect 5675 5455 5700 5490
rect 5550 5450 5700 5455
rect 5800 5545 6200 5550
rect 5800 5510 5825 5545
rect 5925 5510 6075 5545
rect 6175 5510 6200 5545
rect 5800 5490 6200 5510
rect 5800 5455 5825 5490
rect 5925 5455 6075 5490
rect 6175 5455 6200 5490
rect 5800 5450 6200 5455
rect 6300 5545 6450 5550
rect 6300 5510 6325 5545
rect 6425 5510 6450 5545
rect 6300 5490 6450 5510
rect 6300 5455 6325 5490
rect 6425 5455 6450 5490
rect 6300 5450 6450 5455
rect 6550 5545 6700 5550
rect 6550 5510 6575 5545
rect 6675 5510 6700 5545
rect 6550 5490 6700 5510
rect 6550 5455 6575 5490
rect 6675 5455 6700 5490
rect 6550 5450 6700 5455
rect 6800 5545 6950 5550
rect 6800 5510 6825 5545
rect 6925 5510 6950 5545
rect 6800 5490 6950 5510
rect 6800 5455 6825 5490
rect 6925 5455 6950 5490
rect 6800 5450 6950 5455
rect 7050 5545 7200 5550
rect 7050 5510 7075 5545
rect 7175 5510 7200 5545
rect 7050 5490 7200 5510
rect 7050 5455 7075 5490
rect 7175 5455 7200 5490
rect 7050 5450 7200 5455
rect 7300 5545 7450 5550
rect 7300 5510 7325 5545
rect 7425 5510 7450 5545
rect 7300 5490 7450 5510
rect 7300 5455 7325 5490
rect 7425 5455 7450 5490
rect 7300 5450 7450 5455
rect 7550 5545 7700 5550
rect 7550 5510 7575 5545
rect 7675 5510 7700 5545
rect 7550 5490 7700 5510
rect 7550 5455 7575 5490
rect 7675 5455 7700 5490
rect 7550 5450 7700 5455
rect 7800 5545 8000 5550
rect 7800 5510 7825 5545
rect 7925 5510 8000 5545
rect 7800 5490 8000 5510
rect 7800 5455 7825 5490
rect 7925 5455 8000 5490
rect 7800 5450 8000 5455
rect 0 5440 60 5450
rect 190 5440 310 5450
rect 440 5440 560 5450
rect 690 5440 810 5450
rect 940 5440 1060 5450
rect 1190 5440 1310 5450
rect 1440 5440 1560 5450
rect 1690 5440 1810 5450
rect 1940 5440 2060 5450
rect 2190 5440 2310 5450
rect 2440 5440 2560 5450
rect 2690 5440 2810 5450
rect 2940 5440 3060 5450
rect 3190 5440 3310 5450
rect 3440 5440 3560 5450
rect 3690 5440 3810 5450
rect 3940 5440 4060 5450
rect 4190 5440 4310 5450
rect 4440 5440 4560 5450
rect 4690 5440 4810 5450
rect 4940 5440 5060 5450
rect 5190 5440 5310 5450
rect 5440 5440 5560 5450
rect 5690 5440 5810 5450
rect 5940 5440 6060 5450
rect 6190 5440 6310 5450
rect 6440 5440 6560 5450
rect 6690 5440 6810 5450
rect 6940 5440 7060 5450
rect 7190 5440 7310 5450
rect 7440 5440 7560 5450
rect 7690 5440 7810 5450
rect 7940 5440 8000 5450
rect 0 5425 50 5440
rect 0 5325 10 5425
rect 45 5325 50 5425
rect 0 5310 50 5325
rect 200 5425 300 5440
rect 200 5325 205 5425
rect 240 5325 260 5425
rect 295 5325 300 5425
rect 200 5310 300 5325
rect 450 5425 550 5440
rect 450 5325 455 5425
rect 490 5325 510 5425
rect 545 5325 550 5425
rect 450 5310 550 5325
rect 700 5425 800 5440
rect 700 5325 705 5425
rect 740 5325 760 5425
rect 795 5325 800 5425
rect 700 5310 800 5325
rect 950 5425 1050 5440
rect 950 5325 955 5425
rect 990 5325 1010 5425
rect 1045 5325 1050 5425
rect 950 5310 1050 5325
rect 1200 5425 1300 5440
rect 1200 5325 1205 5425
rect 1240 5325 1260 5425
rect 1295 5325 1300 5425
rect 1200 5310 1300 5325
rect 1450 5425 1550 5440
rect 1450 5325 1455 5425
rect 1490 5325 1510 5425
rect 1545 5325 1550 5425
rect 1450 5310 1550 5325
rect 1700 5425 1800 5440
rect 1700 5325 1705 5425
rect 1740 5325 1760 5425
rect 1795 5325 1800 5425
rect 1700 5310 1800 5325
rect 1950 5425 2050 5440
rect 1950 5325 1955 5425
rect 1990 5325 2010 5425
rect 2045 5325 2050 5425
rect 1950 5310 2050 5325
rect 2200 5425 2300 5440
rect 2200 5325 2205 5425
rect 2240 5325 2260 5425
rect 2295 5325 2300 5425
rect 2200 5310 2300 5325
rect 2450 5425 2550 5440
rect 2450 5325 2455 5425
rect 2490 5325 2510 5425
rect 2545 5325 2550 5425
rect 2450 5310 2550 5325
rect 2700 5425 2800 5440
rect 2700 5325 2705 5425
rect 2740 5325 2760 5425
rect 2795 5325 2800 5425
rect 2700 5310 2800 5325
rect 2950 5425 3050 5440
rect 2950 5325 2955 5425
rect 2990 5325 3010 5425
rect 3045 5325 3050 5425
rect 2950 5310 3050 5325
rect 3200 5425 3300 5440
rect 3200 5325 3205 5425
rect 3240 5325 3260 5425
rect 3295 5325 3300 5425
rect 3200 5310 3300 5325
rect 3450 5425 3550 5440
rect 3450 5325 3455 5425
rect 3490 5325 3510 5425
rect 3545 5325 3550 5425
rect 3450 5310 3550 5325
rect 3700 5425 3800 5440
rect 3700 5325 3705 5425
rect 3740 5325 3760 5425
rect 3795 5325 3800 5425
rect 3700 5310 3800 5325
rect 3950 5425 4050 5440
rect 3950 5325 3955 5425
rect 3990 5325 4010 5425
rect 4045 5325 4050 5425
rect 3950 5310 4050 5325
rect 4200 5425 4300 5440
rect 4200 5325 4205 5425
rect 4240 5325 4260 5425
rect 4295 5325 4300 5425
rect 4200 5310 4300 5325
rect 4450 5425 4550 5440
rect 4450 5325 4455 5425
rect 4490 5325 4510 5425
rect 4545 5325 4550 5425
rect 4450 5310 4550 5325
rect 4700 5425 4800 5440
rect 4700 5325 4705 5425
rect 4740 5325 4760 5425
rect 4795 5325 4800 5425
rect 4700 5310 4800 5325
rect 4950 5425 5050 5440
rect 4950 5325 4955 5425
rect 4990 5325 5010 5425
rect 5045 5325 5050 5425
rect 4950 5310 5050 5325
rect 5200 5425 5300 5440
rect 5200 5325 5205 5425
rect 5240 5325 5260 5425
rect 5295 5325 5300 5425
rect 5200 5310 5300 5325
rect 5450 5425 5550 5440
rect 5450 5325 5455 5425
rect 5490 5325 5510 5425
rect 5545 5325 5550 5425
rect 5450 5310 5550 5325
rect 5700 5425 5800 5440
rect 5700 5325 5705 5425
rect 5740 5325 5760 5425
rect 5795 5325 5800 5425
rect 5700 5310 5800 5325
rect 5950 5425 6050 5440
rect 5950 5325 5955 5425
rect 5990 5325 6010 5425
rect 6045 5325 6050 5425
rect 5950 5310 6050 5325
rect 6200 5425 6300 5440
rect 6200 5325 6205 5425
rect 6240 5325 6260 5425
rect 6295 5325 6300 5425
rect 6200 5310 6300 5325
rect 6450 5425 6550 5440
rect 6450 5325 6455 5425
rect 6490 5325 6510 5425
rect 6545 5325 6550 5425
rect 6450 5310 6550 5325
rect 6700 5425 6800 5440
rect 6700 5325 6705 5425
rect 6740 5325 6760 5425
rect 6795 5325 6800 5425
rect 6700 5310 6800 5325
rect 6950 5425 7050 5440
rect 6950 5325 6955 5425
rect 6990 5325 7010 5425
rect 7045 5325 7050 5425
rect 6950 5310 7050 5325
rect 7200 5425 7300 5440
rect 7200 5325 7205 5425
rect 7240 5325 7260 5425
rect 7295 5325 7300 5425
rect 7200 5310 7300 5325
rect 7450 5425 7550 5440
rect 7450 5325 7455 5425
rect 7490 5325 7510 5425
rect 7545 5325 7550 5425
rect 7450 5310 7550 5325
rect 7700 5425 7800 5440
rect 7700 5325 7705 5425
rect 7740 5325 7760 5425
rect 7795 5325 7800 5425
rect 7700 5310 7800 5325
rect 7950 5425 8000 5440
rect 7950 5325 7955 5425
rect 7990 5325 8000 5425
rect 7950 5310 8000 5325
rect 0 5300 60 5310
rect 190 5300 310 5310
rect 440 5300 560 5310
rect 690 5300 810 5310
rect 940 5300 1060 5310
rect 1190 5300 1310 5310
rect 1440 5300 1560 5310
rect 1690 5300 1810 5310
rect 1940 5300 2060 5310
rect 2190 5300 2310 5310
rect 2440 5300 2560 5310
rect 2690 5300 2810 5310
rect 2940 5300 3060 5310
rect 3190 5300 3310 5310
rect 3440 5300 3560 5310
rect 3690 5300 3810 5310
rect 3940 5300 4060 5310
rect 4190 5300 4310 5310
rect 4440 5300 4560 5310
rect 4690 5300 4810 5310
rect 4940 5300 5060 5310
rect 5190 5300 5310 5310
rect 5440 5300 5560 5310
rect 5690 5300 5810 5310
rect 5940 5300 6060 5310
rect 6190 5300 6310 5310
rect 6440 5300 6560 5310
rect 6690 5300 6810 5310
rect 6940 5300 7060 5310
rect 7190 5300 7310 5310
rect 7440 5300 7560 5310
rect 7690 5300 7810 5310
rect 7940 5300 8000 5310
rect 0 5295 200 5300
rect 0 5260 75 5295
rect 175 5260 200 5295
rect 0 5240 200 5260
rect 0 5205 75 5240
rect 175 5205 200 5240
rect 0 5200 200 5205
rect 300 5295 450 5300
rect 300 5260 325 5295
rect 425 5260 450 5295
rect 300 5240 450 5260
rect 300 5205 325 5240
rect 425 5205 450 5240
rect 300 5200 450 5205
rect 550 5295 700 5300
rect 550 5260 575 5295
rect 675 5260 700 5295
rect 550 5240 700 5260
rect 550 5205 575 5240
rect 675 5205 700 5240
rect 550 5200 700 5205
rect 800 5295 1200 5300
rect 800 5260 825 5295
rect 925 5260 1075 5295
rect 1175 5260 1200 5295
rect 800 5240 1200 5260
rect 800 5205 825 5240
rect 925 5205 1075 5240
rect 1175 5205 1200 5240
rect 800 5200 1200 5205
rect 1300 5295 1450 5300
rect 1300 5260 1325 5295
rect 1425 5260 1450 5295
rect 1300 5240 1450 5260
rect 1300 5205 1325 5240
rect 1425 5205 1450 5240
rect 1300 5200 1450 5205
rect 1550 5295 1700 5300
rect 1550 5260 1575 5295
rect 1675 5260 1700 5295
rect 1550 5240 1700 5260
rect 1550 5205 1575 5240
rect 1675 5205 1700 5240
rect 1550 5200 1700 5205
rect 1800 5295 2200 5300
rect 1800 5260 1825 5295
rect 1925 5260 2075 5295
rect 2175 5260 2200 5295
rect 1800 5240 2200 5260
rect 1800 5205 1825 5240
rect 1925 5205 2075 5240
rect 2175 5205 2200 5240
rect 1800 5200 2200 5205
rect 2300 5295 2450 5300
rect 2300 5260 2325 5295
rect 2425 5260 2450 5295
rect 2300 5240 2450 5260
rect 2300 5205 2325 5240
rect 2425 5205 2450 5240
rect 2300 5200 2450 5205
rect 2550 5295 2700 5300
rect 2550 5260 2575 5295
rect 2675 5260 2700 5295
rect 2550 5240 2700 5260
rect 2550 5205 2575 5240
rect 2675 5205 2700 5240
rect 2550 5200 2700 5205
rect 2800 5295 3200 5300
rect 2800 5260 2825 5295
rect 2925 5260 3075 5295
rect 3175 5260 3200 5295
rect 2800 5240 3200 5260
rect 2800 5205 2825 5240
rect 2925 5205 3075 5240
rect 3175 5205 3200 5240
rect 2800 5200 3200 5205
rect 3300 5295 3450 5300
rect 3300 5260 3325 5295
rect 3425 5260 3450 5295
rect 3300 5240 3450 5260
rect 3300 5205 3325 5240
rect 3425 5205 3450 5240
rect 3300 5200 3450 5205
rect 3550 5295 3700 5300
rect 3550 5260 3575 5295
rect 3675 5260 3700 5295
rect 3550 5240 3700 5260
rect 3550 5205 3575 5240
rect 3675 5205 3700 5240
rect 3550 5200 3700 5205
rect 3800 5295 4200 5300
rect 3800 5260 3825 5295
rect 3925 5260 4075 5295
rect 4175 5260 4200 5295
rect 3800 5240 4200 5260
rect 3800 5205 3825 5240
rect 3925 5205 4075 5240
rect 4175 5205 4200 5240
rect 3800 5200 4200 5205
rect 4300 5295 4450 5300
rect 4300 5260 4325 5295
rect 4425 5260 4450 5295
rect 4300 5240 4450 5260
rect 4300 5205 4325 5240
rect 4425 5205 4450 5240
rect 4300 5200 4450 5205
rect 4550 5295 4700 5300
rect 4550 5260 4575 5295
rect 4675 5260 4700 5295
rect 4550 5240 4700 5260
rect 4550 5205 4575 5240
rect 4675 5205 4700 5240
rect 4550 5200 4700 5205
rect 4800 5295 5200 5300
rect 4800 5260 4825 5295
rect 4925 5260 5075 5295
rect 5175 5260 5200 5295
rect 4800 5240 5200 5260
rect 4800 5205 4825 5240
rect 4925 5205 5075 5240
rect 5175 5205 5200 5240
rect 4800 5200 5200 5205
rect 5300 5295 5450 5300
rect 5300 5260 5325 5295
rect 5425 5260 5450 5295
rect 5300 5240 5450 5260
rect 5300 5205 5325 5240
rect 5425 5205 5450 5240
rect 5300 5200 5450 5205
rect 5550 5295 5700 5300
rect 5550 5260 5575 5295
rect 5675 5260 5700 5295
rect 5550 5240 5700 5260
rect 5550 5205 5575 5240
rect 5675 5205 5700 5240
rect 5550 5200 5700 5205
rect 5800 5295 6200 5300
rect 5800 5260 5825 5295
rect 5925 5260 6075 5295
rect 6175 5260 6200 5295
rect 5800 5240 6200 5260
rect 5800 5205 5825 5240
rect 5925 5205 6075 5240
rect 6175 5205 6200 5240
rect 5800 5200 6200 5205
rect 6300 5295 6450 5300
rect 6300 5260 6325 5295
rect 6425 5260 6450 5295
rect 6300 5240 6450 5260
rect 6300 5205 6325 5240
rect 6425 5205 6450 5240
rect 6300 5200 6450 5205
rect 6550 5295 6700 5300
rect 6550 5260 6575 5295
rect 6675 5260 6700 5295
rect 6550 5240 6700 5260
rect 6550 5205 6575 5240
rect 6675 5205 6700 5240
rect 6550 5200 6700 5205
rect 6800 5295 7200 5300
rect 6800 5260 6825 5295
rect 6925 5260 7075 5295
rect 7175 5260 7200 5295
rect 6800 5240 7200 5260
rect 6800 5205 6825 5240
rect 6925 5205 7075 5240
rect 7175 5205 7200 5240
rect 6800 5200 7200 5205
rect 7300 5295 7450 5300
rect 7300 5260 7325 5295
rect 7425 5260 7450 5295
rect 7300 5240 7450 5260
rect 7300 5205 7325 5240
rect 7425 5205 7450 5240
rect 7300 5200 7450 5205
rect 7550 5295 7700 5300
rect 7550 5260 7575 5295
rect 7675 5260 7700 5295
rect 7550 5240 7700 5260
rect 7550 5205 7575 5240
rect 7675 5205 7700 5240
rect 7550 5200 7700 5205
rect 7800 5295 8000 5300
rect 7800 5260 7825 5295
rect 7925 5260 8000 5295
rect 7800 5240 8000 5260
rect 7800 5205 7825 5240
rect 7925 5205 8000 5240
rect 7800 5200 8000 5205
rect 0 5190 60 5200
rect 190 5190 310 5200
rect 440 5190 560 5200
rect 690 5190 810 5200
rect 940 5190 1060 5200
rect 1190 5190 1310 5200
rect 1440 5190 1560 5200
rect 1690 5190 1810 5200
rect 1940 5190 2060 5200
rect 2190 5190 2310 5200
rect 2440 5190 2560 5200
rect 2690 5190 2810 5200
rect 2940 5190 3060 5200
rect 3190 5190 3310 5200
rect 3440 5190 3560 5200
rect 3690 5190 3810 5200
rect 3940 5190 4060 5200
rect 4190 5190 4310 5200
rect 4440 5190 4560 5200
rect 4690 5190 4810 5200
rect 4940 5190 5060 5200
rect 5190 5190 5310 5200
rect 5440 5190 5560 5200
rect 5690 5190 5810 5200
rect 5940 5190 6060 5200
rect 6190 5190 6310 5200
rect 6440 5190 6560 5200
rect 6690 5190 6810 5200
rect 6940 5190 7060 5200
rect 7190 5190 7310 5200
rect 7440 5190 7560 5200
rect 7690 5190 7810 5200
rect 7940 5190 8000 5200
rect 0 5175 50 5190
rect 0 5075 10 5175
rect 45 5075 50 5175
rect 0 5060 50 5075
rect 200 5175 300 5190
rect 200 5075 205 5175
rect 240 5075 260 5175
rect 295 5075 300 5175
rect 200 5060 300 5075
rect 450 5175 550 5190
rect 450 5075 455 5175
rect 490 5075 510 5175
rect 545 5075 550 5175
rect 450 5060 550 5075
rect 700 5175 800 5190
rect 700 5075 705 5175
rect 740 5075 760 5175
rect 795 5075 800 5175
rect 700 5060 800 5075
rect 950 5175 1050 5190
rect 950 5075 955 5175
rect 990 5075 1010 5175
rect 1045 5075 1050 5175
rect 950 5060 1050 5075
rect 1200 5175 1300 5190
rect 1200 5075 1205 5175
rect 1240 5075 1260 5175
rect 1295 5075 1300 5175
rect 1200 5060 1300 5075
rect 1450 5175 1550 5190
rect 1450 5075 1455 5175
rect 1490 5075 1510 5175
rect 1545 5075 1550 5175
rect 1450 5060 1550 5075
rect 1700 5175 1800 5190
rect 1700 5075 1705 5175
rect 1740 5075 1760 5175
rect 1795 5075 1800 5175
rect 1700 5060 1800 5075
rect 1950 5175 2050 5190
rect 1950 5075 1955 5175
rect 1990 5075 2010 5175
rect 2045 5075 2050 5175
rect 1950 5060 2050 5075
rect 2200 5175 2300 5190
rect 2200 5075 2205 5175
rect 2240 5075 2260 5175
rect 2295 5075 2300 5175
rect 2200 5060 2300 5075
rect 2450 5175 2550 5190
rect 2450 5075 2455 5175
rect 2490 5075 2510 5175
rect 2545 5075 2550 5175
rect 2450 5060 2550 5075
rect 2700 5175 2800 5190
rect 2700 5075 2705 5175
rect 2740 5075 2760 5175
rect 2795 5075 2800 5175
rect 2700 5060 2800 5075
rect 2950 5175 3050 5190
rect 2950 5075 2955 5175
rect 2990 5075 3010 5175
rect 3045 5075 3050 5175
rect 2950 5060 3050 5075
rect 3200 5175 3300 5190
rect 3200 5075 3205 5175
rect 3240 5075 3260 5175
rect 3295 5075 3300 5175
rect 3200 5060 3300 5075
rect 3450 5175 3550 5190
rect 3450 5075 3455 5175
rect 3490 5075 3510 5175
rect 3545 5075 3550 5175
rect 3450 5060 3550 5075
rect 3700 5175 3800 5190
rect 3700 5075 3705 5175
rect 3740 5075 3760 5175
rect 3795 5075 3800 5175
rect 3700 5060 3800 5075
rect 3950 5175 4050 5190
rect 3950 5075 3955 5175
rect 3990 5075 4010 5175
rect 4045 5075 4050 5175
rect 3950 5060 4050 5075
rect 4200 5175 4300 5190
rect 4200 5075 4205 5175
rect 4240 5075 4260 5175
rect 4295 5075 4300 5175
rect 4200 5060 4300 5075
rect 4450 5175 4550 5190
rect 4450 5075 4455 5175
rect 4490 5075 4510 5175
rect 4545 5075 4550 5175
rect 4450 5060 4550 5075
rect 4700 5175 4800 5190
rect 4700 5075 4705 5175
rect 4740 5075 4760 5175
rect 4795 5075 4800 5175
rect 4700 5060 4800 5075
rect 4950 5175 5050 5190
rect 4950 5075 4955 5175
rect 4990 5075 5010 5175
rect 5045 5075 5050 5175
rect 4950 5060 5050 5075
rect 5200 5175 5300 5190
rect 5200 5075 5205 5175
rect 5240 5075 5260 5175
rect 5295 5075 5300 5175
rect 5200 5060 5300 5075
rect 5450 5175 5550 5190
rect 5450 5075 5455 5175
rect 5490 5075 5510 5175
rect 5545 5075 5550 5175
rect 5450 5060 5550 5075
rect 5700 5175 5800 5190
rect 5700 5075 5705 5175
rect 5740 5075 5760 5175
rect 5795 5075 5800 5175
rect 5700 5060 5800 5075
rect 5950 5175 6050 5190
rect 5950 5075 5955 5175
rect 5990 5075 6010 5175
rect 6045 5075 6050 5175
rect 5950 5060 6050 5075
rect 6200 5175 6300 5190
rect 6200 5075 6205 5175
rect 6240 5075 6260 5175
rect 6295 5075 6300 5175
rect 6200 5060 6300 5075
rect 6450 5175 6550 5190
rect 6450 5075 6455 5175
rect 6490 5075 6510 5175
rect 6545 5075 6550 5175
rect 6450 5060 6550 5075
rect 6700 5175 6800 5190
rect 6700 5075 6705 5175
rect 6740 5075 6760 5175
rect 6795 5075 6800 5175
rect 6700 5060 6800 5075
rect 6950 5175 7050 5190
rect 6950 5075 6955 5175
rect 6990 5075 7010 5175
rect 7045 5075 7050 5175
rect 6950 5060 7050 5075
rect 7200 5175 7300 5190
rect 7200 5075 7205 5175
rect 7240 5075 7260 5175
rect 7295 5075 7300 5175
rect 7200 5060 7300 5075
rect 7450 5175 7550 5190
rect 7450 5075 7455 5175
rect 7490 5075 7510 5175
rect 7545 5075 7550 5175
rect 7450 5060 7550 5075
rect 7700 5175 7800 5190
rect 7700 5075 7705 5175
rect 7740 5075 7760 5175
rect 7795 5075 7800 5175
rect 7700 5060 7800 5075
rect 7950 5175 8000 5190
rect 7950 5075 7955 5175
rect 7990 5075 8000 5175
rect 7950 5060 8000 5075
rect 0 5050 60 5060
rect 190 5050 310 5060
rect 440 5050 560 5060
rect 690 5050 810 5060
rect 940 5050 1060 5060
rect 1190 5050 1310 5060
rect 1440 5050 1560 5060
rect 1690 5050 1810 5060
rect 1940 5050 2060 5060
rect 2190 5050 2310 5060
rect 2440 5050 2560 5060
rect 2690 5050 2810 5060
rect 2940 5050 3060 5060
rect 3190 5050 3310 5060
rect 3440 5050 3560 5060
rect 3690 5050 3810 5060
rect 3940 5050 4060 5060
rect 4190 5050 4310 5060
rect 4440 5050 4560 5060
rect 4690 5050 4810 5060
rect 4940 5050 5060 5060
rect 5190 5050 5310 5060
rect 5440 5050 5560 5060
rect 5690 5050 5810 5060
rect 5940 5050 6060 5060
rect 6190 5050 6310 5060
rect 6440 5050 6560 5060
rect 6690 5050 6810 5060
rect 6940 5050 7060 5060
rect 7190 5050 7310 5060
rect 7440 5050 7560 5060
rect 7690 5050 7810 5060
rect 7940 5050 8000 5060
rect 0 5045 450 5050
rect 0 5010 75 5045
rect 175 5010 325 5045
rect 425 5010 450 5045
rect 0 4990 450 5010
rect 0 4955 75 4990
rect 175 4955 325 4990
rect 425 4955 450 4990
rect 0 4950 450 4955
rect 550 5045 1450 5050
rect 550 5010 575 5045
rect 675 5010 825 5045
rect 925 5010 1075 5045
rect 1175 5010 1325 5045
rect 1425 5010 1450 5045
rect 550 4990 1450 5010
rect 550 4955 575 4990
rect 675 4955 825 4990
rect 925 4955 1075 4990
rect 1175 4955 1325 4990
rect 1425 4955 1450 4990
rect 550 4950 1450 4955
rect 1550 5045 2450 5050
rect 1550 5010 1575 5045
rect 1675 5010 1825 5045
rect 1925 5010 2075 5045
rect 2175 5010 2325 5045
rect 2425 5010 2450 5045
rect 1550 4990 2450 5010
rect 1550 4955 1575 4990
rect 1675 4955 1825 4990
rect 1925 4955 2075 4990
rect 2175 4955 2325 4990
rect 2425 4955 2450 4990
rect 1550 4950 2450 4955
rect 2550 5045 3450 5050
rect 2550 5010 2575 5045
rect 2675 5010 2825 5045
rect 2925 5010 3075 5045
rect 3175 5010 3325 5045
rect 3425 5010 3450 5045
rect 2550 4990 3450 5010
rect 2550 4955 2575 4990
rect 2675 4955 2825 4990
rect 2925 4955 3075 4990
rect 3175 4955 3325 4990
rect 3425 4955 3450 4990
rect 2550 4950 3450 4955
rect 3550 5045 4450 5050
rect 3550 5010 3575 5045
rect 3675 5010 3825 5045
rect 3925 5010 4075 5045
rect 4175 5010 4325 5045
rect 4425 5010 4450 5045
rect 3550 4990 4450 5010
rect 3550 4955 3575 4990
rect 3675 4955 3825 4990
rect 3925 4955 4075 4990
rect 4175 4955 4325 4990
rect 4425 4955 4450 4990
rect 3550 4950 4450 4955
rect 4550 5045 5450 5050
rect 4550 5010 4575 5045
rect 4675 5010 4825 5045
rect 4925 5010 5075 5045
rect 5175 5010 5325 5045
rect 5425 5010 5450 5045
rect 4550 4990 5450 5010
rect 4550 4955 4575 4990
rect 4675 4955 4825 4990
rect 4925 4955 5075 4990
rect 5175 4955 5325 4990
rect 5425 4955 5450 4990
rect 4550 4950 5450 4955
rect 5550 5045 6450 5050
rect 5550 5010 5575 5045
rect 5675 5010 5825 5045
rect 5925 5010 6075 5045
rect 6175 5010 6325 5045
rect 6425 5010 6450 5045
rect 5550 4990 6450 5010
rect 5550 4955 5575 4990
rect 5675 4955 5825 4990
rect 5925 4955 6075 4990
rect 6175 4955 6325 4990
rect 6425 4955 6450 4990
rect 5550 4950 6450 4955
rect 6550 5045 7450 5050
rect 6550 5010 6575 5045
rect 6675 5010 6825 5045
rect 6925 5010 7075 5045
rect 7175 5010 7325 5045
rect 7425 5010 7450 5045
rect 6550 4990 7450 5010
rect 6550 4955 6575 4990
rect 6675 4955 6825 4990
rect 6925 4955 7075 4990
rect 7175 4955 7325 4990
rect 7425 4955 7450 4990
rect 6550 4950 7450 4955
rect 7550 5045 8000 5050
rect 7550 5010 7575 5045
rect 7675 5010 7825 5045
rect 7925 5010 8000 5045
rect 7550 4990 8000 5010
rect 7550 4955 7575 4990
rect 7675 4955 7825 4990
rect 7925 4955 8000 4990
rect 7550 4950 8000 4955
rect 0 4940 60 4950
rect 190 4940 310 4950
rect 440 4940 560 4950
rect 690 4940 810 4950
rect 940 4940 1060 4950
rect 1190 4940 1310 4950
rect 1440 4940 1560 4950
rect 1690 4940 1810 4950
rect 1940 4940 2060 4950
rect 2190 4940 2310 4950
rect 2440 4940 2560 4950
rect 2690 4940 2810 4950
rect 2940 4940 3060 4950
rect 3190 4940 3310 4950
rect 3440 4940 3560 4950
rect 3690 4940 3810 4950
rect 3940 4940 4060 4950
rect 4190 4940 4310 4950
rect 4440 4940 4560 4950
rect 4690 4940 4810 4950
rect 4940 4940 5060 4950
rect 5190 4940 5310 4950
rect 5440 4940 5560 4950
rect 5690 4940 5810 4950
rect 5940 4940 6060 4950
rect 6190 4940 6310 4950
rect 6440 4940 6560 4950
rect 6690 4940 6810 4950
rect 6940 4940 7060 4950
rect 7190 4940 7310 4950
rect 7440 4940 7560 4950
rect 7690 4940 7810 4950
rect 7940 4940 8000 4950
rect 0 4925 50 4940
rect 0 4825 10 4925
rect 45 4825 50 4925
rect 0 4810 50 4825
rect 200 4925 300 4940
rect 200 4825 205 4925
rect 240 4825 260 4925
rect 295 4825 300 4925
rect 200 4810 300 4825
rect 450 4925 550 4940
rect 450 4825 455 4925
rect 490 4825 510 4925
rect 545 4825 550 4925
rect 450 4810 550 4825
rect 700 4925 800 4940
rect 700 4825 705 4925
rect 740 4825 760 4925
rect 795 4825 800 4925
rect 700 4810 800 4825
rect 950 4925 1050 4940
rect 950 4825 955 4925
rect 990 4825 1010 4925
rect 1045 4825 1050 4925
rect 950 4810 1050 4825
rect 1200 4925 1300 4940
rect 1200 4825 1205 4925
rect 1240 4825 1260 4925
rect 1295 4825 1300 4925
rect 1200 4810 1300 4825
rect 1450 4925 1550 4940
rect 1450 4825 1455 4925
rect 1490 4825 1510 4925
rect 1545 4825 1550 4925
rect 1450 4810 1550 4825
rect 1700 4925 1800 4940
rect 1700 4825 1705 4925
rect 1740 4825 1760 4925
rect 1795 4825 1800 4925
rect 1700 4810 1800 4825
rect 1950 4925 2050 4940
rect 1950 4825 1955 4925
rect 1990 4825 2010 4925
rect 2045 4825 2050 4925
rect 1950 4810 2050 4825
rect 2200 4925 2300 4940
rect 2200 4825 2205 4925
rect 2240 4825 2260 4925
rect 2295 4825 2300 4925
rect 2200 4810 2300 4825
rect 2450 4925 2550 4940
rect 2450 4825 2455 4925
rect 2490 4825 2510 4925
rect 2545 4825 2550 4925
rect 2450 4810 2550 4825
rect 2700 4925 2800 4940
rect 2700 4825 2705 4925
rect 2740 4825 2760 4925
rect 2795 4825 2800 4925
rect 2700 4810 2800 4825
rect 2950 4925 3050 4940
rect 2950 4825 2955 4925
rect 2990 4825 3010 4925
rect 3045 4825 3050 4925
rect 2950 4810 3050 4825
rect 3200 4925 3300 4940
rect 3200 4825 3205 4925
rect 3240 4825 3260 4925
rect 3295 4825 3300 4925
rect 3200 4810 3300 4825
rect 3450 4925 3550 4940
rect 3450 4825 3455 4925
rect 3490 4825 3510 4925
rect 3545 4825 3550 4925
rect 3450 4810 3550 4825
rect 3700 4925 3800 4940
rect 3700 4825 3705 4925
rect 3740 4825 3760 4925
rect 3795 4825 3800 4925
rect 3700 4810 3800 4825
rect 3950 4925 4050 4940
rect 3950 4825 3955 4925
rect 3990 4825 4010 4925
rect 4045 4825 4050 4925
rect 3950 4810 4050 4825
rect 4200 4925 4300 4940
rect 4200 4825 4205 4925
rect 4240 4825 4260 4925
rect 4295 4825 4300 4925
rect 4200 4810 4300 4825
rect 4450 4925 4550 4940
rect 4450 4825 4455 4925
rect 4490 4825 4510 4925
rect 4545 4825 4550 4925
rect 4450 4810 4550 4825
rect 4700 4925 4800 4940
rect 4700 4825 4705 4925
rect 4740 4825 4760 4925
rect 4795 4825 4800 4925
rect 4700 4810 4800 4825
rect 4950 4925 5050 4940
rect 4950 4825 4955 4925
rect 4990 4825 5010 4925
rect 5045 4825 5050 4925
rect 4950 4810 5050 4825
rect 5200 4925 5300 4940
rect 5200 4825 5205 4925
rect 5240 4825 5260 4925
rect 5295 4825 5300 4925
rect 5200 4810 5300 4825
rect 5450 4925 5550 4940
rect 5450 4825 5455 4925
rect 5490 4825 5510 4925
rect 5545 4825 5550 4925
rect 5450 4810 5550 4825
rect 5700 4925 5800 4940
rect 5700 4825 5705 4925
rect 5740 4825 5760 4925
rect 5795 4825 5800 4925
rect 5700 4810 5800 4825
rect 5950 4925 6050 4940
rect 5950 4825 5955 4925
rect 5990 4825 6010 4925
rect 6045 4825 6050 4925
rect 5950 4810 6050 4825
rect 6200 4925 6300 4940
rect 6200 4825 6205 4925
rect 6240 4825 6260 4925
rect 6295 4825 6300 4925
rect 6200 4810 6300 4825
rect 6450 4925 6550 4940
rect 6450 4825 6455 4925
rect 6490 4825 6510 4925
rect 6545 4825 6550 4925
rect 6450 4810 6550 4825
rect 6700 4925 6800 4940
rect 6700 4825 6705 4925
rect 6740 4825 6760 4925
rect 6795 4825 6800 4925
rect 6700 4810 6800 4825
rect 6950 4925 7050 4940
rect 6950 4825 6955 4925
rect 6990 4825 7010 4925
rect 7045 4825 7050 4925
rect 6950 4810 7050 4825
rect 7200 4925 7300 4940
rect 7200 4825 7205 4925
rect 7240 4825 7260 4925
rect 7295 4825 7300 4925
rect 7200 4810 7300 4825
rect 7450 4925 7550 4940
rect 7450 4825 7455 4925
rect 7490 4825 7510 4925
rect 7545 4825 7550 4925
rect 7450 4810 7550 4825
rect 7700 4925 7800 4940
rect 7700 4825 7705 4925
rect 7740 4825 7760 4925
rect 7795 4825 7800 4925
rect 7700 4810 7800 4825
rect 7950 4925 8000 4940
rect 7950 4825 7955 4925
rect 7990 4825 8000 4925
rect 7950 4810 8000 4825
rect 0 4800 60 4810
rect 190 4800 310 4810
rect 440 4800 560 4810
rect 690 4800 810 4810
rect 940 4800 1060 4810
rect 1190 4800 1310 4810
rect 1440 4800 1560 4810
rect 1690 4800 1810 4810
rect 1940 4800 2060 4810
rect 2190 4800 2310 4810
rect 2440 4800 2560 4810
rect 2690 4800 2810 4810
rect 2940 4800 3060 4810
rect 3190 4800 3310 4810
rect 3440 4800 3560 4810
rect 3690 4800 3810 4810
rect 3940 4800 4060 4810
rect 4190 4800 4310 4810
rect 4440 4800 4560 4810
rect 4690 4800 4810 4810
rect 4940 4800 5060 4810
rect 5190 4800 5310 4810
rect 5440 4800 5560 4810
rect 5690 4800 5810 4810
rect 5940 4800 6060 4810
rect 6190 4800 6310 4810
rect 6440 4800 6560 4810
rect 6690 4800 6810 4810
rect 6940 4800 7060 4810
rect 7190 4800 7310 4810
rect 7440 4800 7560 4810
rect 7690 4800 7810 4810
rect 7940 4800 8000 4810
rect 0 4795 200 4800
rect 0 4760 75 4795
rect 175 4760 200 4795
rect 0 4740 200 4760
rect 0 4705 75 4740
rect 175 4705 200 4740
rect 0 4700 200 4705
rect 300 4795 450 4800
rect 300 4760 325 4795
rect 425 4760 450 4795
rect 300 4740 450 4760
rect 300 4705 325 4740
rect 425 4705 450 4740
rect 300 4700 450 4705
rect 550 4795 700 4800
rect 550 4760 575 4795
rect 675 4760 700 4795
rect 550 4740 700 4760
rect 550 4705 575 4740
rect 675 4705 700 4740
rect 550 4700 700 4705
rect 800 4795 1200 4800
rect 800 4760 825 4795
rect 925 4760 1075 4795
rect 1175 4760 1200 4795
rect 800 4740 1200 4760
rect 800 4705 825 4740
rect 925 4705 1075 4740
rect 1175 4705 1200 4740
rect 800 4700 1200 4705
rect 1300 4795 1450 4800
rect 1300 4760 1325 4795
rect 1425 4760 1450 4795
rect 1300 4740 1450 4760
rect 1300 4705 1325 4740
rect 1425 4705 1450 4740
rect 1300 4700 1450 4705
rect 1550 4795 1700 4800
rect 1550 4760 1575 4795
rect 1675 4760 1700 4795
rect 1550 4740 1700 4760
rect 1550 4705 1575 4740
rect 1675 4705 1700 4740
rect 1550 4700 1700 4705
rect 1800 4795 2200 4800
rect 1800 4760 1825 4795
rect 1925 4760 2075 4795
rect 2175 4760 2200 4795
rect 1800 4740 2200 4760
rect 1800 4705 1825 4740
rect 1925 4705 2075 4740
rect 2175 4705 2200 4740
rect 1800 4700 2200 4705
rect 2300 4795 2450 4800
rect 2300 4760 2325 4795
rect 2425 4760 2450 4795
rect 2300 4740 2450 4760
rect 2300 4705 2325 4740
rect 2425 4705 2450 4740
rect 2300 4700 2450 4705
rect 2550 4795 2700 4800
rect 2550 4760 2575 4795
rect 2675 4760 2700 4795
rect 2550 4740 2700 4760
rect 2550 4705 2575 4740
rect 2675 4705 2700 4740
rect 2550 4700 2700 4705
rect 2800 4795 3200 4800
rect 2800 4760 2825 4795
rect 2925 4760 3075 4795
rect 3175 4760 3200 4795
rect 2800 4740 3200 4760
rect 2800 4705 2825 4740
rect 2925 4705 3075 4740
rect 3175 4705 3200 4740
rect 2800 4700 3200 4705
rect 3300 4795 3450 4800
rect 3300 4760 3325 4795
rect 3425 4760 3450 4795
rect 3300 4740 3450 4760
rect 3300 4705 3325 4740
rect 3425 4705 3450 4740
rect 3300 4700 3450 4705
rect 3550 4795 3700 4800
rect 3550 4760 3575 4795
rect 3675 4760 3700 4795
rect 3550 4740 3700 4760
rect 3550 4705 3575 4740
rect 3675 4705 3700 4740
rect 3550 4700 3700 4705
rect 3800 4795 4200 4800
rect 3800 4760 3825 4795
rect 3925 4760 4075 4795
rect 4175 4760 4200 4795
rect 3800 4740 4200 4760
rect 3800 4705 3825 4740
rect 3925 4705 4075 4740
rect 4175 4705 4200 4740
rect 3800 4700 4200 4705
rect 4300 4795 4450 4800
rect 4300 4760 4325 4795
rect 4425 4760 4450 4795
rect 4300 4740 4450 4760
rect 4300 4705 4325 4740
rect 4425 4705 4450 4740
rect 4300 4700 4450 4705
rect 4550 4795 4700 4800
rect 4550 4760 4575 4795
rect 4675 4760 4700 4795
rect 4550 4740 4700 4760
rect 4550 4705 4575 4740
rect 4675 4705 4700 4740
rect 4550 4700 4700 4705
rect 4800 4795 5200 4800
rect 4800 4760 4825 4795
rect 4925 4760 5075 4795
rect 5175 4760 5200 4795
rect 4800 4740 5200 4760
rect 4800 4705 4825 4740
rect 4925 4705 5075 4740
rect 5175 4705 5200 4740
rect 4800 4700 5200 4705
rect 5300 4795 5450 4800
rect 5300 4760 5325 4795
rect 5425 4760 5450 4795
rect 5300 4740 5450 4760
rect 5300 4705 5325 4740
rect 5425 4705 5450 4740
rect 5300 4700 5450 4705
rect 5550 4795 5700 4800
rect 5550 4760 5575 4795
rect 5675 4760 5700 4795
rect 5550 4740 5700 4760
rect 5550 4705 5575 4740
rect 5675 4705 5700 4740
rect 5550 4700 5700 4705
rect 5800 4795 6200 4800
rect 5800 4760 5825 4795
rect 5925 4760 6075 4795
rect 6175 4760 6200 4795
rect 5800 4740 6200 4760
rect 5800 4705 5825 4740
rect 5925 4705 6075 4740
rect 6175 4705 6200 4740
rect 5800 4700 6200 4705
rect 6300 4795 6450 4800
rect 6300 4760 6325 4795
rect 6425 4760 6450 4795
rect 6300 4740 6450 4760
rect 6300 4705 6325 4740
rect 6425 4705 6450 4740
rect 6300 4700 6450 4705
rect 6550 4795 6700 4800
rect 6550 4760 6575 4795
rect 6675 4760 6700 4795
rect 6550 4740 6700 4760
rect 6550 4705 6575 4740
rect 6675 4705 6700 4740
rect 6550 4700 6700 4705
rect 6800 4795 7200 4800
rect 6800 4760 6825 4795
rect 6925 4760 7075 4795
rect 7175 4760 7200 4795
rect 6800 4740 7200 4760
rect 6800 4705 6825 4740
rect 6925 4705 7075 4740
rect 7175 4705 7200 4740
rect 6800 4700 7200 4705
rect 7300 4795 7450 4800
rect 7300 4760 7325 4795
rect 7425 4760 7450 4795
rect 7300 4740 7450 4760
rect 7300 4705 7325 4740
rect 7425 4705 7450 4740
rect 7300 4700 7450 4705
rect 7550 4795 7700 4800
rect 7550 4760 7575 4795
rect 7675 4760 7700 4795
rect 7550 4740 7700 4760
rect 7550 4705 7575 4740
rect 7675 4705 7700 4740
rect 7550 4700 7700 4705
rect 7800 4795 8000 4800
rect 7800 4760 7825 4795
rect 7925 4760 8000 4795
rect 7800 4740 8000 4760
rect 7800 4705 7825 4740
rect 7925 4705 8000 4740
rect 7800 4700 8000 4705
rect 0 4690 60 4700
rect 190 4690 310 4700
rect 440 4690 560 4700
rect 690 4690 810 4700
rect 940 4690 1060 4700
rect 1190 4690 1310 4700
rect 1440 4690 1560 4700
rect 1690 4690 1810 4700
rect 1940 4690 2060 4700
rect 2190 4690 2310 4700
rect 2440 4690 2560 4700
rect 2690 4690 2810 4700
rect 2940 4690 3060 4700
rect 3190 4690 3310 4700
rect 3440 4690 3560 4700
rect 3690 4690 3810 4700
rect 3940 4690 4060 4700
rect 4190 4690 4310 4700
rect 4440 4690 4560 4700
rect 4690 4690 4810 4700
rect 4940 4690 5060 4700
rect 5190 4690 5310 4700
rect 5440 4690 5560 4700
rect 5690 4690 5810 4700
rect 5940 4690 6060 4700
rect 6190 4690 6310 4700
rect 6440 4690 6560 4700
rect 6690 4690 6810 4700
rect 6940 4690 7060 4700
rect 7190 4690 7310 4700
rect 7440 4690 7560 4700
rect 7690 4690 7810 4700
rect 7940 4690 8000 4700
rect 0 4675 50 4690
rect 0 4575 10 4675
rect 45 4575 50 4675
rect 0 4560 50 4575
rect 200 4675 300 4690
rect 200 4575 205 4675
rect 240 4575 260 4675
rect 295 4575 300 4675
rect 200 4560 300 4575
rect 450 4675 550 4690
rect 450 4575 455 4675
rect 490 4575 510 4675
rect 545 4575 550 4675
rect 450 4560 550 4575
rect 700 4675 800 4690
rect 700 4575 705 4675
rect 740 4575 760 4675
rect 795 4575 800 4675
rect 700 4560 800 4575
rect 950 4675 1050 4690
rect 950 4575 955 4675
rect 990 4575 1010 4675
rect 1045 4575 1050 4675
rect 950 4560 1050 4575
rect 1200 4675 1300 4690
rect 1200 4575 1205 4675
rect 1240 4575 1260 4675
rect 1295 4575 1300 4675
rect 1200 4560 1300 4575
rect 1450 4675 1550 4690
rect 1450 4575 1455 4675
rect 1490 4575 1510 4675
rect 1545 4575 1550 4675
rect 1450 4560 1550 4575
rect 1700 4675 1800 4690
rect 1700 4575 1705 4675
rect 1740 4575 1760 4675
rect 1795 4575 1800 4675
rect 1700 4560 1800 4575
rect 1950 4675 2050 4690
rect 1950 4575 1955 4675
rect 1990 4575 2010 4675
rect 2045 4575 2050 4675
rect 1950 4560 2050 4575
rect 2200 4675 2300 4690
rect 2200 4575 2205 4675
rect 2240 4575 2260 4675
rect 2295 4575 2300 4675
rect 2200 4560 2300 4575
rect 2450 4675 2550 4690
rect 2450 4575 2455 4675
rect 2490 4575 2510 4675
rect 2545 4575 2550 4675
rect 2450 4560 2550 4575
rect 2700 4675 2800 4690
rect 2700 4575 2705 4675
rect 2740 4575 2760 4675
rect 2795 4575 2800 4675
rect 2700 4560 2800 4575
rect 2950 4675 3050 4690
rect 2950 4575 2955 4675
rect 2990 4575 3010 4675
rect 3045 4575 3050 4675
rect 2950 4560 3050 4575
rect 3200 4675 3300 4690
rect 3200 4575 3205 4675
rect 3240 4575 3260 4675
rect 3295 4575 3300 4675
rect 3200 4560 3300 4575
rect 3450 4675 3550 4690
rect 3450 4575 3455 4675
rect 3490 4575 3510 4675
rect 3545 4575 3550 4675
rect 3450 4560 3550 4575
rect 3700 4675 3800 4690
rect 3700 4575 3705 4675
rect 3740 4575 3760 4675
rect 3795 4575 3800 4675
rect 3700 4560 3800 4575
rect 3950 4675 4050 4690
rect 3950 4575 3955 4675
rect 3990 4575 4010 4675
rect 4045 4575 4050 4675
rect 3950 4560 4050 4575
rect 4200 4675 4300 4690
rect 4200 4575 4205 4675
rect 4240 4575 4260 4675
rect 4295 4575 4300 4675
rect 4200 4560 4300 4575
rect 4450 4675 4550 4690
rect 4450 4575 4455 4675
rect 4490 4575 4510 4675
rect 4545 4575 4550 4675
rect 4450 4560 4550 4575
rect 4700 4675 4800 4690
rect 4700 4575 4705 4675
rect 4740 4575 4760 4675
rect 4795 4575 4800 4675
rect 4700 4560 4800 4575
rect 4950 4675 5050 4690
rect 4950 4575 4955 4675
rect 4990 4575 5010 4675
rect 5045 4575 5050 4675
rect 4950 4560 5050 4575
rect 5200 4675 5300 4690
rect 5200 4575 5205 4675
rect 5240 4575 5260 4675
rect 5295 4575 5300 4675
rect 5200 4560 5300 4575
rect 5450 4675 5550 4690
rect 5450 4575 5455 4675
rect 5490 4575 5510 4675
rect 5545 4575 5550 4675
rect 5450 4560 5550 4575
rect 5700 4675 5800 4690
rect 5700 4575 5705 4675
rect 5740 4575 5760 4675
rect 5795 4575 5800 4675
rect 5700 4560 5800 4575
rect 5950 4675 6050 4690
rect 5950 4575 5955 4675
rect 5990 4575 6010 4675
rect 6045 4575 6050 4675
rect 5950 4560 6050 4575
rect 6200 4675 6300 4690
rect 6200 4575 6205 4675
rect 6240 4575 6260 4675
rect 6295 4575 6300 4675
rect 6200 4560 6300 4575
rect 6450 4675 6550 4690
rect 6450 4575 6455 4675
rect 6490 4575 6510 4675
rect 6545 4575 6550 4675
rect 6450 4560 6550 4575
rect 6700 4675 6800 4690
rect 6700 4575 6705 4675
rect 6740 4575 6760 4675
rect 6795 4575 6800 4675
rect 6700 4560 6800 4575
rect 6950 4675 7050 4690
rect 6950 4575 6955 4675
rect 6990 4575 7010 4675
rect 7045 4575 7050 4675
rect 6950 4560 7050 4575
rect 7200 4675 7300 4690
rect 7200 4575 7205 4675
rect 7240 4575 7260 4675
rect 7295 4575 7300 4675
rect 7200 4560 7300 4575
rect 7450 4675 7550 4690
rect 7450 4575 7455 4675
rect 7490 4575 7510 4675
rect 7545 4575 7550 4675
rect 7450 4560 7550 4575
rect 7700 4675 7800 4690
rect 7700 4575 7705 4675
rect 7740 4575 7760 4675
rect 7795 4575 7800 4675
rect 7700 4560 7800 4575
rect 7950 4675 8000 4690
rect 7950 4575 7955 4675
rect 7990 4575 8000 4675
rect 7950 4560 8000 4575
rect 0 4550 60 4560
rect 190 4550 310 4560
rect 440 4550 560 4560
rect 690 4550 810 4560
rect 940 4550 1060 4560
rect 1190 4550 1310 4560
rect 1440 4550 1560 4560
rect 1690 4550 1810 4560
rect 1940 4550 2060 4560
rect 2190 4550 2310 4560
rect 2440 4550 2560 4560
rect 2690 4550 2810 4560
rect 2940 4550 3060 4560
rect 3190 4550 3310 4560
rect 3440 4550 3560 4560
rect 3690 4550 3810 4560
rect 3940 4550 4060 4560
rect 4190 4550 4310 4560
rect 4440 4550 4560 4560
rect 4690 4550 4810 4560
rect 4940 4550 5060 4560
rect 5190 4550 5310 4560
rect 5440 4550 5560 4560
rect 5690 4550 5810 4560
rect 5940 4550 6060 4560
rect 6190 4550 6310 4560
rect 6440 4550 6560 4560
rect 6690 4550 6810 4560
rect 6940 4550 7060 4560
rect 7190 4550 7310 4560
rect 7440 4550 7560 4560
rect 7690 4550 7810 4560
rect 7940 4550 8000 4560
rect 0 4545 200 4550
rect 0 4510 75 4545
rect 175 4510 200 4545
rect 0 4490 200 4510
rect 0 4455 75 4490
rect 175 4455 200 4490
rect 0 4450 200 4455
rect 300 4545 450 4550
rect 300 4510 325 4545
rect 425 4510 450 4545
rect 300 4490 450 4510
rect 300 4455 325 4490
rect 425 4455 450 4490
rect 300 4450 450 4455
rect 550 4545 700 4550
rect 550 4510 575 4545
rect 675 4510 700 4545
rect 550 4490 700 4510
rect 550 4455 575 4490
rect 675 4455 700 4490
rect 550 4450 700 4455
rect 800 4545 950 4550
rect 800 4510 825 4545
rect 925 4510 950 4545
rect 800 4490 950 4510
rect 800 4455 825 4490
rect 925 4455 950 4490
rect 800 4450 950 4455
rect 1050 4545 1200 4550
rect 1050 4510 1075 4545
rect 1175 4510 1200 4545
rect 1050 4490 1200 4510
rect 1050 4455 1075 4490
rect 1175 4455 1200 4490
rect 1050 4450 1200 4455
rect 1300 4545 1450 4550
rect 1300 4510 1325 4545
rect 1425 4510 1450 4545
rect 1300 4490 1450 4510
rect 1300 4455 1325 4490
rect 1425 4455 1450 4490
rect 1300 4450 1450 4455
rect 1550 4545 1700 4550
rect 1550 4510 1575 4545
rect 1675 4510 1700 4545
rect 1550 4490 1700 4510
rect 1550 4455 1575 4490
rect 1675 4455 1700 4490
rect 1550 4450 1700 4455
rect 1800 4545 2200 4550
rect 1800 4510 1825 4545
rect 1925 4510 2075 4545
rect 2175 4510 2200 4545
rect 1800 4490 2200 4510
rect 1800 4455 1825 4490
rect 1925 4455 2075 4490
rect 2175 4455 2200 4490
rect 1800 4450 2200 4455
rect 2300 4545 2450 4550
rect 2300 4510 2325 4545
rect 2425 4510 2450 4545
rect 2300 4490 2450 4510
rect 2300 4455 2325 4490
rect 2425 4455 2450 4490
rect 2300 4450 2450 4455
rect 2550 4545 2700 4550
rect 2550 4510 2575 4545
rect 2675 4510 2700 4545
rect 2550 4490 2700 4510
rect 2550 4455 2575 4490
rect 2675 4455 2700 4490
rect 2550 4450 2700 4455
rect 2800 4545 2950 4550
rect 2800 4510 2825 4545
rect 2925 4510 2950 4545
rect 2800 4490 2950 4510
rect 2800 4455 2825 4490
rect 2925 4455 2950 4490
rect 2800 4450 2950 4455
rect 3050 4545 3200 4550
rect 3050 4510 3075 4545
rect 3175 4510 3200 4545
rect 3050 4490 3200 4510
rect 3050 4455 3075 4490
rect 3175 4455 3200 4490
rect 3050 4450 3200 4455
rect 3300 4545 3450 4550
rect 3300 4510 3325 4545
rect 3425 4510 3450 4545
rect 3300 4490 3450 4510
rect 3300 4455 3325 4490
rect 3425 4455 3450 4490
rect 3300 4450 3450 4455
rect 3550 4545 3700 4550
rect 3550 4510 3575 4545
rect 3675 4510 3700 4545
rect 3550 4490 3700 4510
rect 3550 4455 3575 4490
rect 3675 4455 3700 4490
rect 3550 4450 3700 4455
rect 3800 4545 4200 4550
rect 3800 4510 3825 4545
rect 3925 4510 4075 4545
rect 4175 4510 4200 4545
rect 3800 4490 4200 4510
rect 3800 4455 3825 4490
rect 3925 4455 4075 4490
rect 4175 4455 4200 4490
rect 3800 4450 4200 4455
rect 4300 4545 4450 4550
rect 4300 4510 4325 4545
rect 4425 4510 4450 4545
rect 4300 4490 4450 4510
rect 4300 4455 4325 4490
rect 4425 4455 4450 4490
rect 4300 4450 4450 4455
rect 4550 4545 4700 4550
rect 4550 4510 4575 4545
rect 4675 4510 4700 4545
rect 4550 4490 4700 4510
rect 4550 4455 4575 4490
rect 4675 4455 4700 4490
rect 4550 4450 4700 4455
rect 4800 4545 4950 4550
rect 4800 4510 4825 4545
rect 4925 4510 4950 4545
rect 4800 4490 4950 4510
rect 4800 4455 4825 4490
rect 4925 4455 4950 4490
rect 4800 4450 4950 4455
rect 5050 4545 5200 4550
rect 5050 4510 5075 4545
rect 5175 4510 5200 4545
rect 5050 4490 5200 4510
rect 5050 4455 5075 4490
rect 5175 4455 5200 4490
rect 5050 4450 5200 4455
rect 5300 4545 5450 4550
rect 5300 4510 5325 4545
rect 5425 4510 5450 4545
rect 5300 4490 5450 4510
rect 5300 4455 5325 4490
rect 5425 4455 5450 4490
rect 5300 4450 5450 4455
rect 5550 4545 5700 4550
rect 5550 4510 5575 4545
rect 5675 4510 5700 4545
rect 5550 4490 5700 4510
rect 5550 4455 5575 4490
rect 5675 4455 5700 4490
rect 5550 4450 5700 4455
rect 5800 4545 6200 4550
rect 5800 4510 5825 4545
rect 5925 4510 6075 4545
rect 6175 4510 6200 4545
rect 5800 4490 6200 4510
rect 5800 4455 5825 4490
rect 5925 4455 6075 4490
rect 6175 4455 6200 4490
rect 5800 4450 6200 4455
rect 6300 4545 6450 4550
rect 6300 4510 6325 4545
rect 6425 4510 6450 4545
rect 6300 4490 6450 4510
rect 6300 4455 6325 4490
rect 6425 4455 6450 4490
rect 6300 4450 6450 4455
rect 6550 4545 6700 4550
rect 6550 4510 6575 4545
rect 6675 4510 6700 4545
rect 6550 4490 6700 4510
rect 6550 4455 6575 4490
rect 6675 4455 6700 4490
rect 6550 4450 6700 4455
rect 6800 4545 6950 4550
rect 6800 4510 6825 4545
rect 6925 4510 6950 4545
rect 6800 4490 6950 4510
rect 6800 4455 6825 4490
rect 6925 4455 6950 4490
rect 6800 4450 6950 4455
rect 7050 4545 7200 4550
rect 7050 4510 7075 4545
rect 7175 4510 7200 4545
rect 7050 4490 7200 4510
rect 7050 4455 7075 4490
rect 7175 4455 7200 4490
rect 7050 4450 7200 4455
rect 7300 4545 7450 4550
rect 7300 4510 7325 4545
rect 7425 4510 7450 4545
rect 7300 4490 7450 4510
rect 7300 4455 7325 4490
rect 7425 4455 7450 4490
rect 7300 4450 7450 4455
rect 7550 4545 7700 4550
rect 7550 4510 7575 4545
rect 7675 4510 7700 4545
rect 7550 4490 7700 4510
rect 7550 4455 7575 4490
rect 7675 4455 7700 4490
rect 7550 4450 7700 4455
rect 7800 4545 8000 4550
rect 7800 4510 7825 4545
rect 7925 4510 8000 4545
rect 7800 4490 8000 4510
rect 7800 4455 7825 4490
rect 7925 4455 8000 4490
rect 7800 4450 8000 4455
rect 0 4440 60 4450
rect 190 4440 310 4450
rect 440 4440 560 4450
rect 690 4440 810 4450
rect 940 4440 1060 4450
rect 1190 4440 1310 4450
rect 1440 4440 1560 4450
rect 1690 4440 1810 4450
rect 1940 4440 2060 4450
rect 2190 4440 2310 4450
rect 2440 4440 2560 4450
rect 2690 4440 2810 4450
rect 2940 4440 3060 4450
rect 3190 4440 3310 4450
rect 3440 4440 3560 4450
rect 3690 4440 3810 4450
rect 3940 4440 4060 4450
rect 4190 4440 4310 4450
rect 4440 4440 4560 4450
rect 4690 4440 4810 4450
rect 4940 4440 5060 4450
rect 5190 4440 5310 4450
rect 5440 4440 5560 4450
rect 5690 4440 5810 4450
rect 5940 4440 6060 4450
rect 6190 4440 6310 4450
rect 6440 4440 6560 4450
rect 6690 4440 6810 4450
rect 6940 4440 7060 4450
rect 7190 4440 7310 4450
rect 7440 4440 7560 4450
rect 7690 4440 7810 4450
rect 7940 4440 8000 4450
rect 0 4425 50 4440
rect 0 4325 10 4425
rect 45 4325 50 4425
rect 0 4310 50 4325
rect 200 4425 300 4440
rect 200 4325 205 4425
rect 240 4325 260 4425
rect 295 4325 300 4425
rect 200 4310 300 4325
rect 450 4425 550 4440
rect 450 4325 455 4425
rect 490 4325 510 4425
rect 545 4325 550 4425
rect 450 4310 550 4325
rect 700 4425 800 4440
rect 700 4325 705 4425
rect 740 4325 760 4425
rect 795 4325 800 4425
rect 700 4310 800 4325
rect 950 4425 1050 4440
rect 950 4325 955 4425
rect 990 4325 1010 4425
rect 1045 4325 1050 4425
rect 950 4310 1050 4325
rect 1200 4425 1300 4440
rect 1200 4325 1205 4425
rect 1240 4325 1260 4425
rect 1295 4325 1300 4425
rect 1200 4310 1300 4325
rect 1450 4425 1550 4440
rect 1450 4325 1455 4425
rect 1490 4325 1510 4425
rect 1545 4325 1550 4425
rect 1450 4310 1550 4325
rect 1700 4425 1800 4440
rect 1700 4325 1705 4425
rect 1740 4325 1760 4425
rect 1795 4325 1800 4425
rect 1700 4310 1800 4325
rect 1950 4425 2050 4440
rect 1950 4325 1955 4425
rect 1990 4325 2010 4425
rect 2045 4325 2050 4425
rect 1950 4310 2050 4325
rect 2200 4425 2300 4440
rect 2200 4325 2205 4425
rect 2240 4325 2260 4425
rect 2295 4325 2300 4425
rect 2200 4310 2300 4325
rect 2450 4425 2550 4440
rect 2450 4325 2455 4425
rect 2490 4325 2510 4425
rect 2545 4325 2550 4425
rect 2450 4310 2550 4325
rect 2700 4425 2800 4440
rect 2700 4325 2705 4425
rect 2740 4325 2760 4425
rect 2795 4325 2800 4425
rect 2700 4310 2800 4325
rect 2950 4425 3050 4440
rect 2950 4325 2955 4425
rect 2990 4325 3010 4425
rect 3045 4325 3050 4425
rect 2950 4310 3050 4325
rect 3200 4425 3300 4440
rect 3200 4325 3205 4425
rect 3240 4325 3260 4425
rect 3295 4325 3300 4425
rect 3200 4310 3300 4325
rect 3450 4425 3550 4440
rect 3450 4325 3455 4425
rect 3490 4325 3510 4425
rect 3545 4325 3550 4425
rect 3450 4310 3550 4325
rect 3700 4425 3800 4440
rect 3700 4325 3705 4425
rect 3740 4325 3760 4425
rect 3795 4325 3800 4425
rect 3700 4310 3800 4325
rect 3950 4425 4050 4440
rect 3950 4325 3955 4425
rect 3990 4325 4010 4425
rect 4045 4325 4050 4425
rect 3950 4310 4050 4325
rect 4200 4425 4300 4440
rect 4200 4325 4205 4425
rect 4240 4325 4260 4425
rect 4295 4325 4300 4425
rect 4200 4310 4300 4325
rect 4450 4425 4550 4440
rect 4450 4325 4455 4425
rect 4490 4325 4510 4425
rect 4545 4325 4550 4425
rect 4450 4310 4550 4325
rect 4700 4425 4800 4440
rect 4700 4325 4705 4425
rect 4740 4325 4760 4425
rect 4795 4325 4800 4425
rect 4700 4310 4800 4325
rect 4950 4425 5050 4440
rect 4950 4325 4955 4425
rect 4990 4325 5010 4425
rect 5045 4325 5050 4425
rect 4950 4310 5050 4325
rect 5200 4425 5300 4440
rect 5200 4325 5205 4425
rect 5240 4325 5260 4425
rect 5295 4325 5300 4425
rect 5200 4310 5300 4325
rect 5450 4425 5550 4440
rect 5450 4325 5455 4425
rect 5490 4325 5510 4425
rect 5545 4325 5550 4425
rect 5450 4310 5550 4325
rect 5700 4425 5800 4440
rect 5700 4325 5705 4425
rect 5740 4325 5760 4425
rect 5795 4325 5800 4425
rect 5700 4310 5800 4325
rect 5950 4425 6050 4440
rect 5950 4325 5955 4425
rect 5990 4325 6010 4425
rect 6045 4325 6050 4425
rect 5950 4310 6050 4325
rect 6200 4425 6300 4440
rect 6200 4325 6205 4425
rect 6240 4325 6260 4425
rect 6295 4325 6300 4425
rect 6200 4310 6300 4325
rect 6450 4425 6550 4440
rect 6450 4325 6455 4425
rect 6490 4325 6510 4425
rect 6545 4325 6550 4425
rect 6450 4310 6550 4325
rect 6700 4425 6800 4440
rect 6700 4325 6705 4425
rect 6740 4325 6760 4425
rect 6795 4325 6800 4425
rect 6700 4310 6800 4325
rect 6950 4425 7050 4440
rect 6950 4325 6955 4425
rect 6990 4325 7010 4425
rect 7045 4325 7050 4425
rect 6950 4310 7050 4325
rect 7200 4425 7300 4440
rect 7200 4325 7205 4425
rect 7240 4325 7260 4425
rect 7295 4325 7300 4425
rect 7200 4310 7300 4325
rect 7450 4425 7550 4440
rect 7450 4325 7455 4425
rect 7490 4325 7510 4425
rect 7545 4325 7550 4425
rect 7450 4310 7550 4325
rect 7700 4425 7800 4440
rect 7700 4325 7705 4425
rect 7740 4325 7760 4425
rect 7795 4325 7800 4425
rect 7700 4310 7800 4325
rect 7950 4425 8000 4440
rect 7950 4325 7955 4425
rect 7990 4325 8000 4425
rect 7950 4310 8000 4325
rect 0 4300 60 4310
rect 190 4300 310 4310
rect 440 4300 560 4310
rect 690 4300 810 4310
rect 940 4300 1060 4310
rect 1190 4300 1310 4310
rect 1440 4300 1560 4310
rect 1690 4300 1810 4310
rect 1940 4300 2060 4310
rect 2190 4300 2310 4310
rect 2440 4300 2560 4310
rect 2690 4300 2810 4310
rect 2940 4300 3060 4310
rect 3190 4300 3310 4310
rect 3440 4300 3560 4310
rect 3690 4300 3810 4310
rect 3940 4300 4060 4310
rect 4190 4300 4310 4310
rect 4440 4300 4560 4310
rect 4690 4300 4810 4310
rect 4940 4300 5060 4310
rect 5190 4300 5310 4310
rect 5440 4300 5560 4310
rect 5690 4300 5810 4310
rect 5940 4300 6060 4310
rect 6190 4300 6310 4310
rect 6440 4300 6560 4310
rect 6690 4300 6810 4310
rect 6940 4300 7060 4310
rect 7190 4300 7310 4310
rect 7440 4300 7560 4310
rect 7690 4300 7810 4310
rect 7940 4300 8000 4310
rect 0 4295 200 4300
rect 0 4260 75 4295
rect 175 4260 200 4295
rect 0 4240 200 4260
rect 0 4205 75 4240
rect 175 4205 200 4240
rect 0 4200 200 4205
rect 300 4295 450 4300
rect 300 4260 325 4295
rect 425 4260 450 4295
rect 300 4240 450 4260
rect 300 4205 325 4240
rect 425 4205 450 4240
rect 300 4200 450 4205
rect 550 4295 700 4300
rect 550 4260 575 4295
rect 675 4260 700 4295
rect 550 4240 700 4260
rect 550 4205 575 4240
rect 675 4205 700 4240
rect 550 4200 700 4205
rect 800 4295 1200 4300
rect 800 4260 825 4295
rect 925 4260 1075 4295
rect 1175 4260 1200 4295
rect 800 4240 1200 4260
rect 800 4205 825 4240
rect 925 4205 1075 4240
rect 1175 4205 1200 4240
rect 800 4200 1200 4205
rect 1300 4295 1450 4300
rect 1300 4260 1325 4295
rect 1425 4260 1450 4295
rect 1300 4240 1450 4260
rect 1300 4205 1325 4240
rect 1425 4205 1450 4240
rect 1300 4200 1450 4205
rect 1550 4295 1700 4300
rect 1550 4260 1575 4295
rect 1675 4260 1700 4295
rect 1550 4240 1700 4260
rect 1550 4205 1575 4240
rect 1675 4205 1700 4240
rect 1550 4200 1700 4205
rect 1800 4295 2200 4300
rect 1800 4260 1825 4295
rect 1925 4260 2075 4295
rect 2175 4260 2200 4295
rect 1800 4240 2200 4260
rect 1800 4205 1825 4240
rect 1925 4205 2075 4240
rect 2175 4205 2200 4240
rect 1800 4200 2200 4205
rect 2300 4295 2450 4300
rect 2300 4260 2325 4295
rect 2425 4260 2450 4295
rect 2300 4240 2450 4260
rect 2300 4205 2325 4240
rect 2425 4205 2450 4240
rect 2300 4200 2450 4205
rect 2550 4295 2700 4300
rect 2550 4260 2575 4295
rect 2675 4260 2700 4295
rect 2550 4240 2700 4260
rect 2550 4205 2575 4240
rect 2675 4205 2700 4240
rect 2550 4200 2700 4205
rect 2800 4295 3200 4300
rect 2800 4260 2825 4295
rect 2925 4260 3075 4295
rect 3175 4260 3200 4295
rect 2800 4240 3200 4260
rect 2800 4205 2825 4240
rect 2925 4205 3075 4240
rect 3175 4205 3200 4240
rect 2800 4200 3200 4205
rect 3300 4295 3450 4300
rect 3300 4260 3325 4295
rect 3425 4260 3450 4295
rect 3300 4240 3450 4260
rect 3300 4205 3325 4240
rect 3425 4205 3450 4240
rect 3300 4200 3450 4205
rect 3550 4295 3700 4300
rect 3550 4260 3575 4295
rect 3675 4260 3700 4295
rect 3550 4240 3700 4260
rect 3550 4205 3575 4240
rect 3675 4205 3700 4240
rect 3550 4200 3700 4205
rect 3800 4295 4200 4300
rect 3800 4260 3825 4295
rect 3925 4260 4075 4295
rect 4175 4260 4200 4295
rect 3800 4240 4200 4260
rect 3800 4205 3825 4240
rect 3925 4205 4075 4240
rect 4175 4205 4200 4240
rect 3800 4200 4200 4205
rect 4300 4295 4450 4300
rect 4300 4260 4325 4295
rect 4425 4260 4450 4295
rect 4300 4240 4450 4260
rect 4300 4205 4325 4240
rect 4425 4205 4450 4240
rect 4300 4200 4450 4205
rect 4550 4295 4700 4300
rect 4550 4260 4575 4295
rect 4675 4260 4700 4295
rect 4550 4240 4700 4260
rect 4550 4205 4575 4240
rect 4675 4205 4700 4240
rect 4550 4200 4700 4205
rect 4800 4295 5200 4300
rect 4800 4260 4825 4295
rect 4925 4260 5075 4295
rect 5175 4260 5200 4295
rect 4800 4240 5200 4260
rect 4800 4205 4825 4240
rect 4925 4205 5075 4240
rect 5175 4205 5200 4240
rect 4800 4200 5200 4205
rect 5300 4295 5450 4300
rect 5300 4260 5325 4295
rect 5425 4260 5450 4295
rect 5300 4240 5450 4260
rect 5300 4205 5325 4240
rect 5425 4205 5450 4240
rect 5300 4200 5450 4205
rect 5550 4295 5700 4300
rect 5550 4260 5575 4295
rect 5675 4260 5700 4295
rect 5550 4240 5700 4260
rect 5550 4205 5575 4240
rect 5675 4205 5700 4240
rect 5550 4200 5700 4205
rect 5800 4295 6200 4300
rect 5800 4260 5825 4295
rect 5925 4260 6075 4295
rect 6175 4260 6200 4295
rect 5800 4240 6200 4260
rect 5800 4205 5825 4240
rect 5925 4205 6075 4240
rect 6175 4205 6200 4240
rect 5800 4200 6200 4205
rect 6300 4295 6450 4300
rect 6300 4260 6325 4295
rect 6425 4260 6450 4295
rect 6300 4240 6450 4260
rect 6300 4205 6325 4240
rect 6425 4205 6450 4240
rect 6300 4200 6450 4205
rect 6550 4295 6700 4300
rect 6550 4260 6575 4295
rect 6675 4260 6700 4295
rect 6550 4240 6700 4260
rect 6550 4205 6575 4240
rect 6675 4205 6700 4240
rect 6550 4200 6700 4205
rect 6800 4295 7200 4300
rect 6800 4260 6825 4295
rect 6925 4260 7075 4295
rect 7175 4260 7200 4295
rect 6800 4240 7200 4260
rect 6800 4205 6825 4240
rect 6925 4205 7075 4240
rect 7175 4205 7200 4240
rect 6800 4200 7200 4205
rect 7300 4295 7450 4300
rect 7300 4260 7325 4295
rect 7425 4260 7450 4295
rect 7300 4240 7450 4260
rect 7300 4205 7325 4240
rect 7425 4205 7450 4240
rect 7300 4200 7450 4205
rect 7550 4295 7700 4300
rect 7550 4260 7575 4295
rect 7675 4260 7700 4295
rect 7550 4240 7700 4260
rect 7550 4205 7575 4240
rect 7675 4205 7700 4240
rect 7550 4200 7700 4205
rect 7800 4295 8000 4300
rect 7800 4260 7825 4295
rect 7925 4260 8000 4295
rect 7800 4240 8000 4260
rect 7800 4205 7825 4240
rect 7925 4205 8000 4240
rect 7800 4200 8000 4205
rect 0 4190 60 4200
rect 190 4190 310 4200
rect 440 4190 560 4200
rect 690 4190 810 4200
rect 940 4190 1060 4200
rect 1190 4190 1310 4200
rect 1440 4190 1560 4200
rect 1690 4190 1810 4200
rect 1940 4190 2060 4200
rect 2190 4190 2310 4200
rect 2440 4190 2560 4200
rect 2690 4190 2810 4200
rect 2940 4190 3060 4200
rect 3190 4190 3310 4200
rect 3440 4190 3560 4200
rect 3690 4190 3810 4200
rect 3940 4190 4060 4200
rect 4190 4190 4310 4200
rect 4440 4190 4560 4200
rect 4690 4190 4810 4200
rect 4940 4190 5060 4200
rect 5190 4190 5310 4200
rect 5440 4190 5560 4200
rect 5690 4190 5810 4200
rect 5940 4190 6060 4200
rect 6190 4190 6310 4200
rect 6440 4190 6560 4200
rect 6690 4190 6810 4200
rect 6940 4190 7060 4200
rect 7190 4190 7310 4200
rect 7440 4190 7560 4200
rect 7690 4190 7810 4200
rect 7940 4190 8000 4200
rect 0 4175 50 4190
rect 0 4075 10 4175
rect 45 4075 50 4175
rect 0 4060 50 4075
rect 200 4175 300 4190
rect 200 4075 205 4175
rect 240 4075 260 4175
rect 295 4075 300 4175
rect 200 4060 300 4075
rect 450 4175 550 4190
rect 450 4075 455 4175
rect 490 4075 510 4175
rect 545 4075 550 4175
rect 450 4060 550 4075
rect 700 4175 800 4190
rect 700 4075 705 4175
rect 740 4075 760 4175
rect 795 4075 800 4175
rect 700 4060 800 4075
rect 950 4175 1050 4190
rect 950 4075 955 4175
rect 990 4075 1010 4175
rect 1045 4075 1050 4175
rect 950 4060 1050 4075
rect 1200 4175 1300 4190
rect 1200 4075 1205 4175
rect 1240 4075 1260 4175
rect 1295 4075 1300 4175
rect 1200 4060 1300 4075
rect 1450 4175 1550 4190
rect 1450 4075 1455 4175
rect 1490 4075 1510 4175
rect 1545 4075 1550 4175
rect 1450 4060 1550 4075
rect 1700 4175 1800 4190
rect 1700 4075 1705 4175
rect 1740 4075 1760 4175
rect 1795 4075 1800 4175
rect 1700 4060 1800 4075
rect 1950 4175 2050 4190
rect 1950 4075 1955 4175
rect 1990 4075 2010 4175
rect 2045 4075 2050 4175
rect 1950 4060 2050 4075
rect 2200 4175 2300 4190
rect 2200 4075 2205 4175
rect 2240 4075 2260 4175
rect 2295 4075 2300 4175
rect 2200 4060 2300 4075
rect 2450 4175 2550 4190
rect 2450 4075 2455 4175
rect 2490 4075 2510 4175
rect 2545 4075 2550 4175
rect 2450 4060 2550 4075
rect 2700 4175 2800 4190
rect 2700 4075 2705 4175
rect 2740 4075 2760 4175
rect 2795 4075 2800 4175
rect 2700 4060 2800 4075
rect 2950 4175 3050 4190
rect 2950 4075 2955 4175
rect 2990 4075 3010 4175
rect 3045 4075 3050 4175
rect 2950 4060 3050 4075
rect 3200 4175 3300 4190
rect 3200 4075 3205 4175
rect 3240 4075 3260 4175
rect 3295 4075 3300 4175
rect 3200 4060 3300 4075
rect 3450 4175 3550 4190
rect 3450 4075 3455 4175
rect 3490 4075 3510 4175
rect 3545 4075 3550 4175
rect 3450 4060 3550 4075
rect 3700 4175 3800 4190
rect 3700 4075 3705 4175
rect 3740 4075 3760 4175
rect 3795 4075 3800 4175
rect 3700 4060 3800 4075
rect 3950 4175 4050 4190
rect 3950 4075 3955 4175
rect 3990 4075 4010 4175
rect 4045 4075 4050 4175
rect 3950 4060 4050 4075
rect 4200 4175 4300 4190
rect 4200 4075 4205 4175
rect 4240 4075 4260 4175
rect 4295 4075 4300 4175
rect 4200 4060 4300 4075
rect 4450 4175 4550 4190
rect 4450 4075 4455 4175
rect 4490 4075 4510 4175
rect 4545 4075 4550 4175
rect 4450 4060 4550 4075
rect 4700 4175 4800 4190
rect 4700 4075 4705 4175
rect 4740 4075 4760 4175
rect 4795 4075 4800 4175
rect 4700 4060 4800 4075
rect 4950 4175 5050 4190
rect 4950 4075 4955 4175
rect 4990 4075 5010 4175
rect 5045 4075 5050 4175
rect 4950 4060 5050 4075
rect 5200 4175 5300 4190
rect 5200 4075 5205 4175
rect 5240 4075 5260 4175
rect 5295 4075 5300 4175
rect 5200 4060 5300 4075
rect 5450 4175 5550 4190
rect 5450 4075 5455 4175
rect 5490 4075 5510 4175
rect 5545 4075 5550 4175
rect 5450 4060 5550 4075
rect 5700 4175 5800 4190
rect 5700 4075 5705 4175
rect 5740 4075 5760 4175
rect 5795 4075 5800 4175
rect 5700 4060 5800 4075
rect 5950 4175 6050 4190
rect 5950 4075 5955 4175
rect 5990 4075 6010 4175
rect 6045 4075 6050 4175
rect 5950 4060 6050 4075
rect 6200 4175 6300 4190
rect 6200 4075 6205 4175
rect 6240 4075 6260 4175
rect 6295 4075 6300 4175
rect 6200 4060 6300 4075
rect 6450 4175 6550 4190
rect 6450 4075 6455 4175
rect 6490 4075 6510 4175
rect 6545 4075 6550 4175
rect 6450 4060 6550 4075
rect 6700 4175 6800 4190
rect 6700 4075 6705 4175
rect 6740 4075 6760 4175
rect 6795 4075 6800 4175
rect 6700 4060 6800 4075
rect 6950 4175 7050 4190
rect 6950 4075 6955 4175
rect 6990 4075 7010 4175
rect 7045 4075 7050 4175
rect 6950 4060 7050 4075
rect 7200 4175 7300 4190
rect 7200 4075 7205 4175
rect 7240 4075 7260 4175
rect 7295 4075 7300 4175
rect 7200 4060 7300 4075
rect 7450 4175 7550 4190
rect 7450 4075 7455 4175
rect 7490 4075 7510 4175
rect 7545 4075 7550 4175
rect 7450 4060 7550 4075
rect 7700 4175 7800 4190
rect 7700 4075 7705 4175
rect 7740 4075 7760 4175
rect 7795 4075 7800 4175
rect 7700 4060 7800 4075
rect 7950 4175 8000 4190
rect 7950 4075 7955 4175
rect 7990 4075 8000 4175
rect 7950 4060 8000 4075
rect 0 4050 60 4060
rect 190 4050 310 4060
rect 440 4050 560 4060
rect 690 4050 810 4060
rect 940 4050 1060 4060
rect 1190 4050 1310 4060
rect 1440 4050 1560 4060
rect 1690 4050 1810 4060
rect 1940 4050 2060 4060
rect 2190 4050 2310 4060
rect 2440 4050 2560 4060
rect 2690 4050 2810 4060
rect 2940 4050 3060 4060
rect 3190 4050 3310 4060
rect 3440 4050 3560 4060
rect 3690 4050 3810 4060
rect 3940 4050 4060 4060
rect 4190 4050 4310 4060
rect 4440 4050 4560 4060
rect 4690 4050 4810 4060
rect 4940 4050 5060 4060
rect 5190 4050 5310 4060
rect 5440 4050 5560 4060
rect 5690 4050 5810 4060
rect 5940 4050 6060 4060
rect 6190 4050 6310 4060
rect 6440 4050 6560 4060
rect 6690 4050 6810 4060
rect 6940 4050 7060 4060
rect 7190 4050 7310 4060
rect 7440 4050 7560 4060
rect 7690 4050 7810 4060
rect 7940 4050 8000 4060
rect 0 4045 8000 4050
rect 0 4010 75 4045
rect 175 4010 325 4045
rect 425 4010 575 4045
rect 675 4010 825 4045
rect 925 4010 1075 4045
rect 1175 4010 1325 4045
rect 1425 4010 1575 4045
rect 1675 4010 1825 4045
rect 1925 4010 2075 4045
rect 2175 4010 2325 4045
rect 2425 4010 2575 4045
rect 2675 4010 2825 4045
rect 2925 4010 3075 4045
rect 3175 4010 3325 4045
rect 3425 4010 3575 4045
rect 3675 4010 3825 4045
rect 3925 4010 4075 4045
rect 4175 4010 4325 4045
rect 4425 4010 4575 4045
rect 4675 4010 4825 4045
rect 4925 4010 5075 4045
rect 5175 4010 5325 4045
rect 5425 4010 5575 4045
rect 5675 4010 5825 4045
rect 5925 4010 6075 4045
rect 6175 4010 6325 4045
rect 6425 4010 6575 4045
rect 6675 4010 6825 4045
rect 6925 4010 7075 4045
rect 7175 4010 7325 4045
rect 7425 4010 7575 4045
rect 7675 4010 7825 4045
rect 7925 4010 8000 4045
rect 0 3990 8000 4010
rect 0 3955 75 3990
rect 175 3955 325 3990
rect 425 3955 575 3990
rect 675 3955 825 3990
rect 925 3955 1075 3990
rect 1175 3955 1325 3990
rect 1425 3955 1575 3990
rect 1675 3955 1825 3990
rect 1925 3955 2075 3990
rect 2175 3955 2325 3990
rect 2425 3955 2575 3990
rect 2675 3955 2825 3990
rect 2925 3955 3075 3990
rect 3175 3955 3325 3990
rect 3425 3955 3575 3990
rect 3675 3955 3825 3990
rect 3925 3955 4075 3990
rect 4175 3955 4325 3990
rect 4425 3955 4575 3990
rect 4675 3955 4825 3990
rect 4925 3955 5075 3990
rect 5175 3955 5325 3990
rect 5425 3955 5575 3990
rect 5675 3955 5825 3990
rect 5925 3955 6075 3990
rect 6175 3955 6325 3990
rect 6425 3955 6575 3990
rect 6675 3955 6825 3990
rect 6925 3955 7075 3990
rect 7175 3955 7325 3990
rect 7425 3955 7575 3990
rect 7675 3955 7825 3990
rect 7925 3955 8000 3990
rect 0 3950 8000 3955
rect 0 3940 60 3950
rect 190 3940 310 3950
rect 440 3940 560 3950
rect 690 3940 810 3950
rect 940 3940 1060 3950
rect 1190 3940 1310 3950
rect 1440 3940 1560 3950
rect 1690 3940 1810 3950
rect 1940 3940 2060 3950
rect 2190 3940 2310 3950
rect 2440 3940 2560 3950
rect 2690 3940 2810 3950
rect 2940 3940 3060 3950
rect 3190 3940 3310 3950
rect 3440 3940 3560 3950
rect 3690 3940 3810 3950
rect 3940 3940 4060 3950
rect 4190 3940 4310 3950
rect 4440 3940 4560 3950
rect 4690 3940 4810 3950
rect 4940 3940 5060 3950
rect 5190 3940 5310 3950
rect 5440 3940 5560 3950
rect 5690 3940 5810 3950
rect 5940 3940 6060 3950
rect 6190 3940 6310 3950
rect 6440 3940 6560 3950
rect 6690 3940 6810 3950
rect 6940 3940 7060 3950
rect 7190 3940 7310 3950
rect 7440 3940 7560 3950
rect 7690 3940 7810 3950
rect 7940 3940 8000 3950
rect 0 3925 50 3940
rect 0 3825 10 3925
rect 45 3825 50 3925
rect 0 3810 50 3825
rect 200 3925 300 3940
rect 200 3825 205 3925
rect 240 3825 260 3925
rect 295 3825 300 3925
rect 200 3810 300 3825
rect 450 3925 550 3940
rect 450 3825 455 3925
rect 490 3825 510 3925
rect 545 3825 550 3925
rect 450 3810 550 3825
rect 700 3925 800 3940
rect 700 3825 705 3925
rect 740 3825 760 3925
rect 795 3825 800 3925
rect 700 3810 800 3825
rect 950 3925 1050 3940
rect 950 3825 955 3925
rect 990 3825 1010 3925
rect 1045 3825 1050 3925
rect 950 3810 1050 3825
rect 1200 3925 1300 3940
rect 1200 3825 1205 3925
rect 1240 3825 1260 3925
rect 1295 3825 1300 3925
rect 1200 3810 1300 3825
rect 1450 3925 1550 3940
rect 1450 3825 1455 3925
rect 1490 3825 1510 3925
rect 1545 3825 1550 3925
rect 1450 3810 1550 3825
rect 1700 3925 1800 3940
rect 1700 3825 1705 3925
rect 1740 3825 1760 3925
rect 1795 3825 1800 3925
rect 1700 3810 1800 3825
rect 1950 3925 2050 3940
rect 1950 3825 1955 3925
rect 1990 3825 2010 3925
rect 2045 3825 2050 3925
rect 1950 3810 2050 3825
rect 2200 3925 2300 3940
rect 2200 3825 2205 3925
rect 2240 3825 2260 3925
rect 2295 3825 2300 3925
rect 2200 3810 2300 3825
rect 2450 3925 2550 3940
rect 2450 3825 2455 3925
rect 2490 3825 2510 3925
rect 2545 3825 2550 3925
rect 2450 3810 2550 3825
rect 2700 3925 2800 3940
rect 2700 3825 2705 3925
rect 2740 3825 2760 3925
rect 2795 3825 2800 3925
rect 2700 3810 2800 3825
rect 2950 3925 3050 3940
rect 2950 3825 2955 3925
rect 2990 3825 3010 3925
rect 3045 3825 3050 3925
rect 2950 3810 3050 3825
rect 3200 3925 3300 3940
rect 3200 3825 3205 3925
rect 3240 3825 3260 3925
rect 3295 3825 3300 3925
rect 3200 3810 3300 3825
rect 3450 3925 3550 3940
rect 3450 3825 3455 3925
rect 3490 3825 3510 3925
rect 3545 3825 3550 3925
rect 3450 3810 3550 3825
rect 3700 3925 3800 3940
rect 3700 3825 3705 3925
rect 3740 3825 3760 3925
rect 3795 3825 3800 3925
rect 3700 3810 3800 3825
rect 3950 3925 4050 3940
rect 3950 3825 3955 3925
rect 3990 3825 4010 3925
rect 4045 3825 4050 3925
rect 3950 3810 4050 3825
rect 4200 3925 4300 3940
rect 4200 3825 4205 3925
rect 4240 3825 4260 3925
rect 4295 3825 4300 3925
rect 4200 3810 4300 3825
rect 4450 3925 4550 3940
rect 4450 3825 4455 3925
rect 4490 3825 4510 3925
rect 4545 3825 4550 3925
rect 4450 3810 4550 3825
rect 4700 3925 4800 3940
rect 4700 3825 4705 3925
rect 4740 3825 4760 3925
rect 4795 3825 4800 3925
rect 4700 3810 4800 3825
rect 4950 3925 5050 3940
rect 4950 3825 4955 3925
rect 4990 3825 5010 3925
rect 5045 3825 5050 3925
rect 4950 3810 5050 3825
rect 5200 3925 5300 3940
rect 5200 3825 5205 3925
rect 5240 3825 5260 3925
rect 5295 3825 5300 3925
rect 5200 3810 5300 3825
rect 5450 3925 5550 3940
rect 5450 3825 5455 3925
rect 5490 3825 5510 3925
rect 5545 3825 5550 3925
rect 5450 3810 5550 3825
rect 5700 3925 5800 3940
rect 5700 3825 5705 3925
rect 5740 3825 5760 3925
rect 5795 3825 5800 3925
rect 5700 3810 5800 3825
rect 5950 3925 6050 3940
rect 5950 3825 5955 3925
rect 5990 3825 6010 3925
rect 6045 3825 6050 3925
rect 5950 3810 6050 3825
rect 6200 3925 6300 3940
rect 6200 3825 6205 3925
rect 6240 3825 6260 3925
rect 6295 3825 6300 3925
rect 6200 3810 6300 3825
rect 6450 3925 6550 3940
rect 6450 3825 6455 3925
rect 6490 3825 6510 3925
rect 6545 3825 6550 3925
rect 6450 3810 6550 3825
rect 6700 3925 6800 3940
rect 6700 3825 6705 3925
rect 6740 3825 6760 3925
rect 6795 3825 6800 3925
rect 6700 3810 6800 3825
rect 6950 3925 7050 3940
rect 6950 3825 6955 3925
rect 6990 3825 7010 3925
rect 7045 3825 7050 3925
rect 6950 3810 7050 3825
rect 7200 3925 7300 3940
rect 7200 3825 7205 3925
rect 7240 3825 7260 3925
rect 7295 3825 7300 3925
rect 7200 3810 7300 3825
rect 7450 3925 7550 3940
rect 7450 3825 7455 3925
rect 7490 3825 7510 3925
rect 7545 3825 7550 3925
rect 7450 3810 7550 3825
rect 7700 3925 7800 3940
rect 7700 3825 7705 3925
rect 7740 3825 7760 3925
rect 7795 3825 7800 3925
rect 7700 3810 7800 3825
rect 7950 3925 8000 3940
rect 7950 3825 7955 3925
rect 7990 3825 8000 3925
rect 7950 3810 8000 3825
rect 0 3800 60 3810
rect 190 3800 310 3810
rect 440 3800 560 3810
rect 690 3800 810 3810
rect 940 3800 1060 3810
rect 1190 3800 1310 3810
rect 1440 3800 1560 3810
rect 1690 3800 1810 3810
rect 1940 3800 2060 3810
rect 2190 3800 2310 3810
rect 2440 3800 2560 3810
rect 2690 3800 2810 3810
rect 2940 3800 3060 3810
rect 3190 3800 3310 3810
rect 3440 3800 3560 3810
rect 3690 3800 3810 3810
rect 3940 3800 4060 3810
rect 4190 3800 4310 3810
rect 4440 3800 4560 3810
rect 4690 3800 4810 3810
rect 4940 3800 5060 3810
rect 5190 3800 5310 3810
rect 5440 3800 5560 3810
rect 5690 3800 5810 3810
rect 5940 3800 6060 3810
rect 6190 3800 6310 3810
rect 6440 3800 6560 3810
rect 6690 3800 6810 3810
rect 6940 3800 7060 3810
rect 7190 3800 7310 3810
rect 7440 3800 7560 3810
rect 7690 3800 7810 3810
rect 7940 3800 8000 3810
rect 0 3795 200 3800
rect 0 3760 75 3795
rect 175 3760 200 3795
rect 0 3740 200 3760
rect 0 3705 75 3740
rect 175 3705 200 3740
rect 0 3700 200 3705
rect 300 3795 450 3800
rect 300 3760 325 3795
rect 425 3760 450 3795
rect 300 3740 450 3760
rect 300 3705 325 3740
rect 425 3705 450 3740
rect 300 3700 450 3705
rect 550 3795 700 3800
rect 550 3760 575 3795
rect 675 3760 700 3795
rect 550 3740 700 3760
rect 550 3705 575 3740
rect 675 3705 700 3740
rect 550 3700 700 3705
rect 800 3795 1200 3800
rect 800 3760 825 3795
rect 925 3760 1075 3795
rect 1175 3760 1200 3795
rect 800 3740 1200 3760
rect 800 3705 825 3740
rect 925 3705 1075 3740
rect 1175 3705 1200 3740
rect 800 3700 1200 3705
rect 1300 3795 1450 3800
rect 1300 3760 1325 3795
rect 1425 3760 1450 3795
rect 1300 3740 1450 3760
rect 1300 3705 1325 3740
rect 1425 3705 1450 3740
rect 1300 3700 1450 3705
rect 1550 3795 1700 3800
rect 1550 3760 1575 3795
rect 1675 3760 1700 3795
rect 1550 3740 1700 3760
rect 1550 3705 1575 3740
rect 1675 3705 1700 3740
rect 1550 3700 1700 3705
rect 1800 3795 2200 3800
rect 1800 3760 1825 3795
rect 1925 3760 2075 3795
rect 2175 3760 2200 3795
rect 1800 3740 2200 3760
rect 1800 3705 1825 3740
rect 1925 3705 2075 3740
rect 2175 3705 2200 3740
rect 1800 3700 2200 3705
rect 2300 3795 2450 3800
rect 2300 3760 2325 3795
rect 2425 3760 2450 3795
rect 2300 3740 2450 3760
rect 2300 3705 2325 3740
rect 2425 3705 2450 3740
rect 2300 3700 2450 3705
rect 2550 3795 2700 3800
rect 2550 3760 2575 3795
rect 2675 3760 2700 3795
rect 2550 3740 2700 3760
rect 2550 3705 2575 3740
rect 2675 3705 2700 3740
rect 2550 3700 2700 3705
rect 2800 3795 3200 3800
rect 2800 3760 2825 3795
rect 2925 3760 3075 3795
rect 3175 3760 3200 3795
rect 2800 3740 3200 3760
rect 2800 3705 2825 3740
rect 2925 3705 3075 3740
rect 3175 3705 3200 3740
rect 2800 3700 3200 3705
rect 3300 3795 3450 3800
rect 3300 3760 3325 3795
rect 3425 3760 3450 3795
rect 3300 3740 3450 3760
rect 3300 3705 3325 3740
rect 3425 3705 3450 3740
rect 3300 3700 3450 3705
rect 3550 3795 3700 3800
rect 3550 3760 3575 3795
rect 3675 3760 3700 3795
rect 3550 3740 3700 3760
rect 3550 3705 3575 3740
rect 3675 3705 3700 3740
rect 3550 3700 3700 3705
rect 3800 3795 4200 3800
rect 3800 3760 3825 3795
rect 3925 3760 4075 3795
rect 4175 3760 4200 3795
rect 3800 3740 4200 3760
rect 3800 3705 3825 3740
rect 3925 3705 4075 3740
rect 4175 3705 4200 3740
rect 3800 3700 4200 3705
rect 4300 3795 4450 3800
rect 4300 3760 4325 3795
rect 4425 3760 4450 3795
rect 4300 3740 4450 3760
rect 4300 3705 4325 3740
rect 4425 3705 4450 3740
rect 4300 3700 4450 3705
rect 4550 3795 4700 3800
rect 4550 3760 4575 3795
rect 4675 3760 4700 3795
rect 4550 3740 4700 3760
rect 4550 3705 4575 3740
rect 4675 3705 4700 3740
rect 4550 3700 4700 3705
rect 4800 3795 5200 3800
rect 4800 3760 4825 3795
rect 4925 3760 5075 3795
rect 5175 3760 5200 3795
rect 4800 3740 5200 3760
rect 4800 3705 4825 3740
rect 4925 3705 5075 3740
rect 5175 3705 5200 3740
rect 4800 3700 5200 3705
rect 5300 3795 5450 3800
rect 5300 3760 5325 3795
rect 5425 3760 5450 3795
rect 5300 3740 5450 3760
rect 5300 3705 5325 3740
rect 5425 3705 5450 3740
rect 5300 3700 5450 3705
rect 5550 3795 5700 3800
rect 5550 3760 5575 3795
rect 5675 3760 5700 3795
rect 5550 3740 5700 3760
rect 5550 3705 5575 3740
rect 5675 3705 5700 3740
rect 5550 3700 5700 3705
rect 5800 3795 6200 3800
rect 5800 3760 5825 3795
rect 5925 3760 6075 3795
rect 6175 3760 6200 3795
rect 5800 3740 6200 3760
rect 5800 3705 5825 3740
rect 5925 3705 6075 3740
rect 6175 3705 6200 3740
rect 5800 3700 6200 3705
rect 6300 3795 6450 3800
rect 6300 3760 6325 3795
rect 6425 3760 6450 3795
rect 6300 3740 6450 3760
rect 6300 3705 6325 3740
rect 6425 3705 6450 3740
rect 6300 3700 6450 3705
rect 6550 3795 6700 3800
rect 6550 3760 6575 3795
rect 6675 3760 6700 3795
rect 6550 3740 6700 3760
rect 6550 3705 6575 3740
rect 6675 3705 6700 3740
rect 6550 3700 6700 3705
rect 6800 3795 7200 3800
rect 6800 3760 6825 3795
rect 6925 3760 7075 3795
rect 7175 3760 7200 3795
rect 6800 3740 7200 3760
rect 6800 3705 6825 3740
rect 6925 3705 7075 3740
rect 7175 3705 7200 3740
rect 6800 3700 7200 3705
rect 7300 3795 7450 3800
rect 7300 3760 7325 3795
rect 7425 3760 7450 3795
rect 7300 3740 7450 3760
rect 7300 3705 7325 3740
rect 7425 3705 7450 3740
rect 7300 3700 7450 3705
rect 7550 3795 7700 3800
rect 7550 3760 7575 3795
rect 7675 3760 7700 3795
rect 7550 3740 7700 3760
rect 7550 3705 7575 3740
rect 7675 3705 7700 3740
rect 7550 3700 7700 3705
rect 7800 3795 8000 3800
rect 7800 3760 7825 3795
rect 7925 3760 8000 3795
rect 7800 3740 8000 3760
rect 7800 3705 7825 3740
rect 7925 3705 8000 3740
rect 7800 3700 8000 3705
rect 0 3690 60 3700
rect 190 3690 310 3700
rect 440 3690 560 3700
rect 690 3690 810 3700
rect 940 3690 1060 3700
rect 1190 3690 1310 3700
rect 1440 3690 1560 3700
rect 1690 3690 1810 3700
rect 1940 3690 2060 3700
rect 2190 3690 2310 3700
rect 2440 3690 2560 3700
rect 2690 3690 2810 3700
rect 2940 3690 3060 3700
rect 3190 3690 3310 3700
rect 3440 3690 3560 3700
rect 3690 3690 3810 3700
rect 3940 3690 4060 3700
rect 4190 3690 4310 3700
rect 4440 3690 4560 3700
rect 4690 3690 4810 3700
rect 4940 3690 5060 3700
rect 5190 3690 5310 3700
rect 5440 3690 5560 3700
rect 5690 3690 5810 3700
rect 5940 3690 6060 3700
rect 6190 3690 6310 3700
rect 6440 3690 6560 3700
rect 6690 3690 6810 3700
rect 6940 3690 7060 3700
rect 7190 3690 7310 3700
rect 7440 3690 7560 3700
rect 7690 3690 7810 3700
rect 7940 3690 8000 3700
rect 0 3675 50 3690
rect 0 3575 10 3675
rect 45 3575 50 3675
rect 0 3560 50 3575
rect 200 3675 300 3690
rect 200 3575 205 3675
rect 240 3575 260 3675
rect 295 3575 300 3675
rect 200 3560 300 3575
rect 450 3675 550 3690
rect 450 3575 455 3675
rect 490 3575 510 3675
rect 545 3575 550 3675
rect 450 3560 550 3575
rect 700 3675 800 3690
rect 700 3575 705 3675
rect 740 3575 760 3675
rect 795 3575 800 3675
rect 700 3560 800 3575
rect 950 3675 1050 3690
rect 950 3575 955 3675
rect 990 3575 1010 3675
rect 1045 3575 1050 3675
rect 950 3560 1050 3575
rect 1200 3675 1300 3690
rect 1200 3575 1205 3675
rect 1240 3575 1260 3675
rect 1295 3575 1300 3675
rect 1200 3560 1300 3575
rect 1450 3675 1550 3690
rect 1450 3575 1455 3675
rect 1490 3575 1510 3675
rect 1545 3575 1550 3675
rect 1450 3560 1550 3575
rect 1700 3675 1800 3690
rect 1700 3575 1705 3675
rect 1740 3575 1760 3675
rect 1795 3575 1800 3675
rect 1700 3560 1800 3575
rect 1950 3675 2050 3690
rect 1950 3575 1955 3675
rect 1990 3575 2010 3675
rect 2045 3575 2050 3675
rect 1950 3560 2050 3575
rect 2200 3675 2300 3690
rect 2200 3575 2205 3675
rect 2240 3575 2260 3675
rect 2295 3575 2300 3675
rect 2200 3560 2300 3575
rect 2450 3675 2550 3690
rect 2450 3575 2455 3675
rect 2490 3575 2510 3675
rect 2545 3575 2550 3675
rect 2450 3560 2550 3575
rect 2700 3675 2800 3690
rect 2700 3575 2705 3675
rect 2740 3575 2760 3675
rect 2795 3575 2800 3675
rect 2700 3560 2800 3575
rect 2950 3675 3050 3690
rect 2950 3575 2955 3675
rect 2990 3575 3010 3675
rect 3045 3575 3050 3675
rect 2950 3560 3050 3575
rect 3200 3675 3300 3690
rect 3200 3575 3205 3675
rect 3240 3575 3260 3675
rect 3295 3575 3300 3675
rect 3200 3560 3300 3575
rect 3450 3675 3550 3690
rect 3450 3575 3455 3675
rect 3490 3575 3510 3675
rect 3545 3575 3550 3675
rect 3450 3560 3550 3575
rect 3700 3675 3800 3690
rect 3700 3575 3705 3675
rect 3740 3575 3760 3675
rect 3795 3575 3800 3675
rect 3700 3560 3800 3575
rect 3950 3675 4050 3690
rect 3950 3575 3955 3675
rect 3990 3575 4010 3675
rect 4045 3575 4050 3675
rect 3950 3560 4050 3575
rect 4200 3675 4300 3690
rect 4200 3575 4205 3675
rect 4240 3575 4260 3675
rect 4295 3575 4300 3675
rect 4200 3560 4300 3575
rect 4450 3675 4550 3690
rect 4450 3575 4455 3675
rect 4490 3575 4510 3675
rect 4545 3575 4550 3675
rect 4450 3560 4550 3575
rect 4700 3675 4800 3690
rect 4700 3575 4705 3675
rect 4740 3575 4760 3675
rect 4795 3575 4800 3675
rect 4700 3560 4800 3575
rect 4950 3675 5050 3690
rect 4950 3575 4955 3675
rect 4990 3575 5010 3675
rect 5045 3575 5050 3675
rect 4950 3560 5050 3575
rect 5200 3675 5300 3690
rect 5200 3575 5205 3675
rect 5240 3575 5260 3675
rect 5295 3575 5300 3675
rect 5200 3560 5300 3575
rect 5450 3675 5550 3690
rect 5450 3575 5455 3675
rect 5490 3575 5510 3675
rect 5545 3575 5550 3675
rect 5450 3560 5550 3575
rect 5700 3675 5800 3690
rect 5700 3575 5705 3675
rect 5740 3575 5760 3675
rect 5795 3575 5800 3675
rect 5700 3560 5800 3575
rect 5950 3675 6050 3690
rect 5950 3575 5955 3675
rect 5990 3575 6010 3675
rect 6045 3575 6050 3675
rect 5950 3560 6050 3575
rect 6200 3675 6300 3690
rect 6200 3575 6205 3675
rect 6240 3575 6260 3675
rect 6295 3575 6300 3675
rect 6200 3560 6300 3575
rect 6450 3675 6550 3690
rect 6450 3575 6455 3675
rect 6490 3575 6510 3675
rect 6545 3575 6550 3675
rect 6450 3560 6550 3575
rect 6700 3675 6800 3690
rect 6700 3575 6705 3675
rect 6740 3575 6760 3675
rect 6795 3575 6800 3675
rect 6700 3560 6800 3575
rect 6950 3675 7050 3690
rect 6950 3575 6955 3675
rect 6990 3575 7010 3675
rect 7045 3575 7050 3675
rect 6950 3560 7050 3575
rect 7200 3675 7300 3690
rect 7200 3575 7205 3675
rect 7240 3575 7260 3675
rect 7295 3575 7300 3675
rect 7200 3560 7300 3575
rect 7450 3675 7550 3690
rect 7450 3575 7455 3675
rect 7490 3575 7510 3675
rect 7545 3575 7550 3675
rect 7450 3560 7550 3575
rect 7700 3675 7800 3690
rect 7700 3575 7705 3675
rect 7740 3575 7760 3675
rect 7795 3575 7800 3675
rect 7700 3560 7800 3575
rect 7950 3675 8000 3690
rect 7950 3575 7955 3675
rect 7990 3575 8000 3675
rect 7950 3560 8000 3575
rect 0 3550 60 3560
rect 190 3550 310 3560
rect 440 3550 560 3560
rect 690 3550 810 3560
rect 940 3550 1060 3560
rect 1190 3550 1310 3560
rect 1440 3550 1560 3560
rect 1690 3550 1810 3560
rect 1940 3550 2060 3560
rect 2190 3550 2310 3560
rect 2440 3550 2560 3560
rect 2690 3550 2810 3560
rect 2940 3550 3060 3560
rect 3190 3550 3310 3560
rect 3440 3550 3560 3560
rect 3690 3550 3810 3560
rect 3940 3550 4060 3560
rect 4190 3550 4310 3560
rect 4440 3550 4560 3560
rect 4690 3550 4810 3560
rect 4940 3550 5060 3560
rect 5190 3550 5310 3560
rect 5440 3550 5560 3560
rect 5690 3550 5810 3560
rect 5940 3550 6060 3560
rect 6190 3550 6310 3560
rect 6440 3550 6560 3560
rect 6690 3550 6810 3560
rect 6940 3550 7060 3560
rect 7190 3550 7310 3560
rect 7440 3550 7560 3560
rect 7690 3550 7810 3560
rect 7940 3550 8000 3560
rect 0 3545 200 3550
rect 0 3510 75 3545
rect 175 3510 200 3545
rect 0 3490 200 3510
rect 0 3455 75 3490
rect 175 3455 200 3490
rect 0 3450 200 3455
rect 300 3545 450 3550
rect 300 3510 325 3545
rect 425 3510 450 3545
rect 300 3490 450 3510
rect 300 3455 325 3490
rect 425 3455 450 3490
rect 300 3450 450 3455
rect 550 3545 700 3550
rect 550 3510 575 3545
rect 675 3510 700 3545
rect 550 3490 700 3510
rect 550 3455 575 3490
rect 675 3455 700 3490
rect 550 3450 700 3455
rect 800 3545 950 3550
rect 800 3510 825 3545
rect 925 3510 950 3545
rect 800 3490 950 3510
rect 800 3455 825 3490
rect 925 3455 950 3490
rect 800 3450 950 3455
rect 1050 3545 1200 3550
rect 1050 3510 1075 3545
rect 1175 3510 1200 3545
rect 1050 3490 1200 3510
rect 1050 3455 1075 3490
rect 1175 3455 1200 3490
rect 1050 3450 1200 3455
rect 1300 3545 1450 3550
rect 1300 3510 1325 3545
rect 1425 3510 1450 3545
rect 1300 3490 1450 3510
rect 1300 3455 1325 3490
rect 1425 3455 1450 3490
rect 1300 3450 1450 3455
rect 1550 3545 1700 3550
rect 1550 3510 1575 3545
rect 1675 3510 1700 3545
rect 1550 3490 1700 3510
rect 1550 3455 1575 3490
rect 1675 3455 1700 3490
rect 1550 3450 1700 3455
rect 1800 3545 2200 3550
rect 1800 3510 1825 3545
rect 1925 3510 2075 3545
rect 2175 3510 2200 3545
rect 1800 3490 2200 3510
rect 1800 3455 1825 3490
rect 1925 3455 2075 3490
rect 2175 3455 2200 3490
rect 1800 3450 2200 3455
rect 2300 3545 2450 3550
rect 2300 3510 2325 3545
rect 2425 3510 2450 3545
rect 2300 3490 2450 3510
rect 2300 3455 2325 3490
rect 2425 3455 2450 3490
rect 2300 3450 2450 3455
rect 2550 3545 2700 3550
rect 2550 3510 2575 3545
rect 2675 3510 2700 3545
rect 2550 3490 2700 3510
rect 2550 3455 2575 3490
rect 2675 3455 2700 3490
rect 2550 3450 2700 3455
rect 2800 3545 2950 3550
rect 2800 3510 2825 3545
rect 2925 3510 2950 3545
rect 2800 3490 2950 3510
rect 2800 3455 2825 3490
rect 2925 3455 2950 3490
rect 2800 3450 2950 3455
rect 3050 3545 3200 3550
rect 3050 3510 3075 3545
rect 3175 3510 3200 3545
rect 3050 3490 3200 3510
rect 3050 3455 3075 3490
rect 3175 3455 3200 3490
rect 3050 3450 3200 3455
rect 3300 3545 3450 3550
rect 3300 3510 3325 3545
rect 3425 3510 3450 3545
rect 3300 3490 3450 3510
rect 3300 3455 3325 3490
rect 3425 3455 3450 3490
rect 3300 3450 3450 3455
rect 3550 3545 3700 3550
rect 3550 3510 3575 3545
rect 3675 3510 3700 3545
rect 3550 3490 3700 3510
rect 3550 3455 3575 3490
rect 3675 3455 3700 3490
rect 3550 3450 3700 3455
rect 3800 3545 4200 3550
rect 3800 3510 3825 3545
rect 3925 3510 4075 3545
rect 4175 3510 4200 3545
rect 3800 3490 4200 3510
rect 3800 3455 3825 3490
rect 3925 3455 4075 3490
rect 4175 3455 4200 3490
rect 3800 3450 4200 3455
rect 4300 3545 4450 3550
rect 4300 3510 4325 3545
rect 4425 3510 4450 3545
rect 4300 3490 4450 3510
rect 4300 3455 4325 3490
rect 4425 3455 4450 3490
rect 4300 3450 4450 3455
rect 4550 3545 4700 3550
rect 4550 3510 4575 3545
rect 4675 3510 4700 3545
rect 4550 3490 4700 3510
rect 4550 3455 4575 3490
rect 4675 3455 4700 3490
rect 4550 3450 4700 3455
rect 4800 3545 4950 3550
rect 4800 3510 4825 3545
rect 4925 3510 4950 3545
rect 4800 3490 4950 3510
rect 4800 3455 4825 3490
rect 4925 3455 4950 3490
rect 4800 3450 4950 3455
rect 5050 3545 5200 3550
rect 5050 3510 5075 3545
rect 5175 3510 5200 3545
rect 5050 3490 5200 3510
rect 5050 3455 5075 3490
rect 5175 3455 5200 3490
rect 5050 3450 5200 3455
rect 5300 3545 5450 3550
rect 5300 3510 5325 3545
rect 5425 3510 5450 3545
rect 5300 3490 5450 3510
rect 5300 3455 5325 3490
rect 5425 3455 5450 3490
rect 5300 3450 5450 3455
rect 5550 3545 5700 3550
rect 5550 3510 5575 3545
rect 5675 3510 5700 3545
rect 5550 3490 5700 3510
rect 5550 3455 5575 3490
rect 5675 3455 5700 3490
rect 5550 3450 5700 3455
rect 5800 3545 6200 3550
rect 5800 3510 5825 3545
rect 5925 3510 6075 3545
rect 6175 3510 6200 3545
rect 5800 3490 6200 3510
rect 5800 3455 5825 3490
rect 5925 3455 6075 3490
rect 6175 3455 6200 3490
rect 5800 3450 6200 3455
rect 6300 3545 6450 3550
rect 6300 3510 6325 3545
rect 6425 3510 6450 3545
rect 6300 3490 6450 3510
rect 6300 3455 6325 3490
rect 6425 3455 6450 3490
rect 6300 3450 6450 3455
rect 6550 3545 6700 3550
rect 6550 3510 6575 3545
rect 6675 3510 6700 3545
rect 6550 3490 6700 3510
rect 6550 3455 6575 3490
rect 6675 3455 6700 3490
rect 6550 3450 6700 3455
rect 6800 3545 6950 3550
rect 6800 3510 6825 3545
rect 6925 3510 6950 3545
rect 6800 3490 6950 3510
rect 6800 3455 6825 3490
rect 6925 3455 6950 3490
rect 6800 3450 6950 3455
rect 7050 3545 7200 3550
rect 7050 3510 7075 3545
rect 7175 3510 7200 3545
rect 7050 3490 7200 3510
rect 7050 3455 7075 3490
rect 7175 3455 7200 3490
rect 7050 3450 7200 3455
rect 7300 3545 7450 3550
rect 7300 3510 7325 3545
rect 7425 3510 7450 3545
rect 7300 3490 7450 3510
rect 7300 3455 7325 3490
rect 7425 3455 7450 3490
rect 7300 3450 7450 3455
rect 7550 3545 7700 3550
rect 7550 3510 7575 3545
rect 7675 3510 7700 3545
rect 7550 3490 7700 3510
rect 7550 3455 7575 3490
rect 7675 3455 7700 3490
rect 7550 3450 7700 3455
rect 7800 3545 8000 3550
rect 7800 3510 7825 3545
rect 7925 3510 8000 3545
rect 7800 3490 8000 3510
rect 7800 3455 7825 3490
rect 7925 3455 8000 3490
rect 7800 3450 8000 3455
rect 0 3440 60 3450
rect 190 3440 310 3450
rect 440 3440 560 3450
rect 690 3440 810 3450
rect 940 3440 1060 3450
rect 1190 3440 1310 3450
rect 1440 3440 1560 3450
rect 1690 3440 1810 3450
rect 1940 3440 2060 3450
rect 2190 3440 2310 3450
rect 2440 3440 2560 3450
rect 2690 3440 2810 3450
rect 2940 3440 3060 3450
rect 3190 3440 3310 3450
rect 3440 3440 3560 3450
rect 3690 3440 3810 3450
rect 3940 3440 4060 3450
rect 4190 3440 4310 3450
rect 4440 3440 4560 3450
rect 4690 3440 4810 3450
rect 4940 3440 5060 3450
rect 5190 3440 5310 3450
rect 5440 3440 5560 3450
rect 5690 3440 5810 3450
rect 5940 3440 6060 3450
rect 6190 3440 6310 3450
rect 6440 3440 6560 3450
rect 6690 3440 6810 3450
rect 6940 3440 7060 3450
rect 7190 3440 7310 3450
rect 7440 3440 7560 3450
rect 7690 3440 7810 3450
rect 7940 3440 8000 3450
rect 0 3425 50 3440
rect 0 3325 10 3425
rect 45 3325 50 3425
rect 0 3310 50 3325
rect 200 3425 300 3440
rect 200 3325 205 3425
rect 240 3325 260 3425
rect 295 3325 300 3425
rect 200 3310 300 3325
rect 450 3425 550 3440
rect 450 3325 455 3425
rect 490 3325 510 3425
rect 545 3325 550 3425
rect 450 3310 550 3325
rect 700 3425 800 3440
rect 700 3325 705 3425
rect 740 3325 760 3425
rect 795 3325 800 3425
rect 700 3310 800 3325
rect 950 3425 1050 3440
rect 950 3325 955 3425
rect 990 3325 1010 3425
rect 1045 3325 1050 3425
rect 950 3310 1050 3325
rect 1200 3425 1300 3440
rect 1200 3325 1205 3425
rect 1240 3325 1260 3425
rect 1295 3325 1300 3425
rect 1200 3310 1300 3325
rect 1450 3425 1550 3440
rect 1450 3325 1455 3425
rect 1490 3325 1510 3425
rect 1545 3325 1550 3425
rect 1450 3310 1550 3325
rect 1700 3425 1800 3440
rect 1700 3325 1705 3425
rect 1740 3325 1760 3425
rect 1795 3325 1800 3425
rect 1700 3310 1800 3325
rect 1950 3425 2050 3440
rect 1950 3325 1955 3425
rect 1990 3325 2010 3425
rect 2045 3325 2050 3425
rect 1950 3310 2050 3325
rect 2200 3425 2300 3440
rect 2200 3325 2205 3425
rect 2240 3325 2260 3425
rect 2295 3325 2300 3425
rect 2200 3310 2300 3325
rect 2450 3425 2550 3440
rect 2450 3325 2455 3425
rect 2490 3325 2510 3425
rect 2545 3325 2550 3425
rect 2450 3310 2550 3325
rect 2700 3425 2800 3440
rect 2700 3325 2705 3425
rect 2740 3325 2760 3425
rect 2795 3325 2800 3425
rect 2700 3310 2800 3325
rect 2950 3425 3050 3440
rect 2950 3325 2955 3425
rect 2990 3325 3010 3425
rect 3045 3325 3050 3425
rect 2950 3310 3050 3325
rect 3200 3425 3300 3440
rect 3200 3325 3205 3425
rect 3240 3325 3260 3425
rect 3295 3325 3300 3425
rect 3200 3310 3300 3325
rect 3450 3425 3550 3440
rect 3450 3325 3455 3425
rect 3490 3325 3510 3425
rect 3545 3325 3550 3425
rect 3450 3310 3550 3325
rect 3700 3425 3800 3440
rect 3700 3325 3705 3425
rect 3740 3325 3760 3425
rect 3795 3325 3800 3425
rect 3700 3310 3800 3325
rect 3950 3425 4050 3440
rect 3950 3325 3955 3425
rect 3990 3325 4010 3425
rect 4045 3325 4050 3425
rect 3950 3310 4050 3325
rect 4200 3425 4300 3440
rect 4200 3325 4205 3425
rect 4240 3325 4260 3425
rect 4295 3325 4300 3425
rect 4200 3310 4300 3325
rect 4450 3425 4550 3440
rect 4450 3325 4455 3425
rect 4490 3325 4510 3425
rect 4545 3325 4550 3425
rect 4450 3310 4550 3325
rect 4700 3425 4800 3440
rect 4700 3325 4705 3425
rect 4740 3325 4760 3425
rect 4795 3325 4800 3425
rect 4700 3310 4800 3325
rect 4950 3425 5050 3440
rect 4950 3325 4955 3425
rect 4990 3325 5010 3425
rect 5045 3325 5050 3425
rect 4950 3310 5050 3325
rect 5200 3425 5300 3440
rect 5200 3325 5205 3425
rect 5240 3325 5260 3425
rect 5295 3325 5300 3425
rect 5200 3310 5300 3325
rect 5450 3425 5550 3440
rect 5450 3325 5455 3425
rect 5490 3325 5510 3425
rect 5545 3325 5550 3425
rect 5450 3310 5550 3325
rect 5700 3425 5800 3440
rect 5700 3325 5705 3425
rect 5740 3325 5760 3425
rect 5795 3325 5800 3425
rect 5700 3310 5800 3325
rect 5950 3425 6050 3440
rect 5950 3325 5955 3425
rect 5990 3325 6010 3425
rect 6045 3325 6050 3425
rect 5950 3310 6050 3325
rect 6200 3425 6300 3440
rect 6200 3325 6205 3425
rect 6240 3325 6260 3425
rect 6295 3325 6300 3425
rect 6200 3310 6300 3325
rect 6450 3425 6550 3440
rect 6450 3325 6455 3425
rect 6490 3325 6510 3425
rect 6545 3325 6550 3425
rect 6450 3310 6550 3325
rect 6700 3425 6800 3440
rect 6700 3325 6705 3425
rect 6740 3325 6760 3425
rect 6795 3325 6800 3425
rect 6700 3310 6800 3325
rect 6950 3425 7050 3440
rect 6950 3325 6955 3425
rect 6990 3325 7010 3425
rect 7045 3325 7050 3425
rect 6950 3310 7050 3325
rect 7200 3425 7300 3440
rect 7200 3325 7205 3425
rect 7240 3325 7260 3425
rect 7295 3325 7300 3425
rect 7200 3310 7300 3325
rect 7450 3425 7550 3440
rect 7450 3325 7455 3425
rect 7490 3325 7510 3425
rect 7545 3325 7550 3425
rect 7450 3310 7550 3325
rect 7700 3425 7800 3440
rect 7700 3325 7705 3425
rect 7740 3325 7760 3425
rect 7795 3325 7800 3425
rect 7700 3310 7800 3325
rect 7950 3425 8000 3440
rect 7950 3325 7955 3425
rect 7990 3325 8000 3425
rect 7950 3310 8000 3325
rect 0 3300 60 3310
rect 190 3300 310 3310
rect 440 3300 560 3310
rect 690 3300 810 3310
rect 940 3300 1060 3310
rect 1190 3300 1310 3310
rect 1440 3300 1560 3310
rect 1690 3300 1810 3310
rect 1940 3300 2060 3310
rect 2190 3300 2310 3310
rect 2440 3300 2560 3310
rect 2690 3300 2810 3310
rect 2940 3300 3060 3310
rect 3190 3300 3310 3310
rect 3440 3300 3560 3310
rect 3690 3300 3810 3310
rect 3940 3300 4060 3310
rect 4190 3300 4310 3310
rect 4440 3300 4560 3310
rect 4690 3300 4810 3310
rect 4940 3300 5060 3310
rect 5190 3300 5310 3310
rect 5440 3300 5560 3310
rect 5690 3300 5810 3310
rect 5940 3300 6060 3310
rect 6190 3300 6310 3310
rect 6440 3300 6560 3310
rect 6690 3300 6810 3310
rect 6940 3300 7060 3310
rect 7190 3300 7310 3310
rect 7440 3300 7560 3310
rect 7690 3300 7810 3310
rect 7940 3300 8000 3310
rect 0 3295 200 3300
rect 0 3260 75 3295
rect 175 3260 200 3295
rect 0 3240 200 3260
rect 0 3205 75 3240
rect 175 3205 200 3240
rect 0 3200 200 3205
rect 300 3295 450 3300
rect 300 3260 325 3295
rect 425 3260 450 3295
rect 300 3240 450 3260
rect 300 3205 325 3240
rect 425 3205 450 3240
rect 300 3200 450 3205
rect 550 3295 700 3300
rect 550 3260 575 3295
rect 675 3260 700 3295
rect 550 3240 700 3260
rect 550 3205 575 3240
rect 675 3205 700 3240
rect 550 3200 700 3205
rect 800 3295 1200 3300
rect 800 3260 825 3295
rect 925 3260 1075 3295
rect 1175 3260 1200 3295
rect 800 3240 1200 3260
rect 800 3205 825 3240
rect 925 3205 1075 3240
rect 1175 3205 1200 3240
rect 800 3200 1200 3205
rect 1300 3295 1450 3300
rect 1300 3260 1325 3295
rect 1425 3260 1450 3295
rect 1300 3240 1450 3260
rect 1300 3205 1325 3240
rect 1425 3205 1450 3240
rect 1300 3200 1450 3205
rect 1550 3295 1700 3300
rect 1550 3260 1575 3295
rect 1675 3260 1700 3295
rect 1550 3240 1700 3260
rect 1550 3205 1575 3240
rect 1675 3205 1700 3240
rect 1550 3200 1700 3205
rect 1800 3295 2200 3300
rect 1800 3260 1825 3295
rect 1925 3260 2075 3295
rect 2175 3260 2200 3295
rect 1800 3240 2200 3260
rect 1800 3205 1825 3240
rect 1925 3205 2075 3240
rect 2175 3205 2200 3240
rect 1800 3200 2200 3205
rect 2300 3295 2450 3300
rect 2300 3260 2325 3295
rect 2425 3260 2450 3295
rect 2300 3240 2450 3260
rect 2300 3205 2325 3240
rect 2425 3205 2450 3240
rect 2300 3200 2450 3205
rect 2550 3295 2700 3300
rect 2550 3260 2575 3295
rect 2675 3260 2700 3295
rect 2550 3240 2700 3260
rect 2550 3205 2575 3240
rect 2675 3205 2700 3240
rect 2550 3200 2700 3205
rect 2800 3295 3200 3300
rect 2800 3260 2825 3295
rect 2925 3260 3075 3295
rect 3175 3260 3200 3295
rect 2800 3240 3200 3260
rect 2800 3205 2825 3240
rect 2925 3205 3075 3240
rect 3175 3205 3200 3240
rect 2800 3200 3200 3205
rect 3300 3295 3450 3300
rect 3300 3260 3325 3295
rect 3425 3260 3450 3295
rect 3300 3240 3450 3260
rect 3300 3205 3325 3240
rect 3425 3205 3450 3240
rect 3300 3200 3450 3205
rect 3550 3295 3700 3300
rect 3550 3260 3575 3295
rect 3675 3260 3700 3295
rect 3550 3240 3700 3260
rect 3550 3205 3575 3240
rect 3675 3205 3700 3240
rect 3550 3200 3700 3205
rect 3800 3295 4200 3300
rect 3800 3260 3825 3295
rect 3925 3260 4075 3295
rect 4175 3260 4200 3295
rect 3800 3240 4200 3260
rect 3800 3205 3825 3240
rect 3925 3205 4075 3240
rect 4175 3205 4200 3240
rect 3800 3200 4200 3205
rect 4300 3295 4450 3300
rect 4300 3260 4325 3295
rect 4425 3260 4450 3295
rect 4300 3240 4450 3260
rect 4300 3205 4325 3240
rect 4425 3205 4450 3240
rect 4300 3200 4450 3205
rect 4550 3295 4700 3300
rect 4550 3260 4575 3295
rect 4675 3260 4700 3295
rect 4550 3240 4700 3260
rect 4550 3205 4575 3240
rect 4675 3205 4700 3240
rect 4550 3200 4700 3205
rect 4800 3295 5200 3300
rect 4800 3260 4825 3295
rect 4925 3260 5075 3295
rect 5175 3260 5200 3295
rect 4800 3240 5200 3260
rect 4800 3205 4825 3240
rect 4925 3205 5075 3240
rect 5175 3205 5200 3240
rect 4800 3200 5200 3205
rect 5300 3295 5450 3300
rect 5300 3260 5325 3295
rect 5425 3260 5450 3295
rect 5300 3240 5450 3260
rect 5300 3205 5325 3240
rect 5425 3205 5450 3240
rect 5300 3200 5450 3205
rect 5550 3295 5700 3300
rect 5550 3260 5575 3295
rect 5675 3260 5700 3295
rect 5550 3240 5700 3260
rect 5550 3205 5575 3240
rect 5675 3205 5700 3240
rect 5550 3200 5700 3205
rect 5800 3295 6200 3300
rect 5800 3260 5825 3295
rect 5925 3260 6075 3295
rect 6175 3260 6200 3295
rect 5800 3240 6200 3260
rect 5800 3205 5825 3240
rect 5925 3205 6075 3240
rect 6175 3205 6200 3240
rect 5800 3200 6200 3205
rect 6300 3295 6450 3300
rect 6300 3260 6325 3295
rect 6425 3260 6450 3295
rect 6300 3240 6450 3260
rect 6300 3205 6325 3240
rect 6425 3205 6450 3240
rect 6300 3200 6450 3205
rect 6550 3295 6700 3300
rect 6550 3260 6575 3295
rect 6675 3260 6700 3295
rect 6550 3240 6700 3260
rect 6550 3205 6575 3240
rect 6675 3205 6700 3240
rect 6550 3200 6700 3205
rect 6800 3295 7200 3300
rect 6800 3260 6825 3295
rect 6925 3260 7075 3295
rect 7175 3260 7200 3295
rect 6800 3240 7200 3260
rect 6800 3205 6825 3240
rect 6925 3205 7075 3240
rect 7175 3205 7200 3240
rect 6800 3200 7200 3205
rect 7300 3295 7450 3300
rect 7300 3260 7325 3295
rect 7425 3260 7450 3295
rect 7300 3240 7450 3260
rect 7300 3205 7325 3240
rect 7425 3205 7450 3240
rect 7300 3200 7450 3205
rect 7550 3295 7700 3300
rect 7550 3260 7575 3295
rect 7675 3260 7700 3295
rect 7550 3240 7700 3260
rect 7550 3205 7575 3240
rect 7675 3205 7700 3240
rect 7550 3200 7700 3205
rect 7800 3295 8000 3300
rect 7800 3260 7825 3295
rect 7925 3260 8000 3295
rect 7800 3240 8000 3260
rect 7800 3205 7825 3240
rect 7925 3205 8000 3240
rect 7800 3200 8000 3205
rect 0 3190 60 3200
rect 190 3190 310 3200
rect 440 3190 560 3200
rect 690 3190 810 3200
rect 940 3190 1060 3200
rect 1190 3190 1310 3200
rect 1440 3190 1560 3200
rect 1690 3190 1810 3200
rect 1940 3190 2060 3200
rect 2190 3190 2310 3200
rect 2440 3190 2560 3200
rect 2690 3190 2810 3200
rect 2940 3190 3060 3200
rect 3190 3190 3310 3200
rect 3440 3190 3560 3200
rect 3690 3190 3810 3200
rect 3940 3190 4060 3200
rect 4190 3190 4310 3200
rect 4440 3190 4560 3200
rect 4690 3190 4810 3200
rect 4940 3190 5060 3200
rect 5190 3190 5310 3200
rect 5440 3190 5560 3200
rect 5690 3190 5810 3200
rect 5940 3190 6060 3200
rect 6190 3190 6310 3200
rect 6440 3190 6560 3200
rect 6690 3190 6810 3200
rect 6940 3190 7060 3200
rect 7190 3190 7310 3200
rect 7440 3190 7560 3200
rect 7690 3190 7810 3200
rect 7940 3190 8000 3200
rect 0 3175 50 3190
rect 0 3075 10 3175
rect 45 3075 50 3175
rect 0 3060 50 3075
rect 200 3175 300 3190
rect 200 3075 205 3175
rect 240 3075 260 3175
rect 295 3075 300 3175
rect 200 3060 300 3075
rect 450 3175 550 3190
rect 450 3075 455 3175
rect 490 3075 510 3175
rect 545 3075 550 3175
rect 450 3060 550 3075
rect 700 3175 800 3190
rect 700 3075 705 3175
rect 740 3075 760 3175
rect 795 3075 800 3175
rect 700 3060 800 3075
rect 950 3175 1050 3190
rect 950 3075 955 3175
rect 990 3075 1010 3175
rect 1045 3075 1050 3175
rect 950 3060 1050 3075
rect 1200 3175 1300 3190
rect 1200 3075 1205 3175
rect 1240 3075 1260 3175
rect 1295 3075 1300 3175
rect 1200 3060 1300 3075
rect 1450 3175 1550 3190
rect 1450 3075 1455 3175
rect 1490 3075 1510 3175
rect 1545 3075 1550 3175
rect 1450 3060 1550 3075
rect 1700 3175 1800 3190
rect 1700 3075 1705 3175
rect 1740 3075 1760 3175
rect 1795 3075 1800 3175
rect 1700 3060 1800 3075
rect 1950 3175 2050 3190
rect 1950 3075 1955 3175
rect 1990 3075 2010 3175
rect 2045 3075 2050 3175
rect 1950 3060 2050 3075
rect 2200 3175 2300 3190
rect 2200 3075 2205 3175
rect 2240 3075 2260 3175
rect 2295 3075 2300 3175
rect 2200 3060 2300 3075
rect 2450 3175 2550 3190
rect 2450 3075 2455 3175
rect 2490 3075 2510 3175
rect 2545 3075 2550 3175
rect 2450 3060 2550 3075
rect 2700 3175 2800 3190
rect 2700 3075 2705 3175
rect 2740 3075 2760 3175
rect 2795 3075 2800 3175
rect 2700 3060 2800 3075
rect 2950 3175 3050 3190
rect 2950 3075 2955 3175
rect 2990 3075 3010 3175
rect 3045 3075 3050 3175
rect 2950 3060 3050 3075
rect 3200 3175 3300 3190
rect 3200 3075 3205 3175
rect 3240 3075 3260 3175
rect 3295 3075 3300 3175
rect 3200 3060 3300 3075
rect 3450 3175 3550 3190
rect 3450 3075 3455 3175
rect 3490 3075 3510 3175
rect 3545 3075 3550 3175
rect 3450 3060 3550 3075
rect 3700 3175 3800 3190
rect 3700 3075 3705 3175
rect 3740 3075 3760 3175
rect 3795 3075 3800 3175
rect 3700 3060 3800 3075
rect 3950 3175 4050 3190
rect 3950 3075 3955 3175
rect 3990 3075 4010 3175
rect 4045 3075 4050 3175
rect 3950 3060 4050 3075
rect 4200 3175 4300 3190
rect 4200 3075 4205 3175
rect 4240 3075 4260 3175
rect 4295 3075 4300 3175
rect 4200 3060 4300 3075
rect 4450 3175 4550 3190
rect 4450 3075 4455 3175
rect 4490 3075 4510 3175
rect 4545 3075 4550 3175
rect 4450 3060 4550 3075
rect 4700 3175 4800 3190
rect 4700 3075 4705 3175
rect 4740 3075 4760 3175
rect 4795 3075 4800 3175
rect 4700 3060 4800 3075
rect 4950 3175 5050 3190
rect 4950 3075 4955 3175
rect 4990 3075 5010 3175
rect 5045 3075 5050 3175
rect 4950 3060 5050 3075
rect 5200 3175 5300 3190
rect 5200 3075 5205 3175
rect 5240 3075 5260 3175
rect 5295 3075 5300 3175
rect 5200 3060 5300 3075
rect 5450 3175 5550 3190
rect 5450 3075 5455 3175
rect 5490 3075 5510 3175
rect 5545 3075 5550 3175
rect 5450 3060 5550 3075
rect 5700 3175 5800 3190
rect 5700 3075 5705 3175
rect 5740 3075 5760 3175
rect 5795 3075 5800 3175
rect 5700 3060 5800 3075
rect 5950 3175 6050 3190
rect 5950 3075 5955 3175
rect 5990 3075 6010 3175
rect 6045 3075 6050 3175
rect 5950 3060 6050 3075
rect 6200 3175 6300 3190
rect 6200 3075 6205 3175
rect 6240 3075 6260 3175
rect 6295 3075 6300 3175
rect 6200 3060 6300 3075
rect 6450 3175 6550 3190
rect 6450 3075 6455 3175
rect 6490 3075 6510 3175
rect 6545 3075 6550 3175
rect 6450 3060 6550 3075
rect 6700 3175 6800 3190
rect 6700 3075 6705 3175
rect 6740 3075 6760 3175
rect 6795 3075 6800 3175
rect 6700 3060 6800 3075
rect 6950 3175 7050 3190
rect 6950 3075 6955 3175
rect 6990 3075 7010 3175
rect 7045 3075 7050 3175
rect 6950 3060 7050 3075
rect 7200 3175 7300 3190
rect 7200 3075 7205 3175
rect 7240 3075 7260 3175
rect 7295 3075 7300 3175
rect 7200 3060 7300 3075
rect 7450 3175 7550 3190
rect 7450 3075 7455 3175
rect 7490 3075 7510 3175
rect 7545 3075 7550 3175
rect 7450 3060 7550 3075
rect 7700 3175 7800 3190
rect 7700 3075 7705 3175
rect 7740 3075 7760 3175
rect 7795 3075 7800 3175
rect 7700 3060 7800 3075
rect 7950 3175 8000 3190
rect 7950 3075 7955 3175
rect 7990 3075 8000 3175
rect 7950 3060 8000 3075
rect 0 3050 60 3060
rect 190 3050 310 3060
rect 440 3050 560 3060
rect 690 3050 810 3060
rect 940 3050 1060 3060
rect 1190 3050 1310 3060
rect 1440 3050 1560 3060
rect 1690 3050 1810 3060
rect 1940 3050 2060 3060
rect 2190 3050 2310 3060
rect 2440 3050 2560 3060
rect 2690 3050 2810 3060
rect 2940 3050 3060 3060
rect 3190 3050 3310 3060
rect 3440 3050 3560 3060
rect 3690 3050 3810 3060
rect 3940 3050 4060 3060
rect 4190 3050 4310 3060
rect 4440 3050 4560 3060
rect 4690 3050 4810 3060
rect 4940 3050 5060 3060
rect 5190 3050 5310 3060
rect 5440 3050 5560 3060
rect 5690 3050 5810 3060
rect 5940 3050 6060 3060
rect 6190 3050 6310 3060
rect 6440 3050 6560 3060
rect 6690 3050 6810 3060
rect 6940 3050 7060 3060
rect 7190 3050 7310 3060
rect 7440 3050 7560 3060
rect 7690 3050 7810 3060
rect 7940 3050 8000 3060
rect 0 3045 450 3050
rect 0 3010 75 3045
rect 175 3010 325 3045
rect 425 3010 450 3045
rect 0 2990 450 3010
rect 0 2955 75 2990
rect 175 2955 325 2990
rect 425 2955 450 2990
rect 0 2950 450 2955
rect 550 3045 1450 3050
rect 550 3010 575 3045
rect 675 3010 825 3045
rect 925 3010 1075 3045
rect 1175 3010 1325 3045
rect 1425 3010 1450 3045
rect 550 2990 1450 3010
rect 550 2955 575 2990
rect 675 2955 825 2990
rect 925 2955 1075 2990
rect 1175 2955 1325 2990
rect 1425 2955 1450 2990
rect 550 2950 1450 2955
rect 1550 3045 2450 3050
rect 1550 3010 1575 3045
rect 1675 3010 1825 3045
rect 1925 3010 2075 3045
rect 2175 3010 2325 3045
rect 2425 3010 2450 3045
rect 1550 2990 2450 3010
rect 1550 2955 1575 2990
rect 1675 2955 1825 2990
rect 1925 2955 2075 2990
rect 2175 2955 2325 2990
rect 2425 2955 2450 2990
rect 1550 2950 2450 2955
rect 2550 3045 3450 3050
rect 2550 3010 2575 3045
rect 2675 3010 2825 3045
rect 2925 3010 3075 3045
rect 3175 3010 3325 3045
rect 3425 3010 3450 3045
rect 2550 2990 3450 3010
rect 2550 2955 2575 2990
rect 2675 2955 2825 2990
rect 2925 2955 3075 2990
rect 3175 2955 3325 2990
rect 3425 2955 3450 2990
rect 2550 2950 3450 2955
rect 3550 3045 4450 3050
rect 3550 3010 3575 3045
rect 3675 3010 3825 3045
rect 3925 3010 4075 3045
rect 4175 3010 4325 3045
rect 4425 3010 4450 3045
rect 3550 2990 4450 3010
rect 3550 2955 3575 2990
rect 3675 2955 3825 2990
rect 3925 2955 4075 2990
rect 4175 2955 4325 2990
rect 4425 2955 4450 2990
rect 3550 2950 4450 2955
rect 4550 3045 5450 3050
rect 4550 3010 4575 3045
rect 4675 3010 4825 3045
rect 4925 3010 5075 3045
rect 5175 3010 5325 3045
rect 5425 3010 5450 3045
rect 4550 2990 5450 3010
rect 4550 2955 4575 2990
rect 4675 2955 4825 2990
rect 4925 2955 5075 2990
rect 5175 2955 5325 2990
rect 5425 2955 5450 2990
rect 4550 2950 5450 2955
rect 5550 3045 6450 3050
rect 5550 3010 5575 3045
rect 5675 3010 5825 3045
rect 5925 3010 6075 3045
rect 6175 3010 6325 3045
rect 6425 3010 6450 3045
rect 5550 2990 6450 3010
rect 5550 2955 5575 2990
rect 5675 2955 5825 2990
rect 5925 2955 6075 2990
rect 6175 2955 6325 2990
rect 6425 2955 6450 2990
rect 5550 2950 6450 2955
rect 6550 3045 7450 3050
rect 6550 3010 6575 3045
rect 6675 3010 6825 3045
rect 6925 3010 7075 3045
rect 7175 3010 7325 3045
rect 7425 3010 7450 3045
rect 6550 2990 7450 3010
rect 6550 2955 6575 2990
rect 6675 2955 6825 2990
rect 6925 2955 7075 2990
rect 7175 2955 7325 2990
rect 7425 2955 7450 2990
rect 6550 2950 7450 2955
rect 7550 3045 8000 3050
rect 7550 3010 7575 3045
rect 7675 3010 7825 3045
rect 7925 3010 8000 3045
rect 7550 2990 8000 3010
rect 7550 2955 7575 2990
rect 7675 2955 7825 2990
rect 7925 2955 8000 2990
rect 7550 2950 8000 2955
rect 0 2940 60 2950
rect 190 2940 310 2950
rect 440 2940 560 2950
rect 690 2940 810 2950
rect 940 2940 1060 2950
rect 1190 2940 1310 2950
rect 1440 2940 1560 2950
rect 1690 2940 1810 2950
rect 1940 2940 2060 2950
rect 2190 2940 2310 2950
rect 2440 2940 2560 2950
rect 2690 2940 2810 2950
rect 2940 2940 3060 2950
rect 3190 2940 3310 2950
rect 3440 2940 3560 2950
rect 3690 2940 3810 2950
rect 3940 2940 4060 2950
rect 4190 2940 4310 2950
rect 4440 2940 4560 2950
rect 4690 2940 4810 2950
rect 4940 2940 5060 2950
rect 5190 2940 5310 2950
rect 5440 2940 5560 2950
rect 5690 2940 5810 2950
rect 5940 2940 6060 2950
rect 6190 2940 6310 2950
rect 6440 2940 6560 2950
rect 6690 2940 6810 2950
rect 6940 2940 7060 2950
rect 7190 2940 7310 2950
rect 7440 2940 7560 2950
rect 7690 2940 7810 2950
rect 7940 2940 8000 2950
rect 0 2925 50 2940
rect 0 2825 10 2925
rect 45 2825 50 2925
rect 0 2810 50 2825
rect 200 2925 300 2940
rect 200 2825 205 2925
rect 240 2825 260 2925
rect 295 2825 300 2925
rect 200 2810 300 2825
rect 450 2925 550 2940
rect 450 2825 455 2925
rect 490 2825 510 2925
rect 545 2825 550 2925
rect 450 2810 550 2825
rect 700 2925 800 2940
rect 700 2825 705 2925
rect 740 2825 760 2925
rect 795 2825 800 2925
rect 700 2810 800 2825
rect 950 2925 1050 2940
rect 950 2825 955 2925
rect 990 2825 1010 2925
rect 1045 2825 1050 2925
rect 950 2810 1050 2825
rect 1200 2925 1300 2940
rect 1200 2825 1205 2925
rect 1240 2825 1260 2925
rect 1295 2825 1300 2925
rect 1200 2810 1300 2825
rect 1450 2925 1550 2940
rect 1450 2825 1455 2925
rect 1490 2825 1510 2925
rect 1545 2825 1550 2925
rect 1450 2810 1550 2825
rect 1700 2925 1800 2940
rect 1700 2825 1705 2925
rect 1740 2825 1760 2925
rect 1795 2825 1800 2925
rect 1700 2810 1800 2825
rect 1950 2925 2050 2940
rect 1950 2825 1955 2925
rect 1990 2825 2010 2925
rect 2045 2825 2050 2925
rect 1950 2810 2050 2825
rect 2200 2925 2300 2940
rect 2200 2825 2205 2925
rect 2240 2825 2260 2925
rect 2295 2825 2300 2925
rect 2200 2810 2300 2825
rect 2450 2925 2550 2940
rect 2450 2825 2455 2925
rect 2490 2825 2510 2925
rect 2545 2825 2550 2925
rect 2450 2810 2550 2825
rect 2700 2925 2800 2940
rect 2700 2825 2705 2925
rect 2740 2825 2760 2925
rect 2795 2825 2800 2925
rect 2700 2810 2800 2825
rect 2950 2925 3050 2940
rect 2950 2825 2955 2925
rect 2990 2825 3010 2925
rect 3045 2825 3050 2925
rect 2950 2810 3050 2825
rect 3200 2925 3300 2940
rect 3200 2825 3205 2925
rect 3240 2825 3260 2925
rect 3295 2825 3300 2925
rect 3200 2810 3300 2825
rect 3450 2925 3550 2940
rect 3450 2825 3455 2925
rect 3490 2825 3510 2925
rect 3545 2825 3550 2925
rect 3450 2810 3550 2825
rect 3700 2925 3800 2940
rect 3700 2825 3705 2925
rect 3740 2825 3760 2925
rect 3795 2825 3800 2925
rect 3700 2810 3800 2825
rect 3950 2925 4050 2940
rect 3950 2825 3955 2925
rect 3990 2825 4010 2925
rect 4045 2825 4050 2925
rect 3950 2810 4050 2825
rect 4200 2925 4300 2940
rect 4200 2825 4205 2925
rect 4240 2825 4260 2925
rect 4295 2825 4300 2925
rect 4200 2810 4300 2825
rect 4450 2925 4550 2940
rect 4450 2825 4455 2925
rect 4490 2825 4510 2925
rect 4545 2825 4550 2925
rect 4450 2810 4550 2825
rect 4700 2925 4800 2940
rect 4700 2825 4705 2925
rect 4740 2825 4760 2925
rect 4795 2825 4800 2925
rect 4700 2810 4800 2825
rect 4950 2925 5050 2940
rect 4950 2825 4955 2925
rect 4990 2825 5010 2925
rect 5045 2825 5050 2925
rect 4950 2810 5050 2825
rect 5200 2925 5300 2940
rect 5200 2825 5205 2925
rect 5240 2825 5260 2925
rect 5295 2825 5300 2925
rect 5200 2810 5300 2825
rect 5450 2925 5550 2940
rect 5450 2825 5455 2925
rect 5490 2825 5510 2925
rect 5545 2825 5550 2925
rect 5450 2810 5550 2825
rect 5700 2925 5800 2940
rect 5700 2825 5705 2925
rect 5740 2825 5760 2925
rect 5795 2825 5800 2925
rect 5700 2810 5800 2825
rect 5950 2925 6050 2940
rect 5950 2825 5955 2925
rect 5990 2825 6010 2925
rect 6045 2825 6050 2925
rect 5950 2810 6050 2825
rect 6200 2925 6300 2940
rect 6200 2825 6205 2925
rect 6240 2825 6260 2925
rect 6295 2825 6300 2925
rect 6200 2810 6300 2825
rect 6450 2925 6550 2940
rect 6450 2825 6455 2925
rect 6490 2825 6510 2925
rect 6545 2825 6550 2925
rect 6450 2810 6550 2825
rect 6700 2925 6800 2940
rect 6700 2825 6705 2925
rect 6740 2825 6760 2925
rect 6795 2825 6800 2925
rect 6700 2810 6800 2825
rect 6950 2925 7050 2940
rect 6950 2825 6955 2925
rect 6990 2825 7010 2925
rect 7045 2825 7050 2925
rect 6950 2810 7050 2825
rect 7200 2925 7300 2940
rect 7200 2825 7205 2925
rect 7240 2825 7260 2925
rect 7295 2825 7300 2925
rect 7200 2810 7300 2825
rect 7450 2925 7550 2940
rect 7450 2825 7455 2925
rect 7490 2825 7510 2925
rect 7545 2825 7550 2925
rect 7450 2810 7550 2825
rect 7700 2925 7800 2940
rect 7700 2825 7705 2925
rect 7740 2825 7760 2925
rect 7795 2825 7800 2925
rect 7700 2810 7800 2825
rect 7950 2925 8000 2940
rect 7950 2825 7955 2925
rect 7990 2825 8000 2925
rect 7950 2810 8000 2825
rect 0 2800 60 2810
rect 190 2800 310 2810
rect 440 2800 560 2810
rect 690 2800 810 2810
rect 940 2800 1060 2810
rect 1190 2800 1310 2810
rect 1440 2800 1560 2810
rect 1690 2800 1810 2810
rect 1940 2800 2060 2810
rect 2190 2800 2310 2810
rect 2440 2800 2560 2810
rect 2690 2800 2810 2810
rect 2940 2800 3060 2810
rect 3190 2800 3310 2810
rect 3440 2800 3560 2810
rect 3690 2800 3810 2810
rect 3940 2800 4060 2810
rect 4190 2800 4310 2810
rect 4440 2800 4560 2810
rect 4690 2800 4810 2810
rect 4940 2800 5060 2810
rect 5190 2800 5310 2810
rect 5440 2800 5560 2810
rect 5690 2800 5810 2810
rect 5940 2800 6060 2810
rect 6190 2800 6310 2810
rect 6440 2800 6560 2810
rect 6690 2800 6810 2810
rect 6940 2800 7060 2810
rect 7190 2800 7310 2810
rect 7440 2800 7560 2810
rect 7690 2800 7810 2810
rect 7940 2800 8000 2810
rect 0 2795 200 2800
rect 0 2760 75 2795
rect 175 2760 200 2795
rect 0 2740 200 2760
rect 0 2705 75 2740
rect 175 2705 200 2740
rect 0 2700 200 2705
rect 300 2795 450 2800
rect 300 2760 325 2795
rect 425 2760 450 2795
rect 300 2740 450 2760
rect 300 2705 325 2740
rect 425 2705 450 2740
rect 300 2700 450 2705
rect 550 2795 700 2800
rect 550 2760 575 2795
rect 675 2760 700 2795
rect 550 2740 700 2760
rect 550 2705 575 2740
rect 675 2705 700 2740
rect 550 2700 700 2705
rect 800 2795 1200 2800
rect 800 2760 825 2795
rect 925 2760 1075 2795
rect 1175 2760 1200 2795
rect 800 2740 1200 2760
rect 800 2705 825 2740
rect 925 2705 1075 2740
rect 1175 2705 1200 2740
rect 800 2700 1200 2705
rect 1300 2795 1450 2800
rect 1300 2760 1325 2795
rect 1425 2760 1450 2795
rect 1300 2740 1450 2760
rect 1300 2705 1325 2740
rect 1425 2705 1450 2740
rect 1300 2700 1450 2705
rect 1550 2795 1700 2800
rect 1550 2760 1575 2795
rect 1675 2760 1700 2795
rect 1550 2740 1700 2760
rect 1550 2705 1575 2740
rect 1675 2705 1700 2740
rect 1550 2700 1700 2705
rect 1800 2795 2200 2800
rect 1800 2760 1825 2795
rect 1925 2760 2075 2795
rect 2175 2760 2200 2795
rect 1800 2740 2200 2760
rect 1800 2705 1825 2740
rect 1925 2705 2075 2740
rect 2175 2705 2200 2740
rect 1800 2700 2200 2705
rect 2300 2795 2450 2800
rect 2300 2760 2325 2795
rect 2425 2760 2450 2795
rect 2300 2740 2450 2760
rect 2300 2705 2325 2740
rect 2425 2705 2450 2740
rect 2300 2700 2450 2705
rect 2550 2795 2700 2800
rect 2550 2760 2575 2795
rect 2675 2760 2700 2795
rect 2550 2740 2700 2760
rect 2550 2705 2575 2740
rect 2675 2705 2700 2740
rect 2550 2700 2700 2705
rect 2800 2795 3200 2800
rect 2800 2760 2825 2795
rect 2925 2760 3075 2795
rect 3175 2760 3200 2795
rect 2800 2740 3200 2760
rect 2800 2705 2825 2740
rect 2925 2705 3075 2740
rect 3175 2705 3200 2740
rect 2800 2700 3200 2705
rect 3300 2795 3450 2800
rect 3300 2760 3325 2795
rect 3425 2760 3450 2795
rect 3300 2740 3450 2760
rect 3300 2705 3325 2740
rect 3425 2705 3450 2740
rect 3300 2700 3450 2705
rect 3550 2795 3700 2800
rect 3550 2760 3575 2795
rect 3675 2760 3700 2795
rect 3550 2740 3700 2760
rect 3550 2705 3575 2740
rect 3675 2705 3700 2740
rect 3550 2700 3700 2705
rect 3800 2795 4200 2800
rect 3800 2760 3825 2795
rect 3925 2760 4075 2795
rect 4175 2760 4200 2795
rect 3800 2740 4200 2760
rect 3800 2705 3825 2740
rect 3925 2705 4075 2740
rect 4175 2705 4200 2740
rect 3800 2700 4200 2705
rect 4300 2795 4450 2800
rect 4300 2760 4325 2795
rect 4425 2760 4450 2795
rect 4300 2740 4450 2760
rect 4300 2705 4325 2740
rect 4425 2705 4450 2740
rect 4300 2700 4450 2705
rect 4550 2795 4700 2800
rect 4550 2760 4575 2795
rect 4675 2760 4700 2795
rect 4550 2740 4700 2760
rect 4550 2705 4575 2740
rect 4675 2705 4700 2740
rect 4550 2700 4700 2705
rect 4800 2795 5200 2800
rect 4800 2760 4825 2795
rect 4925 2760 5075 2795
rect 5175 2760 5200 2795
rect 4800 2740 5200 2760
rect 4800 2705 4825 2740
rect 4925 2705 5075 2740
rect 5175 2705 5200 2740
rect 4800 2700 5200 2705
rect 5300 2795 5450 2800
rect 5300 2760 5325 2795
rect 5425 2760 5450 2795
rect 5300 2740 5450 2760
rect 5300 2705 5325 2740
rect 5425 2705 5450 2740
rect 5300 2700 5450 2705
rect 5550 2795 5700 2800
rect 5550 2760 5575 2795
rect 5675 2760 5700 2795
rect 5550 2740 5700 2760
rect 5550 2705 5575 2740
rect 5675 2705 5700 2740
rect 5550 2700 5700 2705
rect 5800 2795 6200 2800
rect 5800 2760 5825 2795
rect 5925 2760 6075 2795
rect 6175 2760 6200 2795
rect 5800 2740 6200 2760
rect 5800 2705 5825 2740
rect 5925 2705 6075 2740
rect 6175 2705 6200 2740
rect 5800 2700 6200 2705
rect 6300 2795 6450 2800
rect 6300 2760 6325 2795
rect 6425 2760 6450 2795
rect 6300 2740 6450 2760
rect 6300 2705 6325 2740
rect 6425 2705 6450 2740
rect 6300 2700 6450 2705
rect 6550 2795 6700 2800
rect 6550 2760 6575 2795
rect 6675 2760 6700 2795
rect 6550 2740 6700 2760
rect 6550 2705 6575 2740
rect 6675 2705 6700 2740
rect 6550 2700 6700 2705
rect 6800 2795 7200 2800
rect 6800 2760 6825 2795
rect 6925 2760 7075 2795
rect 7175 2760 7200 2795
rect 6800 2740 7200 2760
rect 6800 2705 6825 2740
rect 6925 2705 7075 2740
rect 7175 2705 7200 2740
rect 6800 2700 7200 2705
rect 7300 2795 7450 2800
rect 7300 2760 7325 2795
rect 7425 2760 7450 2795
rect 7300 2740 7450 2760
rect 7300 2705 7325 2740
rect 7425 2705 7450 2740
rect 7300 2700 7450 2705
rect 7550 2795 7700 2800
rect 7550 2760 7575 2795
rect 7675 2760 7700 2795
rect 7550 2740 7700 2760
rect 7550 2705 7575 2740
rect 7675 2705 7700 2740
rect 7550 2700 7700 2705
rect 7800 2795 8000 2800
rect 7800 2760 7825 2795
rect 7925 2760 8000 2795
rect 7800 2740 8000 2760
rect 7800 2705 7825 2740
rect 7925 2705 8000 2740
rect 7800 2700 8000 2705
rect 0 2690 60 2700
rect 190 2690 310 2700
rect 440 2690 560 2700
rect 690 2690 810 2700
rect 940 2690 1060 2700
rect 1190 2690 1310 2700
rect 1440 2690 1560 2700
rect 1690 2690 1810 2700
rect 1940 2690 2060 2700
rect 2190 2690 2310 2700
rect 2440 2690 2560 2700
rect 2690 2690 2810 2700
rect 2940 2690 3060 2700
rect 3190 2690 3310 2700
rect 3440 2690 3560 2700
rect 3690 2690 3810 2700
rect 3940 2690 4060 2700
rect 4190 2690 4310 2700
rect 4440 2690 4560 2700
rect 4690 2690 4810 2700
rect 4940 2690 5060 2700
rect 5190 2690 5310 2700
rect 5440 2690 5560 2700
rect 5690 2690 5810 2700
rect 5940 2690 6060 2700
rect 6190 2690 6310 2700
rect 6440 2690 6560 2700
rect 6690 2690 6810 2700
rect 6940 2690 7060 2700
rect 7190 2690 7310 2700
rect 7440 2690 7560 2700
rect 7690 2690 7810 2700
rect 7940 2690 8000 2700
rect 0 2675 50 2690
rect 0 2575 10 2675
rect 45 2575 50 2675
rect 0 2560 50 2575
rect 200 2675 300 2690
rect 200 2575 205 2675
rect 240 2575 260 2675
rect 295 2575 300 2675
rect 200 2560 300 2575
rect 450 2675 550 2690
rect 450 2575 455 2675
rect 490 2575 510 2675
rect 545 2575 550 2675
rect 450 2560 550 2575
rect 700 2675 800 2690
rect 700 2575 705 2675
rect 740 2575 760 2675
rect 795 2575 800 2675
rect 700 2560 800 2575
rect 950 2675 1050 2690
rect 950 2575 955 2675
rect 990 2575 1010 2675
rect 1045 2575 1050 2675
rect 950 2560 1050 2575
rect 1200 2675 1300 2690
rect 1200 2575 1205 2675
rect 1240 2575 1260 2675
rect 1295 2575 1300 2675
rect 1200 2560 1300 2575
rect 1450 2675 1550 2690
rect 1450 2575 1455 2675
rect 1490 2575 1510 2675
rect 1545 2575 1550 2675
rect 1450 2560 1550 2575
rect 1700 2675 1800 2690
rect 1700 2575 1705 2675
rect 1740 2575 1760 2675
rect 1795 2575 1800 2675
rect 1700 2560 1800 2575
rect 1950 2675 2050 2690
rect 1950 2575 1955 2675
rect 1990 2575 2010 2675
rect 2045 2575 2050 2675
rect 1950 2560 2050 2575
rect 2200 2675 2300 2690
rect 2200 2575 2205 2675
rect 2240 2575 2260 2675
rect 2295 2575 2300 2675
rect 2200 2560 2300 2575
rect 2450 2675 2550 2690
rect 2450 2575 2455 2675
rect 2490 2575 2510 2675
rect 2545 2575 2550 2675
rect 2450 2560 2550 2575
rect 2700 2675 2800 2690
rect 2700 2575 2705 2675
rect 2740 2575 2760 2675
rect 2795 2575 2800 2675
rect 2700 2560 2800 2575
rect 2950 2675 3050 2690
rect 2950 2575 2955 2675
rect 2990 2575 3010 2675
rect 3045 2575 3050 2675
rect 2950 2560 3050 2575
rect 3200 2675 3300 2690
rect 3200 2575 3205 2675
rect 3240 2575 3260 2675
rect 3295 2575 3300 2675
rect 3200 2560 3300 2575
rect 3450 2675 3550 2690
rect 3450 2575 3455 2675
rect 3490 2575 3510 2675
rect 3545 2575 3550 2675
rect 3450 2560 3550 2575
rect 3700 2675 3800 2690
rect 3700 2575 3705 2675
rect 3740 2575 3760 2675
rect 3795 2575 3800 2675
rect 3700 2560 3800 2575
rect 3950 2675 4050 2690
rect 3950 2575 3955 2675
rect 3990 2575 4010 2675
rect 4045 2575 4050 2675
rect 3950 2560 4050 2575
rect 4200 2675 4300 2690
rect 4200 2575 4205 2675
rect 4240 2575 4260 2675
rect 4295 2575 4300 2675
rect 4200 2560 4300 2575
rect 4450 2675 4550 2690
rect 4450 2575 4455 2675
rect 4490 2575 4510 2675
rect 4545 2575 4550 2675
rect 4450 2560 4550 2575
rect 4700 2675 4800 2690
rect 4700 2575 4705 2675
rect 4740 2575 4760 2675
rect 4795 2575 4800 2675
rect 4700 2560 4800 2575
rect 4950 2675 5050 2690
rect 4950 2575 4955 2675
rect 4990 2575 5010 2675
rect 5045 2575 5050 2675
rect 4950 2560 5050 2575
rect 5200 2675 5300 2690
rect 5200 2575 5205 2675
rect 5240 2575 5260 2675
rect 5295 2575 5300 2675
rect 5200 2560 5300 2575
rect 5450 2675 5550 2690
rect 5450 2575 5455 2675
rect 5490 2575 5510 2675
rect 5545 2575 5550 2675
rect 5450 2560 5550 2575
rect 5700 2675 5800 2690
rect 5700 2575 5705 2675
rect 5740 2575 5760 2675
rect 5795 2575 5800 2675
rect 5700 2560 5800 2575
rect 5950 2675 6050 2690
rect 5950 2575 5955 2675
rect 5990 2575 6010 2675
rect 6045 2575 6050 2675
rect 5950 2560 6050 2575
rect 6200 2675 6300 2690
rect 6200 2575 6205 2675
rect 6240 2575 6260 2675
rect 6295 2575 6300 2675
rect 6200 2560 6300 2575
rect 6450 2675 6550 2690
rect 6450 2575 6455 2675
rect 6490 2575 6510 2675
rect 6545 2575 6550 2675
rect 6450 2560 6550 2575
rect 6700 2675 6800 2690
rect 6700 2575 6705 2675
rect 6740 2575 6760 2675
rect 6795 2575 6800 2675
rect 6700 2560 6800 2575
rect 6950 2675 7050 2690
rect 6950 2575 6955 2675
rect 6990 2575 7010 2675
rect 7045 2575 7050 2675
rect 6950 2560 7050 2575
rect 7200 2675 7300 2690
rect 7200 2575 7205 2675
rect 7240 2575 7260 2675
rect 7295 2575 7300 2675
rect 7200 2560 7300 2575
rect 7450 2675 7550 2690
rect 7450 2575 7455 2675
rect 7490 2575 7510 2675
rect 7545 2575 7550 2675
rect 7450 2560 7550 2575
rect 7700 2675 7800 2690
rect 7700 2575 7705 2675
rect 7740 2575 7760 2675
rect 7795 2575 7800 2675
rect 7700 2560 7800 2575
rect 7950 2675 8000 2690
rect 7950 2575 7955 2675
rect 7990 2575 8000 2675
rect 7950 2560 8000 2575
rect 0 2550 60 2560
rect 190 2550 310 2560
rect 440 2550 560 2560
rect 690 2550 810 2560
rect 940 2550 1060 2560
rect 1190 2550 1310 2560
rect 1440 2550 1560 2560
rect 1690 2550 1810 2560
rect 1940 2550 2060 2560
rect 2190 2550 2310 2560
rect 2440 2550 2560 2560
rect 2690 2550 2810 2560
rect 2940 2550 3060 2560
rect 3190 2550 3310 2560
rect 3440 2550 3560 2560
rect 3690 2550 3810 2560
rect 3940 2550 4060 2560
rect 4190 2550 4310 2560
rect 4440 2550 4560 2560
rect 4690 2550 4810 2560
rect 4940 2550 5060 2560
rect 5190 2550 5310 2560
rect 5440 2550 5560 2560
rect 5690 2550 5810 2560
rect 5940 2550 6060 2560
rect 6190 2550 6310 2560
rect 6440 2550 6560 2560
rect 6690 2550 6810 2560
rect 6940 2550 7060 2560
rect 7190 2550 7310 2560
rect 7440 2550 7560 2560
rect 7690 2550 7810 2560
rect 7940 2550 8000 2560
rect 0 2545 200 2550
rect 0 2510 75 2545
rect 175 2510 200 2545
rect 0 2490 200 2510
rect 0 2455 75 2490
rect 175 2455 200 2490
rect 0 2450 200 2455
rect 300 2545 450 2550
rect 300 2510 325 2545
rect 425 2510 450 2545
rect 300 2490 450 2510
rect 300 2455 325 2490
rect 425 2455 450 2490
rect 300 2450 450 2455
rect 550 2545 700 2550
rect 550 2510 575 2545
rect 675 2510 700 2545
rect 550 2490 700 2510
rect 550 2455 575 2490
rect 675 2455 700 2490
rect 550 2450 700 2455
rect 800 2545 950 2550
rect 800 2510 825 2545
rect 925 2510 950 2545
rect 800 2490 950 2510
rect 800 2455 825 2490
rect 925 2455 950 2490
rect 800 2450 950 2455
rect 1050 2545 1200 2550
rect 1050 2510 1075 2545
rect 1175 2510 1200 2545
rect 1050 2490 1200 2510
rect 1050 2455 1075 2490
rect 1175 2455 1200 2490
rect 1050 2450 1200 2455
rect 1300 2545 1450 2550
rect 1300 2510 1325 2545
rect 1425 2510 1450 2545
rect 1300 2490 1450 2510
rect 1300 2455 1325 2490
rect 1425 2455 1450 2490
rect 1300 2450 1450 2455
rect 1550 2545 1700 2550
rect 1550 2510 1575 2545
rect 1675 2510 1700 2545
rect 1550 2490 1700 2510
rect 1550 2455 1575 2490
rect 1675 2455 1700 2490
rect 1550 2450 1700 2455
rect 1800 2545 2200 2550
rect 1800 2510 1825 2545
rect 1925 2510 2075 2545
rect 2175 2510 2200 2545
rect 1800 2490 2200 2510
rect 1800 2455 1825 2490
rect 1925 2455 2075 2490
rect 2175 2455 2200 2490
rect 1800 2450 2200 2455
rect 2300 2545 2450 2550
rect 2300 2510 2325 2545
rect 2425 2510 2450 2545
rect 2300 2490 2450 2510
rect 2300 2455 2325 2490
rect 2425 2455 2450 2490
rect 2300 2450 2450 2455
rect 2550 2545 2700 2550
rect 2550 2510 2575 2545
rect 2675 2510 2700 2545
rect 2550 2490 2700 2510
rect 2550 2455 2575 2490
rect 2675 2455 2700 2490
rect 2550 2450 2700 2455
rect 2800 2545 2950 2550
rect 2800 2510 2825 2545
rect 2925 2510 2950 2545
rect 2800 2490 2950 2510
rect 2800 2455 2825 2490
rect 2925 2455 2950 2490
rect 2800 2450 2950 2455
rect 3050 2545 3200 2550
rect 3050 2510 3075 2545
rect 3175 2510 3200 2545
rect 3050 2490 3200 2510
rect 3050 2455 3075 2490
rect 3175 2455 3200 2490
rect 3050 2450 3200 2455
rect 3300 2545 3450 2550
rect 3300 2510 3325 2545
rect 3425 2510 3450 2545
rect 3300 2490 3450 2510
rect 3300 2455 3325 2490
rect 3425 2455 3450 2490
rect 3300 2450 3450 2455
rect 3550 2545 3700 2550
rect 3550 2510 3575 2545
rect 3675 2510 3700 2545
rect 3550 2490 3700 2510
rect 3550 2455 3575 2490
rect 3675 2455 3700 2490
rect 3550 2450 3700 2455
rect 3800 2545 4200 2550
rect 3800 2510 3825 2545
rect 3925 2510 4075 2545
rect 4175 2510 4200 2545
rect 3800 2490 4200 2510
rect 3800 2455 3825 2490
rect 3925 2455 4075 2490
rect 4175 2455 4200 2490
rect 3800 2450 4200 2455
rect 4300 2545 4450 2550
rect 4300 2510 4325 2545
rect 4425 2510 4450 2545
rect 4300 2490 4450 2510
rect 4300 2455 4325 2490
rect 4425 2455 4450 2490
rect 4300 2450 4450 2455
rect 4550 2545 4700 2550
rect 4550 2510 4575 2545
rect 4675 2510 4700 2545
rect 4550 2490 4700 2510
rect 4550 2455 4575 2490
rect 4675 2455 4700 2490
rect 4550 2450 4700 2455
rect 4800 2545 4950 2550
rect 4800 2510 4825 2545
rect 4925 2510 4950 2545
rect 4800 2490 4950 2510
rect 4800 2455 4825 2490
rect 4925 2455 4950 2490
rect 4800 2450 4950 2455
rect 5050 2545 5200 2550
rect 5050 2510 5075 2545
rect 5175 2510 5200 2545
rect 5050 2490 5200 2510
rect 5050 2455 5075 2490
rect 5175 2455 5200 2490
rect 5050 2450 5200 2455
rect 5300 2545 5450 2550
rect 5300 2510 5325 2545
rect 5425 2510 5450 2545
rect 5300 2490 5450 2510
rect 5300 2455 5325 2490
rect 5425 2455 5450 2490
rect 5300 2450 5450 2455
rect 5550 2545 5700 2550
rect 5550 2510 5575 2545
rect 5675 2510 5700 2545
rect 5550 2490 5700 2510
rect 5550 2455 5575 2490
rect 5675 2455 5700 2490
rect 5550 2450 5700 2455
rect 5800 2545 6200 2550
rect 5800 2510 5825 2545
rect 5925 2510 6075 2545
rect 6175 2510 6200 2545
rect 5800 2490 6200 2510
rect 5800 2455 5825 2490
rect 5925 2455 6075 2490
rect 6175 2455 6200 2490
rect 5800 2450 6200 2455
rect 6300 2545 6450 2550
rect 6300 2510 6325 2545
rect 6425 2510 6450 2545
rect 6300 2490 6450 2510
rect 6300 2455 6325 2490
rect 6425 2455 6450 2490
rect 6300 2450 6450 2455
rect 6550 2545 6700 2550
rect 6550 2510 6575 2545
rect 6675 2510 6700 2545
rect 6550 2490 6700 2510
rect 6550 2455 6575 2490
rect 6675 2455 6700 2490
rect 6550 2450 6700 2455
rect 6800 2545 6950 2550
rect 6800 2510 6825 2545
rect 6925 2510 6950 2545
rect 6800 2490 6950 2510
rect 6800 2455 6825 2490
rect 6925 2455 6950 2490
rect 6800 2450 6950 2455
rect 7050 2545 7200 2550
rect 7050 2510 7075 2545
rect 7175 2510 7200 2545
rect 7050 2490 7200 2510
rect 7050 2455 7075 2490
rect 7175 2455 7200 2490
rect 7050 2450 7200 2455
rect 7300 2545 7450 2550
rect 7300 2510 7325 2545
rect 7425 2510 7450 2545
rect 7300 2490 7450 2510
rect 7300 2455 7325 2490
rect 7425 2455 7450 2490
rect 7300 2450 7450 2455
rect 7550 2545 7700 2550
rect 7550 2510 7575 2545
rect 7675 2510 7700 2545
rect 7550 2490 7700 2510
rect 7550 2455 7575 2490
rect 7675 2455 7700 2490
rect 7550 2450 7700 2455
rect 7800 2545 8000 2550
rect 7800 2510 7825 2545
rect 7925 2510 8000 2545
rect 7800 2490 8000 2510
rect 7800 2455 7825 2490
rect 7925 2455 8000 2490
rect 7800 2450 8000 2455
rect 0 2440 60 2450
rect 190 2440 310 2450
rect 440 2440 560 2450
rect 690 2440 810 2450
rect 940 2440 1060 2450
rect 1190 2440 1310 2450
rect 1440 2440 1560 2450
rect 1690 2440 1810 2450
rect 1940 2440 2060 2450
rect 2190 2440 2310 2450
rect 2440 2440 2560 2450
rect 2690 2440 2810 2450
rect 2940 2440 3060 2450
rect 3190 2440 3310 2450
rect 3440 2440 3560 2450
rect 3690 2440 3810 2450
rect 3940 2440 4060 2450
rect 4190 2440 4310 2450
rect 4440 2440 4560 2450
rect 4690 2440 4810 2450
rect 4940 2440 5060 2450
rect 5190 2440 5310 2450
rect 5440 2440 5560 2450
rect 5690 2440 5810 2450
rect 5940 2440 6060 2450
rect 6190 2440 6310 2450
rect 6440 2440 6560 2450
rect 6690 2440 6810 2450
rect 6940 2440 7060 2450
rect 7190 2440 7310 2450
rect 7440 2440 7560 2450
rect 7690 2440 7810 2450
rect 7940 2440 8000 2450
rect 0 2425 50 2440
rect 0 2325 10 2425
rect 45 2325 50 2425
rect 0 2310 50 2325
rect 200 2425 300 2440
rect 200 2325 205 2425
rect 240 2325 260 2425
rect 295 2325 300 2425
rect 200 2310 300 2325
rect 450 2425 550 2440
rect 450 2325 455 2425
rect 490 2325 510 2425
rect 545 2325 550 2425
rect 450 2310 550 2325
rect 700 2425 800 2440
rect 700 2325 705 2425
rect 740 2325 760 2425
rect 795 2325 800 2425
rect 700 2310 800 2325
rect 950 2425 1050 2440
rect 950 2325 955 2425
rect 990 2325 1010 2425
rect 1045 2325 1050 2425
rect 950 2310 1050 2325
rect 1200 2425 1300 2440
rect 1200 2325 1205 2425
rect 1240 2325 1260 2425
rect 1295 2325 1300 2425
rect 1200 2310 1300 2325
rect 1450 2425 1550 2440
rect 1450 2325 1455 2425
rect 1490 2325 1510 2425
rect 1545 2325 1550 2425
rect 1450 2310 1550 2325
rect 1700 2425 1800 2440
rect 1700 2325 1705 2425
rect 1740 2325 1760 2425
rect 1795 2325 1800 2425
rect 1700 2310 1800 2325
rect 1950 2425 2050 2440
rect 1950 2325 1955 2425
rect 1990 2325 2010 2425
rect 2045 2325 2050 2425
rect 1950 2310 2050 2325
rect 2200 2425 2300 2440
rect 2200 2325 2205 2425
rect 2240 2325 2260 2425
rect 2295 2325 2300 2425
rect 2200 2310 2300 2325
rect 2450 2425 2550 2440
rect 2450 2325 2455 2425
rect 2490 2325 2510 2425
rect 2545 2325 2550 2425
rect 2450 2310 2550 2325
rect 2700 2425 2800 2440
rect 2700 2325 2705 2425
rect 2740 2325 2760 2425
rect 2795 2325 2800 2425
rect 2700 2310 2800 2325
rect 2950 2425 3050 2440
rect 2950 2325 2955 2425
rect 2990 2325 3010 2425
rect 3045 2325 3050 2425
rect 2950 2310 3050 2325
rect 3200 2425 3300 2440
rect 3200 2325 3205 2425
rect 3240 2325 3260 2425
rect 3295 2325 3300 2425
rect 3200 2310 3300 2325
rect 3450 2425 3550 2440
rect 3450 2325 3455 2425
rect 3490 2325 3510 2425
rect 3545 2325 3550 2425
rect 3450 2310 3550 2325
rect 3700 2425 3800 2440
rect 3700 2325 3705 2425
rect 3740 2325 3760 2425
rect 3795 2325 3800 2425
rect 3700 2310 3800 2325
rect 3950 2425 4050 2440
rect 3950 2325 3955 2425
rect 3990 2325 4010 2425
rect 4045 2325 4050 2425
rect 3950 2310 4050 2325
rect 4200 2425 4300 2440
rect 4200 2325 4205 2425
rect 4240 2325 4260 2425
rect 4295 2325 4300 2425
rect 4200 2310 4300 2325
rect 4450 2425 4550 2440
rect 4450 2325 4455 2425
rect 4490 2325 4510 2425
rect 4545 2325 4550 2425
rect 4450 2310 4550 2325
rect 4700 2425 4800 2440
rect 4700 2325 4705 2425
rect 4740 2325 4760 2425
rect 4795 2325 4800 2425
rect 4700 2310 4800 2325
rect 4950 2425 5050 2440
rect 4950 2325 4955 2425
rect 4990 2325 5010 2425
rect 5045 2325 5050 2425
rect 4950 2310 5050 2325
rect 5200 2425 5300 2440
rect 5200 2325 5205 2425
rect 5240 2325 5260 2425
rect 5295 2325 5300 2425
rect 5200 2310 5300 2325
rect 5450 2425 5550 2440
rect 5450 2325 5455 2425
rect 5490 2325 5510 2425
rect 5545 2325 5550 2425
rect 5450 2310 5550 2325
rect 5700 2425 5800 2440
rect 5700 2325 5705 2425
rect 5740 2325 5760 2425
rect 5795 2325 5800 2425
rect 5700 2310 5800 2325
rect 5950 2425 6050 2440
rect 5950 2325 5955 2425
rect 5990 2325 6010 2425
rect 6045 2325 6050 2425
rect 5950 2310 6050 2325
rect 6200 2425 6300 2440
rect 6200 2325 6205 2425
rect 6240 2325 6260 2425
rect 6295 2325 6300 2425
rect 6200 2310 6300 2325
rect 6450 2425 6550 2440
rect 6450 2325 6455 2425
rect 6490 2325 6510 2425
rect 6545 2325 6550 2425
rect 6450 2310 6550 2325
rect 6700 2425 6800 2440
rect 6700 2325 6705 2425
rect 6740 2325 6760 2425
rect 6795 2325 6800 2425
rect 6700 2310 6800 2325
rect 6950 2425 7050 2440
rect 6950 2325 6955 2425
rect 6990 2325 7010 2425
rect 7045 2325 7050 2425
rect 6950 2310 7050 2325
rect 7200 2425 7300 2440
rect 7200 2325 7205 2425
rect 7240 2325 7260 2425
rect 7295 2325 7300 2425
rect 7200 2310 7300 2325
rect 7450 2425 7550 2440
rect 7450 2325 7455 2425
rect 7490 2325 7510 2425
rect 7545 2325 7550 2425
rect 7450 2310 7550 2325
rect 7700 2425 7800 2440
rect 7700 2325 7705 2425
rect 7740 2325 7760 2425
rect 7795 2325 7800 2425
rect 7700 2310 7800 2325
rect 7950 2425 8000 2440
rect 7950 2325 7955 2425
rect 7990 2325 8000 2425
rect 7950 2310 8000 2325
rect 0 2300 60 2310
rect 190 2300 310 2310
rect 440 2300 560 2310
rect 690 2300 810 2310
rect 940 2300 1060 2310
rect 1190 2300 1310 2310
rect 1440 2300 1560 2310
rect 1690 2300 1810 2310
rect 1940 2300 2060 2310
rect 2190 2300 2310 2310
rect 2440 2300 2560 2310
rect 2690 2300 2810 2310
rect 2940 2300 3060 2310
rect 3190 2300 3310 2310
rect 3440 2300 3560 2310
rect 3690 2300 3810 2310
rect 3940 2300 4060 2310
rect 4190 2300 4310 2310
rect 4440 2300 4560 2310
rect 4690 2300 4810 2310
rect 4940 2300 5060 2310
rect 5190 2300 5310 2310
rect 5440 2300 5560 2310
rect 5690 2300 5810 2310
rect 5940 2300 6060 2310
rect 6190 2300 6310 2310
rect 6440 2300 6560 2310
rect 6690 2300 6810 2310
rect 6940 2300 7060 2310
rect 7190 2300 7310 2310
rect 7440 2300 7560 2310
rect 7690 2300 7810 2310
rect 7940 2300 8000 2310
rect 0 2295 200 2300
rect 0 2260 75 2295
rect 175 2260 200 2295
rect 0 2240 200 2260
rect 0 2205 75 2240
rect 175 2205 200 2240
rect 0 2200 200 2205
rect 300 2295 450 2300
rect 300 2260 325 2295
rect 425 2260 450 2295
rect 300 2240 450 2260
rect 300 2205 325 2240
rect 425 2205 450 2240
rect 300 2200 450 2205
rect 550 2295 700 2300
rect 550 2260 575 2295
rect 675 2260 700 2295
rect 550 2240 700 2260
rect 550 2205 575 2240
rect 675 2205 700 2240
rect 550 2200 700 2205
rect 800 2295 1200 2300
rect 800 2260 825 2295
rect 925 2260 1075 2295
rect 1175 2260 1200 2295
rect 800 2240 1200 2260
rect 800 2205 825 2240
rect 925 2205 1075 2240
rect 1175 2205 1200 2240
rect 800 2200 1200 2205
rect 1300 2295 1450 2300
rect 1300 2260 1325 2295
rect 1425 2260 1450 2295
rect 1300 2240 1450 2260
rect 1300 2205 1325 2240
rect 1425 2205 1450 2240
rect 1300 2200 1450 2205
rect 1550 2295 1700 2300
rect 1550 2260 1575 2295
rect 1675 2260 1700 2295
rect 1550 2240 1700 2260
rect 1550 2205 1575 2240
rect 1675 2205 1700 2240
rect 1550 2200 1700 2205
rect 1800 2295 2200 2300
rect 1800 2260 1825 2295
rect 1925 2260 2075 2295
rect 2175 2260 2200 2295
rect 1800 2240 2200 2260
rect 1800 2205 1825 2240
rect 1925 2205 2075 2240
rect 2175 2205 2200 2240
rect 1800 2200 2200 2205
rect 2300 2295 2450 2300
rect 2300 2260 2325 2295
rect 2425 2260 2450 2295
rect 2300 2240 2450 2260
rect 2300 2205 2325 2240
rect 2425 2205 2450 2240
rect 2300 2200 2450 2205
rect 2550 2295 2700 2300
rect 2550 2260 2575 2295
rect 2675 2260 2700 2295
rect 2550 2240 2700 2260
rect 2550 2205 2575 2240
rect 2675 2205 2700 2240
rect 2550 2200 2700 2205
rect 2800 2295 3200 2300
rect 2800 2260 2825 2295
rect 2925 2260 3075 2295
rect 3175 2260 3200 2295
rect 2800 2240 3200 2260
rect 2800 2205 2825 2240
rect 2925 2205 3075 2240
rect 3175 2205 3200 2240
rect 2800 2200 3200 2205
rect 3300 2295 3450 2300
rect 3300 2260 3325 2295
rect 3425 2260 3450 2295
rect 3300 2240 3450 2260
rect 3300 2205 3325 2240
rect 3425 2205 3450 2240
rect 3300 2200 3450 2205
rect 3550 2295 3700 2300
rect 3550 2260 3575 2295
rect 3675 2260 3700 2295
rect 3550 2240 3700 2260
rect 3550 2205 3575 2240
rect 3675 2205 3700 2240
rect 3550 2200 3700 2205
rect 3800 2295 4200 2300
rect 3800 2260 3825 2295
rect 3925 2260 4075 2295
rect 4175 2260 4200 2295
rect 3800 2240 4200 2260
rect 3800 2205 3825 2240
rect 3925 2205 4075 2240
rect 4175 2205 4200 2240
rect 3800 2200 4200 2205
rect 4300 2295 4450 2300
rect 4300 2260 4325 2295
rect 4425 2260 4450 2295
rect 4300 2240 4450 2260
rect 4300 2205 4325 2240
rect 4425 2205 4450 2240
rect 4300 2200 4450 2205
rect 4550 2295 4700 2300
rect 4550 2260 4575 2295
rect 4675 2260 4700 2295
rect 4550 2240 4700 2260
rect 4550 2205 4575 2240
rect 4675 2205 4700 2240
rect 4550 2200 4700 2205
rect 4800 2295 5200 2300
rect 4800 2260 4825 2295
rect 4925 2260 5075 2295
rect 5175 2260 5200 2295
rect 4800 2240 5200 2260
rect 4800 2205 4825 2240
rect 4925 2205 5075 2240
rect 5175 2205 5200 2240
rect 4800 2200 5200 2205
rect 5300 2295 5450 2300
rect 5300 2260 5325 2295
rect 5425 2260 5450 2295
rect 5300 2240 5450 2260
rect 5300 2205 5325 2240
rect 5425 2205 5450 2240
rect 5300 2200 5450 2205
rect 5550 2295 5700 2300
rect 5550 2260 5575 2295
rect 5675 2260 5700 2295
rect 5550 2240 5700 2260
rect 5550 2205 5575 2240
rect 5675 2205 5700 2240
rect 5550 2200 5700 2205
rect 5800 2295 6200 2300
rect 5800 2260 5825 2295
rect 5925 2260 6075 2295
rect 6175 2260 6200 2295
rect 5800 2240 6200 2260
rect 5800 2205 5825 2240
rect 5925 2205 6075 2240
rect 6175 2205 6200 2240
rect 5800 2200 6200 2205
rect 6300 2295 6450 2300
rect 6300 2260 6325 2295
rect 6425 2260 6450 2295
rect 6300 2240 6450 2260
rect 6300 2205 6325 2240
rect 6425 2205 6450 2240
rect 6300 2200 6450 2205
rect 6550 2295 6700 2300
rect 6550 2260 6575 2295
rect 6675 2260 6700 2295
rect 6550 2240 6700 2260
rect 6550 2205 6575 2240
rect 6675 2205 6700 2240
rect 6550 2200 6700 2205
rect 6800 2295 7200 2300
rect 6800 2260 6825 2295
rect 6925 2260 7075 2295
rect 7175 2260 7200 2295
rect 6800 2240 7200 2260
rect 6800 2205 6825 2240
rect 6925 2205 7075 2240
rect 7175 2205 7200 2240
rect 6800 2200 7200 2205
rect 7300 2295 7450 2300
rect 7300 2260 7325 2295
rect 7425 2260 7450 2295
rect 7300 2240 7450 2260
rect 7300 2205 7325 2240
rect 7425 2205 7450 2240
rect 7300 2200 7450 2205
rect 7550 2295 7700 2300
rect 7550 2260 7575 2295
rect 7675 2260 7700 2295
rect 7550 2240 7700 2260
rect 7550 2205 7575 2240
rect 7675 2205 7700 2240
rect 7550 2200 7700 2205
rect 7800 2295 8000 2300
rect 7800 2260 7825 2295
rect 7925 2260 8000 2295
rect 7800 2240 8000 2260
rect 7800 2205 7825 2240
rect 7925 2205 8000 2240
rect 7800 2200 8000 2205
rect 0 2190 60 2200
rect 190 2190 310 2200
rect 440 2190 560 2200
rect 690 2190 810 2200
rect 940 2190 1060 2200
rect 1190 2190 1310 2200
rect 1440 2190 1560 2200
rect 1690 2190 1810 2200
rect 1940 2190 2060 2200
rect 2190 2190 2310 2200
rect 2440 2190 2560 2200
rect 2690 2190 2810 2200
rect 2940 2190 3060 2200
rect 3190 2190 3310 2200
rect 3440 2190 3560 2200
rect 3690 2190 3810 2200
rect 3940 2190 4060 2200
rect 4190 2190 4310 2200
rect 4440 2190 4560 2200
rect 4690 2190 4810 2200
rect 4940 2190 5060 2200
rect 5190 2190 5310 2200
rect 5440 2190 5560 2200
rect 5690 2190 5810 2200
rect 5940 2190 6060 2200
rect 6190 2190 6310 2200
rect 6440 2190 6560 2200
rect 6690 2190 6810 2200
rect 6940 2190 7060 2200
rect 7190 2190 7310 2200
rect 7440 2190 7560 2200
rect 7690 2190 7810 2200
rect 7940 2190 8000 2200
rect 0 2175 50 2190
rect 0 2075 10 2175
rect 45 2075 50 2175
rect 0 2060 50 2075
rect 200 2175 300 2190
rect 200 2075 205 2175
rect 240 2075 260 2175
rect 295 2075 300 2175
rect 200 2060 300 2075
rect 450 2175 550 2190
rect 450 2075 455 2175
rect 490 2075 510 2175
rect 545 2075 550 2175
rect 450 2060 550 2075
rect 700 2175 800 2190
rect 700 2075 705 2175
rect 740 2075 760 2175
rect 795 2075 800 2175
rect 700 2060 800 2075
rect 950 2175 1050 2190
rect 950 2075 955 2175
rect 990 2075 1010 2175
rect 1045 2075 1050 2175
rect 950 2060 1050 2075
rect 1200 2175 1300 2190
rect 1200 2075 1205 2175
rect 1240 2075 1260 2175
rect 1295 2075 1300 2175
rect 1200 2060 1300 2075
rect 1450 2175 1550 2190
rect 1450 2075 1455 2175
rect 1490 2075 1510 2175
rect 1545 2075 1550 2175
rect 1450 2060 1550 2075
rect 1700 2175 1800 2190
rect 1700 2075 1705 2175
rect 1740 2075 1760 2175
rect 1795 2075 1800 2175
rect 1700 2060 1800 2075
rect 1950 2175 2050 2190
rect 1950 2075 1955 2175
rect 1990 2075 2010 2175
rect 2045 2075 2050 2175
rect 1950 2060 2050 2075
rect 2200 2175 2300 2190
rect 2200 2075 2205 2175
rect 2240 2075 2260 2175
rect 2295 2075 2300 2175
rect 2200 2060 2300 2075
rect 2450 2175 2550 2190
rect 2450 2075 2455 2175
rect 2490 2075 2510 2175
rect 2545 2075 2550 2175
rect 2450 2060 2550 2075
rect 2700 2175 2800 2190
rect 2700 2075 2705 2175
rect 2740 2075 2760 2175
rect 2795 2075 2800 2175
rect 2700 2060 2800 2075
rect 2950 2175 3050 2190
rect 2950 2075 2955 2175
rect 2990 2075 3010 2175
rect 3045 2075 3050 2175
rect 2950 2060 3050 2075
rect 3200 2175 3300 2190
rect 3200 2075 3205 2175
rect 3240 2075 3260 2175
rect 3295 2075 3300 2175
rect 3200 2060 3300 2075
rect 3450 2175 3550 2190
rect 3450 2075 3455 2175
rect 3490 2075 3510 2175
rect 3545 2075 3550 2175
rect 3450 2060 3550 2075
rect 3700 2175 3800 2190
rect 3700 2075 3705 2175
rect 3740 2075 3760 2175
rect 3795 2075 3800 2175
rect 3700 2060 3800 2075
rect 3950 2175 4050 2190
rect 3950 2075 3955 2175
rect 3990 2075 4010 2175
rect 4045 2075 4050 2175
rect 3950 2060 4050 2075
rect 4200 2175 4300 2190
rect 4200 2075 4205 2175
rect 4240 2075 4260 2175
rect 4295 2075 4300 2175
rect 4200 2060 4300 2075
rect 4450 2175 4550 2190
rect 4450 2075 4455 2175
rect 4490 2075 4510 2175
rect 4545 2075 4550 2175
rect 4450 2060 4550 2075
rect 4700 2175 4800 2190
rect 4700 2075 4705 2175
rect 4740 2075 4760 2175
rect 4795 2075 4800 2175
rect 4700 2060 4800 2075
rect 4950 2175 5050 2190
rect 4950 2075 4955 2175
rect 4990 2075 5010 2175
rect 5045 2075 5050 2175
rect 4950 2060 5050 2075
rect 5200 2175 5300 2190
rect 5200 2075 5205 2175
rect 5240 2075 5260 2175
rect 5295 2075 5300 2175
rect 5200 2060 5300 2075
rect 5450 2175 5550 2190
rect 5450 2075 5455 2175
rect 5490 2075 5510 2175
rect 5545 2075 5550 2175
rect 5450 2060 5550 2075
rect 5700 2175 5800 2190
rect 5700 2075 5705 2175
rect 5740 2075 5760 2175
rect 5795 2075 5800 2175
rect 5700 2060 5800 2075
rect 5950 2175 6050 2190
rect 5950 2075 5955 2175
rect 5990 2075 6010 2175
rect 6045 2075 6050 2175
rect 5950 2060 6050 2075
rect 6200 2175 6300 2190
rect 6200 2075 6205 2175
rect 6240 2075 6260 2175
rect 6295 2075 6300 2175
rect 6200 2060 6300 2075
rect 6450 2175 6550 2190
rect 6450 2075 6455 2175
rect 6490 2075 6510 2175
rect 6545 2075 6550 2175
rect 6450 2060 6550 2075
rect 6700 2175 6800 2190
rect 6700 2075 6705 2175
rect 6740 2075 6760 2175
rect 6795 2075 6800 2175
rect 6700 2060 6800 2075
rect 6950 2175 7050 2190
rect 6950 2075 6955 2175
rect 6990 2075 7010 2175
rect 7045 2075 7050 2175
rect 6950 2060 7050 2075
rect 7200 2175 7300 2190
rect 7200 2075 7205 2175
rect 7240 2075 7260 2175
rect 7295 2075 7300 2175
rect 7200 2060 7300 2075
rect 7450 2175 7550 2190
rect 7450 2075 7455 2175
rect 7490 2075 7510 2175
rect 7545 2075 7550 2175
rect 7450 2060 7550 2075
rect 7700 2175 7800 2190
rect 7700 2075 7705 2175
rect 7740 2075 7760 2175
rect 7795 2075 7800 2175
rect 7700 2060 7800 2075
rect 7950 2175 8000 2190
rect 7950 2075 7955 2175
rect 7990 2075 8000 2175
rect 7950 2060 8000 2075
rect 0 2050 60 2060
rect 190 2050 310 2060
rect 440 2050 560 2060
rect 690 2050 810 2060
rect 940 2050 1060 2060
rect 1190 2050 1310 2060
rect 1440 2050 1560 2060
rect 1690 2050 1810 2060
rect 1940 2050 2060 2060
rect 2190 2050 2310 2060
rect 2440 2050 2560 2060
rect 2690 2050 2810 2060
rect 2940 2050 3060 2060
rect 3190 2050 3310 2060
rect 3440 2050 3560 2060
rect 3690 2050 3810 2060
rect 3940 2050 4060 2060
rect 4190 2050 4310 2060
rect 4440 2050 4560 2060
rect 4690 2050 4810 2060
rect 4940 2050 5060 2060
rect 5190 2050 5310 2060
rect 5440 2050 5560 2060
rect 5690 2050 5810 2060
rect 5940 2050 6060 2060
rect 6190 2050 6310 2060
rect 6440 2050 6560 2060
rect 6690 2050 6810 2060
rect 6940 2050 7060 2060
rect 7190 2050 7310 2060
rect 7440 2050 7560 2060
rect 7690 2050 7810 2060
rect 7940 2050 8000 2060
rect 0 2045 8000 2050
rect 0 2010 75 2045
rect 175 2010 325 2045
rect 425 2010 575 2045
rect 675 2010 825 2045
rect 925 2010 1075 2045
rect 1175 2010 1325 2045
rect 1425 2010 1575 2045
rect 1675 2010 1825 2045
rect 1925 2010 2075 2045
rect 2175 2010 2325 2045
rect 2425 2010 2575 2045
rect 2675 2010 2825 2045
rect 2925 2010 3075 2045
rect 3175 2010 3325 2045
rect 3425 2010 3575 2045
rect 3675 2010 3825 2045
rect 3925 2010 4075 2045
rect 4175 2010 4325 2045
rect 4425 2010 4575 2045
rect 4675 2010 4825 2045
rect 4925 2010 5075 2045
rect 5175 2010 5325 2045
rect 5425 2010 5575 2045
rect 5675 2010 5825 2045
rect 5925 2010 6075 2045
rect 6175 2010 6325 2045
rect 6425 2010 6575 2045
rect 6675 2010 6825 2045
rect 6925 2010 7075 2045
rect 7175 2010 7325 2045
rect 7425 2010 7575 2045
rect 7675 2010 7825 2045
rect 7925 2010 8000 2045
rect 0 1990 8000 2010
rect 0 1955 75 1990
rect 175 1955 325 1990
rect 425 1955 575 1990
rect 675 1955 825 1990
rect 925 1955 1075 1990
rect 1175 1955 1325 1990
rect 1425 1955 1575 1990
rect 1675 1955 1825 1990
rect 1925 1955 2075 1990
rect 2175 1955 2325 1990
rect 2425 1955 2575 1990
rect 2675 1955 2825 1990
rect 2925 1955 3075 1990
rect 3175 1955 3325 1990
rect 3425 1955 3575 1990
rect 3675 1955 3825 1990
rect 3925 1955 4075 1990
rect 4175 1955 4325 1990
rect 4425 1955 4575 1990
rect 4675 1955 4825 1990
rect 4925 1955 5075 1990
rect 5175 1955 5325 1990
rect 5425 1955 5575 1990
rect 5675 1955 5825 1990
rect 5925 1955 6075 1990
rect 6175 1955 6325 1990
rect 6425 1955 6575 1990
rect 6675 1955 6825 1990
rect 6925 1955 7075 1990
rect 7175 1955 7325 1990
rect 7425 1955 7575 1990
rect 7675 1955 7825 1990
rect 7925 1955 8000 1990
rect 0 1950 8000 1955
rect 0 1940 60 1950
rect 190 1940 310 1950
rect 440 1940 560 1950
rect 690 1940 810 1950
rect 940 1940 1060 1950
rect 1190 1940 1310 1950
rect 1440 1940 1560 1950
rect 1690 1940 1810 1950
rect 1940 1940 2060 1950
rect 2190 1940 2310 1950
rect 2440 1940 2560 1950
rect 2690 1940 2810 1950
rect 2940 1940 3060 1950
rect 3190 1940 3310 1950
rect 3440 1940 3560 1950
rect 3690 1940 3810 1950
rect 3940 1940 4060 1950
rect 4190 1940 4310 1950
rect 4440 1940 4560 1950
rect 4690 1940 4810 1950
rect 4940 1940 5060 1950
rect 5190 1940 5310 1950
rect 5440 1940 5560 1950
rect 5690 1940 5810 1950
rect 5940 1940 6060 1950
rect 6190 1940 6310 1950
rect 6440 1940 6560 1950
rect 6690 1940 6810 1950
rect 6940 1940 7060 1950
rect 7190 1940 7310 1950
rect 7440 1940 7560 1950
rect 7690 1940 7810 1950
rect 7940 1940 8000 1950
rect 0 1925 50 1940
rect 0 1825 10 1925
rect 45 1825 50 1925
rect 0 1810 50 1825
rect 200 1925 300 1940
rect 200 1825 205 1925
rect 240 1825 260 1925
rect 295 1825 300 1925
rect 200 1810 300 1825
rect 450 1925 550 1940
rect 450 1825 455 1925
rect 490 1825 510 1925
rect 545 1825 550 1925
rect 450 1810 550 1825
rect 700 1925 800 1940
rect 700 1825 705 1925
rect 740 1825 760 1925
rect 795 1825 800 1925
rect 700 1810 800 1825
rect 950 1925 1050 1940
rect 950 1825 955 1925
rect 990 1825 1010 1925
rect 1045 1825 1050 1925
rect 950 1810 1050 1825
rect 1200 1925 1300 1940
rect 1200 1825 1205 1925
rect 1240 1825 1260 1925
rect 1295 1825 1300 1925
rect 1200 1810 1300 1825
rect 1450 1925 1550 1940
rect 1450 1825 1455 1925
rect 1490 1825 1510 1925
rect 1545 1825 1550 1925
rect 1450 1810 1550 1825
rect 1700 1925 1800 1940
rect 1700 1825 1705 1925
rect 1740 1825 1760 1925
rect 1795 1825 1800 1925
rect 1700 1810 1800 1825
rect 1950 1925 2050 1940
rect 1950 1825 1955 1925
rect 1990 1825 2010 1925
rect 2045 1825 2050 1925
rect 1950 1810 2050 1825
rect 2200 1925 2300 1940
rect 2200 1825 2205 1925
rect 2240 1825 2260 1925
rect 2295 1825 2300 1925
rect 2200 1810 2300 1825
rect 2450 1925 2550 1940
rect 2450 1825 2455 1925
rect 2490 1825 2510 1925
rect 2545 1825 2550 1925
rect 2450 1810 2550 1825
rect 2700 1925 2800 1940
rect 2700 1825 2705 1925
rect 2740 1825 2760 1925
rect 2795 1825 2800 1925
rect 2700 1810 2800 1825
rect 2950 1925 3050 1940
rect 2950 1825 2955 1925
rect 2990 1825 3010 1925
rect 3045 1825 3050 1925
rect 2950 1810 3050 1825
rect 3200 1925 3300 1940
rect 3200 1825 3205 1925
rect 3240 1825 3260 1925
rect 3295 1825 3300 1925
rect 3200 1810 3300 1825
rect 3450 1925 3550 1940
rect 3450 1825 3455 1925
rect 3490 1825 3510 1925
rect 3545 1825 3550 1925
rect 3450 1810 3550 1825
rect 3700 1925 3800 1940
rect 3700 1825 3705 1925
rect 3740 1825 3760 1925
rect 3795 1825 3800 1925
rect 3700 1810 3800 1825
rect 3950 1925 4050 1940
rect 3950 1825 3955 1925
rect 3990 1825 4010 1925
rect 4045 1825 4050 1925
rect 3950 1810 4050 1825
rect 4200 1925 4300 1940
rect 4200 1825 4205 1925
rect 4240 1825 4260 1925
rect 4295 1825 4300 1925
rect 4200 1810 4300 1825
rect 4450 1925 4550 1940
rect 4450 1825 4455 1925
rect 4490 1825 4510 1925
rect 4545 1825 4550 1925
rect 4450 1810 4550 1825
rect 4700 1925 4800 1940
rect 4700 1825 4705 1925
rect 4740 1825 4760 1925
rect 4795 1825 4800 1925
rect 4700 1810 4800 1825
rect 4950 1925 5050 1940
rect 4950 1825 4955 1925
rect 4990 1825 5010 1925
rect 5045 1825 5050 1925
rect 4950 1810 5050 1825
rect 5200 1925 5300 1940
rect 5200 1825 5205 1925
rect 5240 1825 5260 1925
rect 5295 1825 5300 1925
rect 5200 1810 5300 1825
rect 5450 1925 5550 1940
rect 5450 1825 5455 1925
rect 5490 1825 5510 1925
rect 5545 1825 5550 1925
rect 5450 1810 5550 1825
rect 5700 1925 5800 1940
rect 5700 1825 5705 1925
rect 5740 1825 5760 1925
rect 5795 1825 5800 1925
rect 5700 1810 5800 1825
rect 5950 1925 6050 1940
rect 5950 1825 5955 1925
rect 5990 1825 6010 1925
rect 6045 1825 6050 1925
rect 5950 1810 6050 1825
rect 6200 1925 6300 1940
rect 6200 1825 6205 1925
rect 6240 1825 6260 1925
rect 6295 1825 6300 1925
rect 6200 1810 6300 1825
rect 6450 1925 6550 1940
rect 6450 1825 6455 1925
rect 6490 1825 6510 1925
rect 6545 1825 6550 1925
rect 6450 1810 6550 1825
rect 6700 1925 6800 1940
rect 6700 1825 6705 1925
rect 6740 1825 6760 1925
rect 6795 1825 6800 1925
rect 6700 1810 6800 1825
rect 6950 1925 7050 1940
rect 6950 1825 6955 1925
rect 6990 1825 7010 1925
rect 7045 1825 7050 1925
rect 6950 1810 7050 1825
rect 7200 1925 7300 1940
rect 7200 1825 7205 1925
rect 7240 1825 7260 1925
rect 7295 1825 7300 1925
rect 7200 1810 7300 1825
rect 7450 1925 7550 1940
rect 7450 1825 7455 1925
rect 7490 1825 7510 1925
rect 7545 1825 7550 1925
rect 7450 1810 7550 1825
rect 7700 1925 7800 1940
rect 7700 1825 7705 1925
rect 7740 1825 7760 1925
rect 7795 1825 7800 1925
rect 7700 1810 7800 1825
rect 7950 1925 8000 1940
rect 7950 1825 7955 1925
rect 7990 1825 8000 1925
rect 7950 1810 8000 1825
rect 0 1800 60 1810
rect 190 1800 310 1810
rect 440 1800 560 1810
rect 690 1800 810 1810
rect 940 1800 1060 1810
rect 1190 1800 1310 1810
rect 1440 1800 1560 1810
rect 1690 1800 1810 1810
rect 1940 1800 2060 1810
rect 2190 1800 2310 1810
rect 2440 1800 2560 1810
rect 2690 1800 2810 1810
rect 2940 1800 3060 1810
rect 3190 1800 3310 1810
rect 3440 1800 3560 1810
rect 3690 1800 3810 1810
rect 3940 1800 4060 1810
rect 4190 1800 4310 1810
rect 4440 1800 4560 1810
rect 4690 1800 4810 1810
rect 4940 1800 5060 1810
rect 5190 1800 5310 1810
rect 5440 1800 5560 1810
rect 5690 1800 5810 1810
rect 5940 1800 6060 1810
rect 6190 1800 6310 1810
rect 6440 1800 6560 1810
rect 6690 1800 6810 1810
rect 6940 1800 7060 1810
rect 7190 1800 7310 1810
rect 7440 1800 7560 1810
rect 7690 1800 7810 1810
rect 7940 1800 8000 1810
rect 0 1795 200 1800
rect 0 1760 75 1795
rect 175 1760 200 1795
rect 0 1740 200 1760
rect 0 1705 75 1740
rect 175 1705 200 1740
rect 0 1700 200 1705
rect 300 1795 450 1800
rect 300 1760 325 1795
rect 425 1760 450 1795
rect 300 1740 450 1760
rect 300 1705 325 1740
rect 425 1705 450 1740
rect 300 1700 450 1705
rect 550 1795 700 1800
rect 550 1760 575 1795
rect 675 1760 700 1795
rect 550 1740 700 1760
rect 550 1705 575 1740
rect 675 1705 700 1740
rect 550 1700 700 1705
rect 800 1795 1200 1800
rect 800 1760 825 1795
rect 925 1760 1075 1795
rect 1175 1760 1200 1795
rect 800 1740 1200 1760
rect 800 1705 825 1740
rect 925 1705 1075 1740
rect 1175 1705 1200 1740
rect 800 1700 1200 1705
rect 1300 1795 1450 1800
rect 1300 1760 1325 1795
rect 1425 1760 1450 1795
rect 1300 1740 1450 1760
rect 1300 1705 1325 1740
rect 1425 1705 1450 1740
rect 1300 1700 1450 1705
rect 1550 1795 1700 1800
rect 1550 1760 1575 1795
rect 1675 1760 1700 1795
rect 1550 1740 1700 1760
rect 1550 1705 1575 1740
rect 1675 1705 1700 1740
rect 1550 1700 1700 1705
rect 1800 1795 2200 1800
rect 1800 1760 1825 1795
rect 1925 1760 2075 1795
rect 2175 1760 2200 1795
rect 1800 1740 2200 1760
rect 1800 1705 1825 1740
rect 1925 1705 2075 1740
rect 2175 1705 2200 1740
rect 1800 1700 2200 1705
rect 2300 1795 2450 1800
rect 2300 1760 2325 1795
rect 2425 1760 2450 1795
rect 2300 1740 2450 1760
rect 2300 1705 2325 1740
rect 2425 1705 2450 1740
rect 2300 1700 2450 1705
rect 2550 1795 2700 1800
rect 2550 1760 2575 1795
rect 2675 1760 2700 1795
rect 2550 1740 2700 1760
rect 2550 1705 2575 1740
rect 2675 1705 2700 1740
rect 2550 1700 2700 1705
rect 2800 1795 3200 1800
rect 2800 1760 2825 1795
rect 2925 1760 3075 1795
rect 3175 1760 3200 1795
rect 2800 1740 3200 1760
rect 2800 1705 2825 1740
rect 2925 1705 3075 1740
rect 3175 1705 3200 1740
rect 2800 1700 3200 1705
rect 3300 1795 3450 1800
rect 3300 1760 3325 1795
rect 3425 1760 3450 1795
rect 3300 1740 3450 1760
rect 3300 1705 3325 1740
rect 3425 1705 3450 1740
rect 3300 1700 3450 1705
rect 3550 1795 3700 1800
rect 3550 1760 3575 1795
rect 3675 1760 3700 1795
rect 3550 1740 3700 1760
rect 3550 1705 3575 1740
rect 3675 1705 3700 1740
rect 3550 1700 3700 1705
rect 3800 1795 4200 1800
rect 3800 1760 3825 1795
rect 3925 1760 4075 1795
rect 4175 1760 4200 1795
rect 3800 1740 4200 1760
rect 3800 1705 3825 1740
rect 3925 1705 4075 1740
rect 4175 1705 4200 1740
rect 3800 1700 4200 1705
rect 4300 1795 4450 1800
rect 4300 1760 4325 1795
rect 4425 1760 4450 1795
rect 4300 1740 4450 1760
rect 4300 1705 4325 1740
rect 4425 1705 4450 1740
rect 4300 1700 4450 1705
rect 4550 1795 4700 1800
rect 4550 1760 4575 1795
rect 4675 1760 4700 1795
rect 4550 1740 4700 1760
rect 4550 1705 4575 1740
rect 4675 1705 4700 1740
rect 4550 1700 4700 1705
rect 4800 1795 5200 1800
rect 4800 1760 4825 1795
rect 4925 1760 5075 1795
rect 5175 1760 5200 1795
rect 4800 1740 5200 1760
rect 4800 1705 4825 1740
rect 4925 1705 5075 1740
rect 5175 1705 5200 1740
rect 4800 1700 5200 1705
rect 5300 1795 5450 1800
rect 5300 1760 5325 1795
rect 5425 1760 5450 1795
rect 5300 1740 5450 1760
rect 5300 1705 5325 1740
rect 5425 1705 5450 1740
rect 5300 1700 5450 1705
rect 5550 1795 5700 1800
rect 5550 1760 5575 1795
rect 5675 1760 5700 1795
rect 5550 1740 5700 1760
rect 5550 1705 5575 1740
rect 5675 1705 5700 1740
rect 5550 1700 5700 1705
rect 5800 1795 6200 1800
rect 5800 1760 5825 1795
rect 5925 1760 6075 1795
rect 6175 1760 6200 1795
rect 5800 1740 6200 1760
rect 5800 1705 5825 1740
rect 5925 1705 6075 1740
rect 6175 1705 6200 1740
rect 5800 1700 6200 1705
rect 6300 1795 6450 1800
rect 6300 1760 6325 1795
rect 6425 1760 6450 1795
rect 6300 1740 6450 1760
rect 6300 1705 6325 1740
rect 6425 1705 6450 1740
rect 6300 1700 6450 1705
rect 6550 1795 6700 1800
rect 6550 1760 6575 1795
rect 6675 1760 6700 1795
rect 6550 1740 6700 1760
rect 6550 1705 6575 1740
rect 6675 1705 6700 1740
rect 6550 1700 6700 1705
rect 6800 1795 7200 1800
rect 6800 1760 6825 1795
rect 6925 1760 7075 1795
rect 7175 1760 7200 1795
rect 6800 1740 7200 1760
rect 6800 1705 6825 1740
rect 6925 1705 7075 1740
rect 7175 1705 7200 1740
rect 6800 1700 7200 1705
rect 7300 1795 7450 1800
rect 7300 1760 7325 1795
rect 7425 1760 7450 1795
rect 7300 1740 7450 1760
rect 7300 1705 7325 1740
rect 7425 1705 7450 1740
rect 7300 1700 7450 1705
rect 7550 1795 7700 1800
rect 7550 1760 7575 1795
rect 7675 1760 7700 1795
rect 7550 1740 7700 1760
rect 7550 1705 7575 1740
rect 7675 1705 7700 1740
rect 7550 1700 7700 1705
rect 7800 1795 8000 1800
rect 7800 1760 7825 1795
rect 7925 1760 8000 1795
rect 7800 1740 8000 1760
rect 7800 1705 7825 1740
rect 7925 1705 8000 1740
rect 7800 1700 8000 1705
rect 0 1690 60 1700
rect 190 1690 310 1700
rect 440 1690 560 1700
rect 690 1690 810 1700
rect 940 1690 1060 1700
rect 1190 1690 1310 1700
rect 1440 1690 1560 1700
rect 1690 1690 1810 1700
rect 1940 1690 2060 1700
rect 2190 1690 2310 1700
rect 2440 1690 2560 1700
rect 2690 1690 2810 1700
rect 2940 1690 3060 1700
rect 3190 1690 3310 1700
rect 3440 1690 3560 1700
rect 3690 1690 3810 1700
rect 3940 1690 4060 1700
rect 4190 1690 4310 1700
rect 4440 1690 4560 1700
rect 4690 1690 4810 1700
rect 4940 1690 5060 1700
rect 5190 1690 5310 1700
rect 5440 1690 5560 1700
rect 5690 1690 5810 1700
rect 5940 1690 6060 1700
rect 6190 1690 6310 1700
rect 6440 1690 6560 1700
rect 6690 1690 6810 1700
rect 6940 1690 7060 1700
rect 7190 1690 7310 1700
rect 7440 1690 7560 1700
rect 7690 1690 7810 1700
rect 7940 1690 8000 1700
rect 0 1675 50 1690
rect 0 1575 10 1675
rect 45 1575 50 1675
rect 0 1560 50 1575
rect 200 1675 300 1690
rect 200 1575 205 1675
rect 240 1575 260 1675
rect 295 1575 300 1675
rect 200 1560 300 1575
rect 450 1675 550 1690
rect 450 1575 455 1675
rect 490 1575 510 1675
rect 545 1575 550 1675
rect 450 1560 550 1575
rect 700 1675 800 1690
rect 700 1575 705 1675
rect 740 1575 760 1675
rect 795 1575 800 1675
rect 700 1560 800 1575
rect 950 1675 1050 1690
rect 950 1575 955 1675
rect 990 1575 1010 1675
rect 1045 1575 1050 1675
rect 950 1560 1050 1575
rect 1200 1675 1300 1690
rect 1200 1575 1205 1675
rect 1240 1575 1260 1675
rect 1295 1575 1300 1675
rect 1200 1560 1300 1575
rect 1450 1675 1550 1690
rect 1450 1575 1455 1675
rect 1490 1575 1510 1675
rect 1545 1575 1550 1675
rect 1450 1560 1550 1575
rect 1700 1675 1800 1690
rect 1700 1575 1705 1675
rect 1740 1575 1760 1675
rect 1795 1575 1800 1675
rect 1700 1560 1800 1575
rect 1950 1675 2050 1690
rect 1950 1575 1955 1675
rect 1990 1575 2010 1675
rect 2045 1575 2050 1675
rect 1950 1560 2050 1575
rect 2200 1675 2300 1690
rect 2200 1575 2205 1675
rect 2240 1575 2260 1675
rect 2295 1575 2300 1675
rect 2200 1560 2300 1575
rect 2450 1675 2550 1690
rect 2450 1575 2455 1675
rect 2490 1575 2510 1675
rect 2545 1575 2550 1675
rect 2450 1560 2550 1575
rect 2700 1675 2800 1690
rect 2700 1575 2705 1675
rect 2740 1575 2760 1675
rect 2795 1575 2800 1675
rect 2700 1560 2800 1575
rect 2950 1675 3050 1690
rect 2950 1575 2955 1675
rect 2990 1575 3010 1675
rect 3045 1575 3050 1675
rect 2950 1560 3050 1575
rect 3200 1675 3300 1690
rect 3200 1575 3205 1675
rect 3240 1575 3260 1675
rect 3295 1575 3300 1675
rect 3200 1560 3300 1575
rect 3450 1675 3550 1690
rect 3450 1575 3455 1675
rect 3490 1575 3510 1675
rect 3545 1575 3550 1675
rect 3450 1560 3550 1575
rect 3700 1675 3800 1690
rect 3700 1575 3705 1675
rect 3740 1575 3760 1675
rect 3795 1575 3800 1675
rect 3700 1560 3800 1575
rect 3950 1675 4050 1690
rect 3950 1575 3955 1675
rect 3990 1575 4010 1675
rect 4045 1575 4050 1675
rect 3950 1560 4050 1575
rect 4200 1675 4300 1690
rect 4200 1575 4205 1675
rect 4240 1575 4260 1675
rect 4295 1575 4300 1675
rect 4200 1560 4300 1575
rect 4450 1675 4550 1690
rect 4450 1575 4455 1675
rect 4490 1575 4510 1675
rect 4545 1575 4550 1675
rect 4450 1560 4550 1575
rect 4700 1675 4800 1690
rect 4700 1575 4705 1675
rect 4740 1575 4760 1675
rect 4795 1575 4800 1675
rect 4700 1560 4800 1575
rect 4950 1675 5050 1690
rect 4950 1575 4955 1675
rect 4990 1575 5010 1675
rect 5045 1575 5050 1675
rect 4950 1560 5050 1575
rect 5200 1675 5300 1690
rect 5200 1575 5205 1675
rect 5240 1575 5260 1675
rect 5295 1575 5300 1675
rect 5200 1560 5300 1575
rect 5450 1675 5550 1690
rect 5450 1575 5455 1675
rect 5490 1575 5510 1675
rect 5545 1575 5550 1675
rect 5450 1560 5550 1575
rect 5700 1675 5800 1690
rect 5700 1575 5705 1675
rect 5740 1575 5760 1675
rect 5795 1575 5800 1675
rect 5700 1560 5800 1575
rect 5950 1675 6050 1690
rect 5950 1575 5955 1675
rect 5990 1575 6010 1675
rect 6045 1575 6050 1675
rect 5950 1560 6050 1575
rect 6200 1675 6300 1690
rect 6200 1575 6205 1675
rect 6240 1575 6260 1675
rect 6295 1575 6300 1675
rect 6200 1560 6300 1575
rect 6450 1675 6550 1690
rect 6450 1575 6455 1675
rect 6490 1575 6510 1675
rect 6545 1575 6550 1675
rect 6450 1560 6550 1575
rect 6700 1675 6800 1690
rect 6700 1575 6705 1675
rect 6740 1575 6760 1675
rect 6795 1575 6800 1675
rect 6700 1560 6800 1575
rect 6950 1675 7050 1690
rect 6950 1575 6955 1675
rect 6990 1575 7010 1675
rect 7045 1575 7050 1675
rect 6950 1560 7050 1575
rect 7200 1675 7300 1690
rect 7200 1575 7205 1675
rect 7240 1575 7260 1675
rect 7295 1575 7300 1675
rect 7200 1560 7300 1575
rect 7450 1675 7550 1690
rect 7450 1575 7455 1675
rect 7490 1575 7510 1675
rect 7545 1575 7550 1675
rect 7450 1560 7550 1575
rect 7700 1675 7800 1690
rect 7700 1575 7705 1675
rect 7740 1575 7760 1675
rect 7795 1575 7800 1675
rect 7700 1560 7800 1575
rect 7950 1675 8000 1690
rect 7950 1575 7955 1675
rect 7990 1575 8000 1675
rect 7950 1560 8000 1575
rect 0 1550 60 1560
rect 190 1550 310 1560
rect 440 1550 560 1560
rect 690 1550 810 1560
rect 940 1550 1060 1560
rect 1190 1550 1310 1560
rect 1440 1550 1560 1560
rect 1690 1550 1810 1560
rect 1940 1550 2060 1560
rect 2190 1550 2310 1560
rect 2440 1550 2560 1560
rect 2690 1550 2810 1560
rect 2940 1550 3060 1560
rect 3190 1550 3310 1560
rect 3440 1550 3560 1560
rect 3690 1550 3810 1560
rect 3940 1550 4060 1560
rect 4190 1550 4310 1560
rect 4440 1550 4560 1560
rect 4690 1550 4810 1560
rect 4940 1550 5060 1560
rect 5190 1550 5310 1560
rect 5440 1550 5560 1560
rect 5690 1550 5810 1560
rect 5940 1550 6060 1560
rect 6190 1550 6310 1560
rect 6440 1550 6560 1560
rect 6690 1550 6810 1560
rect 6940 1550 7060 1560
rect 7190 1550 7310 1560
rect 7440 1550 7560 1560
rect 7690 1550 7810 1560
rect 7940 1550 8000 1560
rect 0 1545 200 1550
rect 0 1510 75 1545
rect 175 1510 200 1545
rect 0 1490 200 1510
rect 0 1455 75 1490
rect 175 1455 200 1490
rect 0 1450 200 1455
rect 300 1545 450 1550
rect 300 1510 325 1545
rect 425 1510 450 1545
rect 300 1490 450 1510
rect 300 1455 325 1490
rect 425 1455 450 1490
rect 300 1450 450 1455
rect 550 1545 700 1550
rect 550 1510 575 1545
rect 675 1510 700 1545
rect 550 1490 700 1510
rect 550 1455 575 1490
rect 675 1455 700 1490
rect 550 1450 700 1455
rect 800 1545 950 1550
rect 800 1510 825 1545
rect 925 1510 950 1545
rect 800 1490 950 1510
rect 800 1455 825 1490
rect 925 1455 950 1490
rect 800 1450 950 1455
rect 1050 1545 1200 1550
rect 1050 1510 1075 1545
rect 1175 1510 1200 1545
rect 1050 1490 1200 1510
rect 1050 1455 1075 1490
rect 1175 1455 1200 1490
rect 1050 1450 1200 1455
rect 1300 1545 1450 1550
rect 1300 1510 1325 1545
rect 1425 1510 1450 1545
rect 1300 1490 1450 1510
rect 1300 1455 1325 1490
rect 1425 1455 1450 1490
rect 1300 1450 1450 1455
rect 1550 1545 1700 1550
rect 1550 1510 1575 1545
rect 1675 1510 1700 1545
rect 1550 1490 1700 1510
rect 1550 1455 1575 1490
rect 1675 1455 1700 1490
rect 1550 1450 1700 1455
rect 1800 1545 2200 1550
rect 1800 1510 1825 1545
rect 1925 1510 2075 1545
rect 2175 1510 2200 1545
rect 1800 1490 2200 1510
rect 1800 1455 1825 1490
rect 1925 1455 2075 1490
rect 2175 1455 2200 1490
rect 1800 1450 2200 1455
rect 2300 1545 2450 1550
rect 2300 1510 2325 1545
rect 2425 1510 2450 1545
rect 2300 1490 2450 1510
rect 2300 1455 2325 1490
rect 2425 1455 2450 1490
rect 2300 1450 2450 1455
rect 2550 1545 2700 1550
rect 2550 1510 2575 1545
rect 2675 1510 2700 1545
rect 2550 1490 2700 1510
rect 2550 1455 2575 1490
rect 2675 1455 2700 1490
rect 2550 1450 2700 1455
rect 2800 1545 2950 1550
rect 2800 1510 2825 1545
rect 2925 1510 2950 1545
rect 2800 1490 2950 1510
rect 2800 1455 2825 1490
rect 2925 1455 2950 1490
rect 2800 1450 2950 1455
rect 3050 1545 3200 1550
rect 3050 1510 3075 1545
rect 3175 1510 3200 1545
rect 3050 1490 3200 1510
rect 3050 1455 3075 1490
rect 3175 1455 3200 1490
rect 3050 1450 3200 1455
rect 3300 1545 3450 1550
rect 3300 1510 3325 1545
rect 3425 1510 3450 1545
rect 3300 1490 3450 1510
rect 3300 1455 3325 1490
rect 3425 1455 3450 1490
rect 3300 1450 3450 1455
rect 3550 1545 3700 1550
rect 3550 1510 3575 1545
rect 3675 1510 3700 1545
rect 3550 1490 3700 1510
rect 3550 1455 3575 1490
rect 3675 1455 3700 1490
rect 3550 1450 3700 1455
rect 3800 1545 4200 1550
rect 3800 1510 3825 1545
rect 3925 1510 4075 1545
rect 4175 1510 4200 1545
rect 3800 1490 4200 1510
rect 3800 1455 3825 1490
rect 3925 1455 4075 1490
rect 4175 1455 4200 1490
rect 3800 1450 4200 1455
rect 4300 1545 4450 1550
rect 4300 1510 4325 1545
rect 4425 1510 4450 1545
rect 4300 1490 4450 1510
rect 4300 1455 4325 1490
rect 4425 1455 4450 1490
rect 4300 1450 4450 1455
rect 4550 1545 4700 1550
rect 4550 1510 4575 1545
rect 4675 1510 4700 1545
rect 4550 1490 4700 1510
rect 4550 1455 4575 1490
rect 4675 1455 4700 1490
rect 4550 1450 4700 1455
rect 4800 1545 4950 1550
rect 4800 1510 4825 1545
rect 4925 1510 4950 1545
rect 4800 1490 4950 1510
rect 4800 1455 4825 1490
rect 4925 1455 4950 1490
rect 4800 1450 4950 1455
rect 5050 1545 5200 1550
rect 5050 1510 5075 1545
rect 5175 1510 5200 1545
rect 5050 1490 5200 1510
rect 5050 1455 5075 1490
rect 5175 1455 5200 1490
rect 5050 1450 5200 1455
rect 5300 1545 5450 1550
rect 5300 1510 5325 1545
rect 5425 1510 5450 1545
rect 5300 1490 5450 1510
rect 5300 1455 5325 1490
rect 5425 1455 5450 1490
rect 5300 1450 5450 1455
rect 5550 1545 5700 1550
rect 5550 1510 5575 1545
rect 5675 1510 5700 1545
rect 5550 1490 5700 1510
rect 5550 1455 5575 1490
rect 5675 1455 5700 1490
rect 5550 1450 5700 1455
rect 5800 1545 6200 1550
rect 5800 1510 5825 1545
rect 5925 1510 6075 1545
rect 6175 1510 6200 1545
rect 5800 1490 6200 1510
rect 5800 1455 5825 1490
rect 5925 1455 6075 1490
rect 6175 1455 6200 1490
rect 5800 1450 6200 1455
rect 6300 1545 6450 1550
rect 6300 1510 6325 1545
rect 6425 1510 6450 1545
rect 6300 1490 6450 1510
rect 6300 1455 6325 1490
rect 6425 1455 6450 1490
rect 6300 1450 6450 1455
rect 6550 1545 6700 1550
rect 6550 1510 6575 1545
rect 6675 1510 6700 1545
rect 6550 1490 6700 1510
rect 6550 1455 6575 1490
rect 6675 1455 6700 1490
rect 6550 1450 6700 1455
rect 6800 1545 6950 1550
rect 6800 1510 6825 1545
rect 6925 1510 6950 1545
rect 6800 1490 6950 1510
rect 6800 1455 6825 1490
rect 6925 1455 6950 1490
rect 6800 1450 6950 1455
rect 7050 1545 7200 1550
rect 7050 1510 7075 1545
rect 7175 1510 7200 1545
rect 7050 1490 7200 1510
rect 7050 1455 7075 1490
rect 7175 1455 7200 1490
rect 7050 1450 7200 1455
rect 7300 1545 7450 1550
rect 7300 1510 7325 1545
rect 7425 1510 7450 1545
rect 7300 1490 7450 1510
rect 7300 1455 7325 1490
rect 7425 1455 7450 1490
rect 7300 1450 7450 1455
rect 7550 1545 7700 1550
rect 7550 1510 7575 1545
rect 7675 1510 7700 1545
rect 7550 1490 7700 1510
rect 7550 1455 7575 1490
rect 7675 1455 7700 1490
rect 7550 1450 7700 1455
rect 7800 1545 8000 1550
rect 7800 1510 7825 1545
rect 7925 1510 8000 1545
rect 7800 1490 8000 1510
rect 7800 1455 7825 1490
rect 7925 1455 8000 1490
rect 7800 1450 8000 1455
rect 0 1440 60 1450
rect 190 1440 310 1450
rect 440 1440 560 1450
rect 690 1440 810 1450
rect 940 1440 1060 1450
rect 1190 1440 1310 1450
rect 1440 1440 1560 1450
rect 1690 1440 1810 1450
rect 1940 1440 2060 1450
rect 2190 1440 2310 1450
rect 2440 1440 2560 1450
rect 2690 1440 2810 1450
rect 2940 1440 3060 1450
rect 3190 1440 3310 1450
rect 3440 1440 3560 1450
rect 3690 1440 3810 1450
rect 3940 1440 4060 1450
rect 4190 1440 4310 1450
rect 4440 1440 4560 1450
rect 4690 1440 4810 1450
rect 4940 1440 5060 1450
rect 5190 1440 5310 1450
rect 5440 1440 5560 1450
rect 5690 1440 5810 1450
rect 5940 1440 6060 1450
rect 6190 1440 6310 1450
rect 6440 1440 6560 1450
rect 6690 1440 6810 1450
rect 6940 1440 7060 1450
rect 7190 1440 7310 1450
rect 7440 1440 7560 1450
rect 7690 1440 7810 1450
rect 7940 1440 8000 1450
rect 0 1425 50 1440
rect 0 1325 10 1425
rect 45 1325 50 1425
rect 0 1310 50 1325
rect 200 1425 300 1440
rect 200 1325 205 1425
rect 240 1325 260 1425
rect 295 1325 300 1425
rect 200 1310 300 1325
rect 450 1425 550 1440
rect 450 1325 455 1425
rect 490 1325 510 1425
rect 545 1325 550 1425
rect 450 1310 550 1325
rect 700 1425 800 1440
rect 700 1325 705 1425
rect 740 1325 760 1425
rect 795 1325 800 1425
rect 700 1310 800 1325
rect 950 1425 1050 1440
rect 950 1325 955 1425
rect 990 1325 1010 1425
rect 1045 1325 1050 1425
rect 950 1310 1050 1325
rect 1200 1425 1300 1440
rect 1200 1325 1205 1425
rect 1240 1325 1260 1425
rect 1295 1325 1300 1425
rect 1200 1310 1300 1325
rect 1450 1425 1550 1440
rect 1450 1325 1455 1425
rect 1490 1325 1510 1425
rect 1545 1325 1550 1425
rect 1450 1310 1550 1325
rect 1700 1425 1800 1440
rect 1700 1325 1705 1425
rect 1740 1325 1760 1425
rect 1795 1325 1800 1425
rect 1700 1310 1800 1325
rect 1950 1425 2050 1440
rect 1950 1325 1955 1425
rect 1990 1325 2010 1425
rect 2045 1325 2050 1425
rect 1950 1310 2050 1325
rect 2200 1425 2300 1440
rect 2200 1325 2205 1425
rect 2240 1325 2260 1425
rect 2295 1325 2300 1425
rect 2200 1310 2300 1325
rect 2450 1425 2550 1440
rect 2450 1325 2455 1425
rect 2490 1325 2510 1425
rect 2545 1325 2550 1425
rect 2450 1310 2550 1325
rect 2700 1425 2800 1440
rect 2700 1325 2705 1425
rect 2740 1325 2760 1425
rect 2795 1325 2800 1425
rect 2700 1310 2800 1325
rect 2950 1425 3050 1440
rect 2950 1325 2955 1425
rect 2990 1325 3010 1425
rect 3045 1325 3050 1425
rect 2950 1310 3050 1325
rect 3200 1425 3300 1440
rect 3200 1325 3205 1425
rect 3240 1325 3260 1425
rect 3295 1325 3300 1425
rect 3200 1310 3300 1325
rect 3450 1425 3550 1440
rect 3450 1325 3455 1425
rect 3490 1325 3510 1425
rect 3545 1325 3550 1425
rect 3450 1310 3550 1325
rect 3700 1425 3800 1440
rect 3700 1325 3705 1425
rect 3740 1325 3760 1425
rect 3795 1325 3800 1425
rect 3700 1310 3800 1325
rect 3950 1425 4050 1440
rect 3950 1325 3955 1425
rect 3990 1325 4010 1425
rect 4045 1325 4050 1425
rect 3950 1310 4050 1325
rect 4200 1425 4300 1440
rect 4200 1325 4205 1425
rect 4240 1325 4260 1425
rect 4295 1325 4300 1425
rect 4200 1310 4300 1325
rect 4450 1425 4550 1440
rect 4450 1325 4455 1425
rect 4490 1325 4510 1425
rect 4545 1325 4550 1425
rect 4450 1310 4550 1325
rect 4700 1425 4800 1440
rect 4700 1325 4705 1425
rect 4740 1325 4760 1425
rect 4795 1325 4800 1425
rect 4700 1310 4800 1325
rect 4950 1425 5050 1440
rect 4950 1325 4955 1425
rect 4990 1325 5010 1425
rect 5045 1325 5050 1425
rect 4950 1310 5050 1325
rect 5200 1425 5300 1440
rect 5200 1325 5205 1425
rect 5240 1325 5260 1425
rect 5295 1325 5300 1425
rect 5200 1310 5300 1325
rect 5450 1425 5550 1440
rect 5450 1325 5455 1425
rect 5490 1325 5510 1425
rect 5545 1325 5550 1425
rect 5450 1310 5550 1325
rect 5700 1425 5800 1440
rect 5700 1325 5705 1425
rect 5740 1325 5760 1425
rect 5795 1325 5800 1425
rect 5700 1310 5800 1325
rect 5950 1425 6050 1440
rect 5950 1325 5955 1425
rect 5990 1325 6010 1425
rect 6045 1325 6050 1425
rect 5950 1310 6050 1325
rect 6200 1425 6300 1440
rect 6200 1325 6205 1425
rect 6240 1325 6260 1425
rect 6295 1325 6300 1425
rect 6200 1310 6300 1325
rect 6450 1425 6550 1440
rect 6450 1325 6455 1425
rect 6490 1325 6510 1425
rect 6545 1325 6550 1425
rect 6450 1310 6550 1325
rect 6700 1425 6800 1440
rect 6700 1325 6705 1425
rect 6740 1325 6760 1425
rect 6795 1325 6800 1425
rect 6700 1310 6800 1325
rect 6950 1425 7050 1440
rect 6950 1325 6955 1425
rect 6990 1325 7010 1425
rect 7045 1325 7050 1425
rect 6950 1310 7050 1325
rect 7200 1425 7300 1440
rect 7200 1325 7205 1425
rect 7240 1325 7260 1425
rect 7295 1325 7300 1425
rect 7200 1310 7300 1325
rect 7450 1425 7550 1440
rect 7450 1325 7455 1425
rect 7490 1325 7510 1425
rect 7545 1325 7550 1425
rect 7450 1310 7550 1325
rect 7700 1425 7800 1440
rect 7700 1325 7705 1425
rect 7740 1325 7760 1425
rect 7795 1325 7800 1425
rect 7700 1310 7800 1325
rect 7950 1425 8000 1440
rect 7950 1325 7955 1425
rect 7990 1325 8000 1425
rect 7950 1310 8000 1325
rect 0 1300 60 1310
rect 190 1300 310 1310
rect 440 1300 560 1310
rect 690 1300 810 1310
rect 940 1300 1060 1310
rect 1190 1300 1310 1310
rect 1440 1300 1560 1310
rect 1690 1300 1810 1310
rect 1940 1300 2060 1310
rect 2190 1300 2310 1310
rect 2440 1300 2560 1310
rect 2690 1300 2810 1310
rect 2940 1300 3060 1310
rect 3190 1300 3310 1310
rect 3440 1300 3560 1310
rect 3690 1300 3810 1310
rect 3940 1300 4060 1310
rect 4190 1300 4310 1310
rect 4440 1300 4560 1310
rect 4690 1300 4810 1310
rect 4940 1300 5060 1310
rect 5190 1300 5310 1310
rect 5440 1300 5560 1310
rect 5690 1300 5810 1310
rect 5940 1300 6060 1310
rect 6190 1300 6310 1310
rect 6440 1300 6560 1310
rect 6690 1300 6810 1310
rect 6940 1300 7060 1310
rect 7190 1300 7310 1310
rect 7440 1300 7560 1310
rect 7690 1300 7810 1310
rect 7940 1300 8000 1310
rect 0 1295 200 1300
rect 0 1260 75 1295
rect 175 1260 200 1295
rect 0 1240 200 1260
rect 0 1205 75 1240
rect 175 1205 200 1240
rect 0 1200 200 1205
rect 300 1295 450 1300
rect 300 1260 325 1295
rect 425 1260 450 1295
rect 300 1240 450 1260
rect 300 1205 325 1240
rect 425 1205 450 1240
rect 300 1200 450 1205
rect 550 1295 700 1300
rect 550 1260 575 1295
rect 675 1260 700 1295
rect 550 1240 700 1260
rect 550 1205 575 1240
rect 675 1205 700 1240
rect 550 1200 700 1205
rect 800 1295 1200 1300
rect 800 1260 825 1295
rect 925 1260 1075 1295
rect 1175 1260 1200 1295
rect 800 1240 1200 1260
rect 800 1205 825 1240
rect 925 1205 1075 1240
rect 1175 1205 1200 1240
rect 800 1200 1200 1205
rect 1300 1295 1450 1300
rect 1300 1260 1325 1295
rect 1425 1260 1450 1295
rect 1300 1240 1450 1260
rect 1300 1205 1325 1240
rect 1425 1205 1450 1240
rect 1300 1200 1450 1205
rect 1550 1295 1700 1300
rect 1550 1260 1575 1295
rect 1675 1260 1700 1295
rect 1550 1240 1700 1260
rect 1550 1205 1575 1240
rect 1675 1205 1700 1240
rect 1550 1200 1700 1205
rect 1800 1295 2200 1300
rect 1800 1260 1825 1295
rect 1925 1260 2075 1295
rect 2175 1260 2200 1295
rect 1800 1240 2200 1260
rect 1800 1205 1825 1240
rect 1925 1205 2075 1240
rect 2175 1205 2200 1240
rect 1800 1200 2200 1205
rect 2300 1295 2450 1300
rect 2300 1260 2325 1295
rect 2425 1260 2450 1295
rect 2300 1240 2450 1260
rect 2300 1205 2325 1240
rect 2425 1205 2450 1240
rect 2300 1200 2450 1205
rect 2550 1295 2700 1300
rect 2550 1260 2575 1295
rect 2675 1260 2700 1295
rect 2550 1240 2700 1260
rect 2550 1205 2575 1240
rect 2675 1205 2700 1240
rect 2550 1200 2700 1205
rect 2800 1295 3200 1300
rect 2800 1260 2825 1295
rect 2925 1260 3075 1295
rect 3175 1260 3200 1295
rect 2800 1240 3200 1260
rect 2800 1205 2825 1240
rect 2925 1205 3075 1240
rect 3175 1205 3200 1240
rect 2800 1200 3200 1205
rect 3300 1295 3450 1300
rect 3300 1260 3325 1295
rect 3425 1260 3450 1295
rect 3300 1240 3450 1260
rect 3300 1205 3325 1240
rect 3425 1205 3450 1240
rect 3300 1200 3450 1205
rect 3550 1295 3700 1300
rect 3550 1260 3575 1295
rect 3675 1260 3700 1295
rect 3550 1240 3700 1260
rect 3550 1205 3575 1240
rect 3675 1205 3700 1240
rect 3550 1200 3700 1205
rect 3800 1295 4200 1300
rect 3800 1260 3825 1295
rect 3925 1260 4075 1295
rect 4175 1260 4200 1295
rect 3800 1240 4200 1260
rect 3800 1205 3825 1240
rect 3925 1205 4075 1240
rect 4175 1205 4200 1240
rect 3800 1200 4200 1205
rect 4300 1295 4450 1300
rect 4300 1260 4325 1295
rect 4425 1260 4450 1295
rect 4300 1240 4450 1260
rect 4300 1205 4325 1240
rect 4425 1205 4450 1240
rect 4300 1200 4450 1205
rect 4550 1295 4700 1300
rect 4550 1260 4575 1295
rect 4675 1260 4700 1295
rect 4550 1240 4700 1260
rect 4550 1205 4575 1240
rect 4675 1205 4700 1240
rect 4550 1200 4700 1205
rect 4800 1295 5200 1300
rect 4800 1260 4825 1295
rect 4925 1260 5075 1295
rect 5175 1260 5200 1295
rect 4800 1240 5200 1260
rect 4800 1205 4825 1240
rect 4925 1205 5075 1240
rect 5175 1205 5200 1240
rect 4800 1200 5200 1205
rect 5300 1295 5450 1300
rect 5300 1260 5325 1295
rect 5425 1260 5450 1295
rect 5300 1240 5450 1260
rect 5300 1205 5325 1240
rect 5425 1205 5450 1240
rect 5300 1200 5450 1205
rect 5550 1295 5700 1300
rect 5550 1260 5575 1295
rect 5675 1260 5700 1295
rect 5550 1240 5700 1260
rect 5550 1205 5575 1240
rect 5675 1205 5700 1240
rect 5550 1200 5700 1205
rect 5800 1295 6200 1300
rect 5800 1260 5825 1295
rect 5925 1260 6075 1295
rect 6175 1260 6200 1295
rect 5800 1240 6200 1260
rect 5800 1205 5825 1240
rect 5925 1205 6075 1240
rect 6175 1205 6200 1240
rect 5800 1200 6200 1205
rect 6300 1295 6450 1300
rect 6300 1260 6325 1295
rect 6425 1260 6450 1295
rect 6300 1240 6450 1260
rect 6300 1205 6325 1240
rect 6425 1205 6450 1240
rect 6300 1200 6450 1205
rect 6550 1295 6700 1300
rect 6550 1260 6575 1295
rect 6675 1260 6700 1295
rect 6550 1240 6700 1260
rect 6550 1205 6575 1240
rect 6675 1205 6700 1240
rect 6550 1200 6700 1205
rect 6800 1295 7200 1300
rect 6800 1260 6825 1295
rect 6925 1260 7075 1295
rect 7175 1260 7200 1295
rect 6800 1240 7200 1260
rect 6800 1205 6825 1240
rect 6925 1205 7075 1240
rect 7175 1205 7200 1240
rect 6800 1200 7200 1205
rect 7300 1295 7450 1300
rect 7300 1260 7325 1295
rect 7425 1260 7450 1295
rect 7300 1240 7450 1260
rect 7300 1205 7325 1240
rect 7425 1205 7450 1240
rect 7300 1200 7450 1205
rect 7550 1295 7700 1300
rect 7550 1260 7575 1295
rect 7675 1260 7700 1295
rect 7550 1240 7700 1260
rect 7550 1205 7575 1240
rect 7675 1205 7700 1240
rect 7550 1200 7700 1205
rect 7800 1295 8000 1300
rect 7800 1260 7825 1295
rect 7925 1260 8000 1295
rect 7800 1240 8000 1260
rect 7800 1205 7825 1240
rect 7925 1205 8000 1240
rect 7800 1200 8000 1205
rect 0 1190 60 1200
rect 190 1190 310 1200
rect 440 1190 560 1200
rect 690 1190 810 1200
rect 940 1190 1060 1200
rect 1190 1190 1310 1200
rect 1440 1190 1560 1200
rect 1690 1190 1810 1200
rect 1940 1190 2060 1200
rect 2190 1190 2310 1200
rect 2440 1190 2560 1200
rect 2690 1190 2810 1200
rect 2940 1190 3060 1200
rect 3190 1190 3310 1200
rect 3440 1190 3560 1200
rect 3690 1190 3810 1200
rect 3940 1190 4060 1200
rect 4190 1190 4310 1200
rect 4440 1190 4560 1200
rect 4690 1190 4810 1200
rect 4940 1190 5060 1200
rect 5190 1190 5310 1200
rect 5440 1190 5560 1200
rect 5690 1190 5810 1200
rect 5940 1190 6060 1200
rect 6190 1190 6310 1200
rect 6440 1190 6560 1200
rect 6690 1190 6810 1200
rect 6940 1190 7060 1200
rect 7190 1190 7310 1200
rect 7440 1190 7560 1200
rect 7690 1190 7810 1200
rect 7940 1190 8000 1200
rect 0 1175 50 1190
rect 0 1075 10 1175
rect 45 1075 50 1175
rect 0 1060 50 1075
rect 200 1175 300 1190
rect 200 1075 205 1175
rect 240 1075 260 1175
rect 295 1075 300 1175
rect 200 1060 300 1075
rect 450 1175 550 1190
rect 450 1075 455 1175
rect 490 1075 510 1175
rect 545 1075 550 1175
rect 450 1060 550 1075
rect 700 1175 800 1190
rect 700 1075 705 1175
rect 740 1075 760 1175
rect 795 1075 800 1175
rect 700 1060 800 1075
rect 950 1175 1050 1190
rect 950 1075 955 1175
rect 990 1075 1010 1175
rect 1045 1075 1050 1175
rect 950 1060 1050 1075
rect 1200 1175 1300 1190
rect 1200 1075 1205 1175
rect 1240 1075 1260 1175
rect 1295 1075 1300 1175
rect 1200 1060 1300 1075
rect 1450 1175 1550 1190
rect 1450 1075 1455 1175
rect 1490 1075 1510 1175
rect 1545 1075 1550 1175
rect 1450 1060 1550 1075
rect 1700 1175 1800 1190
rect 1700 1075 1705 1175
rect 1740 1075 1760 1175
rect 1795 1075 1800 1175
rect 1700 1060 1800 1075
rect 1950 1175 2050 1190
rect 1950 1075 1955 1175
rect 1990 1075 2010 1175
rect 2045 1075 2050 1175
rect 1950 1060 2050 1075
rect 2200 1175 2300 1190
rect 2200 1075 2205 1175
rect 2240 1075 2260 1175
rect 2295 1075 2300 1175
rect 2200 1060 2300 1075
rect 2450 1175 2550 1190
rect 2450 1075 2455 1175
rect 2490 1075 2510 1175
rect 2545 1075 2550 1175
rect 2450 1060 2550 1075
rect 2700 1175 2800 1190
rect 2700 1075 2705 1175
rect 2740 1075 2760 1175
rect 2795 1075 2800 1175
rect 2700 1060 2800 1075
rect 2950 1175 3050 1190
rect 2950 1075 2955 1175
rect 2990 1075 3010 1175
rect 3045 1075 3050 1175
rect 2950 1060 3050 1075
rect 3200 1175 3300 1190
rect 3200 1075 3205 1175
rect 3240 1075 3260 1175
rect 3295 1075 3300 1175
rect 3200 1060 3300 1075
rect 3450 1175 3550 1190
rect 3450 1075 3455 1175
rect 3490 1075 3510 1175
rect 3545 1075 3550 1175
rect 3450 1060 3550 1075
rect 3700 1175 3800 1190
rect 3700 1075 3705 1175
rect 3740 1075 3760 1175
rect 3795 1075 3800 1175
rect 3700 1060 3800 1075
rect 3950 1175 4050 1190
rect 3950 1075 3955 1175
rect 3990 1075 4010 1175
rect 4045 1075 4050 1175
rect 3950 1060 4050 1075
rect 4200 1175 4300 1190
rect 4200 1075 4205 1175
rect 4240 1075 4260 1175
rect 4295 1075 4300 1175
rect 4200 1060 4300 1075
rect 4450 1175 4550 1190
rect 4450 1075 4455 1175
rect 4490 1075 4510 1175
rect 4545 1075 4550 1175
rect 4450 1060 4550 1075
rect 4700 1175 4800 1190
rect 4700 1075 4705 1175
rect 4740 1075 4760 1175
rect 4795 1075 4800 1175
rect 4700 1060 4800 1075
rect 4950 1175 5050 1190
rect 4950 1075 4955 1175
rect 4990 1075 5010 1175
rect 5045 1075 5050 1175
rect 4950 1060 5050 1075
rect 5200 1175 5300 1190
rect 5200 1075 5205 1175
rect 5240 1075 5260 1175
rect 5295 1075 5300 1175
rect 5200 1060 5300 1075
rect 5450 1175 5550 1190
rect 5450 1075 5455 1175
rect 5490 1075 5510 1175
rect 5545 1075 5550 1175
rect 5450 1060 5550 1075
rect 5700 1175 5800 1190
rect 5700 1075 5705 1175
rect 5740 1075 5760 1175
rect 5795 1075 5800 1175
rect 5700 1060 5800 1075
rect 5950 1175 6050 1190
rect 5950 1075 5955 1175
rect 5990 1075 6010 1175
rect 6045 1075 6050 1175
rect 5950 1060 6050 1075
rect 6200 1175 6300 1190
rect 6200 1075 6205 1175
rect 6240 1075 6260 1175
rect 6295 1075 6300 1175
rect 6200 1060 6300 1075
rect 6450 1175 6550 1190
rect 6450 1075 6455 1175
rect 6490 1075 6510 1175
rect 6545 1075 6550 1175
rect 6450 1060 6550 1075
rect 6700 1175 6800 1190
rect 6700 1075 6705 1175
rect 6740 1075 6760 1175
rect 6795 1075 6800 1175
rect 6700 1060 6800 1075
rect 6950 1175 7050 1190
rect 6950 1075 6955 1175
rect 6990 1075 7010 1175
rect 7045 1075 7050 1175
rect 6950 1060 7050 1075
rect 7200 1175 7300 1190
rect 7200 1075 7205 1175
rect 7240 1075 7260 1175
rect 7295 1075 7300 1175
rect 7200 1060 7300 1075
rect 7450 1175 7550 1190
rect 7450 1075 7455 1175
rect 7490 1075 7510 1175
rect 7545 1075 7550 1175
rect 7450 1060 7550 1075
rect 7700 1175 7800 1190
rect 7700 1075 7705 1175
rect 7740 1075 7760 1175
rect 7795 1075 7800 1175
rect 7700 1060 7800 1075
rect 7950 1175 8000 1190
rect 7950 1075 7955 1175
rect 7990 1075 8000 1175
rect 7950 1060 8000 1075
rect 0 1050 60 1060
rect 190 1050 310 1060
rect 440 1050 560 1060
rect 690 1050 810 1060
rect 940 1050 1060 1060
rect 1190 1050 1310 1060
rect 1440 1050 1560 1060
rect 1690 1050 1810 1060
rect 1940 1050 2060 1060
rect 2190 1050 2310 1060
rect 2440 1050 2560 1060
rect 2690 1050 2810 1060
rect 2940 1050 3060 1060
rect 3190 1050 3310 1060
rect 3440 1050 3560 1060
rect 3690 1050 3810 1060
rect 3940 1050 4060 1060
rect 4190 1050 4310 1060
rect 4440 1050 4560 1060
rect 4690 1050 4810 1060
rect 4940 1050 5060 1060
rect 5190 1050 5310 1060
rect 5440 1050 5560 1060
rect 5690 1050 5810 1060
rect 5940 1050 6060 1060
rect 6190 1050 6310 1060
rect 6440 1050 6560 1060
rect 6690 1050 6810 1060
rect 6940 1050 7060 1060
rect 7190 1050 7310 1060
rect 7440 1050 7560 1060
rect 7690 1050 7810 1060
rect 7940 1050 8000 1060
rect 0 1045 450 1050
rect 0 1010 75 1045
rect 175 1010 325 1045
rect 425 1010 450 1045
rect 0 990 450 1010
rect 0 955 75 990
rect 175 955 325 990
rect 425 955 450 990
rect 0 950 450 955
rect 550 1045 1450 1050
rect 550 1010 575 1045
rect 675 1010 825 1045
rect 925 1010 1075 1045
rect 1175 1010 1325 1045
rect 1425 1010 1450 1045
rect 550 990 1450 1010
rect 550 955 575 990
rect 675 955 825 990
rect 925 955 1075 990
rect 1175 955 1325 990
rect 1425 955 1450 990
rect 550 950 1450 955
rect 1550 1045 2450 1050
rect 1550 1010 1575 1045
rect 1675 1010 1825 1045
rect 1925 1010 2075 1045
rect 2175 1010 2325 1045
rect 2425 1010 2450 1045
rect 1550 990 2450 1010
rect 1550 955 1575 990
rect 1675 955 1825 990
rect 1925 955 2075 990
rect 2175 955 2325 990
rect 2425 955 2450 990
rect 1550 950 2450 955
rect 2550 1045 3450 1050
rect 2550 1010 2575 1045
rect 2675 1010 2825 1045
rect 2925 1010 3075 1045
rect 3175 1010 3325 1045
rect 3425 1010 3450 1045
rect 2550 990 3450 1010
rect 2550 955 2575 990
rect 2675 955 2825 990
rect 2925 955 3075 990
rect 3175 955 3325 990
rect 3425 955 3450 990
rect 2550 950 3450 955
rect 3550 1045 4450 1050
rect 3550 1010 3575 1045
rect 3675 1010 3825 1045
rect 3925 1010 4075 1045
rect 4175 1010 4325 1045
rect 4425 1010 4450 1045
rect 3550 990 4450 1010
rect 3550 955 3575 990
rect 3675 955 3825 990
rect 3925 955 4075 990
rect 4175 955 4325 990
rect 4425 955 4450 990
rect 3550 950 4450 955
rect 4550 1045 5450 1050
rect 4550 1010 4575 1045
rect 4675 1010 4825 1045
rect 4925 1010 5075 1045
rect 5175 1010 5325 1045
rect 5425 1010 5450 1045
rect 4550 990 5450 1010
rect 4550 955 4575 990
rect 4675 955 4825 990
rect 4925 955 5075 990
rect 5175 955 5325 990
rect 5425 955 5450 990
rect 4550 950 5450 955
rect 5550 1045 6450 1050
rect 5550 1010 5575 1045
rect 5675 1010 5825 1045
rect 5925 1010 6075 1045
rect 6175 1010 6325 1045
rect 6425 1010 6450 1045
rect 5550 990 6450 1010
rect 5550 955 5575 990
rect 5675 955 5825 990
rect 5925 955 6075 990
rect 6175 955 6325 990
rect 6425 955 6450 990
rect 5550 950 6450 955
rect 6550 1045 7450 1050
rect 6550 1010 6575 1045
rect 6675 1010 6825 1045
rect 6925 1010 7075 1045
rect 7175 1010 7325 1045
rect 7425 1010 7450 1045
rect 6550 990 7450 1010
rect 6550 955 6575 990
rect 6675 955 6825 990
rect 6925 955 7075 990
rect 7175 955 7325 990
rect 7425 955 7450 990
rect 6550 950 7450 955
rect 7550 1045 8000 1050
rect 7550 1010 7575 1045
rect 7675 1010 7825 1045
rect 7925 1010 8000 1045
rect 7550 990 8000 1010
rect 7550 955 7575 990
rect 7675 955 7825 990
rect 7925 955 8000 990
rect 7550 950 8000 955
rect 0 940 60 950
rect 190 940 310 950
rect 440 940 560 950
rect 690 940 810 950
rect 940 940 1060 950
rect 1190 940 1310 950
rect 1440 940 1560 950
rect 1690 940 1810 950
rect 1940 940 2060 950
rect 2190 940 2310 950
rect 2440 940 2560 950
rect 2690 940 2810 950
rect 2940 940 3060 950
rect 3190 940 3310 950
rect 3440 940 3560 950
rect 3690 940 3810 950
rect 3940 940 4060 950
rect 4190 940 4310 950
rect 4440 940 4560 950
rect 4690 940 4810 950
rect 4940 940 5060 950
rect 5190 940 5310 950
rect 5440 940 5560 950
rect 5690 940 5810 950
rect 5940 940 6060 950
rect 6190 940 6310 950
rect 6440 940 6560 950
rect 6690 940 6810 950
rect 6940 940 7060 950
rect 7190 940 7310 950
rect 7440 940 7560 950
rect 7690 940 7810 950
rect 7940 940 8000 950
rect 0 925 50 940
rect 0 825 10 925
rect 45 825 50 925
rect 0 810 50 825
rect 200 925 300 940
rect 200 825 205 925
rect 240 825 260 925
rect 295 825 300 925
rect 200 810 300 825
rect 450 925 550 940
rect 450 825 455 925
rect 490 825 510 925
rect 545 825 550 925
rect 450 810 550 825
rect 700 925 800 940
rect 700 825 705 925
rect 740 825 760 925
rect 795 825 800 925
rect 700 810 800 825
rect 950 925 1050 940
rect 950 825 955 925
rect 990 825 1010 925
rect 1045 825 1050 925
rect 950 810 1050 825
rect 1200 925 1300 940
rect 1200 825 1205 925
rect 1240 825 1260 925
rect 1295 825 1300 925
rect 1200 810 1300 825
rect 1450 925 1550 940
rect 1450 825 1455 925
rect 1490 825 1510 925
rect 1545 825 1550 925
rect 1450 810 1550 825
rect 1700 925 1800 940
rect 1700 825 1705 925
rect 1740 825 1760 925
rect 1795 825 1800 925
rect 1700 810 1800 825
rect 1950 925 2050 940
rect 1950 825 1955 925
rect 1990 825 2010 925
rect 2045 825 2050 925
rect 1950 810 2050 825
rect 2200 925 2300 940
rect 2200 825 2205 925
rect 2240 825 2260 925
rect 2295 825 2300 925
rect 2200 810 2300 825
rect 2450 925 2550 940
rect 2450 825 2455 925
rect 2490 825 2510 925
rect 2545 825 2550 925
rect 2450 810 2550 825
rect 2700 925 2800 940
rect 2700 825 2705 925
rect 2740 825 2760 925
rect 2795 825 2800 925
rect 2700 810 2800 825
rect 2950 925 3050 940
rect 2950 825 2955 925
rect 2990 825 3010 925
rect 3045 825 3050 925
rect 2950 810 3050 825
rect 3200 925 3300 940
rect 3200 825 3205 925
rect 3240 825 3260 925
rect 3295 825 3300 925
rect 3200 810 3300 825
rect 3450 925 3550 940
rect 3450 825 3455 925
rect 3490 825 3510 925
rect 3545 825 3550 925
rect 3450 810 3550 825
rect 3700 925 3800 940
rect 3700 825 3705 925
rect 3740 825 3760 925
rect 3795 825 3800 925
rect 3700 810 3800 825
rect 3950 925 4050 940
rect 3950 825 3955 925
rect 3990 825 4010 925
rect 4045 825 4050 925
rect 3950 810 4050 825
rect 4200 925 4300 940
rect 4200 825 4205 925
rect 4240 825 4260 925
rect 4295 825 4300 925
rect 4200 810 4300 825
rect 4450 925 4550 940
rect 4450 825 4455 925
rect 4490 825 4510 925
rect 4545 825 4550 925
rect 4450 810 4550 825
rect 4700 925 4800 940
rect 4700 825 4705 925
rect 4740 825 4760 925
rect 4795 825 4800 925
rect 4700 810 4800 825
rect 4950 925 5050 940
rect 4950 825 4955 925
rect 4990 825 5010 925
rect 5045 825 5050 925
rect 4950 810 5050 825
rect 5200 925 5300 940
rect 5200 825 5205 925
rect 5240 825 5260 925
rect 5295 825 5300 925
rect 5200 810 5300 825
rect 5450 925 5550 940
rect 5450 825 5455 925
rect 5490 825 5510 925
rect 5545 825 5550 925
rect 5450 810 5550 825
rect 5700 925 5800 940
rect 5700 825 5705 925
rect 5740 825 5760 925
rect 5795 825 5800 925
rect 5700 810 5800 825
rect 5950 925 6050 940
rect 5950 825 5955 925
rect 5990 825 6010 925
rect 6045 825 6050 925
rect 5950 810 6050 825
rect 6200 925 6300 940
rect 6200 825 6205 925
rect 6240 825 6260 925
rect 6295 825 6300 925
rect 6200 810 6300 825
rect 6450 925 6550 940
rect 6450 825 6455 925
rect 6490 825 6510 925
rect 6545 825 6550 925
rect 6450 810 6550 825
rect 6700 925 6800 940
rect 6700 825 6705 925
rect 6740 825 6760 925
rect 6795 825 6800 925
rect 6700 810 6800 825
rect 6950 925 7050 940
rect 6950 825 6955 925
rect 6990 825 7010 925
rect 7045 825 7050 925
rect 6950 810 7050 825
rect 7200 925 7300 940
rect 7200 825 7205 925
rect 7240 825 7260 925
rect 7295 825 7300 925
rect 7200 810 7300 825
rect 7450 925 7550 940
rect 7450 825 7455 925
rect 7490 825 7510 925
rect 7545 825 7550 925
rect 7450 810 7550 825
rect 7700 925 7800 940
rect 7700 825 7705 925
rect 7740 825 7760 925
rect 7795 825 7800 925
rect 7700 810 7800 825
rect 7950 925 8000 940
rect 7950 825 7955 925
rect 7990 825 8000 925
rect 7950 810 8000 825
rect 0 800 60 810
rect 190 800 310 810
rect 440 800 560 810
rect 690 800 810 810
rect 940 800 1060 810
rect 1190 800 1310 810
rect 1440 800 1560 810
rect 1690 800 1810 810
rect 1940 800 2060 810
rect 2190 800 2310 810
rect 2440 800 2560 810
rect 2690 800 2810 810
rect 2940 800 3060 810
rect 3190 800 3310 810
rect 3440 800 3560 810
rect 3690 800 3810 810
rect 3940 800 4060 810
rect 4190 800 4310 810
rect 4440 800 4560 810
rect 4690 800 4810 810
rect 4940 800 5060 810
rect 5190 800 5310 810
rect 5440 800 5560 810
rect 5690 800 5810 810
rect 5940 800 6060 810
rect 6190 800 6310 810
rect 6440 800 6560 810
rect 6690 800 6810 810
rect 6940 800 7060 810
rect 7190 800 7310 810
rect 7440 800 7560 810
rect 7690 800 7810 810
rect 7940 800 8000 810
rect 0 795 200 800
rect 0 760 75 795
rect 175 760 200 795
rect 0 740 200 760
rect 0 705 75 740
rect 175 705 200 740
rect 0 700 200 705
rect 300 795 450 800
rect 300 760 325 795
rect 425 760 450 795
rect 300 740 450 760
rect 300 705 325 740
rect 425 705 450 740
rect 300 700 450 705
rect 550 795 700 800
rect 550 760 575 795
rect 675 760 700 795
rect 550 740 700 760
rect 550 705 575 740
rect 675 705 700 740
rect 550 700 700 705
rect 800 795 1200 800
rect 800 760 825 795
rect 925 760 1075 795
rect 1175 760 1200 795
rect 800 740 1200 760
rect 800 705 825 740
rect 925 705 1075 740
rect 1175 705 1200 740
rect 800 700 1200 705
rect 1300 795 1450 800
rect 1300 760 1325 795
rect 1425 760 1450 795
rect 1300 740 1450 760
rect 1300 705 1325 740
rect 1425 705 1450 740
rect 1300 700 1450 705
rect 1550 795 1700 800
rect 1550 760 1575 795
rect 1675 760 1700 795
rect 1550 740 1700 760
rect 1550 705 1575 740
rect 1675 705 1700 740
rect 1550 700 1700 705
rect 1800 795 2200 800
rect 1800 760 1825 795
rect 1925 760 2075 795
rect 2175 760 2200 795
rect 1800 740 2200 760
rect 1800 705 1825 740
rect 1925 705 2075 740
rect 2175 705 2200 740
rect 1800 700 2200 705
rect 2300 795 2450 800
rect 2300 760 2325 795
rect 2425 760 2450 795
rect 2300 740 2450 760
rect 2300 705 2325 740
rect 2425 705 2450 740
rect 2300 700 2450 705
rect 2550 795 2700 800
rect 2550 760 2575 795
rect 2675 760 2700 795
rect 2550 740 2700 760
rect 2550 705 2575 740
rect 2675 705 2700 740
rect 2550 700 2700 705
rect 2800 795 3200 800
rect 2800 760 2825 795
rect 2925 760 3075 795
rect 3175 760 3200 795
rect 2800 740 3200 760
rect 2800 705 2825 740
rect 2925 705 3075 740
rect 3175 705 3200 740
rect 2800 700 3200 705
rect 3300 795 3450 800
rect 3300 760 3325 795
rect 3425 760 3450 795
rect 3300 740 3450 760
rect 3300 705 3325 740
rect 3425 705 3450 740
rect 3300 700 3450 705
rect 3550 795 3700 800
rect 3550 760 3575 795
rect 3675 760 3700 795
rect 3550 740 3700 760
rect 3550 705 3575 740
rect 3675 705 3700 740
rect 3550 700 3700 705
rect 3800 795 4200 800
rect 3800 760 3825 795
rect 3925 760 4075 795
rect 4175 760 4200 795
rect 3800 740 4200 760
rect 3800 705 3825 740
rect 3925 705 4075 740
rect 4175 705 4200 740
rect 3800 700 4200 705
rect 4300 795 4450 800
rect 4300 760 4325 795
rect 4425 760 4450 795
rect 4300 740 4450 760
rect 4300 705 4325 740
rect 4425 705 4450 740
rect 4300 700 4450 705
rect 4550 795 4700 800
rect 4550 760 4575 795
rect 4675 760 4700 795
rect 4550 740 4700 760
rect 4550 705 4575 740
rect 4675 705 4700 740
rect 4550 700 4700 705
rect 4800 795 5200 800
rect 4800 760 4825 795
rect 4925 760 5075 795
rect 5175 760 5200 795
rect 4800 740 5200 760
rect 4800 705 4825 740
rect 4925 705 5075 740
rect 5175 705 5200 740
rect 4800 700 5200 705
rect 5300 795 5450 800
rect 5300 760 5325 795
rect 5425 760 5450 795
rect 5300 740 5450 760
rect 5300 705 5325 740
rect 5425 705 5450 740
rect 5300 700 5450 705
rect 5550 795 5700 800
rect 5550 760 5575 795
rect 5675 760 5700 795
rect 5550 740 5700 760
rect 5550 705 5575 740
rect 5675 705 5700 740
rect 5550 700 5700 705
rect 5800 795 6200 800
rect 5800 760 5825 795
rect 5925 760 6075 795
rect 6175 760 6200 795
rect 5800 740 6200 760
rect 5800 705 5825 740
rect 5925 705 6075 740
rect 6175 705 6200 740
rect 5800 700 6200 705
rect 6300 795 6450 800
rect 6300 760 6325 795
rect 6425 760 6450 795
rect 6300 740 6450 760
rect 6300 705 6325 740
rect 6425 705 6450 740
rect 6300 700 6450 705
rect 6550 795 6700 800
rect 6550 760 6575 795
rect 6675 760 6700 795
rect 6550 740 6700 760
rect 6550 705 6575 740
rect 6675 705 6700 740
rect 6550 700 6700 705
rect 6800 795 7200 800
rect 6800 760 6825 795
rect 6925 760 7075 795
rect 7175 760 7200 795
rect 6800 740 7200 760
rect 6800 705 6825 740
rect 6925 705 7075 740
rect 7175 705 7200 740
rect 6800 700 7200 705
rect 7300 795 7450 800
rect 7300 760 7325 795
rect 7425 760 7450 795
rect 7300 740 7450 760
rect 7300 705 7325 740
rect 7425 705 7450 740
rect 7300 700 7450 705
rect 7550 795 7700 800
rect 7550 760 7575 795
rect 7675 760 7700 795
rect 7550 740 7700 760
rect 7550 705 7575 740
rect 7675 705 7700 740
rect 7550 700 7700 705
rect 7800 795 8000 800
rect 7800 760 7825 795
rect 7925 760 8000 795
rect 7800 740 8000 760
rect 7800 705 7825 740
rect 7925 705 8000 740
rect 7800 700 8000 705
rect 0 690 60 700
rect 190 690 310 700
rect 440 690 560 700
rect 690 690 810 700
rect 940 690 1060 700
rect 1190 690 1310 700
rect 1440 690 1560 700
rect 1690 690 1810 700
rect 1940 690 2060 700
rect 2190 690 2310 700
rect 2440 690 2560 700
rect 2690 690 2810 700
rect 2940 690 3060 700
rect 3190 690 3310 700
rect 3440 690 3560 700
rect 3690 690 3810 700
rect 3940 690 4060 700
rect 4190 690 4310 700
rect 4440 690 4560 700
rect 4690 690 4810 700
rect 4940 690 5060 700
rect 5190 690 5310 700
rect 5440 690 5560 700
rect 5690 690 5810 700
rect 5940 690 6060 700
rect 6190 690 6310 700
rect 6440 690 6560 700
rect 6690 690 6810 700
rect 6940 690 7060 700
rect 7190 690 7310 700
rect 7440 690 7560 700
rect 7690 690 7810 700
rect 7940 690 8000 700
rect 0 675 50 690
rect 0 575 10 675
rect 45 575 50 675
rect 0 560 50 575
rect 200 675 300 690
rect 200 575 205 675
rect 240 575 260 675
rect 295 575 300 675
rect 200 560 300 575
rect 450 675 550 690
rect 450 575 455 675
rect 490 575 510 675
rect 545 575 550 675
rect 450 560 550 575
rect 700 675 800 690
rect 700 575 705 675
rect 740 575 760 675
rect 795 575 800 675
rect 700 560 800 575
rect 950 675 1050 690
rect 950 575 955 675
rect 990 575 1010 675
rect 1045 575 1050 675
rect 950 560 1050 575
rect 1200 675 1300 690
rect 1200 575 1205 675
rect 1240 575 1260 675
rect 1295 575 1300 675
rect 1200 560 1300 575
rect 1450 675 1550 690
rect 1450 575 1455 675
rect 1490 575 1510 675
rect 1545 575 1550 675
rect 1450 560 1550 575
rect 1700 675 1800 690
rect 1700 575 1705 675
rect 1740 575 1760 675
rect 1795 575 1800 675
rect 1700 560 1800 575
rect 1950 675 2050 690
rect 1950 575 1955 675
rect 1990 575 2010 675
rect 2045 575 2050 675
rect 1950 560 2050 575
rect 2200 675 2300 690
rect 2200 575 2205 675
rect 2240 575 2260 675
rect 2295 575 2300 675
rect 2200 560 2300 575
rect 2450 675 2550 690
rect 2450 575 2455 675
rect 2490 575 2510 675
rect 2545 575 2550 675
rect 2450 560 2550 575
rect 2700 675 2800 690
rect 2700 575 2705 675
rect 2740 575 2760 675
rect 2795 575 2800 675
rect 2700 560 2800 575
rect 2950 675 3050 690
rect 2950 575 2955 675
rect 2990 575 3010 675
rect 3045 575 3050 675
rect 2950 560 3050 575
rect 3200 675 3300 690
rect 3200 575 3205 675
rect 3240 575 3260 675
rect 3295 575 3300 675
rect 3200 560 3300 575
rect 3450 675 3550 690
rect 3450 575 3455 675
rect 3490 575 3510 675
rect 3545 575 3550 675
rect 3450 560 3550 575
rect 3700 675 3800 690
rect 3700 575 3705 675
rect 3740 575 3760 675
rect 3795 575 3800 675
rect 3700 560 3800 575
rect 3950 675 4050 690
rect 3950 575 3955 675
rect 3990 575 4010 675
rect 4045 575 4050 675
rect 3950 560 4050 575
rect 4200 675 4300 690
rect 4200 575 4205 675
rect 4240 575 4260 675
rect 4295 575 4300 675
rect 4200 560 4300 575
rect 4450 675 4550 690
rect 4450 575 4455 675
rect 4490 575 4510 675
rect 4545 575 4550 675
rect 4450 560 4550 575
rect 4700 675 4800 690
rect 4700 575 4705 675
rect 4740 575 4760 675
rect 4795 575 4800 675
rect 4700 560 4800 575
rect 4950 675 5050 690
rect 4950 575 4955 675
rect 4990 575 5010 675
rect 5045 575 5050 675
rect 4950 560 5050 575
rect 5200 675 5300 690
rect 5200 575 5205 675
rect 5240 575 5260 675
rect 5295 575 5300 675
rect 5200 560 5300 575
rect 5450 675 5550 690
rect 5450 575 5455 675
rect 5490 575 5510 675
rect 5545 575 5550 675
rect 5450 560 5550 575
rect 5700 675 5800 690
rect 5700 575 5705 675
rect 5740 575 5760 675
rect 5795 575 5800 675
rect 5700 560 5800 575
rect 5950 675 6050 690
rect 5950 575 5955 675
rect 5990 575 6010 675
rect 6045 575 6050 675
rect 5950 560 6050 575
rect 6200 675 6300 690
rect 6200 575 6205 675
rect 6240 575 6260 675
rect 6295 575 6300 675
rect 6200 560 6300 575
rect 6450 675 6550 690
rect 6450 575 6455 675
rect 6490 575 6510 675
rect 6545 575 6550 675
rect 6450 560 6550 575
rect 6700 675 6800 690
rect 6700 575 6705 675
rect 6740 575 6760 675
rect 6795 575 6800 675
rect 6700 560 6800 575
rect 6950 675 7050 690
rect 6950 575 6955 675
rect 6990 575 7010 675
rect 7045 575 7050 675
rect 6950 560 7050 575
rect 7200 675 7300 690
rect 7200 575 7205 675
rect 7240 575 7260 675
rect 7295 575 7300 675
rect 7200 560 7300 575
rect 7450 675 7550 690
rect 7450 575 7455 675
rect 7490 575 7510 675
rect 7545 575 7550 675
rect 7450 560 7550 575
rect 7700 675 7800 690
rect 7700 575 7705 675
rect 7740 575 7760 675
rect 7795 575 7800 675
rect 7700 560 7800 575
rect 7950 675 8000 690
rect 7950 575 7955 675
rect 7990 575 8000 675
rect 7950 560 8000 575
rect 0 550 60 560
rect 190 550 310 560
rect 440 550 560 560
rect 690 550 810 560
rect 940 550 1060 560
rect 1190 550 1310 560
rect 1440 550 1560 560
rect 1690 550 1810 560
rect 1940 550 2060 560
rect 2190 550 2310 560
rect 2440 550 2560 560
rect 2690 550 2810 560
rect 2940 550 3060 560
rect 3190 550 3310 560
rect 3440 550 3560 560
rect 3690 550 3810 560
rect 3940 550 4060 560
rect 4190 550 4310 560
rect 4440 550 4560 560
rect 4690 550 4810 560
rect 4940 550 5060 560
rect 5190 550 5310 560
rect 5440 550 5560 560
rect 5690 550 5810 560
rect 5940 550 6060 560
rect 6190 550 6310 560
rect 6440 550 6560 560
rect 6690 550 6810 560
rect 6940 550 7060 560
rect 7190 550 7310 560
rect 7440 550 7560 560
rect 7690 550 7810 560
rect 7940 550 8000 560
rect 0 545 200 550
rect 0 510 75 545
rect 175 510 200 545
rect 0 490 200 510
rect 0 455 75 490
rect 175 455 200 490
rect 0 450 200 455
rect 300 545 450 550
rect 300 510 325 545
rect 425 510 450 545
rect 300 490 450 510
rect 300 455 325 490
rect 425 455 450 490
rect 300 450 450 455
rect 550 545 700 550
rect 550 510 575 545
rect 675 510 700 545
rect 550 490 700 510
rect 550 455 575 490
rect 675 455 700 490
rect 550 450 700 455
rect 800 545 950 550
rect 800 510 825 545
rect 925 510 950 545
rect 800 490 950 510
rect 800 455 825 490
rect 925 455 950 490
rect 800 450 950 455
rect 1050 545 1200 550
rect 1050 510 1075 545
rect 1175 510 1200 545
rect 1050 490 1200 510
rect 1050 455 1075 490
rect 1175 455 1200 490
rect 1050 450 1200 455
rect 1300 545 1450 550
rect 1300 510 1325 545
rect 1425 510 1450 545
rect 1300 490 1450 510
rect 1300 455 1325 490
rect 1425 455 1450 490
rect 1300 450 1450 455
rect 1550 545 1700 550
rect 1550 510 1575 545
rect 1675 510 1700 545
rect 1550 490 1700 510
rect 1550 455 1575 490
rect 1675 455 1700 490
rect 1550 450 1700 455
rect 1800 545 2200 550
rect 1800 510 1825 545
rect 1925 510 2075 545
rect 2175 510 2200 545
rect 1800 490 2200 510
rect 1800 455 1825 490
rect 1925 455 2075 490
rect 2175 455 2200 490
rect 1800 450 2200 455
rect 2300 545 2450 550
rect 2300 510 2325 545
rect 2425 510 2450 545
rect 2300 490 2450 510
rect 2300 455 2325 490
rect 2425 455 2450 490
rect 2300 450 2450 455
rect 2550 545 2700 550
rect 2550 510 2575 545
rect 2675 510 2700 545
rect 2550 490 2700 510
rect 2550 455 2575 490
rect 2675 455 2700 490
rect 2550 450 2700 455
rect 2800 545 2950 550
rect 2800 510 2825 545
rect 2925 510 2950 545
rect 2800 490 2950 510
rect 2800 455 2825 490
rect 2925 455 2950 490
rect 2800 450 2950 455
rect 3050 545 3200 550
rect 3050 510 3075 545
rect 3175 510 3200 545
rect 3050 490 3200 510
rect 3050 455 3075 490
rect 3175 455 3200 490
rect 3050 450 3200 455
rect 3300 545 3450 550
rect 3300 510 3325 545
rect 3425 510 3450 545
rect 3300 490 3450 510
rect 3300 455 3325 490
rect 3425 455 3450 490
rect 3300 450 3450 455
rect 3550 545 3700 550
rect 3550 510 3575 545
rect 3675 510 3700 545
rect 3550 490 3700 510
rect 3550 455 3575 490
rect 3675 455 3700 490
rect 3550 450 3700 455
rect 3800 545 4200 550
rect 3800 510 3825 545
rect 3925 510 4075 545
rect 4175 510 4200 545
rect 3800 490 4200 510
rect 3800 455 3825 490
rect 3925 455 4075 490
rect 4175 455 4200 490
rect 3800 450 4200 455
rect 4300 545 4450 550
rect 4300 510 4325 545
rect 4425 510 4450 545
rect 4300 490 4450 510
rect 4300 455 4325 490
rect 4425 455 4450 490
rect 4300 450 4450 455
rect 4550 545 4700 550
rect 4550 510 4575 545
rect 4675 510 4700 545
rect 4550 490 4700 510
rect 4550 455 4575 490
rect 4675 455 4700 490
rect 4550 450 4700 455
rect 4800 545 4950 550
rect 4800 510 4825 545
rect 4925 510 4950 545
rect 4800 490 4950 510
rect 4800 455 4825 490
rect 4925 455 4950 490
rect 4800 450 4950 455
rect 5050 545 5200 550
rect 5050 510 5075 545
rect 5175 510 5200 545
rect 5050 490 5200 510
rect 5050 455 5075 490
rect 5175 455 5200 490
rect 5050 450 5200 455
rect 5300 545 5450 550
rect 5300 510 5325 545
rect 5425 510 5450 545
rect 5300 490 5450 510
rect 5300 455 5325 490
rect 5425 455 5450 490
rect 5300 450 5450 455
rect 5550 545 5700 550
rect 5550 510 5575 545
rect 5675 510 5700 545
rect 5550 490 5700 510
rect 5550 455 5575 490
rect 5675 455 5700 490
rect 5550 450 5700 455
rect 5800 545 6200 550
rect 5800 510 5825 545
rect 5925 510 6075 545
rect 6175 510 6200 545
rect 5800 490 6200 510
rect 5800 455 5825 490
rect 5925 455 6075 490
rect 6175 455 6200 490
rect 5800 450 6200 455
rect 6300 545 6450 550
rect 6300 510 6325 545
rect 6425 510 6450 545
rect 6300 490 6450 510
rect 6300 455 6325 490
rect 6425 455 6450 490
rect 6300 450 6450 455
rect 6550 545 6700 550
rect 6550 510 6575 545
rect 6675 510 6700 545
rect 6550 490 6700 510
rect 6550 455 6575 490
rect 6675 455 6700 490
rect 6550 450 6700 455
rect 6800 545 6950 550
rect 6800 510 6825 545
rect 6925 510 6950 545
rect 6800 490 6950 510
rect 6800 455 6825 490
rect 6925 455 6950 490
rect 6800 450 6950 455
rect 7050 545 7200 550
rect 7050 510 7075 545
rect 7175 510 7200 545
rect 7050 490 7200 510
rect 7050 455 7075 490
rect 7175 455 7200 490
rect 7050 450 7200 455
rect 7300 545 7450 550
rect 7300 510 7325 545
rect 7425 510 7450 545
rect 7300 490 7450 510
rect 7300 455 7325 490
rect 7425 455 7450 490
rect 7300 450 7450 455
rect 7550 545 7700 550
rect 7550 510 7575 545
rect 7675 510 7700 545
rect 7550 490 7700 510
rect 7550 455 7575 490
rect 7675 455 7700 490
rect 7550 450 7700 455
rect 7800 545 8000 550
rect 7800 510 7825 545
rect 7925 510 8000 545
rect 7800 490 8000 510
rect 7800 455 7825 490
rect 7925 455 8000 490
rect 7800 450 8000 455
rect 0 440 60 450
rect 190 440 310 450
rect 440 440 560 450
rect 690 440 810 450
rect 940 440 1060 450
rect 1190 440 1310 450
rect 1440 440 1560 450
rect 1690 440 1810 450
rect 1940 440 2060 450
rect 2190 440 2310 450
rect 2440 440 2560 450
rect 2690 440 2810 450
rect 2940 440 3060 450
rect 3190 440 3310 450
rect 3440 440 3560 450
rect 3690 440 3810 450
rect 3940 440 4060 450
rect 4190 440 4310 450
rect 4440 440 4560 450
rect 4690 440 4810 450
rect 4940 440 5060 450
rect 5190 440 5310 450
rect 5440 440 5560 450
rect 5690 440 5810 450
rect 5940 440 6060 450
rect 6190 440 6310 450
rect 6440 440 6560 450
rect 6690 440 6810 450
rect 6940 440 7060 450
rect 7190 440 7310 450
rect 7440 440 7560 450
rect 7690 440 7810 450
rect 7940 440 8000 450
rect 0 425 50 440
rect 0 325 10 425
rect 45 325 50 425
rect 0 310 50 325
rect 200 425 300 440
rect 200 325 205 425
rect 240 325 260 425
rect 295 325 300 425
rect 200 310 300 325
rect 450 425 550 440
rect 450 325 455 425
rect 490 325 510 425
rect 545 325 550 425
rect 450 310 550 325
rect 700 425 800 440
rect 700 325 705 425
rect 740 325 760 425
rect 795 325 800 425
rect 700 310 800 325
rect 950 425 1050 440
rect 950 325 955 425
rect 990 325 1010 425
rect 1045 325 1050 425
rect 950 310 1050 325
rect 1200 425 1300 440
rect 1200 325 1205 425
rect 1240 325 1260 425
rect 1295 325 1300 425
rect 1200 310 1300 325
rect 1450 425 1550 440
rect 1450 325 1455 425
rect 1490 325 1510 425
rect 1545 325 1550 425
rect 1450 310 1550 325
rect 1700 425 1800 440
rect 1700 325 1705 425
rect 1740 325 1760 425
rect 1795 325 1800 425
rect 1700 310 1800 325
rect 1950 425 2050 440
rect 1950 325 1955 425
rect 1990 325 2010 425
rect 2045 325 2050 425
rect 1950 310 2050 325
rect 2200 425 2300 440
rect 2200 325 2205 425
rect 2240 325 2260 425
rect 2295 325 2300 425
rect 2200 310 2300 325
rect 2450 425 2550 440
rect 2450 325 2455 425
rect 2490 325 2510 425
rect 2545 325 2550 425
rect 2450 310 2550 325
rect 2700 425 2800 440
rect 2700 325 2705 425
rect 2740 325 2760 425
rect 2795 325 2800 425
rect 2700 310 2800 325
rect 2950 425 3050 440
rect 2950 325 2955 425
rect 2990 325 3010 425
rect 3045 325 3050 425
rect 2950 310 3050 325
rect 3200 425 3300 440
rect 3200 325 3205 425
rect 3240 325 3260 425
rect 3295 325 3300 425
rect 3200 310 3300 325
rect 3450 425 3550 440
rect 3450 325 3455 425
rect 3490 325 3510 425
rect 3545 325 3550 425
rect 3450 310 3550 325
rect 3700 425 3800 440
rect 3700 325 3705 425
rect 3740 325 3760 425
rect 3795 325 3800 425
rect 3700 310 3800 325
rect 3950 425 4050 440
rect 3950 325 3955 425
rect 3990 325 4010 425
rect 4045 325 4050 425
rect 3950 310 4050 325
rect 4200 425 4300 440
rect 4200 325 4205 425
rect 4240 325 4260 425
rect 4295 325 4300 425
rect 4200 310 4300 325
rect 4450 425 4550 440
rect 4450 325 4455 425
rect 4490 325 4510 425
rect 4545 325 4550 425
rect 4450 310 4550 325
rect 4700 425 4800 440
rect 4700 325 4705 425
rect 4740 325 4760 425
rect 4795 325 4800 425
rect 4700 310 4800 325
rect 4950 425 5050 440
rect 4950 325 4955 425
rect 4990 325 5010 425
rect 5045 325 5050 425
rect 4950 310 5050 325
rect 5200 425 5300 440
rect 5200 325 5205 425
rect 5240 325 5260 425
rect 5295 325 5300 425
rect 5200 310 5300 325
rect 5450 425 5550 440
rect 5450 325 5455 425
rect 5490 325 5510 425
rect 5545 325 5550 425
rect 5450 310 5550 325
rect 5700 425 5800 440
rect 5700 325 5705 425
rect 5740 325 5760 425
rect 5795 325 5800 425
rect 5700 310 5800 325
rect 5950 425 6050 440
rect 5950 325 5955 425
rect 5990 325 6010 425
rect 6045 325 6050 425
rect 5950 310 6050 325
rect 6200 425 6300 440
rect 6200 325 6205 425
rect 6240 325 6260 425
rect 6295 325 6300 425
rect 6200 310 6300 325
rect 6450 425 6550 440
rect 6450 325 6455 425
rect 6490 325 6510 425
rect 6545 325 6550 425
rect 6450 310 6550 325
rect 6700 425 6800 440
rect 6700 325 6705 425
rect 6740 325 6760 425
rect 6795 325 6800 425
rect 6700 310 6800 325
rect 6950 425 7050 440
rect 6950 325 6955 425
rect 6990 325 7010 425
rect 7045 325 7050 425
rect 6950 310 7050 325
rect 7200 425 7300 440
rect 7200 325 7205 425
rect 7240 325 7260 425
rect 7295 325 7300 425
rect 7200 310 7300 325
rect 7450 425 7550 440
rect 7450 325 7455 425
rect 7490 325 7510 425
rect 7545 325 7550 425
rect 7450 310 7550 325
rect 7700 425 7800 440
rect 7700 325 7705 425
rect 7740 325 7760 425
rect 7795 325 7800 425
rect 7700 310 7800 325
rect 7950 425 8000 440
rect 7950 325 7955 425
rect 7990 325 8000 425
rect 7950 310 8000 325
rect 0 300 60 310
rect 190 300 310 310
rect 440 300 560 310
rect 690 300 810 310
rect 940 300 1060 310
rect 1190 300 1310 310
rect 1440 300 1560 310
rect 1690 300 1810 310
rect 1940 300 2060 310
rect 2190 300 2310 310
rect 2440 300 2560 310
rect 2690 300 2810 310
rect 2940 300 3060 310
rect 3190 300 3310 310
rect 3440 300 3560 310
rect 3690 300 3810 310
rect 3940 300 4060 310
rect 4190 300 4310 310
rect 4440 300 4560 310
rect 4690 300 4810 310
rect 4940 300 5060 310
rect 5190 300 5310 310
rect 5440 300 5560 310
rect 5690 300 5810 310
rect 5940 300 6060 310
rect 6190 300 6310 310
rect 6440 300 6560 310
rect 6690 300 6810 310
rect 6940 300 7060 310
rect 7190 300 7310 310
rect 7440 300 7560 310
rect 7690 300 7810 310
rect 7940 300 8000 310
rect 0 295 200 300
rect 0 260 75 295
rect 175 260 200 295
rect 0 240 200 260
rect 0 205 75 240
rect 175 205 200 240
rect 0 200 200 205
rect 300 295 450 300
rect 300 260 325 295
rect 425 260 450 295
rect 300 240 450 260
rect 300 205 325 240
rect 425 205 450 240
rect 300 200 450 205
rect 550 295 700 300
rect 550 260 575 295
rect 675 260 700 295
rect 550 240 700 260
rect 550 205 575 240
rect 675 205 700 240
rect 550 200 700 205
rect 800 295 1200 300
rect 800 260 825 295
rect 925 260 1075 295
rect 1175 260 1200 295
rect 800 240 1200 260
rect 800 205 825 240
rect 925 205 1075 240
rect 1175 205 1200 240
rect 800 200 1200 205
rect 1300 295 1450 300
rect 1300 260 1325 295
rect 1425 260 1450 295
rect 1300 240 1450 260
rect 1300 205 1325 240
rect 1425 205 1450 240
rect 1300 200 1450 205
rect 1550 295 1700 300
rect 1550 260 1575 295
rect 1675 260 1700 295
rect 1550 240 1700 260
rect 1550 205 1575 240
rect 1675 205 1700 240
rect 1550 200 1700 205
rect 1800 295 2200 300
rect 1800 260 1825 295
rect 1925 260 2075 295
rect 2175 260 2200 295
rect 1800 240 2200 260
rect 1800 205 1825 240
rect 1925 205 2075 240
rect 2175 205 2200 240
rect 1800 200 2200 205
rect 2300 295 2450 300
rect 2300 260 2325 295
rect 2425 260 2450 295
rect 2300 240 2450 260
rect 2300 205 2325 240
rect 2425 205 2450 240
rect 2300 200 2450 205
rect 2550 295 2700 300
rect 2550 260 2575 295
rect 2675 260 2700 295
rect 2550 240 2700 260
rect 2550 205 2575 240
rect 2675 205 2700 240
rect 2550 200 2700 205
rect 2800 295 3200 300
rect 2800 260 2825 295
rect 2925 260 3075 295
rect 3175 260 3200 295
rect 2800 240 3200 260
rect 2800 205 2825 240
rect 2925 205 3075 240
rect 3175 205 3200 240
rect 2800 200 3200 205
rect 3300 295 3450 300
rect 3300 260 3325 295
rect 3425 260 3450 295
rect 3300 240 3450 260
rect 3300 205 3325 240
rect 3425 205 3450 240
rect 3300 200 3450 205
rect 3550 295 3700 300
rect 3550 260 3575 295
rect 3675 260 3700 295
rect 3550 240 3700 260
rect 3550 205 3575 240
rect 3675 205 3700 240
rect 3550 200 3700 205
rect 3800 295 4200 300
rect 3800 260 3825 295
rect 3925 260 4075 295
rect 4175 260 4200 295
rect 3800 240 4200 260
rect 3800 205 3825 240
rect 3925 205 4075 240
rect 4175 205 4200 240
rect 3800 200 4200 205
rect 4300 295 4450 300
rect 4300 260 4325 295
rect 4425 260 4450 295
rect 4300 240 4450 260
rect 4300 205 4325 240
rect 4425 205 4450 240
rect 4300 200 4450 205
rect 4550 295 4700 300
rect 4550 260 4575 295
rect 4675 260 4700 295
rect 4550 240 4700 260
rect 4550 205 4575 240
rect 4675 205 4700 240
rect 4550 200 4700 205
rect 4800 295 5200 300
rect 4800 260 4825 295
rect 4925 260 5075 295
rect 5175 260 5200 295
rect 4800 240 5200 260
rect 4800 205 4825 240
rect 4925 205 5075 240
rect 5175 205 5200 240
rect 4800 200 5200 205
rect 5300 295 5450 300
rect 5300 260 5325 295
rect 5425 260 5450 295
rect 5300 240 5450 260
rect 5300 205 5325 240
rect 5425 205 5450 240
rect 5300 200 5450 205
rect 5550 295 5700 300
rect 5550 260 5575 295
rect 5675 260 5700 295
rect 5550 240 5700 260
rect 5550 205 5575 240
rect 5675 205 5700 240
rect 5550 200 5700 205
rect 5800 295 6200 300
rect 5800 260 5825 295
rect 5925 260 6075 295
rect 6175 260 6200 295
rect 5800 240 6200 260
rect 5800 205 5825 240
rect 5925 205 6075 240
rect 6175 205 6200 240
rect 5800 200 6200 205
rect 6300 295 6450 300
rect 6300 260 6325 295
rect 6425 260 6450 295
rect 6300 240 6450 260
rect 6300 205 6325 240
rect 6425 205 6450 240
rect 6300 200 6450 205
rect 6550 295 6700 300
rect 6550 260 6575 295
rect 6675 260 6700 295
rect 6550 240 6700 260
rect 6550 205 6575 240
rect 6675 205 6700 240
rect 6550 200 6700 205
rect 6800 295 7200 300
rect 6800 260 6825 295
rect 6925 260 7075 295
rect 7175 260 7200 295
rect 6800 240 7200 260
rect 6800 205 6825 240
rect 6925 205 7075 240
rect 7175 205 7200 240
rect 6800 200 7200 205
rect 7300 295 7450 300
rect 7300 260 7325 295
rect 7425 260 7450 295
rect 7300 240 7450 260
rect 7300 205 7325 240
rect 7425 205 7450 240
rect 7300 200 7450 205
rect 7550 295 7700 300
rect 7550 260 7575 295
rect 7675 260 7700 295
rect 7550 240 7700 260
rect 7550 205 7575 240
rect 7675 205 7700 240
rect 7550 200 7700 205
rect 7800 295 8000 300
rect 7800 260 7825 295
rect 7925 260 8000 295
rect 7800 240 8000 260
rect 7800 205 7825 240
rect 7925 205 8000 240
rect 7800 200 8000 205
rect 0 190 60 200
rect 190 190 310 200
rect 440 190 560 200
rect 690 190 810 200
rect 940 190 1060 200
rect 1190 190 1310 200
rect 1440 190 1560 200
rect 1690 190 1810 200
rect 1940 190 2060 200
rect 2190 190 2310 200
rect 2440 190 2560 200
rect 2690 190 2810 200
rect 2940 190 3060 200
rect 3190 190 3310 200
rect 3440 190 3560 200
rect 3690 190 3810 200
rect 3940 190 4060 200
rect 4190 190 4310 200
rect 4440 190 4560 200
rect 4690 190 4810 200
rect 4940 190 5060 200
rect 5190 190 5310 200
rect 5440 190 5560 200
rect 5690 190 5810 200
rect 5940 190 6060 200
rect 6190 190 6310 200
rect 6440 190 6560 200
rect 6690 190 6810 200
rect 6940 190 7060 200
rect 7190 190 7310 200
rect 7440 190 7560 200
rect 7690 190 7810 200
rect 7940 190 8000 200
rect 0 175 50 190
rect 0 75 10 175
rect 45 75 50 175
rect 0 60 50 75
rect 200 175 300 190
rect 200 75 205 175
rect 240 75 260 175
rect 295 75 300 175
rect 200 60 300 75
rect 450 175 550 190
rect 450 75 455 175
rect 490 75 510 175
rect 545 75 550 175
rect 450 60 550 75
rect 700 175 800 190
rect 700 75 705 175
rect 740 75 760 175
rect 795 75 800 175
rect 700 60 800 75
rect 950 175 1050 190
rect 950 75 955 175
rect 990 75 1010 175
rect 1045 75 1050 175
rect 950 60 1050 75
rect 1200 175 1300 190
rect 1200 75 1205 175
rect 1240 75 1260 175
rect 1295 75 1300 175
rect 1200 60 1300 75
rect 1450 175 1550 190
rect 1450 75 1455 175
rect 1490 75 1510 175
rect 1545 75 1550 175
rect 1450 60 1550 75
rect 1700 175 1800 190
rect 1700 75 1705 175
rect 1740 75 1760 175
rect 1795 75 1800 175
rect 1700 60 1800 75
rect 1950 175 2050 190
rect 1950 75 1955 175
rect 1990 75 2010 175
rect 2045 75 2050 175
rect 1950 60 2050 75
rect 2200 175 2300 190
rect 2200 75 2205 175
rect 2240 75 2260 175
rect 2295 75 2300 175
rect 2200 60 2300 75
rect 2450 175 2550 190
rect 2450 75 2455 175
rect 2490 75 2510 175
rect 2545 75 2550 175
rect 2450 60 2550 75
rect 2700 175 2800 190
rect 2700 75 2705 175
rect 2740 75 2760 175
rect 2795 75 2800 175
rect 2700 60 2800 75
rect 2950 175 3050 190
rect 2950 75 2955 175
rect 2990 75 3010 175
rect 3045 75 3050 175
rect 2950 60 3050 75
rect 3200 175 3300 190
rect 3200 75 3205 175
rect 3240 75 3260 175
rect 3295 75 3300 175
rect 3200 60 3300 75
rect 3450 175 3550 190
rect 3450 75 3455 175
rect 3490 75 3510 175
rect 3545 75 3550 175
rect 3450 60 3550 75
rect 3700 175 3800 190
rect 3700 75 3705 175
rect 3740 75 3760 175
rect 3795 75 3800 175
rect 3700 60 3800 75
rect 3950 175 4050 190
rect 3950 75 3955 175
rect 3990 75 4010 175
rect 4045 75 4050 175
rect 3950 60 4050 75
rect 4200 175 4300 190
rect 4200 75 4205 175
rect 4240 75 4260 175
rect 4295 75 4300 175
rect 4200 60 4300 75
rect 4450 175 4550 190
rect 4450 75 4455 175
rect 4490 75 4510 175
rect 4545 75 4550 175
rect 4450 60 4550 75
rect 4700 175 4800 190
rect 4700 75 4705 175
rect 4740 75 4760 175
rect 4795 75 4800 175
rect 4700 60 4800 75
rect 4950 175 5050 190
rect 4950 75 4955 175
rect 4990 75 5010 175
rect 5045 75 5050 175
rect 4950 60 5050 75
rect 5200 175 5300 190
rect 5200 75 5205 175
rect 5240 75 5260 175
rect 5295 75 5300 175
rect 5200 60 5300 75
rect 5450 175 5550 190
rect 5450 75 5455 175
rect 5490 75 5510 175
rect 5545 75 5550 175
rect 5450 60 5550 75
rect 5700 175 5800 190
rect 5700 75 5705 175
rect 5740 75 5760 175
rect 5795 75 5800 175
rect 5700 60 5800 75
rect 5950 175 6050 190
rect 5950 75 5955 175
rect 5990 75 6010 175
rect 6045 75 6050 175
rect 5950 60 6050 75
rect 6200 175 6300 190
rect 6200 75 6205 175
rect 6240 75 6260 175
rect 6295 75 6300 175
rect 6200 60 6300 75
rect 6450 175 6550 190
rect 6450 75 6455 175
rect 6490 75 6510 175
rect 6545 75 6550 175
rect 6450 60 6550 75
rect 6700 175 6800 190
rect 6700 75 6705 175
rect 6740 75 6760 175
rect 6795 75 6800 175
rect 6700 60 6800 75
rect 6950 175 7050 190
rect 6950 75 6955 175
rect 6990 75 7010 175
rect 7045 75 7050 175
rect 6950 60 7050 75
rect 7200 175 7300 190
rect 7200 75 7205 175
rect 7240 75 7260 175
rect 7295 75 7300 175
rect 7200 60 7300 75
rect 7450 175 7550 190
rect 7450 75 7455 175
rect 7490 75 7510 175
rect 7545 75 7550 175
rect 7450 60 7550 75
rect 7700 175 7800 190
rect 7700 75 7705 175
rect 7740 75 7760 175
rect 7795 75 7800 175
rect 7700 60 7800 75
rect 7950 175 8000 190
rect 7950 75 7955 175
rect 7990 75 8000 175
rect 7950 60 8000 75
rect 0 50 60 60
rect 190 50 310 60
rect 440 50 560 60
rect 690 50 810 60
rect 940 50 1060 60
rect 1190 50 1310 60
rect 1440 50 1560 60
rect 1690 50 1810 60
rect 1940 50 2060 60
rect 2190 50 2310 60
rect 2440 50 2560 60
rect 2690 50 2810 60
rect 2940 50 3060 60
rect 3190 50 3310 60
rect 3440 50 3560 60
rect 3690 50 3810 60
rect 3940 50 4060 60
rect 4190 50 4310 60
rect 4440 50 4560 60
rect 4690 50 4810 60
rect 4940 50 5060 60
rect 5190 50 5310 60
rect 5440 50 5560 60
rect 5690 50 5810 60
rect 5940 50 6060 60
rect 6190 50 6310 60
rect 6440 50 6560 60
rect 6690 50 6810 60
rect 6940 50 7060 60
rect 7190 50 7310 60
rect 7440 50 7560 60
rect 7690 50 7810 60
rect 7940 50 8000 60
rect 0 45 8000 50
rect 0 10 75 45
rect 175 10 325 45
rect 425 10 575 45
rect 675 10 825 45
rect 925 10 1075 45
rect 1175 10 1325 45
rect 1425 10 1575 45
rect 1675 10 1825 45
rect 1925 10 2075 45
rect 2175 10 2325 45
rect 2425 10 2575 45
rect 2675 10 2825 45
rect 2925 10 3075 45
rect 3175 10 3325 45
rect 3425 10 3575 45
rect 3675 10 3825 45
rect 3925 10 4075 45
rect 4175 10 4325 45
rect 4425 10 4575 45
rect 4675 10 4825 45
rect 4925 10 5075 45
rect 5175 10 5325 45
rect 5425 10 5575 45
rect 5675 10 5825 45
rect 5925 10 6075 45
rect 6175 10 6325 45
rect 6425 10 6575 45
rect 6675 10 6825 45
rect 6925 10 7075 45
rect 7175 10 7325 45
rect 7425 10 7575 45
rect 7675 10 7825 45
rect 7925 10 8000 45
rect 0 0 8000 10
<< via3 >>
rect 200 7700 300 7800
rect 450 7700 550 7800
rect 700 7700 800 7800
rect 1200 7700 1300 7800
rect 1450 7700 1550 7800
rect 1700 7700 1800 7800
rect 2200 7700 2300 7800
rect 2450 7700 2550 7800
rect 2700 7700 2800 7800
rect 3200 7700 3300 7800
rect 3450 7700 3550 7800
rect 3700 7700 3800 7800
rect 4200 7700 4300 7800
rect 4450 7700 4550 7800
rect 4700 7700 4800 7800
rect 5200 7700 5300 7800
rect 5450 7700 5550 7800
rect 5700 7700 5800 7800
rect 6200 7700 6300 7800
rect 6450 7700 6550 7800
rect 6700 7700 6800 7800
rect 7200 7700 7300 7800
rect 7450 7700 7550 7800
rect 7700 7700 7800 7800
rect 200 7450 300 7550
rect 450 7450 550 7550
rect 700 7450 800 7550
rect 950 7450 1050 7550
rect 1200 7450 1300 7550
rect 1450 7450 1550 7550
rect 1700 7450 1800 7550
rect 2200 7450 2300 7550
rect 2450 7450 2550 7550
rect 2700 7450 2800 7550
rect 2950 7450 3050 7550
rect 3200 7450 3300 7550
rect 3450 7450 3550 7550
rect 3700 7450 3800 7550
rect 4200 7450 4300 7550
rect 4450 7450 4550 7550
rect 4700 7450 4800 7550
rect 4950 7450 5050 7550
rect 5200 7450 5300 7550
rect 5450 7450 5550 7550
rect 5700 7450 5800 7550
rect 6200 7450 6300 7550
rect 6450 7450 6550 7550
rect 6700 7450 6800 7550
rect 6950 7450 7050 7550
rect 7200 7450 7300 7550
rect 7450 7450 7550 7550
rect 7700 7450 7800 7550
rect 200 7200 300 7300
rect 450 7200 550 7300
rect 700 7200 800 7300
rect 1200 7200 1300 7300
rect 1450 7200 1550 7300
rect 1700 7200 1800 7300
rect 2200 7200 2300 7300
rect 2450 7200 2550 7300
rect 2700 7200 2800 7300
rect 3200 7200 3300 7300
rect 3450 7200 3550 7300
rect 3700 7200 3800 7300
rect 4200 7200 4300 7300
rect 4450 7200 4550 7300
rect 4700 7200 4800 7300
rect 5200 7200 5300 7300
rect 5450 7200 5550 7300
rect 5700 7200 5800 7300
rect 6200 7200 6300 7300
rect 6450 7200 6550 7300
rect 6700 7200 6800 7300
rect 7200 7200 7300 7300
rect 7450 7200 7550 7300
rect 7700 7200 7800 7300
rect 450 6950 550 7050
rect 1450 6950 1550 7050
rect 2450 6950 2550 7050
rect 3450 6950 3550 7050
rect 4450 6950 4550 7050
rect 5450 6950 5550 7050
rect 6450 6950 6550 7050
rect 7450 6950 7550 7050
rect 200 6700 300 6800
rect 450 6700 550 6800
rect 700 6700 800 6800
rect 1200 6700 1300 6800
rect 1450 6700 1550 6800
rect 1700 6700 1800 6800
rect 2200 6700 2300 6800
rect 2450 6700 2550 6800
rect 2700 6700 2800 6800
rect 3200 6700 3300 6800
rect 3450 6700 3550 6800
rect 3700 6700 3800 6800
rect 4200 6700 4300 6800
rect 4450 6700 4550 6800
rect 4700 6700 4800 6800
rect 5200 6700 5300 6800
rect 5450 6700 5550 6800
rect 5700 6700 5800 6800
rect 6200 6700 6300 6800
rect 6450 6700 6550 6800
rect 6700 6700 6800 6800
rect 7200 6700 7300 6800
rect 7450 6700 7550 6800
rect 7700 6700 7800 6800
rect 200 6450 300 6550
rect 450 6450 550 6550
rect 700 6450 800 6550
rect 950 6450 1050 6550
rect 1200 6450 1300 6550
rect 1450 6450 1550 6550
rect 1700 6450 1800 6550
rect 2200 6450 2300 6550
rect 2450 6450 2550 6550
rect 2700 6450 2800 6550
rect 2950 6450 3050 6550
rect 3200 6450 3300 6550
rect 3450 6450 3550 6550
rect 3700 6450 3800 6550
rect 4200 6450 4300 6550
rect 4450 6450 4550 6550
rect 4700 6450 4800 6550
rect 4950 6450 5050 6550
rect 5200 6450 5300 6550
rect 5450 6450 5550 6550
rect 5700 6450 5800 6550
rect 6200 6450 6300 6550
rect 6450 6450 6550 6550
rect 6700 6450 6800 6550
rect 6950 6450 7050 6550
rect 7200 6450 7300 6550
rect 7450 6450 7550 6550
rect 7700 6450 7800 6550
rect 200 6200 300 6300
rect 450 6200 550 6300
rect 700 6200 800 6300
rect 1200 6200 1300 6300
rect 1450 6200 1550 6300
rect 1700 6200 1800 6300
rect 2200 6200 2300 6300
rect 2450 6200 2550 6300
rect 2700 6200 2800 6300
rect 3200 6200 3300 6300
rect 3450 6200 3550 6300
rect 3700 6200 3800 6300
rect 4200 6200 4300 6300
rect 4450 6200 4550 6300
rect 4700 6200 4800 6300
rect 5200 6200 5300 6300
rect 5450 6200 5550 6300
rect 5700 6200 5800 6300
rect 6200 6200 6300 6300
rect 6450 6200 6550 6300
rect 6700 6200 6800 6300
rect 7200 6200 7300 6300
rect 7450 6200 7550 6300
rect 7700 6200 7800 6300
rect 200 5700 300 5800
rect 450 5700 550 5800
rect 700 5700 800 5800
rect 1200 5700 1300 5800
rect 1450 5700 1550 5800
rect 1700 5700 1800 5800
rect 2200 5700 2300 5800
rect 2450 5700 2550 5800
rect 2700 5700 2800 5800
rect 3200 5700 3300 5800
rect 3450 5700 3550 5800
rect 3700 5700 3800 5800
rect 4200 5700 4300 5800
rect 4450 5700 4550 5800
rect 4700 5700 4800 5800
rect 5200 5700 5300 5800
rect 5450 5700 5550 5800
rect 5700 5700 5800 5800
rect 6200 5700 6300 5800
rect 6450 5700 6550 5800
rect 6700 5700 6800 5800
rect 7200 5700 7300 5800
rect 7450 5700 7550 5800
rect 7700 5700 7800 5800
rect 200 5450 300 5550
rect 450 5450 550 5550
rect 700 5450 800 5550
rect 950 5450 1050 5550
rect 1200 5450 1300 5550
rect 1450 5450 1550 5550
rect 1700 5450 1800 5550
rect 2200 5450 2300 5550
rect 2450 5450 2550 5550
rect 2700 5450 2800 5550
rect 2950 5450 3050 5550
rect 3200 5450 3300 5550
rect 3450 5450 3550 5550
rect 3700 5450 3800 5550
rect 4200 5450 4300 5550
rect 4450 5450 4550 5550
rect 4700 5450 4800 5550
rect 4950 5450 5050 5550
rect 5200 5450 5300 5550
rect 5450 5450 5550 5550
rect 5700 5450 5800 5550
rect 6200 5450 6300 5550
rect 6450 5450 6550 5550
rect 6700 5450 6800 5550
rect 6950 5450 7050 5550
rect 7200 5450 7300 5550
rect 7450 5450 7550 5550
rect 7700 5450 7800 5550
rect 200 5200 300 5300
rect 450 5200 550 5300
rect 700 5200 800 5300
rect 1200 5200 1300 5300
rect 1450 5200 1550 5300
rect 1700 5200 1800 5300
rect 2200 5200 2300 5300
rect 2450 5200 2550 5300
rect 2700 5200 2800 5300
rect 3200 5200 3300 5300
rect 3450 5200 3550 5300
rect 3700 5200 3800 5300
rect 4200 5200 4300 5300
rect 4450 5200 4550 5300
rect 4700 5200 4800 5300
rect 5200 5200 5300 5300
rect 5450 5200 5550 5300
rect 5700 5200 5800 5300
rect 6200 5200 6300 5300
rect 6450 5200 6550 5300
rect 6700 5200 6800 5300
rect 7200 5200 7300 5300
rect 7450 5200 7550 5300
rect 7700 5200 7800 5300
rect 450 4950 550 5050
rect 1450 4950 1550 5050
rect 2450 4950 2550 5050
rect 3450 4950 3550 5050
rect 4450 4950 4550 5050
rect 5450 4950 5550 5050
rect 6450 4950 6550 5050
rect 7450 4950 7550 5050
rect 200 4700 300 4800
rect 450 4700 550 4800
rect 700 4700 800 4800
rect 1200 4700 1300 4800
rect 1450 4700 1550 4800
rect 1700 4700 1800 4800
rect 2200 4700 2300 4800
rect 2450 4700 2550 4800
rect 2700 4700 2800 4800
rect 3200 4700 3300 4800
rect 3450 4700 3550 4800
rect 3700 4700 3800 4800
rect 4200 4700 4300 4800
rect 4450 4700 4550 4800
rect 4700 4700 4800 4800
rect 5200 4700 5300 4800
rect 5450 4700 5550 4800
rect 5700 4700 5800 4800
rect 6200 4700 6300 4800
rect 6450 4700 6550 4800
rect 6700 4700 6800 4800
rect 7200 4700 7300 4800
rect 7450 4700 7550 4800
rect 7700 4700 7800 4800
rect 200 4450 300 4550
rect 450 4450 550 4550
rect 700 4450 800 4550
rect 950 4450 1050 4550
rect 1200 4450 1300 4550
rect 1450 4450 1550 4550
rect 1700 4450 1800 4550
rect 2200 4450 2300 4550
rect 2450 4450 2550 4550
rect 2700 4450 2800 4550
rect 2950 4450 3050 4550
rect 3200 4450 3300 4550
rect 3450 4450 3550 4550
rect 3700 4450 3800 4550
rect 4200 4450 4300 4550
rect 4450 4450 4550 4550
rect 4700 4450 4800 4550
rect 4950 4450 5050 4550
rect 5200 4450 5300 4550
rect 5450 4450 5550 4550
rect 5700 4450 5800 4550
rect 6200 4450 6300 4550
rect 6450 4450 6550 4550
rect 6700 4450 6800 4550
rect 6950 4450 7050 4550
rect 7200 4450 7300 4550
rect 7450 4450 7550 4550
rect 7700 4450 7800 4550
rect 200 4200 300 4300
rect 450 4200 550 4300
rect 700 4200 800 4300
rect 1200 4200 1300 4300
rect 1450 4200 1550 4300
rect 1700 4200 1800 4300
rect 2200 4200 2300 4300
rect 2450 4200 2550 4300
rect 2700 4200 2800 4300
rect 3200 4200 3300 4300
rect 3450 4200 3550 4300
rect 3700 4200 3800 4300
rect 4200 4200 4300 4300
rect 4450 4200 4550 4300
rect 4700 4200 4800 4300
rect 5200 4200 5300 4300
rect 5450 4200 5550 4300
rect 5700 4200 5800 4300
rect 6200 4200 6300 4300
rect 6450 4200 6550 4300
rect 6700 4200 6800 4300
rect 7200 4200 7300 4300
rect 7450 4200 7550 4300
rect 7700 4200 7800 4300
rect 200 3700 300 3800
rect 450 3700 550 3800
rect 700 3700 800 3800
rect 1200 3700 1300 3800
rect 1450 3700 1550 3800
rect 1700 3700 1800 3800
rect 2200 3700 2300 3800
rect 2450 3700 2550 3800
rect 2700 3700 2800 3800
rect 3200 3700 3300 3800
rect 3450 3700 3550 3800
rect 3700 3700 3800 3800
rect 4200 3700 4300 3800
rect 4450 3700 4550 3800
rect 4700 3700 4800 3800
rect 5200 3700 5300 3800
rect 5450 3700 5550 3800
rect 5700 3700 5800 3800
rect 6200 3700 6300 3800
rect 6450 3700 6550 3800
rect 6700 3700 6800 3800
rect 7200 3700 7300 3800
rect 7450 3700 7550 3800
rect 7700 3700 7800 3800
rect 200 3450 300 3550
rect 450 3450 550 3550
rect 700 3450 800 3550
rect 950 3450 1050 3550
rect 1200 3450 1300 3550
rect 1450 3450 1550 3550
rect 1700 3450 1800 3550
rect 2200 3450 2300 3550
rect 2450 3450 2550 3550
rect 2700 3450 2800 3550
rect 2950 3450 3050 3550
rect 3200 3450 3300 3550
rect 3450 3450 3550 3550
rect 3700 3450 3800 3550
rect 4200 3450 4300 3550
rect 4450 3450 4550 3550
rect 4700 3450 4800 3550
rect 4950 3450 5050 3550
rect 5200 3450 5300 3550
rect 5450 3450 5550 3550
rect 5700 3450 5800 3550
rect 6200 3450 6300 3550
rect 6450 3450 6550 3550
rect 6700 3450 6800 3550
rect 6950 3450 7050 3550
rect 7200 3450 7300 3550
rect 7450 3450 7550 3550
rect 7700 3450 7800 3550
rect 200 3200 300 3300
rect 450 3200 550 3300
rect 700 3200 800 3300
rect 1200 3200 1300 3300
rect 1450 3200 1550 3300
rect 1700 3200 1800 3300
rect 2200 3200 2300 3300
rect 2450 3200 2550 3300
rect 2700 3200 2800 3300
rect 3200 3200 3300 3300
rect 3450 3200 3550 3300
rect 3700 3200 3800 3300
rect 4200 3200 4300 3300
rect 4450 3200 4550 3300
rect 4700 3200 4800 3300
rect 5200 3200 5300 3300
rect 5450 3200 5550 3300
rect 5700 3200 5800 3300
rect 6200 3200 6300 3300
rect 6450 3200 6550 3300
rect 6700 3200 6800 3300
rect 7200 3200 7300 3300
rect 7450 3200 7550 3300
rect 7700 3200 7800 3300
rect 450 2950 550 3050
rect 1450 2950 1550 3050
rect 2450 2950 2550 3050
rect 3450 2950 3550 3050
rect 4450 2950 4550 3050
rect 5450 2950 5550 3050
rect 6450 2950 6550 3050
rect 7450 2950 7550 3050
rect 200 2700 300 2800
rect 450 2700 550 2800
rect 700 2700 800 2800
rect 1200 2700 1300 2800
rect 1450 2700 1550 2800
rect 1700 2700 1800 2800
rect 2200 2700 2300 2800
rect 2450 2700 2550 2800
rect 2700 2700 2800 2800
rect 3200 2700 3300 2800
rect 3450 2700 3550 2800
rect 3700 2700 3800 2800
rect 4200 2700 4300 2800
rect 4450 2700 4550 2800
rect 4700 2700 4800 2800
rect 5200 2700 5300 2800
rect 5450 2700 5550 2800
rect 5700 2700 5800 2800
rect 6200 2700 6300 2800
rect 6450 2700 6550 2800
rect 6700 2700 6800 2800
rect 7200 2700 7300 2800
rect 7450 2700 7550 2800
rect 7700 2700 7800 2800
rect 200 2450 300 2550
rect 450 2450 550 2550
rect 700 2450 800 2550
rect 950 2450 1050 2550
rect 1200 2450 1300 2550
rect 1450 2450 1550 2550
rect 1700 2450 1800 2550
rect 2200 2450 2300 2550
rect 2450 2450 2550 2550
rect 2700 2450 2800 2550
rect 2950 2450 3050 2550
rect 3200 2450 3300 2550
rect 3450 2450 3550 2550
rect 3700 2450 3800 2550
rect 4200 2450 4300 2550
rect 4450 2450 4550 2550
rect 4700 2450 4800 2550
rect 4950 2450 5050 2550
rect 5200 2450 5300 2550
rect 5450 2450 5550 2550
rect 5700 2450 5800 2550
rect 6200 2450 6300 2550
rect 6450 2450 6550 2550
rect 6700 2450 6800 2550
rect 6950 2450 7050 2550
rect 7200 2450 7300 2550
rect 7450 2450 7550 2550
rect 7700 2450 7800 2550
rect 200 2200 300 2300
rect 450 2200 550 2300
rect 700 2200 800 2300
rect 1200 2200 1300 2300
rect 1450 2200 1550 2300
rect 1700 2200 1800 2300
rect 2200 2200 2300 2300
rect 2450 2200 2550 2300
rect 2700 2200 2800 2300
rect 3200 2200 3300 2300
rect 3450 2200 3550 2300
rect 3700 2200 3800 2300
rect 4200 2200 4300 2300
rect 4450 2200 4550 2300
rect 4700 2200 4800 2300
rect 5200 2200 5300 2300
rect 5450 2200 5550 2300
rect 5700 2200 5800 2300
rect 6200 2200 6300 2300
rect 6450 2200 6550 2300
rect 6700 2200 6800 2300
rect 7200 2200 7300 2300
rect 7450 2200 7550 2300
rect 7700 2200 7800 2300
rect 200 1700 300 1800
rect 450 1700 550 1800
rect 700 1700 800 1800
rect 1200 1700 1300 1800
rect 1450 1700 1550 1800
rect 1700 1700 1800 1800
rect 2200 1700 2300 1800
rect 2450 1700 2550 1800
rect 2700 1700 2800 1800
rect 3200 1700 3300 1800
rect 3450 1700 3550 1800
rect 3700 1700 3800 1800
rect 4200 1700 4300 1800
rect 4450 1700 4550 1800
rect 4700 1700 4800 1800
rect 5200 1700 5300 1800
rect 5450 1700 5550 1800
rect 5700 1700 5800 1800
rect 6200 1700 6300 1800
rect 6450 1700 6550 1800
rect 6700 1700 6800 1800
rect 7200 1700 7300 1800
rect 7450 1700 7550 1800
rect 7700 1700 7800 1800
rect 200 1450 300 1550
rect 450 1450 550 1550
rect 700 1450 800 1550
rect 950 1450 1050 1550
rect 1200 1450 1300 1550
rect 1450 1450 1550 1550
rect 1700 1450 1800 1550
rect 2200 1450 2300 1550
rect 2450 1450 2550 1550
rect 2700 1450 2800 1550
rect 2950 1450 3050 1550
rect 3200 1450 3300 1550
rect 3450 1450 3550 1550
rect 3700 1450 3800 1550
rect 4200 1450 4300 1550
rect 4450 1450 4550 1550
rect 4700 1450 4800 1550
rect 4950 1450 5050 1550
rect 5200 1450 5300 1550
rect 5450 1450 5550 1550
rect 5700 1450 5800 1550
rect 6200 1450 6300 1550
rect 6450 1450 6550 1550
rect 6700 1450 6800 1550
rect 6950 1450 7050 1550
rect 7200 1450 7300 1550
rect 7450 1450 7550 1550
rect 7700 1450 7800 1550
rect 200 1200 300 1300
rect 450 1200 550 1300
rect 700 1200 800 1300
rect 1200 1200 1300 1300
rect 1450 1200 1550 1300
rect 1700 1200 1800 1300
rect 2200 1200 2300 1300
rect 2450 1200 2550 1300
rect 2700 1200 2800 1300
rect 3200 1200 3300 1300
rect 3450 1200 3550 1300
rect 3700 1200 3800 1300
rect 4200 1200 4300 1300
rect 4450 1200 4550 1300
rect 4700 1200 4800 1300
rect 5200 1200 5300 1300
rect 5450 1200 5550 1300
rect 5700 1200 5800 1300
rect 6200 1200 6300 1300
rect 6450 1200 6550 1300
rect 6700 1200 6800 1300
rect 7200 1200 7300 1300
rect 7450 1200 7550 1300
rect 7700 1200 7800 1300
rect 450 950 550 1050
rect 1450 950 1550 1050
rect 2450 950 2550 1050
rect 3450 950 3550 1050
rect 4450 950 4550 1050
rect 5450 950 5550 1050
rect 6450 950 6550 1050
rect 7450 950 7550 1050
rect 200 700 300 800
rect 450 700 550 800
rect 700 700 800 800
rect 1200 700 1300 800
rect 1450 700 1550 800
rect 1700 700 1800 800
rect 2200 700 2300 800
rect 2450 700 2550 800
rect 2700 700 2800 800
rect 3200 700 3300 800
rect 3450 700 3550 800
rect 3700 700 3800 800
rect 4200 700 4300 800
rect 4450 700 4550 800
rect 4700 700 4800 800
rect 5200 700 5300 800
rect 5450 700 5550 800
rect 5700 700 5800 800
rect 6200 700 6300 800
rect 6450 700 6550 800
rect 6700 700 6800 800
rect 7200 700 7300 800
rect 7450 700 7550 800
rect 7700 700 7800 800
rect 200 450 300 550
rect 450 450 550 550
rect 700 450 800 550
rect 950 450 1050 550
rect 1200 450 1300 550
rect 1450 450 1550 550
rect 1700 450 1800 550
rect 2200 450 2300 550
rect 2450 450 2550 550
rect 2700 450 2800 550
rect 2950 450 3050 550
rect 3200 450 3300 550
rect 3450 450 3550 550
rect 3700 450 3800 550
rect 4200 450 4300 550
rect 4450 450 4550 550
rect 4700 450 4800 550
rect 4950 450 5050 550
rect 5200 450 5300 550
rect 5450 450 5550 550
rect 5700 450 5800 550
rect 6200 450 6300 550
rect 6450 450 6550 550
rect 6700 450 6800 550
rect 6950 450 7050 550
rect 7200 450 7300 550
rect 7450 450 7550 550
rect 7700 450 7800 550
rect 200 200 300 300
rect 450 200 550 300
rect 700 200 800 300
rect 1200 200 1300 300
rect 1450 200 1550 300
rect 1700 200 1800 300
rect 2200 200 2300 300
rect 2450 200 2550 300
rect 2700 200 2800 300
rect 3200 200 3300 300
rect 3450 200 3550 300
rect 3700 200 3800 300
rect 4200 200 4300 300
rect 4450 200 4550 300
rect 4700 200 4800 300
rect 5200 200 5300 300
rect 5450 200 5550 300
rect 5700 200 5800 300
rect 6200 200 6300 300
rect 6450 200 6550 300
rect 6700 200 6800 300
rect 7200 200 7300 300
rect 7450 200 7550 300
rect 7700 200 7800 300
<< metal4 >>
rect 260 7820 740 8000
rect 1260 7820 1740 8000
rect 2260 7820 2740 8000
rect 3260 7820 3740 8000
rect 4260 7820 4740 8000
rect 5260 7820 5740 8000
rect 6260 7820 6740 8000
rect 7260 7820 7740 8000
rect 180 7800 820 7820
rect 180 7740 200 7800
rect 0 7700 200 7740
rect 300 7700 450 7800
rect 550 7700 700 7800
rect 800 7740 820 7800
rect 1180 7800 1820 7820
rect 1180 7740 1200 7800
rect 800 7700 1200 7740
rect 1300 7700 1450 7800
rect 1550 7700 1700 7800
rect 1800 7740 1820 7800
rect 2180 7800 2820 7820
rect 2180 7740 2200 7800
rect 1800 7700 2200 7740
rect 2300 7700 2450 7800
rect 2550 7700 2700 7800
rect 2800 7740 2820 7800
rect 3180 7800 3820 7820
rect 3180 7740 3200 7800
rect 2800 7700 3200 7740
rect 3300 7700 3450 7800
rect 3550 7700 3700 7800
rect 3800 7740 3820 7800
rect 4180 7800 4820 7820
rect 4180 7740 4200 7800
rect 3800 7700 4200 7740
rect 4300 7700 4450 7800
rect 4550 7700 4700 7800
rect 4800 7740 4820 7800
rect 5180 7800 5820 7820
rect 5180 7740 5200 7800
rect 4800 7700 5200 7740
rect 5300 7700 5450 7800
rect 5550 7700 5700 7800
rect 5800 7740 5820 7800
rect 6180 7800 6820 7820
rect 6180 7740 6200 7800
rect 5800 7700 6200 7740
rect 6300 7700 6450 7800
rect 6550 7700 6700 7800
rect 6800 7740 6820 7800
rect 7180 7800 7820 7820
rect 7180 7740 7200 7800
rect 6800 7700 7200 7740
rect 7300 7700 7450 7800
rect 7550 7700 7700 7800
rect 7800 7740 7820 7800
rect 7800 7700 8000 7740
rect 0 7550 8000 7700
rect 0 7450 200 7550
rect 300 7450 450 7550
rect 550 7450 700 7550
rect 800 7450 950 7550
rect 1050 7450 1200 7550
rect 1300 7450 1450 7550
rect 1550 7450 1700 7550
rect 1800 7450 2200 7550
rect 2300 7450 2450 7550
rect 2550 7450 2700 7550
rect 2800 7450 2950 7550
rect 3050 7450 3200 7550
rect 3300 7450 3450 7550
rect 3550 7450 3700 7550
rect 3800 7450 4200 7550
rect 4300 7450 4450 7550
rect 4550 7450 4700 7550
rect 4800 7450 4950 7550
rect 5050 7450 5200 7550
rect 5300 7450 5450 7550
rect 5550 7450 5700 7550
rect 5800 7450 6200 7550
rect 6300 7450 6450 7550
rect 6550 7450 6700 7550
rect 6800 7450 6950 7550
rect 7050 7450 7200 7550
rect 7300 7450 7450 7550
rect 7550 7450 7700 7550
rect 7800 7450 8000 7550
rect 0 7300 8000 7450
rect 0 7260 200 7300
rect 180 7200 200 7260
rect 300 7200 450 7300
rect 550 7200 700 7300
rect 800 7260 1200 7300
rect 800 7200 820 7260
rect 180 7180 820 7200
rect 1180 7200 1200 7260
rect 1300 7200 1450 7300
rect 1550 7200 1700 7300
rect 1800 7260 2200 7300
rect 1800 7200 1820 7260
rect 1180 7180 1820 7200
rect 2180 7200 2200 7260
rect 2300 7200 2450 7300
rect 2550 7200 2700 7300
rect 2800 7260 3200 7300
rect 2800 7200 2820 7260
rect 2180 7180 2820 7200
rect 3180 7200 3200 7260
rect 3300 7200 3450 7300
rect 3550 7200 3700 7300
rect 3800 7260 4200 7300
rect 3800 7200 3820 7260
rect 3180 7180 3820 7200
rect 4180 7200 4200 7260
rect 4300 7200 4450 7300
rect 4550 7200 4700 7300
rect 4800 7260 5200 7300
rect 4800 7200 4820 7260
rect 4180 7180 4820 7200
rect 5180 7200 5200 7260
rect 5300 7200 5450 7300
rect 5550 7200 5700 7300
rect 5800 7260 6200 7300
rect 5800 7200 5820 7260
rect 5180 7180 5820 7200
rect 6180 7200 6200 7260
rect 6300 7200 6450 7300
rect 6550 7200 6700 7300
rect 6800 7260 7200 7300
rect 6800 7200 6820 7260
rect 6180 7180 6820 7200
rect 7180 7200 7200 7260
rect 7300 7200 7450 7300
rect 7550 7200 7700 7300
rect 7800 7260 8000 7300
rect 7800 7200 7820 7260
rect 7180 7180 7820 7200
rect 260 7050 740 7180
rect 260 6950 450 7050
rect 550 6950 740 7050
rect 260 6820 740 6950
rect 1260 7050 1740 7180
rect 1260 6950 1450 7050
rect 1550 6950 1740 7050
rect 1260 6820 1740 6950
rect 2260 7050 2740 7180
rect 2260 6950 2450 7050
rect 2550 6950 2740 7050
rect 2260 6820 2740 6950
rect 3260 7050 3740 7180
rect 3260 6950 3450 7050
rect 3550 6950 3740 7050
rect 3260 6820 3740 6950
rect 4260 7050 4740 7180
rect 4260 6950 4450 7050
rect 4550 6950 4740 7050
rect 4260 6820 4740 6950
rect 5260 7050 5740 7180
rect 5260 6950 5450 7050
rect 5550 6950 5740 7050
rect 5260 6820 5740 6950
rect 6260 7050 6740 7180
rect 6260 6950 6450 7050
rect 6550 6950 6740 7050
rect 6260 6820 6740 6950
rect 7260 7050 7740 7180
rect 7260 6950 7450 7050
rect 7550 6950 7740 7050
rect 7260 6820 7740 6950
rect 180 6800 820 6820
rect 180 6740 200 6800
rect 0 6700 200 6740
rect 300 6700 450 6800
rect 550 6700 700 6800
rect 800 6740 820 6800
rect 1180 6800 1820 6820
rect 1180 6740 1200 6800
rect 800 6700 1200 6740
rect 1300 6700 1450 6800
rect 1550 6700 1700 6800
rect 1800 6740 1820 6800
rect 2180 6800 2820 6820
rect 2180 6740 2200 6800
rect 1800 6700 2200 6740
rect 2300 6700 2450 6800
rect 2550 6700 2700 6800
rect 2800 6740 2820 6800
rect 3180 6800 3820 6820
rect 3180 6740 3200 6800
rect 2800 6700 3200 6740
rect 3300 6700 3450 6800
rect 3550 6700 3700 6800
rect 3800 6740 3820 6800
rect 4180 6800 4820 6820
rect 4180 6740 4200 6800
rect 3800 6700 4200 6740
rect 4300 6700 4450 6800
rect 4550 6700 4700 6800
rect 4800 6740 4820 6800
rect 5180 6800 5820 6820
rect 5180 6740 5200 6800
rect 4800 6700 5200 6740
rect 5300 6700 5450 6800
rect 5550 6700 5700 6800
rect 5800 6740 5820 6800
rect 6180 6800 6820 6820
rect 6180 6740 6200 6800
rect 5800 6700 6200 6740
rect 6300 6700 6450 6800
rect 6550 6700 6700 6800
rect 6800 6740 6820 6800
rect 7180 6800 7820 6820
rect 7180 6740 7200 6800
rect 6800 6700 7200 6740
rect 7300 6700 7450 6800
rect 7550 6700 7700 6800
rect 7800 6740 7820 6800
rect 7800 6700 8000 6740
rect 0 6550 8000 6700
rect 0 6450 200 6550
rect 300 6450 450 6550
rect 550 6450 700 6550
rect 800 6450 950 6550
rect 1050 6450 1200 6550
rect 1300 6450 1450 6550
rect 1550 6450 1700 6550
rect 1800 6450 2200 6550
rect 2300 6450 2450 6550
rect 2550 6450 2700 6550
rect 2800 6450 2950 6550
rect 3050 6450 3200 6550
rect 3300 6450 3450 6550
rect 3550 6450 3700 6550
rect 3800 6450 4200 6550
rect 4300 6450 4450 6550
rect 4550 6450 4700 6550
rect 4800 6450 4950 6550
rect 5050 6450 5200 6550
rect 5300 6450 5450 6550
rect 5550 6450 5700 6550
rect 5800 6450 6200 6550
rect 6300 6450 6450 6550
rect 6550 6450 6700 6550
rect 6800 6450 6950 6550
rect 7050 6450 7200 6550
rect 7300 6450 7450 6550
rect 7550 6450 7700 6550
rect 7800 6450 8000 6550
rect 0 6300 8000 6450
rect 0 6260 200 6300
rect 180 6200 200 6260
rect 300 6200 450 6300
rect 550 6200 700 6300
rect 800 6260 1200 6300
rect 800 6200 820 6260
rect 180 6180 820 6200
rect 1180 6200 1200 6260
rect 1300 6200 1450 6300
rect 1550 6200 1700 6300
rect 1800 6260 2200 6300
rect 1800 6200 1820 6260
rect 1180 6180 1820 6200
rect 2180 6200 2200 6260
rect 2300 6200 2450 6300
rect 2550 6200 2700 6300
rect 2800 6260 3200 6300
rect 2800 6200 2820 6260
rect 2180 6180 2820 6200
rect 3180 6200 3200 6260
rect 3300 6200 3450 6300
rect 3550 6200 3700 6300
rect 3800 6260 4200 6300
rect 3800 6200 3820 6260
rect 3180 6180 3820 6200
rect 4180 6200 4200 6260
rect 4300 6200 4450 6300
rect 4550 6200 4700 6300
rect 4800 6260 5200 6300
rect 4800 6200 4820 6260
rect 4180 6180 4820 6200
rect 5180 6200 5200 6260
rect 5300 6200 5450 6300
rect 5550 6200 5700 6300
rect 5800 6260 6200 6300
rect 5800 6200 5820 6260
rect 5180 6180 5820 6200
rect 6180 6200 6200 6260
rect 6300 6200 6450 6300
rect 6550 6200 6700 6300
rect 6800 6260 7200 6300
rect 6800 6200 6820 6260
rect 6180 6180 6820 6200
rect 7180 6200 7200 6260
rect 7300 6200 7450 6300
rect 7550 6200 7700 6300
rect 7800 6260 8000 6300
rect 7800 6200 7820 6260
rect 7180 6180 7820 6200
rect 260 5820 740 6180
rect 1260 5820 1740 6180
rect 2260 5820 2740 6180
rect 3260 5820 3740 6180
rect 4260 5820 4740 6180
rect 5260 5820 5740 6180
rect 6260 5820 6740 6180
rect 7260 5820 7740 6180
rect 180 5800 820 5820
rect 180 5740 200 5800
rect 0 5700 200 5740
rect 300 5700 450 5800
rect 550 5700 700 5800
rect 800 5740 820 5800
rect 1180 5800 1820 5820
rect 1180 5740 1200 5800
rect 800 5700 1200 5740
rect 1300 5700 1450 5800
rect 1550 5700 1700 5800
rect 1800 5740 1820 5800
rect 2180 5800 2820 5820
rect 2180 5740 2200 5800
rect 1800 5700 2200 5740
rect 2300 5700 2450 5800
rect 2550 5700 2700 5800
rect 2800 5740 2820 5800
rect 3180 5800 3820 5820
rect 3180 5740 3200 5800
rect 2800 5700 3200 5740
rect 3300 5700 3450 5800
rect 3550 5700 3700 5800
rect 3800 5740 3820 5800
rect 4180 5800 4820 5820
rect 4180 5740 4200 5800
rect 3800 5700 4200 5740
rect 4300 5700 4450 5800
rect 4550 5700 4700 5800
rect 4800 5740 4820 5800
rect 5180 5800 5820 5820
rect 5180 5740 5200 5800
rect 4800 5700 5200 5740
rect 5300 5700 5450 5800
rect 5550 5700 5700 5800
rect 5800 5740 5820 5800
rect 6180 5800 6820 5820
rect 6180 5740 6200 5800
rect 5800 5700 6200 5740
rect 6300 5700 6450 5800
rect 6550 5700 6700 5800
rect 6800 5740 6820 5800
rect 7180 5800 7820 5820
rect 7180 5740 7200 5800
rect 6800 5700 7200 5740
rect 7300 5700 7450 5800
rect 7550 5700 7700 5800
rect 7800 5740 7820 5800
rect 7800 5700 8000 5740
rect 0 5550 8000 5700
rect 0 5450 200 5550
rect 300 5450 450 5550
rect 550 5450 700 5550
rect 800 5450 950 5550
rect 1050 5450 1200 5550
rect 1300 5450 1450 5550
rect 1550 5450 1700 5550
rect 1800 5450 2200 5550
rect 2300 5450 2450 5550
rect 2550 5450 2700 5550
rect 2800 5450 2950 5550
rect 3050 5450 3200 5550
rect 3300 5450 3450 5550
rect 3550 5450 3700 5550
rect 3800 5450 4200 5550
rect 4300 5450 4450 5550
rect 4550 5450 4700 5550
rect 4800 5450 4950 5550
rect 5050 5450 5200 5550
rect 5300 5450 5450 5550
rect 5550 5450 5700 5550
rect 5800 5450 6200 5550
rect 6300 5450 6450 5550
rect 6550 5450 6700 5550
rect 6800 5450 6950 5550
rect 7050 5450 7200 5550
rect 7300 5450 7450 5550
rect 7550 5450 7700 5550
rect 7800 5450 8000 5550
rect 0 5300 8000 5450
rect 0 5260 200 5300
rect 180 5200 200 5260
rect 300 5200 450 5300
rect 550 5200 700 5300
rect 800 5260 1200 5300
rect 800 5200 820 5260
rect 180 5180 820 5200
rect 1180 5200 1200 5260
rect 1300 5200 1450 5300
rect 1550 5200 1700 5300
rect 1800 5260 2200 5300
rect 1800 5200 1820 5260
rect 1180 5180 1820 5200
rect 2180 5200 2200 5260
rect 2300 5200 2450 5300
rect 2550 5200 2700 5300
rect 2800 5260 3200 5300
rect 2800 5200 2820 5260
rect 2180 5180 2820 5200
rect 3180 5200 3200 5260
rect 3300 5200 3450 5300
rect 3550 5200 3700 5300
rect 3800 5260 4200 5300
rect 3800 5200 3820 5260
rect 3180 5180 3820 5200
rect 4180 5200 4200 5260
rect 4300 5200 4450 5300
rect 4550 5200 4700 5300
rect 4800 5260 5200 5300
rect 4800 5200 4820 5260
rect 4180 5180 4820 5200
rect 5180 5200 5200 5260
rect 5300 5200 5450 5300
rect 5550 5200 5700 5300
rect 5800 5260 6200 5300
rect 5800 5200 5820 5260
rect 5180 5180 5820 5200
rect 6180 5200 6200 5260
rect 6300 5200 6450 5300
rect 6550 5200 6700 5300
rect 6800 5260 7200 5300
rect 6800 5200 6820 5260
rect 6180 5180 6820 5200
rect 7180 5200 7200 5260
rect 7300 5200 7450 5300
rect 7550 5200 7700 5300
rect 7800 5260 8000 5300
rect 7800 5200 7820 5260
rect 7180 5180 7820 5200
rect 260 5050 740 5180
rect 260 4950 450 5050
rect 550 4950 740 5050
rect 260 4820 740 4950
rect 1260 5050 1740 5180
rect 1260 4950 1450 5050
rect 1550 4950 1740 5050
rect 1260 4820 1740 4950
rect 2260 5050 2740 5180
rect 2260 4950 2450 5050
rect 2550 4950 2740 5050
rect 2260 4820 2740 4950
rect 3260 5050 3740 5180
rect 3260 4950 3450 5050
rect 3550 4950 3740 5050
rect 3260 4820 3740 4950
rect 4260 5050 4740 5180
rect 4260 4950 4450 5050
rect 4550 4950 4740 5050
rect 4260 4820 4740 4950
rect 5260 5050 5740 5180
rect 5260 4950 5450 5050
rect 5550 4950 5740 5050
rect 5260 4820 5740 4950
rect 6260 5050 6740 5180
rect 6260 4950 6450 5050
rect 6550 4950 6740 5050
rect 6260 4820 6740 4950
rect 7260 5050 7740 5180
rect 7260 4950 7450 5050
rect 7550 4950 7740 5050
rect 7260 4820 7740 4950
rect 180 4800 820 4820
rect 180 4740 200 4800
rect 0 4700 200 4740
rect 300 4700 450 4800
rect 550 4700 700 4800
rect 800 4740 820 4800
rect 1180 4800 1820 4820
rect 1180 4740 1200 4800
rect 800 4700 1200 4740
rect 1300 4700 1450 4800
rect 1550 4700 1700 4800
rect 1800 4740 1820 4800
rect 2180 4800 2820 4820
rect 2180 4740 2200 4800
rect 1800 4700 2200 4740
rect 2300 4700 2450 4800
rect 2550 4700 2700 4800
rect 2800 4740 2820 4800
rect 3180 4800 3820 4820
rect 3180 4740 3200 4800
rect 2800 4700 3200 4740
rect 3300 4700 3450 4800
rect 3550 4700 3700 4800
rect 3800 4740 3820 4800
rect 4180 4800 4820 4820
rect 4180 4740 4200 4800
rect 3800 4700 4200 4740
rect 4300 4700 4450 4800
rect 4550 4700 4700 4800
rect 4800 4740 4820 4800
rect 5180 4800 5820 4820
rect 5180 4740 5200 4800
rect 4800 4700 5200 4740
rect 5300 4700 5450 4800
rect 5550 4700 5700 4800
rect 5800 4740 5820 4800
rect 6180 4800 6820 4820
rect 6180 4740 6200 4800
rect 5800 4700 6200 4740
rect 6300 4700 6450 4800
rect 6550 4700 6700 4800
rect 6800 4740 6820 4800
rect 7180 4800 7820 4820
rect 7180 4740 7200 4800
rect 6800 4700 7200 4740
rect 7300 4700 7450 4800
rect 7550 4700 7700 4800
rect 7800 4740 7820 4800
rect 7800 4700 8000 4740
rect 0 4550 8000 4700
rect 0 4450 200 4550
rect 300 4450 450 4550
rect 550 4450 700 4550
rect 800 4450 950 4550
rect 1050 4450 1200 4550
rect 1300 4450 1450 4550
rect 1550 4450 1700 4550
rect 1800 4450 2200 4550
rect 2300 4450 2450 4550
rect 2550 4450 2700 4550
rect 2800 4450 2950 4550
rect 3050 4450 3200 4550
rect 3300 4450 3450 4550
rect 3550 4450 3700 4550
rect 3800 4450 4200 4550
rect 4300 4450 4450 4550
rect 4550 4450 4700 4550
rect 4800 4450 4950 4550
rect 5050 4450 5200 4550
rect 5300 4450 5450 4550
rect 5550 4450 5700 4550
rect 5800 4450 6200 4550
rect 6300 4450 6450 4550
rect 6550 4450 6700 4550
rect 6800 4450 6950 4550
rect 7050 4450 7200 4550
rect 7300 4450 7450 4550
rect 7550 4450 7700 4550
rect 7800 4450 8000 4550
rect 0 4300 8000 4450
rect 0 4260 200 4300
rect 180 4200 200 4260
rect 300 4200 450 4300
rect 550 4200 700 4300
rect 800 4260 1200 4300
rect 800 4200 820 4260
rect 180 4180 820 4200
rect 1180 4200 1200 4260
rect 1300 4200 1450 4300
rect 1550 4200 1700 4300
rect 1800 4260 2200 4300
rect 1800 4200 1820 4260
rect 1180 4180 1820 4200
rect 2180 4200 2200 4260
rect 2300 4200 2450 4300
rect 2550 4200 2700 4300
rect 2800 4260 3200 4300
rect 2800 4200 2820 4260
rect 2180 4180 2820 4200
rect 3180 4200 3200 4260
rect 3300 4200 3450 4300
rect 3550 4200 3700 4300
rect 3800 4260 4200 4300
rect 3800 4200 3820 4260
rect 3180 4180 3820 4200
rect 4180 4200 4200 4260
rect 4300 4200 4450 4300
rect 4550 4200 4700 4300
rect 4800 4260 5200 4300
rect 4800 4200 4820 4260
rect 4180 4180 4820 4200
rect 5180 4200 5200 4260
rect 5300 4200 5450 4300
rect 5550 4200 5700 4300
rect 5800 4260 6200 4300
rect 5800 4200 5820 4260
rect 5180 4180 5820 4200
rect 6180 4200 6200 4260
rect 6300 4200 6450 4300
rect 6550 4200 6700 4300
rect 6800 4260 7200 4300
rect 6800 4200 6820 4260
rect 6180 4180 6820 4200
rect 7180 4200 7200 4260
rect 7300 4200 7450 4300
rect 7550 4200 7700 4300
rect 7800 4260 8000 4300
rect 7800 4200 7820 4260
rect 7180 4180 7820 4200
rect 260 3820 740 4180
rect 1260 3820 1740 4180
rect 2260 3820 2740 4180
rect 3260 3820 3740 4180
rect 4260 3820 4740 4180
rect 5260 3820 5740 4180
rect 6260 3820 6740 4180
rect 7260 3820 7740 4180
rect 180 3800 820 3820
rect 180 3740 200 3800
rect 0 3700 200 3740
rect 300 3700 450 3800
rect 550 3700 700 3800
rect 800 3740 820 3800
rect 1180 3800 1820 3820
rect 1180 3740 1200 3800
rect 800 3700 1200 3740
rect 1300 3700 1450 3800
rect 1550 3700 1700 3800
rect 1800 3740 1820 3800
rect 2180 3800 2820 3820
rect 2180 3740 2200 3800
rect 1800 3700 2200 3740
rect 2300 3700 2450 3800
rect 2550 3700 2700 3800
rect 2800 3740 2820 3800
rect 3180 3800 3820 3820
rect 3180 3740 3200 3800
rect 2800 3700 3200 3740
rect 3300 3700 3450 3800
rect 3550 3700 3700 3800
rect 3800 3740 3820 3800
rect 4180 3800 4820 3820
rect 4180 3740 4200 3800
rect 3800 3700 4200 3740
rect 4300 3700 4450 3800
rect 4550 3700 4700 3800
rect 4800 3740 4820 3800
rect 5180 3800 5820 3820
rect 5180 3740 5200 3800
rect 4800 3700 5200 3740
rect 5300 3700 5450 3800
rect 5550 3700 5700 3800
rect 5800 3740 5820 3800
rect 6180 3800 6820 3820
rect 6180 3740 6200 3800
rect 5800 3700 6200 3740
rect 6300 3700 6450 3800
rect 6550 3700 6700 3800
rect 6800 3740 6820 3800
rect 7180 3800 7820 3820
rect 7180 3740 7200 3800
rect 6800 3700 7200 3740
rect 7300 3700 7450 3800
rect 7550 3700 7700 3800
rect 7800 3740 7820 3800
rect 7800 3700 8000 3740
rect 0 3550 8000 3700
rect 0 3450 200 3550
rect 300 3450 450 3550
rect 550 3450 700 3550
rect 800 3450 950 3550
rect 1050 3450 1200 3550
rect 1300 3450 1450 3550
rect 1550 3450 1700 3550
rect 1800 3450 2200 3550
rect 2300 3450 2450 3550
rect 2550 3450 2700 3550
rect 2800 3450 2950 3550
rect 3050 3450 3200 3550
rect 3300 3450 3450 3550
rect 3550 3450 3700 3550
rect 3800 3450 4200 3550
rect 4300 3450 4450 3550
rect 4550 3450 4700 3550
rect 4800 3450 4950 3550
rect 5050 3450 5200 3550
rect 5300 3450 5450 3550
rect 5550 3450 5700 3550
rect 5800 3450 6200 3550
rect 6300 3450 6450 3550
rect 6550 3450 6700 3550
rect 6800 3450 6950 3550
rect 7050 3450 7200 3550
rect 7300 3450 7450 3550
rect 7550 3450 7700 3550
rect 7800 3450 8000 3550
rect 0 3300 8000 3450
rect 0 3260 200 3300
rect 180 3200 200 3260
rect 300 3200 450 3300
rect 550 3200 700 3300
rect 800 3260 1200 3300
rect 800 3200 820 3260
rect 180 3180 820 3200
rect 1180 3200 1200 3260
rect 1300 3200 1450 3300
rect 1550 3200 1700 3300
rect 1800 3260 2200 3300
rect 1800 3200 1820 3260
rect 1180 3180 1820 3200
rect 2180 3200 2200 3260
rect 2300 3200 2450 3300
rect 2550 3200 2700 3300
rect 2800 3260 3200 3300
rect 2800 3200 2820 3260
rect 2180 3180 2820 3200
rect 3180 3200 3200 3260
rect 3300 3200 3450 3300
rect 3550 3200 3700 3300
rect 3800 3260 4200 3300
rect 3800 3200 3820 3260
rect 3180 3180 3820 3200
rect 4180 3200 4200 3260
rect 4300 3200 4450 3300
rect 4550 3200 4700 3300
rect 4800 3260 5200 3300
rect 4800 3200 4820 3260
rect 4180 3180 4820 3200
rect 5180 3200 5200 3260
rect 5300 3200 5450 3300
rect 5550 3200 5700 3300
rect 5800 3260 6200 3300
rect 5800 3200 5820 3260
rect 5180 3180 5820 3200
rect 6180 3200 6200 3260
rect 6300 3200 6450 3300
rect 6550 3200 6700 3300
rect 6800 3260 7200 3300
rect 6800 3200 6820 3260
rect 6180 3180 6820 3200
rect 7180 3200 7200 3260
rect 7300 3200 7450 3300
rect 7550 3200 7700 3300
rect 7800 3260 8000 3300
rect 7800 3200 7820 3260
rect 7180 3180 7820 3200
rect 260 3050 740 3180
rect 260 2950 450 3050
rect 550 2950 740 3050
rect 260 2820 740 2950
rect 1260 3050 1740 3180
rect 1260 2950 1450 3050
rect 1550 2950 1740 3050
rect 1260 2820 1740 2950
rect 2260 3050 2740 3180
rect 2260 2950 2450 3050
rect 2550 2950 2740 3050
rect 2260 2820 2740 2950
rect 3260 3050 3740 3180
rect 3260 2950 3450 3050
rect 3550 2950 3740 3050
rect 3260 2820 3740 2950
rect 4260 3050 4740 3180
rect 4260 2950 4450 3050
rect 4550 2950 4740 3050
rect 4260 2820 4740 2950
rect 5260 3050 5740 3180
rect 5260 2950 5450 3050
rect 5550 2950 5740 3050
rect 5260 2820 5740 2950
rect 6260 3050 6740 3180
rect 6260 2950 6450 3050
rect 6550 2950 6740 3050
rect 6260 2820 6740 2950
rect 7260 3050 7740 3180
rect 7260 2950 7450 3050
rect 7550 2950 7740 3050
rect 7260 2820 7740 2950
rect 180 2800 820 2820
rect 180 2740 200 2800
rect 0 2700 200 2740
rect 300 2700 450 2800
rect 550 2700 700 2800
rect 800 2740 820 2800
rect 1180 2800 1820 2820
rect 1180 2740 1200 2800
rect 800 2700 1200 2740
rect 1300 2700 1450 2800
rect 1550 2700 1700 2800
rect 1800 2740 1820 2800
rect 2180 2800 2820 2820
rect 2180 2740 2200 2800
rect 1800 2700 2200 2740
rect 2300 2700 2450 2800
rect 2550 2700 2700 2800
rect 2800 2740 2820 2800
rect 3180 2800 3820 2820
rect 3180 2740 3200 2800
rect 2800 2700 3200 2740
rect 3300 2700 3450 2800
rect 3550 2700 3700 2800
rect 3800 2740 3820 2800
rect 4180 2800 4820 2820
rect 4180 2740 4200 2800
rect 3800 2700 4200 2740
rect 4300 2700 4450 2800
rect 4550 2700 4700 2800
rect 4800 2740 4820 2800
rect 5180 2800 5820 2820
rect 5180 2740 5200 2800
rect 4800 2700 5200 2740
rect 5300 2700 5450 2800
rect 5550 2700 5700 2800
rect 5800 2740 5820 2800
rect 6180 2800 6820 2820
rect 6180 2740 6200 2800
rect 5800 2700 6200 2740
rect 6300 2700 6450 2800
rect 6550 2700 6700 2800
rect 6800 2740 6820 2800
rect 7180 2800 7820 2820
rect 7180 2740 7200 2800
rect 6800 2700 7200 2740
rect 7300 2700 7450 2800
rect 7550 2700 7700 2800
rect 7800 2740 7820 2800
rect 7800 2700 8000 2740
rect 0 2550 8000 2700
rect 0 2450 200 2550
rect 300 2450 450 2550
rect 550 2450 700 2550
rect 800 2450 950 2550
rect 1050 2450 1200 2550
rect 1300 2450 1450 2550
rect 1550 2450 1700 2550
rect 1800 2450 2200 2550
rect 2300 2450 2450 2550
rect 2550 2450 2700 2550
rect 2800 2450 2950 2550
rect 3050 2450 3200 2550
rect 3300 2450 3450 2550
rect 3550 2450 3700 2550
rect 3800 2450 4200 2550
rect 4300 2450 4450 2550
rect 4550 2450 4700 2550
rect 4800 2450 4950 2550
rect 5050 2450 5200 2550
rect 5300 2450 5450 2550
rect 5550 2450 5700 2550
rect 5800 2450 6200 2550
rect 6300 2450 6450 2550
rect 6550 2450 6700 2550
rect 6800 2450 6950 2550
rect 7050 2450 7200 2550
rect 7300 2450 7450 2550
rect 7550 2450 7700 2550
rect 7800 2450 8000 2550
rect 0 2300 8000 2450
rect 0 2260 200 2300
rect 180 2200 200 2260
rect 300 2200 450 2300
rect 550 2200 700 2300
rect 800 2260 1200 2300
rect 800 2200 820 2260
rect 180 2180 820 2200
rect 1180 2200 1200 2260
rect 1300 2200 1450 2300
rect 1550 2200 1700 2300
rect 1800 2260 2200 2300
rect 1800 2200 1820 2260
rect 1180 2180 1820 2200
rect 2180 2200 2200 2260
rect 2300 2200 2450 2300
rect 2550 2200 2700 2300
rect 2800 2260 3200 2300
rect 2800 2200 2820 2260
rect 2180 2180 2820 2200
rect 3180 2200 3200 2260
rect 3300 2200 3450 2300
rect 3550 2200 3700 2300
rect 3800 2260 4200 2300
rect 3800 2200 3820 2260
rect 3180 2180 3820 2200
rect 4180 2200 4200 2260
rect 4300 2200 4450 2300
rect 4550 2200 4700 2300
rect 4800 2260 5200 2300
rect 4800 2200 4820 2260
rect 4180 2180 4820 2200
rect 5180 2200 5200 2260
rect 5300 2200 5450 2300
rect 5550 2200 5700 2300
rect 5800 2260 6200 2300
rect 5800 2200 5820 2260
rect 5180 2180 5820 2200
rect 6180 2200 6200 2260
rect 6300 2200 6450 2300
rect 6550 2200 6700 2300
rect 6800 2260 7200 2300
rect 6800 2200 6820 2260
rect 6180 2180 6820 2200
rect 7180 2200 7200 2260
rect 7300 2200 7450 2300
rect 7550 2200 7700 2300
rect 7800 2260 8000 2300
rect 7800 2200 7820 2260
rect 7180 2180 7820 2200
rect 260 1820 740 2180
rect 1260 1820 1740 2180
rect 2260 1820 2740 2180
rect 3260 1820 3740 2180
rect 4260 1820 4740 2180
rect 5260 1820 5740 2180
rect 6260 1820 6740 2180
rect 7260 1820 7740 2180
rect 180 1800 820 1820
rect 180 1740 200 1800
rect 0 1700 200 1740
rect 300 1700 450 1800
rect 550 1700 700 1800
rect 800 1740 820 1800
rect 1180 1800 1820 1820
rect 1180 1740 1200 1800
rect 800 1700 1200 1740
rect 1300 1700 1450 1800
rect 1550 1700 1700 1800
rect 1800 1740 1820 1800
rect 2180 1800 2820 1820
rect 2180 1740 2200 1800
rect 1800 1700 2200 1740
rect 2300 1700 2450 1800
rect 2550 1700 2700 1800
rect 2800 1740 2820 1800
rect 3180 1800 3820 1820
rect 3180 1740 3200 1800
rect 2800 1700 3200 1740
rect 3300 1700 3450 1800
rect 3550 1700 3700 1800
rect 3800 1740 3820 1800
rect 4180 1800 4820 1820
rect 4180 1740 4200 1800
rect 3800 1700 4200 1740
rect 4300 1700 4450 1800
rect 4550 1700 4700 1800
rect 4800 1740 4820 1800
rect 5180 1800 5820 1820
rect 5180 1740 5200 1800
rect 4800 1700 5200 1740
rect 5300 1700 5450 1800
rect 5550 1700 5700 1800
rect 5800 1740 5820 1800
rect 6180 1800 6820 1820
rect 6180 1740 6200 1800
rect 5800 1700 6200 1740
rect 6300 1700 6450 1800
rect 6550 1700 6700 1800
rect 6800 1740 6820 1800
rect 7180 1800 7820 1820
rect 7180 1740 7200 1800
rect 6800 1700 7200 1740
rect 7300 1700 7450 1800
rect 7550 1700 7700 1800
rect 7800 1740 7820 1800
rect 7800 1700 8000 1740
rect 0 1550 8000 1700
rect 0 1450 200 1550
rect 300 1450 450 1550
rect 550 1450 700 1550
rect 800 1450 950 1550
rect 1050 1450 1200 1550
rect 1300 1450 1450 1550
rect 1550 1450 1700 1550
rect 1800 1450 2200 1550
rect 2300 1450 2450 1550
rect 2550 1450 2700 1550
rect 2800 1450 2950 1550
rect 3050 1450 3200 1550
rect 3300 1450 3450 1550
rect 3550 1450 3700 1550
rect 3800 1450 4200 1550
rect 4300 1450 4450 1550
rect 4550 1450 4700 1550
rect 4800 1450 4950 1550
rect 5050 1450 5200 1550
rect 5300 1450 5450 1550
rect 5550 1450 5700 1550
rect 5800 1450 6200 1550
rect 6300 1450 6450 1550
rect 6550 1450 6700 1550
rect 6800 1450 6950 1550
rect 7050 1450 7200 1550
rect 7300 1450 7450 1550
rect 7550 1450 7700 1550
rect 7800 1450 8000 1550
rect 0 1300 8000 1450
rect 0 1260 200 1300
rect 180 1200 200 1260
rect 300 1200 450 1300
rect 550 1200 700 1300
rect 800 1260 1200 1300
rect 800 1200 820 1260
rect 180 1180 820 1200
rect 1180 1200 1200 1260
rect 1300 1200 1450 1300
rect 1550 1200 1700 1300
rect 1800 1260 2200 1300
rect 1800 1200 1820 1260
rect 1180 1180 1820 1200
rect 2180 1200 2200 1260
rect 2300 1200 2450 1300
rect 2550 1200 2700 1300
rect 2800 1260 3200 1300
rect 2800 1200 2820 1260
rect 2180 1180 2820 1200
rect 3180 1200 3200 1260
rect 3300 1200 3450 1300
rect 3550 1200 3700 1300
rect 3800 1260 4200 1300
rect 3800 1200 3820 1260
rect 3180 1180 3820 1200
rect 4180 1200 4200 1260
rect 4300 1200 4450 1300
rect 4550 1200 4700 1300
rect 4800 1260 5200 1300
rect 4800 1200 4820 1260
rect 4180 1180 4820 1200
rect 5180 1200 5200 1260
rect 5300 1200 5450 1300
rect 5550 1200 5700 1300
rect 5800 1260 6200 1300
rect 5800 1200 5820 1260
rect 5180 1180 5820 1200
rect 6180 1200 6200 1260
rect 6300 1200 6450 1300
rect 6550 1200 6700 1300
rect 6800 1260 7200 1300
rect 6800 1200 6820 1260
rect 6180 1180 6820 1200
rect 7180 1200 7200 1260
rect 7300 1200 7450 1300
rect 7550 1200 7700 1300
rect 7800 1260 8000 1300
rect 7800 1200 7820 1260
rect 7180 1180 7820 1200
rect 260 1050 740 1180
rect 260 950 450 1050
rect 550 950 740 1050
rect 260 820 740 950
rect 1260 1050 1740 1180
rect 1260 950 1450 1050
rect 1550 950 1740 1050
rect 1260 820 1740 950
rect 2260 1050 2740 1180
rect 2260 950 2450 1050
rect 2550 950 2740 1050
rect 2260 820 2740 950
rect 3260 1050 3740 1180
rect 3260 950 3450 1050
rect 3550 950 3740 1050
rect 3260 820 3740 950
rect 4260 1050 4740 1180
rect 4260 950 4450 1050
rect 4550 950 4740 1050
rect 4260 820 4740 950
rect 5260 1050 5740 1180
rect 5260 950 5450 1050
rect 5550 950 5740 1050
rect 5260 820 5740 950
rect 6260 1050 6740 1180
rect 6260 950 6450 1050
rect 6550 950 6740 1050
rect 6260 820 6740 950
rect 7260 1050 7740 1180
rect 7260 950 7450 1050
rect 7550 950 7740 1050
rect 7260 820 7740 950
rect 180 800 820 820
rect 180 740 200 800
rect 0 700 200 740
rect 300 700 450 800
rect 550 700 700 800
rect 800 740 820 800
rect 1180 800 1820 820
rect 1180 740 1200 800
rect 800 700 1200 740
rect 1300 700 1450 800
rect 1550 700 1700 800
rect 1800 740 1820 800
rect 2180 800 2820 820
rect 2180 740 2200 800
rect 1800 700 2200 740
rect 2300 700 2450 800
rect 2550 700 2700 800
rect 2800 740 2820 800
rect 3180 800 3820 820
rect 3180 740 3200 800
rect 2800 700 3200 740
rect 3300 700 3450 800
rect 3550 700 3700 800
rect 3800 740 3820 800
rect 4180 800 4820 820
rect 4180 740 4200 800
rect 3800 700 4200 740
rect 4300 700 4450 800
rect 4550 700 4700 800
rect 4800 740 4820 800
rect 5180 800 5820 820
rect 5180 740 5200 800
rect 4800 700 5200 740
rect 5300 700 5450 800
rect 5550 700 5700 800
rect 5800 740 5820 800
rect 6180 800 6820 820
rect 6180 740 6200 800
rect 5800 700 6200 740
rect 6300 700 6450 800
rect 6550 700 6700 800
rect 6800 740 6820 800
rect 7180 800 7820 820
rect 7180 740 7200 800
rect 6800 700 7200 740
rect 7300 700 7450 800
rect 7550 700 7700 800
rect 7800 740 7820 800
rect 7800 700 8000 740
rect 0 550 8000 700
rect 0 450 200 550
rect 300 450 450 550
rect 550 450 700 550
rect 800 450 950 550
rect 1050 450 1200 550
rect 1300 450 1450 550
rect 1550 450 1700 550
rect 1800 450 2200 550
rect 2300 450 2450 550
rect 2550 450 2700 550
rect 2800 450 2950 550
rect 3050 450 3200 550
rect 3300 450 3450 550
rect 3550 450 3700 550
rect 3800 450 4200 550
rect 4300 450 4450 550
rect 4550 450 4700 550
rect 4800 450 4950 550
rect 5050 450 5200 550
rect 5300 450 5450 550
rect 5550 450 5700 550
rect 5800 450 6200 550
rect 6300 450 6450 550
rect 6550 450 6700 550
rect 6800 450 6950 550
rect 7050 450 7200 550
rect 7300 450 7450 550
rect 7550 450 7700 550
rect 7800 450 8000 550
rect 0 300 8000 450
rect 0 260 200 300
rect 180 200 200 260
rect 300 200 450 300
rect 550 200 700 300
rect 800 260 1200 300
rect 800 200 820 260
rect 180 180 820 200
rect 1180 200 1200 260
rect 1300 200 1450 300
rect 1550 200 1700 300
rect 1800 260 2200 300
rect 1800 200 1820 260
rect 1180 180 1820 200
rect 2180 200 2200 260
rect 2300 200 2450 300
rect 2550 200 2700 300
rect 2800 260 3200 300
rect 2800 200 2820 260
rect 2180 180 2820 200
rect 3180 200 3200 260
rect 3300 200 3450 300
rect 3550 200 3700 300
rect 3800 260 4200 300
rect 3800 200 3820 260
rect 3180 180 3820 200
rect 4180 200 4200 260
rect 4300 200 4450 300
rect 4550 200 4700 300
rect 4800 260 5200 300
rect 4800 200 4820 260
rect 4180 180 4820 200
rect 5180 200 5200 260
rect 5300 200 5450 300
rect 5550 200 5700 300
rect 5800 260 6200 300
rect 5800 200 5820 260
rect 5180 180 5820 200
rect 6180 200 6200 260
rect 6300 200 6450 300
rect 6550 200 6700 300
rect 6800 260 7200 300
rect 6800 200 6820 260
rect 6180 180 6820 200
rect 7180 200 7200 260
rect 7300 200 7450 300
rect 7550 200 7700 300
rect 7800 260 8000 300
rect 7800 200 7820 260
rect 7180 180 7820 200
rect 260 0 740 180
rect 1260 0 1740 180
rect 2260 0 2740 180
rect 3260 0 3740 180
rect 4260 0 4740 180
rect 5260 0 5740 180
rect 6260 0 6740 180
rect 7260 0 7740 180
<< end >>
