magic
tech sky130B
magscale 1 2
timestamp 1661911784
<< pwell >>
rect -6860 16066 -5174 17128
rect -2100 7400 -1486 8886
rect -194 8517 1020 8520
rect -194 8512 1069 8517
rect -194 8490 1166 8512
rect -200 7419 1176 8490
rect -200 7370 1138 7419
rect 1151 7370 1176 7419
rect -200 7344 1176 7370
rect -200 7330 -124 7344
rect -114 7330 1176 7344
rect -194 7320 1166 7330
rect -1300 5640 -686 7126
rect -4400 -2100 -3678 -590
rect 0 -740 1030 460
<< nmos >>
rect -6666 16092 -6636 17102
rect -6580 16092 -6550 17102
rect -6272 16092 -6242 17102
rect -6186 16092 -6156 17102
rect -5878 16092 -5848 17102
rect -5792 16092 -5762 17102
rect -5484 16092 -5454 17102
rect -5398 16092 -5368 17102
rect -1 7481 29 8491
rect 85 7481 115 8491
rect 171 7481 201 8491
rect 257 7481 287 8491
rect 343 7481 373 8491
rect 429 7481 459 8491
rect 515 7481 545 8491
rect 601 7481 631 8491
rect 687 7481 717 8491
rect 773 7481 803 8491
rect 859 7481 889 8491
rect 945 7481 975 8491
rect 203 -711 233 299
rect 289 -711 319 299
rect 375 -711 405 299
rect 461 -711 491 299
rect 547 -711 577 299
rect 633 -711 663 299
rect 719 -711 749 299
rect 805 -711 835 299
<< ndiff >>
rect -6722 17090 -6666 17102
rect -6722 17056 -6711 17090
rect -6677 17056 -6666 17090
rect -6722 17022 -6666 17056
rect -6722 16988 -6711 17022
rect -6677 16988 -6666 17022
rect -6722 16954 -6666 16988
rect -6722 16920 -6711 16954
rect -6677 16920 -6666 16954
rect -6722 16886 -6666 16920
rect -6722 16852 -6711 16886
rect -6677 16852 -6666 16886
rect -6722 16818 -6666 16852
rect -6722 16784 -6711 16818
rect -6677 16784 -6666 16818
rect -6722 16750 -6666 16784
rect -6722 16716 -6711 16750
rect -6677 16716 -6666 16750
rect -6722 16682 -6666 16716
rect -6722 16648 -6711 16682
rect -6677 16648 -6666 16682
rect -6722 16614 -6666 16648
rect -6722 16580 -6711 16614
rect -6677 16580 -6666 16614
rect -6722 16546 -6666 16580
rect -6722 16512 -6711 16546
rect -6677 16512 -6666 16546
rect -6722 16478 -6666 16512
rect -6722 16444 -6711 16478
rect -6677 16444 -6666 16478
rect -6722 16410 -6666 16444
rect -6722 16376 -6711 16410
rect -6677 16376 -6666 16410
rect -6722 16342 -6666 16376
rect -6722 16308 -6711 16342
rect -6677 16308 -6666 16342
rect -6722 16274 -6666 16308
rect -6722 16240 -6711 16274
rect -6677 16240 -6666 16274
rect -6722 16206 -6666 16240
rect -6722 16172 -6711 16206
rect -6677 16172 -6666 16206
rect -6722 16138 -6666 16172
rect -6722 16104 -6711 16138
rect -6677 16104 -6666 16138
rect -6722 16092 -6666 16104
rect -6636 17090 -6580 17102
rect -6636 17056 -6625 17090
rect -6591 17056 -6580 17090
rect -6636 17022 -6580 17056
rect -6636 16988 -6625 17022
rect -6591 16988 -6580 17022
rect -6636 16954 -6580 16988
rect -6636 16920 -6625 16954
rect -6591 16920 -6580 16954
rect -6636 16886 -6580 16920
rect -6636 16852 -6625 16886
rect -6591 16852 -6580 16886
rect -6636 16818 -6580 16852
rect -6636 16784 -6625 16818
rect -6591 16784 -6580 16818
rect -6636 16750 -6580 16784
rect -6636 16716 -6625 16750
rect -6591 16716 -6580 16750
rect -6636 16682 -6580 16716
rect -6636 16648 -6625 16682
rect -6591 16648 -6580 16682
rect -6636 16614 -6580 16648
rect -6636 16580 -6625 16614
rect -6591 16580 -6580 16614
rect -6636 16546 -6580 16580
rect -6636 16512 -6625 16546
rect -6591 16512 -6580 16546
rect -6636 16478 -6580 16512
rect -6636 16444 -6625 16478
rect -6591 16444 -6580 16478
rect -6636 16410 -6580 16444
rect -6636 16376 -6625 16410
rect -6591 16376 -6580 16410
rect -6636 16342 -6580 16376
rect -6636 16308 -6625 16342
rect -6591 16308 -6580 16342
rect -6636 16274 -6580 16308
rect -6636 16240 -6625 16274
rect -6591 16240 -6580 16274
rect -6636 16206 -6580 16240
rect -6636 16172 -6625 16206
rect -6591 16172 -6580 16206
rect -6636 16138 -6580 16172
rect -6636 16104 -6625 16138
rect -6591 16104 -6580 16138
rect -6636 16092 -6580 16104
rect -6550 17090 -6494 17102
rect -6550 17056 -6539 17090
rect -6505 17056 -6494 17090
rect -6550 17022 -6494 17056
rect -6550 16988 -6539 17022
rect -6505 16988 -6494 17022
rect -6550 16954 -6494 16988
rect -6550 16920 -6539 16954
rect -6505 16920 -6494 16954
rect -6550 16886 -6494 16920
rect -6550 16852 -6539 16886
rect -6505 16852 -6494 16886
rect -6550 16818 -6494 16852
rect -6550 16784 -6539 16818
rect -6505 16784 -6494 16818
rect -6550 16750 -6494 16784
rect -6550 16716 -6539 16750
rect -6505 16716 -6494 16750
rect -6550 16682 -6494 16716
rect -6550 16648 -6539 16682
rect -6505 16648 -6494 16682
rect -6550 16614 -6494 16648
rect -6550 16580 -6539 16614
rect -6505 16580 -6494 16614
rect -6550 16546 -6494 16580
rect -6550 16512 -6539 16546
rect -6505 16512 -6494 16546
rect -6550 16478 -6494 16512
rect -6550 16444 -6539 16478
rect -6505 16444 -6494 16478
rect -6550 16410 -6494 16444
rect -6550 16376 -6539 16410
rect -6505 16376 -6494 16410
rect -6550 16342 -6494 16376
rect -6550 16308 -6539 16342
rect -6505 16308 -6494 16342
rect -6550 16274 -6494 16308
rect -6550 16240 -6539 16274
rect -6505 16240 -6494 16274
rect -6550 16206 -6494 16240
rect -6550 16172 -6539 16206
rect -6505 16172 -6494 16206
rect -6550 16138 -6494 16172
rect -6550 16104 -6539 16138
rect -6505 16104 -6494 16138
rect -6550 16092 -6494 16104
rect -6328 17090 -6272 17102
rect -6328 17056 -6317 17090
rect -6283 17056 -6272 17090
rect -6328 17022 -6272 17056
rect -6328 16988 -6317 17022
rect -6283 16988 -6272 17022
rect -6328 16954 -6272 16988
rect -6328 16920 -6317 16954
rect -6283 16920 -6272 16954
rect -6328 16886 -6272 16920
rect -6328 16852 -6317 16886
rect -6283 16852 -6272 16886
rect -6328 16818 -6272 16852
rect -6328 16784 -6317 16818
rect -6283 16784 -6272 16818
rect -6328 16750 -6272 16784
rect -6328 16716 -6317 16750
rect -6283 16716 -6272 16750
rect -6328 16682 -6272 16716
rect -6328 16648 -6317 16682
rect -6283 16648 -6272 16682
rect -6328 16614 -6272 16648
rect -6328 16580 -6317 16614
rect -6283 16580 -6272 16614
rect -6328 16546 -6272 16580
rect -6328 16512 -6317 16546
rect -6283 16512 -6272 16546
rect -6328 16478 -6272 16512
rect -6328 16444 -6317 16478
rect -6283 16444 -6272 16478
rect -6328 16410 -6272 16444
rect -6328 16376 -6317 16410
rect -6283 16376 -6272 16410
rect -6328 16342 -6272 16376
rect -6328 16308 -6317 16342
rect -6283 16308 -6272 16342
rect -6328 16274 -6272 16308
rect -6328 16240 -6317 16274
rect -6283 16240 -6272 16274
rect -6328 16206 -6272 16240
rect -6328 16172 -6317 16206
rect -6283 16172 -6272 16206
rect -6328 16138 -6272 16172
rect -6328 16104 -6317 16138
rect -6283 16104 -6272 16138
rect -6328 16092 -6272 16104
rect -6242 17090 -6186 17102
rect -6242 17056 -6231 17090
rect -6197 17056 -6186 17090
rect -6242 17022 -6186 17056
rect -6242 16988 -6231 17022
rect -6197 16988 -6186 17022
rect -6242 16954 -6186 16988
rect -6242 16920 -6231 16954
rect -6197 16920 -6186 16954
rect -6242 16886 -6186 16920
rect -6242 16852 -6231 16886
rect -6197 16852 -6186 16886
rect -6242 16818 -6186 16852
rect -6242 16784 -6231 16818
rect -6197 16784 -6186 16818
rect -6242 16750 -6186 16784
rect -6242 16716 -6231 16750
rect -6197 16716 -6186 16750
rect -6242 16682 -6186 16716
rect -6242 16648 -6231 16682
rect -6197 16648 -6186 16682
rect -6242 16614 -6186 16648
rect -6242 16580 -6231 16614
rect -6197 16580 -6186 16614
rect -6242 16546 -6186 16580
rect -6242 16512 -6231 16546
rect -6197 16512 -6186 16546
rect -6242 16478 -6186 16512
rect -6242 16444 -6231 16478
rect -6197 16444 -6186 16478
rect -6242 16410 -6186 16444
rect -6242 16376 -6231 16410
rect -6197 16376 -6186 16410
rect -6242 16342 -6186 16376
rect -6242 16308 -6231 16342
rect -6197 16308 -6186 16342
rect -6242 16274 -6186 16308
rect -6242 16240 -6231 16274
rect -6197 16240 -6186 16274
rect -6242 16206 -6186 16240
rect -6242 16172 -6231 16206
rect -6197 16172 -6186 16206
rect -6242 16138 -6186 16172
rect -6242 16104 -6231 16138
rect -6197 16104 -6186 16138
rect -6242 16092 -6186 16104
rect -6156 17090 -6100 17102
rect -6156 17056 -6145 17090
rect -6111 17056 -6100 17090
rect -6156 17022 -6100 17056
rect -6156 16988 -6145 17022
rect -6111 16988 -6100 17022
rect -6156 16954 -6100 16988
rect -6156 16920 -6145 16954
rect -6111 16920 -6100 16954
rect -6156 16886 -6100 16920
rect -6156 16852 -6145 16886
rect -6111 16852 -6100 16886
rect -6156 16818 -6100 16852
rect -6156 16784 -6145 16818
rect -6111 16784 -6100 16818
rect -6156 16750 -6100 16784
rect -6156 16716 -6145 16750
rect -6111 16716 -6100 16750
rect -6156 16682 -6100 16716
rect -6156 16648 -6145 16682
rect -6111 16648 -6100 16682
rect -6156 16614 -6100 16648
rect -6156 16580 -6145 16614
rect -6111 16580 -6100 16614
rect -6156 16546 -6100 16580
rect -6156 16512 -6145 16546
rect -6111 16512 -6100 16546
rect -6156 16478 -6100 16512
rect -6156 16444 -6145 16478
rect -6111 16444 -6100 16478
rect -6156 16410 -6100 16444
rect -6156 16376 -6145 16410
rect -6111 16376 -6100 16410
rect -6156 16342 -6100 16376
rect -6156 16308 -6145 16342
rect -6111 16308 -6100 16342
rect -6156 16274 -6100 16308
rect -6156 16240 -6145 16274
rect -6111 16240 -6100 16274
rect -6156 16206 -6100 16240
rect -6156 16172 -6145 16206
rect -6111 16172 -6100 16206
rect -6156 16138 -6100 16172
rect -6156 16104 -6145 16138
rect -6111 16104 -6100 16138
rect -6156 16092 -6100 16104
rect -5934 17090 -5878 17102
rect -5934 17056 -5923 17090
rect -5889 17056 -5878 17090
rect -5934 17022 -5878 17056
rect -5934 16988 -5923 17022
rect -5889 16988 -5878 17022
rect -5934 16954 -5878 16988
rect -5934 16920 -5923 16954
rect -5889 16920 -5878 16954
rect -5934 16886 -5878 16920
rect -5934 16852 -5923 16886
rect -5889 16852 -5878 16886
rect -5934 16818 -5878 16852
rect -5934 16784 -5923 16818
rect -5889 16784 -5878 16818
rect -5934 16750 -5878 16784
rect -5934 16716 -5923 16750
rect -5889 16716 -5878 16750
rect -5934 16682 -5878 16716
rect -5934 16648 -5923 16682
rect -5889 16648 -5878 16682
rect -5934 16614 -5878 16648
rect -5934 16580 -5923 16614
rect -5889 16580 -5878 16614
rect -5934 16546 -5878 16580
rect -5934 16512 -5923 16546
rect -5889 16512 -5878 16546
rect -5934 16478 -5878 16512
rect -5934 16444 -5923 16478
rect -5889 16444 -5878 16478
rect -5934 16410 -5878 16444
rect -5934 16376 -5923 16410
rect -5889 16376 -5878 16410
rect -5934 16342 -5878 16376
rect -5934 16308 -5923 16342
rect -5889 16308 -5878 16342
rect -5934 16274 -5878 16308
rect -5934 16240 -5923 16274
rect -5889 16240 -5878 16274
rect -5934 16206 -5878 16240
rect -5934 16172 -5923 16206
rect -5889 16172 -5878 16206
rect -5934 16138 -5878 16172
rect -5934 16104 -5923 16138
rect -5889 16104 -5878 16138
rect -5934 16092 -5878 16104
rect -5848 17090 -5792 17102
rect -5848 17056 -5837 17090
rect -5803 17056 -5792 17090
rect -5848 17022 -5792 17056
rect -5848 16988 -5837 17022
rect -5803 16988 -5792 17022
rect -5848 16954 -5792 16988
rect -5848 16920 -5837 16954
rect -5803 16920 -5792 16954
rect -5848 16886 -5792 16920
rect -5848 16852 -5837 16886
rect -5803 16852 -5792 16886
rect -5848 16818 -5792 16852
rect -5848 16784 -5837 16818
rect -5803 16784 -5792 16818
rect -5848 16750 -5792 16784
rect -5848 16716 -5837 16750
rect -5803 16716 -5792 16750
rect -5848 16682 -5792 16716
rect -5848 16648 -5837 16682
rect -5803 16648 -5792 16682
rect -5848 16614 -5792 16648
rect -5848 16580 -5837 16614
rect -5803 16580 -5792 16614
rect -5848 16546 -5792 16580
rect -5848 16512 -5837 16546
rect -5803 16512 -5792 16546
rect -5848 16478 -5792 16512
rect -5848 16444 -5837 16478
rect -5803 16444 -5792 16478
rect -5848 16410 -5792 16444
rect -5848 16376 -5837 16410
rect -5803 16376 -5792 16410
rect -5848 16342 -5792 16376
rect -5848 16308 -5837 16342
rect -5803 16308 -5792 16342
rect -5848 16274 -5792 16308
rect -5848 16240 -5837 16274
rect -5803 16240 -5792 16274
rect -5848 16206 -5792 16240
rect -5848 16172 -5837 16206
rect -5803 16172 -5792 16206
rect -5848 16138 -5792 16172
rect -5848 16104 -5837 16138
rect -5803 16104 -5792 16138
rect -5848 16092 -5792 16104
rect -5762 17090 -5706 17102
rect -5762 17056 -5751 17090
rect -5717 17056 -5706 17090
rect -5762 17022 -5706 17056
rect -5762 16988 -5751 17022
rect -5717 16988 -5706 17022
rect -5762 16954 -5706 16988
rect -5762 16920 -5751 16954
rect -5717 16920 -5706 16954
rect -5762 16886 -5706 16920
rect -5762 16852 -5751 16886
rect -5717 16852 -5706 16886
rect -5762 16818 -5706 16852
rect -5762 16784 -5751 16818
rect -5717 16784 -5706 16818
rect -5762 16750 -5706 16784
rect -5762 16716 -5751 16750
rect -5717 16716 -5706 16750
rect -5762 16682 -5706 16716
rect -5762 16648 -5751 16682
rect -5717 16648 -5706 16682
rect -5762 16614 -5706 16648
rect -5762 16580 -5751 16614
rect -5717 16580 -5706 16614
rect -5762 16546 -5706 16580
rect -5762 16512 -5751 16546
rect -5717 16512 -5706 16546
rect -5762 16478 -5706 16512
rect -5762 16444 -5751 16478
rect -5717 16444 -5706 16478
rect -5762 16410 -5706 16444
rect -5762 16376 -5751 16410
rect -5717 16376 -5706 16410
rect -5762 16342 -5706 16376
rect -5762 16308 -5751 16342
rect -5717 16308 -5706 16342
rect -5762 16274 -5706 16308
rect -5762 16240 -5751 16274
rect -5717 16240 -5706 16274
rect -5762 16206 -5706 16240
rect -5762 16172 -5751 16206
rect -5717 16172 -5706 16206
rect -5762 16138 -5706 16172
rect -5762 16104 -5751 16138
rect -5717 16104 -5706 16138
rect -5762 16092 -5706 16104
rect -5540 17090 -5484 17102
rect -5540 17056 -5529 17090
rect -5495 17056 -5484 17090
rect -5540 17022 -5484 17056
rect -5540 16988 -5529 17022
rect -5495 16988 -5484 17022
rect -5540 16954 -5484 16988
rect -5540 16920 -5529 16954
rect -5495 16920 -5484 16954
rect -5540 16886 -5484 16920
rect -5540 16852 -5529 16886
rect -5495 16852 -5484 16886
rect -5540 16818 -5484 16852
rect -5540 16784 -5529 16818
rect -5495 16784 -5484 16818
rect -5540 16750 -5484 16784
rect -5540 16716 -5529 16750
rect -5495 16716 -5484 16750
rect -5540 16682 -5484 16716
rect -5540 16648 -5529 16682
rect -5495 16648 -5484 16682
rect -5540 16614 -5484 16648
rect -5540 16580 -5529 16614
rect -5495 16580 -5484 16614
rect -5540 16546 -5484 16580
rect -5540 16512 -5529 16546
rect -5495 16512 -5484 16546
rect -5540 16478 -5484 16512
rect -5540 16444 -5529 16478
rect -5495 16444 -5484 16478
rect -5540 16410 -5484 16444
rect -5540 16376 -5529 16410
rect -5495 16376 -5484 16410
rect -5540 16342 -5484 16376
rect -5540 16308 -5529 16342
rect -5495 16308 -5484 16342
rect -5540 16274 -5484 16308
rect -5540 16240 -5529 16274
rect -5495 16240 -5484 16274
rect -5540 16206 -5484 16240
rect -5540 16172 -5529 16206
rect -5495 16172 -5484 16206
rect -5540 16138 -5484 16172
rect -5540 16104 -5529 16138
rect -5495 16104 -5484 16138
rect -5540 16092 -5484 16104
rect -5454 17090 -5398 17102
rect -5454 17056 -5443 17090
rect -5409 17056 -5398 17090
rect -5454 17022 -5398 17056
rect -5454 16988 -5443 17022
rect -5409 16988 -5398 17022
rect -5454 16954 -5398 16988
rect -5454 16920 -5443 16954
rect -5409 16920 -5398 16954
rect -5454 16886 -5398 16920
rect -5454 16852 -5443 16886
rect -5409 16852 -5398 16886
rect -5454 16818 -5398 16852
rect -5454 16784 -5443 16818
rect -5409 16784 -5398 16818
rect -5454 16750 -5398 16784
rect -5454 16716 -5443 16750
rect -5409 16716 -5398 16750
rect -5454 16682 -5398 16716
rect -5454 16648 -5443 16682
rect -5409 16648 -5398 16682
rect -5454 16614 -5398 16648
rect -5454 16580 -5443 16614
rect -5409 16580 -5398 16614
rect -5454 16546 -5398 16580
rect -5454 16512 -5443 16546
rect -5409 16512 -5398 16546
rect -5454 16478 -5398 16512
rect -5454 16444 -5443 16478
rect -5409 16444 -5398 16478
rect -5454 16410 -5398 16444
rect -5454 16376 -5443 16410
rect -5409 16376 -5398 16410
rect -5454 16342 -5398 16376
rect -5454 16308 -5443 16342
rect -5409 16308 -5398 16342
rect -5454 16274 -5398 16308
rect -5454 16240 -5443 16274
rect -5409 16240 -5398 16274
rect -5454 16206 -5398 16240
rect -5454 16172 -5443 16206
rect -5409 16172 -5398 16206
rect -5454 16138 -5398 16172
rect -5454 16104 -5443 16138
rect -5409 16104 -5398 16138
rect -5454 16092 -5398 16104
rect -5368 17090 -5312 17102
rect -5368 17056 -5357 17090
rect -5323 17056 -5312 17090
rect -5368 17022 -5312 17056
rect -5368 16988 -5357 17022
rect -5323 16988 -5312 17022
rect -5368 16954 -5312 16988
rect -5368 16920 -5357 16954
rect -5323 16920 -5312 16954
rect -5368 16886 -5312 16920
rect -5368 16852 -5357 16886
rect -5323 16852 -5312 16886
rect -5368 16818 -5312 16852
rect -5368 16784 -5357 16818
rect -5323 16784 -5312 16818
rect -5368 16750 -5312 16784
rect -5368 16716 -5357 16750
rect -5323 16716 -5312 16750
rect -5368 16682 -5312 16716
rect -5368 16648 -5357 16682
rect -5323 16648 -5312 16682
rect -5368 16614 -5312 16648
rect -5368 16580 -5357 16614
rect -5323 16580 -5312 16614
rect -5368 16546 -5312 16580
rect -5368 16512 -5357 16546
rect -5323 16512 -5312 16546
rect -5368 16478 -5312 16512
rect -5368 16444 -5357 16478
rect -5323 16444 -5312 16478
rect -5368 16410 -5312 16444
rect -5368 16376 -5357 16410
rect -5323 16376 -5312 16410
rect -5368 16342 -5312 16376
rect -5368 16308 -5357 16342
rect -5323 16308 -5312 16342
rect -5368 16274 -5312 16308
rect -5368 16240 -5357 16274
rect -5323 16240 -5312 16274
rect -5368 16206 -5312 16240
rect -5368 16172 -5357 16206
rect -5323 16172 -5312 16206
rect -5368 16138 -5312 16172
rect -5368 16104 -5357 16138
rect -5323 16104 -5312 16138
rect -5368 16092 -5312 16104
rect -57 8479 -1 8491
rect -57 8445 -46 8479
rect -12 8445 -1 8479
rect -57 8411 -1 8445
rect -57 8377 -46 8411
rect -12 8377 -1 8411
rect -57 8343 -1 8377
rect -57 8309 -46 8343
rect -12 8309 -1 8343
rect -57 8275 -1 8309
rect -57 8241 -46 8275
rect -12 8241 -1 8275
rect -57 8207 -1 8241
rect -57 8173 -46 8207
rect -12 8173 -1 8207
rect -57 8139 -1 8173
rect -57 8105 -46 8139
rect -12 8105 -1 8139
rect -57 8071 -1 8105
rect -57 8037 -46 8071
rect -12 8037 -1 8071
rect -57 8003 -1 8037
rect -57 7969 -46 8003
rect -12 7969 -1 8003
rect -57 7935 -1 7969
rect -57 7901 -46 7935
rect -12 7901 -1 7935
rect -57 7867 -1 7901
rect -57 7833 -46 7867
rect -12 7833 -1 7867
rect -57 7799 -1 7833
rect -57 7765 -46 7799
rect -12 7765 -1 7799
rect -57 7731 -1 7765
rect -57 7697 -46 7731
rect -12 7697 -1 7731
rect -57 7663 -1 7697
rect -57 7629 -46 7663
rect -12 7629 -1 7663
rect -57 7595 -1 7629
rect -57 7561 -46 7595
rect -12 7561 -1 7595
rect -57 7527 -1 7561
rect -57 7493 -46 7527
rect -12 7493 -1 7527
rect -57 7481 -1 7493
rect 29 8479 85 8491
rect 29 8445 40 8479
rect 74 8445 85 8479
rect 29 8411 85 8445
rect 29 8377 40 8411
rect 74 8377 85 8411
rect 29 8343 85 8377
rect 29 8309 40 8343
rect 74 8309 85 8343
rect 29 8275 85 8309
rect 29 8241 40 8275
rect 74 8241 85 8275
rect 29 8207 85 8241
rect 29 8173 40 8207
rect 74 8173 85 8207
rect 29 8139 85 8173
rect 29 8105 40 8139
rect 74 8105 85 8139
rect 29 8071 85 8105
rect 29 8037 40 8071
rect 74 8037 85 8071
rect 29 8003 85 8037
rect 29 7969 40 8003
rect 74 7969 85 8003
rect 29 7935 85 7969
rect 29 7901 40 7935
rect 74 7901 85 7935
rect 29 7867 85 7901
rect 29 7833 40 7867
rect 74 7833 85 7867
rect 29 7799 85 7833
rect 29 7765 40 7799
rect 74 7765 85 7799
rect 29 7731 85 7765
rect 29 7697 40 7731
rect 74 7697 85 7731
rect 29 7663 85 7697
rect 29 7629 40 7663
rect 74 7629 85 7663
rect 29 7595 85 7629
rect 29 7561 40 7595
rect 74 7561 85 7595
rect 29 7527 85 7561
rect 29 7493 40 7527
rect 74 7493 85 7527
rect 29 7481 85 7493
rect 115 8479 171 8491
rect 115 8445 126 8479
rect 160 8445 171 8479
rect 115 8411 171 8445
rect 115 8377 126 8411
rect 160 8377 171 8411
rect 115 8343 171 8377
rect 115 8309 126 8343
rect 160 8309 171 8343
rect 115 8275 171 8309
rect 115 8241 126 8275
rect 160 8241 171 8275
rect 115 8207 171 8241
rect 115 8173 126 8207
rect 160 8173 171 8207
rect 115 8139 171 8173
rect 115 8105 126 8139
rect 160 8105 171 8139
rect 115 8071 171 8105
rect 115 8037 126 8071
rect 160 8037 171 8071
rect 115 8003 171 8037
rect 115 7969 126 8003
rect 160 7969 171 8003
rect 115 7935 171 7969
rect 115 7901 126 7935
rect 160 7901 171 7935
rect 115 7867 171 7901
rect 115 7833 126 7867
rect 160 7833 171 7867
rect 115 7799 171 7833
rect 115 7765 126 7799
rect 160 7765 171 7799
rect 115 7731 171 7765
rect 115 7697 126 7731
rect 160 7697 171 7731
rect 115 7663 171 7697
rect 115 7629 126 7663
rect 160 7629 171 7663
rect 115 7595 171 7629
rect 115 7561 126 7595
rect 160 7561 171 7595
rect 115 7527 171 7561
rect 115 7493 126 7527
rect 160 7493 171 7527
rect 115 7481 171 7493
rect 201 8479 257 8491
rect 201 8445 212 8479
rect 246 8445 257 8479
rect 201 8411 257 8445
rect 201 8377 212 8411
rect 246 8377 257 8411
rect 201 8343 257 8377
rect 201 8309 212 8343
rect 246 8309 257 8343
rect 201 8275 257 8309
rect 201 8241 212 8275
rect 246 8241 257 8275
rect 201 8207 257 8241
rect 201 8173 212 8207
rect 246 8173 257 8207
rect 201 8139 257 8173
rect 201 8105 212 8139
rect 246 8105 257 8139
rect 201 8071 257 8105
rect 201 8037 212 8071
rect 246 8037 257 8071
rect 201 8003 257 8037
rect 201 7969 212 8003
rect 246 7969 257 8003
rect 201 7935 257 7969
rect 201 7901 212 7935
rect 246 7901 257 7935
rect 201 7867 257 7901
rect 201 7833 212 7867
rect 246 7833 257 7867
rect 201 7799 257 7833
rect 201 7765 212 7799
rect 246 7765 257 7799
rect 201 7731 257 7765
rect 201 7697 212 7731
rect 246 7697 257 7731
rect 201 7663 257 7697
rect 201 7629 212 7663
rect 246 7629 257 7663
rect 201 7595 257 7629
rect 201 7561 212 7595
rect 246 7561 257 7595
rect 201 7527 257 7561
rect 201 7493 212 7527
rect 246 7493 257 7527
rect 201 7481 257 7493
rect 287 8479 343 8491
rect 287 8445 298 8479
rect 332 8445 343 8479
rect 287 8411 343 8445
rect 287 8377 298 8411
rect 332 8377 343 8411
rect 287 8343 343 8377
rect 287 8309 298 8343
rect 332 8309 343 8343
rect 287 8275 343 8309
rect 287 8241 298 8275
rect 332 8241 343 8275
rect 287 8207 343 8241
rect 287 8173 298 8207
rect 332 8173 343 8207
rect 287 8139 343 8173
rect 287 8105 298 8139
rect 332 8105 343 8139
rect 287 8071 343 8105
rect 287 8037 298 8071
rect 332 8037 343 8071
rect 287 8003 343 8037
rect 287 7969 298 8003
rect 332 7969 343 8003
rect 287 7935 343 7969
rect 287 7901 298 7935
rect 332 7901 343 7935
rect 287 7867 343 7901
rect 287 7833 298 7867
rect 332 7833 343 7867
rect 287 7799 343 7833
rect 287 7765 298 7799
rect 332 7765 343 7799
rect 287 7731 343 7765
rect 287 7697 298 7731
rect 332 7697 343 7731
rect 287 7663 343 7697
rect 287 7629 298 7663
rect 332 7629 343 7663
rect 287 7595 343 7629
rect 287 7561 298 7595
rect 332 7561 343 7595
rect 287 7527 343 7561
rect 287 7493 298 7527
rect 332 7493 343 7527
rect 287 7481 343 7493
rect 373 8479 429 8491
rect 373 8445 384 8479
rect 418 8445 429 8479
rect 373 8411 429 8445
rect 373 8377 384 8411
rect 418 8377 429 8411
rect 373 8343 429 8377
rect 373 8309 384 8343
rect 418 8309 429 8343
rect 373 8275 429 8309
rect 373 8241 384 8275
rect 418 8241 429 8275
rect 373 8207 429 8241
rect 373 8173 384 8207
rect 418 8173 429 8207
rect 373 8139 429 8173
rect 373 8105 384 8139
rect 418 8105 429 8139
rect 373 8071 429 8105
rect 373 8037 384 8071
rect 418 8037 429 8071
rect 373 8003 429 8037
rect 373 7969 384 8003
rect 418 7969 429 8003
rect 373 7935 429 7969
rect 373 7901 384 7935
rect 418 7901 429 7935
rect 373 7867 429 7901
rect 373 7833 384 7867
rect 418 7833 429 7867
rect 373 7799 429 7833
rect 373 7765 384 7799
rect 418 7765 429 7799
rect 373 7731 429 7765
rect 373 7697 384 7731
rect 418 7697 429 7731
rect 373 7663 429 7697
rect 373 7629 384 7663
rect 418 7629 429 7663
rect 373 7595 429 7629
rect 373 7561 384 7595
rect 418 7561 429 7595
rect 373 7527 429 7561
rect 373 7493 384 7527
rect 418 7493 429 7527
rect 373 7481 429 7493
rect 459 8479 515 8491
rect 459 8445 470 8479
rect 504 8445 515 8479
rect 459 8411 515 8445
rect 459 8377 470 8411
rect 504 8377 515 8411
rect 459 8343 515 8377
rect 459 8309 470 8343
rect 504 8309 515 8343
rect 459 8275 515 8309
rect 459 8241 470 8275
rect 504 8241 515 8275
rect 459 8207 515 8241
rect 459 8173 470 8207
rect 504 8173 515 8207
rect 459 8139 515 8173
rect 459 8105 470 8139
rect 504 8105 515 8139
rect 459 8071 515 8105
rect 459 8037 470 8071
rect 504 8037 515 8071
rect 459 8003 515 8037
rect 459 7969 470 8003
rect 504 7969 515 8003
rect 459 7935 515 7969
rect 459 7901 470 7935
rect 504 7901 515 7935
rect 459 7867 515 7901
rect 459 7833 470 7867
rect 504 7833 515 7867
rect 459 7799 515 7833
rect 459 7765 470 7799
rect 504 7765 515 7799
rect 459 7731 515 7765
rect 459 7697 470 7731
rect 504 7697 515 7731
rect 459 7663 515 7697
rect 459 7629 470 7663
rect 504 7629 515 7663
rect 459 7595 515 7629
rect 459 7561 470 7595
rect 504 7561 515 7595
rect 459 7527 515 7561
rect 459 7493 470 7527
rect 504 7493 515 7527
rect 459 7481 515 7493
rect 545 8479 601 8491
rect 545 8445 556 8479
rect 590 8445 601 8479
rect 545 8411 601 8445
rect 545 8377 556 8411
rect 590 8377 601 8411
rect 545 8343 601 8377
rect 545 8309 556 8343
rect 590 8309 601 8343
rect 545 8275 601 8309
rect 545 8241 556 8275
rect 590 8241 601 8275
rect 545 8207 601 8241
rect 545 8173 556 8207
rect 590 8173 601 8207
rect 545 8139 601 8173
rect 545 8105 556 8139
rect 590 8105 601 8139
rect 545 8071 601 8105
rect 545 8037 556 8071
rect 590 8037 601 8071
rect 545 8003 601 8037
rect 545 7969 556 8003
rect 590 7969 601 8003
rect 545 7935 601 7969
rect 545 7901 556 7935
rect 590 7901 601 7935
rect 545 7867 601 7901
rect 545 7833 556 7867
rect 590 7833 601 7867
rect 545 7799 601 7833
rect 545 7765 556 7799
rect 590 7765 601 7799
rect 545 7731 601 7765
rect 545 7697 556 7731
rect 590 7697 601 7731
rect 545 7663 601 7697
rect 545 7629 556 7663
rect 590 7629 601 7663
rect 545 7595 601 7629
rect 545 7561 556 7595
rect 590 7561 601 7595
rect 545 7527 601 7561
rect 545 7493 556 7527
rect 590 7493 601 7527
rect 545 7481 601 7493
rect 631 8479 687 8491
rect 631 8445 642 8479
rect 676 8445 687 8479
rect 631 8411 687 8445
rect 631 8377 642 8411
rect 676 8377 687 8411
rect 631 8343 687 8377
rect 631 8309 642 8343
rect 676 8309 687 8343
rect 631 8275 687 8309
rect 631 8241 642 8275
rect 676 8241 687 8275
rect 631 8207 687 8241
rect 631 8173 642 8207
rect 676 8173 687 8207
rect 631 8139 687 8173
rect 631 8105 642 8139
rect 676 8105 687 8139
rect 631 8071 687 8105
rect 631 8037 642 8071
rect 676 8037 687 8071
rect 631 8003 687 8037
rect 631 7969 642 8003
rect 676 7969 687 8003
rect 631 7935 687 7969
rect 631 7901 642 7935
rect 676 7901 687 7935
rect 631 7867 687 7901
rect 631 7833 642 7867
rect 676 7833 687 7867
rect 631 7799 687 7833
rect 631 7765 642 7799
rect 676 7765 687 7799
rect 631 7731 687 7765
rect 631 7697 642 7731
rect 676 7697 687 7731
rect 631 7663 687 7697
rect 631 7629 642 7663
rect 676 7629 687 7663
rect 631 7595 687 7629
rect 631 7561 642 7595
rect 676 7561 687 7595
rect 631 7527 687 7561
rect 631 7493 642 7527
rect 676 7493 687 7527
rect 631 7481 687 7493
rect 717 8479 773 8491
rect 717 8445 728 8479
rect 762 8445 773 8479
rect 717 8411 773 8445
rect 717 8377 728 8411
rect 762 8377 773 8411
rect 717 8343 773 8377
rect 717 8309 728 8343
rect 762 8309 773 8343
rect 717 8275 773 8309
rect 717 8241 728 8275
rect 762 8241 773 8275
rect 717 8207 773 8241
rect 717 8173 728 8207
rect 762 8173 773 8207
rect 717 8139 773 8173
rect 717 8105 728 8139
rect 762 8105 773 8139
rect 717 8071 773 8105
rect 717 8037 728 8071
rect 762 8037 773 8071
rect 717 8003 773 8037
rect 717 7969 728 8003
rect 762 7969 773 8003
rect 717 7935 773 7969
rect 717 7901 728 7935
rect 762 7901 773 7935
rect 717 7867 773 7901
rect 717 7833 728 7867
rect 762 7833 773 7867
rect 717 7799 773 7833
rect 717 7765 728 7799
rect 762 7765 773 7799
rect 717 7731 773 7765
rect 717 7697 728 7731
rect 762 7697 773 7731
rect 717 7663 773 7697
rect 717 7629 728 7663
rect 762 7629 773 7663
rect 717 7595 773 7629
rect 717 7561 728 7595
rect 762 7561 773 7595
rect 717 7527 773 7561
rect 717 7493 728 7527
rect 762 7493 773 7527
rect 717 7481 773 7493
rect 803 8479 859 8491
rect 803 8445 814 8479
rect 848 8445 859 8479
rect 803 8411 859 8445
rect 803 8377 814 8411
rect 848 8377 859 8411
rect 803 8343 859 8377
rect 803 8309 814 8343
rect 848 8309 859 8343
rect 803 8275 859 8309
rect 803 8241 814 8275
rect 848 8241 859 8275
rect 803 8207 859 8241
rect 803 8173 814 8207
rect 848 8173 859 8207
rect 803 8139 859 8173
rect 803 8105 814 8139
rect 848 8105 859 8139
rect 803 8071 859 8105
rect 803 8037 814 8071
rect 848 8037 859 8071
rect 803 8003 859 8037
rect 803 7969 814 8003
rect 848 7969 859 8003
rect 803 7935 859 7969
rect 803 7901 814 7935
rect 848 7901 859 7935
rect 803 7867 859 7901
rect 803 7833 814 7867
rect 848 7833 859 7867
rect 803 7799 859 7833
rect 803 7765 814 7799
rect 848 7765 859 7799
rect 803 7731 859 7765
rect 803 7697 814 7731
rect 848 7697 859 7731
rect 803 7663 859 7697
rect 803 7629 814 7663
rect 848 7629 859 7663
rect 803 7595 859 7629
rect 803 7561 814 7595
rect 848 7561 859 7595
rect 803 7527 859 7561
rect 803 7493 814 7527
rect 848 7493 859 7527
rect 803 7481 859 7493
rect 889 8479 945 8491
rect 889 8445 900 8479
rect 934 8445 945 8479
rect 889 8411 945 8445
rect 889 8377 900 8411
rect 934 8377 945 8411
rect 889 8343 945 8377
rect 889 8309 900 8343
rect 934 8309 945 8343
rect 889 8275 945 8309
rect 889 8241 900 8275
rect 934 8241 945 8275
rect 889 8207 945 8241
rect 889 8173 900 8207
rect 934 8173 945 8207
rect 889 8139 945 8173
rect 889 8105 900 8139
rect 934 8105 945 8139
rect 889 8071 945 8105
rect 889 8037 900 8071
rect 934 8037 945 8071
rect 889 8003 945 8037
rect 889 7969 900 8003
rect 934 7969 945 8003
rect 889 7935 945 7969
rect 889 7901 900 7935
rect 934 7901 945 7935
rect 889 7867 945 7901
rect 889 7833 900 7867
rect 934 7833 945 7867
rect 889 7799 945 7833
rect 889 7765 900 7799
rect 934 7765 945 7799
rect 889 7731 945 7765
rect 889 7697 900 7731
rect 934 7697 945 7731
rect 889 7663 945 7697
rect 889 7629 900 7663
rect 934 7629 945 7663
rect 889 7595 945 7629
rect 889 7561 900 7595
rect 934 7561 945 7595
rect 889 7527 945 7561
rect 889 7493 900 7527
rect 934 7493 945 7527
rect 889 7481 945 7493
rect 975 8479 1031 8491
rect 975 8445 986 8479
rect 1020 8445 1031 8479
rect 975 8411 1031 8445
rect 975 8377 986 8411
rect 1020 8377 1031 8411
rect 975 8343 1031 8377
rect 975 8309 986 8343
rect 1020 8309 1031 8343
rect 975 8275 1031 8309
rect 975 8241 986 8275
rect 1020 8241 1031 8275
rect 975 8207 1031 8241
rect 975 8173 986 8207
rect 1020 8173 1031 8207
rect 975 8139 1031 8173
rect 975 8105 986 8139
rect 1020 8105 1031 8139
rect 975 8071 1031 8105
rect 975 8037 986 8071
rect 1020 8037 1031 8071
rect 975 8003 1031 8037
rect 975 7969 986 8003
rect 1020 7969 1031 8003
rect 975 7935 1031 7969
rect 975 7901 986 7935
rect 1020 7901 1031 7935
rect 975 7867 1031 7901
rect 975 7833 986 7867
rect 1020 7833 1031 7867
rect 975 7799 1031 7833
rect 975 7765 986 7799
rect 1020 7765 1031 7799
rect 975 7731 1031 7765
rect 975 7697 986 7731
rect 1020 7697 1031 7731
rect 975 7663 1031 7697
rect 975 7629 986 7663
rect 1020 7629 1031 7663
rect 975 7595 1031 7629
rect 975 7561 986 7595
rect 1020 7561 1031 7595
rect 975 7527 1031 7561
rect 975 7493 986 7527
rect 1020 7493 1031 7527
rect 975 7481 1031 7493
rect 147 287 203 299
rect 147 253 158 287
rect 192 253 203 287
rect 147 219 203 253
rect 147 185 158 219
rect 192 185 203 219
rect 147 151 203 185
rect 147 117 158 151
rect 192 117 203 151
rect 147 83 203 117
rect 147 49 158 83
rect 192 49 203 83
rect 147 15 203 49
rect 147 -19 158 15
rect 192 -19 203 15
rect 147 -53 203 -19
rect 147 -87 158 -53
rect 192 -87 203 -53
rect 147 -121 203 -87
rect 147 -155 158 -121
rect 192 -155 203 -121
rect 147 -189 203 -155
rect 147 -223 158 -189
rect 192 -223 203 -189
rect 147 -257 203 -223
rect 147 -291 158 -257
rect 192 -291 203 -257
rect 147 -325 203 -291
rect 147 -359 158 -325
rect 192 -359 203 -325
rect 147 -393 203 -359
rect 147 -427 158 -393
rect 192 -427 203 -393
rect 147 -461 203 -427
rect 147 -495 158 -461
rect 192 -495 203 -461
rect 147 -529 203 -495
rect 147 -563 158 -529
rect 192 -563 203 -529
rect 147 -597 203 -563
rect 147 -631 158 -597
rect 192 -631 203 -597
rect 147 -665 203 -631
rect 147 -699 158 -665
rect 192 -699 203 -665
rect 147 -711 203 -699
rect 233 287 289 299
rect 233 253 244 287
rect 278 253 289 287
rect 233 219 289 253
rect 233 185 244 219
rect 278 185 289 219
rect 233 151 289 185
rect 233 117 244 151
rect 278 117 289 151
rect 233 83 289 117
rect 233 49 244 83
rect 278 49 289 83
rect 233 15 289 49
rect 233 -19 244 15
rect 278 -19 289 15
rect 233 -53 289 -19
rect 233 -87 244 -53
rect 278 -87 289 -53
rect 233 -121 289 -87
rect 233 -155 244 -121
rect 278 -155 289 -121
rect 233 -189 289 -155
rect 233 -223 244 -189
rect 278 -223 289 -189
rect 233 -257 289 -223
rect 233 -291 244 -257
rect 278 -291 289 -257
rect 233 -325 289 -291
rect 233 -359 244 -325
rect 278 -359 289 -325
rect 233 -393 289 -359
rect 233 -427 244 -393
rect 278 -427 289 -393
rect 233 -461 289 -427
rect 233 -495 244 -461
rect 278 -495 289 -461
rect 233 -529 289 -495
rect 233 -563 244 -529
rect 278 -563 289 -529
rect 233 -597 289 -563
rect 233 -631 244 -597
rect 278 -631 289 -597
rect 233 -665 289 -631
rect 233 -699 244 -665
rect 278 -699 289 -665
rect 233 -711 289 -699
rect 319 287 375 299
rect 319 253 330 287
rect 364 253 375 287
rect 319 219 375 253
rect 319 185 330 219
rect 364 185 375 219
rect 319 151 375 185
rect 319 117 330 151
rect 364 117 375 151
rect 319 83 375 117
rect 319 49 330 83
rect 364 49 375 83
rect 319 15 375 49
rect 319 -19 330 15
rect 364 -19 375 15
rect 319 -53 375 -19
rect 319 -87 330 -53
rect 364 -87 375 -53
rect 319 -121 375 -87
rect 319 -155 330 -121
rect 364 -155 375 -121
rect 319 -189 375 -155
rect 319 -223 330 -189
rect 364 -223 375 -189
rect 319 -257 375 -223
rect 319 -291 330 -257
rect 364 -291 375 -257
rect 319 -325 375 -291
rect 319 -359 330 -325
rect 364 -359 375 -325
rect 319 -393 375 -359
rect 319 -427 330 -393
rect 364 -427 375 -393
rect 319 -461 375 -427
rect 319 -495 330 -461
rect 364 -495 375 -461
rect 319 -529 375 -495
rect 319 -563 330 -529
rect 364 -563 375 -529
rect 319 -597 375 -563
rect 319 -631 330 -597
rect 364 -631 375 -597
rect 319 -665 375 -631
rect 319 -699 330 -665
rect 364 -699 375 -665
rect 319 -711 375 -699
rect 405 287 461 299
rect 405 253 416 287
rect 450 253 461 287
rect 405 219 461 253
rect 405 185 416 219
rect 450 185 461 219
rect 405 151 461 185
rect 405 117 416 151
rect 450 117 461 151
rect 405 83 461 117
rect 405 49 416 83
rect 450 49 461 83
rect 405 15 461 49
rect 405 -19 416 15
rect 450 -19 461 15
rect 405 -53 461 -19
rect 405 -87 416 -53
rect 450 -87 461 -53
rect 405 -121 461 -87
rect 405 -155 416 -121
rect 450 -155 461 -121
rect 405 -189 461 -155
rect 405 -223 416 -189
rect 450 -223 461 -189
rect 405 -257 461 -223
rect 405 -291 416 -257
rect 450 -291 461 -257
rect 405 -325 461 -291
rect 405 -359 416 -325
rect 450 -359 461 -325
rect 405 -393 461 -359
rect 405 -427 416 -393
rect 450 -427 461 -393
rect 405 -461 461 -427
rect 405 -495 416 -461
rect 450 -495 461 -461
rect 405 -529 461 -495
rect 405 -563 416 -529
rect 450 -563 461 -529
rect 405 -597 461 -563
rect 405 -631 416 -597
rect 450 -631 461 -597
rect 405 -665 461 -631
rect 405 -699 416 -665
rect 450 -699 461 -665
rect 405 -711 461 -699
rect 491 287 547 299
rect 491 253 502 287
rect 536 253 547 287
rect 491 219 547 253
rect 491 185 502 219
rect 536 185 547 219
rect 491 151 547 185
rect 491 117 502 151
rect 536 117 547 151
rect 491 83 547 117
rect 491 49 502 83
rect 536 49 547 83
rect 491 15 547 49
rect 491 -19 502 15
rect 536 -19 547 15
rect 491 -53 547 -19
rect 491 -87 502 -53
rect 536 -87 547 -53
rect 491 -121 547 -87
rect 491 -155 502 -121
rect 536 -155 547 -121
rect 491 -189 547 -155
rect 491 -223 502 -189
rect 536 -223 547 -189
rect 491 -257 547 -223
rect 491 -291 502 -257
rect 536 -291 547 -257
rect 491 -325 547 -291
rect 491 -359 502 -325
rect 536 -359 547 -325
rect 491 -393 547 -359
rect 491 -427 502 -393
rect 536 -427 547 -393
rect 491 -461 547 -427
rect 491 -495 502 -461
rect 536 -495 547 -461
rect 491 -529 547 -495
rect 491 -563 502 -529
rect 536 -563 547 -529
rect 491 -597 547 -563
rect 491 -631 502 -597
rect 536 -631 547 -597
rect 491 -665 547 -631
rect 491 -699 502 -665
rect 536 -699 547 -665
rect 491 -711 547 -699
rect 577 287 633 299
rect 577 253 588 287
rect 622 253 633 287
rect 577 219 633 253
rect 577 185 588 219
rect 622 185 633 219
rect 577 151 633 185
rect 577 117 588 151
rect 622 117 633 151
rect 577 83 633 117
rect 577 49 588 83
rect 622 49 633 83
rect 577 15 633 49
rect 577 -19 588 15
rect 622 -19 633 15
rect 577 -53 633 -19
rect 577 -87 588 -53
rect 622 -87 633 -53
rect 577 -121 633 -87
rect 577 -155 588 -121
rect 622 -155 633 -121
rect 577 -189 633 -155
rect 577 -223 588 -189
rect 622 -223 633 -189
rect 577 -257 633 -223
rect 577 -291 588 -257
rect 622 -291 633 -257
rect 577 -325 633 -291
rect 577 -359 588 -325
rect 622 -359 633 -325
rect 577 -393 633 -359
rect 577 -427 588 -393
rect 622 -427 633 -393
rect 577 -461 633 -427
rect 577 -495 588 -461
rect 622 -495 633 -461
rect 577 -529 633 -495
rect 577 -563 588 -529
rect 622 -563 633 -529
rect 577 -597 633 -563
rect 577 -631 588 -597
rect 622 -631 633 -597
rect 577 -665 633 -631
rect 577 -699 588 -665
rect 622 -699 633 -665
rect 577 -711 633 -699
rect 663 287 719 299
rect 663 253 674 287
rect 708 253 719 287
rect 663 219 719 253
rect 663 185 674 219
rect 708 185 719 219
rect 663 151 719 185
rect 663 117 674 151
rect 708 117 719 151
rect 663 83 719 117
rect 663 49 674 83
rect 708 49 719 83
rect 663 15 719 49
rect 663 -19 674 15
rect 708 -19 719 15
rect 663 -53 719 -19
rect 663 -87 674 -53
rect 708 -87 719 -53
rect 663 -121 719 -87
rect 663 -155 674 -121
rect 708 -155 719 -121
rect 663 -189 719 -155
rect 663 -223 674 -189
rect 708 -223 719 -189
rect 663 -257 719 -223
rect 663 -291 674 -257
rect 708 -291 719 -257
rect 663 -325 719 -291
rect 663 -359 674 -325
rect 708 -359 719 -325
rect 663 -393 719 -359
rect 663 -427 674 -393
rect 708 -427 719 -393
rect 663 -461 719 -427
rect 663 -495 674 -461
rect 708 -495 719 -461
rect 663 -529 719 -495
rect 663 -563 674 -529
rect 708 -563 719 -529
rect 663 -597 719 -563
rect 663 -631 674 -597
rect 708 -631 719 -597
rect 663 -665 719 -631
rect 663 -699 674 -665
rect 708 -699 719 -665
rect 663 -711 719 -699
rect 749 287 805 299
rect 749 253 760 287
rect 794 253 805 287
rect 749 219 805 253
rect 749 185 760 219
rect 794 185 805 219
rect 749 151 805 185
rect 749 117 760 151
rect 794 117 805 151
rect 749 83 805 117
rect 749 49 760 83
rect 794 49 805 83
rect 749 15 805 49
rect 749 -19 760 15
rect 794 -19 805 15
rect 749 -53 805 -19
rect 749 -87 760 -53
rect 794 -87 805 -53
rect 749 -121 805 -87
rect 749 -155 760 -121
rect 794 -155 805 -121
rect 749 -189 805 -155
rect 749 -223 760 -189
rect 794 -223 805 -189
rect 749 -257 805 -223
rect 749 -291 760 -257
rect 794 -291 805 -257
rect 749 -325 805 -291
rect 749 -359 760 -325
rect 794 -359 805 -325
rect 749 -393 805 -359
rect 749 -427 760 -393
rect 794 -427 805 -393
rect 749 -461 805 -427
rect 749 -495 760 -461
rect 794 -495 805 -461
rect 749 -529 805 -495
rect 749 -563 760 -529
rect 794 -563 805 -529
rect 749 -597 805 -563
rect 749 -631 760 -597
rect 794 -631 805 -597
rect 749 -665 805 -631
rect 749 -699 760 -665
rect 794 -699 805 -665
rect 749 -711 805 -699
rect 835 287 891 299
rect 835 253 846 287
rect 880 253 891 287
rect 835 219 891 253
rect 835 185 846 219
rect 880 185 891 219
rect 835 151 891 185
rect 835 117 846 151
rect 880 117 891 151
rect 835 83 891 117
rect 835 49 846 83
rect 880 49 891 83
rect 835 15 891 49
rect 835 -19 846 15
rect 880 -19 891 15
rect 835 -53 891 -19
rect 835 -87 846 -53
rect 880 -87 891 -53
rect 835 -121 891 -87
rect 835 -155 846 -121
rect 880 -155 891 -121
rect 835 -189 891 -155
rect 835 -223 846 -189
rect 880 -223 891 -189
rect 835 -257 891 -223
rect 835 -291 846 -257
rect 880 -291 891 -257
rect 835 -325 891 -291
rect 835 -359 846 -325
rect 880 -359 891 -325
rect 835 -393 891 -359
rect 835 -427 846 -393
rect 880 -427 891 -393
rect 835 -461 891 -427
rect 835 -495 846 -461
rect 880 -495 891 -461
rect 835 -529 891 -495
rect 835 -563 846 -529
rect 880 -563 891 -529
rect 835 -597 891 -563
rect 835 -631 846 -597
rect 880 -631 891 -597
rect 835 -665 891 -631
rect 835 -699 846 -665
rect 880 -699 891 -665
rect 835 -711 891 -699
<< ndiffc >>
rect -6711 17056 -6677 17090
rect -6711 16988 -6677 17022
rect -6711 16920 -6677 16954
rect -6711 16852 -6677 16886
rect -6711 16784 -6677 16818
rect -6711 16716 -6677 16750
rect -6711 16648 -6677 16682
rect -6711 16580 -6677 16614
rect -6711 16512 -6677 16546
rect -6711 16444 -6677 16478
rect -6711 16376 -6677 16410
rect -6711 16308 -6677 16342
rect -6711 16240 -6677 16274
rect -6711 16172 -6677 16206
rect -6711 16104 -6677 16138
rect -6625 17056 -6591 17090
rect -6625 16988 -6591 17022
rect -6625 16920 -6591 16954
rect -6625 16852 -6591 16886
rect -6625 16784 -6591 16818
rect -6625 16716 -6591 16750
rect -6625 16648 -6591 16682
rect -6625 16580 -6591 16614
rect -6625 16512 -6591 16546
rect -6625 16444 -6591 16478
rect -6625 16376 -6591 16410
rect -6625 16308 -6591 16342
rect -6625 16240 -6591 16274
rect -6625 16172 -6591 16206
rect -6625 16104 -6591 16138
rect -6539 17056 -6505 17090
rect -6539 16988 -6505 17022
rect -6539 16920 -6505 16954
rect -6539 16852 -6505 16886
rect -6539 16784 -6505 16818
rect -6539 16716 -6505 16750
rect -6539 16648 -6505 16682
rect -6539 16580 -6505 16614
rect -6539 16512 -6505 16546
rect -6539 16444 -6505 16478
rect -6539 16376 -6505 16410
rect -6539 16308 -6505 16342
rect -6539 16240 -6505 16274
rect -6539 16172 -6505 16206
rect -6539 16104 -6505 16138
rect -6317 17056 -6283 17090
rect -6317 16988 -6283 17022
rect -6317 16920 -6283 16954
rect -6317 16852 -6283 16886
rect -6317 16784 -6283 16818
rect -6317 16716 -6283 16750
rect -6317 16648 -6283 16682
rect -6317 16580 -6283 16614
rect -6317 16512 -6283 16546
rect -6317 16444 -6283 16478
rect -6317 16376 -6283 16410
rect -6317 16308 -6283 16342
rect -6317 16240 -6283 16274
rect -6317 16172 -6283 16206
rect -6317 16104 -6283 16138
rect -6231 17056 -6197 17090
rect -6231 16988 -6197 17022
rect -6231 16920 -6197 16954
rect -6231 16852 -6197 16886
rect -6231 16784 -6197 16818
rect -6231 16716 -6197 16750
rect -6231 16648 -6197 16682
rect -6231 16580 -6197 16614
rect -6231 16512 -6197 16546
rect -6231 16444 -6197 16478
rect -6231 16376 -6197 16410
rect -6231 16308 -6197 16342
rect -6231 16240 -6197 16274
rect -6231 16172 -6197 16206
rect -6231 16104 -6197 16138
rect -6145 17056 -6111 17090
rect -6145 16988 -6111 17022
rect -6145 16920 -6111 16954
rect -6145 16852 -6111 16886
rect -6145 16784 -6111 16818
rect -6145 16716 -6111 16750
rect -6145 16648 -6111 16682
rect -6145 16580 -6111 16614
rect -6145 16512 -6111 16546
rect -6145 16444 -6111 16478
rect -6145 16376 -6111 16410
rect -6145 16308 -6111 16342
rect -6145 16240 -6111 16274
rect -6145 16172 -6111 16206
rect -6145 16104 -6111 16138
rect -5923 17056 -5889 17090
rect -5923 16988 -5889 17022
rect -5923 16920 -5889 16954
rect -5923 16852 -5889 16886
rect -5923 16784 -5889 16818
rect -5923 16716 -5889 16750
rect -5923 16648 -5889 16682
rect -5923 16580 -5889 16614
rect -5923 16512 -5889 16546
rect -5923 16444 -5889 16478
rect -5923 16376 -5889 16410
rect -5923 16308 -5889 16342
rect -5923 16240 -5889 16274
rect -5923 16172 -5889 16206
rect -5923 16104 -5889 16138
rect -5837 17056 -5803 17090
rect -5837 16988 -5803 17022
rect -5837 16920 -5803 16954
rect -5837 16852 -5803 16886
rect -5837 16784 -5803 16818
rect -5837 16716 -5803 16750
rect -5837 16648 -5803 16682
rect -5837 16580 -5803 16614
rect -5837 16512 -5803 16546
rect -5837 16444 -5803 16478
rect -5837 16376 -5803 16410
rect -5837 16308 -5803 16342
rect -5837 16240 -5803 16274
rect -5837 16172 -5803 16206
rect -5837 16104 -5803 16138
rect -5751 17056 -5717 17090
rect -5751 16988 -5717 17022
rect -5751 16920 -5717 16954
rect -5751 16852 -5717 16886
rect -5751 16784 -5717 16818
rect -5751 16716 -5717 16750
rect -5751 16648 -5717 16682
rect -5751 16580 -5717 16614
rect -5751 16512 -5717 16546
rect -5751 16444 -5717 16478
rect -5751 16376 -5717 16410
rect -5751 16308 -5717 16342
rect -5751 16240 -5717 16274
rect -5751 16172 -5717 16206
rect -5751 16104 -5717 16138
rect -5529 17056 -5495 17090
rect -5529 16988 -5495 17022
rect -5529 16920 -5495 16954
rect -5529 16852 -5495 16886
rect -5529 16784 -5495 16818
rect -5529 16716 -5495 16750
rect -5529 16648 -5495 16682
rect -5529 16580 -5495 16614
rect -5529 16512 -5495 16546
rect -5529 16444 -5495 16478
rect -5529 16376 -5495 16410
rect -5529 16308 -5495 16342
rect -5529 16240 -5495 16274
rect -5529 16172 -5495 16206
rect -5529 16104 -5495 16138
rect -5443 17056 -5409 17090
rect -5443 16988 -5409 17022
rect -5443 16920 -5409 16954
rect -5443 16852 -5409 16886
rect -5443 16784 -5409 16818
rect -5443 16716 -5409 16750
rect -5443 16648 -5409 16682
rect -5443 16580 -5409 16614
rect -5443 16512 -5409 16546
rect -5443 16444 -5409 16478
rect -5443 16376 -5409 16410
rect -5443 16308 -5409 16342
rect -5443 16240 -5409 16274
rect -5443 16172 -5409 16206
rect -5443 16104 -5409 16138
rect -5357 17056 -5323 17090
rect -5357 16988 -5323 17022
rect -5357 16920 -5323 16954
rect -5357 16852 -5323 16886
rect -5357 16784 -5323 16818
rect -5357 16716 -5323 16750
rect -5357 16648 -5323 16682
rect -5357 16580 -5323 16614
rect -5357 16512 -5323 16546
rect -5357 16444 -5323 16478
rect -5357 16376 -5323 16410
rect -5357 16308 -5323 16342
rect -5357 16240 -5323 16274
rect -5357 16172 -5323 16206
rect -5357 16104 -5323 16138
rect -46 8445 -12 8479
rect -46 8377 -12 8411
rect -46 8309 -12 8343
rect -46 8241 -12 8275
rect -46 8173 -12 8207
rect -46 8105 -12 8139
rect -46 8037 -12 8071
rect -46 7969 -12 8003
rect -46 7901 -12 7935
rect -46 7833 -12 7867
rect -46 7765 -12 7799
rect -46 7697 -12 7731
rect -46 7629 -12 7663
rect -46 7561 -12 7595
rect -46 7493 -12 7527
rect 40 8445 74 8479
rect 40 8377 74 8411
rect 40 8309 74 8343
rect 40 8241 74 8275
rect 40 8173 74 8207
rect 40 8105 74 8139
rect 40 8037 74 8071
rect 40 7969 74 8003
rect 40 7901 74 7935
rect 40 7833 74 7867
rect 40 7765 74 7799
rect 40 7697 74 7731
rect 40 7629 74 7663
rect 40 7561 74 7595
rect 40 7493 74 7527
rect 126 8445 160 8479
rect 126 8377 160 8411
rect 126 8309 160 8343
rect 126 8241 160 8275
rect 126 8173 160 8207
rect 126 8105 160 8139
rect 126 8037 160 8071
rect 126 7969 160 8003
rect 126 7901 160 7935
rect 126 7833 160 7867
rect 126 7765 160 7799
rect 126 7697 160 7731
rect 126 7629 160 7663
rect 126 7561 160 7595
rect 126 7493 160 7527
rect 212 8445 246 8479
rect 212 8377 246 8411
rect 212 8309 246 8343
rect 212 8241 246 8275
rect 212 8173 246 8207
rect 212 8105 246 8139
rect 212 8037 246 8071
rect 212 7969 246 8003
rect 212 7901 246 7935
rect 212 7833 246 7867
rect 212 7765 246 7799
rect 212 7697 246 7731
rect 212 7629 246 7663
rect 212 7561 246 7595
rect 212 7493 246 7527
rect 298 8445 332 8479
rect 298 8377 332 8411
rect 298 8309 332 8343
rect 298 8241 332 8275
rect 298 8173 332 8207
rect 298 8105 332 8139
rect 298 8037 332 8071
rect 298 7969 332 8003
rect 298 7901 332 7935
rect 298 7833 332 7867
rect 298 7765 332 7799
rect 298 7697 332 7731
rect 298 7629 332 7663
rect 298 7561 332 7595
rect 298 7493 332 7527
rect 384 8445 418 8479
rect 384 8377 418 8411
rect 384 8309 418 8343
rect 384 8241 418 8275
rect 384 8173 418 8207
rect 384 8105 418 8139
rect 384 8037 418 8071
rect 384 7969 418 8003
rect 384 7901 418 7935
rect 384 7833 418 7867
rect 384 7765 418 7799
rect 384 7697 418 7731
rect 384 7629 418 7663
rect 384 7561 418 7595
rect 384 7493 418 7527
rect 470 8445 504 8479
rect 470 8377 504 8411
rect 470 8309 504 8343
rect 470 8241 504 8275
rect 470 8173 504 8207
rect 470 8105 504 8139
rect 470 8037 504 8071
rect 470 7969 504 8003
rect 470 7901 504 7935
rect 470 7833 504 7867
rect 470 7765 504 7799
rect 470 7697 504 7731
rect 470 7629 504 7663
rect 470 7561 504 7595
rect 470 7493 504 7527
rect 556 8445 590 8479
rect 556 8377 590 8411
rect 556 8309 590 8343
rect 556 8241 590 8275
rect 556 8173 590 8207
rect 556 8105 590 8139
rect 556 8037 590 8071
rect 556 7969 590 8003
rect 556 7901 590 7935
rect 556 7833 590 7867
rect 556 7765 590 7799
rect 556 7697 590 7731
rect 556 7629 590 7663
rect 556 7561 590 7595
rect 556 7493 590 7527
rect 642 8445 676 8479
rect 642 8377 676 8411
rect 642 8309 676 8343
rect 642 8241 676 8275
rect 642 8173 676 8207
rect 642 8105 676 8139
rect 642 8037 676 8071
rect 642 7969 676 8003
rect 642 7901 676 7935
rect 642 7833 676 7867
rect 642 7765 676 7799
rect 642 7697 676 7731
rect 642 7629 676 7663
rect 642 7561 676 7595
rect 642 7493 676 7527
rect 728 8445 762 8479
rect 728 8377 762 8411
rect 728 8309 762 8343
rect 728 8241 762 8275
rect 728 8173 762 8207
rect 728 8105 762 8139
rect 728 8037 762 8071
rect 728 7969 762 8003
rect 728 7901 762 7935
rect 728 7833 762 7867
rect 728 7765 762 7799
rect 728 7697 762 7731
rect 728 7629 762 7663
rect 728 7561 762 7595
rect 728 7493 762 7527
rect 814 8445 848 8479
rect 814 8377 848 8411
rect 814 8309 848 8343
rect 814 8241 848 8275
rect 814 8173 848 8207
rect 814 8105 848 8139
rect 814 8037 848 8071
rect 814 7969 848 8003
rect 814 7901 848 7935
rect 814 7833 848 7867
rect 814 7765 848 7799
rect 814 7697 848 7731
rect 814 7629 848 7663
rect 814 7561 848 7595
rect 814 7493 848 7527
rect 900 8445 934 8479
rect 900 8377 934 8411
rect 900 8309 934 8343
rect 900 8241 934 8275
rect 900 8173 934 8207
rect 900 8105 934 8139
rect 900 8037 934 8071
rect 900 7969 934 8003
rect 900 7901 934 7935
rect 900 7833 934 7867
rect 900 7765 934 7799
rect 900 7697 934 7731
rect 900 7629 934 7663
rect 900 7561 934 7595
rect 900 7493 934 7527
rect 986 8445 1020 8479
rect 986 8377 1020 8411
rect 986 8309 1020 8343
rect 986 8241 1020 8275
rect 986 8173 1020 8207
rect 986 8105 1020 8139
rect 986 8037 1020 8071
rect 986 7969 1020 8003
rect 986 7901 1020 7935
rect 986 7833 1020 7867
rect 986 7765 1020 7799
rect 986 7697 1020 7731
rect 986 7629 1020 7663
rect 986 7561 1020 7595
rect 986 7493 1020 7527
rect 158 253 192 287
rect 158 185 192 219
rect 158 117 192 151
rect 158 49 192 83
rect 158 -19 192 15
rect 158 -87 192 -53
rect 158 -155 192 -121
rect 158 -223 192 -189
rect 158 -291 192 -257
rect 158 -359 192 -325
rect 158 -427 192 -393
rect 158 -495 192 -461
rect 158 -563 192 -529
rect 158 -631 192 -597
rect 158 -699 192 -665
rect 244 253 278 287
rect 244 185 278 219
rect 244 117 278 151
rect 244 49 278 83
rect 244 -19 278 15
rect 244 -87 278 -53
rect 244 -155 278 -121
rect 244 -223 278 -189
rect 244 -291 278 -257
rect 244 -359 278 -325
rect 244 -427 278 -393
rect 244 -495 278 -461
rect 244 -563 278 -529
rect 244 -631 278 -597
rect 244 -699 278 -665
rect 330 253 364 287
rect 330 185 364 219
rect 330 117 364 151
rect 330 49 364 83
rect 330 -19 364 15
rect 330 -87 364 -53
rect 330 -155 364 -121
rect 330 -223 364 -189
rect 330 -291 364 -257
rect 330 -359 364 -325
rect 330 -427 364 -393
rect 330 -495 364 -461
rect 330 -563 364 -529
rect 330 -631 364 -597
rect 330 -699 364 -665
rect 416 253 450 287
rect 416 185 450 219
rect 416 117 450 151
rect 416 49 450 83
rect 416 -19 450 15
rect 416 -87 450 -53
rect 416 -155 450 -121
rect 416 -223 450 -189
rect 416 -291 450 -257
rect 416 -359 450 -325
rect 416 -427 450 -393
rect 416 -495 450 -461
rect 416 -563 450 -529
rect 416 -631 450 -597
rect 416 -699 450 -665
rect 502 253 536 287
rect 502 185 536 219
rect 502 117 536 151
rect 502 49 536 83
rect 502 -19 536 15
rect 502 -87 536 -53
rect 502 -155 536 -121
rect 502 -223 536 -189
rect 502 -291 536 -257
rect 502 -359 536 -325
rect 502 -427 536 -393
rect 502 -495 536 -461
rect 502 -563 536 -529
rect 502 -631 536 -597
rect 502 -699 536 -665
rect 588 253 622 287
rect 588 185 622 219
rect 588 117 622 151
rect 588 49 622 83
rect 588 -19 622 15
rect 588 -87 622 -53
rect 588 -155 622 -121
rect 588 -223 622 -189
rect 588 -291 622 -257
rect 588 -359 622 -325
rect 588 -427 622 -393
rect 588 -495 622 -461
rect 588 -563 622 -529
rect 588 -631 622 -597
rect 588 -699 622 -665
rect 674 253 708 287
rect 674 185 708 219
rect 674 117 708 151
rect 674 49 708 83
rect 674 -19 708 15
rect 674 -87 708 -53
rect 674 -155 708 -121
rect 674 -223 708 -189
rect 674 -291 708 -257
rect 674 -359 708 -325
rect 674 -427 708 -393
rect 674 -495 708 -461
rect 674 -563 708 -529
rect 674 -631 708 -597
rect 674 -699 708 -665
rect 760 253 794 287
rect 760 185 794 219
rect 760 117 794 151
rect 760 49 794 83
rect 760 -19 794 15
rect 760 -87 794 -53
rect 760 -155 794 -121
rect 760 -223 794 -189
rect 760 -291 794 -257
rect 760 -359 794 -325
rect 760 -427 794 -393
rect 760 -495 794 -461
rect 760 -563 794 -529
rect 760 -631 794 -597
rect 760 -699 794 -665
rect 846 253 880 287
rect 846 185 880 219
rect 846 117 880 151
rect 846 49 880 83
rect 846 -19 880 15
rect 846 -87 880 -53
rect 846 -155 880 -121
rect 846 -223 880 -189
rect 846 -291 880 -257
rect 846 -359 880 -325
rect 846 -427 880 -393
rect 846 -495 880 -461
rect 846 -563 880 -529
rect 846 -631 880 -597
rect 846 -699 880 -665
<< psubdiff >>
rect -6834 17056 -6776 17102
rect -6834 17022 -6822 17056
rect -6788 17022 -6776 17056
rect -6834 16988 -6776 17022
rect -6834 16954 -6822 16988
rect -6788 16954 -6776 16988
rect -6834 16920 -6776 16954
rect -6834 16886 -6822 16920
rect -6788 16886 -6776 16920
rect -6834 16852 -6776 16886
rect -6834 16818 -6822 16852
rect -6788 16818 -6776 16852
rect -6834 16784 -6776 16818
rect -6834 16750 -6822 16784
rect -6788 16750 -6776 16784
rect -6834 16716 -6776 16750
rect -6834 16682 -6822 16716
rect -6788 16682 -6776 16716
rect -6834 16648 -6776 16682
rect -6834 16614 -6822 16648
rect -6788 16614 -6776 16648
rect -6834 16580 -6776 16614
rect -6834 16546 -6822 16580
rect -6788 16546 -6776 16580
rect -6834 16512 -6776 16546
rect -6834 16478 -6822 16512
rect -6788 16478 -6776 16512
rect -6834 16444 -6776 16478
rect -6834 16410 -6822 16444
rect -6788 16410 -6776 16444
rect -6834 16376 -6776 16410
rect -6834 16342 -6822 16376
rect -6788 16342 -6776 16376
rect -6834 16308 -6776 16342
rect -6834 16274 -6822 16308
rect -6788 16274 -6776 16308
rect -6834 16240 -6776 16274
rect -6834 16206 -6822 16240
rect -6788 16206 -6776 16240
rect -6834 16172 -6776 16206
rect -6834 16138 -6822 16172
rect -6788 16138 -6776 16172
rect -6834 16092 -6776 16138
rect -6440 17056 -6382 17102
rect -6440 17022 -6428 17056
rect -6394 17022 -6382 17056
rect -6440 16988 -6382 17022
rect -6440 16954 -6428 16988
rect -6394 16954 -6382 16988
rect -6440 16920 -6382 16954
rect -6440 16886 -6428 16920
rect -6394 16886 -6382 16920
rect -6440 16852 -6382 16886
rect -6440 16818 -6428 16852
rect -6394 16818 -6382 16852
rect -6440 16784 -6382 16818
rect -6440 16750 -6428 16784
rect -6394 16750 -6382 16784
rect -6440 16716 -6382 16750
rect -6440 16682 -6428 16716
rect -6394 16682 -6382 16716
rect -6440 16648 -6382 16682
rect -6440 16614 -6428 16648
rect -6394 16614 -6382 16648
rect -6440 16580 -6382 16614
rect -6440 16546 -6428 16580
rect -6394 16546 -6382 16580
rect -6440 16512 -6382 16546
rect -6440 16478 -6428 16512
rect -6394 16478 -6382 16512
rect -6440 16444 -6382 16478
rect -6440 16410 -6428 16444
rect -6394 16410 -6382 16444
rect -6440 16376 -6382 16410
rect -6440 16342 -6428 16376
rect -6394 16342 -6382 16376
rect -6440 16308 -6382 16342
rect -6440 16274 -6428 16308
rect -6394 16274 -6382 16308
rect -6440 16240 -6382 16274
rect -6440 16206 -6428 16240
rect -6394 16206 -6382 16240
rect -6440 16172 -6382 16206
rect -6440 16138 -6428 16172
rect -6394 16138 -6382 16172
rect -6440 16092 -6382 16138
rect -6046 17056 -5988 17102
rect -6046 17022 -6034 17056
rect -6000 17022 -5988 17056
rect -6046 16988 -5988 17022
rect -6046 16954 -6034 16988
rect -6000 16954 -5988 16988
rect -6046 16920 -5988 16954
rect -6046 16886 -6034 16920
rect -6000 16886 -5988 16920
rect -6046 16852 -5988 16886
rect -6046 16818 -6034 16852
rect -6000 16818 -5988 16852
rect -6046 16784 -5988 16818
rect -6046 16750 -6034 16784
rect -6000 16750 -5988 16784
rect -6046 16716 -5988 16750
rect -6046 16682 -6034 16716
rect -6000 16682 -5988 16716
rect -6046 16648 -5988 16682
rect -6046 16614 -6034 16648
rect -6000 16614 -5988 16648
rect -6046 16580 -5988 16614
rect -6046 16546 -6034 16580
rect -6000 16546 -5988 16580
rect -6046 16512 -5988 16546
rect -6046 16478 -6034 16512
rect -6000 16478 -5988 16512
rect -6046 16444 -5988 16478
rect -6046 16410 -6034 16444
rect -6000 16410 -5988 16444
rect -6046 16376 -5988 16410
rect -6046 16342 -6034 16376
rect -6000 16342 -5988 16376
rect -6046 16308 -5988 16342
rect -6046 16274 -6034 16308
rect -6000 16274 -5988 16308
rect -6046 16240 -5988 16274
rect -6046 16206 -6034 16240
rect -6000 16206 -5988 16240
rect -6046 16172 -5988 16206
rect -6046 16138 -6034 16172
rect -6000 16138 -5988 16172
rect -6046 16092 -5988 16138
rect -5652 17056 -5594 17102
rect -5652 17022 -5640 17056
rect -5606 17022 -5594 17056
rect -5652 16988 -5594 17022
rect -5652 16954 -5640 16988
rect -5606 16954 -5594 16988
rect -5652 16920 -5594 16954
rect -5652 16886 -5640 16920
rect -5606 16886 -5594 16920
rect -5652 16852 -5594 16886
rect -5652 16818 -5640 16852
rect -5606 16818 -5594 16852
rect -5652 16784 -5594 16818
rect -5652 16750 -5640 16784
rect -5606 16750 -5594 16784
rect -5652 16716 -5594 16750
rect -5652 16682 -5640 16716
rect -5606 16682 -5594 16716
rect -5652 16648 -5594 16682
rect -5652 16614 -5640 16648
rect -5606 16614 -5594 16648
rect -5652 16580 -5594 16614
rect -5652 16546 -5640 16580
rect -5606 16546 -5594 16580
rect -5652 16512 -5594 16546
rect -5652 16478 -5640 16512
rect -5606 16478 -5594 16512
rect -5652 16444 -5594 16478
rect -5652 16410 -5640 16444
rect -5606 16410 -5594 16444
rect -5652 16376 -5594 16410
rect -5652 16342 -5640 16376
rect -5606 16342 -5594 16376
rect -5652 16308 -5594 16342
rect -5652 16274 -5640 16308
rect -5606 16274 -5594 16308
rect -5652 16240 -5594 16274
rect -5652 16206 -5640 16240
rect -5606 16206 -5594 16240
rect -5652 16172 -5594 16206
rect -5652 16138 -5640 16172
rect -5606 16138 -5594 16172
rect -5652 16092 -5594 16138
rect -5258 17056 -5200 17102
rect -5258 17022 -5246 17056
rect -5212 17022 -5200 17056
rect -5258 16988 -5200 17022
rect -5258 16954 -5246 16988
rect -5212 16954 -5200 16988
rect -5258 16920 -5200 16954
rect -5258 16886 -5246 16920
rect -5212 16886 -5200 16920
rect -5258 16852 -5200 16886
rect -5258 16818 -5246 16852
rect -5212 16818 -5200 16852
rect -5258 16784 -5200 16818
rect -5258 16750 -5246 16784
rect -5212 16750 -5200 16784
rect -5258 16716 -5200 16750
rect -5258 16682 -5246 16716
rect -5212 16682 -5200 16716
rect -5258 16648 -5200 16682
rect -5258 16614 -5246 16648
rect -5212 16614 -5200 16648
rect -5258 16580 -5200 16614
rect -5258 16546 -5246 16580
rect -5212 16546 -5200 16580
rect -5258 16512 -5200 16546
rect -5258 16478 -5246 16512
rect -5212 16478 -5200 16512
rect -5258 16444 -5200 16478
rect -5258 16410 -5246 16444
rect -5212 16410 -5200 16444
rect -5258 16376 -5200 16410
rect -5258 16342 -5246 16376
rect -5212 16342 -5200 16376
rect -5258 16308 -5200 16342
rect -5258 16274 -5246 16308
rect -5212 16274 -5200 16308
rect -5258 16240 -5200 16274
rect -5258 16206 -5246 16240
rect -5212 16206 -5200 16240
rect -5258 16172 -5200 16206
rect -5258 16138 -5246 16172
rect -5212 16138 -5200 16172
rect -5258 16092 -5200 16138
rect -2064 8816 -1968 8850
rect -1618 8816 -1522 8850
rect -2064 8754 -2030 8816
rect -1556 8754 -1522 8816
rect -2064 7470 -2030 7532
rect -1556 7470 -1522 7532
rect -2064 7436 -1968 7470
rect -1618 7436 -1522 7470
rect -194 8454 -124 8490
rect -194 8420 -174 8454
rect -140 8420 -124 8454
rect -194 8384 -124 8420
rect -194 8350 -174 8384
rect -140 8350 -124 8384
rect -194 8314 -124 8350
rect -194 8280 -174 8314
rect -140 8280 -124 8314
rect -194 8244 -124 8280
rect -194 8210 -174 8244
rect -140 8210 -124 8244
rect -194 8174 -124 8210
rect -194 8140 -174 8174
rect -140 8140 -124 8174
rect -194 8104 -124 8140
rect -194 8070 -174 8104
rect -140 8070 -124 8104
rect -194 8034 -124 8070
rect -194 8000 -174 8034
rect -140 8000 -124 8034
rect -194 7964 -124 8000
rect -194 7930 -174 7964
rect -140 7930 -124 7964
rect -194 7894 -124 7930
rect -194 7860 -174 7894
rect -140 7860 -124 7894
rect -194 7824 -124 7860
rect -194 7790 -174 7824
rect -140 7790 -124 7824
rect -194 7754 -124 7790
rect -194 7720 -174 7754
rect -140 7720 -124 7754
rect -194 7684 -124 7720
rect -194 7650 -174 7684
rect -140 7650 -124 7684
rect -194 7614 -124 7650
rect -194 7580 -174 7614
rect -140 7580 -124 7614
rect -194 7544 -124 7580
rect -194 7510 -174 7544
rect -140 7510 -124 7544
rect -194 7474 -124 7510
rect 1096 8454 1176 8490
rect 1096 8420 1116 8454
rect 1150 8420 1176 8454
rect 1096 8384 1176 8420
rect 1096 8350 1116 8384
rect 1150 8350 1176 8384
rect 1096 8314 1176 8350
rect 1096 8280 1116 8314
rect 1150 8280 1176 8314
rect 1096 8244 1176 8280
rect 1096 8210 1116 8244
rect 1150 8210 1176 8244
rect 1096 8174 1176 8210
rect 1096 8140 1116 8174
rect 1150 8140 1176 8174
rect 1096 8104 1176 8140
rect 1096 8070 1116 8104
rect 1150 8070 1176 8104
rect 1096 8034 1176 8070
rect 1096 8000 1116 8034
rect 1150 8000 1176 8034
rect 1096 7964 1176 8000
rect 1096 7930 1116 7964
rect 1150 7930 1176 7964
rect 1096 7894 1176 7930
rect 1096 7860 1116 7894
rect 1150 7860 1176 7894
rect 1096 7824 1176 7860
rect 1096 7790 1116 7824
rect 1150 7790 1176 7824
rect 1096 7754 1176 7790
rect 1096 7720 1116 7754
rect 1150 7720 1176 7754
rect 1096 7684 1176 7720
rect 1096 7650 1116 7684
rect 1150 7650 1176 7684
rect 1096 7614 1176 7650
rect 1096 7580 1116 7614
rect 1150 7580 1176 7614
rect 1096 7544 1176 7580
rect 1096 7510 1116 7544
rect 1150 7510 1176 7544
rect -194 7440 -174 7474
rect -140 7440 -124 7474
rect -194 7410 -124 7440
rect 1096 7474 1176 7510
rect 1096 7440 1116 7474
rect 1150 7440 1176 7474
rect 1096 7410 1176 7440
rect -194 7384 1176 7410
rect -194 7350 -94 7384
rect -60 7350 -24 7384
rect 10 7350 46 7384
rect 80 7350 116 7384
rect 150 7350 186 7384
rect 220 7350 256 7384
rect 290 7350 326 7384
rect 360 7350 396 7384
rect 430 7350 466 7384
rect 500 7350 536 7384
rect 570 7350 606 7384
rect 640 7350 676 7384
rect 710 7350 746 7384
rect 780 7350 816 7384
rect 850 7350 886 7384
rect 920 7350 956 7384
rect 990 7350 1026 7384
rect 1060 7350 1176 7384
rect -194 7330 1176 7350
rect -1264 7056 -1168 7090
rect -818 7056 -722 7090
rect -1264 6994 -1230 7056
rect -756 6994 -722 7056
rect -1264 5710 -1230 5772
rect -756 5710 -722 5772
rect -1264 5676 -1168 5710
rect -818 5676 -722 5710
rect 10 430 1030 450
rect 10 390 50 430
rect 990 390 1030 430
rect 10 370 1030 390
rect 10 340 80 370
rect 10 306 30 340
rect 64 306 80 340
rect 10 270 80 306
rect 947 340 1027 370
rect 947 306 967 340
rect 1001 306 1027 340
rect 10 236 30 270
rect 64 236 80 270
rect 10 200 80 236
rect 10 166 30 200
rect 64 166 80 200
rect 10 130 80 166
rect 10 96 30 130
rect 64 96 80 130
rect 10 60 80 96
rect 10 26 30 60
rect 64 26 80 60
rect 10 -10 80 26
rect 10 -44 30 -10
rect 64 -44 80 -10
rect 10 -80 80 -44
rect 10 -114 30 -80
rect 64 -114 80 -80
rect 10 -150 80 -114
rect 10 -184 30 -150
rect 64 -184 80 -150
rect 10 -220 80 -184
rect 10 -254 30 -220
rect 64 -254 80 -220
rect 10 -290 80 -254
rect 10 -324 30 -290
rect 64 -324 80 -290
rect 10 -360 80 -324
rect 10 -394 30 -360
rect 64 -394 80 -360
rect 10 -430 80 -394
rect 10 -464 30 -430
rect 64 -464 80 -430
rect 10 -500 80 -464
rect 10 -534 30 -500
rect 64 -534 80 -500
rect 10 -570 80 -534
rect 10 -604 30 -570
rect 64 -604 80 -570
rect -4364 -660 -4268 -626
rect -3810 -660 -3714 -626
rect -4364 -722 -4330 -660
rect -3748 -722 -3714 -660
rect 10 -640 80 -604
rect 10 -674 30 -640
rect 64 -674 80 -640
rect 10 -710 80 -674
rect 947 270 1027 306
rect 947 236 967 270
rect 1001 236 1027 270
rect 947 200 1027 236
rect 947 166 967 200
rect 1001 166 1027 200
rect 947 130 1027 166
rect 947 96 967 130
rect 1001 96 1027 130
rect 947 60 1027 96
rect 947 26 967 60
rect 1001 26 1027 60
rect 947 -10 1027 26
rect 947 -44 967 -10
rect 1001 -44 1027 -10
rect 947 -80 1027 -44
rect 947 -114 967 -80
rect 1001 -114 1027 -80
rect 947 -150 1027 -114
rect 947 -184 967 -150
rect 1001 -184 1027 -150
rect 947 -220 1027 -184
rect 947 -254 967 -220
rect 1001 -254 1027 -220
rect 947 -290 1027 -254
rect 947 -324 967 -290
rect 1001 -324 1027 -290
rect 947 -360 1027 -324
rect 947 -394 967 -360
rect 1001 -394 1027 -360
rect 947 -430 1027 -394
rect 947 -464 967 -430
rect 1001 -464 1027 -430
rect 947 -500 1027 -464
rect 947 -534 967 -500
rect 1001 -534 1027 -500
rect 947 -570 1027 -534
rect 947 -604 967 -570
rect 1001 -604 1027 -570
rect 947 -640 1027 -604
rect 947 -674 967 -640
rect 1001 -674 1027 -640
rect 947 -710 1027 -674
rect -4364 -2030 -4330 -1968
rect -3748 -2030 -3714 -1968
rect -4364 -2064 -4268 -2030
rect -3810 -2064 -3714 -2030
<< psubdiffcont >>
rect -6822 17022 -6788 17056
rect -6822 16954 -6788 16988
rect -6822 16886 -6788 16920
rect -6822 16818 -6788 16852
rect -6822 16750 -6788 16784
rect -6822 16682 -6788 16716
rect -6822 16614 -6788 16648
rect -6822 16546 -6788 16580
rect -6822 16478 -6788 16512
rect -6822 16410 -6788 16444
rect -6822 16342 -6788 16376
rect -6822 16274 -6788 16308
rect -6822 16206 -6788 16240
rect -6822 16138 -6788 16172
rect -6428 17022 -6394 17056
rect -6428 16954 -6394 16988
rect -6428 16886 -6394 16920
rect -6428 16818 -6394 16852
rect -6428 16750 -6394 16784
rect -6428 16682 -6394 16716
rect -6428 16614 -6394 16648
rect -6428 16546 -6394 16580
rect -6428 16478 -6394 16512
rect -6428 16410 -6394 16444
rect -6428 16342 -6394 16376
rect -6428 16274 -6394 16308
rect -6428 16206 -6394 16240
rect -6428 16138 -6394 16172
rect -6034 17022 -6000 17056
rect -6034 16954 -6000 16988
rect -6034 16886 -6000 16920
rect -6034 16818 -6000 16852
rect -6034 16750 -6000 16784
rect -6034 16682 -6000 16716
rect -6034 16614 -6000 16648
rect -6034 16546 -6000 16580
rect -6034 16478 -6000 16512
rect -6034 16410 -6000 16444
rect -6034 16342 -6000 16376
rect -6034 16274 -6000 16308
rect -6034 16206 -6000 16240
rect -6034 16138 -6000 16172
rect -5640 17022 -5606 17056
rect -5640 16954 -5606 16988
rect -5640 16886 -5606 16920
rect -5640 16818 -5606 16852
rect -5640 16750 -5606 16784
rect -5640 16682 -5606 16716
rect -5640 16614 -5606 16648
rect -5640 16546 -5606 16580
rect -5640 16478 -5606 16512
rect -5640 16410 -5606 16444
rect -5640 16342 -5606 16376
rect -5640 16274 -5606 16308
rect -5640 16206 -5606 16240
rect -5640 16138 -5606 16172
rect -5246 17022 -5212 17056
rect -5246 16954 -5212 16988
rect -5246 16886 -5212 16920
rect -5246 16818 -5212 16852
rect -5246 16750 -5212 16784
rect -5246 16682 -5212 16716
rect -5246 16614 -5212 16648
rect -5246 16546 -5212 16580
rect -5246 16478 -5212 16512
rect -5246 16410 -5212 16444
rect -5246 16342 -5212 16376
rect -5246 16274 -5212 16308
rect -5246 16206 -5212 16240
rect -5246 16138 -5212 16172
rect -1968 8816 -1618 8850
rect -2064 7532 -2030 8754
rect -1556 7532 -1522 8754
rect -1968 7436 -1618 7470
rect -174 8420 -140 8454
rect -174 8350 -140 8384
rect -174 8280 -140 8314
rect -174 8210 -140 8244
rect -174 8140 -140 8174
rect -174 8070 -140 8104
rect -174 8000 -140 8034
rect -174 7930 -140 7964
rect -174 7860 -140 7894
rect -174 7790 -140 7824
rect -174 7720 -140 7754
rect -174 7650 -140 7684
rect -174 7580 -140 7614
rect -174 7510 -140 7544
rect 1116 8420 1150 8454
rect 1116 8350 1150 8384
rect 1116 8280 1150 8314
rect 1116 8210 1150 8244
rect 1116 8140 1150 8174
rect 1116 8070 1150 8104
rect 1116 8000 1150 8034
rect 1116 7930 1150 7964
rect 1116 7860 1150 7894
rect 1116 7790 1150 7824
rect 1116 7720 1150 7754
rect 1116 7650 1150 7684
rect 1116 7580 1150 7614
rect 1116 7510 1150 7544
rect -174 7440 -140 7474
rect 1116 7440 1150 7474
rect -94 7350 -60 7384
rect -24 7350 10 7384
rect 46 7350 80 7384
rect 116 7350 150 7384
rect 186 7350 220 7384
rect 256 7350 290 7384
rect 326 7350 360 7384
rect 396 7350 430 7384
rect 466 7350 500 7384
rect 536 7350 570 7384
rect 606 7350 640 7384
rect 676 7350 710 7384
rect 746 7350 780 7384
rect 816 7350 850 7384
rect 886 7350 920 7384
rect 956 7350 990 7384
rect 1026 7350 1060 7384
rect -1168 7056 -818 7090
rect -1264 5772 -1230 6994
rect -756 5772 -722 6994
rect -1168 5676 -818 5710
rect 50 390 990 430
rect 30 306 64 340
rect 967 306 1001 340
rect 30 236 64 270
rect 30 166 64 200
rect 30 96 64 130
rect 30 26 64 60
rect 30 -44 64 -10
rect 30 -114 64 -80
rect 30 -184 64 -150
rect 30 -254 64 -220
rect 30 -324 64 -290
rect 30 -394 64 -360
rect 30 -464 64 -430
rect 30 -534 64 -500
rect 30 -604 64 -570
rect -4268 -660 -3810 -626
rect -4364 -1968 -4330 -722
rect 30 -674 64 -640
rect 967 236 1001 270
rect 967 166 1001 200
rect 967 96 1001 130
rect 967 26 1001 60
rect 967 -44 1001 -10
rect 967 -114 1001 -80
rect 967 -184 1001 -150
rect 967 -254 1001 -220
rect 967 -324 1001 -290
rect 967 -394 1001 -360
rect 967 -464 1001 -430
rect 967 -534 1001 -500
rect 967 -604 1001 -570
rect 967 -674 1001 -640
rect -3748 -1968 -3714 -722
rect -4268 -2064 -3810 -2030
<< poly >>
rect -6709 17174 -6507 17194
rect -6709 17140 -6693 17174
rect -6659 17140 -6625 17174
rect -6591 17140 -6557 17174
rect -6523 17140 -6507 17174
rect -6709 17124 -6507 17140
rect -6315 17174 -6113 17194
rect -6315 17140 -6299 17174
rect -6265 17140 -6231 17174
rect -6197 17140 -6163 17174
rect -6129 17140 -6113 17174
rect -6315 17124 -6113 17140
rect -5921 17174 -5719 17194
rect -5921 17140 -5905 17174
rect -5871 17140 -5837 17174
rect -5803 17140 -5769 17174
rect -5735 17140 -5719 17174
rect -5921 17124 -5719 17140
rect -5527 17174 -5325 17194
rect -5527 17140 -5511 17174
rect -5477 17140 -5443 17174
rect -5409 17140 -5375 17174
rect -5341 17140 -5325 17174
rect -5527 17124 -5325 17140
rect -6666 17102 -6636 17124
rect -6580 17102 -6550 17124
rect -6272 17102 -6242 17124
rect -6186 17102 -6156 17124
rect -5878 17102 -5848 17124
rect -5792 17102 -5762 17124
rect -5484 17102 -5454 17124
rect -5398 17102 -5368 17124
rect -6666 16070 -6636 16092
rect -6580 16070 -6550 16092
rect -6272 16070 -6242 16092
rect -6186 16070 -6156 16092
rect -5878 16070 -5848 16092
rect -5792 16070 -5762 16092
rect -5484 16070 -5454 16092
rect -5398 16070 -5368 16092
rect -6709 16054 -6507 16070
rect -6709 16020 -6693 16054
rect -6659 16020 -6625 16054
rect -6591 16020 -6557 16054
rect -6523 16020 -6507 16054
rect -6709 16000 -6507 16020
rect -6315 16054 -6113 16070
rect -6315 16020 -6299 16054
rect -6265 16020 -6231 16054
rect -6197 16020 -6163 16054
rect -6129 16020 -6113 16054
rect -6315 16000 -6113 16020
rect -5921 16054 -5719 16070
rect -5921 16020 -5905 16054
rect -5871 16020 -5837 16054
rect -5803 16020 -5769 16054
rect -5735 16020 -5719 16054
rect -5921 16000 -5719 16020
rect -5527 16054 -5325 16070
rect -5527 16020 -5511 16054
rect -5477 16020 -5443 16054
rect -5409 16020 -5375 16054
rect -5341 16020 -5325 16054
rect -5527 16000 -5325 16020
rect -1718 8704 -1652 8720
rect -1718 8670 -1702 8704
rect -1668 8670 -1652 8704
rect -1718 8647 -1652 8670
rect -1934 7616 -1868 7639
rect -1934 7582 -1918 7616
rect -1884 7582 -1868 7616
rect -1934 7566 -1868 7582
rect -26 8563 1021 8583
rect -26 8529 -10 8563
rect 24 8529 58 8563
rect 92 8529 126 8563
rect 160 8529 194 8563
rect 228 8529 262 8563
rect 296 8529 330 8563
rect 364 8529 402 8563
rect 436 8529 470 8563
rect 504 8529 538 8563
rect 572 8529 606 8563
rect 640 8529 674 8563
rect 708 8529 746 8563
rect 780 8529 814 8563
rect 848 8529 882 8563
rect 916 8529 1021 8563
rect -26 8513 1021 8529
rect -1 8491 29 8513
rect 85 8491 115 8513
rect 171 8491 201 8513
rect 257 8491 287 8513
rect 343 8491 373 8513
rect 429 8491 459 8513
rect 515 8491 545 8513
rect 601 8491 631 8513
rect 687 8491 717 8513
rect 773 8491 803 8513
rect 859 8491 889 8513
rect 945 8491 975 8513
rect -1 7455 29 7481
rect 85 7455 115 7481
rect 171 7455 201 7481
rect 257 7455 287 7481
rect -1 7425 287 7455
rect 343 7455 373 7481
rect 429 7455 459 7481
rect 515 7455 545 7481
rect 601 7455 631 7481
rect 343 7425 631 7455
rect 687 7455 717 7481
rect 773 7455 803 7481
rect 859 7455 889 7481
rect 945 7455 975 7481
rect 687 7425 975 7455
rect -918 6944 -852 6960
rect -918 6910 -902 6944
rect -868 6910 -852 6944
rect -918 6887 -852 6910
rect -1134 5856 -1068 5879
rect -1134 5822 -1118 5856
rect -1084 5822 -1068 5856
rect -1134 5806 -1068 5822
rect 203 325 491 355
rect 203 299 233 325
rect 289 299 319 325
rect 375 299 405 325
rect 461 299 491 325
rect 547 325 835 355
rect 547 299 577 325
rect 633 299 663 325
rect 719 299 749 325
rect 805 299 835 325
rect -4234 -773 -4168 -757
rect -4234 -807 -4218 -773
rect -4184 -807 -4168 -773
rect -4234 -830 -4168 -807
rect -3910 -773 -3844 -757
rect -3910 -807 -3894 -773
rect -3860 -807 -3844 -773
rect -3910 -830 -3844 -807
rect 203 -733 233 -711
rect 289 -733 319 -711
rect 375 -733 405 -711
rect 461 -733 491 -711
rect 547 -733 577 -711
rect 633 -733 663 -711
rect 719 -733 749 -711
rect 805 -733 835 -711
rect 178 -749 881 -733
rect 178 -783 194 -749
rect 228 -783 262 -749
rect 296 -783 330 -749
rect 364 -783 398 -749
rect 432 -783 466 -749
rect 500 -783 534 -749
rect 568 -783 606 -749
rect 640 -783 674 -749
rect 708 -783 742 -749
rect 776 -783 810 -749
rect 844 -783 881 -749
rect 178 -803 881 -783
<< polycont >>
rect -6693 17140 -6659 17174
rect -6625 17140 -6591 17174
rect -6557 17140 -6523 17174
rect -6299 17140 -6265 17174
rect -6231 17140 -6197 17174
rect -6163 17140 -6129 17174
rect -5905 17140 -5871 17174
rect -5837 17140 -5803 17174
rect -5769 17140 -5735 17174
rect -5511 17140 -5477 17174
rect -5443 17140 -5409 17174
rect -5375 17140 -5341 17174
rect -6693 16020 -6659 16054
rect -6625 16020 -6591 16054
rect -6557 16020 -6523 16054
rect -6299 16020 -6265 16054
rect -6231 16020 -6197 16054
rect -6163 16020 -6129 16054
rect -5905 16020 -5871 16054
rect -5837 16020 -5803 16054
rect -5769 16020 -5735 16054
rect -5511 16020 -5477 16054
rect -5443 16020 -5409 16054
rect -5375 16020 -5341 16054
rect -1702 8670 -1668 8704
rect -1918 7582 -1884 7616
rect -10 8529 24 8563
rect 58 8529 92 8563
rect 126 8529 160 8563
rect 194 8529 228 8563
rect 262 8529 296 8563
rect 330 8529 364 8563
rect 402 8529 436 8563
rect 470 8529 504 8563
rect 538 8529 572 8563
rect 606 8529 640 8563
rect 674 8529 708 8563
rect 746 8529 780 8563
rect 814 8529 848 8563
rect 882 8529 916 8563
rect -902 6910 -868 6944
rect -1118 5822 -1084 5856
rect -4218 -807 -4184 -773
rect -3894 -807 -3860 -773
rect 194 -783 228 -749
rect 262 -783 296 -749
rect 330 -783 364 -749
rect 398 -783 432 -749
rect 466 -783 500 -749
rect 534 -783 568 -749
rect 606 -783 640 -749
rect 674 -783 708 -749
rect 742 -783 776 -749
rect 810 -783 844 -749
<< npolyres >>
rect -1934 8477 -1760 8543
rect -1934 7639 -1868 8477
rect -1826 7809 -1760 8477
rect -1718 7809 -1652 8647
rect -1826 7743 -1652 7809
rect -1134 6717 -960 6783
rect -1134 5879 -1068 6717
rect -1026 6049 -960 6717
rect -918 6049 -852 6887
rect -1026 5983 -852 6049
rect -4234 -1868 -4168 -830
rect -4126 -1000 -3952 -934
rect -4126 -1868 -4060 -1000
rect -4234 -1934 -4060 -1868
rect -4018 -1868 -3952 -1000
rect -3910 -1868 -3844 -830
rect -4018 -1934 -3844 -1868
<< locali >>
rect -6709 17140 -6697 17174
rect -6659 17140 -6625 17174
rect -6591 17140 -6557 17174
rect -6519 17140 -6507 17174
rect -6315 17140 -6303 17174
rect -6265 17140 -6231 17174
rect -6197 17140 -6163 17174
rect -6125 17140 -6113 17174
rect -5921 17140 -5909 17174
rect -5871 17140 -5837 17174
rect -5803 17140 -5769 17174
rect -5731 17140 -5719 17174
rect -5527 17140 -5515 17174
rect -5477 17140 -5443 17174
rect -5409 17140 -5375 17174
rect -5337 17140 -5325 17174
rect -6711 17090 -6677 17106
rect -6822 17010 -6788 17022
rect -6822 16938 -6788 16954
rect -6822 16866 -6788 16886
rect -6822 16794 -6788 16818
rect -6822 16722 -6788 16750
rect -6822 16650 -6788 16682
rect -6822 16580 -6788 16614
rect -6822 16512 -6788 16544
rect -6822 16444 -6788 16472
rect -6822 16376 -6788 16400
rect -6822 16308 -6788 16328
rect -6822 16240 -6788 16256
rect -6822 16172 -6788 16184
rect -6711 17022 -6677 17048
rect -6711 16954 -6677 16976
rect -6711 16886 -6677 16904
rect -6711 16818 -6677 16832
rect -6711 16750 -6677 16760
rect -6711 16682 -6677 16688
rect -6711 16614 -6677 16616
rect -6711 16578 -6677 16580
rect -6711 16506 -6677 16512
rect -6711 16434 -6677 16444
rect -6711 16362 -6677 16376
rect -6711 16290 -6677 16308
rect -6711 16218 -6677 16240
rect -6711 16146 -6677 16172
rect -6711 16088 -6677 16104
rect -6625 17090 -6591 17106
rect -6625 17022 -6591 17048
rect -6625 16954 -6591 16976
rect -6625 16886 -6591 16904
rect -6625 16818 -6591 16832
rect -6625 16750 -6591 16760
rect -6625 16682 -6591 16688
rect -6625 16614 -6591 16616
rect -6625 16578 -6591 16580
rect -6625 16506 -6591 16512
rect -6625 16434 -6591 16444
rect -6625 16362 -6591 16376
rect -6625 16290 -6591 16308
rect -6625 16218 -6591 16240
rect -6625 16146 -6591 16172
rect -6625 16088 -6591 16104
rect -6539 17090 -6505 17106
rect -6317 17090 -6283 17106
rect -6539 17022 -6505 17048
rect -6539 16954 -6505 16976
rect -6539 16886 -6505 16904
rect -6539 16818 -6505 16832
rect -6539 16750 -6505 16760
rect -6539 16682 -6505 16688
rect -6539 16614 -6505 16616
rect -6539 16578 -6505 16580
rect -6539 16506 -6505 16512
rect -6539 16434 -6505 16444
rect -6539 16362 -6505 16376
rect -6539 16290 -6505 16308
rect -6539 16218 -6505 16240
rect -6539 16146 -6505 16172
rect -6428 17010 -6394 17022
rect -6428 16938 -6394 16954
rect -6428 16866 -6394 16886
rect -6428 16794 -6394 16818
rect -6428 16722 -6394 16750
rect -6428 16650 -6394 16682
rect -6428 16580 -6394 16614
rect -6428 16512 -6394 16544
rect -6428 16444 -6394 16472
rect -6428 16376 -6394 16400
rect -6428 16308 -6394 16328
rect -6428 16240 -6394 16256
rect -6428 16172 -6394 16184
rect -6317 17022 -6283 17048
rect -6317 16954 -6283 16976
rect -6317 16886 -6283 16904
rect -6317 16818 -6283 16832
rect -6317 16750 -6283 16760
rect -6317 16682 -6283 16688
rect -6317 16614 -6283 16616
rect -6317 16578 -6283 16580
rect -6317 16506 -6283 16512
rect -6317 16434 -6283 16444
rect -6317 16362 -6283 16376
rect -6317 16290 -6283 16308
rect -6317 16218 -6283 16240
rect -6317 16146 -6283 16172
rect -6539 16088 -6505 16104
rect -6317 16088 -6283 16104
rect -6231 17090 -6197 17106
rect -6231 17022 -6197 17048
rect -6231 16954 -6197 16976
rect -6231 16886 -6197 16904
rect -6231 16818 -6197 16832
rect -6231 16750 -6197 16760
rect -6231 16682 -6197 16688
rect -6231 16614 -6197 16616
rect -6231 16578 -6197 16580
rect -6231 16506 -6197 16512
rect -6231 16434 -6197 16444
rect -6231 16362 -6197 16376
rect -6231 16290 -6197 16308
rect -6231 16218 -6197 16240
rect -6231 16146 -6197 16172
rect -6231 16088 -6197 16104
rect -6145 17090 -6111 17106
rect -5923 17090 -5889 17106
rect -6145 17022 -6111 17048
rect -6145 16954 -6111 16976
rect -6145 16886 -6111 16904
rect -6145 16818 -6111 16832
rect -6145 16750 -6111 16760
rect -6145 16682 -6111 16688
rect -6145 16614 -6111 16616
rect -6145 16578 -6111 16580
rect -6145 16506 -6111 16512
rect -6145 16434 -6111 16444
rect -6145 16362 -6111 16376
rect -6145 16290 -6111 16308
rect -6145 16218 -6111 16240
rect -6145 16146 -6111 16172
rect -6034 17010 -6000 17022
rect -6034 16938 -6000 16954
rect -6034 16866 -6000 16886
rect -6034 16794 -6000 16818
rect -6034 16722 -6000 16750
rect -6034 16650 -6000 16682
rect -6034 16580 -6000 16614
rect -6034 16512 -6000 16544
rect -6034 16444 -6000 16472
rect -6034 16376 -6000 16400
rect -6034 16308 -6000 16328
rect -6034 16240 -6000 16256
rect -6034 16172 -6000 16184
rect -5923 17022 -5889 17048
rect -5923 16954 -5889 16976
rect -5923 16886 -5889 16904
rect -5923 16818 -5889 16832
rect -5923 16750 -5889 16760
rect -5923 16682 -5889 16688
rect -5923 16614 -5889 16616
rect -5923 16578 -5889 16580
rect -5923 16506 -5889 16512
rect -5923 16434 -5889 16444
rect -5923 16362 -5889 16376
rect -5923 16290 -5889 16308
rect -5923 16218 -5889 16240
rect -5923 16146 -5889 16172
rect -6145 16088 -6111 16104
rect -5923 16088 -5889 16104
rect -5837 17090 -5803 17106
rect -5837 17022 -5803 17048
rect -5837 16954 -5803 16976
rect -5837 16886 -5803 16904
rect -5837 16818 -5803 16832
rect -5837 16750 -5803 16760
rect -5837 16682 -5803 16688
rect -5837 16614 -5803 16616
rect -5837 16578 -5803 16580
rect -5837 16506 -5803 16512
rect -5837 16434 -5803 16444
rect -5837 16362 -5803 16376
rect -5837 16290 -5803 16308
rect -5837 16218 -5803 16240
rect -5837 16146 -5803 16172
rect -5837 16088 -5803 16104
rect -5751 17090 -5717 17106
rect -5529 17090 -5495 17106
rect -5751 17022 -5717 17048
rect -5751 16954 -5717 16976
rect -5751 16886 -5717 16904
rect -5751 16818 -5717 16832
rect -5751 16750 -5717 16760
rect -5751 16682 -5717 16688
rect -5751 16614 -5717 16616
rect -5751 16578 -5717 16580
rect -5751 16506 -5717 16512
rect -5751 16434 -5717 16444
rect -5751 16362 -5717 16376
rect -5751 16290 -5717 16308
rect -5751 16218 -5717 16240
rect -5751 16146 -5717 16172
rect -5640 17010 -5606 17022
rect -5640 16938 -5606 16954
rect -5640 16866 -5606 16886
rect -5640 16794 -5606 16818
rect -5640 16722 -5606 16750
rect -5640 16650 -5606 16682
rect -5640 16580 -5606 16614
rect -5640 16512 -5606 16544
rect -5640 16444 -5606 16472
rect -5640 16376 -5606 16400
rect -5640 16308 -5606 16328
rect -5640 16240 -5606 16256
rect -5640 16172 -5606 16184
rect -5529 17022 -5495 17048
rect -5529 16954 -5495 16976
rect -5529 16886 -5495 16904
rect -5529 16818 -5495 16832
rect -5529 16750 -5495 16760
rect -5529 16682 -5495 16688
rect -5529 16614 -5495 16616
rect -5529 16578 -5495 16580
rect -5529 16506 -5495 16512
rect -5529 16434 -5495 16444
rect -5529 16362 -5495 16376
rect -5529 16290 -5495 16308
rect -5529 16218 -5495 16240
rect -5529 16146 -5495 16172
rect -5751 16088 -5717 16104
rect -5529 16088 -5495 16104
rect -5443 17090 -5409 17106
rect -5443 17022 -5409 17048
rect -5443 16954 -5409 16976
rect -5443 16886 -5409 16904
rect -5443 16818 -5409 16832
rect -5443 16750 -5409 16760
rect -5443 16682 -5409 16688
rect -5443 16614 -5409 16616
rect -5443 16578 -5409 16580
rect -5443 16506 -5409 16512
rect -5443 16434 -5409 16444
rect -5443 16362 -5409 16376
rect -5443 16290 -5409 16308
rect -5443 16218 -5409 16240
rect -5443 16146 -5409 16172
rect -5443 16088 -5409 16104
rect -5357 17090 -5323 17106
rect -5357 17022 -5323 17048
rect -5357 16954 -5323 16976
rect -5357 16886 -5323 16904
rect -5357 16818 -5323 16832
rect -5357 16750 -5323 16760
rect -5357 16682 -5323 16688
rect -5357 16614 -5323 16616
rect -5357 16578 -5323 16580
rect -5357 16506 -5323 16512
rect -5357 16434 -5323 16444
rect -5357 16362 -5323 16376
rect -5357 16290 -5323 16308
rect -5357 16218 -5323 16240
rect -5357 16146 -5323 16172
rect -5246 17010 -5212 17022
rect -5246 16938 -5212 16954
rect -5246 16866 -5212 16886
rect -5246 16794 -5212 16818
rect -5246 16722 -5212 16750
rect -5246 16650 -5212 16682
rect -5246 16580 -5212 16614
rect -5246 16512 -5212 16544
rect -5246 16444 -5212 16472
rect -5246 16376 -5212 16400
rect -5246 16308 -5212 16328
rect -5246 16240 -5212 16256
rect -5246 16172 -5212 16184
rect -5357 16088 -5323 16104
rect -6709 16020 -6697 16054
rect -6659 16020 -6625 16054
rect -6591 16020 -6557 16054
rect -6519 16020 -6507 16054
rect -6315 16020 -6303 16054
rect -6265 16020 -6231 16054
rect -6197 16020 -6163 16054
rect -6125 16020 -6113 16054
rect -5921 16020 -5909 16054
rect -5871 16020 -5837 16054
rect -5803 16020 -5769 16054
rect -5731 16020 -5719 16054
rect -5527 16020 -5515 16054
rect -5477 16020 -5443 16054
rect -5409 16020 -5375 16054
rect -5337 16020 -5325 16054
rect -2064 8816 -1968 8850
rect -1618 8816 -1450 8850
rect -2064 8754 -2030 8816
rect -1556 8754 -1450 8816
rect -2064 7470 -2030 7532
rect -1560 7532 -1556 8500
rect -1522 8500 -1450 8754
rect -26 8529 -10 8563
rect 24 8529 54 8563
rect 92 8529 126 8563
rect 160 8529 194 8563
rect 232 8529 262 8563
rect 296 8529 330 8563
rect 364 8529 398 8563
rect 436 8529 470 8563
rect 504 8529 538 8563
rect 576 8529 606 8563
rect 640 8529 674 8563
rect 708 8529 742 8563
rect 780 8529 814 8563
rect 848 8529 882 8563
rect 920 8529 1020 8563
rect -1522 8480 -1400 8500
rect -1560 7470 -1540 7532
rect -2064 7436 -1968 7470
rect -1618 7436 -1540 7470
rect -2050 7360 -1540 7436
rect -1420 7360 -1400 8480
rect -46 8479 -12 8495
rect -2050 7350 -1400 7360
rect -1560 7340 -1400 7350
rect -184 8454 -134 8470
rect -184 8420 -174 8454
rect -140 8420 -134 8454
rect -184 8384 -134 8420
rect -184 8340 -174 8384
rect -140 8340 -134 8384
rect -184 8314 -134 8340
rect -184 8260 -174 8314
rect -140 8260 -134 8314
rect -184 8244 -134 8260
rect -184 8180 -174 8244
rect -140 8180 -134 8244
rect -184 8174 -134 8180
rect -184 8140 -174 8174
rect -140 8140 -134 8174
rect -184 8134 -134 8140
rect -184 8070 -174 8134
rect -140 8070 -134 8134
rect -184 8054 -134 8070
rect -184 8000 -174 8054
rect -140 8000 -134 8054
rect -184 7974 -134 8000
rect -184 7930 -174 7974
rect -140 7930 -134 7974
rect -184 7894 -134 7930
rect -184 7860 -174 7894
rect -140 7860 -134 7894
rect -184 7824 -134 7860
rect -184 7780 -174 7824
rect -140 7780 -134 7824
rect -184 7754 -134 7780
rect -184 7700 -174 7754
rect -140 7700 -134 7754
rect -184 7684 -134 7700
rect -184 7620 -174 7684
rect -140 7620 -134 7684
rect -184 7614 -134 7620
rect -184 7580 -174 7614
rect -140 7580 -134 7614
rect -184 7574 -134 7580
rect -184 7510 -174 7574
rect -140 7510 -134 7574
rect -184 7494 -134 7510
rect -184 7440 -174 7494
rect -140 7440 -134 7494
rect -46 8411 -12 8437
rect -46 8343 -12 8365
rect -46 8275 -12 8293
rect -46 8207 -12 8221
rect -46 8139 -12 8149
rect -46 8071 -12 8077
rect -46 8003 -12 8005
rect -46 7967 -12 7969
rect -46 7895 -12 7901
rect -46 7823 -12 7833
rect -46 7751 -12 7765
rect -46 7679 -12 7697
rect -46 7607 -12 7629
rect -46 7535 -12 7561
rect -46 7477 -12 7493
rect 40 8479 74 8495
rect 40 8411 74 8437
rect 40 8343 74 8365
rect 40 8275 74 8293
rect 40 8207 74 8221
rect 40 8139 74 8149
rect 40 8071 74 8077
rect 40 8003 74 8005
rect 40 7967 74 7969
rect 40 7895 74 7901
rect 40 7823 74 7833
rect 40 7751 74 7765
rect 40 7679 74 7697
rect 40 7607 74 7629
rect 40 7535 74 7561
rect 40 7477 74 7493
rect 126 8479 160 8495
rect 126 8411 160 8437
rect 126 8343 160 8365
rect 126 8275 160 8293
rect 126 8207 160 8221
rect 126 8139 160 8149
rect 126 8071 160 8077
rect 126 8003 160 8005
rect 126 7967 160 7969
rect 126 7895 160 7901
rect 126 7823 160 7833
rect 126 7751 160 7765
rect 126 7679 160 7697
rect 126 7607 160 7629
rect 126 7535 160 7561
rect 126 7477 160 7493
rect 212 8479 246 8495
rect 212 8411 246 8437
rect 212 8343 246 8365
rect 212 8275 246 8293
rect 212 8207 246 8221
rect 212 8139 246 8149
rect 212 8071 246 8077
rect 212 8003 246 8005
rect 212 7967 246 7969
rect 212 7895 246 7901
rect 212 7823 246 7833
rect 212 7751 246 7765
rect 212 7679 246 7697
rect 212 7607 246 7629
rect 212 7535 246 7561
rect 212 7477 246 7493
rect 298 8479 332 8495
rect 298 8411 332 8437
rect 298 8343 332 8365
rect 298 8275 332 8293
rect 298 8207 332 8221
rect 298 8139 332 8149
rect 298 8071 332 8077
rect 298 8003 332 8005
rect 298 7967 332 7969
rect 298 7895 332 7901
rect 298 7823 332 7833
rect 298 7751 332 7765
rect 298 7679 332 7697
rect 298 7607 332 7629
rect 298 7535 332 7561
rect 298 7477 332 7493
rect 384 8479 418 8495
rect 384 8411 418 8437
rect 384 8343 418 8365
rect 384 8275 418 8293
rect 384 8207 418 8221
rect 384 8139 418 8149
rect 384 8071 418 8077
rect 384 8003 418 8005
rect 384 7967 418 7969
rect 384 7895 418 7901
rect 384 7823 418 7833
rect 384 7751 418 7765
rect 384 7679 418 7697
rect 384 7607 418 7629
rect 384 7535 418 7561
rect 384 7477 418 7493
rect 470 8479 504 8495
rect 470 8411 504 8437
rect 470 8343 504 8365
rect 470 8275 504 8293
rect 470 8207 504 8221
rect 470 8139 504 8149
rect 470 8071 504 8077
rect 470 8003 504 8005
rect 470 7967 504 7969
rect 470 7895 504 7901
rect 470 7823 504 7833
rect 470 7751 504 7765
rect 470 7679 504 7697
rect 470 7607 504 7629
rect 470 7535 504 7561
rect 470 7477 504 7493
rect 556 8479 590 8495
rect 556 8411 590 8437
rect 556 8343 590 8365
rect 556 8275 590 8293
rect 556 8207 590 8221
rect 556 8139 590 8149
rect 556 8071 590 8077
rect 556 8003 590 8005
rect 556 7967 590 7969
rect 556 7895 590 7901
rect 556 7823 590 7833
rect 556 7751 590 7765
rect 556 7679 590 7697
rect 556 7607 590 7629
rect 556 7535 590 7561
rect 556 7477 590 7493
rect 642 8479 676 8495
rect 642 8411 676 8437
rect 642 8343 676 8365
rect 642 8275 676 8293
rect 642 8207 676 8221
rect 642 8139 676 8149
rect 642 8071 676 8077
rect 642 8003 676 8005
rect 642 7967 676 7969
rect 642 7895 676 7901
rect 642 7823 676 7833
rect 642 7751 676 7765
rect 642 7679 676 7697
rect 642 7607 676 7629
rect 642 7535 676 7561
rect 642 7477 676 7493
rect 728 8479 762 8495
rect 728 8411 762 8437
rect 728 8343 762 8365
rect 728 8275 762 8293
rect 728 8207 762 8221
rect 728 8139 762 8149
rect 728 8071 762 8077
rect 728 8003 762 8005
rect 728 7967 762 7969
rect 728 7895 762 7901
rect 728 7823 762 7833
rect 728 7751 762 7765
rect 728 7679 762 7697
rect 728 7607 762 7629
rect 728 7535 762 7561
rect 728 7477 762 7493
rect 814 8479 848 8495
rect 814 8411 848 8437
rect 814 8343 848 8365
rect 814 8275 848 8293
rect 814 8207 848 8221
rect 814 8139 848 8149
rect 814 8071 848 8077
rect 814 8003 848 8005
rect 814 7967 848 7969
rect 814 7895 848 7901
rect 814 7823 848 7833
rect 814 7751 848 7765
rect 814 7679 848 7697
rect 814 7607 848 7629
rect 814 7535 848 7561
rect 814 7477 848 7493
rect 900 8479 934 8495
rect 900 8411 934 8437
rect 900 8343 934 8365
rect 900 8275 934 8293
rect 900 8207 934 8221
rect 900 8139 934 8149
rect 900 8071 934 8077
rect 900 8003 934 8005
rect 900 7967 934 7969
rect 900 7895 934 7901
rect 900 7823 934 7833
rect 900 7751 934 7765
rect 900 7679 934 7697
rect 900 7607 934 7629
rect 900 7535 934 7561
rect 900 7477 934 7493
rect 986 8479 1020 8495
rect 986 8411 1020 8437
rect 986 8343 1020 8365
rect 986 8275 1020 8293
rect 986 8207 1020 8221
rect 986 8139 1020 8149
rect 986 8071 1020 8077
rect 986 8003 1020 8005
rect 986 7967 1020 7969
rect 986 7895 1020 7901
rect 986 7823 1020 7833
rect 986 7751 1020 7765
rect 986 7679 1020 7697
rect 986 7607 1020 7629
rect 986 7535 1020 7561
rect 986 7477 1020 7493
rect 1106 8454 1166 8470
rect 1106 8420 1116 8454
rect 1150 8420 1166 8454
rect 1106 8384 1166 8420
rect 1106 8340 1116 8384
rect 1150 8340 1166 8384
rect 1106 8314 1166 8340
rect 1106 8260 1116 8314
rect 1150 8260 1166 8314
rect 1106 8244 1166 8260
rect 1106 8180 1116 8244
rect 1150 8180 1166 8244
rect 1106 8174 1166 8180
rect 1106 8140 1116 8174
rect 1150 8140 1166 8174
rect 1106 8134 1166 8140
rect 1106 8070 1116 8134
rect 1150 8070 1166 8134
rect 1106 8054 1166 8070
rect 1106 8000 1116 8054
rect 1150 8000 1166 8054
rect 1106 7974 1166 8000
rect 1106 7930 1116 7974
rect 1150 7930 1166 7974
rect 1106 7894 1166 7930
rect 1106 7860 1116 7894
rect 1150 7860 1166 7894
rect 1106 7824 1166 7860
rect 1106 7780 1116 7824
rect 1150 7780 1166 7824
rect 1106 7754 1166 7780
rect 1106 7700 1116 7754
rect 1150 7700 1166 7754
rect 1106 7684 1166 7700
rect 1106 7620 1116 7684
rect 1150 7620 1166 7684
rect 1106 7614 1166 7620
rect 1106 7580 1116 7614
rect 1150 7580 1166 7614
rect 1106 7574 1166 7580
rect 1106 7510 1116 7574
rect 1150 7510 1166 7574
rect 1106 7494 1166 7510
rect -184 7400 -134 7440
rect 1106 7440 1116 7494
rect 1150 7440 1166 7494
rect 1106 7400 1166 7440
rect -184 7384 1166 7400
rect -184 7350 -94 7384
rect -60 7350 -24 7384
rect 10 7350 46 7384
rect 80 7350 116 7384
rect 150 7350 186 7384
rect 220 7350 256 7384
rect 290 7350 326 7384
rect 360 7350 396 7384
rect 430 7350 466 7384
rect 500 7350 536 7384
rect 570 7350 606 7384
rect 640 7350 676 7384
rect 710 7350 746 7384
rect 780 7350 816 7384
rect 850 7350 886 7384
rect 920 7350 956 7384
rect 990 7350 1026 7384
rect 1060 7350 1166 7384
rect -184 7340 1166 7350
rect -1264 7080 -1168 7090
rect -1400 7060 -1168 7080
rect -1400 5700 -1380 7060
rect -1260 7056 -1168 7060
rect -818 7056 -722 7090
rect -1260 6994 -1230 7056
rect -756 6994 -722 7056
rect -1260 5710 -1230 5772
rect -756 5710 -722 5772
rect -1260 5700 -1168 5710
rect -1400 5680 -1168 5700
rect -1264 5676 -1168 5680
rect -818 5676 -722 5710
rect 20 430 1017 440
rect 20 390 50 430
rect 990 390 1017 430
rect 20 380 1017 390
rect 20 340 70 380
rect 20 286 30 340
rect 64 286 70 340
rect 957 340 1017 380
rect 20 270 70 286
rect 20 206 30 270
rect 64 206 70 270
rect 20 200 70 206
rect 20 166 30 200
rect 64 166 70 200
rect 20 160 70 166
rect 20 96 30 160
rect 64 96 70 160
rect 20 80 70 96
rect 20 26 30 80
rect 64 26 70 80
rect 20 0 70 26
rect 20 -44 30 0
rect 64 -44 70 0
rect 20 -80 70 -44
rect 20 -114 30 -80
rect 64 -114 70 -80
rect 20 -150 70 -114
rect 20 -194 30 -150
rect 64 -194 70 -150
rect 20 -220 70 -194
rect 20 -274 30 -220
rect 64 -274 70 -220
rect 20 -290 70 -274
rect 20 -354 30 -290
rect 64 -354 70 -290
rect 20 -360 70 -354
rect 20 -394 30 -360
rect 64 -394 70 -360
rect 20 -400 70 -394
rect 20 -464 30 -400
rect 64 -464 70 -400
rect 20 -480 70 -464
rect 20 -534 30 -480
rect 64 -534 70 -480
rect 20 -560 70 -534
rect 20 -604 30 -560
rect 64 -604 70 -560
rect -4560 -630 -4400 -620
rect -4364 -630 -4268 -626
rect -4560 -640 -4268 -630
rect -4560 -2220 -4540 -640
rect -4420 -660 -4268 -640
rect -3810 -660 -3714 -626
rect -4420 -722 -4330 -660
rect -4420 -1968 -4364 -722
rect -3748 -722 -3714 -660
rect 20 -640 70 -604
rect 20 -674 30 -640
rect 64 -674 70 -640
rect 20 -690 70 -674
rect 158 287 192 303
rect 158 219 192 245
rect 158 151 192 173
rect 158 83 192 101
rect 158 15 192 29
rect 158 -53 192 -43
rect 158 -121 192 -115
rect 158 -189 192 -187
rect 158 -225 192 -223
rect 158 -297 192 -291
rect 158 -369 192 -359
rect 158 -441 192 -427
rect 158 -513 192 -495
rect 158 -585 192 -563
rect 158 -657 192 -631
rect 158 -715 192 -699
rect 244 287 278 303
rect 244 219 278 245
rect 244 151 278 173
rect 244 83 278 101
rect 244 15 278 29
rect 244 -53 278 -43
rect 244 -121 278 -115
rect 244 -189 278 -187
rect 244 -225 278 -223
rect 244 -297 278 -291
rect 244 -369 278 -359
rect 244 -441 278 -427
rect 244 -513 278 -495
rect 244 -585 278 -563
rect 244 -657 278 -631
rect 244 -715 278 -699
rect 330 287 364 303
rect 330 219 364 245
rect 330 151 364 173
rect 330 83 364 101
rect 330 15 364 29
rect 330 -53 364 -43
rect 330 -121 364 -115
rect 330 -189 364 -187
rect 330 -225 364 -223
rect 330 -297 364 -291
rect 330 -369 364 -359
rect 330 -441 364 -427
rect 330 -513 364 -495
rect 330 -585 364 -563
rect 330 -657 364 -631
rect 330 -715 364 -699
rect 416 287 450 303
rect 416 219 450 245
rect 416 151 450 173
rect 416 83 450 101
rect 416 15 450 29
rect 416 -53 450 -43
rect 416 -121 450 -115
rect 416 -189 450 -187
rect 416 -225 450 -223
rect 416 -297 450 -291
rect 416 -369 450 -359
rect 416 -441 450 -427
rect 416 -513 450 -495
rect 416 -585 450 -563
rect 416 -657 450 -631
rect 416 -715 450 -699
rect 502 287 536 303
rect 502 219 536 245
rect 502 151 536 173
rect 502 83 536 101
rect 502 15 536 29
rect 502 -53 536 -43
rect 502 -121 536 -115
rect 502 -189 536 -187
rect 502 -225 536 -223
rect 502 -297 536 -291
rect 502 -369 536 -359
rect 502 -441 536 -427
rect 502 -513 536 -495
rect 502 -585 536 -563
rect 502 -657 536 -631
rect 502 -715 536 -699
rect 588 287 622 303
rect 588 219 622 245
rect 588 151 622 173
rect 588 83 622 101
rect 588 15 622 29
rect 588 -53 622 -43
rect 588 -121 622 -115
rect 588 -189 622 -187
rect 588 -225 622 -223
rect 588 -297 622 -291
rect 588 -369 622 -359
rect 588 -441 622 -427
rect 588 -513 622 -495
rect 588 -585 622 -563
rect 588 -657 622 -631
rect 588 -715 622 -699
rect 674 287 708 303
rect 674 219 708 245
rect 674 151 708 173
rect 674 83 708 101
rect 674 15 708 29
rect 674 -53 708 -43
rect 674 -121 708 -115
rect 674 -189 708 -187
rect 674 -225 708 -223
rect 674 -297 708 -291
rect 674 -369 708 -359
rect 674 -441 708 -427
rect 674 -513 708 -495
rect 674 -585 708 -563
rect 674 -657 708 -631
rect 674 -715 708 -699
rect 760 287 794 303
rect 760 219 794 245
rect 760 151 794 173
rect 760 83 794 101
rect 760 15 794 29
rect 760 -53 794 -43
rect 760 -121 794 -115
rect 760 -189 794 -187
rect 760 -225 794 -223
rect 760 -297 794 -291
rect 760 -369 794 -359
rect 760 -441 794 -427
rect 760 -513 794 -495
rect 760 -585 794 -563
rect 760 -657 794 -631
rect 760 -715 794 -699
rect 846 287 880 303
rect 846 219 880 245
rect 846 151 880 173
rect 846 83 880 101
rect 846 15 880 29
rect 846 -53 880 -43
rect 846 -121 880 -115
rect 846 -189 880 -187
rect 846 -225 880 -223
rect 846 -297 880 -291
rect 846 -369 880 -359
rect 846 -441 880 -427
rect 846 -513 880 -495
rect 846 -585 880 -563
rect 846 -657 880 -631
rect 957 286 967 340
rect 1001 286 1017 340
rect 957 270 1017 286
rect 957 206 967 270
rect 1001 206 1017 270
rect 957 200 1017 206
rect 957 166 967 200
rect 1001 166 1017 200
rect 957 160 1017 166
rect 957 96 967 160
rect 1001 96 1017 160
rect 957 80 1017 96
rect 957 26 967 80
rect 1001 26 1017 80
rect 957 0 1017 26
rect 957 -44 967 0
rect 1001 -44 1017 0
rect 957 -80 1017 -44
rect 957 -114 967 -80
rect 1001 -114 1017 -80
rect 957 -150 1017 -114
rect 957 -194 967 -150
rect 1001 -194 1017 -150
rect 957 -220 1017 -194
rect 957 -274 967 -220
rect 1001 -274 1017 -220
rect 957 -290 1017 -274
rect 957 -354 967 -290
rect 1001 -354 1017 -290
rect 957 -360 1017 -354
rect 957 -394 967 -360
rect 1001 -394 1017 -360
rect 957 -400 1017 -394
rect 957 -464 967 -400
rect 1001 -464 1017 -400
rect 957 -480 1017 -464
rect 957 -534 967 -480
rect 1001 -534 1017 -480
rect 957 -560 1017 -534
rect 957 -604 967 -560
rect 1001 -604 1017 -560
rect 957 -640 1017 -604
rect 957 -674 967 -640
rect 1001 -674 1017 -640
rect 957 -690 1017 -674
rect 846 -715 880 -699
rect -4420 -2030 -4330 -1968
rect 178 -783 194 -749
rect 228 -783 258 -749
rect 296 -783 330 -749
rect 364 -783 398 -749
rect 436 -783 466 -749
rect 500 -783 534 -749
rect 568 -783 602 -749
rect 640 -783 674 -749
rect 708 -783 742 -749
rect 780 -783 810 -749
rect 844 -783 871 -749
rect -3748 -2030 -3714 -1968
rect -4420 -2060 -4268 -2030
rect -3810 -2060 -3714 -2030
rect -3740 -2064 -3714 -2060
rect -3740 -2220 -3720 -2064
rect -4560 -2240 -3720 -2220
<< viali >>
rect -6697 17140 -6693 17174
rect -6693 17140 -6663 17174
rect -6625 17140 -6591 17174
rect -6553 17140 -6523 17174
rect -6523 17140 -6519 17174
rect -6303 17140 -6299 17174
rect -6299 17140 -6269 17174
rect -6231 17140 -6197 17174
rect -6159 17140 -6129 17174
rect -6129 17140 -6125 17174
rect -5909 17140 -5905 17174
rect -5905 17140 -5875 17174
rect -5837 17140 -5803 17174
rect -5765 17140 -5735 17174
rect -5735 17140 -5731 17174
rect -5515 17140 -5511 17174
rect -5511 17140 -5481 17174
rect -5443 17140 -5409 17174
rect -5371 17140 -5341 17174
rect -5341 17140 -5337 17174
rect -6822 17056 -6788 17082
rect -6822 17048 -6788 17056
rect -6822 16988 -6788 17010
rect -6822 16976 -6788 16988
rect -6822 16920 -6788 16938
rect -6822 16904 -6788 16920
rect -6822 16852 -6788 16866
rect -6822 16832 -6788 16852
rect -6822 16784 -6788 16794
rect -6822 16760 -6788 16784
rect -6822 16716 -6788 16722
rect -6822 16688 -6788 16716
rect -6822 16648 -6788 16650
rect -6822 16616 -6788 16648
rect -6822 16546 -6788 16578
rect -6822 16544 -6788 16546
rect -6822 16478 -6788 16506
rect -6822 16472 -6788 16478
rect -6822 16410 -6788 16434
rect -6822 16400 -6788 16410
rect -6822 16342 -6788 16362
rect -6822 16328 -6788 16342
rect -6822 16274 -6788 16290
rect -6822 16256 -6788 16274
rect -6822 16206 -6788 16218
rect -6822 16184 -6788 16206
rect -6822 16138 -6788 16146
rect -6822 16112 -6788 16138
rect -6711 17056 -6677 17082
rect -6711 17048 -6677 17056
rect -6711 16988 -6677 17010
rect -6711 16976 -6677 16988
rect -6711 16920 -6677 16938
rect -6711 16904 -6677 16920
rect -6711 16852 -6677 16866
rect -6711 16832 -6677 16852
rect -6711 16784 -6677 16794
rect -6711 16760 -6677 16784
rect -6711 16716 -6677 16722
rect -6711 16688 -6677 16716
rect -6711 16648 -6677 16650
rect -6711 16616 -6677 16648
rect -6711 16546 -6677 16578
rect -6711 16544 -6677 16546
rect -6711 16478 -6677 16506
rect -6711 16472 -6677 16478
rect -6711 16410 -6677 16434
rect -6711 16400 -6677 16410
rect -6711 16342 -6677 16362
rect -6711 16328 -6677 16342
rect -6711 16274 -6677 16290
rect -6711 16256 -6677 16274
rect -6711 16206 -6677 16218
rect -6711 16184 -6677 16206
rect -6711 16138 -6677 16146
rect -6711 16112 -6677 16138
rect -6625 17056 -6591 17082
rect -6625 17048 -6591 17056
rect -6625 16988 -6591 17010
rect -6625 16976 -6591 16988
rect -6625 16920 -6591 16938
rect -6625 16904 -6591 16920
rect -6625 16852 -6591 16866
rect -6625 16832 -6591 16852
rect -6625 16784 -6591 16794
rect -6625 16760 -6591 16784
rect -6625 16716 -6591 16722
rect -6625 16688 -6591 16716
rect -6625 16648 -6591 16650
rect -6625 16616 -6591 16648
rect -6625 16546 -6591 16578
rect -6625 16544 -6591 16546
rect -6625 16478 -6591 16506
rect -6625 16472 -6591 16478
rect -6625 16410 -6591 16434
rect -6625 16400 -6591 16410
rect -6625 16342 -6591 16362
rect -6625 16328 -6591 16342
rect -6625 16274 -6591 16290
rect -6625 16256 -6591 16274
rect -6625 16206 -6591 16218
rect -6625 16184 -6591 16206
rect -6625 16138 -6591 16146
rect -6625 16112 -6591 16138
rect -6539 17056 -6505 17082
rect -6539 17048 -6505 17056
rect -6539 16988 -6505 17010
rect -6539 16976 -6505 16988
rect -6539 16920 -6505 16938
rect -6539 16904 -6505 16920
rect -6539 16852 -6505 16866
rect -6539 16832 -6505 16852
rect -6539 16784 -6505 16794
rect -6539 16760 -6505 16784
rect -6539 16716 -6505 16722
rect -6539 16688 -6505 16716
rect -6539 16648 -6505 16650
rect -6539 16616 -6505 16648
rect -6539 16546 -6505 16578
rect -6539 16544 -6505 16546
rect -6539 16478 -6505 16506
rect -6539 16472 -6505 16478
rect -6539 16410 -6505 16434
rect -6539 16400 -6505 16410
rect -6539 16342 -6505 16362
rect -6539 16328 -6505 16342
rect -6539 16274 -6505 16290
rect -6539 16256 -6505 16274
rect -6539 16206 -6505 16218
rect -6539 16184 -6505 16206
rect -6539 16138 -6505 16146
rect -6539 16112 -6505 16138
rect -6428 17056 -6394 17082
rect -6428 17048 -6394 17056
rect -6428 16988 -6394 17010
rect -6428 16976 -6394 16988
rect -6428 16920 -6394 16938
rect -6428 16904 -6394 16920
rect -6428 16852 -6394 16866
rect -6428 16832 -6394 16852
rect -6428 16784 -6394 16794
rect -6428 16760 -6394 16784
rect -6428 16716 -6394 16722
rect -6428 16688 -6394 16716
rect -6428 16648 -6394 16650
rect -6428 16616 -6394 16648
rect -6428 16546 -6394 16578
rect -6428 16544 -6394 16546
rect -6428 16478 -6394 16506
rect -6428 16472 -6394 16478
rect -6428 16410 -6394 16434
rect -6428 16400 -6394 16410
rect -6428 16342 -6394 16362
rect -6428 16328 -6394 16342
rect -6428 16274 -6394 16290
rect -6428 16256 -6394 16274
rect -6428 16206 -6394 16218
rect -6428 16184 -6394 16206
rect -6428 16138 -6394 16146
rect -6428 16112 -6394 16138
rect -6317 17056 -6283 17082
rect -6317 17048 -6283 17056
rect -6317 16988 -6283 17010
rect -6317 16976 -6283 16988
rect -6317 16920 -6283 16938
rect -6317 16904 -6283 16920
rect -6317 16852 -6283 16866
rect -6317 16832 -6283 16852
rect -6317 16784 -6283 16794
rect -6317 16760 -6283 16784
rect -6317 16716 -6283 16722
rect -6317 16688 -6283 16716
rect -6317 16648 -6283 16650
rect -6317 16616 -6283 16648
rect -6317 16546 -6283 16578
rect -6317 16544 -6283 16546
rect -6317 16478 -6283 16506
rect -6317 16472 -6283 16478
rect -6317 16410 -6283 16434
rect -6317 16400 -6283 16410
rect -6317 16342 -6283 16362
rect -6317 16328 -6283 16342
rect -6317 16274 -6283 16290
rect -6317 16256 -6283 16274
rect -6317 16206 -6283 16218
rect -6317 16184 -6283 16206
rect -6317 16138 -6283 16146
rect -6317 16112 -6283 16138
rect -6231 17056 -6197 17082
rect -6231 17048 -6197 17056
rect -6231 16988 -6197 17010
rect -6231 16976 -6197 16988
rect -6231 16920 -6197 16938
rect -6231 16904 -6197 16920
rect -6231 16852 -6197 16866
rect -6231 16832 -6197 16852
rect -6231 16784 -6197 16794
rect -6231 16760 -6197 16784
rect -6231 16716 -6197 16722
rect -6231 16688 -6197 16716
rect -6231 16648 -6197 16650
rect -6231 16616 -6197 16648
rect -6231 16546 -6197 16578
rect -6231 16544 -6197 16546
rect -6231 16478 -6197 16506
rect -6231 16472 -6197 16478
rect -6231 16410 -6197 16434
rect -6231 16400 -6197 16410
rect -6231 16342 -6197 16362
rect -6231 16328 -6197 16342
rect -6231 16274 -6197 16290
rect -6231 16256 -6197 16274
rect -6231 16206 -6197 16218
rect -6231 16184 -6197 16206
rect -6231 16138 -6197 16146
rect -6231 16112 -6197 16138
rect -6145 17056 -6111 17082
rect -6145 17048 -6111 17056
rect -6145 16988 -6111 17010
rect -6145 16976 -6111 16988
rect -6145 16920 -6111 16938
rect -6145 16904 -6111 16920
rect -6145 16852 -6111 16866
rect -6145 16832 -6111 16852
rect -6145 16784 -6111 16794
rect -6145 16760 -6111 16784
rect -6145 16716 -6111 16722
rect -6145 16688 -6111 16716
rect -6145 16648 -6111 16650
rect -6145 16616 -6111 16648
rect -6145 16546 -6111 16578
rect -6145 16544 -6111 16546
rect -6145 16478 -6111 16506
rect -6145 16472 -6111 16478
rect -6145 16410 -6111 16434
rect -6145 16400 -6111 16410
rect -6145 16342 -6111 16362
rect -6145 16328 -6111 16342
rect -6145 16274 -6111 16290
rect -6145 16256 -6111 16274
rect -6145 16206 -6111 16218
rect -6145 16184 -6111 16206
rect -6145 16138 -6111 16146
rect -6145 16112 -6111 16138
rect -6034 17056 -6000 17082
rect -6034 17048 -6000 17056
rect -6034 16988 -6000 17010
rect -6034 16976 -6000 16988
rect -6034 16920 -6000 16938
rect -6034 16904 -6000 16920
rect -6034 16852 -6000 16866
rect -6034 16832 -6000 16852
rect -6034 16784 -6000 16794
rect -6034 16760 -6000 16784
rect -6034 16716 -6000 16722
rect -6034 16688 -6000 16716
rect -6034 16648 -6000 16650
rect -6034 16616 -6000 16648
rect -6034 16546 -6000 16578
rect -6034 16544 -6000 16546
rect -6034 16478 -6000 16506
rect -6034 16472 -6000 16478
rect -6034 16410 -6000 16434
rect -6034 16400 -6000 16410
rect -6034 16342 -6000 16362
rect -6034 16328 -6000 16342
rect -6034 16274 -6000 16290
rect -6034 16256 -6000 16274
rect -6034 16206 -6000 16218
rect -6034 16184 -6000 16206
rect -6034 16138 -6000 16146
rect -6034 16112 -6000 16138
rect -5923 17056 -5889 17082
rect -5923 17048 -5889 17056
rect -5923 16988 -5889 17010
rect -5923 16976 -5889 16988
rect -5923 16920 -5889 16938
rect -5923 16904 -5889 16920
rect -5923 16852 -5889 16866
rect -5923 16832 -5889 16852
rect -5923 16784 -5889 16794
rect -5923 16760 -5889 16784
rect -5923 16716 -5889 16722
rect -5923 16688 -5889 16716
rect -5923 16648 -5889 16650
rect -5923 16616 -5889 16648
rect -5923 16546 -5889 16578
rect -5923 16544 -5889 16546
rect -5923 16478 -5889 16506
rect -5923 16472 -5889 16478
rect -5923 16410 -5889 16434
rect -5923 16400 -5889 16410
rect -5923 16342 -5889 16362
rect -5923 16328 -5889 16342
rect -5923 16274 -5889 16290
rect -5923 16256 -5889 16274
rect -5923 16206 -5889 16218
rect -5923 16184 -5889 16206
rect -5923 16138 -5889 16146
rect -5923 16112 -5889 16138
rect -5837 17056 -5803 17082
rect -5837 17048 -5803 17056
rect -5837 16988 -5803 17010
rect -5837 16976 -5803 16988
rect -5837 16920 -5803 16938
rect -5837 16904 -5803 16920
rect -5837 16852 -5803 16866
rect -5837 16832 -5803 16852
rect -5837 16784 -5803 16794
rect -5837 16760 -5803 16784
rect -5837 16716 -5803 16722
rect -5837 16688 -5803 16716
rect -5837 16648 -5803 16650
rect -5837 16616 -5803 16648
rect -5837 16546 -5803 16578
rect -5837 16544 -5803 16546
rect -5837 16478 -5803 16506
rect -5837 16472 -5803 16478
rect -5837 16410 -5803 16434
rect -5837 16400 -5803 16410
rect -5837 16342 -5803 16362
rect -5837 16328 -5803 16342
rect -5837 16274 -5803 16290
rect -5837 16256 -5803 16274
rect -5837 16206 -5803 16218
rect -5837 16184 -5803 16206
rect -5837 16138 -5803 16146
rect -5837 16112 -5803 16138
rect -5751 17056 -5717 17082
rect -5751 17048 -5717 17056
rect -5751 16988 -5717 17010
rect -5751 16976 -5717 16988
rect -5751 16920 -5717 16938
rect -5751 16904 -5717 16920
rect -5751 16852 -5717 16866
rect -5751 16832 -5717 16852
rect -5751 16784 -5717 16794
rect -5751 16760 -5717 16784
rect -5751 16716 -5717 16722
rect -5751 16688 -5717 16716
rect -5751 16648 -5717 16650
rect -5751 16616 -5717 16648
rect -5751 16546 -5717 16578
rect -5751 16544 -5717 16546
rect -5751 16478 -5717 16506
rect -5751 16472 -5717 16478
rect -5751 16410 -5717 16434
rect -5751 16400 -5717 16410
rect -5751 16342 -5717 16362
rect -5751 16328 -5717 16342
rect -5751 16274 -5717 16290
rect -5751 16256 -5717 16274
rect -5751 16206 -5717 16218
rect -5751 16184 -5717 16206
rect -5751 16138 -5717 16146
rect -5751 16112 -5717 16138
rect -5640 17056 -5606 17082
rect -5640 17048 -5606 17056
rect -5640 16988 -5606 17010
rect -5640 16976 -5606 16988
rect -5640 16920 -5606 16938
rect -5640 16904 -5606 16920
rect -5640 16852 -5606 16866
rect -5640 16832 -5606 16852
rect -5640 16784 -5606 16794
rect -5640 16760 -5606 16784
rect -5640 16716 -5606 16722
rect -5640 16688 -5606 16716
rect -5640 16648 -5606 16650
rect -5640 16616 -5606 16648
rect -5640 16546 -5606 16578
rect -5640 16544 -5606 16546
rect -5640 16478 -5606 16506
rect -5640 16472 -5606 16478
rect -5640 16410 -5606 16434
rect -5640 16400 -5606 16410
rect -5640 16342 -5606 16362
rect -5640 16328 -5606 16342
rect -5640 16274 -5606 16290
rect -5640 16256 -5606 16274
rect -5640 16206 -5606 16218
rect -5640 16184 -5606 16206
rect -5640 16138 -5606 16146
rect -5640 16112 -5606 16138
rect -5529 17056 -5495 17082
rect -5529 17048 -5495 17056
rect -5529 16988 -5495 17010
rect -5529 16976 -5495 16988
rect -5529 16920 -5495 16938
rect -5529 16904 -5495 16920
rect -5529 16852 -5495 16866
rect -5529 16832 -5495 16852
rect -5529 16784 -5495 16794
rect -5529 16760 -5495 16784
rect -5529 16716 -5495 16722
rect -5529 16688 -5495 16716
rect -5529 16648 -5495 16650
rect -5529 16616 -5495 16648
rect -5529 16546 -5495 16578
rect -5529 16544 -5495 16546
rect -5529 16478 -5495 16506
rect -5529 16472 -5495 16478
rect -5529 16410 -5495 16434
rect -5529 16400 -5495 16410
rect -5529 16342 -5495 16362
rect -5529 16328 -5495 16342
rect -5529 16274 -5495 16290
rect -5529 16256 -5495 16274
rect -5529 16206 -5495 16218
rect -5529 16184 -5495 16206
rect -5529 16138 -5495 16146
rect -5529 16112 -5495 16138
rect -5443 17056 -5409 17082
rect -5443 17048 -5409 17056
rect -5443 16988 -5409 17010
rect -5443 16976 -5409 16988
rect -5443 16920 -5409 16938
rect -5443 16904 -5409 16920
rect -5443 16852 -5409 16866
rect -5443 16832 -5409 16852
rect -5443 16784 -5409 16794
rect -5443 16760 -5409 16784
rect -5443 16716 -5409 16722
rect -5443 16688 -5409 16716
rect -5443 16648 -5409 16650
rect -5443 16616 -5409 16648
rect -5443 16546 -5409 16578
rect -5443 16544 -5409 16546
rect -5443 16478 -5409 16506
rect -5443 16472 -5409 16478
rect -5443 16410 -5409 16434
rect -5443 16400 -5409 16410
rect -5443 16342 -5409 16362
rect -5443 16328 -5409 16342
rect -5443 16274 -5409 16290
rect -5443 16256 -5409 16274
rect -5443 16206 -5409 16218
rect -5443 16184 -5409 16206
rect -5443 16138 -5409 16146
rect -5443 16112 -5409 16138
rect -5357 17056 -5323 17082
rect -5357 17048 -5323 17056
rect -5357 16988 -5323 17010
rect -5357 16976 -5323 16988
rect -5357 16920 -5323 16938
rect -5357 16904 -5323 16920
rect -5357 16852 -5323 16866
rect -5357 16832 -5323 16852
rect -5357 16784 -5323 16794
rect -5357 16760 -5323 16784
rect -5357 16716 -5323 16722
rect -5357 16688 -5323 16716
rect -5357 16648 -5323 16650
rect -5357 16616 -5323 16648
rect -5357 16546 -5323 16578
rect -5357 16544 -5323 16546
rect -5357 16478 -5323 16506
rect -5357 16472 -5323 16478
rect -5357 16410 -5323 16434
rect -5357 16400 -5323 16410
rect -5357 16342 -5323 16362
rect -5357 16328 -5323 16342
rect -5357 16274 -5323 16290
rect -5357 16256 -5323 16274
rect -5357 16206 -5323 16218
rect -5357 16184 -5323 16206
rect -5357 16138 -5323 16146
rect -5357 16112 -5323 16138
rect -5246 17056 -5212 17082
rect -5246 17048 -5212 17056
rect -5246 16988 -5212 17010
rect -5246 16976 -5212 16988
rect -5246 16920 -5212 16938
rect -5246 16904 -5212 16920
rect -5246 16852 -5212 16866
rect -5246 16832 -5212 16852
rect -5246 16784 -5212 16794
rect -5246 16760 -5212 16784
rect -5246 16716 -5212 16722
rect -5246 16688 -5212 16716
rect -5246 16648 -5212 16650
rect -5246 16616 -5212 16648
rect -5246 16546 -5212 16578
rect -5246 16544 -5212 16546
rect -5246 16478 -5212 16506
rect -5246 16472 -5212 16478
rect -5246 16410 -5212 16434
rect -5246 16400 -5212 16410
rect -5246 16342 -5212 16362
rect -5246 16328 -5212 16342
rect -5246 16274 -5212 16290
rect -5246 16256 -5212 16274
rect -5246 16206 -5212 16218
rect -5246 16184 -5212 16206
rect -5246 16138 -5212 16146
rect -5246 16112 -5212 16138
rect -6697 16020 -6693 16054
rect -6693 16020 -6663 16054
rect -6625 16020 -6591 16054
rect -6553 16020 -6523 16054
rect -6523 16020 -6519 16054
rect -6303 16020 -6299 16054
rect -6299 16020 -6269 16054
rect -6231 16020 -6197 16054
rect -6159 16020 -6129 16054
rect -6129 16020 -6125 16054
rect -5909 16020 -5905 16054
rect -5905 16020 -5875 16054
rect -5837 16020 -5803 16054
rect -5765 16020 -5735 16054
rect -5735 16020 -5731 16054
rect -5515 16020 -5511 16054
rect -5511 16020 -5481 16054
rect -5443 16020 -5409 16054
rect -5371 16020 -5341 16054
rect -5341 16020 -5337 16054
rect -1740 8704 -1620 8760
rect -1740 8670 -1702 8704
rect -1702 8670 -1668 8704
rect -1668 8670 -1620 8704
rect -1740 8640 -1620 8670
rect -1960 7616 -1840 7660
rect -1960 7582 -1918 7616
rect -1918 7582 -1884 7616
rect -1884 7582 -1840 7616
rect -1960 7540 -1840 7582
rect 54 8529 58 8563
rect 58 8529 88 8563
rect 126 8529 160 8563
rect 198 8529 228 8563
rect 228 8529 232 8563
rect 398 8529 402 8563
rect 402 8529 432 8563
rect 470 8529 504 8563
rect 542 8529 572 8563
rect 572 8529 576 8563
rect 742 8529 746 8563
rect 746 8529 776 8563
rect 814 8529 848 8563
rect 886 8529 916 8563
rect 916 8529 920 8563
rect -1540 7532 -1522 8480
rect -1522 7532 -1420 8480
rect -1540 7360 -1420 7532
rect -174 8420 -140 8454
rect -174 8350 -140 8374
rect -174 8340 -140 8350
rect -174 8280 -140 8294
rect -174 8260 -140 8280
rect -174 8210 -140 8214
rect -174 8180 -140 8210
rect -174 8104 -140 8134
rect -174 8100 -140 8104
rect -174 8034 -140 8054
rect -174 8020 -140 8034
rect -174 7964 -140 7974
rect -174 7940 -140 7964
rect -174 7860 -140 7894
rect -174 7790 -140 7814
rect -174 7780 -140 7790
rect -174 7720 -140 7734
rect -174 7700 -140 7720
rect -174 7650 -140 7654
rect -174 7620 -140 7650
rect -174 7544 -140 7574
rect -174 7540 -140 7544
rect -174 7474 -140 7494
rect -174 7460 -140 7474
rect -46 8445 -12 8471
rect -46 8437 -12 8445
rect -46 8377 -12 8399
rect -46 8365 -12 8377
rect -46 8309 -12 8327
rect -46 8293 -12 8309
rect -46 8241 -12 8255
rect -46 8221 -12 8241
rect -46 8173 -12 8183
rect -46 8149 -12 8173
rect -46 8105 -12 8111
rect -46 8077 -12 8105
rect -46 8037 -12 8039
rect -46 8005 -12 8037
rect -46 7935 -12 7967
rect -46 7933 -12 7935
rect -46 7867 -12 7895
rect -46 7861 -12 7867
rect -46 7799 -12 7823
rect -46 7789 -12 7799
rect -46 7731 -12 7751
rect -46 7717 -12 7731
rect -46 7663 -12 7679
rect -46 7645 -12 7663
rect -46 7595 -12 7607
rect -46 7573 -12 7595
rect -46 7527 -12 7535
rect -46 7501 -12 7527
rect 40 8445 74 8471
rect 40 8437 74 8445
rect 40 8377 74 8399
rect 40 8365 74 8377
rect 40 8309 74 8327
rect 40 8293 74 8309
rect 40 8241 74 8255
rect 40 8221 74 8241
rect 40 8173 74 8183
rect 40 8149 74 8173
rect 40 8105 74 8111
rect 40 8077 74 8105
rect 40 8037 74 8039
rect 40 8005 74 8037
rect 40 7935 74 7967
rect 40 7933 74 7935
rect 40 7867 74 7895
rect 40 7861 74 7867
rect 40 7799 74 7823
rect 40 7789 74 7799
rect 40 7731 74 7751
rect 40 7717 74 7731
rect 40 7663 74 7679
rect 40 7645 74 7663
rect 40 7595 74 7607
rect 40 7573 74 7595
rect 40 7527 74 7535
rect 40 7501 74 7527
rect 126 8445 160 8471
rect 126 8437 160 8445
rect 126 8377 160 8399
rect 126 8365 160 8377
rect 126 8309 160 8327
rect 126 8293 160 8309
rect 126 8241 160 8255
rect 126 8221 160 8241
rect 126 8173 160 8183
rect 126 8149 160 8173
rect 126 8105 160 8111
rect 126 8077 160 8105
rect 126 8037 160 8039
rect 126 8005 160 8037
rect 126 7935 160 7967
rect 126 7933 160 7935
rect 126 7867 160 7895
rect 126 7861 160 7867
rect 126 7799 160 7823
rect 126 7789 160 7799
rect 126 7731 160 7751
rect 126 7717 160 7731
rect 126 7663 160 7679
rect 126 7645 160 7663
rect 126 7595 160 7607
rect 126 7573 160 7595
rect 126 7527 160 7535
rect 126 7501 160 7527
rect 212 8445 246 8471
rect 212 8437 246 8445
rect 212 8377 246 8399
rect 212 8365 246 8377
rect 212 8309 246 8327
rect 212 8293 246 8309
rect 212 8241 246 8255
rect 212 8221 246 8241
rect 212 8173 246 8183
rect 212 8149 246 8173
rect 212 8105 246 8111
rect 212 8077 246 8105
rect 212 8037 246 8039
rect 212 8005 246 8037
rect 212 7935 246 7967
rect 212 7933 246 7935
rect 212 7867 246 7895
rect 212 7861 246 7867
rect 212 7799 246 7823
rect 212 7789 246 7799
rect 212 7731 246 7751
rect 212 7717 246 7731
rect 212 7663 246 7679
rect 212 7645 246 7663
rect 212 7595 246 7607
rect 212 7573 246 7595
rect 212 7527 246 7535
rect 212 7501 246 7527
rect 298 8445 332 8471
rect 298 8437 332 8445
rect 298 8377 332 8399
rect 298 8365 332 8377
rect 298 8309 332 8327
rect 298 8293 332 8309
rect 298 8241 332 8255
rect 298 8221 332 8241
rect 298 8173 332 8183
rect 298 8149 332 8173
rect 298 8105 332 8111
rect 298 8077 332 8105
rect 298 8037 332 8039
rect 298 8005 332 8037
rect 298 7935 332 7967
rect 298 7933 332 7935
rect 298 7867 332 7895
rect 298 7861 332 7867
rect 298 7799 332 7823
rect 298 7789 332 7799
rect 298 7731 332 7751
rect 298 7717 332 7731
rect 298 7663 332 7679
rect 298 7645 332 7663
rect 298 7595 332 7607
rect 298 7573 332 7595
rect 298 7527 332 7535
rect 298 7501 332 7527
rect 384 8445 418 8471
rect 384 8437 418 8445
rect 384 8377 418 8399
rect 384 8365 418 8377
rect 384 8309 418 8327
rect 384 8293 418 8309
rect 384 8241 418 8255
rect 384 8221 418 8241
rect 384 8173 418 8183
rect 384 8149 418 8173
rect 384 8105 418 8111
rect 384 8077 418 8105
rect 384 8037 418 8039
rect 384 8005 418 8037
rect 384 7935 418 7967
rect 384 7933 418 7935
rect 384 7867 418 7895
rect 384 7861 418 7867
rect 384 7799 418 7823
rect 384 7789 418 7799
rect 384 7731 418 7751
rect 384 7717 418 7731
rect 384 7663 418 7679
rect 384 7645 418 7663
rect 384 7595 418 7607
rect 384 7573 418 7595
rect 384 7527 418 7535
rect 384 7501 418 7527
rect 470 8445 504 8471
rect 470 8437 504 8445
rect 470 8377 504 8399
rect 470 8365 504 8377
rect 470 8309 504 8327
rect 470 8293 504 8309
rect 470 8241 504 8255
rect 470 8221 504 8241
rect 470 8173 504 8183
rect 470 8149 504 8173
rect 470 8105 504 8111
rect 470 8077 504 8105
rect 470 8037 504 8039
rect 470 8005 504 8037
rect 470 7935 504 7967
rect 470 7933 504 7935
rect 470 7867 504 7895
rect 470 7861 504 7867
rect 470 7799 504 7823
rect 470 7789 504 7799
rect 470 7731 504 7751
rect 470 7717 504 7731
rect 470 7663 504 7679
rect 470 7645 504 7663
rect 470 7595 504 7607
rect 470 7573 504 7595
rect 470 7527 504 7535
rect 470 7501 504 7527
rect 556 8445 590 8471
rect 556 8437 590 8445
rect 556 8377 590 8399
rect 556 8365 590 8377
rect 556 8309 590 8327
rect 556 8293 590 8309
rect 556 8241 590 8255
rect 556 8221 590 8241
rect 556 8173 590 8183
rect 556 8149 590 8173
rect 556 8105 590 8111
rect 556 8077 590 8105
rect 556 8037 590 8039
rect 556 8005 590 8037
rect 556 7935 590 7967
rect 556 7933 590 7935
rect 556 7867 590 7895
rect 556 7861 590 7867
rect 556 7799 590 7823
rect 556 7789 590 7799
rect 556 7731 590 7751
rect 556 7717 590 7731
rect 556 7663 590 7679
rect 556 7645 590 7663
rect 556 7595 590 7607
rect 556 7573 590 7595
rect 556 7527 590 7535
rect 556 7501 590 7527
rect 642 8445 676 8471
rect 642 8437 676 8445
rect 642 8377 676 8399
rect 642 8365 676 8377
rect 642 8309 676 8327
rect 642 8293 676 8309
rect 642 8241 676 8255
rect 642 8221 676 8241
rect 642 8173 676 8183
rect 642 8149 676 8173
rect 642 8105 676 8111
rect 642 8077 676 8105
rect 642 8037 676 8039
rect 642 8005 676 8037
rect 642 7935 676 7967
rect 642 7933 676 7935
rect 642 7867 676 7895
rect 642 7861 676 7867
rect 642 7799 676 7823
rect 642 7789 676 7799
rect 642 7731 676 7751
rect 642 7717 676 7731
rect 642 7663 676 7679
rect 642 7645 676 7663
rect 642 7595 676 7607
rect 642 7573 676 7595
rect 642 7527 676 7535
rect 642 7501 676 7527
rect 728 8445 762 8471
rect 728 8437 762 8445
rect 728 8377 762 8399
rect 728 8365 762 8377
rect 728 8309 762 8327
rect 728 8293 762 8309
rect 728 8241 762 8255
rect 728 8221 762 8241
rect 728 8173 762 8183
rect 728 8149 762 8173
rect 728 8105 762 8111
rect 728 8077 762 8105
rect 728 8037 762 8039
rect 728 8005 762 8037
rect 728 7935 762 7967
rect 728 7933 762 7935
rect 728 7867 762 7895
rect 728 7861 762 7867
rect 728 7799 762 7823
rect 728 7789 762 7799
rect 728 7731 762 7751
rect 728 7717 762 7731
rect 728 7663 762 7679
rect 728 7645 762 7663
rect 728 7595 762 7607
rect 728 7573 762 7595
rect 728 7527 762 7535
rect 728 7501 762 7527
rect 814 8445 848 8471
rect 814 8437 848 8445
rect 814 8377 848 8399
rect 814 8365 848 8377
rect 814 8309 848 8327
rect 814 8293 848 8309
rect 814 8241 848 8255
rect 814 8221 848 8241
rect 814 8173 848 8183
rect 814 8149 848 8173
rect 814 8105 848 8111
rect 814 8077 848 8105
rect 814 8037 848 8039
rect 814 8005 848 8037
rect 814 7935 848 7967
rect 814 7933 848 7935
rect 814 7867 848 7895
rect 814 7861 848 7867
rect 814 7799 848 7823
rect 814 7789 848 7799
rect 814 7731 848 7751
rect 814 7717 848 7731
rect 814 7663 848 7679
rect 814 7645 848 7663
rect 814 7595 848 7607
rect 814 7573 848 7595
rect 814 7527 848 7535
rect 814 7501 848 7527
rect 900 8445 934 8471
rect 900 8437 934 8445
rect 900 8377 934 8399
rect 900 8365 934 8377
rect 900 8309 934 8327
rect 900 8293 934 8309
rect 900 8241 934 8255
rect 900 8221 934 8241
rect 900 8173 934 8183
rect 900 8149 934 8173
rect 900 8105 934 8111
rect 900 8077 934 8105
rect 900 8037 934 8039
rect 900 8005 934 8037
rect 900 7935 934 7967
rect 900 7933 934 7935
rect 900 7867 934 7895
rect 900 7861 934 7867
rect 900 7799 934 7823
rect 900 7789 934 7799
rect 900 7731 934 7751
rect 900 7717 934 7731
rect 900 7663 934 7679
rect 900 7645 934 7663
rect 900 7595 934 7607
rect 900 7573 934 7595
rect 900 7527 934 7535
rect 900 7501 934 7527
rect 986 8445 1020 8471
rect 986 8437 1020 8445
rect 986 8377 1020 8399
rect 986 8365 1020 8377
rect 986 8309 1020 8327
rect 986 8293 1020 8309
rect 986 8241 1020 8255
rect 986 8221 1020 8241
rect 986 8173 1020 8183
rect 986 8149 1020 8173
rect 986 8105 1020 8111
rect 986 8077 1020 8105
rect 986 8037 1020 8039
rect 986 8005 1020 8037
rect 986 7935 1020 7967
rect 986 7933 1020 7935
rect 986 7867 1020 7895
rect 986 7861 1020 7867
rect 986 7799 1020 7823
rect 986 7789 1020 7799
rect 986 7731 1020 7751
rect 986 7717 1020 7731
rect 986 7663 1020 7679
rect 986 7645 1020 7663
rect 986 7595 1020 7607
rect 986 7573 1020 7595
rect 986 7527 1020 7535
rect 986 7501 1020 7527
rect 1116 8420 1150 8454
rect 1116 8350 1150 8374
rect 1116 8340 1150 8350
rect 1116 8280 1150 8294
rect 1116 8260 1150 8280
rect 1116 8210 1150 8214
rect 1116 8180 1150 8210
rect 1116 8104 1150 8134
rect 1116 8100 1150 8104
rect 1116 8034 1150 8054
rect 1116 8020 1150 8034
rect 1116 7964 1150 7974
rect 1116 7940 1150 7964
rect 1116 7860 1150 7894
rect 1116 7790 1150 7814
rect 1116 7780 1150 7790
rect 1116 7720 1150 7734
rect 1116 7700 1150 7720
rect 1116 7650 1150 7654
rect 1116 7620 1150 7650
rect 1116 7544 1150 7574
rect 1116 7540 1150 7544
rect 1116 7474 1150 7494
rect 1116 7460 1150 7474
rect -1380 6994 -1260 7060
rect -1380 5772 -1264 6994
rect -1264 5772 -1260 6994
rect -960 6944 -840 7000
rect -960 6910 -902 6944
rect -902 6910 -868 6944
rect -868 6910 -840 6944
rect -960 6880 -840 6910
rect -1160 5856 -1040 5900
rect -1160 5822 -1118 5856
rect -1118 5822 -1084 5856
rect -1084 5822 -1040 5856
rect -1160 5780 -1040 5822
rect -1380 5700 -1260 5772
rect 30 306 64 320
rect 30 286 64 306
rect 30 236 64 240
rect 30 206 64 236
rect 30 130 64 160
rect 30 126 64 130
rect 30 60 64 80
rect 30 46 64 60
rect 30 -10 64 0
rect 30 -34 64 -10
rect 30 -114 64 -80
rect 30 -184 64 -160
rect 30 -194 64 -184
rect 30 -254 64 -240
rect 30 -274 64 -254
rect 30 -324 64 -320
rect 30 -354 64 -324
rect 30 -430 64 -400
rect 30 -434 64 -430
rect 30 -500 64 -480
rect 30 -514 64 -500
rect 30 -570 64 -560
rect 30 -594 64 -570
rect -4540 -2060 -4420 -640
rect -4260 -773 -4140 -720
rect -4260 -807 -4218 -773
rect -4218 -807 -4184 -773
rect -4184 -807 -4140 -773
rect -4260 -860 -4140 -807
rect -3940 -773 -3820 -720
rect -3940 -807 -3894 -773
rect -3894 -807 -3860 -773
rect -3860 -807 -3820 -773
rect -3940 -860 -3820 -807
rect 30 -674 64 -640
rect 158 253 192 279
rect 158 245 192 253
rect 158 185 192 207
rect 158 173 192 185
rect 158 117 192 135
rect 158 101 192 117
rect 158 49 192 63
rect 158 29 192 49
rect 158 -19 192 -9
rect 158 -43 192 -19
rect 158 -87 192 -81
rect 158 -115 192 -87
rect 158 -155 192 -153
rect 158 -187 192 -155
rect 158 -257 192 -225
rect 158 -259 192 -257
rect 158 -325 192 -297
rect 158 -331 192 -325
rect 158 -393 192 -369
rect 158 -403 192 -393
rect 158 -461 192 -441
rect 158 -475 192 -461
rect 158 -529 192 -513
rect 158 -547 192 -529
rect 158 -597 192 -585
rect 158 -619 192 -597
rect 158 -665 192 -657
rect 158 -691 192 -665
rect 244 253 278 279
rect 244 245 278 253
rect 244 185 278 207
rect 244 173 278 185
rect 244 117 278 135
rect 244 101 278 117
rect 244 49 278 63
rect 244 29 278 49
rect 244 -19 278 -9
rect 244 -43 278 -19
rect 244 -87 278 -81
rect 244 -115 278 -87
rect 244 -155 278 -153
rect 244 -187 278 -155
rect 244 -257 278 -225
rect 244 -259 278 -257
rect 244 -325 278 -297
rect 244 -331 278 -325
rect 244 -393 278 -369
rect 244 -403 278 -393
rect 244 -461 278 -441
rect 244 -475 278 -461
rect 244 -529 278 -513
rect 244 -547 278 -529
rect 244 -597 278 -585
rect 244 -619 278 -597
rect 244 -665 278 -657
rect 244 -691 278 -665
rect 330 253 364 279
rect 330 245 364 253
rect 330 185 364 207
rect 330 173 364 185
rect 330 117 364 135
rect 330 101 364 117
rect 330 49 364 63
rect 330 29 364 49
rect 330 -19 364 -9
rect 330 -43 364 -19
rect 330 -87 364 -81
rect 330 -115 364 -87
rect 330 -155 364 -153
rect 330 -187 364 -155
rect 330 -257 364 -225
rect 330 -259 364 -257
rect 330 -325 364 -297
rect 330 -331 364 -325
rect 330 -393 364 -369
rect 330 -403 364 -393
rect 330 -461 364 -441
rect 330 -475 364 -461
rect 330 -529 364 -513
rect 330 -547 364 -529
rect 330 -597 364 -585
rect 330 -619 364 -597
rect 330 -665 364 -657
rect 330 -691 364 -665
rect 416 253 450 279
rect 416 245 450 253
rect 416 185 450 207
rect 416 173 450 185
rect 416 117 450 135
rect 416 101 450 117
rect 416 49 450 63
rect 416 29 450 49
rect 416 -19 450 -9
rect 416 -43 450 -19
rect 416 -87 450 -81
rect 416 -115 450 -87
rect 416 -155 450 -153
rect 416 -187 450 -155
rect 416 -257 450 -225
rect 416 -259 450 -257
rect 416 -325 450 -297
rect 416 -331 450 -325
rect 416 -393 450 -369
rect 416 -403 450 -393
rect 416 -461 450 -441
rect 416 -475 450 -461
rect 416 -529 450 -513
rect 416 -547 450 -529
rect 416 -597 450 -585
rect 416 -619 450 -597
rect 416 -665 450 -657
rect 416 -691 450 -665
rect 502 253 536 279
rect 502 245 536 253
rect 502 185 536 207
rect 502 173 536 185
rect 502 117 536 135
rect 502 101 536 117
rect 502 49 536 63
rect 502 29 536 49
rect 502 -19 536 -9
rect 502 -43 536 -19
rect 502 -87 536 -81
rect 502 -115 536 -87
rect 502 -155 536 -153
rect 502 -187 536 -155
rect 502 -257 536 -225
rect 502 -259 536 -257
rect 502 -325 536 -297
rect 502 -331 536 -325
rect 502 -393 536 -369
rect 502 -403 536 -393
rect 502 -461 536 -441
rect 502 -475 536 -461
rect 502 -529 536 -513
rect 502 -547 536 -529
rect 502 -597 536 -585
rect 502 -619 536 -597
rect 502 -665 536 -657
rect 502 -691 536 -665
rect 588 253 622 279
rect 588 245 622 253
rect 588 185 622 207
rect 588 173 622 185
rect 588 117 622 135
rect 588 101 622 117
rect 588 49 622 63
rect 588 29 622 49
rect 588 -19 622 -9
rect 588 -43 622 -19
rect 588 -87 622 -81
rect 588 -115 622 -87
rect 588 -155 622 -153
rect 588 -187 622 -155
rect 588 -257 622 -225
rect 588 -259 622 -257
rect 588 -325 622 -297
rect 588 -331 622 -325
rect 588 -393 622 -369
rect 588 -403 622 -393
rect 588 -461 622 -441
rect 588 -475 622 -461
rect 588 -529 622 -513
rect 588 -547 622 -529
rect 588 -597 622 -585
rect 588 -619 622 -597
rect 588 -665 622 -657
rect 588 -691 622 -665
rect 674 253 708 279
rect 674 245 708 253
rect 674 185 708 207
rect 674 173 708 185
rect 674 117 708 135
rect 674 101 708 117
rect 674 49 708 63
rect 674 29 708 49
rect 674 -19 708 -9
rect 674 -43 708 -19
rect 674 -87 708 -81
rect 674 -115 708 -87
rect 674 -155 708 -153
rect 674 -187 708 -155
rect 674 -257 708 -225
rect 674 -259 708 -257
rect 674 -325 708 -297
rect 674 -331 708 -325
rect 674 -393 708 -369
rect 674 -403 708 -393
rect 674 -461 708 -441
rect 674 -475 708 -461
rect 674 -529 708 -513
rect 674 -547 708 -529
rect 674 -597 708 -585
rect 674 -619 708 -597
rect 674 -665 708 -657
rect 674 -691 708 -665
rect 760 253 794 279
rect 760 245 794 253
rect 760 185 794 207
rect 760 173 794 185
rect 760 117 794 135
rect 760 101 794 117
rect 760 49 794 63
rect 760 29 794 49
rect 760 -19 794 -9
rect 760 -43 794 -19
rect 760 -87 794 -81
rect 760 -115 794 -87
rect 760 -155 794 -153
rect 760 -187 794 -155
rect 760 -257 794 -225
rect 760 -259 794 -257
rect 760 -325 794 -297
rect 760 -331 794 -325
rect 760 -393 794 -369
rect 760 -403 794 -393
rect 760 -461 794 -441
rect 760 -475 794 -461
rect 760 -529 794 -513
rect 760 -547 794 -529
rect 760 -597 794 -585
rect 760 -619 794 -597
rect 760 -665 794 -657
rect 760 -691 794 -665
rect 846 253 880 279
rect 846 245 880 253
rect 846 185 880 207
rect 846 173 880 185
rect 846 117 880 135
rect 846 101 880 117
rect 846 49 880 63
rect 846 29 880 49
rect 846 -19 880 -9
rect 846 -43 880 -19
rect 846 -87 880 -81
rect 846 -115 880 -87
rect 846 -155 880 -153
rect 846 -187 880 -155
rect 846 -257 880 -225
rect 846 -259 880 -257
rect 846 -325 880 -297
rect 846 -331 880 -325
rect 846 -393 880 -369
rect 846 -403 880 -393
rect 846 -461 880 -441
rect 846 -475 880 -461
rect 846 -529 880 -513
rect 846 -547 880 -529
rect 846 -597 880 -585
rect 846 -619 880 -597
rect 846 -665 880 -657
rect 846 -691 880 -665
rect 967 306 1001 320
rect 967 286 1001 306
rect 967 236 1001 240
rect 967 206 1001 236
rect 967 130 1001 160
rect 967 126 1001 130
rect 967 60 1001 80
rect 967 46 1001 60
rect 967 -10 1001 0
rect 967 -34 1001 -10
rect 967 -114 1001 -80
rect 967 -184 1001 -160
rect 967 -194 1001 -184
rect 967 -254 1001 -240
rect 967 -274 1001 -254
rect 967 -324 1001 -320
rect 967 -354 1001 -324
rect 967 -430 1001 -400
rect 967 -434 1001 -430
rect 967 -500 1001 -480
rect 967 -514 1001 -500
rect 967 -570 1001 -560
rect 967 -594 1001 -570
rect 967 -674 1001 -640
rect 258 -783 262 -749
rect 262 -783 292 -749
rect 330 -783 364 -749
rect 402 -783 432 -749
rect 432 -783 436 -749
rect 602 -783 606 -749
rect 606 -783 636 -749
rect 674 -783 708 -749
rect 746 -783 776 -749
rect 776 -783 780 -749
rect -4540 -2064 -4268 -2060
rect -4268 -2064 -3810 -2060
rect -3810 -2064 -3740 -2060
rect -4540 -2220 -3740 -2064
<< metal1 >>
rect -6840 17094 -6780 17280
rect -6720 17240 -6500 17260
rect -6720 17160 -6700 17240
rect -6520 17174 -6500 17240
rect -6720 17140 -6697 17160
rect -6663 17140 -6625 17160
rect -6591 17140 -6553 17160
rect -6519 17140 -6500 17174
rect -6709 17128 -6507 17140
rect -6840 17082 -6776 17094
rect -6840 17048 -6822 17082
rect -6788 17048 -6776 17082
rect -6840 17010 -6776 17048
rect -6840 16976 -6822 17010
rect -6788 16976 -6776 17010
rect -6840 16938 -6776 16976
rect -6840 16904 -6822 16938
rect -6788 16904 -6776 16938
rect -6840 16866 -6776 16904
rect -6840 16832 -6822 16866
rect -6788 16832 -6776 16866
rect -6840 16794 -6776 16832
rect -6840 16760 -6822 16794
rect -6788 16760 -6776 16794
rect -6840 16722 -6776 16760
rect -6840 16688 -6822 16722
rect -6788 16688 -6776 16722
rect -6840 16650 -6776 16688
rect -6840 16616 -6822 16650
rect -6788 16616 -6776 16650
rect -6840 16578 -6776 16616
rect -6840 16544 -6822 16578
rect -6788 16544 -6776 16578
rect -6840 16506 -6776 16544
rect -6840 16472 -6822 16506
rect -6788 16472 -6776 16506
rect -6840 16434 -6776 16472
rect -6840 16400 -6822 16434
rect -6788 16400 -6776 16434
rect -6840 16362 -6776 16400
rect -6840 16328 -6822 16362
rect -6788 16328 -6776 16362
rect -6840 16290 -6776 16328
rect -6840 16256 -6822 16290
rect -6788 16256 -6776 16290
rect -6840 16218 -6776 16256
rect -6840 16184 -6822 16218
rect -6788 16184 -6776 16218
rect -6840 16146 -6776 16184
rect -6840 16112 -6822 16146
rect -6788 16112 -6776 16146
rect -6840 16100 -6776 16112
rect -6720 17082 -6668 17094
rect -6720 17048 -6711 17082
rect -6677 17048 -6668 17082
rect -6720 17010 -6668 17048
rect -6720 16976 -6711 17010
rect -6677 16976 -6668 17010
rect -6720 16938 -6668 16976
rect -6720 16904 -6711 16938
rect -6677 16904 -6668 16938
rect -6720 16866 -6668 16904
rect -6720 16832 -6711 16866
rect -6677 16832 -6668 16866
rect -6720 16794 -6668 16832
rect -6720 16760 -6711 16794
rect -6677 16760 -6668 16794
rect -6720 16722 -6668 16760
rect -6720 16688 -6711 16722
rect -6677 16688 -6668 16722
rect -6720 16650 -6668 16688
rect -6720 16616 -6711 16650
rect -6677 16616 -6668 16650
rect -6720 16578 -6668 16616
rect -6720 16544 -6711 16578
rect -6677 16544 -6668 16578
rect -6720 16542 -6668 16544
rect -6720 16478 -6711 16490
rect -6677 16478 -6668 16490
rect -6720 16414 -6711 16426
rect -6677 16414 -6668 16426
rect -6720 16350 -6711 16362
rect -6677 16350 -6668 16362
rect -6720 16290 -6668 16298
rect -6720 16286 -6711 16290
rect -6677 16286 -6668 16290
rect -6720 16222 -6668 16234
rect -6720 16158 -6668 16170
rect -6720 16100 -6668 16106
rect -6634 17088 -6582 17094
rect -6634 17024 -6582 17036
rect -6634 16960 -6582 16972
rect -6634 16904 -6625 16908
rect -6591 16904 -6582 16908
rect -6634 16896 -6582 16904
rect -6634 16832 -6625 16844
rect -6591 16832 -6582 16844
rect -6634 16768 -6625 16780
rect -6591 16768 -6582 16780
rect -6634 16704 -6625 16716
rect -6591 16704 -6582 16716
rect -6634 16650 -6582 16652
rect -6634 16616 -6625 16650
rect -6591 16616 -6582 16650
rect -6634 16578 -6582 16616
rect -6634 16544 -6625 16578
rect -6591 16544 -6582 16578
rect -6634 16506 -6582 16544
rect -6634 16472 -6625 16506
rect -6591 16472 -6582 16506
rect -6634 16434 -6582 16472
rect -6634 16400 -6625 16434
rect -6591 16400 -6582 16434
rect -6634 16362 -6582 16400
rect -6634 16328 -6625 16362
rect -6591 16328 -6582 16362
rect -6634 16290 -6582 16328
rect -6634 16256 -6625 16290
rect -6591 16256 -6582 16290
rect -6634 16218 -6582 16256
rect -6634 16184 -6625 16218
rect -6591 16184 -6582 16218
rect -6634 16146 -6582 16184
rect -6634 16112 -6625 16146
rect -6591 16112 -6582 16146
rect -6634 16100 -6582 16112
rect -6548 17082 -6496 17094
rect -6548 17048 -6539 17082
rect -6505 17048 -6496 17082
rect -6548 17010 -6496 17048
rect -6548 16976 -6539 17010
rect -6505 16976 -6496 17010
rect -6548 16938 -6496 16976
rect -6548 16904 -6539 16938
rect -6505 16904 -6496 16938
rect -6548 16866 -6496 16904
rect -6548 16832 -6539 16866
rect -6505 16832 -6496 16866
rect -6548 16794 -6496 16832
rect -6548 16760 -6539 16794
rect -6505 16760 -6496 16794
rect -6548 16722 -6496 16760
rect -6548 16688 -6539 16722
rect -6505 16688 -6496 16722
rect -6548 16650 -6496 16688
rect -6548 16616 -6539 16650
rect -6505 16616 -6496 16650
rect -6548 16578 -6496 16616
rect -6548 16544 -6539 16578
rect -6505 16544 -6496 16578
rect -6548 16542 -6496 16544
rect -6548 16478 -6539 16490
rect -6505 16478 -6496 16490
rect -6548 16414 -6539 16426
rect -6505 16414 -6496 16426
rect -6548 16350 -6539 16362
rect -6505 16350 -6496 16362
rect -6548 16290 -6496 16298
rect -6548 16286 -6539 16290
rect -6505 16286 -6496 16290
rect -6548 16222 -6496 16234
rect -6548 16158 -6496 16170
rect -6548 16100 -6496 16106
rect -6440 17082 -6380 17280
rect -6320 17240 -6100 17260
rect -6320 17174 -6300 17240
rect -6320 17140 -6303 17174
rect -6120 17160 -6100 17240
rect -6269 17140 -6231 17160
rect -6197 17140 -6159 17160
rect -6125 17140 -6100 17160
rect -6315 17128 -6113 17140
rect -6040 17094 -5980 17280
rect -5920 17240 -5700 17260
rect -5920 17194 -5900 17240
rect -5921 17174 -5900 17194
rect -5921 17140 -5909 17174
rect -5720 17160 -5700 17240
rect -5875 17140 -5837 17160
rect -5803 17140 -5765 17160
rect -5731 17140 -5700 17160
rect -5921 17128 -5719 17140
rect -5660 17094 -5600 17280
rect -5540 17240 -5320 17260
rect -5540 17160 -5520 17240
rect -5340 17174 -5320 17240
rect -5540 17140 -5515 17160
rect -5481 17140 -5443 17160
rect -5409 17140 -5371 17160
rect -5337 17140 -5320 17174
rect -5527 17128 -5325 17140
rect -6440 17048 -6428 17082
rect -6394 17048 -6380 17082
rect -6440 17010 -6380 17048
rect -6440 16976 -6428 17010
rect -6394 16976 -6380 17010
rect -6440 16938 -6380 16976
rect -6440 16904 -6428 16938
rect -6394 16904 -6380 16938
rect -6440 16866 -6380 16904
rect -6440 16832 -6428 16866
rect -6394 16832 -6380 16866
rect -6440 16794 -6380 16832
rect -6440 16760 -6428 16794
rect -6394 16760 -6380 16794
rect -6440 16722 -6380 16760
rect -6440 16688 -6428 16722
rect -6394 16688 -6380 16722
rect -6440 16650 -6380 16688
rect -6440 16616 -6428 16650
rect -6394 16616 -6380 16650
rect -6440 16578 -6380 16616
rect -6440 16544 -6428 16578
rect -6394 16544 -6380 16578
rect -6440 16506 -6380 16544
rect -6440 16472 -6428 16506
rect -6394 16472 -6380 16506
rect -6440 16434 -6380 16472
rect -6440 16400 -6428 16434
rect -6394 16400 -6380 16434
rect -6440 16362 -6380 16400
rect -6440 16328 -6428 16362
rect -6394 16328 -6380 16362
rect -6440 16290 -6380 16328
rect -6440 16256 -6428 16290
rect -6394 16256 -6380 16290
rect -6440 16218 -6380 16256
rect -6440 16184 -6428 16218
rect -6394 16184 -6380 16218
rect -6440 16146 -6380 16184
rect -6440 16112 -6428 16146
rect -6394 16112 -6380 16146
rect -6840 15920 -6780 16100
rect -6709 16054 -6507 16066
rect -6709 16020 -6697 16054
rect -6663 16020 -6625 16054
rect -6591 16020 -6553 16054
rect -6519 16020 -6507 16054
rect -6709 16000 -6507 16020
rect -6440 15920 -6380 16112
rect -6326 17082 -6274 17094
rect -6326 17048 -6317 17082
rect -6283 17048 -6274 17082
rect -6326 17010 -6274 17048
rect -6326 16976 -6317 17010
rect -6283 16976 -6274 17010
rect -6326 16938 -6274 16976
rect -6326 16904 -6317 16938
rect -6283 16904 -6274 16938
rect -6326 16866 -6274 16904
rect -6326 16832 -6317 16866
rect -6283 16832 -6274 16866
rect -6326 16794 -6274 16832
rect -6326 16760 -6317 16794
rect -6283 16760 -6274 16794
rect -6326 16722 -6274 16760
rect -6326 16688 -6317 16722
rect -6283 16688 -6274 16722
rect -6326 16650 -6274 16688
rect -6326 16616 -6317 16650
rect -6283 16616 -6274 16650
rect -6326 16578 -6274 16616
rect -6326 16544 -6317 16578
rect -6283 16544 -6274 16578
rect -6326 16542 -6274 16544
rect -6326 16478 -6317 16490
rect -6283 16478 -6274 16490
rect -6326 16414 -6317 16426
rect -6283 16414 -6274 16426
rect -6326 16350 -6317 16362
rect -6283 16350 -6274 16362
rect -6326 16290 -6274 16298
rect -6326 16286 -6317 16290
rect -6283 16286 -6274 16290
rect -6326 16222 -6274 16234
rect -6326 16158 -6274 16170
rect -6326 16100 -6274 16106
rect -6240 17088 -6188 17094
rect -6240 17024 -6188 17036
rect -6240 16960 -6188 16972
rect -6240 16904 -6231 16908
rect -6197 16904 -6188 16908
rect -6240 16896 -6188 16904
rect -6240 16832 -6231 16844
rect -6197 16832 -6188 16844
rect -6240 16768 -6231 16780
rect -6197 16768 -6188 16780
rect -6240 16704 -6231 16716
rect -6197 16704 -6188 16716
rect -6240 16650 -6188 16652
rect -6240 16616 -6231 16650
rect -6197 16616 -6188 16650
rect -6240 16578 -6188 16616
rect -6240 16544 -6231 16578
rect -6197 16544 -6188 16578
rect -6240 16506 -6188 16544
rect -6240 16472 -6231 16506
rect -6197 16472 -6188 16506
rect -6240 16434 -6188 16472
rect -6240 16400 -6231 16434
rect -6197 16400 -6188 16434
rect -6240 16362 -6188 16400
rect -6240 16328 -6231 16362
rect -6197 16328 -6188 16362
rect -6240 16290 -6188 16328
rect -6240 16256 -6231 16290
rect -6197 16256 -6188 16290
rect -6240 16218 -6188 16256
rect -6240 16184 -6231 16218
rect -6197 16184 -6188 16218
rect -6240 16146 -6188 16184
rect -6240 16112 -6231 16146
rect -6197 16112 -6188 16146
rect -6240 16100 -6188 16112
rect -6154 17082 -6102 17094
rect -6154 17048 -6145 17082
rect -6111 17048 -6102 17082
rect -6154 17010 -6102 17048
rect -6154 16976 -6145 17010
rect -6111 16976 -6102 17010
rect -6154 16938 -6102 16976
rect -6154 16904 -6145 16938
rect -6111 16904 -6102 16938
rect -6154 16866 -6102 16904
rect -6154 16832 -6145 16866
rect -6111 16832 -6102 16866
rect -6154 16794 -6102 16832
rect -6154 16760 -6145 16794
rect -6111 16760 -6102 16794
rect -6154 16722 -6102 16760
rect -6154 16688 -6145 16722
rect -6111 16688 -6102 16722
rect -6154 16650 -6102 16688
rect -6154 16616 -6145 16650
rect -6111 16616 -6102 16650
rect -6154 16578 -6102 16616
rect -6154 16544 -6145 16578
rect -6111 16544 -6102 16578
rect -6154 16542 -6102 16544
rect -6154 16478 -6145 16490
rect -6111 16478 -6102 16490
rect -6154 16414 -6145 16426
rect -6111 16414 -6102 16426
rect -6154 16350 -6145 16362
rect -6111 16350 -6102 16362
rect -6154 16290 -6102 16298
rect -6154 16286 -6145 16290
rect -6111 16286 -6102 16290
rect -6154 16222 -6102 16234
rect -6154 16158 -6102 16170
rect -6154 16100 -6102 16106
rect -6046 17082 -5980 17094
rect -6046 17048 -6034 17082
rect -6000 17048 -5980 17082
rect -6046 17010 -5980 17048
rect -6046 16976 -6034 17010
rect -6000 16976 -5980 17010
rect -6046 16938 -5980 16976
rect -6046 16904 -6034 16938
rect -6000 16904 -5980 16938
rect -6046 16866 -5980 16904
rect -6046 16832 -6034 16866
rect -6000 16832 -5980 16866
rect -6046 16794 -5980 16832
rect -6046 16760 -6034 16794
rect -6000 16760 -5980 16794
rect -6046 16722 -5980 16760
rect -6046 16688 -6034 16722
rect -6000 16688 -5980 16722
rect -6046 16650 -5980 16688
rect -6046 16616 -6034 16650
rect -6000 16616 -5980 16650
rect -6046 16578 -5980 16616
rect -6046 16544 -6034 16578
rect -6000 16544 -5980 16578
rect -6046 16506 -5980 16544
rect -6046 16472 -6034 16506
rect -6000 16472 -5980 16506
rect -6046 16434 -5980 16472
rect -6046 16400 -6034 16434
rect -6000 16400 -5980 16434
rect -6046 16362 -5980 16400
rect -6046 16328 -6034 16362
rect -6000 16328 -5980 16362
rect -6046 16290 -5980 16328
rect -6046 16256 -6034 16290
rect -6000 16256 -5980 16290
rect -6046 16218 -5980 16256
rect -6046 16184 -6034 16218
rect -6000 16184 -5980 16218
rect -6046 16146 -5980 16184
rect -6046 16112 -6034 16146
rect -6000 16112 -5980 16146
rect -6046 16100 -5980 16112
rect -5932 17082 -5880 17094
rect -5932 17048 -5923 17082
rect -5889 17048 -5880 17082
rect -5932 17010 -5880 17048
rect -5932 16976 -5923 17010
rect -5889 16976 -5880 17010
rect -5932 16938 -5880 16976
rect -5932 16904 -5923 16938
rect -5889 16904 -5880 16938
rect -5932 16866 -5880 16904
rect -5932 16832 -5923 16866
rect -5889 16832 -5880 16866
rect -5932 16794 -5880 16832
rect -5932 16760 -5923 16794
rect -5889 16760 -5880 16794
rect -5932 16722 -5880 16760
rect -5932 16688 -5923 16722
rect -5889 16688 -5880 16722
rect -5932 16650 -5880 16688
rect -5932 16616 -5923 16650
rect -5889 16616 -5880 16650
rect -5932 16578 -5880 16616
rect -5932 16544 -5923 16578
rect -5889 16544 -5880 16578
rect -5932 16542 -5880 16544
rect -5932 16478 -5923 16490
rect -5889 16478 -5880 16490
rect -5932 16414 -5923 16426
rect -5889 16414 -5880 16426
rect -5932 16350 -5923 16362
rect -5889 16350 -5880 16362
rect -5932 16290 -5880 16298
rect -5932 16286 -5923 16290
rect -5889 16286 -5880 16290
rect -5932 16222 -5880 16234
rect -5932 16158 -5880 16170
rect -5932 16100 -5880 16106
rect -5846 17088 -5794 17094
rect -5846 17024 -5794 17036
rect -5846 16960 -5794 16972
rect -5846 16904 -5837 16908
rect -5803 16904 -5794 16908
rect -5846 16896 -5794 16904
rect -5846 16832 -5837 16844
rect -5803 16832 -5794 16844
rect -5846 16768 -5837 16780
rect -5803 16768 -5794 16780
rect -5846 16704 -5837 16716
rect -5803 16704 -5794 16716
rect -5846 16650 -5794 16652
rect -5846 16616 -5837 16650
rect -5803 16616 -5794 16650
rect -5846 16578 -5794 16616
rect -5846 16544 -5837 16578
rect -5803 16544 -5794 16578
rect -5846 16506 -5794 16544
rect -5846 16472 -5837 16506
rect -5803 16472 -5794 16506
rect -5846 16434 -5794 16472
rect -5846 16400 -5837 16434
rect -5803 16400 -5794 16434
rect -5846 16362 -5794 16400
rect -5846 16328 -5837 16362
rect -5803 16328 -5794 16362
rect -5846 16290 -5794 16328
rect -5846 16256 -5837 16290
rect -5803 16256 -5794 16290
rect -5846 16218 -5794 16256
rect -5846 16184 -5837 16218
rect -5803 16184 -5794 16218
rect -5846 16146 -5794 16184
rect -5846 16112 -5837 16146
rect -5803 16112 -5794 16146
rect -5846 16100 -5794 16112
rect -5760 17082 -5708 17094
rect -5760 17048 -5751 17082
rect -5717 17048 -5708 17082
rect -5760 17010 -5708 17048
rect -5760 16976 -5751 17010
rect -5717 16976 -5708 17010
rect -5760 16938 -5708 16976
rect -5760 16904 -5751 16938
rect -5717 16904 -5708 16938
rect -5760 16866 -5708 16904
rect -5760 16832 -5751 16866
rect -5717 16832 -5708 16866
rect -5760 16794 -5708 16832
rect -5760 16760 -5751 16794
rect -5717 16760 -5708 16794
rect -5760 16722 -5708 16760
rect -5760 16688 -5751 16722
rect -5717 16688 -5708 16722
rect -5760 16650 -5708 16688
rect -5760 16616 -5751 16650
rect -5717 16616 -5708 16650
rect -5760 16578 -5708 16616
rect -5760 16544 -5751 16578
rect -5717 16544 -5708 16578
rect -5760 16542 -5708 16544
rect -5760 16478 -5751 16490
rect -5717 16478 -5708 16490
rect -5760 16414 -5751 16426
rect -5717 16414 -5708 16426
rect -5760 16350 -5751 16362
rect -5717 16350 -5708 16362
rect -5760 16290 -5708 16298
rect -5760 16286 -5751 16290
rect -5717 16286 -5708 16290
rect -5760 16222 -5708 16234
rect -5760 16158 -5708 16170
rect -5760 16100 -5708 16106
rect -5660 17082 -5594 17094
rect -5660 17048 -5640 17082
rect -5606 17048 -5594 17082
rect -5660 17010 -5594 17048
rect -5660 16976 -5640 17010
rect -5606 16976 -5594 17010
rect -5660 16938 -5594 16976
rect -5660 16904 -5640 16938
rect -5606 16904 -5594 16938
rect -5660 16866 -5594 16904
rect -5660 16832 -5640 16866
rect -5606 16832 -5594 16866
rect -5660 16794 -5594 16832
rect -5660 16760 -5640 16794
rect -5606 16760 -5594 16794
rect -5660 16722 -5594 16760
rect -5660 16688 -5640 16722
rect -5606 16688 -5594 16722
rect -5660 16650 -5594 16688
rect -5660 16616 -5640 16650
rect -5606 16616 -5594 16650
rect -5660 16578 -5594 16616
rect -5660 16544 -5640 16578
rect -5606 16544 -5594 16578
rect -5660 16506 -5594 16544
rect -5660 16472 -5640 16506
rect -5606 16472 -5594 16506
rect -5660 16434 -5594 16472
rect -5660 16400 -5640 16434
rect -5606 16400 -5594 16434
rect -5660 16362 -5594 16400
rect -5660 16328 -5640 16362
rect -5606 16328 -5594 16362
rect -5660 16290 -5594 16328
rect -5660 16256 -5640 16290
rect -5606 16256 -5594 16290
rect -5660 16218 -5594 16256
rect -5660 16184 -5640 16218
rect -5606 16184 -5594 16218
rect -5660 16146 -5594 16184
rect -5660 16112 -5640 16146
rect -5606 16112 -5594 16146
rect -5660 16100 -5594 16112
rect -5538 17082 -5486 17094
rect -5538 17048 -5529 17082
rect -5495 17048 -5486 17082
rect -5538 17010 -5486 17048
rect -5538 16976 -5529 17010
rect -5495 16976 -5486 17010
rect -5538 16938 -5486 16976
rect -5538 16904 -5529 16938
rect -5495 16904 -5486 16938
rect -5538 16866 -5486 16904
rect -5538 16832 -5529 16866
rect -5495 16832 -5486 16866
rect -5538 16794 -5486 16832
rect -5538 16760 -5529 16794
rect -5495 16760 -5486 16794
rect -5538 16722 -5486 16760
rect -5538 16688 -5529 16722
rect -5495 16688 -5486 16722
rect -5538 16650 -5486 16688
rect -5538 16616 -5529 16650
rect -5495 16616 -5486 16650
rect -5538 16578 -5486 16616
rect -5538 16544 -5529 16578
rect -5495 16544 -5486 16578
rect -5538 16542 -5486 16544
rect -5538 16478 -5529 16490
rect -5495 16478 -5486 16490
rect -5538 16414 -5529 16426
rect -5495 16414 -5486 16426
rect -5538 16350 -5529 16362
rect -5495 16350 -5486 16362
rect -5538 16290 -5486 16298
rect -5538 16286 -5529 16290
rect -5495 16286 -5486 16290
rect -5538 16222 -5486 16234
rect -5538 16158 -5486 16170
rect -5538 16100 -5486 16106
rect -5452 17088 -5400 17094
rect -5452 17024 -5400 17036
rect -5452 16960 -5400 16972
rect -5452 16904 -5443 16908
rect -5409 16904 -5400 16908
rect -5452 16896 -5400 16904
rect -5452 16832 -5443 16844
rect -5409 16832 -5400 16844
rect -5452 16768 -5443 16780
rect -5409 16768 -5400 16780
rect -5452 16704 -5443 16716
rect -5409 16704 -5400 16716
rect -5452 16650 -5400 16652
rect -5452 16616 -5443 16650
rect -5409 16616 -5400 16650
rect -5452 16578 -5400 16616
rect -5452 16544 -5443 16578
rect -5409 16544 -5400 16578
rect -5452 16506 -5400 16544
rect -5452 16472 -5443 16506
rect -5409 16472 -5400 16506
rect -5452 16434 -5400 16472
rect -5452 16400 -5443 16434
rect -5409 16400 -5400 16434
rect -5452 16362 -5400 16400
rect -5452 16328 -5443 16362
rect -5409 16328 -5400 16362
rect -5452 16290 -5400 16328
rect -5452 16256 -5443 16290
rect -5409 16256 -5400 16290
rect -5452 16218 -5400 16256
rect -5452 16184 -5443 16218
rect -5409 16184 -5400 16218
rect -5452 16146 -5400 16184
rect -5452 16112 -5443 16146
rect -5409 16112 -5400 16146
rect -5452 16100 -5400 16112
rect -5366 17082 -5314 17094
rect -5366 17048 -5357 17082
rect -5323 17048 -5314 17082
rect -5366 17010 -5314 17048
rect -5366 16976 -5357 17010
rect -5323 16976 -5314 17010
rect -5366 16938 -5314 16976
rect -5366 16904 -5357 16938
rect -5323 16904 -5314 16938
rect -5366 16866 -5314 16904
rect -5366 16832 -5357 16866
rect -5323 16832 -5314 16866
rect -5366 16794 -5314 16832
rect -5366 16760 -5357 16794
rect -5323 16760 -5314 16794
rect -5366 16722 -5314 16760
rect -5366 16688 -5357 16722
rect -5323 16688 -5314 16722
rect -5366 16650 -5314 16688
rect -5366 16616 -5357 16650
rect -5323 16616 -5314 16650
rect -5366 16578 -5314 16616
rect -5366 16544 -5357 16578
rect -5323 16544 -5314 16578
rect -5366 16542 -5314 16544
rect -5366 16478 -5357 16490
rect -5323 16478 -5314 16490
rect -5366 16414 -5357 16426
rect -5323 16414 -5314 16426
rect -5366 16350 -5357 16362
rect -5323 16350 -5314 16362
rect -5366 16290 -5314 16298
rect -5366 16286 -5357 16290
rect -5323 16286 -5314 16290
rect -5366 16222 -5314 16234
rect -5366 16158 -5314 16170
rect -5366 16100 -5314 16106
rect -5260 17082 -5200 17280
rect -5260 17048 -5246 17082
rect -5212 17048 -5200 17082
rect -5260 17010 -5200 17048
rect -5260 16976 -5246 17010
rect -5212 16976 -5200 17010
rect -5260 16938 -5200 16976
rect -5260 16904 -5246 16938
rect -5212 16904 -5200 16938
rect -5260 16866 -5200 16904
rect -5260 16832 -5246 16866
rect -5212 16832 -5200 16866
rect -5260 16794 -5200 16832
rect -5260 16760 -5246 16794
rect -5212 16760 -5200 16794
rect -5260 16722 -5200 16760
rect -5260 16688 -5246 16722
rect -5212 16688 -5200 16722
rect -5260 16650 -5200 16688
rect -5260 16616 -5246 16650
rect -5212 16616 -5200 16650
rect -5260 16578 -5200 16616
rect -5260 16544 -5246 16578
rect -5212 16544 -5200 16578
rect -5260 16506 -5200 16544
rect -5260 16472 -5246 16506
rect -5212 16472 -5200 16506
rect -5260 16434 -5200 16472
rect -5260 16400 -5246 16434
rect -5212 16400 -5200 16434
rect -5260 16362 -5200 16400
rect -5260 16328 -5246 16362
rect -5212 16328 -5200 16362
rect -5260 16290 -5200 16328
rect -5260 16256 -5246 16290
rect -5212 16256 -5200 16290
rect -5260 16218 -5200 16256
rect -5260 16184 -5246 16218
rect -5212 16184 -5200 16218
rect -5260 16146 -5200 16184
rect -5260 16112 -5246 16146
rect -5212 16112 -5200 16146
rect -6315 16054 -6113 16066
rect -6315 16020 -6303 16054
rect -6269 16020 -6231 16054
rect -6197 16020 -6159 16054
rect -6125 16020 -6113 16054
rect -6315 16000 -6113 16020
rect -6040 15920 -5980 16100
rect -5921 16054 -5719 16066
rect -5921 16020 -5909 16054
rect -5875 16020 -5837 16054
rect -5803 16020 -5765 16054
rect -5731 16020 -5719 16054
rect -5921 16000 -5719 16020
rect -5660 15920 -5600 16100
rect -5527 16054 -5325 16066
rect -5527 16020 -5515 16054
rect -5481 16020 -5443 16054
rect -5409 16020 -5371 16054
rect -5337 16020 -5325 16054
rect -5527 16000 -5325 16020
rect -5260 15920 -5200 16112
rect -6840 15900 -5200 15920
rect -6840 15820 -6740 15900
rect -6460 15820 -6000 15900
rect -5280 15820 -5200 15900
rect -6840 15800 -5200 15820
rect -1800 8760 1000 8800
rect -4800 8600 -2000 8700
rect -1800 8640 -1740 8760
rect -1620 8680 1000 8760
rect -1620 8640 1016 8680
rect -1800 8620 1016 8640
rect -1800 8600 1004 8620
rect -4800 7800 -4700 8600
rect -4500 8580 -4380 8600
rect -4120 8580 -3880 8600
rect -3620 8580 -3380 8600
rect -3120 8580 -2880 8600
rect -2620 8580 -2380 8600
rect -2120 8580 -2000 8600
rect -4500 8320 -4400 8580
rect -4100 8320 -3900 8580
rect -3600 8320 -3400 8580
rect -3100 8320 -2900 8580
rect -2600 8320 -2400 8580
rect -2100 8320 -2000 8580
rect -30 8563 1004 8600
rect -30 8529 54 8563
rect 88 8529 126 8563
rect 160 8529 198 8563
rect 232 8529 398 8563
rect 432 8529 470 8563
rect 504 8529 542 8563
rect 576 8529 742 8563
rect 776 8529 814 8563
rect 848 8529 886 8563
rect 920 8529 1004 8563
rect -30 8517 1004 8529
rect -4500 8300 -4380 8320
rect -4120 8300 -3880 8320
rect -3620 8300 -3380 8320
rect -3120 8300 -2880 8320
rect -2620 8300 -2380 8320
rect -2120 8300 -2000 8320
rect -4500 8100 -2000 8300
rect -4500 8080 -4380 8100
rect -4120 8080 -3880 8100
rect -3620 8080 -3380 8100
rect -3120 8080 -2880 8100
rect -2620 8080 -2380 8100
rect -2120 8080 -2000 8100
rect -4500 7820 -4400 8080
rect -4100 7820 -3900 8080
rect -3600 7820 -3400 8080
rect -3100 7820 -2900 8080
rect -2600 7820 -2400 8080
rect -2100 7820 -2000 8080
rect -4500 7800 -4380 7820
rect -4120 7800 -3880 7820
rect -3620 7800 -3380 7820
rect -3120 7800 -2880 7820
rect -2620 7800 -2380 7820
rect -2120 7800 -2000 7820
rect -4800 7700 -2000 7800
rect -1560 8490 -150 8500
rect 1100 8490 1800 8500
rect -1560 8480 -124 8490
rect -55 8480 -3 8483
rect -2500 7680 -1800 7700
rect -2500 7600 -1980 7680
rect -2500 7580 -2380 7600
rect -2120 7580 -1980 7600
rect -2500 7320 -2400 7580
rect -2100 7520 -1980 7580
rect -1820 7520 -1800 7680
rect -2100 7500 -1800 7520
rect -2100 7400 -2000 7500
rect -1560 7400 -1540 8480
rect -2100 7360 -1540 7400
rect -1420 8454 -124 8480
rect -1420 8420 -174 8454
rect -140 8420 -124 8454
rect -1420 8400 -124 8420
rect -1420 8300 -1400 8400
rect -700 8374 -124 8400
rect -700 8340 -174 8374
rect -140 8340 -124 8374
rect -700 8300 -124 8340
rect -1420 8294 -124 8300
rect -1420 8260 -174 8294
rect -140 8260 -124 8294
rect -1420 8214 -124 8260
rect -1420 8200 -174 8214
rect -1420 8100 -1400 8200
rect -700 8180 -174 8200
rect -140 8180 -124 8214
rect -700 8134 -124 8180
rect -700 8100 -174 8134
rect -140 8100 -124 8134
rect -1420 8054 -124 8100
rect -1420 8020 -174 8054
rect -140 8020 -124 8054
rect -1420 8000 -124 8020
rect -1420 7900 -1400 8000
rect -700 7974 -124 8000
rect -700 7940 -174 7974
rect -140 7940 -124 7974
rect -700 7900 -124 7940
rect -1420 7894 -124 7900
rect -1420 7860 -174 7894
rect -140 7860 -124 7894
rect -1420 7814 -124 7860
rect -1420 7800 -174 7814
rect -1420 7700 -1400 7800
rect -700 7780 -174 7800
rect -140 7780 -124 7814
rect -700 7734 -124 7780
rect -700 7700 -174 7734
rect -140 7700 -124 7734
rect -1420 7654 -124 7700
rect -1420 7620 -174 7654
rect -140 7620 -124 7654
rect -1420 7600 -124 7620
rect -1420 7500 -1400 7600
rect -700 7574 -124 7600
rect -700 7540 -174 7574
rect -140 7540 -124 7574
rect -700 7500 -124 7540
rect -1420 7494 -124 7500
rect -1420 7460 -174 7494
rect -140 7460 -124 7494
rect -1420 7400 -124 7460
rect -1420 7360 -1240 7400
rect -2100 7320 -1240 7360
rect -194 7330 -124 7400
rect -57 8471 -3 8480
rect -57 8437 -46 8471
rect -12 8437 -3 8471
rect -57 8399 -3 8437
rect -57 8365 -46 8399
rect -12 8365 -3 8399
rect -57 8327 -3 8365
rect -57 8293 -46 8327
rect -12 8293 -3 8327
rect -57 8255 -3 8293
rect -57 8221 -46 8255
rect -12 8221 -3 8255
rect -57 8183 -3 8221
rect -57 8149 -46 8183
rect -12 8149 -3 8183
rect -57 8111 -3 8149
rect -57 8077 -46 8111
rect -12 8077 -3 8111
rect -57 8039 -3 8077
rect -57 8005 -46 8039
rect -12 8005 -3 8039
rect -57 7967 -3 8005
rect -57 7933 -46 7967
rect -12 7933 -3 7967
rect -57 7895 -3 7933
rect -57 7861 -46 7895
rect -12 7861 -3 7895
rect -57 7823 -3 7861
rect -57 7789 -46 7823
rect -12 7789 -3 7823
rect -57 7751 -3 7789
rect -57 7717 -46 7751
rect -12 7717 -3 7751
rect -57 7679 -3 7717
rect -57 7645 -46 7679
rect -12 7645 -3 7679
rect -57 7607 -3 7645
rect -57 7573 -46 7607
rect -12 7573 -3 7607
rect -57 7535 -3 7573
rect -57 7501 -46 7535
rect -12 7501 -3 7535
rect -57 7400 -3 7501
rect 31 8471 83 8483
rect 31 8437 40 8471
rect 74 8437 83 8471
rect 31 8411 83 8437
rect 31 8331 83 8359
rect 31 8255 83 8279
rect 31 8251 40 8255
rect 74 8251 83 8255
rect 31 8183 83 8199
rect 31 8171 40 8183
rect 74 8171 83 8183
rect 31 8111 83 8119
rect 31 8091 40 8111
rect 74 8091 83 8111
rect 31 8011 40 8039
rect 74 8011 83 8039
rect 31 7933 40 7959
rect 74 7933 83 7959
rect 31 7931 83 7933
rect 31 7861 40 7879
rect 74 7861 83 7879
rect 31 7851 83 7861
rect 31 7789 40 7799
rect 74 7789 83 7799
rect 31 7771 83 7789
rect 31 7717 40 7719
rect 74 7717 83 7719
rect 31 7691 83 7717
rect 31 7611 83 7639
rect 31 7535 83 7559
rect 31 7501 40 7535
rect 74 7501 83 7535
rect 31 7489 83 7501
rect 117 8471 169 8483
rect 117 8437 126 8471
rect 160 8437 169 8471
rect 117 8399 169 8437
rect 117 8365 126 8399
rect 160 8365 169 8399
rect 117 8327 169 8365
rect 117 8293 126 8327
rect 160 8293 169 8327
rect 117 8255 169 8293
rect 117 8221 126 8255
rect 160 8221 169 8255
rect 117 8183 169 8221
rect 117 8149 126 8183
rect 160 8149 169 8183
rect 117 8111 169 8149
rect 117 8077 126 8111
rect 160 8077 169 8111
rect 117 8039 169 8077
rect 117 8005 126 8039
rect 160 8005 169 8039
rect 117 7967 169 8005
rect 117 7933 126 7967
rect 160 7933 169 7967
rect 117 7895 169 7933
rect 117 7861 126 7895
rect 160 7861 169 7895
rect 117 7823 169 7861
rect 117 7789 126 7823
rect 160 7789 169 7823
rect 117 7751 169 7789
rect 117 7717 126 7751
rect 160 7717 169 7751
rect 117 7679 169 7717
rect 117 7645 126 7679
rect 160 7645 169 7679
rect 117 7607 169 7645
rect 117 7573 126 7607
rect 160 7573 169 7607
rect 117 7535 169 7573
rect 117 7501 126 7535
rect 160 7501 169 7535
rect 117 7400 169 7501
rect 203 8471 255 8483
rect 203 8437 212 8471
rect 246 8437 255 8471
rect 203 8411 255 8437
rect 203 8331 255 8359
rect 203 8255 255 8279
rect 203 8251 212 8255
rect 246 8251 255 8255
rect 203 8183 255 8199
rect 203 8171 212 8183
rect 246 8171 255 8183
rect 203 8111 255 8119
rect 203 8091 212 8111
rect 246 8091 255 8111
rect 203 8011 212 8039
rect 246 8011 255 8039
rect 203 7933 212 7959
rect 246 7933 255 7959
rect 203 7931 255 7933
rect 203 7861 212 7879
rect 246 7861 255 7879
rect 203 7851 255 7861
rect 203 7789 212 7799
rect 246 7789 255 7799
rect 203 7771 255 7789
rect 203 7717 212 7719
rect 246 7717 255 7719
rect 203 7691 255 7717
rect 203 7611 255 7639
rect 203 7535 255 7559
rect 203 7501 212 7535
rect 246 7501 255 7535
rect 203 7489 255 7501
rect 289 8471 341 8483
rect 289 8437 298 8471
rect 332 8437 341 8471
rect 289 8399 341 8437
rect 289 8365 298 8399
rect 332 8365 341 8399
rect 289 8327 341 8365
rect 289 8293 298 8327
rect 332 8293 341 8327
rect 289 8255 341 8293
rect 289 8221 298 8255
rect 332 8221 341 8255
rect 289 8183 341 8221
rect 289 8149 298 8183
rect 332 8149 341 8183
rect 289 8111 341 8149
rect 289 8077 298 8111
rect 332 8077 341 8111
rect 289 8039 341 8077
rect 289 8005 298 8039
rect 332 8005 341 8039
rect 289 7967 341 8005
rect 289 7933 298 7967
rect 332 7933 341 7967
rect 289 7895 341 7933
rect 289 7861 298 7895
rect 332 7861 341 7895
rect 289 7823 341 7861
rect 289 7789 298 7823
rect 332 7789 341 7823
rect 289 7751 341 7789
rect 289 7717 298 7751
rect 332 7717 341 7751
rect 289 7679 341 7717
rect 289 7645 298 7679
rect 332 7645 341 7679
rect 289 7607 341 7645
rect 289 7573 298 7607
rect 332 7573 341 7607
rect 289 7535 341 7573
rect 289 7501 298 7535
rect 332 7501 341 7535
rect 289 7400 341 7501
rect 375 8471 427 8483
rect 375 8437 384 8471
rect 418 8437 427 8471
rect 375 8411 427 8437
rect 375 8331 427 8359
rect 375 8255 427 8279
rect 375 8251 384 8255
rect 418 8251 427 8255
rect 375 8183 427 8199
rect 375 8171 384 8183
rect 418 8171 427 8183
rect 375 8111 427 8119
rect 375 8091 384 8111
rect 418 8091 427 8111
rect 375 8011 384 8039
rect 418 8011 427 8039
rect 375 7933 384 7959
rect 418 7933 427 7959
rect 375 7931 427 7933
rect 375 7861 384 7879
rect 418 7861 427 7879
rect 375 7851 427 7861
rect 375 7789 384 7799
rect 418 7789 427 7799
rect 375 7771 427 7789
rect 375 7717 384 7719
rect 418 7717 427 7719
rect 375 7691 427 7717
rect 375 7611 427 7639
rect 375 7535 427 7559
rect 375 7501 384 7535
rect 418 7501 427 7535
rect 375 7489 427 7501
rect 461 8471 513 8483
rect 461 8437 470 8471
rect 504 8437 513 8471
rect 461 8399 513 8437
rect 461 8365 470 8399
rect 504 8365 513 8399
rect 461 8327 513 8365
rect 461 8293 470 8327
rect 504 8293 513 8327
rect 461 8255 513 8293
rect 461 8221 470 8255
rect 504 8221 513 8255
rect 461 8183 513 8221
rect 461 8149 470 8183
rect 504 8149 513 8183
rect 461 8111 513 8149
rect 461 8077 470 8111
rect 504 8077 513 8111
rect 461 8039 513 8077
rect 461 8005 470 8039
rect 504 8005 513 8039
rect 461 7967 513 8005
rect 461 7933 470 7967
rect 504 7933 513 7967
rect 461 7895 513 7933
rect 461 7861 470 7895
rect 504 7861 513 7895
rect 461 7823 513 7861
rect 461 7789 470 7823
rect 504 7789 513 7823
rect 461 7751 513 7789
rect 461 7717 470 7751
rect 504 7717 513 7751
rect 461 7679 513 7717
rect 461 7645 470 7679
rect 504 7645 513 7679
rect 461 7607 513 7645
rect 461 7573 470 7607
rect 504 7573 513 7607
rect 461 7535 513 7573
rect 461 7501 470 7535
rect 504 7501 513 7535
rect 461 7400 513 7501
rect 547 8471 599 8483
rect 547 8437 556 8471
rect 590 8437 599 8471
rect 547 8411 599 8437
rect 547 8331 599 8359
rect 547 8255 599 8279
rect 547 8251 556 8255
rect 590 8251 599 8255
rect 547 8183 599 8199
rect 547 8171 556 8183
rect 590 8171 599 8183
rect 547 8111 599 8119
rect 547 8091 556 8111
rect 590 8091 599 8111
rect 547 8011 556 8039
rect 590 8011 599 8039
rect 547 7933 556 7959
rect 590 7933 599 7959
rect 547 7931 599 7933
rect 547 7861 556 7879
rect 590 7861 599 7879
rect 547 7851 599 7861
rect 547 7789 556 7799
rect 590 7789 599 7799
rect 547 7771 599 7789
rect 547 7717 556 7719
rect 590 7717 599 7719
rect 547 7691 599 7717
rect 547 7611 599 7639
rect 547 7535 599 7559
rect 547 7501 556 7535
rect 590 7501 599 7535
rect 547 7489 599 7501
rect 633 8471 685 8483
rect 633 8437 642 8471
rect 676 8437 685 8471
rect 633 8399 685 8437
rect 633 8365 642 8399
rect 676 8365 685 8399
rect 633 8327 685 8365
rect 633 8293 642 8327
rect 676 8293 685 8327
rect 633 8255 685 8293
rect 633 8221 642 8255
rect 676 8221 685 8255
rect 633 8183 685 8221
rect 633 8149 642 8183
rect 676 8149 685 8183
rect 633 8111 685 8149
rect 633 8077 642 8111
rect 676 8077 685 8111
rect 633 8039 685 8077
rect 633 8005 642 8039
rect 676 8005 685 8039
rect 633 7967 685 8005
rect 633 7933 642 7967
rect 676 7933 685 7967
rect 633 7895 685 7933
rect 633 7861 642 7895
rect 676 7861 685 7895
rect 633 7823 685 7861
rect 633 7789 642 7823
rect 676 7789 685 7823
rect 633 7751 685 7789
rect 633 7717 642 7751
rect 676 7717 685 7751
rect 633 7679 685 7717
rect 633 7645 642 7679
rect 676 7645 685 7679
rect 633 7607 685 7645
rect 633 7573 642 7607
rect 676 7573 685 7607
rect 633 7535 685 7573
rect 633 7501 642 7535
rect 676 7501 685 7535
rect 633 7400 685 7501
rect 719 8471 771 8483
rect 719 8437 728 8471
rect 762 8437 771 8471
rect 719 8411 771 8437
rect 719 8331 771 8359
rect 719 8255 771 8279
rect 719 8251 728 8255
rect 762 8251 771 8255
rect 719 8183 771 8199
rect 719 8171 728 8183
rect 762 8171 771 8183
rect 719 8111 771 8119
rect 719 8091 728 8111
rect 762 8091 771 8111
rect 719 8011 728 8039
rect 762 8011 771 8039
rect 719 7933 728 7959
rect 762 7933 771 7959
rect 719 7931 771 7933
rect 719 7861 728 7879
rect 762 7861 771 7879
rect 719 7851 771 7861
rect 719 7789 728 7799
rect 762 7789 771 7799
rect 719 7771 771 7789
rect 719 7717 728 7719
rect 762 7717 771 7719
rect 719 7691 771 7717
rect 719 7611 771 7639
rect 719 7535 771 7559
rect 719 7501 728 7535
rect 762 7501 771 7535
rect 719 7489 771 7501
rect 805 8471 857 8483
rect 805 8437 814 8471
rect 848 8437 857 8471
rect 805 8399 857 8437
rect 805 8365 814 8399
rect 848 8365 857 8399
rect 805 8327 857 8365
rect 805 8293 814 8327
rect 848 8293 857 8327
rect 805 8255 857 8293
rect 805 8221 814 8255
rect 848 8221 857 8255
rect 805 8183 857 8221
rect 805 8149 814 8183
rect 848 8149 857 8183
rect 805 8111 857 8149
rect 805 8077 814 8111
rect 848 8077 857 8111
rect 805 8039 857 8077
rect 805 8005 814 8039
rect 848 8005 857 8039
rect 805 7967 857 8005
rect 805 7933 814 7967
rect 848 7933 857 7967
rect 805 7895 857 7933
rect 805 7861 814 7895
rect 848 7861 857 7895
rect 805 7823 857 7861
rect 805 7789 814 7823
rect 848 7789 857 7823
rect 805 7751 857 7789
rect 805 7717 814 7751
rect 848 7717 857 7751
rect 805 7679 857 7717
rect 805 7645 814 7679
rect 848 7645 857 7679
rect 805 7607 857 7645
rect 805 7573 814 7607
rect 848 7573 857 7607
rect 805 7535 857 7573
rect 805 7501 814 7535
rect 848 7501 857 7535
rect 805 7400 857 7501
rect 891 8471 943 8483
rect 891 8437 900 8471
rect 934 8437 943 8471
rect 891 8411 943 8437
rect 891 8331 943 8359
rect 891 8255 943 8279
rect 891 8251 900 8255
rect 934 8251 943 8255
rect 891 8183 943 8199
rect 891 8171 900 8183
rect 934 8171 943 8183
rect 891 8111 943 8119
rect 891 8091 900 8111
rect 934 8091 943 8111
rect 891 8011 900 8039
rect 934 8011 943 8039
rect 891 7933 900 7959
rect 934 7933 943 7959
rect 891 7931 943 7933
rect 891 7861 900 7879
rect 934 7861 943 7879
rect 891 7851 943 7861
rect 891 7789 900 7799
rect 934 7789 943 7799
rect 891 7771 943 7789
rect 891 7717 900 7719
rect 934 7717 943 7719
rect 891 7691 943 7717
rect 891 7611 943 7639
rect 891 7535 943 7559
rect 891 7501 900 7535
rect 934 7501 943 7535
rect 891 7489 943 7501
rect 977 8480 1029 8483
rect 977 8471 1031 8480
rect 977 8437 986 8471
rect 1020 8437 1031 8471
rect 977 8399 1031 8437
rect 977 8365 986 8399
rect 1020 8365 1031 8399
rect 977 8327 1031 8365
rect 977 8293 986 8327
rect 1020 8293 1031 8327
rect 977 8255 1031 8293
rect 977 8221 986 8255
rect 1020 8221 1031 8255
rect 977 8183 1031 8221
rect 977 8149 986 8183
rect 1020 8149 1031 8183
rect 977 8111 1031 8149
rect 977 8077 986 8111
rect 1020 8077 1031 8111
rect 977 8039 1031 8077
rect 977 8005 986 8039
rect 1020 8005 1031 8039
rect 977 7967 1031 8005
rect 977 7933 986 7967
rect 1020 7933 1031 7967
rect 977 7895 1031 7933
rect 977 7861 986 7895
rect 1020 7861 1031 7895
rect 977 7823 1031 7861
rect 977 7789 986 7823
rect 1020 7789 1031 7823
rect 977 7751 1031 7789
rect 977 7717 986 7751
rect 1020 7717 1031 7751
rect 977 7679 1031 7717
rect 977 7645 986 7679
rect 1020 7645 1031 7679
rect 977 7607 1031 7645
rect 977 7573 986 7607
rect 1020 7573 1031 7607
rect 977 7535 1031 7573
rect 977 7501 986 7535
rect 1020 7501 1031 7535
rect 977 7400 1031 7501
rect -57 7330 -14 7400
rect -2500 7300 -2380 7320
rect -2120 7300 -1240 7320
rect -184 7310 -124 7330
rect -34 7300 -14 7330
rect 996 7330 1031 7400
rect 1096 8454 1800 8490
rect 1096 8420 1116 8454
rect 1150 8420 1800 8454
rect 1096 8374 1800 8420
rect 1096 8340 1116 8374
rect 1150 8340 1800 8374
rect 1096 8294 1800 8340
rect 1096 8260 1116 8294
rect 1150 8260 1800 8294
rect 1096 8214 1800 8260
rect 1096 8180 1116 8214
rect 1150 8180 1800 8214
rect 1096 8134 1800 8180
rect 1096 8100 1116 8134
rect 1150 8100 1800 8134
rect 1096 8054 1800 8100
rect 1096 8020 1116 8054
rect 1150 8020 1800 8054
rect 1096 7974 1800 8020
rect 1096 7940 1116 7974
rect 1150 7940 1800 7974
rect 1096 7894 1800 7940
rect 1096 7860 1116 7894
rect 1150 7860 1800 7894
rect 1096 7814 1800 7860
rect 1096 7780 1116 7814
rect 1150 7780 1800 7814
rect 1096 7734 1800 7780
rect 1096 7700 1116 7734
rect 1150 7700 1800 7734
rect 1096 7654 1800 7700
rect 1096 7620 1116 7654
rect 1150 7620 1800 7654
rect 1096 7574 1800 7620
rect 1096 7540 1116 7574
rect 1150 7540 1800 7574
rect 1096 7494 1800 7540
rect 1096 7460 1116 7494
rect 1150 7460 1800 7494
rect 1096 7330 1800 7460
rect 996 7300 1016 7330
rect -2500 7180 -1240 7300
rect -2500 7110 -2350 7180
rect -2150 7110 -1850 7180
rect -1650 7110 -1240 7180
rect -2500 7100 -1240 7110
rect -2500 7080 -2380 7100
rect -2120 7080 -1880 7100
rect -1620 7080 -1240 7100
rect -2500 7050 -2400 7080
rect -2500 6850 -2480 7050
rect -2410 6850 -2400 7050
rect -2500 6820 -2400 6850
rect -2100 7050 -1900 7080
rect -2100 6850 -2090 7050
rect -2020 6850 -1980 7050
rect -1910 6850 -1900 7050
rect -2100 6820 -1900 6850
rect -1600 7060 -1240 7080
rect -1600 7050 -1380 7060
rect -1600 6850 -1590 7050
rect -1520 6850 -1380 7050
rect -1600 6820 -1380 6850
rect -2500 6800 -2380 6820
rect -2120 6800 -1880 6820
rect -1620 6800 -1380 6820
rect -2500 6790 -1380 6800
rect -2500 6720 -2350 6790
rect -2150 6720 -1850 6790
rect -1650 6720 -1380 6790
rect -2500 6680 -1380 6720
rect -2500 6610 -2350 6680
rect -2150 6610 -1850 6680
rect -1650 6610 -1380 6680
rect -2500 6600 -1380 6610
rect -2500 6580 -2380 6600
rect -2120 6580 -1880 6600
rect -1620 6580 -1380 6600
rect -2500 6550 -2400 6580
rect -2500 6350 -2480 6550
rect -2410 6350 -2400 6550
rect -2500 6320 -2400 6350
rect -2100 6550 -1900 6580
rect -2100 6350 -2090 6550
rect -2020 6350 -1980 6550
rect -1910 6350 -1900 6550
rect -2100 6320 -1900 6350
rect -1600 6550 -1380 6580
rect -1600 6350 -1590 6550
rect -1520 6350 -1380 6550
rect -1600 6320 -1380 6350
rect -2500 6300 -2380 6320
rect -2120 6300 -1880 6320
rect -1620 6300 -1380 6320
rect -2500 6290 -1380 6300
rect -2500 6220 -2350 6290
rect -2150 6220 -1850 6290
rect -1650 6220 -1380 6290
rect -2500 6200 -1380 6220
rect -4000 6180 -1380 6200
rect -4000 6110 -3850 6180
rect -3650 6110 -3350 6180
rect -3150 6110 -2850 6180
rect -2650 6110 -2350 6180
rect -2150 6110 -1850 6180
rect -1650 6110 -1380 6180
rect -4000 6100 -1380 6110
rect -4000 6080 -3880 6100
rect -3620 6080 -3380 6100
rect -3120 6080 -2880 6100
rect -2620 6080 -2380 6100
rect -2120 6080 -1880 6100
rect -1620 6080 -1380 6100
rect -4000 6050 -3900 6080
rect -4000 5850 -3980 6050
rect -3910 5850 -3900 6050
rect -4000 5820 -3900 5850
rect -3600 6050 -3400 6080
rect -3600 5850 -3590 6050
rect -3520 5850 -3480 6050
rect -3410 5850 -3400 6050
rect -3600 5820 -3400 5850
rect -3100 6050 -2900 6080
rect -3100 5850 -3090 6050
rect -3020 5850 -2980 6050
rect -2910 5850 -2900 6050
rect -3100 5820 -2900 5850
rect -2600 6050 -2400 6080
rect -2600 5850 -2590 6050
rect -2520 5850 -2480 6050
rect -2410 5850 -2400 6050
rect -2600 5820 -2400 5850
rect -2100 6050 -1900 6080
rect -2100 5850 -2090 6050
rect -2020 5850 -1980 6050
rect -1910 5850 -1900 6050
rect -2100 5820 -1900 5850
rect -1600 6050 -1380 6080
rect -1600 5850 -1590 6050
rect -1520 5850 -1380 6050
rect -1600 5820 -1380 5850
rect -4000 5800 -3880 5820
rect -3620 5800 -3380 5820
rect -3120 5800 -2880 5820
rect -2620 5800 -2380 5820
rect -2120 5800 -1880 5820
rect -1620 5800 -1380 5820
rect -4000 5790 -1380 5800
rect -4000 5720 -3850 5790
rect -3650 5720 -3350 5790
rect -3150 5720 -2850 5790
rect -2650 5720 -2350 5790
rect -2150 5720 -1850 5790
rect -1650 5720 -1380 5790
rect -4000 5700 -1380 5720
rect -1260 5700 -1240 7060
rect -1000 7020 -800 7040
rect -1000 6860 -980 7020
rect -820 6860 -800 7020
rect -1000 6840 -800 6860
rect 1100 6700 1800 7330
rect 1100 6680 1320 6700
rect 1580 6680 1800 6700
rect 1100 6420 1300 6680
rect 1600 6420 1800 6680
rect 1100 6400 1320 6420
rect 1580 6400 1800 6420
rect 1100 6200 1800 6400
rect 1100 6180 1320 6200
rect 1580 6180 1800 6200
rect -1200 5920 -1000 5940
rect -1200 5760 -1180 5920
rect -1020 5760 -1000 5920
rect 1100 5920 1300 6180
rect 1600 5920 1800 6180
rect 1100 5900 1320 5920
rect 1580 5900 1800 5920
rect 1100 5800 1800 5900
rect -1200 5740 -1000 5760
rect 500 5700 2500 5800
rect -4000 5680 -500 5700
rect -4000 5610 -3850 5680
rect -3650 5610 -3350 5680
rect -3150 5610 -2850 5680
rect -2650 5610 -2350 5680
rect -2150 5610 -500 5680
rect -4000 5600 -500 5610
rect -4000 5580 -3880 5600
rect -3620 5580 -3380 5600
rect -3120 5580 -2880 5600
rect -2620 5580 -2380 5600
rect -2120 5580 -1880 5600
rect -1620 5580 -1380 5600
rect -1120 5580 -880 5600
rect -620 5580 -500 5600
rect -4000 5550 -3900 5580
rect -4000 5350 -3980 5550
rect -3910 5350 -3900 5550
rect -4000 5320 -3900 5350
rect -3600 5550 -3400 5580
rect -3600 5350 -3590 5550
rect -3520 5350 -3480 5550
rect -3410 5350 -3400 5550
rect -3600 5320 -3400 5350
rect -3100 5550 -2900 5580
rect -3100 5350 -3090 5550
rect -3020 5350 -2980 5550
rect -2910 5350 -2900 5550
rect -3100 5320 -2900 5350
rect -2600 5550 -2400 5580
rect -2600 5350 -2590 5550
rect -2520 5350 -2480 5550
rect -2410 5350 -2400 5550
rect -2600 5320 -2400 5350
rect -2100 5550 -1900 5580
rect -2100 5350 -2090 5550
rect -2020 5350 -1900 5550
rect -2100 5320 -1900 5350
rect -1600 5320 -1400 5580
rect -1100 5320 -900 5580
rect -600 5320 -500 5580
rect -4000 5300 -3880 5320
rect -3620 5300 -3380 5320
rect -3120 5300 -2880 5320
rect -2620 5300 -2380 5320
rect -2120 5300 -1880 5320
rect -1620 5300 -1380 5320
rect -1120 5300 -880 5320
rect -620 5300 -500 5320
rect -4000 5290 -500 5300
rect -4000 5220 -3850 5290
rect -3650 5220 -3350 5290
rect -3150 5220 -2850 5290
rect -2650 5220 -2350 5290
rect -2150 5220 -500 5290
rect -4000 5200 -500 5220
rect 500 5680 620 5700
rect 880 5680 1120 5700
rect 1380 5680 1620 5700
rect 1880 5680 2120 5700
rect 2380 5680 2500 5700
rect 500 5420 600 5680
rect 900 5420 1100 5680
rect 1400 5420 1600 5680
rect 1900 5420 2100 5680
rect 2400 5420 2500 5680
rect 500 5400 620 5420
rect 880 5400 1120 5420
rect 1380 5400 1620 5420
rect 1880 5400 2120 5420
rect 2380 5400 2500 5420
rect 500 5200 2500 5400
rect -5500 5100 -3500 5200
rect -5500 5080 -5380 5100
rect -5120 5080 -4880 5100
rect -4620 5080 -4380 5100
rect -4120 5080 -3880 5100
rect -3620 5080 -3500 5100
rect -5500 4820 -5400 5080
rect -5100 4820 -4900 5080
rect -4600 4820 -4400 5080
rect -4100 4820 -3900 5080
rect -3600 4820 -3500 5080
rect -5500 4800 -5380 4820
rect -5120 4800 -4880 4820
rect -4620 4800 -4380 4820
rect -4120 4800 -3880 4820
rect -3620 4800 -3500 4820
rect -5500 4600 -3500 4800
rect -5500 4580 -5380 4600
rect -5120 4580 -4880 4600
rect -4620 4580 -4380 4600
rect -4120 4580 -3880 4600
rect -3620 4580 -3500 4600
rect -5500 4320 -5400 4580
rect -5100 4320 -4900 4580
rect -4600 4320 -4400 4580
rect -4100 4320 -3900 4580
rect -3600 4320 -3500 4580
rect -5500 4300 -5380 4320
rect -5120 4300 -4880 4320
rect -4620 4300 -4380 4320
rect -4120 4300 -3880 4320
rect -3620 4300 -3500 4320
rect -5500 4100 -3500 4300
rect -5500 4080 -5380 4100
rect -5120 4080 -4880 4100
rect -4620 4080 -4380 4100
rect -4120 4080 -3880 4100
rect -3620 4080 -3500 4100
rect -5500 3820 -5400 4080
rect -5100 3820 -4900 4080
rect -4600 3820 -4400 4080
rect -4100 3820 -3900 4080
rect -3600 3820 -3500 4080
rect -5500 3800 -5380 3820
rect -5120 3800 -4880 3820
rect -4620 3800 -4380 3820
rect -4120 3800 -3880 3820
rect -3620 3800 -3500 3820
rect 500 5180 620 5200
rect 880 5180 1120 5200
rect 1380 5180 1620 5200
rect 1880 5180 2120 5200
rect 2380 5180 2500 5200
rect 500 4920 600 5180
rect 900 4920 1100 5180
rect 1400 4920 1600 5180
rect 1900 4920 2100 5180
rect 2400 4920 2500 5180
rect 500 4900 620 4920
rect 880 4900 1120 4920
rect 1380 4900 1620 4920
rect 1880 4900 2120 4920
rect 2380 4900 2500 4920
rect 500 4700 2500 4900
rect 500 4680 620 4700
rect 880 4680 1120 4700
rect 1380 4680 1620 4700
rect 1880 4680 2120 4700
rect 2380 4680 2500 4700
rect 500 4420 600 4680
rect 900 4420 1100 4680
rect 1400 4420 1600 4680
rect 1900 4420 2100 4680
rect 2400 4420 2500 4680
rect 500 4400 620 4420
rect 880 4400 1120 4420
rect 1380 4400 1620 4420
rect 1880 4400 2120 4420
rect 2380 4400 2500 4420
rect 500 4200 2500 4400
rect 500 4180 620 4200
rect 880 4180 1120 4200
rect 1380 4180 1620 4200
rect 1880 4180 2120 4200
rect 2380 4180 2500 4200
rect 500 3920 600 4180
rect 900 3920 1100 4180
rect 1400 3920 1600 4180
rect 1900 3920 2100 4180
rect 2400 3920 2500 4180
rect 500 3900 620 3920
rect 880 3900 1120 3920
rect 1380 3900 1620 3920
rect 1880 3900 2120 3920
rect 2380 3900 2500 3920
rect 500 3800 2500 3900
rect -5500 3600 -3500 3800
rect -5500 3580 -5380 3600
rect -5120 3580 -4880 3600
rect -4620 3580 -4380 3600
rect -4120 3580 -3880 3600
rect -3620 3580 -3500 3600
rect -5500 3320 -5400 3580
rect -5100 3320 -4900 3580
rect -4600 3320 -4400 3580
rect -4100 3320 -3900 3580
rect -3600 3320 -3500 3580
rect -5500 3300 -5380 3320
rect -5120 3300 -4880 3320
rect -4620 3300 -4380 3320
rect -4120 3300 -3880 3320
rect -3620 3300 -3500 3320
rect -5500 3100 -3500 3300
rect -5500 3080 -5380 3100
rect -5120 3080 -4880 3100
rect -4620 3080 -4380 3100
rect -4120 3080 -3880 3100
rect -3620 3080 -3500 3100
rect -5500 2820 -5400 3080
rect -5100 2820 -4900 3080
rect -4600 2820 -4400 3080
rect -4100 2820 -3900 3080
rect -3600 2820 -3500 3080
rect -5500 2800 -5380 2820
rect -5120 2800 -4880 2820
rect -4620 2800 -4380 2820
rect -4120 2800 -3880 2820
rect -3620 2800 -3500 2820
rect -500 3700 2500 3800
rect -500 3680 -380 3700
rect -120 3680 120 3700
rect 380 3680 620 3700
rect 880 3680 1120 3700
rect 1380 3680 1620 3700
rect 1880 3680 2120 3700
rect 2380 3680 2500 3700
rect -500 3420 -400 3680
rect -100 3420 100 3680
rect 400 3420 600 3680
rect 900 3420 1100 3680
rect 1400 3420 1600 3680
rect 1900 3420 2100 3680
rect 2400 3420 2500 3680
rect -500 3400 -380 3420
rect -120 3400 120 3420
rect 380 3400 620 3420
rect 880 3400 1120 3420
rect 1380 3400 1620 3420
rect 1880 3400 2120 3420
rect 2380 3400 2500 3420
rect -500 3200 2500 3400
rect -500 3180 -380 3200
rect -120 3180 120 3200
rect 380 3180 620 3200
rect 880 3180 1120 3200
rect 1380 3180 1620 3200
rect 1880 3180 2120 3200
rect 2380 3180 2500 3200
rect -500 2920 -400 3180
rect -100 2920 100 3180
rect 400 2920 600 3180
rect 900 2920 1100 3180
rect 1400 2920 1600 3180
rect 1900 2920 2100 3180
rect 2400 2920 2500 3180
rect -500 2900 -380 2920
rect -120 2900 120 2920
rect 380 2900 620 2920
rect 880 2900 1120 2920
rect 1380 2900 1620 2920
rect 1880 2900 2120 2920
rect 2380 2900 2500 2920
rect -500 2800 2500 2900
rect -5500 2700 2500 2800
rect -5500 2680 -3380 2700
rect -3120 2680 -2880 2700
rect -2620 2680 -2380 2700
rect -2120 2680 -1880 2700
rect -1620 2680 -1380 2700
rect -1120 2680 -880 2700
rect -620 2680 -380 2700
rect -120 2680 120 2700
rect 380 2680 620 2700
rect 880 2680 1120 2700
rect 1380 2680 1620 2700
rect 1880 2680 2120 2700
rect 2380 2680 2500 2700
rect -5500 2600 -3400 2680
rect -5500 2580 -5380 2600
rect -5120 2580 -4880 2600
rect -4620 2580 -4380 2600
rect -4120 2580 -3880 2600
rect -3620 2580 -3400 2600
rect -5500 2320 -5400 2580
rect -5100 2320 -4900 2580
rect -4600 2320 -4400 2580
rect -4100 2320 -3900 2580
rect -3600 2420 -3400 2580
rect -3100 2420 -2900 2680
rect -2600 2420 -2400 2680
rect -2100 2420 -1900 2680
rect -1600 2420 -1400 2680
rect -1100 2420 -900 2680
rect -600 2420 -400 2680
rect -100 2420 100 2680
rect 400 2420 600 2680
rect 900 2420 1100 2680
rect 1400 2420 1600 2680
rect 1900 2420 2100 2680
rect 2400 2420 2500 2680
rect -3600 2400 -3380 2420
rect -3120 2400 -2880 2420
rect -2620 2400 -2380 2420
rect -2120 2400 -1880 2420
rect -1620 2400 -1380 2420
rect -1120 2400 -880 2420
rect -620 2400 -380 2420
rect -120 2400 120 2420
rect 380 2400 620 2420
rect 880 2400 1120 2420
rect 1380 2400 1620 2420
rect 1880 2400 2120 2420
rect 2380 2400 2500 2420
rect -3600 2320 2500 2400
rect -5500 2300 -5380 2320
rect -5120 2300 -4880 2320
rect -4620 2300 -4380 2320
rect -4120 2300 -3880 2320
rect -3620 2300 2500 2320
rect -5500 2200 2500 2300
rect -5500 2180 -3380 2200
rect -3120 2180 -2880 2200
rect -2620 2180 -2380 2200
rect -2120 2180 -1880 2200
rect -1620 2180 -1380 2200
rect -1120 2180 -880 2200
rect -620 2180 -380 2200
rect -120 2180 120 2200
rect 380 2180 620 2200
rect 880 2180 1120 2200
rect 1380 2180 1620 2200
rect 1880 2180 2120 2200
rect 2380 2180 2500 2200
rect -5500 2100 -3400 2180
rect -5500 2080 -5380 2100
rect -5120 2080 -4880 2100
rect -4620 2080 -4380 2100
rect -4120 2080 -3880 2100
rect -3620 2080 -3400 2100
rect -5500 1820 -5400 2080
rect -5100 1820 -4900 2080
rect -4600 1820 -4400 2080
rect -4100 1820 -3900 2080
rect -3600 1920 -3400 2080
rect -3100 1920 -2900 2180
rect -2600 1920 -2400 2180
rect -2100 1920 -1900 2180
rect -1600 1920 -1400 2180
rect -1100 1920 -900 2180
rect -600 1920 -400 2180
rect -100 1920 100 2180
rect 400 1920 600 2180
rect 900 1920 1100 2180
rect 1400 1920 1600 2180
rect 1900 1920 2100 2180
rect 2400 1920 2500 2180
rect -3600 1900 -3380 1920
rect -3120 1900 -2880 1920
rect -2620 1900 -2380 1920
rect -2120 1900 -1880 1920
rect -1620 1900 -1380 1920
rect -1120 1900 -880 1920
rect -620 1900 -380 1920
rect -120 1900 120 1920
rect 380 1900 620 1920
rect 880 1900 1120 1920
rect 1380 1900 1620 1920
rect 1880 1900 2120 1920
rect 2380 1900 2500 1920
rect -3600 1820 2500 1900
rect -5500 1800 -5380 1820
rect -5120 1800 -4880 1820
rect -4620 1800 -4380 1820
rect -4120 1800 -3880 1820
rect -3620 1800 2500 1820
rect -5500 1600 -3500 1800
rect -5500 1580 -5380 1600
rect -5120 1580 -4880 1600
rect -4620 1580 -4380 1600
rect -4120 1580 -3880 1600
rect -3620 1580 -3500 1600
rect -5500 1320 -5400 1580
rect -5100 1320 -4900 1580
rect -4600 1320 -4400 1580
rect -4100 1320 -3900 1580
rect -3600 1320 -3500 1580
rect -5500 1300 -5380 1320
rect -5120 1300 -4880 1320
rect -4620 1300 -4380 1320
rect -4120 1300 -3880 1320
rect -3620 1300 -3500 1320
rect -5500 1100 -3500 1300
rect -5500 1080 -5380 1100
rect -5120 1080 -4880 1100
rect -4620 1080 -4380 1100
rect -4120 1080 -3880 1100
rect -3620 1080 -3500 1100
rect -5500 820 -5400 1080
rect -5100 820 -4900 1080
rect -4600 820 -4400 1080
rect -4100 820 -3900 1080
rect -3600 820 -3500 1080
rect -5500 800 -5380 820
rect -5120 800 -4880 820
rect -4620 800 -4380 820
rect -4120 800 -3880 820
rect -3620 800 -3500 820
rect -5500 600 -3500 800
rect -5500 580 -5380 600
rect -5120 580 -4880 600
rect -4620 580 -4380 600
rect -4120 580 -3880 600
rect -3620 580 -3500 600
rect -5500 320 -5400 580
rect -5100 320 -4900 580
rect -4600 320 -4400 580
rect -4100 320 -3900 580
rect -3600 320 -3500 580
rect -5500 300 -5380 320
rect -5120 300 -4880 320
rect -4620 300 -4380 320
rect -4120 300 -3880 320
rect -3620 300 -3500 320
rect -700 1700 -200 1800
rect -700 1680 -580 1700
rect -320 1680 -200 1700
rect -700 1420 -600 1680
rect -300 1420 -200 1680
rect -700 1400 -580 1420
rect -320 1400 -200 1420
rect -700 1200 -200 1400
rect -700 1180 -580 1200
rect -320 1180 -200 1200
rect -700 920 -600 1180
rect -300 920 -200 1180
rect -700 900 -580 920
rect -320 900 -200 920
rect -700 700 -200 900
rect -700 680 -580 700
rect -320 680 -200 700
rect -700 420 -600 680
rect -300 420 -200 680
rect 1100 1700 1600 1800
rect 1100 1680 1220 1700
rect 1480 1680 1600 1700
rect 1100 1420 1200 1680
rect 1500 1420 1600 1680
rect 1100 1400 1220 1420
rect 1480 1400 1600 1420
rect 1100 1200 1600 1400
rect 1100 1180 1220 1200
rect 1480 1180 1600 1200
rect 1100 920 1200 1180
rect 1500 920 1600 1180
rect 1100 900 1220 920
rect 1480 900 1600 920
rect 1100 700 1600 900
rect 1100 680 1220 700
rect 1480 680 1600 700
rect -700 400 -580 420
rect -320 400 -200 420
rect -700 300 -200 400
rect 10 320 80 450
rect 150 431 170 460
rect 149 380 170 431
rect 870 450 890 460
rect 870 380 891 450
rect 149 370 891 380
rect 10 300 30 320
rect -5500 100 -3500 300
rect -750 286 30 300
rect 64 286 80 320
rect -750 240 80 286
rect -750 206 30 240
rect 64 206 80 240
rect -750 200 80 206
rect -5500 80 -5380 100
rect -5120 80 -4880 100
rect -4620 80 -4380 100
rect -4120 80 -3880 100
rect -3620 80 -3500 100
rect -5500 -180 -5400 80
rect -5100 -180 -4900 80
rect -4600 -180 -4400 80
rect -4100 -180 -3900 80
rect -3600 -180 -3500 80
rect -5500 -200 -5380 -180
rect -5120 -200 -4880 -180
rect -4620 -200 -4380 -180
rect -4120 -200 -3880 -180
rect -3620 -200 -3500 -180
rect -5500 -300 -3500 -200
rect -1500 160 80 200
rect -1500 126 30 160
rect 64 126 80 160
rect -1500 100 80 126
rect -1500 80 -1380 100
rect -1120 80 80 100
rect -1500 -180 -1400 80
rect -1100 46 30 80
rect 64 46 80 80
rect -1100 0 80 46
rect -1100 -34 30 0
rect 64 -34 80 0
rect -1100 -80 80 -34
rect -1100 -114 30 -80
rect 64 -114 80 -80
rect -1100 -160 80 -114
rect -1100 -180 30 -160
rect -1500 -200 -1380 -180
rect -1120 -194 30 -180
rect 64 -194 80 -160
rect -1120 -200 80 -194
rect -1500 -240 80 -200
rect -1500 -274 30 -240
rect 64 -274 80 -240
rect -5500 -400 -4500 -300
rect -5500 -420 -5380 -400
rect -5120 -420 -4880 -400
rect -4620 -420 -4500 -400
rect -5500 -680 -5400 -420
rect -5100 -680 -4900 -420
rect -4600 -600 -4500 -420
rect -1500 -320 80 -274
rect -1500 -354 30 -320
rect 64 -354 80 -320
rect -1500 -400 80 -354
rect -1500 -420 -1380 -400
rect -1120 -420 30 -400
rect -4600 -640 -4400 -600
rect -4600 -680 -4540 -640
rect -5500 -700 -5380 -680
rect -5120 -700 -4880 -680
rect -4620 -700 -4540 -680
rect -5500 -900 -4540 -700
rect -5500 -920 -5380 -900
rect -5120 -920 -4880 -900
rect -4620 -920 -4540 -900
rect -5500 -1180 -5400 -920
rect -5100 -1180 -4900 -920
rect -4600 -1180 -4540 -920
rect -5500 -1200 -5380 -1180
rect -5120 -1200 -4880 -1180
rect -4620 -1200 -4540 -1180
rect -14500 -1400 -10000 -1300
rect -14500 -1420 -14380 -1400
rect -14120 -1420 -13880 -1400
rect -13620 -1420 -13380 -1400
rect -13120 -1420 -12880 -1400
rect -12620 -1420 -12380 -1400
rect -12120 -1420 -11880 -1400
rect -11620 -1420 -11380 -1400
rect -11120 -1420 -10880 -1400
rect -10620 -1420 -10380 -1400
rect -10120 -1420 -10000 -1400
rect -14500 -1680 -14400 -1420
rect -14100 -1680 -13900 -1420
rect -13600 -1680 -13400 -1420
rect -13100 -1680 -12900 -1420
rect -12600 -1680 -12400 -1420
rect -12100 -1680 -11900 -1420
rect -11600 -1680 -11400 -1420
rect -11100 -1680 -10900 -1420
rect -10600 -1680 -10400 -1420
rect -10100 -1680 -10000 -1420
rect -14500 -1700 -14380 -1680
rect -14120 -1700 -13880 -1680
rect -13620 -1700 -13380 -1680
rect -13120 -1700 -12880 -1680
rect -12620 -1700 -12380 -1680
rect -12120 -1700 -11880 -1680
rect -11620 -1700 -11380 -1680
rect -11120 -1700 -10880 -1680
rect -10620 -1700 -10380 -1680
rect -10120 -1700 -10000 -1680
rect -14500 -1900 -11600 -1700
rect -11400 -1900 -10000 -1700
rect -14500 -1920 -14380 -1900
rect -14120 -1920 -13880 -1900
rect -13620 -1920 -13380 -1900
rect -13120 -1920 -12880 -1900
rect -12620 -1920 -12380 -1900
rect -12120 -1920 -11880 -1900
rect -11620 -1920 -11380 -1900
rect -11120 -1920 -10880 -1900
rect -10620 -1920 -10380 -1900
rect -10120 -1920 -10000 -1900
rect -14500 -2180 -14400 -1920
rect -14100 -2180 -13900 -1920
rect -13600 -2180 -13400 -1920
rect -13100 -2180 -12900 -1920
rect -12600 -2180 -12400 -1920
rect -12100 -2180 -11900 -1920
rect -11600 -2180 -11400 -1920
rect -11100 -2180 -10900 -1920
rect -10600 -2180 -10400 -1920
rect -10100 -2180 -10000 -1920
rect -14500 -2200 -14380 -2180
rect -14120 -2200 -13880 -2180
rect -13620 -2200 -13380 -2180
rect -13120 -2200 -12880 -2180
rect -12620 -2200 -12380 -2180
rect -12120 -2200 -11880 -2180
rect -11620 -2200 -11380 -2180
rect -11120 -2200 -10880 -2180
rect -10620 -2200 -10380 -2180
rect -10120 -2200 -10000 -2180
rect -14500 -2400 -11600 -2200
rect -11400 -2300 -10000 -2200
rect -5500 -1400 -4540 -1200
rect -5500 -1420 -5380 -1400
rect -5120 -1420 -4880 -1400
rect -4620 -1420 -4540 -1400
rect -5500 -1680 -5400 -1420
rect -5100 -1680 -4900 -1420
rect -4600 -1680 -4540 -1420
rect -5500 -1700 -5380 -1680
rect -5120 -1700 -4880 -1680
rect -4620 -1700 -4540 -1680
rect -5500 -1900 -4540 -1700
rect -5500 -1920 -5380 -1900
rect -5120 -1920 -4880 -1900
rect -4620 -1920 -4540 -1900
rect -5500 -2180 -5400 -1920
rect -5100 -2180 -4900 -1920
rect -4600 -2180 -4540 -1920
rect -4420 -2000 -4400 -640
rect -4320 -690 -4120 -670
rect -4320 -890 -4300 -690
rect -4140 -890 -4120 -690
rect -4320 -910 -4120 -890
rect -3980 -690 -3780 -670
rect -3980 -890 -3960 -690
rect -3800 -890 -3780 -690
rect -3980 -910 -3780 -890
rect -1500 -680 -1400 -420
rect -1100 -434 30 -420
rect 64 -434 80 -400
rect -1100 -480 80 -434
rect -1100 -514 30 -480
rect 64 -514 80 -480
rect -1100 -560 80 -514
rect -1100 -594 30 -560
rect 64 -594 80 -560
rect -1100 -640 80 -594
rect -1100 -674 30 -640
rect 64 -674 80 -640
rect -1100 -680 80 -674
rect -1500 -700 -1380 -680
rect -1120 -700 80 -680
rect 147 279 201 370
rect 147 245 158 279
rect 192 245 201 279
rect 147 207 201 245
rect 147 173 158 207
rect 192 173 201 207
rect 147 135 201 173
rect 147 101 158 135
rect 192 101 201 135
rect 147 63 201 101
rect 147 29 158 63
rect 192 29 201 63
rect 147 -9 201 29
rect 147 -43 158 -9
rect 192 -43 201 -9
rect 147 -81 201 -43
rect 147 -115 158 -81
rect 192 -115 201 -81
rect 147 -153 201 -115
rect 147 -187 158 -153
rect 192 -187 201 -153
rect 147 -225 201 -187
rect 147 -259 158 -225
rect 192 -259 201 -225
rect 147 -297 201 -259
rect 147 -331 158 -297
rect 192 -331 201 -297
rect 147 -369 201 -331
rect 147 -403 158 -369
rect 192 -403 201 -369
rect 147 -441 201 -403
rect 147 -475 158 -441
rect 192 -475 201 -441
rect 147 -513 201 -475
rect 147 -547 158 -513
rect 192 -547 201 -513
rect 147 -585 201 -547
rect 147 -619 158 -585
rect 192 -619 201 -585
rect 147 -657 201 -619
rect 147 -691 158 -657
rect 192 -691 201 -657
rect 147 -700 201 -691
rect -1500 -800 -700 -700
rect 10 -710 80 -700
rect 149 -703 201 -700
rect 235 279 287 291
rect 235 245 244 279
rect 278 245 287 279
rect 235 221 287 245
rect 235 141 287 169
rect 235 63 287 89
rect 235 61 244 63
rect 278 61 287 63
rect 235 -9 287 9
rect 235 -19 244 -9
rect 278 -19 287 -9
rect 235 -81 287 -71
rect 235 -99 244 -81
rect 278 -99 287 -81
rect 235 -153 287 -151
rect 235 -179 244 -153
rect 278 -179 287 -153
rect 235 -259 244 -231
rect 278 -259 287 -231
rect 235 -331 244 -311
rect 278 -331 287 -311
rect 235 -339 287 -331
rect 235 -403 244 -391
rect 278 -403 287 -391
rect 235 -419 287 -403
rect 235 -475 244 -471
rect 278 -475 287 -471
rect 235 -499 287 -475
rect 235 -579 287 -551
rect 235 -657 287 -631
rect 235 -691 244 -657
rect 278 -691 287 -657
rect 235 -703 287 -691
rect 321 279 373 370
rect 321 245 330 279
rect 364 245 373 279
rect 321 207 373 245
rect 321 173 330 207
rect 364 173 373 207
rect 321 135 373 173
rect 321 101 330 135
rect 364 101 373 135
rect 321 63 373 101
rect 321 29 330 63
rect 364 29 373 63
rect 321 -9 373 29
rect 321 -43 330 -9
rect 364 -43 373 -9
rect 321 -81 373 -43
rect 321 -115 330 -81
rect 364 -115 373 -81
rect 321 -153 373 -115
rect 321 -187 330 -153
rect 364 -187 373 -153
rect 321 -225 373 -187
rect 321 -259 330 -225
rect 364 -259 373 -225
rect 321 -297 373 -259
rect 321 -331 330 -297
rect 364 -331 373 -297
rect 321 -369 373 -331
rect 321 -403 330 -369
rect 364 -403 373 -369
rect 321 -441 373 -403
rect 321 -475 330 -441
rect 364 -475 373 -441
rect 321 -513 373 -475
rect 321 -547 330 -513
rect 364 -547 373 -513
rect 321 -585 373 -547
rect 321 -619 330 -585
rect 364 -619 373 -585
rect 321 -657 373 -619
rect 321 -691 330 -657
rect 364 -691 373 -657
rect 321 -703 373 -691
rect 407 279 459 291
rect 407 245 416 279
rect 450 245 459 279
rect 407 221 459 245
rect 407 141 459 169
rect 407 63 459 89
rect 407 61 416 63
rect 450 61 459 63
rect 407 -9 459 9
rect 407 -19 416 -9
rect 450 -19 459 -9
rect 407 -81 459 -71
rect 407 -99 416 -81
rect 450 -99 459 -81
rect 407 -153 459 -151
rect 407 -179 416 -153
rect 450 -179 459 -153
rect 407 -259 416 -231
rect 450 -259 459 -231
rect 407 -331 416 -311
rect 450 -331 459 -311
rect 407 -339 459 -331
rect 407 -403 416 -391
rect 450 -403 459 -391
rect 407 -419 459 -403
rect 407 -475 416 -471
rect 450 -475 459 -471
rect 407 -499 459 -475
rect 407 -579 459 -551
rect 407 -657 459 -631
rect 407 -691 416 -657
rect 450 -691 459 -657
rect 407 -703 459 -691
rect 493 279 545 370
rect 493 245 502 279
rect 536 245 545 279
rect 493 207 545 245
rect 493 173 502 207
rect 536 173 545 207
rect 493 135 545 173
rect 493 101 502 135
rect 536 101 545 135
rect 493 63 545 101
rect 493 29 502 63
rect 536 29 545 63
rect 493 -9 545 29
rect 493 -43 502 -9
rect 536 -43 545 -9
rect 493 -81 545 -43
rect 493 -115 502 -81
rect 536 -115 545 -81
rect 493 -153 545 -115
rect 493 -187 502 -153
rect 536 -187 545 -153
rect 493 -225 545 -187
rect 493 -259 502 -225
rect 536 -259 545 -225
rect 493 -297 545 -259
rect 493 -331 502 -297
rect 536 -331 545 -297
rect 493 -369 545 -331
rect 493 -403 502 -369
rect 536 -403 545 -369
rect 493 -441 545 -403
rect 493 -475 502 -441
rect 536 -475 545 -441
rect 493 -513 545 -475
rect 493 -547 502 -513
rect 536 -547 545 -513
rect 493 -585 545 -547
rect 493 -619 502 -585
rect 536 -619 545 -585
rect 493 -657 545 -619
rect 493 -691 502 -657
rect 536 -691 545 -657
rect 493 -703 545 -691
rect 579 279 631 291
rect 579 245 588 279
rect 622 245 631 279
rect 579 221 631 245
rect 579 141 631 169
rect 579 63 631 89
rect 579 61 588 63
rect 622 61 631 63
rect 579 -9 631 9
rect 579 -19 588 -9
rect 622 -19 631 -9
rect 579 -81 631 -71
rect 579 -99 588 -81
rect 622 -99 631 -81
rect 579 -153 631 -151
rect 579 -179 588 -153
rect 622 -179 631 -153
rect 579 -259 588 -231
rect 622 -259 631 -231
rect 579 -331 588 -311
rect 622 -331 631 -311
rect 579 -339 631 -331
rect 579 -403 588 -391
rect 622 -403 631 -391
rect 579 -419 631 -403
rect 579 -475 588 -471
rect 622 -475 631 -471
rect 579 -499 631 -475
rect 579 -579 631 -551
rect 579 -657 631 -631
rect 579 -691 588 -657
rect 622 -691 631 -657
rect 579 -703 631 -691
rect 665 279 717 370
rect 665 245 674 279
rect 708 245 717 279
rect 665 207 717 245
rect 665 173 674 207
rect 708 173 717 207
rect 665 135 717 173
rect 665 101 674 135
rect 708 101 717 135
rect 665 63 717 101
rect 665 29 674 63
rect 708 29 717 63
rect 665 -9 717 29
rect 665 -43 674 -9
rect 708 -43 717 -9
rect 665 -81 717 -43
rect 665 -115 674 -81
rect 708 -115 717 -81
rect 665 -153 717 -115
rect 665 -187 674 -153
rect 708 -187 717 -153
rect 665 -225 717 -187
rect 665 -259 674 -225
rect 708 -259 717 -225
rect 665 -297 717 -259
rect 665 -331 674 -297
rect 708 -331 717 -297
rect 665 -369 717 -331
rect 665 -403 674 -369
rect 708 -403 717 -369
rect 665 -441 717 -403
rect 665 -475 674 -441
rect 708 -475 717 -441
rect 665 -513 717 -475
rect 665 -547 674 -513
rect 708 -547 717 -513
rect 665 -585 717 -547
rect 665 -619 674 -585
rect 708 -619 717 -585
rect 665 -657 717 -619
rect 665 -691 674 -657
rect 708 -691 717 -657
rect 665 -703 717 -691
rect 751 279 803 291
rect 751 245 760 279
rect 794 245 803 279
rect 751 221 803 245
rect 751 141 803 169
rect 751 63 803 89
rect 751 61 760 63
rect 794 61 803 63
rect 751 -9 803 9
rect 751 -19 760 -9
rect 794 -19 803 -9
rect 751 -81 803 -71
rect 751 -99 760 -81
rect 794 -99 803 -81
rect 751 -153 803 -151
rect 751 -179 760 -153
rect 794 -179 803 -153
rect 751 -259 760 -231
rect 794 -259 803 -231
rect 751 -331 760 -311
rect 794 -331 803 -311
rect 751 -339 803 -331
rect 751 -403 760 -391
rect 794 -403 803 -391
rect 751 -419 803 -403
rect 751 -475 760 -471
rect 794 -475 803 -471
rect 751 -499 803 -475
rect 751 -579 803 -551
rect 751 -657 803 -631
rect 751 -691 760 -657
rect 794 -691 803 -657
rect 751 -703 803 -691
rect 837 279 891 370
rect 837 245 846 279
rect 880 245 891 279
rect 837 207 891 245
rect 837 173 846 207
rect 880 173 891 207
rect 837 135 891 173
rect 837 101 846 135
rect 880 101 891 135
rect 837 63 891 101
rect 837 29 846 63
rect 880 29 891 63
rect 837 -9 891 29
rect 837 -43 846 -9
rect 880 -43 891 -9
rect 837 -81 891 -43
rect 837 -115 846 -81
rect 880 -115 891 -81
rect 837 -153 891 -115
rect 837 -187 846 -153
rect 880 -187 891 -153
rect 837 -225 891 -187
rect 837 -259 846 -225
rect 880 -259 891 -225
rect 837 -297 891 -259
rect 837 -331 846 -297
rect 880 -331 891 -297
rect 837 -369 891 -331
rect 837 -403 846 -369
rect 880 -403 891 -369
rect 837 -441 891 -403
rect 837 -475 846 -441
rect 880 -475 891 -441
rect 837 -513 891 -475
rect 837 -547 846 -513
rect 880 -547 891 -513
rect 837 -585 891 -547
rect 837 -619 846 -585
rect 880 -619 891 -585
rect 837 -657 891 -619
rect 837 -691 846 -657
rect 880 -691 891 -657
rect 837 -700 891 -691
rect 947 390 1020 450
rect 1100 420 1200 680
rect 1500 420 1600 680
rect 1100 400 1220 420
rect 1480 400 1600 420
rect 947 320 1017 390
rect 947 286 967 320
rect 1001 300 1017 320
rect 1100 300 1600 400
rect 1001 286 1750 300
rect 947 240 1750 286
rect 947 206 967 240
rect 1001 206 1750 240
rect 947 160 1750 206
rect 947 126 967 160
rect 1001 126 1750 160
rect 947 80 1750 126
rect 947 46 967 80
rect 1001 46 1750 80
rect 947 0 1750 46
rect 947 -34 967 0
rect 1001 -34 1750 0
rect 947 -80 1750 -34
rect 947 -114 967 -80
rect 1001 -114 1750 -80
rect 947 -160 1750 -114
rect 947 -194 967 -160
rect 1001 -194 1750 -160
rect 947 -240 1750 -194
rect 947 -274 967 -240
rect 1001 -274 1750 -240
rect 947 -320 1750 -274
rect 947 -354 967 -320
rect 1001 -354 1750 -320
rect 947 -400 1750 -354
rect 947 -434 967 -400
rect 1001 -434 1750 -400
rect 947 -480 1750 -434
rect 947 -514 967 -480
rect 1001 -514 1750 -480
rect 947 -560 1750 -514
rect 947 -594 967 -560
rect 1001 -594 1750 -560
rect 947 -640 1750 -594
rect 947 -674 967 -640
rect 1001 -674 1750 -640
rect 947 -700 1750 -674
rect 837 -703 889 -700
rect 947 -710 1017 -700
rect 174 -749 864 -737
rect 174 -783 258 -749
rect 292 -783 330 -749
rect 364 -783 402 -749
rect 436 -783 602 -749
rect 636 -783 674 -749
rect 708 -783 746 -749
rect 780 -783 864 -749
rect -1500 -900 -1000 -800
rect 174 -840 864 -783
rect 170 -900 867 -840
rect -1500 -920 -1380 -900
rect -1120 -920 -1000 -900
rect -1500 -1180 -1400 -920
rect -1100 -1180 -1000 -920
rect 200 -1100 300 -900
rect 400 -1100 500 -900
rect 600 -1100 700 -900
rect 800 -1100 900 -900
rect -1500 -1200 -1380 -1180
rect -1120 -1200 -1000 -1180
rect -1500 -1400 -1000 -1200
rect -1500 -1420 -1380 -1400
rect -1120 -1420 -1000 -1400
rect -1500 -1680 -1400 -1420
rect -1100 -1680 -1000 -1420
rect -1500 -1700 -1380 -1680
rect -1120 -1700 -1000 -1680
rect -1500 -1900 -1000 -1700
rect -200 -1200 1300 -1100
rect -200 -1700 -100 -1200
rect 1200 -1700 1300 -1200
rect -200 -1800 1300 -1700
rect -1500 -1920 -1380 -1900
rect -1120 -1920 -1000 -1900
rect -4420 -2060 -3600 -2000
rect -5500 -2200 -5380 -2180
rect -5120 -2200 -4880 -2180
rect -4620 -2200 -4540 -2180
rect -5500 -2220 -4540 -2200
rect -3740 -2220 -3600 -2060
rect -5500 -2300 -3600 -2220
rect -1500 -2180 -1400 -1920
rect -1100 -2180 -1000 -1920
rect -1500 -2200 -1380 -2180
rect -1120 -2200 -1000 -2180
rect -1500 -2300 -1000 -2200
rect -11400 -2400 -1000 -2300
rect -14500 -2420 -14380 -2400
rect -14120 -2420 -13880 -2400
rect -13620 -2420 -13380 -2400
rect -13120 -2420 -12880 -2400
rect -12620 -2420 -12380 -2400
rect -12120 -2420 -11880 -2400
rect -11620 -2420 -11380 -2400
rect -11120 -2420 -10880 -2400
rect -10620 -2420 -10380 -2400
rect -10120 -2420 -9880 -2400
rect -9620 -2420 -9380 -2400
rect -9120 -2420 -8880 -2400
rect -8620 -2420 -8380 -2400
rect -8120 -2420 -7880 -2400
rect -7620 -2420 -7380 -2400
rect -7120 -2420 -6880 -2400
rect -6620 -2420 -6380 -2400
rect -6120 -2420 -5880 -2400
rect -5620 -2420 -5380 -2400
rect -5120 -2420 -4880 -2400
rect -4620 -2420 -4380 -2400
rect -4120 -2420 -3880 -2400
rect -3620 -2420 -3380 -2400
rect -3120 -2420 -2880 -2400
rect -2620 -2420 -2380 -2400
rect -2120 -2420 -1880 -2400
rect -1620 -2420 -1380 -2400
rect -1120 -2420 -1000 -2400
rect -14500 -2680 -14400 -2420
rect -14100 -2680 -13900 -2420
rect -13600 -2680 -13400 -2420
rect -13100 -2680 -12900 -2420
rect -12600 -2680 -12400 -2420
rect -12100 -2680 -11900 -2420
rect -11600 -2680 -11400 -2420
rect -11100 -2680 -10900 -2420
rect -10600 -2680 -10400 -2420
rect -10100 -2680 -9900 -2420
rect -9600 -2680 -9400 -2420
rect -9100 -2680 -8900 -2420
rect -8600 -2680 -8400 -2420
rect -8100 -2680 -7900 -2420
rect -7600 -2680 -7400 -2420
rect -7100 -2680 -6900 -2420
rect -6600 -2680 -6400 -2420
rect -6100 -2680 -5900 -2420
rect -5600 -2680 -5400 -2420
rect -5100 -2680 -4900 -2420
rect -4600 -2680 -4400 -2420
rect -4100 -2680 -3900 -2420
rect -3600 -2680 -3400 -2420
rect -3100 -2680 -2900 -2420
rect -2600 -2680 -2400 -2420
rect -2100 -2680 -1900 -2420
rect -1600 -2680 -1400 -2420
rect -1100 -2680 -1000 -2420
rect -14500 -2700 -14380 -2680
rect -14120 -2700 -13880 -2680
rect -13620 -2700 -13380 -2680
rect -13120 -2700 -12880 -2680
rect -12620 -2700 -12380 -2680
rect -12120 -2700 -11880 -2680
rect -11620 -2700 -11380 -2680
rect -11120 -2700 -10880 -2680
rect -10620 -2700 -10380 -2680
rect -10120 -2700 -9880 -2680
rect -9620 -2700 -9380 -2680
rect -9120 -2700 -8880 -2680
rect -8620 -2700 -8380 -2680
rect -8120 -2700 -7880 -2680
rect -7620 -2700 -7380 -2680
rect -7120 -2700 -6880 -2680
rect -6620 -2700 -6380 -2680
rect -6120 -2700 -5880 -2680
rect -5620 -2700 -5380 -2680
rect -5120 -2700 -4880 -2680
rect -4620 -2700 -4380 -2680
rect -4120 -2700 -3880 -2680
rect -3620 -2700 -3380 -2680
rect -3120 -2700 -2880 -2680
rect -2620 -2700 -2380 -2680
rect -2120 -2700 -1880 -2680
rect -1620 -2700 -1380 -2680
rect -1120 -2700 -1000 -2680
rect -14500 -2900 -11600 -2700
rect -11400 -2900 -1000 -2700
rect -14500 -2920 -14380 -2900
rect -14120 -2920 -13880 -2900
rect -13620 -2920 -13380 -2900
rect -13120 -2920 -12880 -2900
rect -12620 -2920 -12380 -2900
rect -12120 -2920 -11880 -2900
rect -11620 -2920 -11380 -2900
rect -11120 -2920 -10880 -2900
rect -10620 -2920 -10380 -2900
rect -10120 -2920 -9880 -2900
rect -9620 -2920 -9380 -2900
rect -9120 -2920 -8880 -2900
rect -8620 -2920 -8380 -2900
rect -8120 -2920 -7880 -2900
rect -7620 -2920 -7380 -2900
rect -7120 -2920 -6880 -2900
rect -6620 -2920 -6380 -2900
rect -6120 -2920 -5880 -2900
rect -5620 -2920 -5380 -2900
rect -5120 -2920 -4880 -2900
rect -4620 -2920 -4380 -2900
rect -4120 -2920 -3880 -2900
rect -3620 -2920 -3380 -2900
rect -3120 -2920 -2880 -2900
rect -2620 -2920 -2380 -2900
rect -2120 -2920 -1880 -2900
rect -1620 -2920 -1380 -2900
rect -1120 -2920 -1000 -2900
rect -14500 -3180 -14400 -2920
rect -14100 -3180 -13900 -2920
rect -13600 -3180 -13400 -2920
rect -13100 -3180 -12900 -2920
rect -12600 -3180 -12400 -2920
rect -12100 -3180 -11900 -2920
rect -11600 -3180 -11400 -2920
rect -11100 -3180 -10900 -2920
rect -10600 -3180 -10400 -2920
rect -10100 -3180 -9900 -2920
rect -9600 -3180 -9400 -2920
rect -9100 -3180 -8900 -2920
rect -8600 -3180 -8400 -2920
rect -8100 -3180 -7900 -2920
rect -7600 -3180 -7400 -2920
rect -7100 -3180 -6900 -2920
rect -6600 -3180 -6400 -2920
rect -6100 -3180 -5900 -2920
rect -5600 -3180 -5400 -2920
rect -5100 -3180 -4900 -2920
rect -4600 -3180 -4400 -2920
rect -4100 -3180 -3900 -2920
rect -3600 -3180 -3400 -2920
rect -3100 -3180 -2900 -2920
rect -2600 -3180 -2400 -2920
rect -2100 -3180 -1900 -2920
rect -1600 -3180 -1400 -2920
rect -1100 -3180 -1000 -2920
rect -14500 -3200 -14380 -3180
rect -14120 -3200 -13880 -3180
rect -13620 -3200 -13380 -3180
rect -13120 -3200 -12880 -3180
rect -12620 -3200 -12380 -3180
rect -12120 -3200 -11880 -3180
rect -11620 -3200 -11380 -3180
rect -11120 -3200 -10880 -3180
rect -10620 -3200 -10380 -3180
rect -10120 -3200 -9880 -3180
rect -9620 -3200 -9380 -3180
rect -9120 -3200 -8880 -3180
rect -8620 -3200 -8380 -3180
rect -8120 -3200 -7880 -3180
rect -7620 -3200 -7380 -3180
rect -7120 -3200 -6880 -3180
rect -6620 -3200 -6380 -3180
rect -6120 -3200 -5880 -3180
rect -5620 -3200 -5380 -3180
rect -5120 -3200 -4880 -3180
rect -4620 -3200 -4380 -3180
rect -4120 -3200 -3880 -3180
rect -3620 -3200 -3380 -3180
rect -3120 -3200 -2880 -3180
rect -2620 -3200 -2380 -3180
rect -2120 -3200 -1880 -3180
rect -1620 -3200 -1380 -3180
rect -1120 -3200 -1000 -3180
rect -14500 -3300 -1000 -3200
<< via1 >>
rect -6700 17174 -6520 17240
rect -6700 17160 -6697 17174
rect -6697 17160 -6663 17174
rect -6663 17160 -6625 17174
rect -6625 17160 -6591 17174
rect -6591 17160 -6553 17174
rect -6553 17160 -6520 17174
rect -6720 16506 -6668 16542
rect -6720 16490 -6711 16506
rect -6711 16490 -6677 16506
rect -6677 16490 -6668 16506
rect -6720 16472 -6711 16478
rect -6711 16472 -6677 16478
rect -6677 16472 -6668 16478
rect -6720 16434 -6668 16472
rect -6720 16426 -6711 16434
rect -6711 16426 -6677 16434
rect -6677 16426 -6668 16434
rect -6720 16400 -6711 16414
rect -6711 16400 -6677 16414
rect -6677 16400 -6668 16414
rect -6720 16362 -6668 16400
rect -6720 16328 -6711 16350
rect -6711 16328 -6677 16350
rect -6677 16328 -6668 16350
rect -6720 16298 -6668 16328
rect -6720 16256 -6711 16286
rect -6711 16256 -6677 16286
rect -6677 16256 -6668 16286
rect -6720 16234 -6668 16256
rect -6720 16218 -6668 16222
rect -6720 16184 -6711 16218
rect -6711 16184 -6677 16218
rect -6677 16184 -6668 16218
rect -6720 16170 -6668 16184
rect -6720 16146 -6668 16158
rect -6720 16112 -6711 16146
rect -6711 16112 -6677 16146
rect -6677 16112 -6668 16146
rect -6720 16106 -6668 16112
rect -6634 17082 -6582 17088
rect -6634 17048 -6625 17082
rect -6625 17048 -6591 17082
rect -6591 17048 -6582 17082
rect -6634 17036 -6582 17048
rect -6634 17010 -6582 17024
rect -6634 16976 -6625 17010
rect -6625 16976 -6591 17010
rect -6591 16976 -6582 17010
rect -6634 16972 -6582 16976
rect -6634 16938 -6582 16960
rect -6634 16908 -6625 16938
rect -6625 16908 -6591 16938
rect -6591 16908 -6582 16938
rect -6634 16866 -6582 16896
rect -6634 16844 -6625 16866
rect -6625 16844 -6591 16866
rect -6591 16844 -6582 16866
rect -6634 16794 -6582 16832
rect -6634 16780 -6625 16794
rect -6625 16780 -6591 16794
rect -6591 16780 -6582 16794
rect -6634 16760 -6625 16768
rect -6625 16760 -6591 16768
rect -6591 16760 -6582 16768
rect -6634 16722 -6582 16760
rect -6634 16716 -6625 16722
rect -6625 16716 -6591 16722
rect -6591 16716 -6582 16722
rect -6634 16688 -6625 16704
rect -6625 16688 -6591 16704
rect -6591 16688 -6582 16704
rect -6634 16652 -6582 16688
rect -6548 16506 -6496 16542
rect -6548 16490 -6539 16506
rect -6539 16490 -6505 16506
rect -6505 16490 -6496 16506
rect -6548 16472 -6539 16478
rect -6539 16472 -6505 16478
rect -6505 16472 -6496 16478
rect -6548 16434 -6496 16472
rect -6548 16426 -6539 16434
rect -6539 16426 -6505 16434
rect -6505 16426 -6496 16434
rect -6548 16400 -6539 16414
rect -6539 16400 -6505 16414
rect -6505 16400 -6496 16414
rect -6548 16362 -6496 16400
rect -6548 16328 -6539 16350
rect -6539 16328 -6505 16350
rect -6505 16328 -6496 16350
rect -6548 16298 -6496 16328
rect -6548 16256 -6539 16286
rect -6539 16256 -6505 16286
rect -6505 16256 -6496 16286
rect -6548 16234 -6496 16256
rect -6548 16218 -6496 16222
rect -6548 16184 -6539 16218
rect -6539 16184 -6505 16218
rect -6505 16184 -6496 16218
rect -6548 16170 -6496 16184
rect -6548 16146 -6496 16158
rect -6548 16112 -6539 16146
rect -6539 16112 -6505 16146
rect -6505 16112 -6496 16146
rect -6548 16106 -6496 16112
rect -6300 17174 -6120 17240
rect -6300 17160 -6269 17174
rect -6269 17160 -6231 17174
rect -6231 17160 -6197 17174
rect -6197 17160 -6159 17174
rect -6159 17160 -6125 17174
rect -6125 17160 -6120 17174
rect -5900 17174 -5720 17240
rect -5900 17160 -5875 17174
rect -5875 17160 -5837 17174
rect -5837 17160 -5803 17174
rect -5803 17160 -5765 17174
rect -5765 17160 -5731 17174
rect -5731 17160 -5720 17174
rect -5520 17174 -5340 17240
rect -5520 17160 -5515 17174
rect -5515 17160 -5481 17174
rect -5481 17160 -5443 17174
rect -5443 17160 -5409 17174
rect -5409 17160 -5371 17174
rect -5371 17160 -5340 17174
rect -6326 16506 -6274 16542
rect -6326 16490 -6317 16506
rect -6317 16490 -6283 16506
rect -6283 16490 -6274 16506
rect -6326 16472 -6317 16478
rect -6317 16472 -6283 16478
rect -6283 16472 -6274 16478
rect -6326 16434 -6274 16472
rect -6326 16426 -6317 16434
rect -6317 16426 -6283 16434
rect -6283 16426 -6274 16434
rect -6326 16400 -6317 16414
rect -6317 16400 -6283 16414
rect -6283 16400 -6274 16414
rect -6326 16362 -6274 16400
rect -6326 16328 -6317 16350
rect -6317 16328 -6283 16350
rect -6283 16328 -6274 16350
rect -6326 16298 -6274 16328
rect -6326 16256 -6317 16286
rect -6317 16256 -6283 16286
rect -6283 16256 -6274 16286
rect -6326 16234 -6274 16256
rect -6326 16218 -6274 16222
rect -6326 16184 -6317 16218
rect -6317 16184 -6283 16218
rect -6283 16184 -6274 16218
rect -6326 16170 -6274 16184
rect -6326 16146 -6274 16158
rect -6326 16112 -6317 16146
rect -6317 16112 -6283 16146
rect -6283 16112 -6274 16146
rect -6326 16106 -6274 16112
rect -6240 17082 -6188 17088
rect -6240 17048 -6231 17082
rect -6231 17048 -6197 17082
rect -6197 17048 -6188 17082
rect -6240 17036 -6188 17048
rect -6240 17010 -6188 17024
rect -6240 16976 -6231 17010
rect -6231 16976 -6197 17010
rect -6197 16976 -6188 17010
rect -6240 16972 -6188 16976
rect -6240 16938 -6188 16960
rect -6240 16908 -6231 16938
rect -6231 16908 -6197 16938
rect -6197 16908 -6188 16938
rect -6240 16866 -6188 16896
rect -6240 16844 -6231 16866
rect -6231 16844 -6197 16866
rect -6197 16844 -6188 16866
rect -6240 16794 -6188 16832
rect -6240 16780 -6231 16794
rect -6231 16780 -6197 16794
rect -6197 16780 -6188 16794
rect -6240 16760 -6231 16768
rect -6231 16760 -6197 16768
rect -6197 16760 -6188 16768
rect -6240 16722 -6188 16760
rect -6240 16716 -6231 16722
rect -6231 16716 -6197 16722
rect -6197 16716 -6188 16722
rect -6240 16688 -6231 16704
rect -6231 16688 -6197 16704
rect -6197 16688 -6188 16704
rect -6240 16652 -6188 16688
rect -6154 16506 -6102 16542
rect -6154 16490 -6145 16506
rect -6145 16490 -6111 16506
rect -6111 16490 -6102 16506
rect -6154 16472 -6145 16478
rect -6145 16472 -6111 16478
rect -6111 16472 -6102 16478
rect -6154 16434 -6102 16472
rect -6154 16426 -6145 16434
rect -6145 16426 -6111 16434
rect -6111 16426 -6102 16434
rect -6154 16400 -6145 16414
rect -6145 16400 -6111 16414
rect -6111 16400 -6102 16414
rect -6154 16362 -6102 16400
rect -6154 16328 -6145 16350
rect -6145 16328 -6111 16350
rect -6111 16328 -6102 16350
rect -6154 16298 -6102 16328
rect -6154 16256 -6145 16286
rect -6145 16256 -6111 16286
rect -6111 16256 -6102 16286
rect -6154 16234 -6102 16256
rect -6154 16218 -6102 16222
rect -6154 16184 -6145 16218
rect -6145 16184 -6111 16218
rect -6111 16184 -6102 16218
rect -6154 16170 -6102 16184
rect -6154 16146 -6102 16158
rect -6154 16112 -6145 16146
rect -6145 16112 -6111 16146
rect -6111 16112 -6102 16146
rect -6154 16106 -6102 16112
rect -5932 16506 -5880 16542
rect -5932 16490 -5923 16506
rect -5923 16490 -5889 16506
rect -5889 16490 -5880 16506
rect -5932 16472 -5923 16478
rect -5923 16472 -5889 16478
rect -5889 16472 -5880 16478
rect -5932 16434 -5880 16472
rect -5932 16426 -5923 16434
rect -5923 16426 -5889 16434
rect -5889 16426 -5880 16434
rect -5932 16400 -5923 16414
rect -5923 16400 -5889 16414
rect -5889 16400 -5880 16414
rect -5932 16362 -5880 16400
rect -5932 16328 -5923 16350
rect -5923 16328 -5889 16350
rect -5889 16328 -5880 16350
rect -5932 16298 -5880 16328
rect -5932 16256 -5923 16286
rect -5923 16256 -5889 16286
rect -5889 16256 -5880 16286
rect -5932 16234 -5880 16256
rect -5932 16218 -5880 16222
rect -5932 16184 -5923 16218
rect -5923 16184 -5889 16218
rect -5889 16184 -5880 16218
rect -5932 16170 -5880 16184
rect -5932 16146 -5880 16158
rect -5932 16112 -5923 16146
rect -5923 16112 -5889 16146
rect -5889 16112 -5880 16146
rect -5932 16106 -5880 16112
rect -5846 17082 -5794 17088
rect -5846 17048 -5837 17082
rect -5837 17048 -5803 17082
rect -5803 17048 -5794 17082
rect -5846 17036 -5794 17048
rect -5846 17010 -5794 17024
rect -5846 16976 -5837 17010
rect -5837 16976 -5803 17010
rect -5803 16976 -5794 17010
rect -5846 16972 -5794 16976
rect -5846 16938 -5794 16960
rect -5846 16908 -5837 16938
rect -5837 16908 -5803 16938
rect -5803 16908 -5794 16938
rect -5846 16866 -5794 16896
rect -5846 16844 -5837 16866
rect -5837 16844 -5803 16866
rect -5803 16844 -5794 16866
rect -5846 16794 -5794 16832
rect -5846 16780 -5837 16794
rect -5837 16780 -5803 16794
rect -5803 16780 -5794 16794
rect -5846 16760 -5837 16768
rect -5837 16760 -5803 16768
rect -5803 16760 -5794 16768
rect -5846 16722 -5794 16760
rect -5846 16716 -5837 16722
rect -5837 16716 -5803 16722
rect -5803 16716 -5794 16722
rect -5846 16688 -5837 16704
rect -5837 16688 -5803 16704
rect -5803 16688 -5794 16704
rect -5846 16652 -5794 16688
rect -5760 16506 -5708 16542
rect -5760 16490 -5751 16506
rect -5751 16490 -5717 16506
rect -5717 16490 -5708 16506
rect -5760 16472 -5751 16478
rect -5751 16472 -5717 16478
rect -5717 16472 -5708 16478
rect -5760 16434 -5708 16472
rect -5760 16426 -5751 16434
rect -5751 16426 -5717 16434
rect -5717 16426 -5708 16434
rect -5760 16400 -5751 16414
rect -5751 16400 -5717 16414
rect -5717 16400 -5708 16414
rect -5760 16362 -5708 16400
rect -5760 16328 -5751 16350
rect -5751 16328 -5717 16350
rect -5717 16328 -5708 16350
rect -5760 16298 -5708 16328
rect -5760 16256 -5751 16286
rect -5751 16256 -5717 16286
rect -5717 16256 -5708 16286
rect -5760 16234 -5708 16256
rect -5760 16218 -5708 16222
rect -5760 16184 -5751 16218
rect -5751 16184 -5717 16218
rect -5717 16184 -5708 16218
rect -5760 16170 -5708 16184
rect -5760 16146 -5708 16158
rect -5760 16112 -5751 16146
rect -5751 16112 -5717 16146
rect -5717 16112 -5708 16146
rect -5760 16106 -5708 16112
rect -5538 16506 -5486 16542
rect -5538 16490 -5529 16506
rect -5529 16490 -5495 16506
rect -5495 16490 -5486 16506
rect -5538 16472 -5529 16478
rect -5529 16472 -5495 16478
rect -5495 16472 -5486 16478
rect -5538 16434 -5486 16472
rect -5538 16426 -5529 16434
rect -5529 16426 -5495 16434
rect -5495 16426 -5486 16434
rect -5538 16400 -5529 16414
rect -5529 16400 -5495 16414
rect -5495 16400 -5486 16414
rect -5538 16362 -5486 16400
rect -5538 16328 -5529 16350
rect -5529 16328 -5495 16350
rect -5495 16328 -5486 16350
rect -5538 16298 -5486 16328
rect -5538 16256 -5529 16286
rect -5529 16256 -5495 16286
rect -5495 16256 -5486 16286
rect -5538 16234 -5486 16256
rect -5538 16218 -5486 16222
rect -5538 16184 -5529 16218
rect -5529 16184 -5495 16218
rect -5495 16184 -5486 16218
rect -5538 16170 -5486 16184
rect -5538 16146 -5486 16158
rect -5538 16112 -5529 16146
rect -5529 16112 -5495 16146
rect -5495 16112 -5486 16146
rect -5538 16106 -5486 16112
rect -5452 17082 -5400 17088
rect -5452 17048 -5443 17082
rect -5443 17048 -5409 17082
rect -5409 17048 -5400 17082
rect -5452 17036 -5400 17048
rect -5452 17010 -5400 17024
rect -5452 16976 -5443 17010
rect -5443 16976 -5409 17010
rect -5409 16976 -5400 17010
rect -5452 16972 -5400 16976
rect -5452 16938 -5400 16960
rect -5452 16908 -5443 16938
rect -5443 16908 -5409 16938
rect -5409 16908 -5400 16938
rect -5452 16866 -5400 16896
rect -5452 16844 -5443 16866
rect -5443 16844 -5409 16866
rect -5409 16844 -5400 16866
rect -5452 16794 -5400 16832
rect -5452 16780 -5443 16794
rect -5443 16780 -5409 16794
rect -5409 16780 -5400 16794
rect -5452 16760 -5443 16768
rect -5443 16760 -5409 16768
rect -5409 16760 -5400 16768
rect -5452 16722 -5400 16760
rect -5452 16716 -5443 16722
rect -5443 16716 -5409 16722
rect -5409 16716 -5400 16722
rect -5452 16688 -5443 16704
rect -5443 16688 -5409 16704
rect -5409 16688 -5400 16704
rect -5452 16652 -5400 16688
rect -5366 16506 -5314 16542
rect -5366 16490 -5357 16506
rect -5357 16490 -5323 16506
rect -5323 16490 -5314 16506
rect -5366 16472 -5357 16478
rect -5357 16472 -5323 16478
rect -5323 16472 -5314 16478
rect -5366 16434 -5314 16472
rect -5366 16426 -5357 16434
rect -5357 16426 -5323 16434
rect -5323 16426 -5314 16434
rect -5366 16400 -5357 16414
rect -5357 16400 -5323 16414
rect -5323 16400 -5314 16414
rect -5366 16362 -5314 16400
rect -5366 16328 -5357 16350
rect -5357 16328 -5323 16350
rect -5323 16328 -5314 16350
rect -5366 16298 -5314 16328
rect -5366 16256 -5357 16286
rect -5357 16256 -5323 16286
rect -5323 16256 -5314 16286
rect -5366 16234 -5314 16256
rect -5366 16218 -5314 16222
rect -5366 16184 -5357 16218
rect -5357 16184 -5323 16218
rect -5323 16184 -5314 16218
rect -5366 16170 -5314 16184
rect -5366 16146 -5314 16158
rect -5366 16112 -5357 16146
rect -5357 16112 -5323 16146
rect -5323 16112 -5314 16146
rect -5366 16106 -5314 16112
rect -6740 15820 -6460 15900
rect -6000 15820 -5280 15900
rect -4700 7800 -4500 8600
rect -1980 7660 -1820 7680
rect -1980 7540 -1960 7660
rect -1960 7540 -1840 7660
rect -1840 7540 -1820 7660
rect -1980 7520 -1820 7540
rect 31 8399 83 8411
rect 31 8365 40 8399
rect 40 8365 74 8399
rect 74 8365 83 8399
rect 31 8359 83 8365
rect 31 8327 83 8331
rect 31 8293 40 8327
rect 40 8293 74 8327
rect 74 8293 83 8327
rect 31 8279 83 8293
rect 31 8221 40 8251
rect 40 8221 74 8251
rect 74 8221 83 8251
rect 31 8199 83 8221
rect 31 8149 40 8171
rect 40 8149 74 8171
rect 74 8149 83 8171
rect 31 8119 83 8149
rect 31 8077 40 8091
rect 40 8077 74 8091
rect 74 8077 83 8091
rect 31 8039 83 8077
rect 31 8005 40 8011
rect 40 8005 74 8011
rect 74 8005 83 8011
rect 31 7967 83 8005
rect 31 7959 40 7967
rect 40 7959 74 7967
rect 74 7959 83 7967
rect 31 7895 83 7931
rect 31 7879 40 7895
rect 40 7879 74 7895
rect 74 7879 83 7895
rect 31 7823 83 7851
rect 31 7799 40 7823
rect 40 7799 74 7823
rect 74 7799 83 7823
rect 31 7751 83 7771
rect 31 7719 40 7751
rect 40 7719 74 7751
rect 74 7719 83 7751
rect 31 7679 83 7691
rect 31 7645 40 7679
rect 40 7645 74 7679
rect 74 7645 83 7679
rect 31 7639 83 7645
rect 31 7607 83 7611
rect 31 7573 40 7607
rect 40 7573 74 7607
rect 74 7573 83 7607
rect 31 7559 83 7573
rect 203 8399 255 8411
rect 203 8365 212 8399
rect 212 8365 246 8399
rect 246 8365 255 8399
rect 203 8359 255 8365
rect 203 8327 255 8331
rect 203 8293 212 8327
rect 212 8293 246 8327
rect 246 8293 255 8327
rect 203 8279 255 8293
rect 203 8221 212 8251
rect 212 8221 246 8251
rect 246 8221 255 8251
rect 203 8199 255 8221
rect 203 8149 212 8171
rect 212 8149 246 8171
rect 246 8149 255 8171
rect 203 8119 255 8149
rect 203 8077 212 8091
rect 212 8077 246 8091
rect 246 8077 255 8091
rect 203 8039 255 8077
rect 203 8005 212 8011
rect 212 8005 246 8011
rect 246 8005 255 8011
rect 203 7967 255 8005
rect 203 7959 212 7967
rect 212 7959 246 7967
rect 246 7959 255 7967
rect 203 7895 255 7931
rect 203 7879 212 7895
rect 212 7879 246 7895
rect 246 7879 255 7895
rect 203 7823 255 7851
rect 203 7799 212 7823
rect 212 7799 246 7823
rect 246 7799 255 7823
rect 203 7751 255 7771
rect 203 7719 212 7751
rect 212 7719 246 7751
rect 246 7719 255 7751
rect 203 7679 255 7691
rect 203 7645 212 7679
rect 212 7645 246 7679
rect 246 7645 255 7679
rect 203 7639 255 7645
rect 203 7607 255 7611
rect 203 7573 212 7607
rect 212 7573 246 7607
rect 246 7573 255 7607
rect 203 7559 255 7573
rect 375 8399 427 8411
rect 375 8365 384 8399
rect 384 8365 418 8399
rect 418 8365 427 8399
rect 375 8359 427 8365
rect 375 8327 427 8331
rect 375 8293 384 8327
rect 384 8293 418 8327
rect 418 8293 427 8327
rect 375 8279 427 8293
rect 375 8221 384 8251
rect 384 8221 418 8251
rect 418 8221 427 8251
rect 375 8199 427 8221
rect 375 8149 384 8171
rect 384 8149 418 8171
rect 418 8149 427 8171
rect 375 8119 427 8149
rect 375 8077 384 8091
rect 384 8077 418 8091
rect 418 8077 427 8091
rect 375 8039 427 8077
rect 375 8005 384 8011
rect 384 8005 418 8011
rect 418 8005 427 8011
rect 375 7967 427 8005
rect 375 7959 384 7967
rect 384 7959 418 7967
rect 418 7959 427 7967
rect 375 7895 427 7931
rect 375 7879 384 7895
rect 384 7879 418 7895
rect 418 7879 427 7895
rect 375 7823 427 7851
rect 375 7799 384 7823
rect 384 7799 418 7823
rect 418 7799 427 7823
rect 375 7751 427 7771
rect 375 7719 384 7751
rect 384 7719 418 7751
rect 418 7719 427 7751
rect 375 7679 427 7691
rect 375 7645 384 7679
rect 384 7645 418 7679
rect 418 7645 427 7679
rect 375 7639 427 7645
rect 375 7607 427 7611
rect 375 7573 384 7607
rect 384 7573 418 7607
rect 418 7573 427 7607
rect 375 7559 427 7573
rect 547 8399 599 8411
rect 547 8365 556 8399
rect 556 8365 590 8399
rect 590 8365 599 8399
rect 547 8359 599 8365
rect 547 8327 599 8331
rect 547 8293 556 8327
rect 556 8293 590 8327
rect 590 8293 599 8327
rect 547 8279 599 8293
rect 547 8221 556 8251
rect 556 8221 590 8251
rect 590 8221 599 8251
rect 547 8199 599 8221
rect 547 8149 556 8171
rect 556 8149 590 8171
rect 590 8149 599 8171
rect 547 8119 599 8149
rect 547 8077 556 8091
rect 556 8077 590 8091
rect 590 8077 599 8091
rect 547 8039 599 8077
rect 547 8005 556 8011
rect 556 8005 590 8011
rect 590 8005 599 8011
rect 547 7967 599 8005
rect 547 7959 556 7967
rect 556 7959 590 7967
rect 590 7959 599 7967
rect 547 7895 599 7931
rect 547 7879 556 7895
rect 556 7879 590 7895
rect 590 7879 599 7895
rect 547 7823 599 7851
rect 547 7799 556 7823
rect 556 7799 590 7823
rect 590 7799 599 7823
rect 547 7751 599 7771
rect 547 7719 556 7751
rect 556 7719 590 7751
rect 590 7719 599 7751
rect 547 7679 599 7691
rect 547 7645 556 7679
rect 556 7645 590 7679
rect 590 7645 599 7679
rect 547 7639 599 7645
rect 547 7607 599 7611
rect 547 7573 556 7607
rect 556 7573 590 7607
rect 590 7573 599 7607
rect 547 7559 599 7573
rect 719 8399 771 8411
rect 719 8365 728 8399
rect 728 8365 762 8399
rect 762 8365 771 8399
rect 719 8359 771 8365
rect 719 8327 771 8331
rect 719 8293 728 8327
rect 728 8293 762 8327
rect 762 8293 771 8327
rect 719 8279 771 8293
rect 719 8221 728 8251
rect 728 8221 762 8251
rect 762 8221 771 8251
rect 719 8199 771 8221
rect 719 8149 728 8171
rect 728 8149 762 8171
rect 762 8149 771 8171
rect 719 8119 771 8149
rect 719 8077 728 8091
rect 728 8077 762 8091
rect 762 8077 771 8091
rect 719 8039 771 8077
rect 719 8005 728 8011
rect 728 8005 762 8011
rect 762 8005 771 8011
rect 719 7967 771 8005
rect 719 7959 728 7967
rect 728 7959 762 7967
rect 762 7959 771 7967
rect 719 7895 771 7931
rect 719 7879 728 7895
rect 728 7879 762 7895
rect 762 7879 771 7895
rect 719 7823 771 7851
rect 719 7799 728 7823
rect 728 7799 762 7823
rect 762 7799 771 7823
rect 719 7751 771 7771
rect 719 7719 728 7751
rect 728 7719 762 7751
rect 762 7719 771 7751
rect 719 7679 771 7691
rect 719 7645 728 7679
rect 728 7645 762 7679
rect 762 7645 771 7679
rect 719 7639 771 7645
rect 719 7607 771 7611
rect 719 7573 728 7607
rect 728 7573 762 7607
rect 762 7573 771 7607
rect 719 7559 771 7573
rect 891 8399 943 8411
rect 891 8365 900 8399
rect 900 8365 934 8399
rect 934 8365 943 8399
rect 891 8359 943 8365
rect 891 8327 943 8331
rect 891 8293 900 8327
rect 900 8293 934 8327
rect 934 8293 943 8327
rect 891 8279 943 8293
rect 891 8221 900 8251
rect 900 8221 934 8251
rect 934 8221 943 8251
rect 891 8199 943 8221
rect 891 8149 900 8171
rect 900 8149 934 8171
rect 934 8149 943 8171
rect 891 8119 943 8149
rect 891 8077 900 8091
rect 900 8077 934 8091
rect 934 8077 943 8091
rect 891 8039 943 8077
rect 891 8005 900 8011
rect 900 8005 934 8011
rect 934 8005 943 8011
rect 891 7967 943 8005
rect 891 7959 900 7967
rect 900 7959 934 7967
rect 934 7959 943 7967
rect 891 7895 943 7931
rect 891 7879 900 7895
rect 900 7879 934 7895
rect 934 7879 943 7895
rect 891 7823 943 7851
rect 891 7799 900 7823
rect 900 7799 934 7823
rect 934 7799 943 7823
rect 891 7751 943 7771
rect 891 7719 900 7751
rect 900 7719 934 7751
rect 934 7719 943 7751
rect 891 7679 943 7691
rect 891 7645 900 7679
rect 900 7645 934 7679
rect 934 7645 943 7679
rect 891 7639 943 7645
rect 891 7607 943 7611
rect 891 7573 900 7607
rect 900 7573 934 7607
rect 934 7573 943 7607
rect 891 7559 943 7573
rect -14 7300 996 7400
rect -2350 7110 -2150 7180
rect -1850 7110 -1650 7180
rect -2480 6850 -2410 7050
rect -2090 6850 -2020 7050
rect -1980 6850 -1910 7050
rect -1590 6850 -1520 7050
rect -2350 6720 -2150 6790
rect -1850 6720 -1650 6790
rect -2350 6610 -2150 6680
rect -1850 6610 -1650 6680
rect -2480 6350 -2410 6550
rect -2090 6350 -2020 6550
rect -1980 6350 -1910 6550
rect -1590 6350 -1520 6550
rect -2350 6220 -2150 6290
rect -1850 6220 -1650 6290
rect -3850 6110 -3650 6180
rect -3350 6110 -3150 6180
rect -2850 6110 -2650 6180
rect -2350 6110 -2150 6180
rect -1850 6110 -1650 6180
rect -3980 5850 -3910 6050
rect -3590 5850 -3520 6050
rect -3480 5850 -3410 6050
rect -3090 5850 -3020 6050
rect -2980 5850 -2910 6050
rect -2590 5850 -2520 6050
rect -2480 5850 -2410 6050
rect -2090 5850 -2020 6050
rect -1980 5850 -1910 6050
rect -1590 5850 -1520 6050
rect -3850 5720 -3650 5790
rect -3350 5720 -3150 5790
rect -2850 5720 -2650 5790
rect -2350 5720 -2150 5790
rect -1850 5720 -1650 5790
rect -980 7000 -820 7020
rect -980 6880 -960 7000
rect -960 6880 -840 7000
rect -840 6880 -820 7000
rect -980 6860 -820 6880
rect -1180 5900 -1020 5920
rect -1180 5780 -1160 5900
rect -1160 5780 -1040 5900
rect -1040 5780 -1020 5900
rect -1180 5760 -1020 5780
rect -3850 5610 -3650 5680
rect -3350 5610 -3150 5680
rect -2850 5610 -2650 5680
rect -2350 5610 -2150 5680
rect -3980 5350 -3910 5550
rect -3590 5350 -3520 5550
rect -3480 5350 -3410 5550
rect -3090 5350 -3020 5550
rect -2980 5350 -2910 5550
rect -2590 5350 -2520 5550
rect -2480 5350 -2410 5550
rect -2090 5350 -2020 5550
rect -3850 5220 -3650 5290
rect -3350 5220 -3150 5290
rect -2850 5220 -2650 5290
rect -2350 5220 -2150 5290
rect 170 380 870 460
rect -11600 -1900 -11400 -1700
rect -11600 -2400 -11400 -2200
rect -4300 -720 -4140 -690
rect -4300 -860 -4260 -720
rect -4260 -860 -4140 -720
rect -4300 -890 -4140 -860
rect -3960 -720 -3800 -690
rect -3960 -860 -3940 -720
rect -3940 -860 -3820 -720
rect -3820 -860 -3800 -720
rect -3960 -890 -3800 -860
rect 235 207 287 221
rect 235 173 244 207
rect 244 173 278 207
rect 278 173 287 207
rect 235 169 287 173
rect 235 135 287 141
rect 235 101 244 135
rect 244 101 278 135
rect 278 101 287 135
rect 235 89 287 101
rect 235 29 244 61
rect 244 29 278 61
rect 278 29 287 61
rect 235 9 287 29
rect 235 -43 244 -19
rect 244 -43 278 -19
rect 278 -43 287 -19
rect 235 -71 287 -43
rect 235 -115 244 -99
rect 244 -115 278 -99
rect 278 -115 287 -99
rect 235 -151 287 -115
rect 235 -187 244 -179
rect 244 -187 278 -179
rect 278 -187 287 -179
rect 235 -225 287 -187
rect 235 -231 244 -225
rect 244 -231 278 -225
rect 278 -231 287 -225
rect 235 -297 287 -259
rect 235 -311 244 -297
rect 244 -311 278 -297
rect 278 -311 287 -297
rect 235 -369 287 -339
rect 235 -391 244 -369
rect 244 -391 278 -369
rect 278 -391 287 -369
rect 235 -441 287 -419
rect 235 -471 244 -441
rect 244 -471 278 -441
rect 278 -471 287 -441
rect 235 -513 287 -499
rect 235 -547 244 -513
rect 244 -547 278 -513
rect 278 -547 287 -513
rect 235 -551 287 -547
rect 235 -585 287 -579
rect 235 -619 244 -585
rect 244 -619 278 -585
rect 278 -619 287 -585
rect 235 -631 287 -619
rect 407 207 459 221
rect 407 173 416 207
rect 416 173 450 207
rect 450 173 459 207
rect 407 169 459 173
rect 407 135 459 141
rect 407 101 416 135
rect 416 101 450 135
rect 450 101 459 135
rect 407 89 459 101
rect 407 29 416 61
rect 416 29 450 61
rect 450 29 459 61
rect 407 9 459 29
rect 407 -43 416 -19
rect 416 -43 450 -19
rect 450 -43 459 -19
rect 407 -71 459 -43
rect 407 -115 416 -99
rect 416 -115 450 -99
rect 450 -115 459 -99
rect 407 -151 459 -115
rect 407 -187 416 -179
rect 416 -187 450 -179
rect 450 -187 459 -179
rect 407 -225 459 -187
rect 407 -231 416 -225
rect 416 -231 450 -225
rect 450 -231 459 -225
rect 407 -297 459 -259
rect 407 -311 416 -297
rect 416 -311 450 -297
rect 450 -311 459 -297
rect 407 -369 459 -339
rect 407 -391 416 -369
rect 416 -391 450 -369
rect 450 -391 459 -369
rect 407 -441 459 -419
rect 407 -471 416 -441
rect 416 -471 450 -441
rect 450 -471 459 -441
rect 407 -513 459 -499
rect 407 -547 416 -513
rect 416 -547 450 -513
rect 450 -547 459 -513
rect 407 -551 459 -547
rect 407 -585 459 -579
rect 407 -619 416 -585
rect 416 -619 450 -585
rect 450 -619 459 -585
rect 407 -631 459 -619
rect 579 207 631 221
rect 579 173 588 207
rect 588 173 622 207
rect 622 173 631 207
rect 579 169 631 173
rect 579 135 631 141
rect 579 101 588 135
rect 588 101 622 135
rect 622 101 631 135
rect 579 89 631 101
rect 579 29 588 61
rect 588 29 622 61
rect 622 29 631 61
rect 579 9 631 29
rect 579 -43 588 -19
rect 588 -43 622 -19
rect 622 -43 631 -19
rect 579 -71 631 -43
rect 579 -115 588 -99
rect 588 -115 622 -99
rect 622 -115 631 -99
rect 579 -151 631 -115
rect 579 -187 588 -179
rect 588 -187 622 -179
rect 622 -187 631 -179
rect 579 -225 631 -187
rect 579 -231 588 -225
rect 588 -231 622 -225
rect 622 -231 631 -225
rect 579 -297 631 -259
rect 579 -311 588 -297
rect 588 -311 622 -297
rect 622 -311 631 -297
rect 579 -369 631 -339
rect 579 -391 588 -369
rect 588 -391 622 -369
rect 622 -391 631 -369
rect 579 -441 631 -419
rect 579 -471 588 -441
rect 588 -471 622 -441
rect 622 -471 631 -441
rect 579 -513 631 -499
rect 579 -547 588 -513
rect 588 -547 622 -513
rect 622 -547 631 -513
rect 579 -551 631 -547
rect 579 -585 631 -579
rect 579 -619 588 -585
rect 588 -619 622 -585
rect 622 -619 631 -585
rect 579 -631 631 -619
rect 751 207 803 221
rect 751 173 760 207
rect 760 173 794 207
rect 794 173 803 207
rect 751 169 803 173
rect 751 135 803 141
rect 751 101 760 135
rect 760 101 794 135
rect 794 101 803 135
rect 751 89 803 101
rect 751 29 760 61
rect 760 29 794 61
rect 794 29 803 61
rect 751 9 803 29
rect 751 -43 760 -19
rect 760 -43 794 -19
rect 794 -43 803 -19
rect 751 -71 803 -43
rect 751 -115 760 -99
rect 760 -115 794 -99
rect 794 -115 803 -99
rect 751 -151 803 -115
rect 751 -187 760 -179
rect 760 -187 794 -179
rect 794 -187 803 -179
rect 751 -225 803 -187
rect 751 -231 760 -225
rect 760 -231 794 -225
rect 794 -231 803 -225
rect 751 -297 803 -259
rect 751 -311 760 -297
rect 760 -311 794 -297
rect 794 -311 803 -297
rect 751 -369 803 -339
rect 751 -391 760 -369
rect 760 -391 794 -369
rect 794 -391 803 -369
rect 751 -441 803 -419
rect 751 -471 760 -441
rect 760 -471 794 -441
rect 794 -471 803 -441
rect 751 -513 803 -499
rect 751 -547 760 -513
rect 760 -547 794 -513
rect 794 -547 803 -513
rect 751 -551 803 -547
rect 751 -585 803 -579
rect 751 -619 760 -585
rect 760 -619 794 -585
rect 794 -619 803 -585
rect 751 -631 803 -619
rect -100 -1700 1200 -1200
rect -11600 -2900 -11400 -2700
<< metal2 >>
rect -6700 17260 -6600 18600
rect -6300 17260 -6200 18600
rect -5900 17260 -5800 18600
rect -5500 17260 -5400 18600
rect -6720 17240 -6500 17260
rect -6720 17160 -6700 17240
rect -6520 17160 -6500 17240
rect -6720 17140 -6500 17160
rect -6320 17240 -6100 17260
rect -6320 17160 -6300 17240
rect -6120 17160 -6100 17240
rect -6320 17140 -6100 17160
rect -5920 17240 -5700 17260
rect -5920 17160 -5900 17240
rect -5720 17160 -5700 17240
rect -5920 17140 -5700 17160
rect -5540 17240 -5320 17260
rect -5540 17160 -5520 17240
rect -5340 17160 -5320 17240
rect -5540 17140 -5320 17160
rect -4800 17100 -3300 17200
rect -6860 17088 -4700 17100
rect -6860 17036 -6634 17088
rect -6582 17036 -6240 17088
rect -6188 17036 -5846 17088
rect -5794 17036 -5452 17088
rect -5400 17036 -4700 17088
rect -6860 17024 -4700 17036
rect -6860 16972 -6634 17024
rect -6582 16972 -6240 17024
rect -6188 16972 -5846 17024
rect -5794 16972 -5452 17024
rect -5400 16972 -4700 17024
rect -6860 16960 -4700 16972
rect -6860 16908 -6634 16960
rect -6582 16908 -6240 16960
rect -6188 16908 -5846 16960
rect -5794 16908 -5452 16960
rect -5400 16908 -4700 16960
rect -6860 16896 -4700 16908
rect -6860 16844 -6634 16896
rect -6582 16844 -6240 16896
rect -6188 16844 -5846 16896
rect -5794 16844 -5452 16896
rect -5400 16844 -4700 16896
rect -6860 16832 -4700 16844
rect -6860 16780 -6634 16832
rect -6582 16780 -6240 16832
rect -6188 16780 -5846 16832
rect -5794 16780 -5452 16832
rect -5400 16780 -4700 16832
rect -6860 16768 -4700 16780
rect -6860 16716 -6634 16768
rect -6582 16716 -6240 16768
rect -6188 16716 -5846 16768
rect -5794 16716 -5452 16768
rect -5400 16716 -4700 16768
rect -6860 16704 -4700 16716
rect -6860 16652 -6634 16704
rect -6582 16652 -6240 16704
rect -6188 16652 -5846 16704
rect -5794 16652 -5452 16704
rect -5400 16652 -4700 16704
rect -6860 16620 -4700 16652
rect -5000 16600 -4700 16620
rect -3400 16600 -3300 17100
rect -6740 16542 -6480 16560
rect -6740 16490 -6720 16542
rect -6668 16490 -6548 16542
rect -6496 16490 -6480 16542
rect -6740 16478 -6480 16490
rect -6740 16426 -6720 16478
rect -6668 16426 -6548 16478
rect -6496 16426 -6480 16478
rect -6740 16414 -6480 16426
rect -6740 16362 -6720 16414
rect -6668 16362 -6548 16414
rect -6496 16362 -6480 16414
rect -6740 16360 -6480 16362
rect -6920 16350 -6480 16360
rect -6920 16320 -6720 16350
rect -6920 16020 -6900 16320
rect -6780 16298 -6720 16320
rect -6668 16298 -6548 16350
rect -6496 16298 -6480 16350
rect -6780 16286 -6480 16298
rect -6780 16234 -6720 16286
rect -6668 16234 -6548 16286
rect -6496 16234 -6480 16286
rect -6780 16222 -6480 16234
rect -6780 16170 -6720 16222
rect -6668 16170 -6548 16222
rect -6496 16170 -6480 16222
rect -6780 16158 -6480 16170
rect -6780 16106 -6720 16158
rect -6668 16106 -6548 16158
rect -6496 16106 -6480 16158
rect -6780 16020 -6480 16106
rect -6920 16000 -6480 16020
rect -6340 16542 -6080 16560
rect -6340 16490 -6326 16542
rect -6274 16490 -6154 16542
rect -6102 16490 -6080 16542
rect -6340 16478 -6080 16490
rect -6340 16426 -6326 16478
rect -6274 16426 -6154 16478
rect -6102 16426 -6080 16478
rect -6340 16414 -6080 16426
rect -6340 16362 -6326 16414
rect -6274 16362 -6154 16414
rect -6102 16362 -6080 16414
rect -6340 16350 -6080 16362
rect -6340 16298 -6326 16350
rect -6274 16298 -6154 16350
rect -6102 16298 -6080 16350
rect -6340 16286 -6080 16298
rect -6340 16234 -6326 16286
rect -6274 16234 -6154 16286
rect -6102 16234 -6080 16286
rect -6340 16222 -6080 16234
rect -6340 16170 -6326 16222
rect -6274 16170 -6154 16222
rect -6102 16170 -6080 16222
rect -6340 16158 -6080 16170
rect -6340 16106 -6326 16158
rect -6274 16106 -6154 16158
rect -6102 16106 -6080 16158
rect -6760 15900 -6440 15920
rect -6760 15820 -6740 15900
rect -6460 15820 -6440 15900
rect -6760 15800 -6440 15820
rect -6620 15080 -6460 15800
rect -6340 15780 -6080 16106
rect -5940 16542 -5680 16560
rect -5940 16490 -5932 16542
rect -5880 16540 -5760 16542
rect -5708 16540 -5680 16542
rect -5940 16478 -5920 16490
rect -5940 16426 -5932 16478
rect -5940 16414 -5920 16426
rect -5940 16362 -5932 16414
rect -5940 16350 -5920 16362
rect -5940 16298 -5932 16350
rect -5940 16286 -5920 16298
rect -5940 16234 -5932 16286
rect -5940 16222 -5920 16234
rect -5940 16170 -5932 16222
rect -5940 16158 -5920 16170
rect -5940 16106 -5932 16158
rect -5700 16120 -5680 16540
rect -5880 16106 -5760 16120
rect -5708 16106 -5680 16120
rect -5940 16080 -5680 16106
rect -5560 16542 -5300 16560
rect -5560 16490 -5538 16542
rect -5486 16490 -5366 16542
rect -5314 16490 -5300 16542
rect -4800 16500 -3300 16600
rect -5560 16478 -5300 16490
rect -5560 16426 -5538 16478
rect -5486 16426 -5366 16478
rect -5314 16426 -5300 16478
rect -5560 16414 -5300 16426
rect -5560 16362 -5538 16414
rect -5486 16362 -5366 16414
rect -5314 16362 -5300 16414
rect -5560 16360 -5300 16362
rect -5560 16350 -5100 16360
rect -5560 16298 -5538 16350
rect -5486 16298 -5366 16350
rect -5314 16340 -5100 16350
rect -5314 16298 -5260 16340
rect -5560 16286 -5260 16298
rect -5560 16234 -5538 16286
rect -5486 16234 -5366 16286
rect -5314 16234 -5260 16286
rect -5560 16222 -5260 16234
rect -5560 16170 -5538 16222
rect -5486 16170 -5366 16222
rect -5314 16170 -5260 16222
rect -5560 16158 -5260 16170
rect -5560 16106 -5538 16158
rect -5486 16106 -5366 16158
rect -5314 16106 -5260 16158
rect -5560 16020 -5260 16106
rect -5120 16020 -5100 16340
rect -5560 16000 -5100 16020
rect -6020 15900 -5260 15920
rect -6020 15820 -6000 15900
rect -5280 15820 -5260 15900
rect -6020 15800 -5260 15820
rect -6340 15620 -6320 15780
rect -6100 15620 -6080 15780
rect -6340 15600 -6080 15620
rect -5700 15080 -5420 15800
rect -6620 15000 -5420 15080
rect -6700 14400 -5300 15000
rect -9200 14200 -4400 14400
rect -9200 12600 -9000 14200
rect -15200 12400 -9000 12600
rect -15200 11600 -15000 12400
rect -4600 11600 -4400 14200
rect -15200 11400 -4400 11600
rect -15000 8000 -13200 11400
rect -12800 8000 -11800 11400
rect -11400 8000 -10600 11400
rect -10200 8000 -9400 11400
rect -9000 8000 -8200 11400
rect -7800 8000 -7000 11400
rect -6600 8000 -5800 11400
rect -5400 8600 -4400 11400
rect -800 12500 1000 12600
rect -800 9100 -700 12500
rect 900 9100 1000 12500
rect -800 9000 1000 9100
rect -5400 8000 -4700 8600
rect -15000 7800 -4700 8000
rect -4500 8000 -4400 8600
rect -50 8600 1000 9000
rect -50 8520 1036 8600
rect -50 8519 1033 8520
rect -50 8500 1000 8519
rect 31 8411 83 8500
rect 31 8331 83 8359
rect 31 8251 83 8279
rect 31 8171 83 8199
rect 31 8091 83 8119
rect 31 8011 83 8039
rect -4500 7800 -4200 8000
rect -15000 3200 -14800 7800
rect -4400 6200 -4200 7800
rect 31 7931 83 7959
rect 31 7851 83 7879
rect 31 7771 83 7799
rect -2000 7680 -1640 7700
rect -2000 7520 -1980 7680
rect -1660 7520 -1640 7680
rect -2000 7500 -1640 7520
rect 31 7691 83 7719
rect 31 7611 83 7639
rect 31 7489 83 7559
rect 203 8411 255 8500
rect 203 8331 255 8359
rect 203 8251 255 8279
rect 203 8171 255 8199
rect 203 8091 255 8119
rect 203 8011 255 8039
rect 203 7931 255 7959
rect 203 7851 255 7879
rect 203 7771 255 7799
rect 203 7691 255 7719
rect 203 7611 255 7639
rect 203 7489 255 7559
rect 375 8411 427 8500
rect 375 8331 427 8359
rect 375 8251 427 8279
rect 375 8171 427 8199
rect 375 8091 427 8119
rect 375 8011 427 8039
rect 375 7931 427 7959
rect 375 7851 427 7879
rect 375 7771 427 7799
rect 375 7691 427 7719
rect 375 7611 427 7639
rect 375 7489 427 7559
rect 547 8411 599 8500
rect 547 8331 599 8359
rect 547 8251 599 8279
rect 547 8171 599 8199
rect 547 8091 599 8119
rect 547 8011 599 8039
rect 547 7931 599 7959
rect 547 7851 599 7879
rect 547 7771 599 7799
rect 547 7691 599 7719
rect 547 7611 599 7639
rect 547 7489 599 7559
rect 719 8411 771 8500
rect 719 8331 771 8359
rect 719 8251 771 8279
rect 719 8171 771 8199
rect 719 8091 771 8119
rect 719 8011 771 8039
rect 719 7931 771 7959
rect 719 7851 771 7879
rect 719 7771 771 7799
rect 719 7691 771 7719
rect 719 7611 771 7639
rect 719 7489 771 7559
rect 891 8411 943 8500
rect 891 8331 943 8359
rect 891 8251 943 8279
rect 891 8171 943 8199
rect 891 8091 943 8119
rect 891 8011 943 8039
rect 891 7931 943 7959
rect 891 7851 943 7879
rect 891 7771 943 7799
rect 891 7691 943 7719
rect 891 7611 943 7639
rect 891 7489 943 7559
rect -34 7300 -14 7400
rect 996 7300 1016 7400
rect 0 7200 1000 7300
rect -2360 7180 -2140 7200
rect -2360 7110 -2350 7180
rect -2150 7110 -2140 7180
rect -2360 7060 -2140 7110
rect -1860 7180 -1640 7200
rect -1860 7110 -1850 7180
rect -1650 7110 -1640 7180
rect -1860 7060 -1640 7110
rect -2500 7050 -1500 7060
rect -2500 6850 -2480 7050
rect -2410 6850 -2090 7050
rect -2020 6850 -1980 7050
rect -1910 6850 -1590 7050
rect -1520 6850 -1500 7050
rect -2500 6840 -1500 6850
rect -1160 7020 -800 7040
rect -1160 6860 -1140 7020
rect -820 6860 -800 7020
rect -1160 6840 -800 6860
rect -2360 6790 -2140 6840
rect -2360 6720 -2350 6790
rect -2150 6720 -2140 6790
rect -2360 6680 -2140 6720
rect -2360 6610 -2350 6680
rect -2150 6610 -2140 6680
rect -2360 6560 -2140 6610
rect -1860 6790 -1640 6840
rect -1860 6720 -1850 6790
rect -1650 6720 -1640 6790
rect -1860 6680 -1640 6720
rect -1860 6610 -1850 6680
rect -1650 6610 -1640 6680
rect -1860 6560 -1640 6610
rect -2500 6550 -1500 6560
rect -2500 6350 -2480 6550
rect -2410 6350 -2090 6550
rect -2020 6350 -1980 6550
rect -1910 6350 -1590 6550
rect -1520 6350 -1500 6550
rect -2500 6340 -1500 6350
rect 0 6400 100 7200
rect 900 6400 1000 7200
rect -2360 6290 -2140 6340
rect -2360 6220 -2350 6290
rect -2150 6220 -2140 6290
rect -4400 6060 -4000 6200
rect -3860 6180 -3640 6200
rect -3860 6110 -3850 6180
rect -3650 6110 -3640 6180
rect -3860 6060 -3640 6110
rect -3360 6180 -3140 6200
rect -3360 6110 -3350 6180
rect -3150 6110 -3140 6180
rect -3360 6060 -3140 6110
rect -2860 6180 -2640 6200
rect -2860 6110 -2850 6180
rect -2650 6110 -2640 6180
rect -2860 6060 -2640 6110
rect -2360 6180 -2140 6220
rect -2360 6110 -2350 6180
rect -2150 6110 -2140 6180
rect -2360 6060 -2140 6110
rect -1860 6290 -1640 6340
rect 0 6300 1000 6400
rect -1860 6220 -1850 6290
rect -1650 6220 -1640 6290
rect -1860 6180 -1640 6220
rect -1860 6110 -1850 6180
rect -1650 6110 -1640 6180
rect -1860 6060 -1640 6110
rect -4400 6050 -1500 6060
rect -4400 5850 -3980 6050
rect -3910 5850 -3590 6050
rect -3520 5850 -3480 6050
rect -3410 5850 -3090 6050
rect -3020 5850 -2980 6050
rect -2910 5850 -2590 6050
rect -2520 5850 -2480 6050
rect -2410 5850 -2090 6050
rect -2020 5850 -1980 6050
rect -1910 5850 -1590 6050
rect -1520 5850 -1500 6050
rect -4400 5840 -1500 5850
rect -1200 5920 -840 5940
rect -4400 5600 -4000 5840
rect -3860 5790 -3640 5840
rect -3860 5720 -3850 5790
rect -3650 5720 -3640 5790
rect -3860 5680 -3640 5720
rect -3860 5610 -3850 5680
rect -3650 5610 -3640 5680
rect -3860 5600 -3640 5610
rect -4400 5560 -3640 5600
rect -3360 5790 -3140 5840
rect -3360 5720 -3350 5790
rect -3150 5720 -3140 5790
rect -3360 5680 -3140 5720
rect -3360 5610 -3350 5680
rect -3150 5610 -3140 5680
rect -3360 5560 -3140 5610
rect -2860 5790 -2640 5840
rect -2860 5720 -2850 5790
rect -2650 5720 -2640 5790
rect -2860 5680 -2640 5720
rect -2860 5610 -2850 5680
rect -2650 5610 -2640 5680
rect -2860 5560 -2640 5610
rect -2360 5790 -2140 5840
rect -2360 5720 -2350 5790
rect -2150 5720 -2140 5790
rect -2360 5680 -2140 5720
rect -1860 5790 -1640 5840
rect -1860 5720 -1850 5790
rect -1650 5720 -1640 5790
rect -1200 5760 -1180 5920
rect -860 5760 -840 5920
rect -1200 5740 -840 5760
rect -1860 5700 -1640 5720
rect -2360 5610 -2350 5680
rect -2150 5610 -2140 5680
rect -2360 5560 -2140 5610
rect -4400 5550 -2000 5560
rect -4400 5400 -3980 5550
rect -4000 5350 -3980 5400
rect -3910 5350 -3590 5550
rect -3520 5350 -3480 5550
rect -3410 5350 -3090 5550
rect -3020 5350 -2980 5550
rect -2910 5350 -2590 5550
rect -2520 5350 -2480 5550
rect -2410 5350 -2090 5550
rect -2020 5350 -2000 5550
rect -4000 5340 -2000 5350
rect -4000 5290 -3640 5340
rect -4000 5220 -3850 5290
rect -3650 5220 -3640 5290
rect -4000 5200 -3640 5220
rect -3360 5290 -3140 5340
rect -3360 5220 -3350 5290
rect -3150 5220 -3140 5290
rect -3360 5200 -3140 5220
rect -2860 5290 -2640 5340
rect -2860 5220 -2850 5290
rect -2650 5220 -2640 5290
rect -2860 5200 -2640 5220
rect -2360 5290 -2140 5340
rect -2360 5220 -2350 5290
rect -2150 5220 -2140 5290
rect -2360 5200 -2140 5220
rect -4000 3200 -3800 5200
rect -15000 3000 -3800 3200
rect 0 1200 1000 1300
rect 0 500 100 1200
rect 900 500 1000 1200
rect 0 460 1000 500
rect 0 400 170 460
rect 150 380 170 400
rect 870 400 1000 460
rect 870 380 890 400
rect 235 221 287 291
rect 235 141 287 169
rect 235 61 287 89
rect 235 -19 287 9
rect 235 -99 287 -71
rect 235 -179 287 -151
rect 235 -259 287 -231
rect 235 -339 287 -311
rect 235 -419 287 -391
rect 235 -499 287 -471
rect 235 -579 287 -551
rect -4320 -680 -4120 -660
rect -4320 -900 -4300 -680
rect -4140 -900 -4120 -680
rect -4320 -920 -4120 -900
rect -3980 -690 -3780 -670
rect -3980 -890 -3960 -690
rect -3800 -890 -3780 -690
rect 235 -700 287 -631
rect 407 221 459 291
rect 407 141 459 169
rect 407 61 459 89
rect 407 -19 459 9
rect 407 -99 459 -71
rect 407 -179 459 -151
rect 407 -259 459 -231
rect 407 -339 459 -311
rect 407 -419 459 -391
rect 407 -499 459 -471
rect 407 -579 459 -551
rect 407 -700 459 -631
rect 579 221 631 291
rect 579 141 631 169
rect 579 61 631 89
rect 579 -19 631 9
rect 579 -99 631 -71
rect 579 -179 631 -151
rect 579 -259 631 -231
rect 579 -339 631 -311
rect 579 -419 631 -391
rect 579 -499 631 -471
rect 579 -579 631 -551
rect 579 -700 631 -631
rect 751 221 803 291
rect 751 141 803 169
rect 751 61 803 89
rect 751 -19 803 9
rect 751 -99 803 -71
rect 751 -179 803 -151
rect 751 -259 803 -231
rect 751 -339 803 -311
rect 751 -419 803 -391
rect 751 -499 803 -471
rect 751 -579 803 -551
rect 751 -700 803 -631
rect -3980 -910 -3780 -890
rect -800 -1000 1900 -700
rect -12000 -1400 -11000 -1300
rect -12000 -3200 -11900 -1400
rect -11100 -3200 -11000 -1400
rect -12000 -3300 -11000 -3200
rect -800 -2200 -400 -1000
rect -200 -1200 1300 -1100
rect -200 -1700 -100 -1200
rect 1200 -1700 1300 -1200
rect -200 -1800 1300 -1700
rect 1500 -2200 1900 -1000
rect -800 -2300 1900 -2200
rect -800 -4700 -700 -2300
rect 1800 -4700 1900 -2300
rect -800 -4800 1900 -4700
<< via2 >>
rect -4700 16600 -3400 17100
rect -6900 16020 -6780 16320
rect -5920 16490 -5880 16540
rect -5880 16490 -5760 16540
rect -5760 16490 -5708 16540
rect -5708 16490 -5700 16540
rect -5920 16478 -5700 16490
rect -5920 16426 -5880 16478
rect -5880 16426 -5760 16478
rect -5760 16426 -5708 16478
rect -5708 16426 -5700 16478
rect -5920 16414 -5700 16426
rect -5920 16362 -5880 16414
rect -5880 16362 -5760 16414
rect -5760 16362 -5708 16414
rect -5708 16362 -5700 16414
rect -5920 16350 -5700 16362
rect -5920 16298 -5880 16350
rect -5880 16298 -5760 16350
rect -5760 16298 -5708 16350
rect -5708 16298 -5700 16350
rect -5920 16286 -5700 16298
rect -5920 16234 -5880 16286
rect -5880 16234 -5760 16286
rect -5760 16234 -5708 16286
rect -5708 16234 -5700 16286
rect -5920 16222 -5700 16234
rect -5920 16170 -5880 16222
rect -5880 16170 -5760 16222
rect -5760 16170 -5708 16222
rect -5708 16170 -5700 16222
rect -5920 16158 -5700 16170
rect -5920 16120 -5880 16158
rect -5880 16120 -5760 16158
rect -5760 16120 -5708 16158
rect -5708 16120 -5700 16158
rect -5260 16020 -5120 16340
rect -6320 15620 -6100 15780
rect -9000 12400 -4600 14200
rect -15000 11600 -4600 12400
rect -700 9100 900 12500
rect -14800 5400 -4400 7800
rect -1980 7520 -1820 7680
rect -1820 7520 -1660 7680
rect -1140 6860 -980 7020
rect -980 6860 -820 7020
rect 100 6400 900 7200
rect -1180 5760 -1020 5920
rect -1020 5760 -860 5920
rect -14800 3200 -4000 5400
rect 100 500 900 1200
rect -4300 -690 -4140 -680
rect -4300 -890 -4140 -690
rect -4300 -900 -4140 -890
rect -3960 -890 -3800 -690
rect -11900 -1700 -11100 -1400
rect -11900 -1900 -11600 -1700
rect -11600 -1900 -11400 -1700
rect -11400 -1900 -11100 -1700
rect -11900 -2200 -11100 -1900
rect -11900 -2400 -11600 -2200
rect -11600 -2400 -11400 -2200
rect -11400 -2400 -11100 -2200
rect -11900 -2700 -11100 -2400
rect -11900 -2900 -11600 -2700
rect -11600 -2900 -11400 -2700
rect -11400 -2900 -11100 -2700
rect -11900 -3200 -11100 -2900
rect -100 -1700 1200 -1200
rect -700 -4700 1800 -2300
<< metal3 >>
rect -18000 23700 -10400 23800
rect -18000 22400 -17900 23700
rect -10500 22400 -10400 23700
rect -18000 22000 -10400 22400
rect -20600 20000 -10400 22000
rect -20600 19800 -7600 20000
rect -20600 16600 -9000 19800
rect -7800 17600 -7600 19800
rect -4700 18400 1000 18500
rect -7800 16600 -7200 17600
rect -6860 17320 -5180 18400
rect -20600 16400 -7200 16600
rect -5960 16540 -5680 17320
rect -4700 17200 -4300 18400
rect -20600 13000 -10400 16400
rect -6920 16320 -6760 16400
rect -6920 16020 -6900 16320
rect -6780 16020 -6760 16320
rect -5960 16120 -5920 16540
rect -5700 16120 -5680 16540
rect -4800 17100 -4300 17200
rect -4800 16600 -4700 17100
rect 900 16600 1000 18400
rect -4800 16500 1000 16600
rect -5960 16100 -5680 16120
rect -5280 16340 -5100 16360
rect -6920 16000 -6760 16020
rect -5280 16020 -5260 16340
rect -5120 16020 -5100 16340
rect -5280 16000 -5100 16020
rect -7340 15120 -6760 16000
rect -6380 15780 -6080 15800
rect -6380 15620 -6320 15780
rect -6100 15640 -6080 15780
rect -6100 15620 -5800 15640
rect -6380 15160 -5800 15620
rect -5260 14920 -4380 16000
rect -9200 14200 -4400 14400
rect -9200 12600 -9000 14200
rect -18000 12400 -9000 12600
rect -18000 11600 -17800 12400
rect -4600 11600 -4400 14200
rect -18000 11400 -4400 11600
rect -800 12500 1000 12600
rect -800 9380 -700 12500
rect -1160 9100 -700 9380
rect 900 9100 1000 12500
rect -1160 9000 1000 9100
rect -3600 8150 -2600 8200
rect -15000 7800 -4200 8000
rect -15000 3200 -14800 7800
rect -4400 5600 -4200 7800
rect -3600 7850 -3550 8150
rect -2650 7850 -2600 8150
rect -3600 7750 -2600 7850
rect -3600 7700 -1650 7750
rect -3600 7680 -1640 7700
rect -3600 7520 -1980 7680
rect -1660 7520 -1640 7680
rect -3600 7500 -1640 7520
rect -3600 7400 -1650 7500
rect -3600 6000 -2600 7400
rect -1160 7020 -800 9000
rect 2300 8000 6500 8100
rect 2300 7400 2400 8000
rect -1160 6860 -1140 7020
rect -820 6860 -800 7020
rect -1160 6840 -800 6860
rect 0 7200 2400 7400
rect 0 6400 100 7200
rect 900 6600 2400 7200
rect 6400 6600 6500 8000
rect 900 6400 6500 6600
rect 0 6300 6500 6400
rect -1200 5920 200 6000
rect -1200 5760 -1180 5920
rect -860 5900 200 5920
rect -860 5800 -300 5900
rect -860 5760 -840 5800
rect -1200 5740 -840 5760
rect -4400 5400 -3800 5600
rect -4000 3200 -3800 5400
rect -15000 3000 -3800 3200
rect -5600 -50 -3600 2600
rect -3200 600 -800 5200
rect -400 4400 -300 5800
rect 100 4400 200 5900
rect -400 4200 200 4400
rect -3200 100 -3100 600
rect -900 100 -800 600
rect 0 1200 6700 1500
rect 0 500 100 1200
rect 900 500 2400 1200
rect 0 400 2400 500
rect -3200 0 -800 100
rect 2300 0 2400 400
rect 6600 0 6700 1200
rect -5600 -350 -5550 -50
rect -3650 -350 -3600 -50
rect -5600 -400 -3600 -350
rect -4320 -680 -4120 -660
rect -3950 -670 -3650 -400
rect -4320 -900 -4300 -680
rect -4140 -900 -4120 -680
rect -4320 -920 -4120 -900
rect -3980 -680 -3650 -670
rect -3000 -680 -1000 0
rect 2300 -100 6700 0
rect -3980 -690 -1000 -680
rect -3980 -890 -3960 -690
rect -3800 -890 -1000 -690
rect -3980 -910 -1000 -890
rect -3660 -920 -1000 -910
rect -3000 -1100 -1000 -920
rect -3000 -1200 2800 -1100
rect -12000 -1400 -11000 -1300
rect -12000 -3200 -11900 -1400
rect -11100 -3200 -11000 -1400
rect -3000 -1700 -100 -1200
rect 1200 -1700 2800 -1200
rect -3000 -1800 2800 -1700
rect -3000 -2000 -1000 -1800
rect -12000 -3300 -11000 -3200
rect -800 -2300 1900 -2200
rect -800 -4700 -700 -2300
rect 1800 -4700 1900 -2300
rect -800 -4800 1900 -4700
<< via3 >>
rect -17900 22400 -10500 23700
rect -9000 16600 -7800 19800
rect -4300 17100 900 18400
rect -4300 16600 -3400 17100
rect -3400 16600 900 17100
rect -9000 12400 -4600 14200
rect -17800 11600 -15000 12400
rect -15000 11600 -4600 12400
rect -700 9100 900 12500
rect -14800 5400 -4400 7800
rect -3550 7850 -2650 8150
rect 2400 6600 6400 8000
rect -14800 3200 -4000 5400
rect -300 4400 100 5900
rect -3100 100 -900 600
rect 2400 0 6600 1200
rect -5550 -350 -3650 -50
rect -11900 -3200 -11100 -1400
rect -700 -4700 1800 -2300
<< mimcap >>
rect -20500 21800 -10500 21900
rect -20500 13200 -20400 21800
rect -10600 13200 -10500 21800
rect -6820 18340 -5220 18360
rect -6820 17380 -6800 18340
rect -5240 17380 -5220 18340
rect -6820 17360 -5220 17380
rect -7300 15940 -6800 15960
rect -7300 15180 -7280 15940
rect -6820 15180 -6800 15940
rect -5220 15940 -4420 15960
rect -6340 15580 -5840 15600
rect -6340 15220 -6320 15580
rect -5860 15220 -5840 15580
rect -6340 15200 -5840 15220
rect -7300 15160 -6800 15180
rect -5220 14980 -5200 15940
rect -4440 14980 -4420 15940
rect -5220 14960 -4420 14980
rect -20500 13100 -10500 13200
rect -3550 7500 -2650 7550
rect -3550 6100 -3500 7500
rect -2700 6100 -2650 7500
rect -3550 6050 -2650 6100
rect -3150 5100 -850 5150
rect -5550 2500 -3650 2550
rect -5550 300 -5500 2500
rect -3700 300 -3650 2500
rect -3150 1100 -3100 5100
rect -900 1100 -850 5100
rect -3150 1050 -850 1100
rect -5550 250 -3650 300
<< mimcapcontact >>
rect -20400 13200 -10600 21800
rect -6800 17380 -5240 18340
rect -7280 15180 -6820 15940
rect -6320 15220 -5860 15580
rect -5200 14980 -4440 15940
rect -3500 6100 -2700 7500
rect -5500 300 -3700 2500
rect -3100 1100 -900 5100
<< metal4 >>
rect -18000 23700 -10400 23800
rect -18000 22400 -17900 23700
rect -10500 22400 -10400 23700
rect -18000 22300 -10400 22400
rect -20600 21800 -10400 22200
rect -20600 13200 -20400 21800
rect -10600 15600 -10400 21800
rect -9200 19800 -7600 20000
rect -9200 16600 -9000 19800
rect -7800 17600 -7600 19800
rect -3600 18500 1000 23300
rect -4400 18400 1000 18500
rect -6860 18340 -5180 18400
rect -6860 17660 -6800 18340
rect -7340 17600 -6800 17660
rect -7800 17380 -6800 17600
rect -5240 17380 -5180 18340
rect -7800 17320 -5180 17380
rect -7800 16600 -7020 17320
rect -9200 16400 -7020 16600
rect -4400 16600 -4300 18400
rect 900 16600 1000 18400
rect -4400 16500 1000 16600
rect -7340 16180 -4640 16400
rect -7340 16000 -7020 16180
rect -7340 15940 -6760 16000
rect -10600 14400 -8000 15600
rect -7340 15180 -7280 15940
rect -6820 15180 -6760 15940
rect -6020 15640 -5760 16180
rect -7340 15120 -6760 15180
rect -6380 15580 -5760 15640
rect -6380 15220 -6320 15580
rect -5860 15220 -5760 15580
rect -6380 15160 -5760 15220
rect -5260 16000 -4640 16180
rect -5260 15940 -4380 16000
rect -5260 14980 -5200 15940
rect -4440 14980 -4380 15940
rect -5260 14920 -4380 14980
rect -10600 14200 -4400 14400
rect -10600 13200 -9000 14200
rect -20600 12400 -9000 13200
rect -20600 11600 -17800 12400
rect -4600 11600 -4400 14200
rect -20600 11400 -4400 11600
rect -3600 12500 1000 16500
rect -3600 10800 -700 12500
rect -4000 10600 -700 10800
rect -21000 9100 -700 10600
rect 900 9100 1000 12500
rect -21000 9000 1000 9100
rect 2300 10100 6500 10200
rect -3600 8150 -2600 8200
rect -15000 7800 -4200 8000
rect -3600 7850 -3550 8150
rect -2650 7850 -2600 8150
rect -3600 7800 -2600 7850
rect 2300 8000 2600 10100
rect -15000 3200 -14800 7800
rect -4400 7600 -4200 7800
rect -4400 7500 -2600 7600
rect -4400 7300 -3500 7500
rect -4400 7100 -4200 7300
rect -3600 7100 -3500 7300
rect -4400 6900 -3500 7100
rect -4400 6700 -4200 6900
rect -3600 6700 -3500 6900
rect -4400 6500 -3500 6700
rect -4400 6300 -4200 6500
rect -3600 6300 -3500 6500
rect -4400 6100 -3500 6300
rect -2700 6100 -2600 7500
rect 2300 6600 2400 8000
rect 6400 6600 6500 10100
rect 2300 6500 6500 6600
rect -4400 6000 -2600 6100
rect -4400 5600 -4200 6000
rect -400 5900 200 6000
rect -4400 5400 -3800 5600
rect -4000 3200 -3800 5400
rect -400 5200 -300 5900
rect -15000 3000 -3800 3200
rect -5600 2600 -5400 3000
rect -5200 2600 -5000 3000
rect -4800 2600 -4600 3000
rect -4400 2600 -4200 3000
rect -4000 2600 -3800 3000
rect -3200 5100 -300 5200
rect -5600 2500 -3600 2600
rect -5600 300 -5500 2500
rect -3700 300 -3600 2500
rect -3200 1100 -3100 5100
rect -900 4400 -300 5100
rect 100 4400 200 5900
rect -900 4200 200 4400
rect -900 1100 -800 4200
rect -3200 1000 -800 1100
rect 2300 1200 11700 1300
rect -5600 200 -3600 300
rect -3200 600 -800 700
rect -3200 100 -3100 600
rect -900 100 -800 600
rect -3200 0 -800 100
rect 2300 0 2400 1200
rect 6600 0 11700 1200
rect -5600 -50 -3600 0
rect -5600 -350 -5550 -50
rect -3650 -350 -3600 -50
rect -5600 -400 -3600 -350
rect 2300 -600 11700 0
rect -12000 -1400 -11000 -1300
rect -12000 -3200 -11900 -1400
rect -11100 -3200 -11000 -1400
rect -12000 -3300 -11000 -3200
rect -800 -2300 1900 -2200
rect -800 -4700 -700 -2300
rect 1800 -4700 1900 -2300
rect -800 -5000 1900 -4700
<< via4 >>
rect -17900 22400 -10500 23700
rect -3550 7850 -2650 8150
rect 2600 8000 6400 10100
rect -14800 3200 -6200 7800
rect 2600 6900 6400 8000
rect -3100 100 -900 600
rect -5550 -350 -3650 -50
rect -11900 -3200 -11100 -1400
<< mimcap2 >>
rect -20500 21800 -10500 21900
rect -20500 13200 -20400 21800
rect -10600 13200 -10500 21800
rect -20500 13100 -10500 13200
rect -3550 7500 -2650 7550
rect -3550 6100 -3500 7500
rect -2700 6100 -2650 7500
rect -3550 6050 -2650 6100
rect -3150 5100 -850 5150
rect -5550 2500 -3650 2550
rect -5550 300 -5500 2500
rect -3700 300 -3650 2500
rect -3150 1100 -3100 5100
rect -900 1100 -850 5100
rect -3150 1050 -850 1100
rect -5550 250 -3650 300
<< mimcap2contact >>
rect -20400 13200 -10600 21800
rect -3500 6100 -2700 7500
rect -5500 300 -3700 2500
rect -3100 1100 -900 5100
<< metal5 >>
rect -19000 23800 -18400 23900
rect -20600 23700 -10400 23800
rect -20600 22400 -17900 23700
rect -10500 22400 -10400 23700
rect -20600 21800 -10400 22400
rect -20600 13200 -20400 21800
rect -10600 13200 -10400 21800
rect -20600 13000 -10400 13200
rect 2500 10100 6500 10200
rect -3600 8150 -2600 8200
rect -19800 7800 -6000 8000
rect -19800 5800 -14800 7800
rect -19800 3000 -15800 5800
rect -15000 3200 -14800 5800
rect -6200 3200 -6000 7800
rect -3600 7850 -3550 8150
rect -2650 7850 -2600 8150
rect -3600 7500 -2600 7850
rect -3600 6100 -3500 7500
rect -2700 6100 -2600 7500
rect 2500 6900 2600 10100
rect 6400 6900 6500 10100
rect 2500 6800 6500 6900
rect -3600 6000 -2600 6100
rect -15000 3000 -6000 3200
rect -3200 5100 -800 5200
rect -19800 800 -11000 3000
rect -19800 -2000 -15800 800
rect -15000 -1400 -11000 800
rect -5600 2500 -3600 2600
rect -5600 300 -5500 2500
rect -3700 300 -3600 2500
rect -5600 -50 -3600 300
rect -3200 1100 -3100 5100
rect -900 1100 -800 5100
rect -3200 600 -800 1100
rect -3200 100 -3100 600
rect -900 100 -800 600
rect -3200 0 -800 100
rect -5600 -350 -5550 -50
rect -3650 -350 -3600 -50
rect -5600 -400 -3600 -350
rect -15000 -2000 -11900 -1400
rect -19800 -3200 -11900 -2000
rect -11100 -3200 -11000 -1400
rect -800 -3000 1900 -2200
rect -19800 -4200 -11000 -3200
rect -19800 -7000 -15800 -4200
rect -15000 -7000 -11000 -4200
rect -19800 -9200 -11000 -7000
rect -19800 -12000 -15800 -9200
rect -15000 -12000 -11000 -9200
rect -19800 -14200 -11000 -12000
<< labels >>
rlabel metal5 -19800 6700 -15800 8000 1 VLO
rlabel metal5 -19000 23800 -18400 23900 1 VHI
rlabel metal4 -3600 22900 1000 23300 1 VOUT
rlabel metal4 -800 -5000 1900 -4800 1 SS
rlabel metal4 7200 -600 11700 1300 1 D1
rlabel metal4 2300 6500 6500 10200 1 S1
rlabel metal3 -2500 7400 -2200 7740 1 BIAS_TOP
rlabel metal3 -4300 -900 -4200 -700 1 BIAS_BOT
rlabel metal4 -400 4200 200 6000 1 RFB_MID
rlabel metal1 -1800 8600 -1600 8800 1 G_TOP
rlabel metal3 2400 -1800 2800 -1100 1 VIN
rlabel metal2 -5500 18500 -5400 18600 1 G4
rlabel metal2 -5900 18500 -5800 18600 1 G8
rlabel metal2 -6300 18500 -6200 18600 1 G1
rlabel metal2 -6700 18500 -6600 18600 1 G2
<< end >>
