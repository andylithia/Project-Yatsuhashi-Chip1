magic
tech sky130B
magscale 1 2
timestamp 1664070703
<< pwell >>
rect 0 0 5138 6516
rect 7000 0 12138 6516
rect 14000 0 19138 6516
rect 21000 0 26138 6516
rect 0 -7000 5138 -484
rect 7000 -7000 12138 -484
rect 14000 -7000 19138 -484
rect 21000 -7000 26138 -484
<< mvnmos >>
rect 228 258 328 6258
rect 386 258 486 6258
rect 544 258 644 6258
rect 702 258 802 6258
rect 860 258 960 6258
rect 1018 258 1118 6258
rect 1176 258 1276 6258
rect 1334 258 1434 6258
rect 1492 258 1592 6258
rect 1650 258 1750 6258
rect 1808 258 1908 6258
rect 1966 258 2066 6258
rect 2124 258 2224 6258
rect 2282 258 2382 6258
rect 2440 258 2540 6258
rect 2598 258 2698 6258
rect 2756 258 2856 6258
rect 2914 258 3014 6258
rect 3072 258 3172 6258
rect 3230 258 3330 6258
rect 3388 258 3488 6258
rect 3546 258 3646 6258
rect 3704 258 3804 6258
rect 3862 258 3962 6258
rect 4020 258 4120 6258
rect 4178 258 4278 6258
rect 4336 258 4436 6258
rect 4494 258 4594 6258
rect 4652 258 4752 6258
rect 4810 258 4910 6258
rect 7228 258 7328 6258
rect 7386 258 7486 6258
rect 7544 258 7644 6258
rect 7702 258 7802 6258
rect 7860 258 7960 6258
rect 8018 258 8118 6258
rect 8176 258 8276 6258
rect 8334 258 8434 6258
rect 8492 258 8592 6258
rect 8650 258 8750 6258
rect 8808 258 8908 6258
rect 8966 258 9066 6258
rect 9124 258 9224 6258
rect 9282 258 9382 6258
rect 9440 258 9540 6258
rect 9598 258 9698 6258
rect 9756 258 9856 6258
rect 9914 258 10014 6258
rect 10072 258 10172 6258
rect 10230 258 10330 6258
rect 10388 258 10488 6258
rect 10546 258 10646 6258
rect 10704 258 10804 6258
rect 10862 258 10962 6258
rect 11020 258 11120 6258
rect 11178 258 11278 6258
rect 11336 258 11436 6258
rect 11494 258 11594 6258
rect 11652 258 11752 6258
rect 11810 258 11910 6258
rect 14228 258 14328 6258
rect 14386 258 14486 6258
rect 14544 258 14644 6258
rect 14702 258 14802 6258
rect 14860 258 14960 6258
rect 15018 258 15118 6258
rect 15176 258 15276 6258
rect 15334 258 15434 6258
rect 15492 258 15592 6258
rect 15650 258 15750 6258
rect 15808 258 15908 6258
rect 15966 258 16066 6258
rect 16124 258 16224 6258
rect 16282 258 16382 6258
rect 16440 258 16540 6258
rect 16598 258 16698 6258
rect 16756 258 16856 6258
rect 16914 258 17014 6258
rect 17072 258 17172 6258
rect 17230 258 17330 6258
rect 17388 258 17488 6258
rect 17546 258 17646 6258
rect 17704 258 17804 6258
rect 17862 258 17962 6258
rect 18020 258 18120 6258
rect 18178 258 18278 6258
rect 18336 258 18436 6258
rect 18494 258 18594 6258
rect 18652 258 18752 6258
rect 18810 258 18910 6258
rect 21228 258 21328 6258
rect 21386 258 21486 6258
rect 21544 258 21644 6258
rect 21702 258 21802 6258
rect 21860 258 21960 6258
rect 22018 258 22118 6258
rect 22176 258 22276 6258
rect 22334 258 22434 6258
rect 22492 258 22592 6258
rect 22650 258 22750 6258
rect 22808 258 22908 6258
rect 22966 258 23066 6258
rect 23124 258 23224 6258
rect 23282 258 23382 6258
rect 23440 258 23540 6258
rect 23598 258 23698 6258
rect 23756 258 23856 6258
rect 23914 258 24014 6258
rect 24072 258 24172 6258
rect 24230 258 24330 6258
rect 24388 258 24488 6258
rect 24546 258 24646 6258
rect 24704 258 24804 6258
rect 24862 258 24962 6258
rect 25020 258 25120 6258
rect 25178 258 25278 6258
rect 25336 258 25436 6258
rect 25494 258 25594 6258
rect 25652 258 25752 6258
rect 25810 258 25910 6258
rect 228 -6742 328 -742
rect 386 -6742 486 -742
rect 544 -6742 644 -742
rect 702 -6742 802 -742
rect 860 -6742 960 -742
rect 1018 -6742 1118 -742
rect 1176 -6742 1276 -742
rect 1334 -6742 1434 -742
rect 1492 -6742 1592 -742
rect 1650 -6742 1750 -742
rect 1808 -6742 1908 -742
rect 1966 -6742 2066 -742
rect 2124 -6742 2224 -742
rect 2282 -6742 2382 -742
rect 2440 -6742 2540 -742
rect 2598 -6742 2698 -742
rect 2756 -6742 2856 -742
rect 2914 -6742 3014 -742
rect 3072 -6742 3172 -742
rect 3230 -6742 3330 -742
rect 3388 -6742 3488 -742
rect 3546 -6742 3646 -742
rect 3704 -6742 3804 -742
rect 3862 -6742 3962 -742
rect 4020 -6742 4120 -742
rect 4178 -6742 4278 -742
rect 4336 -6742 4436 -742
rect 4494 -6742 4594 -742
rect 4652 -6742 4752 -742
rect 4810 -6742 4910 -742
rect 7228 -6742 7328 -742
rect 7386 -6742 7486 -742
rect 7544 -6742 7644 -742
rect 7702 -6742 7802 -742
rect 7860 -6742 7960 -742
rect 8018 -6742 8118 -742
rect 8176 -6742 8276 -742
rect 8334 -6742 8434 -742
rect 8492 -6742 8592 -742
rect 8650 -6742 8750 -742
rect 8808 -6742 8908 -742
rect 8966 -6742 9066 -742
rect 9124 -6742 9224 -742
rect 9282 -6742 9382 -742
rect 9440 -6742 9540 -742
rect 9598 -6742 9698 -742
rect 9756 -6742 9856 -742
rect 9914 -6742 10014 -742
rect 10072 -6742 10172 -742
rect 10230 -6742 10330 -742
rect 10388 -6742 10488 -742
rect 10546 -6742 10646 -742
rect 10704 -6742 10804 -742
rect 10862 -6742 10962 -742
rect 11020 -6742 11120 -742
rect 11178 -6742 11278 -742
rect 11336 -6742 11436 -742
rect 11494 -6742 11594 -742
rect 11652 -6742 11752 -742
rect 11810 -6742 11910 -742
rect 14228 -6742 14328 -742
rect 14386 -6742 14486 -742
rect 14544 -6742 14644 -742
rect 14702 -6742 14802 -742
rect 14860 -6742 14960 -742
rect 15018 -6742 15118 -742
rect 15176 -6742 15276 -742
rect 15334 -6742 15434 -742
rect 15492 -6742 15592 -742
rect 15650 -6742 15750 -742
rect 15808 -6742 15908 -742
rect 15966 -6742 16066 -742
rect 16124 -6742 16224 -742
rect 16282 -6742 16382 -742
rect 16440 -6742 16540 -742
rect 16598 -6742 16698 -742
rect 16756 -6742 16856 -742
rect 16914 -6742 17014 -742
rect 17072 -6742 17172 -742
rect 17230 -6742 17330 -742
rect 17388 -6742 17488 -742
rect 17546 -6742 17646 -742
rect 17704 -6742 17804 -742
rect 17862 -6742 17962 -742
rect 18020 -6742 18120 -742
rect 18178 -6742 18278 -742
rect 18336 -6742 18436 -742
rect 18494 -6742 18594 -742
rect 18652 -6742 18752 -742
rect 18810 -6742 18910 -742
rect 21228 -6742 21328 -742
rect 21386 -6742 21486 -742
rect 21544 -6742 21644 -742
rect 21702 -6742 21802 -742
rect 21860 -6742 21960 -742
rect 22018 -6742 22118 -742
rect 22176 -6742 22276 -742
rect 22334 -6742 22434 -742
rect 22492 -6742 22592 -742
rect 22650 -6742 22750 -742
rect 22808 -6742 22908 -742
rect 22966 -6742 23066 -742
rect 23124 -6742 23224 -742
rect 23282 -6742 23382 -742
rect 23440 -6742 23540 -742
rect 23598 -6742 23698 -742
rect 23756 -6742 23856 -742
rect 23914 -6742 24014 -742
rect 24072 -6742 24172 -742
rect 24230 -6742 24330 -742
rect 24388 -6742 24488 -742
rect 24546 -6742 24646 -742
rect 24704 -6742 24804 -742
rect 24862 -6742 24962 -742
rect 25020 -6742 25120 -742
rect 25178 -6742 25278 -742
rect 25336 -6742 25436 -742
rect 25494 -6742 25594 -742
rect 25652 -6742 25752 -742
rect 25810 -6742 25910 -742
<< mvndiff >>
rect 170 6246 228 6258
rect 170 270 182 6246
rect 216 270 228 6246
rect 170 258 228 270
rect 328 6246 386 6258
rect 328 270 340 6246
rect 374 270 386 6246
rect 328 258 386 270
rect 486 6246 544 6258
rect 486 270 498 6246
rect 532 270 544 6246
rect 486 258 544 270
rect 644 6246 702 6258
rect 644 270 656 6246
rect 690 270 702 6246
rect 644 258 702 270
rect 802 6246 860 6258
rect 802 270 814 6246
rect 848 270 860 6246
rect 802 258 860 270
rect 960 6246 1018 6258
rect 960 270 972 6246
rect 1006 270 1018 6246
rect 960 258 1018 270
rect 1118 6246 1176 6258
rect 1118 270 1130 6246
rect 1164 270 1176 6246
rect 1118 258 1176 270
rect 1276 6246 1334 6258
rect 1276 270 1288 6246
rect 1322 270 1334 6246
rect 1276 258 1334 270
rect 1434 6246 1492 6258
rect 1434 270 1446 6246
rect 1480 270 1492 6246
rect 1434 258 1492 270
rect 1592 6246 1650 6258
rect 1592 270 1604 6246
rect 1638 270 1650 6246
rect 1592 258 1650 270
rect 1750 6246 1808 6258
rect 1750 270 1762 6246
rect 1796 270 1808 6246
rect 1750 258 1808 270
rect 1908 6246 1966 6258
rect 1908 270 1920 6246
rect 1954 270 1966 6246
rect 1908 258 1966 270
rect 2066 6246 2124 6258
rect 2066 270 2078 6246
rect 2112 270 2124 6246
rect 2066 258 2124 270
rect 2224 6246 2282 6258
rect 2224 270 2236 6246
rect 2270 270 2282 6246
rect 2224 258 2282 270
rect 2382 6246 2440 6258
rect 2382 270 2394 6246
rect 2428 270 2440 6246
rect 2382 258 2440 270
rect 2540 6246 2598 6258
rect 2540 270 2552 6246
rect 2586 270 2598 6246
rect 2540 258 2598 270
rect 2698 6246 2756 6258
rect 2698 270 2710 6246
rect 2744 270 2756 6246
rect 2698 258 2756 270
rect 2856 6246 2914 6258
rect 2856 270 2868 6246
rect 2902 270 2914 6246
rect 2856 258 2914 270
rect 3014 6246 3072 6258
rect 3014 270 3026 6246
rect 3060 270 3072 6246
rect 3014 258 3072 270
rect 3172 6246 3230 6258
rect 3172 270 3184 6246
rect 3218 270 3230 6246
rect 3172 258 3230 270
rect 3330 6246 3388 6258
rect 3330 270 3342 6246
rect 3376 270 3388 6246
rect 3330 258 3388 270
rect 3488 6246 3546 6258
rect 3488 270 3500 6246
rect 3534 270 3546 6246
rect 3488 258 3546 270
rect 3646 6246 3704 6258
rect 3646 270 3658 6246
rect 3692 270 3704 6246
rect 3646 258 3704 270
rect 3804 6246 3862 6258
rect 3804 270 3816 6246
rect 3850 270 3862 6246
rect 3804 258 3862 270
rect 3962 6246 4020 6258
rect 3962 270 3974 6246
rect 4008 270 4020 6246
rect 3962 258 4020 270
rect 4120 6246 4178 6258
rect 4120 270 4132 6246
rect 4166 270 4178 6246
rect 4120 258 4178 270
rect 4278 6246 4336 6258
rect 4278 270 4290 6246
rect 4324 270 4336 6246
rect 4278 258 4336 270
rect 4436 6246 4494 6258
rect 4436 270 4448 6246
rect 4482 270 4494 6246
rect 4436 258 4494 270
rect 4594 6246 4652 6258
rect 4594 270 4606 6246
rect 4640 270 4652 6246
rect 4594 258 4652 270
rect 4752 6246 4810 6258
rect 4752 270 4764 6246
rect 4798 270 4810 6246
rect 4752 258 4810 270
rect 4910 6246 4968 6258
rect 4910 270 4922 6246
rect 4956 270 4968 6246
rect 4910 258 4968 270
rect 7170 6246 7228 6258
rect 7170 270 7182 6246
rect 7216 270 7228 6246
rect 7170 258 7228 270
rect 7328 6246 7386 6258
rect 7328 270 7340 6246
rect 7374 270 7386 6246
rect 7328 258 7386 270
rect 7486 6246 7544 6258
rect 7486 270 7498 6246
rect 7532 270 7544 6246
rect 7486 258 7544 270
rect 7644 6246 7702 6258
rect 7644 270 7656 6246
rect 7690 270 7702 6246
rect 7644 258 7702 270
rect 7802 6246 7860 6258
rect 7802 270 7814 6246
rect 7848 270 7860 6246
rect 7802 258 7860 270
rect 7960 6246 8018 6258
rect 7960 270 7972 6246
rect 8006 270 8018 6246
rect 7960 258 8018 270
rect 8118 6246 8176 6258
rect 8118 270 8130 6246
rect 8164 270 8176 6246
rect 8118 258 8176 270
rect 8276 6246 8334 6258
rect 8276 270 8288 6246
rect 8322 270 8334 6246
rect 8276 258 8334 270
rect 8434 6246 8492 6258
rect 8434 270 8446 6246
rect 8480 270 8492 6246
rect 8434 258 8492 270
rect 8592 6246 8650 6258
rect 8592 270 8604 6246
rect 8638 270 8650 6246
rect 8592 258 8650 270
rect 8750 6246 8808 6258
rect 8750 270 8762 6246
rect 8796 270 8808 6246
rect 8750 258 8808 270
rect 8908 6246 8966 6258
rect 8908 270 8920 6246
rect 8954 270 8966 6246
rect 8908 258 8966 270
rect 9066 6246 9124 6258
rect 9066 270 9078 6246
rect 9112 270 9124 6246
rect 9066 258 9124 270
rect 9224 6246 9282 6258
rect 9224 270 9236 6246
rect 9270 270 9282 6246
rect 9224 258 9282 270
rect 9382 6246 9440 6258
rect 9382 270 9394 6246
rect 9428 270 9440 6246
rect 9382 258 9440 270
rect 9540 6246 9598 6258
rect 9540 270 9552 6246
rect 9586 270 9598 6246
rect 9540 258 9598 270
rect 9698 6246 9756 6258
rect 9698 270 9710 6246
rect 9744 270 9756 6246
rect 9698 258 9756 270
rect 9856 6246 9914 6258
rect 9856 270 9868 6246
rect 9902 270 9914 6246
rect 9856 258 9914 270
rect 10014 6246 10072 6258
rect 10014 270 10026 6246
rect 10060 270 10072 6246
rect 10014 258 10072 270
rect 10172 6246 10230 6258
rect 10172 270 10184 6246
rect 10218 270 10230 6246
rect 10172 258 10230 270
rect 10330 6246 10388 6258
rect 10330 270 10342 6246
rect 10376 270 10388 6246
rect 10330 258 10388 270
rect 10488 6246 10546 6258
rect 10488 270 10500 6246
rect 10534 270 10546 6246
rect 10488 258 10546 270
rect 10646 6246 10704 6258
rect 10646 270 10658 6246
rect 10692 270 10704 6246
rect 10646 258 10704 270
rect 10804 6246 10862 6258
rect 10804 270 10816 6246
rect 10850 270 10862 6246
rect 10804 258 10862 270
rect 10962 6246 11020 6258
rect 10962 270 10974 6246
rect 11008 270 11020 6246
rect 10962 258 11020 270
rect 11120 6246 11178 6258
rect 11120 270 11132 6246
rect 11166 270 11178 6246
rect 11120 258 11178 270
rect 11278 6246 11336 6258
rect 11278 270 11290 6246
rect 11324 270 11336 6246
rect 11278 258 11336 270
rect 11436 6246 11494 6258
rect 11436 270 11448 6246
rect 11482 270 11494 6246
rect 11436 258 11494 270
rect 11594 6246 11652 6258
rect 11594 270 11606 6246
rect 11640 270 11652 6246
rect 11594 258 11652 270
rect 11752 6246 11810 6258
rect 11752 270 11764 6246
rect 11798 270 11810 6246
rect 11752 258 11810 270
rect 11910 6246 11968 6258
rect 11910 270 11922 6246
rect 11956 270 11968 6246
rect 11910 258 11968 270
rect 14170 6246 14228 6258
rect 14170 270 14182 6246
rect 14216 270 14228 6246
rect 14170 258 14228 270
rect 14328 6246 14386 6258
rect 14328 270 14340 6246
rect 14374 270 14386 6246
rect 14328 258 14386 270
rect 14486 6246 14544 6258
rect 14486 270 14498 6246
rect 14532 270 14544 6246
rect 14486 258 14544 270
rect 14644 6246 14702 6258
rect 14644 270 14656 6246
rect 14690 270 14702 6246
rect 14644 258 14702 270
rect 14802 6246 14860 6258
rect 14802 270 14814 6246
rect 14848 270 14860 6246
rect 14802 258 14860 270
rect 14960 6246 15018 6258
rect 14960 270 14972 6246
rect 15006 270 15018 6246
rect 14960 258 15018 270
rect 15118 6246 15176 6258
rect 15118 270 15130 6246
rect 15164 270 15176 6246
rect 15118 258 15176 270
rect 15276 6246 15334 6258
rect 15276 270 15288 6246
rect 15322 270 15334 6246
rect 15276 258 15334 270
rect 15434 6246 15492 6258
rect 15434 270 15446 6246
rect 15480 270 15492 6246
rect 15434 258 15492 270
rect 15592 6246 15650 6258
rect 15592 270 15604 6246
rect 15638 270 15650 6246
rect 15592 258 15650 270
rect 15750 6246 15808 6258
rect 15750 270 15762 6246
rect 15796 270 15808 6246
rect 15750 258 15808 270
rect 15908 6246 15966 6258
rect 15908 270 15920 6246
rect 15954 270 15966 6246
rect 15908 258 15966 270
rect 16066 6246 16124 6258
rect 16066 270 16078 6246
rect 16112 270 16124 6246
rect 16066 258 16124 270
rect 16224 6246 16282 6258
rect 16224 270 16236 6246
rect 16270 270 16282 6246
rect 16224 258 16282 270
rect 16382 6246 16440 6258
rect 16382 270 16394 6246
rect 16428 270 16440 6246
rect 16382 258 16440 270
rect 16540 6246 16598 6258
rect 16540 270 16552 6246
rect 16586 270 16598 6246
rect 16540 258 16598 270
rect 16698 6246 16756 6258
rect 16698 270 16710 6246
rect 16744 270 16756 6246
rect 16698 258 16756 270
rect 16856 6246 16914 6258
rect 16856 270 16868 6246
rect 16902 270 16914 6246
rect 16856 258 16914 270
rect 17014 6246 17072 6258
rect 17014 270 17026 6246
rect 17060 270 17072 6246
rect 17014 258 17072 270
rect 17172 6246 17230 6258
rect 17172 270 17184 6246
rect 17218 270 17230 6246
rect 17172 258 17230 270
rect 17330 6246 17388 6258
rect 17330 270 17342 6246
rect 17376 270 17388 6246
rect 17330 258 17388 270
rect 17488 6246 17546 6258
rect 17488 270 17500 6246
rect 17534 270 17546 6246
rect 17488 258 17546 270
rect 17646 6246 17704 6258
rect 17646 270 17658 6246
rect 17692 270 17704 6246
rect 17646 258 17704 270
rect 17804 6246 17862 6258
rect 17804 270 17816 6246
rect 17850 270 17862 6246
rect 17804 258 17862 270
rect 17962 6246 18020 6258
rect 17962 270 17974 6246
rect 18008 270 18020 6246
rect 17962 258 18020 270
rect 18120 6246 18178 6258
rect 18120 270 18132 6246
rect 18166 270 18178 6246
rect 18120 258 18178 270
rect 18278 6246 18336 6258
rect 18278 270 18290 6246
rect 18324 270 18336 6246
rect 18278 258 18336 270
rect 18436 6246 18494 6258
rect 18436 270 18448 6246
rect 18482 270 18494 6246
rect 18436 258 18494 270
rect 18594 6246 18652 6258
rect 18594 270 18606 6246
rect 18640 270 18652 6246
rect 18594 258 18652 270
rect 18752 6246 18810 6258
rect 18752 270 18764 6246
rect 18798 270 18810 6246
rect 18752 258 18810 270
rect 18910 6246 18968 6258
rect 18910 270 18922 6246
rect 18956 270 18968 6246
rect 18910 258 18968 270
rect 21170 6246 21228 6258
rect 21170 270 21182 6246
rect 21216 270 21228 6246
rect 21170 258 21228 270
rect 21328 6246 21386 6258
rect 21328 270 21340 6246
rect 21374 270 21386 6246
rect 21328 258 21386 270
rect 21486 6246 21544 6258
rect 21486 270 21498 6246
rect 21532 270 21544 6246
rect 21486 258 21544 270
rect 21644 6246 21702 6258
rect 21644 270 21656 6246
rect 21690 270 21702 6246
rect 21644 258 21702 270
rect 21802 6246 21860 6258
rect 21802 270 21814 6246
rect 21848 270 21860 6246
rect 21802 258 21860 270
rect 21960 6246 22018 6258
rect 21960 270 21972 6246
rect 22006 270 22018 6246
rect 21960 258 22018 270
rect 22118 6246 22176 6258
rect 22118 270 22130 6246
rect 22164 270 22176 6246
rect 22118 258 22176 270
rect 22276 6246 22334 6258
rect 22276 270 22288 6246
rect 22322 270 22334 6246
rect 22276 258 22334 270
rect 22434 6246 22492 6258
rect 22434 270 22446 6246
rect 22480 270 22492 6246
rect 22434 258 22492 270
rect 22592 6246 22650 6258
rect 22592 270 22604 6246
rect 22638 270 22650 6246
rect 22592 258 22650 270
rect 22750 6246 22808 6258
rect 22750 270 22762 6246
rect 22796 270 22808 6246
rect 22750 258 22808 270
rect 22908 6246 22966 6258
rect 22908 270 22920 6246
rect 22954 270 22966 6246
rect 22908 258 22966 270
rect 23066 6246 23124 6258
rect 23066 270 23078 6246
rect 23112 270 23124 6246
rect 23066 258 23124 270
rect 23224 6246 23282 6258
rect 23224 270 23236 6246
rect 23270 270 23282 6246
rect 23224 258 23282 270
rect 23382 6246 23440 6258
rect 23382 270 23394 6246
rect 23428 270 23440 6246
rect 23382 258 23440 270
rect 23540 6246 23598 6258
rect 23540 270 23552 6246
rect 23586 270 23598 6246
rect 23540 258 23598 270
rect 23698 6246 23756 6258
rect 23698 270 23710 6246
rect 23744 270 23756 6246
rect 23698 258 23756 270
rect 23856 6246 23914 6258
rect 23856 270 23868 6246
rect 23902 270 23914 6246
rect 23856 258 23914 270
rect 24014 6246 24072 6258
rect 24014 270 24026 6246
rect 24060 270 24072 6246
rect 24014 258 24072 270
rect 24172 6246 24230 6258
rect 24172 270 24184 6246
rect 24218 270 24230 6246
rect 24172 258 24230 270
rect 24330 6246 24388 6258
rect 24330 270 24342 6246
rect 24376 270 24388 6246
rect 24330 258 24388 270
rect 24488 6246 24546 6258
rect 24488 270 24500 6246
rect 24534 270 24546 6246
rect 24488 258 24546 270
rect 24646 6246 24704 6258
rect 24646 270 24658 6246
rect 24692 270 24704 6246
rect 24646 258 24704 270
rect 24804 6246 24862 6258
rect 24804 270 24816 6246
rect 24850 270 24862 6246
rect 24804 258 24862 270
rect 24962 6246 25020 6258
rect 24962 270 24974 6246
rect 25008 270 25020 6246
rect 24962 258 25020 270
rect 25120 6246 25178 6258
rect 25120 270 25132 6246
rect 25166 270 25178 6246
rect 25120 258 25178 270
rect 25278 6246 25336 6258
rect 25278 270 25290 6246
rect 25324 270 25336 6246
rect 25278 258 25336 270
rect 25436 6246 25494 6258
rect 25436 270 25448 6246
rect 25482 270 25494 6246
rect 25436 258 25494 270
rect 25594 6246 25652 6258
rect 25594 270 25606 6246
rect 25640 270 25652 6246
rect 25594 258 25652 270
rect 25752 6246 25810 6258
rect 25752 270 25764 6246
rect 25798 270 25810 6246
rect 25752 258 25810 270
rect 25910 6246 25968 6258
rect 25910 270 25922 6246
rect 25956 270 25968 6246
rect 25910 258 25968 270
rect 170 -754 228 -742
rect 170 -6730 182 -754
rect 216 -6730 228 -754
rect 170 -6742 228 -6730
rect 328 -754 386 -742
rect 328 -6730 340 -754
rect 374 -6730 386 -754
rect 328 -6742 386 -6730
rect 486 -754 544 -742
rect 486 -6730 498 -754
rect 532 -6730 544 -754
rect 486 -6742 544 -6730
rect 644 -754 702 -742
rect 644 -6730 656 -754
rect 690 -6730 702 -754
rect 644 -6742 702 -6730
rect 802 -754 860 -742
rect 802 -6730 814 -754
rect 848 -6730 860 -754
rect 802 -6742 860 -6730
rect 960 -754 1018 -742
rect 960 -6730 972 -754
rect 1006 -6730 1018 -754
rect 960 -6742 1018 -6730
rect 1118 -754 1176 -742
rect 1118 -6730 1130 -754
rect 1164 -6730 1176 -754
rect 1118 -6742 1176 -6730
rect 1276 -754 1334 -742
rect 1276 -6730 1288 -754
rect 1322 -6730 1334 -754
rect 1276 -6742 1334 -6730
rect 1434 -754 1492 -742
rect 1434 -6730 1446 -754
rect 1480 -6730 1492 -754
rect 1434 -6742 1492 -6730
rect 1592 -754 1650 -742
rect 1592 -6730 1604 -754
rect 1638 -6730 1650 -754
rect 1592 -6742 1650 -6730
rect 1750 -754 1808 -742
rect 1750 -6730 1762 -754
rect 1796 -6730 1808 -754
rect 1750 -6742 1808 -6730
rect 1908 -754 1966 -742
rect 1908 -6730 1920 -754
rect 1954 -6730 1966 -754
rect 1908 -6742 1966 -6730
rect 2066 -754 2124 -742
rect 2066 -6730 2078 -754
rect 2112 -6730 2124 -754
rect 2066 -6742 2124 -6730
rect 2224 -754 2282 -742
rect 2224 -6730 2236 -754
rect 2270 -6730 2282 -754
rect 2224 -6742 2282 -6730
rect 2382 -754 2440 -742
rect 2382 -6730 2394 -754
rect 2428 -6730 2440 -754
rect 2382 -6742 2440 -6730
rect 2540 -754 2598 -742
rect 2540 -6730 2552 -754
rect 2586 -6730 2598 -754
rect 2540 -6742 2598 -6730
rect 2698 -754 2756 -742
rect 2698 -6730 2710 -754
rect 2744 -6730 2756 -754
rect 2698 -6742 2756 -6730
rect 2856 -754 2914 -742
rect 2856 -6730 2868 -754
rect 2902 -6730 2914 -754
rect 2856 -6742 2914 -6730
rect 3014 -754 3072 -742
rect 3014 -6730 3026 -754
rect 3060 -6730 3072 -754
rect 3014 -6742 3072 -6730
rect 3172 -754 3230 -742
rect 3172 -6730 3184 -754
rect 3218 -6730 3230 -754
rect 3172 -6742 3230 -6730
rect 3330 -754 3388 -742
rect 3330 -6730 3342 -754
rect 3376 -6730 3388 -754
rect 3330 -6742 3388 -6730
rect 3488 -754 3546 -742
rect 3488 -6730 3500 -754
rect 3534 -6730 3546 -754
rect 3488 -6742 3546 -6730
rect 3646 -754 3704 -742
rect 3646 -6730 3658 -754
rect 3692 -6730 3704 -754
rect 3646 -6742 3704 -6730
rect 3804 -754 3862 -742
rect 3804 -6730 3816 -754
rect 3850 -6730 3862 -754
rect 3804 -6742 3862 -6730
rect 3962 -754 4020 -742
rect 3962 -6730 3974 -754
rect 4008 -6730 4020 -754
rect 3962 -6742 4020 -6730
rect 4120 -754 4178 -742
rect 4120 -6730 4132 -754
rect 4166 -6730 4178 -754
rect 4120 -6742 4178 -6730
rect 4278 -754 4336 -742
rect 4278 -6730 4290 -754
rect 4324 -6730 4336 -754
rect 4278 -6742 4336 -6730
rect 4436 -754 4494 -742
rect 4436 -6730 4448 -754
rect 4482 -6730 4494 -754
rect 4436 -6742 4494 -6730
rect 4594 -754 4652 -742
rect 4594 -6730 4606 -754
rect 4640 -6730 4652 -754
rect 4594 -6742 4652 -6730
rect 4752 -754 4810 -742
rect 4752 -6730 4764 -754
rect 4798 -6730 4810 -754
rect 4752 -6742 4810 -6730
rect 4910 -754 4968 -742
rect 4910 -6730 4922 -754
rect 4956 -6730 4968 -754
rect 4910 -6742 4968 -6730
rect 7170 -754 7228 -742
rect 7170 -6730 7182 -754
rect 7216 -6730 7228 -754
rect 7170 -6742 7228 -6730
rect 7328 -754 7386 -742
rect 7328 -6730 7340 -754
rect 7374 -6730 7386 -754
rect 7328 -6742 7386 -6730
rect 7486 -754 7544 -742
rect 7486 -6730 7498 -754
rect 7532 -6730 7544 -754
rect 7486 -6742 7544 -6730
rect 7644 -754 7702 -742
rect 7644 -6730 7656 -754
rect 7690 -6730 7702 -754
rect 7644 -6742 7702 -6730
rect 7802 -754 7860 -742
rect 7802 -6730 7814 -754
rect 7848 -6730 7860 -754
rect 7802 -6742 7860 -6730
rect 7960 -754 8018 -742
rect 7960 -6730 7972 -754
rect 8006 -6730 8018 -754
rect 7960 -6742 8018 -6730
rect 8118 -754 8176 -742
rect 8118 -6730 8130 -754
rect 8164 -6730 8176 -754
rect 8118 -6742 8176 -6730
rect 8276 -754 8334 -742
rect 8276 -6730 8288 -754
rect 8322 -6730 8334 -754
rect 8276 -6742 8334 -6730
rect 8434 -754 8492 -742
rect 8434 -6730 8446 -754
rect 8480 -6730 8492 -754
rect 8434 -6742 8492 -6730
rect 8592 -754 8650 -742
rect 8592 -6730 8604 -754
rect 8638 -6730 8650 -754
rect 8592 -6742 8650 -6730
rect 8750 -754 8808 -742
rect 8750 -6730 8762 -754
rect 8796 -6730 8808 -754
rect 8750 -6742 8808 -6730
rect 8908 -754 8966 -742
rect 8908 -6730 8920 -754
rect 8954 -6730 8966 -754
rect 8908 -6742 8966 -6730
rect 9066 -754 9124 -742
rect 9066 -6730 9078 -754
rect 9112 -6730 9124 -754
rect 9066 -6742 9124 -6730
rect 9224 -754 9282 -742
rect 9224 -6730 9236 -754
rect 9270 -6730 9282 -754
rect 9224 -6742 9282 -6730
rect 9382 -754 9440 -742
rect 9382 -6730 9394 -754
rect 9428 -6730 9440 -754
rect 9382 -6742 9440 -6730
rect 9540 -754 9598 -742
rect 9540 -6730 9552 -754
rect 9586 -6730 9598 -754
rect 9540 -6742 9598 -6730
rect 9698 -754 9756 -742
rect 9698 -6730 9710 -754
rect 9744 -6730 9756 -754
rect 9698 -6742 9756 -6730
rect 9856 -754 9914 -742
rect 9856 -6730 9868 -754
rect 9902 -6730 9914 -754
rect 9856 -6742 9914 -6730
rect 10014 -754 10072 -742
rect 10014 -6730 10026 -754
rect 10060 -6730 10072 -754
rect 10014 -6742 10072 -6730
rect 10172 -754 10230 -742
rect 10172 -6730 10184 -754
rect 10218 -6730 10230 -754
rect 10172 -6742 10230 -6730
rect 10330 -754 10388 -742
rect 10330 -6730 10342 -754
rect 10376 -6730 10388 -754
rect 10330 -6742 10388 -6730
rect 10488 -754 10546 -742
rect 10488 -6730 10500 -754
rect 10534 -6730 10546 -754
rect 10488 -6742 10546 -6730
rect 10646 -754 10704 -742
rect 10646 -6730 10658 -754
rect 10692 -6730 10704 -754
rect 10646 -6742 10704 -6730
rect 10804 -754 10862 -742
rect 10804 -6730 10816 -754
rect 10850 -6730 10862 -754
rect 10804 -6742 10862 -6730
rect 10962 -754 11020 -742
rect 10962 -6730 10974 -754
rect 11008 -6730 11020 -754
rect 10962 -6742 11020 -6730
rect 11120 -754 11178 -742
rect 11120 -6730 11132 -754
rect 11166 -6730 11178 -754
rect 11120 -6742 11178 -6730
rect 11278 -754 11336 -742
rect 11278 -6730 11290 -754
rect 11324 -6730 11336 -754
rect 11278 -6742 11336 -6730
rect 11436 -754 11494 -742
rect 11436 -6730 11448 -754
rect 11482 -6730 11494 -754
rect 11436 -6742 11494 -6730
rect 11594 -754 11652 -742
rect 11594 -6730 11606 -754
rect 11640 -6730 11652 -754
rect 11594 -6742 11652 -6730
rect 11752 -754 11810 -742
rect 11752 -6730 11764 -754
rect 11798 -6730 11810 -754
rect 11752 -6742 11810 -6730
rect 11910 -754 11968 -742
rect 11910 -6730 11922 -754
rect 11956 -6730 11968 -754
rect 11910 -6742 11968 -6730
rect 14170 -754 14228 -742
rect 14170 -6730 14182 -754
rect 14216 -6730 14228 -754
rect 14170 -6742 14228 -6730
rect 14328 -754 14386 -742
rect 14328 -6730 14340 -754
rect 14374 -6730 14386 -754
rect 14328 -6742 14386 -6730
rect 14486 -754 14544 -742
rect 14486 -6730 14498 -754
rect 14532 -6730 14544 -754
rect 14486 -6742 14544 -6730
rect 14644 -754 14702 -742
rect 14644 -6730 14656 -754
rect 14690 -6730 14702 -754
rect 14644 -6742 14702 -6730
rect 14802 -754 14860 -742
rect 14802 -6730 14814 -754
rect 14848 -6730 14860 -754
rect 14802 -6742 14860 -6730
rect 14960 -754 15018 -742
rect 14960 -6730 14972 -754
rect 15006 -6730 15018 -754
rect 14960 -6742 15018 -6730
rect 15118 -754 15176 -742
rect 15118 -6730 15130 -754
rect 15164 -6730 15176 -754
rect 15118 -6742 15176 -6730
rect 15276 -754 15334 -742
rect 15276 -6730 15288 -754
rect 15322 -6730 15334 -754
rect 15276 -6742 15334 -6730
rect 15434 -754 15492 -742
rect 15434 -6730 15446 -754
rect 15480 -6730 15492 -754
rect 15434 -6742 15492 -6730
rect 15592 -754 15650 -742
rect 15592 -6730 15604 -754
rect 15638 -6730 15650 -754
rect 15592 -6742 15650 -6730
rect 15750 -754 15808 -742
rect 15750 -6730 15762 -754
rect 15796 -6730 15808 -754
rect 15750 -6742 15808 -6730
rect 15908 -754 15966 -742
rect 15908 -6730 15920 -754
rect 15954 -6730 15966 -754
rect 15908 -6742 15966 -6730
rect 16066 -754 16124 -742
rect 16066 -6730 16078 -754
rect 16112 -6730 16124 -754
rect 16066 -6742 16124 -6730
rect 16224 -754 16282 -742
rect 16224 -6730 16236 -754
rect 16270 -6730 16282 -754
rect 16224 -6742 16282 -6730
rect 16382 -754 16440 -742
rect 16382 -6730 16394 -754
rect 16428 -6730 16440 -754
rect 16382 -6742 16440 -6730
rect 16540 -754 16598 -742
rect 16540 -6730 16552 -754
rect 16586 -6730 16598 -754
rect 16540 -6742 16598 -6730
rect 16698 -754 16756 -742
rect 16698 -6730 16710 -754
rect 16744 -6730 16756 -754
rect 16698 -6742 16756 -6730
rect 16856 -754 16914 -742
rect 16856 -6730 16868 -754
rect 16902 -6730 16914 -754
rect 16856 -6742 16914 -6730
rect 17014 -754 17072 -742
rect 17014 -6730 17026 -754
rect 17060 -6730 17072 -754
rect 17014 -6742 17072 -6730
rect 17172 -754 17230 -742
rect 17172 -6730 17184 -754
rect 17218 -6730 17230 -754
rect 17172 -6742 17230 -6730
rect 17330 -754 17388 -742
rect 17330 -6730 17342 -754
rect 17376 -6730 17388 -754
rect 17330 -6742 17388 -6730
rect 17488 -754 17546 -742
rect 17488 -6730 17500 -754
rect 17534 -6730 17546 -754
rect 17488 -6742 17546 -6730
rect 17646 -754 17704 -742
rect 17646 -6730 17658 -754
rect 17692 -6730 17704 -754
rect 17646 -6742 17704 -6730
rect 17804 -754 17862 -742
rect 17804 -6730 17816 -754
rect 17850 -6730 17862 -754
rect 17804 -6742 17862 -6730
rect 17962 -754 18020 -742
rect 17962 -6730 17974 -754
rect 18008 -6730 18020 -754
rect 17962 -6742 18020 -6730
rect 18120 -754 18178 -742
rect 18120 -6730 18132 -754
rect 18166 -6730 18178 -754
rect 18120 -6742 18178 -6730
rect 18278 -754 18336 -742
rect 18278 -6730 18290 -754
rect 18324 -6730 18336 -754
rect 18278 -6742 18336 -6730
rect 18436 -754 18494 -742
rect 18436 -6730 18448 -754
rect 18482 -6730 18494 -754
rect 18436 -6742 18494 -6730
rect 18594 -754 18652 -742
rect 18594 -6730 18606 -754
rect 18640 -6730 18652 -754
rect 18594 -6742 18652 -6730
rect 18752 -754 18810 -742
rect 18752 -6730 18764 -754
rect 18798 -6730 18810 -754
rect 18752 -6742 18810 -6730
rect 18910 -754 18968 -742
rect 18910 -6730 18922 -754
rect 18956 -6730 18968 -754
rect 18910 -6742 18968 -6730
rect 21170 -754 21228 -742
rect 21170 -6730 21182 -754
rect 21216 -6730 21228 -754
rect 21170 -6742 21228 -6730
rect 21328 -754 21386 -742
rect 21328 -6730 21340 -754
rect 21374 -6730 21386 -754
rect 21328 -6742 21386 -6730
rect 21486 -754 21544 -742
rect 21486 -6730 21498 -754
rect 21532 -6730 21544 -754
rect 21486 -6742 21544 -6730
rect 21644 -754 21702 -742
rect 21644 -6730 21656 -754
rect 21690 -6730 21702 -754
rect 21644 -6742 21702 -6730
rect 21802 -754 21860 -742
rect 21802 -6730 21814 -754
rect 21848 -6730 21860 -754
rect 21802 -6742 21860 -6730
rect 21960 -754 22018 -742
rect 21960 -6730 21972 -754
rect 22006 -6730 22018 -754
rect 21960 -6742 22018 -6730
rect 22118 -754 22176 -742
rect 22118 -6730 22130 -754
rect 22164 -6730 22176 -754
rect 22118 -6742 22176 -6730
rect 22276 -754 22334 -742
rect 22276 -6730 22288 -754
rect 22322 -6730 22334 -754
rect 22276 -6742 22334 -6730
rect 22434 -754 22492 -742
rect 22434 -6730 22446 -754
rect 22480 -6730 22492 -754
rect 22434 -6742 22492 -6730
rect 22592 -754 22650 -742
rect 22592 -6730 22604 -754
rect 22638 -6730 22650 -754
rect 22592 -6742 22650 -6730
rect 22750 -754 22808 -742
rect 22750 -6730 22762 -754
rect 22796 -6730 22808 -754
rect 22750 -6742 22808 -6730
rect 22908 -754 22966 -742
rect 22908 -6730 22920 -754
rect 22954 -6730 22966 -754
rect 22908 -6742 22966 -6730
rect 23066 -754 23124 -742
rect 23066 -6730 23078 -754
rect 23112 -6730 23124 -754
rect 23066 -6742 23124 -6730
rect 23224 -754 23282 -742
rect 23224 -6730 23236 -754
rect 23270 -6730 23282 -754
rect 23224 -6742 23282 -6730
rect 23382 -754 23440 -742
rect 23382 -6730 23394 -754
rect 23428 -6730 23440 -754
rect 23382 -6742 23440 -6730
rect 23540 -754 23598 -742
rect 23540 -6730 23552 -754
rect 23586 -6730 23598 -754
rect 23540 -6742 23598 -6730
rect 23698 -754 23756 -742
rect 23698 -6730 23710 -754
rect 23744 -6730 23756 -754
rect 23698 -6742 23756 -6730
rect 23856 -754 23914 -742
rect 23856 -6730 23868 -754
rect 23902 -6730 23914 -754
rect 23856 -6742 23914 -6730
rect 24014 -754 24072 -742
rect 24014 -6730 24026 -754
rect 24060 -6730 24072 -754
rect 24014 -6742 24072 -6730
rect 24172 -754 24230 -742
rect 24172 -6730 24184 -754
rect 24218 -6730 24230 -754
rect 24172 -6742 24230 -6730
rect 24330 -754 24388 -742
rect 24330 -6730 24342 -754
rect 24376 -6730 24388 -754
rect 24330 -6742 24388 -6730
rect 24488 -754 24546 -742
rect 24488 -6730 24500 -754
rect 24534 -6730 24546 -754
rect 24488 -6742 24546 -6730
rect 24646 -754 24704 -742
rect 24646 -6730 24658 -754
rect 24692 -6730 24704 -754
rect 24646 -6742 24704 -6730
rect 24804 -754 24862 -742
rect 24804 -6730 24816 -754
rect 24850 -6730 24862 -754
rect 24804 -6742 24862 -6730
rect 24962 -754 25020 -742
rect 24962 -6730 24974 -754
rect 25008 -6730 25020 -754
rect 24962 -6742 25020 -6730
rect 25120 -754 25178 -742
rect 25120 -6730 25132 -754
rect 25166 -6730 25178 -754
rect 25120 -6742 25178 -6730
rect 25278 -754 25336 -742
rect 25278 -6730 25290 -754
rect 25324 -6730 25336 -754
rect 25278 -6742 25336 -6730
rect 25436 -754 25494 -742
rect 25436 -6730 25448 -754
rect 25482 -6730 25494 -754
rect 25436 -6742 25494 -6730
rect 25594 -754 25652 -742
rect 25594 -6730 25606 -754
rect 25640 -6730 25652 -754
rect 25594 -6742 25652 -6730
rect 25752 -754 25810 -742
rect 25752 -6730 25764 -754
rect 25798 -6730 25810 -754
rect 25752 -6742 25810 -6730
rect 25910 -754 25968 -742
rect 25910 -6730 25922 -754
rect 25956 -6730 25968 -754
rect 25910 -6742 25968 -6730
<< mvndiffc >>
rect 182 270 216 6246
rect 340 270 374 6246
rect 498 270 532 6246
rect 656 270 690 6246
rect 814 270 848 6246
rect 972 270 1006 6246
rect 1130 270 1164 6246
rect 1288 270 1322 6246
rect 1446 270 1480 6246
rect 1604 270 1638 6246
rect 1762 270 1796 6246
rect 1920 270 1954 6246
rect 2078 270 2112 6246
rect 2236 270 2270 6246
rect 2394 270 2428 6246
rect 2552 270 2586 6246
rect 2710 270 2744 6246
rect 2868 270 2902 6246
rect 3026 270 3060 6246
rect 3184 270 3218 6246
rect 3342 270 3376 6246
rect 3500 270 3534 6246
rect 3658 270 3692 6246
rect 3816 270 3850 6246
rect 3974 270 4008 6246
rect 4132 270 4166 6246
rect 4290 270 4324 6246
rect 4448 270 4482 6246
rect 4606 270 4640 6246
rect 4764 270 4798 6246
rect 4922 270 4956 6246
rect 7182 270 7216 6246
rect 7340 270 7374 6246
rect 7498 270 7532 6246
rect 7656 270 7690 6246
rect 7814 270 7848 6246
rect 7972 270 8006 6246
rect 8130 270 8164 6246
rect 8288 270 8322 6246
rect 8446 270 8480 6246
rect 8604 270 8638 6246
rect 8762 270 8796 6246
rect 8920 270 8954 6246
rect 9078 270 9112 6246
rect 9236 270 9270 6246
rect 9394 270 9428 6246
rect 9552 270 9586 6246
rect 9710 270 9744 6246
rect 9868 270 9902 6246
rect 10026 270 10060 6246
rect 10184 270 10218 6246
rect 10342 270 10376 6246
rect 10500 270 10534 6246
rect 10658 270 10692 6246
rect 10816 270 10850 6246
rect 10974 270 11008 6246
rect 11132 270 11166 6246
rect 11290 270 11324 6246
rect 11448 270 11482 6246
rect 11606 270 11640 6246
rect 11764 270 11798 6246
rect 11922 270 11956 6246
rect 14182 270 14216 6246
rect 14340 270 14374 6246
rect 14498 270 14532 6246
rect 14656 270 14690 6246
rect 14814 270 14848 6246
rect 14972 270 15006 6246
rect 15130 270 15164 6246
rect 15288 270 15322 6246
rect 15446 270 15480 6246
rect 15604 270 15638 6246
rect 15762 270 15796 6246
rect 15920 270 15954 6246
rect 16078 270 16112 6246
rect 16236 270 16270 6246
rect 16394 270 16428 6246
rect 16552 270 16586 6246
rect 16710 270 16744 6246
rect 16868 270 16902 6246
rect 17026 270 17060 6246
rect 17184 270 17218 6246
rect 17342 270 17376 6246
rect 17500 270 17534 6246
rect 17658 270 17692 6246
rect 17816 270 17850 6246
rect 17974 270 18008 6246
rect 18132 270 18166 6246
rect 18290 270 18324 6246
rect 18448 270 18482 6246
rect 18606 270 18640 6246
rect 18764 270 18798 6246
rect 18922 270 18956 6246
rect 21182 270 21216 6246
rect 21340 270 21374 6246
rect 21498 270 21532 6246
rect 21656 270 21690 6246
rect 21814 270 21848 6246
rect 21972 270 22006 6246
rect 22130 270 22164 6246
rect 22288 270 22322 6246
rect 22446 270 22480 6246
rect 22604 270 22638 6246
rect 22762 270 22796 6246
rect 22920 270 22954 6246
rect 23078 270 23112 6246
rect 23236 270 23270 6246
rect 23394 270 23428 6246
rect 23552 270 23586 6246
rect 23710 270 23744 6246
rect 23868 270 23902 6246
rect 24026 270 24060 6246
rect 24184 270 24218 6246
rect 24342 270 24376 6246
rect 24500 270 24534 6246
rect 24658 270 24692 6246
rect 24816 270 24850 6246
rect 24974 270 25008 6246
rect 25132 270 25166 6246
rect 25290 270 25324 6246
rect 25448 270 25482 6246
rect 25606 270 25640 6246
rect 25764 270 25798 6246
rect 25922 270 25956 6246
rect 182 -6730 216 -754
rect 340 -6730 374 -754
rect 498 -6730 532 -754
rect 656 -6730 690 -754
rect 814 -6730 848 -754
rect 972 -6730 1006 -754
rect 1130 -6730 1164 -754
rect 1288 -6730 1322 -754
rect 1446 -6730 1480 -754
rect 1604 -6730 1638 -754
rect 1762 -6730 1796 -754
rect 1920 -6730 1954 -754
rect 2078 -6730 2112 -754
rect 2236 -6730 2270 -754
rect 2394 -6730 2428 -754
rect 2552 -6730 2586 -754
rect 2710 -6730 2744 -754
rect 2868 -6730 2902 -754
rect 3026 -6730 3060 -754
rect 3184 -6730 3218 -754
rect 3342 -6730 3376 -754
rect 3500 -6730 3534 -754
rect 3658 -6730 3692 -754
rect 3816 -6730 3850 -754
rect 3974 -6730 4008 -754
rect 4132 -6730 4166 -754
rect 4290 -6730 4324 -754
rect 4448 -6730 4482 -754
rect 4606 -6730 4640 -754
rect 4764 -6730 4798 -754
rect 4922 -6730 4956 -754
rect 7182 -6730 7216 -754
rect 7340 -6730 7374 -754
rect 7498 -6730 7532 -754
rect 7656 -6730 7690 -754
rect 7814 -6730 7848 -754
rect 7972 -6730 8006 -754
rect 8130 -6730 8164 -754
rect 8288 -6730 8322 -754
rect 8446 -6730 8480 -754
rect 8604 -6730 8638 -754
rect 8762 -6730 8796 -754
rect 8920 -6730 8954 -754
rect 9078 -6730 9112 -754
rect 9236 -6730 9270 -754
rect 9394 -6730 9428 -754
rect 9552 -6730 9586 -754
rect 9710 -6730 9744 -754
rect 9868 -6730 9902 -754
rect 10026 -6730 10060 -754
rect 10184 -6730 10218 -754
rect 10342 -6730 10376 -754
rect 10500 -6730 10534 -754
rect 10658 -6730 10692 -754
rect 10816 -6730 10850 -754
rect 10974 -6730 11008 -754
rect 11132 -6730 11166 -754
rect 11290 -6730 11324 -754
rect 11448 -6730 11482 -754
rect 11606 -6730 11640 -754
rect 11764 -6730 11798 -754
rect 11922 -6730 11956 -754
rect 14182 -6730 14216 -754
rect 14340 -6730 14374 -754
rect 14498 -6730 14532 -754
rect 14656 -6730 14690 -754
rect 14814 -6730 14848 -754
rect 14972 -6730 15006 -754
rect 15130 -6730 15164 -754
rect 15288 -6730 15322 -754
rect 15446 -6730 15480 -754
rect 15604 -6730 15638 -754
rect 15762 -6730 15796 -754
rect 15920 -6730 15954 -754
rect 16078 -6730 16112 -754
rect 16236 -6730 16270 -754
rect 16394 -6730 16428 -754
rect 16552 -6730 16586 -754
rect 16710 -6730 16744 -754
rect 16868 -6730 16902 -754
rect 17026 -6730 17060 -754
rect 17184 -6730 17218 -754
rect 17342 -6730 17376 -754
rect 17500 -6730 17534 -754
rect 17658 -6730 17692 -754
rect 17816 -6730 17850 -754
rect 17974 -6730 18008 -754
rect 18132 -6730 18166 -754
rect 18290 -6730 18324 -754
rect 18448 -6730 18482 -754
rect 18606 -6730 18640 -754
rect 18764 -6730 18798 -754
rect 18922 -6730 18956 -754
rect 21182 -6730 21216 -754
rect 21340 -6730 21374 -754
rect 21498 -6730 21532 -754
rect 21656 -6730 21690 -754
rect 21814 -6730 21848 -754
rect 21972 -6730 22006 -754
rect 22130 -6730 22164 -754
rect 22288 -6730 22322 -754
rect 22446 -6730 22480 -754
rect 22604 -6730 22638 -754
rect 22762 -6730 22796 -754
rect 22920 -6730 22954 -754
rect 23078 -6730 23112 -754
rect 23236 -6730 23270 -754
rect 23394 -6730 23428 -754
rect 23552 -6730 23586 -754
rect 23710 -6730 23744 -754
rect 23868 -6730 23902 -754
rect 24026 -6730 24060 -754
rect 24184 -6730 24218 -754
rect 24342 -6730 24376 -754
rect 24500 -6730 24534 -754
rect 24658 -6730 24692 -754
rect 24816 -6730 24850 -754
rect 24974 -6730 25008 -754
rect 25132 -6730 25166 -754
rect 25290 -6730 25324 -754
rect 25448 -6730 25482 -754
rect 25606 -6730 25640 -754
rect 25764 -6730 25798 -754
rect 25922 -6730 25956 -754
<< mvpsubdiff >>
rect 36 6468 5102 6480
rect 36 6434 144 6468
rect 4994 6434 5102 6468
rect 36 6422 5102 6434
rect 36 6372 94 6422
rect 36 144 48 6372
rect 82 144 94 6372
rect 5044 6372 5102 6422
rect 36 94 94 144
rect 5044 144 5056 6372
rect 5090 144 5102 6372
rect 5044 94 5102 144
rect 36 82 5102 94
rect 36 48 144 82
rect 4994 48 5102 82
rect 36 36 5102 48
rect 7036 6468 12102 6480
rect 7036 6434 7144 6468
rect 11994 6434 12102 6468
rect 7036 6422 12102 6434
rect 7036 6372 7094 6422
rect 7036 144 7048 6372
rect 7082 144 7094 6372
rect 12044 6372 12102 6422
rect 7036 94 7094 144
rect 12044 144 12056 6372
rect 12090 144 12102 6372
rect 12044 94 12102 144
rect 7036 82 12102 94
rect 7036 48 7144 82
rect 11994 48 12102 82
rect 7036 36 12102 48
rect 14036 6468 19102 6480
rect 14036 6434 14144 6468
rect 18994 6434 19102 6468
rect 14036 6422 19102 6434
rect 14036 6372 14094 6422
rect 14036 144 14048 6372
rect 14082 144 14094 6372
rect 19044 6372 19102 6422
rect 14036 94 14094 144
rect 19044 144 19056 6372
rect 19090 144 19102 6372
rect 19044 94 19102 144
rect 14036 82 19102 94
rect 14036 48 14144 82
rect 18994 48 19102 82
rect 14036 36 19102 48
rect 21036 6468 26102 6480
rect 21036 6434 21144 6468
rect 25994 6434 26102 6468
rect 21036 6422 26102 6434
rect 21036 6372 21094 6422
rect 21036 144 21048 6372
rect 21082 144 21094 6372
rect 26044 6372 26102 6422
rect 21036 94 21094 144
rect 26044 144 26056 6372
rect 26090 144 26102 6372
rect 26044 94 26102 144
rect 21036 82 26102 94
rect 21036 48 21144 82
rect 25994 48 26102 82
rect 21036 36 26102 48
rect 36 -532 5102 -520
rect 36 -566 144 -532
rect 4994 -566 5102 -532
rect 36 -578 5102 -566
rect 36 -628 94 -578
rect 36 -6856 48 -628
rect 82 -6856 94 -628
rect 5044 -628 5102 -578
rect 36 -6906 94 -6856
rect 5044 -6856 5056 -628
rect 5090 -6856 5102 -628
rect 5044 -6906 5102 -6856
rect 36 -6918 5102 -6906
rect 36 -6952 144 -6918
rect 4994 -6952 5102 -6918
rect 36 -6964 5102 -6952
rect 7036 -532 12102 -520
rect 7036 -566 7144 -532
rect 11994 -566 12102 -532
rect 7036 -578 12102 -566
rect 7036 -628 7094 -578
rect 7036 -6856 7048 -628
rect 7082 -6856 7094 -628
rect 12044 -628 12102 -578
rect 7036 -6906 7094 -6856
rect 12044 -6856 12056 -628
rect 12090 -6856 12102 -628
rect 12044 -6906 12102 -6856
rect 7036 -6918 12102 -6906
rect 7036 -6952 7144 -6918
rect 11994 -6952 12102 -6918
rect 7036 -6964 12102 -6952
rect 14036 -532 19102 -520
rect 14036 -566 14144 -532
rect 18994 -566 19102 -532
rect 14036 -578 19102 -566
rect 14036 -628 14094 -578
rect 14036 -6856 14048 -628
rect 14082 -6856 14094 -628
rect 19044 -628 19102 -578
rect 14036 -6906 14094 -6856
rect 19044 -6856 19056 -628
rect 19090 -6856 19102 -628
rect 19044 -6906 19102 -6856
rect 14036 -6918 19102 -6906
rect 14036 -6952 14144 -6918
rect 18994 -6952 19102 -6918
rect 14036 -6964 19102 -6952
rect 21036 -532 26102 -520
rect 21036 -566 21144 -532
rect 25994 -566 26102 -532
rect 21036 -578 26102 -566
rect 21036 -628 21094 -578
rect 21036 -6856 21048 -628
rect 21082 -6856 21094 -628
rect 26044 -628 26102 -578
rect 21036 -6906 21094 -6856
rect 26044 -6856 26056 -628
rect 26090 -6856 26102 -628
rect 26044 -6906 26102 -6856
rect 21036 -6918 26102 -6906
rect 21036 -6952 21144 -6918
rect 25994 -6952 26102 -6918
rect 21036 -6964 26102 -6952
<< mvpsubdiffcont >>
rect 144 6434 4994 6468
rect 48 144 82 6372
rect 5056 144 5090 6372
rect 144 48 4994 82
rect 7144 6434 11994 6468
rect 7048 144 7082 6372
rect 12056 144 12090 6372
rect 7144 48 11994 82
rect 14144 6434 18994 6468
rect 14048 144 14082 6372
rect 19056 144 19090 6372
rect 14144 48 18994 82
rect 21144 6434 25994 6468
rect 21048 144 21082 6372
rect 26056 144 26090 6372
rect 21144 48 25994 82
rect 144 -566 4994 -532
rect 48 -6856 82 -628
rect 5056 -6856 5090 -628
rect 144 -6952 4994 -6918
rect 7144 -566 11994 -532
rect 7048 -6856 7082 -628
rect 12056 -6856 12090 -628
rect 7144 -6952 11994 -6918
rect 14144 -566 18994 -532
rect 14048 -6856 14082 -628
rect 19056 -6856 19090 -628
rect 14144 -6952 18994 -6918
rect 21144 -566 25994 -532
rect 21048 -6856 21082 -628
rect 26056 -6856 26090 -628
rect 21144 -6952 25994 -6918
<< poly >>
rect 228 6330 328 6346
rect 228 6296 244 6330
rect 312 6296 328 6330
rect 228 6258 328 6296
rect 386 6330 486 6346
rect 386 6296 402 6330
rect 470 6296 486 6330
rect 386 6258 486 6296
rect 544 6330 644 6346
rect 544 6296 560 6330
rect 628 6296 644 6330
rect 544 6258 644 6296
rect 702 6330 802 6346
rect 702 6296 718 6330
rect 786 6296 802 6330
rect 702 6258 802 6296
rect 860 6330 960 6346
rect 860 6296 876 6330
rect 944 6296 960 6330
rect 860 6258 960 6296
rect 1018 6330 1118 6346
rect 1018 6296 1034 6330
rect 1102 6296 1118 6330
rect 1018 6258 1118 6296
rect 1176 6330 1276 6346
rect 1176 6296 1192 6330
rect 1260 6296 1276 6330
rect 1176 6258 1276 6296
rect 1334 6330 1434 6346
rect 1334 6296 1350 6330
rect 1418 6296 1434 6330
rect 1334 6258 1434 6296
rect 1492 6330 1592 6346
rect 1492 6296 1508 6330
rect 1576 6296 1592 6330
rect 1492 6258 1592 6296
rect 1650 6330 1750 6346
rect 1650 6296 1666 6330
rect 1734 6296 1750 6330
rect 1650 6258 1750 6296
rect 1808 6330 1908 6346
rect 1808 6296 1824 6330
rect 1892 6296 1908 6330
rect 1808 6258 1908 6296
rect 1966 6330 2066 6346
rect 1966 6296 1982 6330
rect 2050 6296 2066 6330
rect 1966 6258 2066 6296
rect 2124 6330 2224 6346
rect 2124 6296 2140 6330
rect 2208 6296 2224 6330
rect 2124 6258 2224 6296
rect 2282 6330 2382 6346
rect 2282 6296 2298 6330
rect 2366 6296 2382 6330
rect 2282 6258 2382 6296
rect 2440 6330 2540 6346
rect 2440 6296 2456 6330
rect 2524 6296 2540 6330
rect 2440 6258 2540 6296
rect 2598 6330 2698 6346
rect 2598 6296 2614 6330
rect 2682 6296 2698 6330
rect 2598 6258 2698 6296
rect 2756 6330 2856 6346
rect 2756 6296 2772 6330
rect 2840 6296 2856 6330
rect 2756 6258 2856 6296
rect 2914 6330 3014 6346
rect 2914 6296 2930 6330
rect 2998 6296 3014 6330
rect 2914 6258 3014 6296
rect 3072 6330 3172 6346
rect 3072 6296 3088 6330
rect 3156 6296 3172 6330
rect 3072 6258 3172 6296
rect 3230 6330 3330 6346
rect 3230 6296 3246 6330
rect 3314 6296 3330 6330
rect 3230 6258 3330 6296
rect 3388 6330 3488 6346
rect 3388 6296 3404 6330
rect 3472 6296 3488 6330
rect 3388 6258 3488 6296
rect 3546 6330 3646 6346
rect 3546 6296 3562 6330
rect 3630 6296 3646 6330
rect 3546 6258 3646 6296
rect 3704 6330 3804 6346
rect 3704 6296 3720 6330
rect 3788 6296 3804 6330
rect 3704 6258 3804 6296
rect 3862 6330 3962 6346
rect 3862 6296 3878 6330
rect 3946 6296 3962 6330
rect 3862 6258 3962 6296
rect 4020 6330 4120 6346
rect 4020 6296 4036 6330
rect 4104 6296 4120 6330
rect 4020 6258 4120 6296
rect 4178 6330 4278 6346
rect 4178 6296 4194 6330
rect 4262 6296 4278 6330
rect 4178 6258 4278 6296
rect 4336 6330 4436 6346
rect 4336 6296 4352 6330
rect 4420 6296 4436 6330
rect 4336 6258 4436 6296
rect 4494 6330 4594 6346
rect 4494 6296 4510 6330
rect 4578 6296 4594 6330
rect 4494 6258 4594 6296
rect 4652 6330 4752 6346
rect 4652 6296 4668 6330
rect 4736 6296 4752 6330
rect 4652 6258 4752 6296
rect 4810 6330 4910 6346
rect 4810 6296 4826 6330
rect 4894 6296 4910 6330
rect 4810 6258 4910 6296
rect 228 220 328 258
rect 228 186 244 220
rect 312 186 328 220
rect 228 170 328 186
rect 386 220 486 258
rect 386 186 402 220
rect 470 186 486 220
rect 386 170 486 186
rect 544 220 644 258
rect 544 186 560 220
rect 628 186 644 220
rect 544 170 644 186
rect 702 220 802 258
rect 702 186 718 220
rect 786 186 802 220
rect 702 170 802 186
rect 860 220 960 258
rect 860 186 876 220
rect 944 186 960 220
rect 860 170 960 186
rect 1018 220 1118 258
rect 1018 186 1034 220
rect 1102 186 1118 220
rect 1018 170 1118 186
rect 1176 220 1276 258
rect 1176 186 1192 220
rect 1260 186 1276 220
rect 1176 170 1276 186
rect 1334 220 1434 258
rect 1334 186 1350 220
rect 1418 186 1434 220
rect 1334 170 1434 186
rect 1492 220 1592 258
rect 1492 186 1508 220
rect 1576 186 1592 220
rect 1492 170 1592 186
rect 1650 220 1750 258
rect 1650 186 1666 220
rect 1734 186 1750 220
rect 1650 170 1750 186
rect 1808 220 1908 258
rect 1808 186 1824 220
rect 1892 186 1908 220
rect 1808 170 1908 186
rect 1966 220 2066 258
rect 1966 186 1982 220
rect 2050 186 2066 220
rect 1966 170 2066 186
rect 2124 220 2224 258
rect 2124 186 2140 220
rect 2208 186 2224 220
rect 2124 170 2224 186
rect 2282 220 2382 258
rect 2282 186 2298 220
rect 2366 186 2382 220
rect 2282 170 2382 186
rect 2440 220 2540 258
rect 2440 186 2456 220
rect 2524 186 2540 220
rect 2440 170 2540 186
rect 2598 220 2698 258
rect 2598 186 2614 220
rect 2682 186 2698 220
rect 2598 170 2698 186
rect 2756 220 2856 258
rect 2756 186 2772 220
rect 2840 186 2856 220
rect 2756 170 2856 186
rect 2914 220 3014 258
rect 2914 186 2930 220
rect 2998 186 3014 220
rect 2914 170 3014 186
rect 3072 220 3172 258
rect 3072 186 3088 220
rect 3156 186 3172 220
rect 3072 170 3172 186
rect 3230 220 3330 258
rect 3230 186 3246 220
rect 3314 186 3330 220
rect 3230 170 3330 186
rect 3388 220 3488 258
rect 3388 186 3404 220
rect 3472 186 3488 220
rect 3388 170 3488 186
rect 3546 220 3646 258
rect 3546 186 3562 220
rect 3630 186 3646 220
rect 3546 170 3646 186
rect 3704 220 3804 258
rect 3704 186 3720 220
rect 3788 186 3804 220
rect 3704 170 3804 186
rect 3862 220 3962 258
rect 3862 186 3878 220
rect 3946 186 3962 220
rect 3862 170 3962 186
rect 4020 220 4120 258
rect 4020 186 4036 220
rect 4104 186 4120 220
rect 4020 170 4120 186
rect 4178 220 4278 258
rect 4178 186 4194 220
rect 4262 186 4278 220
rect 4178 170 4278 186
rect 4336 220 4436 258
rect 4336 186 4352 220
rect 4420 186 4436 220
rect 4336 170 4436 186
rect 4494 220 4594 258
rect 4494 186 4510 220
rect 4578 186 4594 220
rect 4494 170 4594 186
rect 4652 220 4752 258
rect 4652 186 4668 220
rect 4736 186 4752 220
rect 4652 170 4752 186
rect 4810 220 4910 258
rect 4810 186 4826 220
rect 4894 186 4910 220
rect 4810 170 4910 186
rect 7228 6330 7328 6346
rect 7228 6296 7244 6330
rect 7312 6296 7328 6330
rect 7228 6258 7328 6296
rect 7386 6330 7486 6346
rect 7386 6296 7402 6330
rect 7470 6296 7486 6330
rect 7386 6258 7486 6296
rect 7544 6330 7644 6346
rect 7544 6296 7560 6330
rect 7628 6296 7644 6330
rect 7544 6258 7644 6296
rect 7702 6330 7802 6346
rect 7702 6296 7718 6330
rect 7786 6296 7802 6330
rect 7702 6258 7802 6296
rect 7860 6330 7960 6346
rect 7860 6296 7876 6330
rect 7944 6296 7960 6330
rect 7860 6258 7960 6296
rect 8018 6330 8118 6346
rect 8018 6296 8034 6330
rect 8102 6296 8118 6330
rect 8018 6258 8118 6296
rect 8176 6330 8276 6346
rect 8176 6296 8192 6330
rect 8260 6296 8276 6330
rect 8176 6258 8276 6296
rect 8334 6330 8434 6346
rect 8334 6296 8350 6330
rect 8418 6296 8434 6330
rect 8334 6258 8434 6296
rect 8492 6330 8592 6346
rect 8492 6296 8508 6330
rect 8576 6296 8592 6330
rect 8492 6258 8592 6296
rect 8650 6330 8750 6346
rect 8650 6296 8666 6330
rect 8734 6296 8750 6330
rect 8650 6258 8750 6296
rect 8808 6330 8908 6346
rect 8808 6296 8824 6330
rect 8892 6296 8908 6330
rect 8808 6258 8908 6296
rect 8966 6330 9066 6346
rect 8966 6296 8982 6330
rect 9050 6296 9066 6330
rect 8966 6258 9066 6296
rect 9124 6330 9224 6346
rect 9124 6296 9140 6330
rect 9208 6296 9224 6330
rect 9124 6258 9224 6296
rect 9282 6330 9382 6346
rect 9282 6296 9298 6330
rect 9366 6296 9382 6330
rect 9282 6258 9382 6296
rect 9440 6330 9540 6346
rect 9440 6296 9456 6330
rect 9524 6296 9540 6330
rect 9440 6258 9540 6296
rect 9598 6330 9698 6346
rect 9598 6296 9614 6330
rect 9682 6296 9698 6330
rect 9598 6258 9698 6296
rect 9756 6330 9856 6346
rect 9756 6296 9772 6330
rect 9840 6296 9856 6330
rect 9756 6258 9856 6296
rect 9914 6330 10014 6346
rect 9914 6296 9930 6330
rect 9998 6296 10014 6330
rect 9914 6258 10014 6296
rect 10072 6330 10172 6346
rect 10072 6296 10088 6330
rect 10156 6296 10172 6330
rect 10072 6258 10172 6296
rect 10230 6330 10330 6346
rect 10230 6296 10246 6330
rect 10314 6296 10330 6330
rect 10230 6258 10330 6296
rect 10388 6330 10488 6346
rect 10388 6296 10404 6330
rect 10472 6296 10488 6330
rect 10388 6258 10488 6296
rect 10546 6330 10646 6346
rect 10546 6296 10562 6330
rect 10630 6296 10646 6330
rect 10546 6258 10646 6296
rect 10704 6330 10804 6346
rect 10704 6296 10720 6330
rect 10788 6296 10804 6330
rect 10704 6258 10804 6296
rect 10862 6330 10962 6346
rect 10862 6296 10878 6330
rect 10946 6296 10962 6330
rect 10862 6258 10962 6296
rect 11020 6330 11120 6346
rect 11020 6296 11036 6330
rect 11104 6296 11120 6330
rect 11020 6258 11120 6296
rect 11178 6330 11278 6346
rect 11178 6296 11194 6330
rect 11262 6296 11278 6330
rect 11178 6258 11278 6296
rect 11336 6330 11436 6346
rect 11336 6296 11352 6330
rect 11420 6296 11436 6330
rect 11336 6258 11436 6296
rect 11494 6330 11594 6346
rect 11494 6296 11510 6330
rect 11578 6296 11594 6330
rect 11494 6258 11594 6296
rect 11652 6330 11752 6346
rect 11652 6296 11668 6330
rect 11736 6296 11752 6330
rect 11652 6258 11752 6296
rect 11810 6330 11910 6346
rect 11810 6296 11826 6330
rect 11894 6296 11910 6330
rect 11810 6258 11910 6296
rect 7228 220 7328 258
rect 7228 186 7244 220
rect 7312 186 7328 220
rect 7228 170 7328 186
rect 7386 220 7486 258
rect 7386 186 7402 220
rect 7470 186 7486 220
rect 7386 170 7486 186
rect 7544 220 7644 258
rect 7544 186 7560 220
rect 7628 186 7644 220
rect 7544 170 7644 186
rect 7702 220 7802 258
rect 7702 186 7718 220
rect 7786 186 7802 220
rect 7702 170 7802 186
rect 7860 220 7960 258
rect 7860 186 7876 220
rect 7944 186 7960 220
rect 7860 170 7960 186
rect 8018 220 8118 258
rect 8018 186 8034 220
rect 8102 186 8118 220
rect 8018 170 8118 186
rect 8176 220 8276 258
rect 8176 186 8192 220
rect 8260 186 8276 220
rect 8176 170 8276 186
rect 8334 220 8434 258
rect 8334 186 8350 220
rect 8418 186 8434 220
rect 8334 170 8434 186
rect 8492 220 8592 258
rect 8492 186 8508 220
rect 8576 186 8592 220
rect 8492 170 8592 186
rect 8650 220 8750 258
rect 8650 186 8666 220
rect 8734 186 8750 220
rect 8650 170 8750 186
rect 8808 220 8908 258
rect 8808 186 8824 220
rect 8892 186 8908 220
rect 8808 170 8908 186
rect 8966 220 9066 258
rect 8966 186 8982 220
rect 9050 186 9066 220
rect 8966 170 9066 186
rect 9124 220 9224 258
rect 9124 186 9140 220
rect 9208 186 9224 220
rect 9124 170 9224 186
rect 9282 220 9382 258
rect 9282 186 9298 220
rect 9366 186 9382 220
rect 9282 170 9382 186
rect 9440 220 9540 258
rect 9440 186 9456 220
rect 9524 186 9540 220
rect 9440 170 9540 186
rect 9598 220 9698 258
rect 9598 186 9614 220
rect 9682 186 9698 220
rect 9598 170 9698 186
rect 9756 220 9856 258
rect 9756 186 9772 220
rect 9840 186 9856 220
rect 9756 170 9856 186
rect 9914 220 10014 258
rect 9914 186 9930 220
rect 9998 186 10014 220
rect 9914 170 10014 186
rect 10072 220 10172 258
rect 10072 186 10088 220
rect 10156 186 10172 220
rect 10072 170 10172 186
rect 10230 220 10330 258
rect 10230 186 10246 220
rect 10314 186 10330 220
rect 10230 170 10330 186
rect 10388 220 10488 258
rect 10388 186 10404 220
rect 10472 186 10488 220
rect 10388 170 10488 186
rect 10546 220 10646 258
rect 10546 186 10562 220
rect 10630 186 10646 220
rect 10546 170 10646 186
rect 10704 220 10804 258
rect 10704 186 10720 220
rect 10788 186 10804 220
rect 10704 170 10804 186
rect 10862 220 10962 258
rect 10862 186 10878 220
rect 10946 186 10962 220
rect 10862 170 10962 186
rect 11020 220 11120 258
rect 11020 186 11036 220
rect 11104 186 11120 220
rect 11020 170 11120 186
rect 11178 220 11278 258
rect 11178 186 11194 220
rect 11262 186 11278 220
rect 11178 170 11278 186
rect 11336 220 11436 258
rect 11336 186 11352 220
rect 11420 186 11436 220
rect 11336 170 11436 186
rect 11494 220 11594 258
rect 11494 186 11510 220
rect 11578 186 11594 220
rect 11494 170 11594 186
rect 11652 220 11752 258
rect 11652 186 11668 220
rect 11736 186 11752 220
rect 11652 170 11752 186
rect 11810 220 11910 258
rect 11810 186 11826 220
rect 11894 186 11910 220
rect 11810 170 11910 186
rect 14228 6330 14328 6346
rect 14228 6296 14244 6330
rect 14312 6296 14328 6330
rect 14228 6258 14328 6296
rect 14386 6330 14486 6346
rect 14386 6296 14402 6330
rect 14470 6296 14486 6330
rect 14386 6258 14486 6296
rect 14544 6330 14644 6346
rect 14544 6296 14560 6330
rect 14628 6296 14644 6330
rect 14544 6258 14644 6296
rect 14702 6330 14802 6346
rect 14702 6296 14718 6330
rect 14786 6296 14802 6330
rect 14702 6258 14802 6296
rect 14860 6330 14960 6346
rect 14860 6296 14876 6330
rect 14944 6296 14960 6330
rect 14860 6258 14960 6296
rect 15018 6330 15118 6346
rect 15018 6296 15034 6330
rect 15102 6296 15118 6330
rect 15018 6258 15118 6296
rect 15176 6330 15276 6346
rect 15176 6296 15192 6330
rect 15260 6296 15276 6330
rect 15176 6258 15276 6296
rect 15334 6330 15434 6346
rect 15334 6296 15350 6330
rect 15418 6296 15434 6330
rect 15334 6258 15434 6296
rect 15492 6330 15592 6346
rect 15492 6296 15508 6330
rect 15576 6296 15592 6330
rect 15492 6258 15592 6296
rect 15650 6330 15750 6346
rect 15650 6296 15666 6330
rect 15734 6296 15750 6330
rect 15650 6258 15750 6296
rect 15808 6330 15908 6346
rect 15808 6296 15824 6330
rect 15892 6296 15908 6330
rect 15808 6258 15908 6296
rect 15966 6330 16066 6346
rect 15966 6296 15982 6330
rect 16050 6296 16066 6330
rect 15966 6258 16066 6296
rect 16124 6330 16224 6346
rect 16124 6296 16140 6330
rect 16208 6296 16224 6330
rect 16124 6258 16224 6296
rect 16282 6330 16382 6346
rect 16282 6296 16298 6330
rect 16366 6296 16382 6330
rect 16282 6258 16382 6296
rect 16440 6330 16540 6346
rect 16440 6296 16456 6330
rect 16524 6296 16540 6330
rect 16440 6258 16540 6296
rect 16598 6330 16698 6346
rect 16598 6296 16614 6330
rect 16682 6296 16698 6330
rect 16598 6258 16698 6296
rect 16756 6330 16856 6346
rect 16756 6296 16772 6330
rect 16840 6296 16856 6330
rect 16756 6258 16856 6296
rect 16914 6330 17014 6346
rect 16914 6296 16930 6330
rect 16998 6296 17014 6330
rect 16914 6258 17014 6296
rect 17072 6330 17172 6346
rect 17072 6296 17088 6330
rect 17156 6296 17172 6330
rect 17072 6258 17172 6296
rect 17230 6330 17330 6346
rect 17230 6296 17246 6330
rect 17314 6296 17330 6330
rect 17230 6258 17330 6296
rect 17388 6330 17488 6346
rect 17388 6296 17404 6330
rect 17472 6296 17488 6330
rect 17388 6258 17488 6296
rect 17546 6330 17646 6346
rect 17546 6296 17562 6330
rect 17630 6296 17646 6330
rect 17546 6258 17646 6296
rect 17704 6330 17804 6346
rect 17704 6296 17720 6330
rect 17788 6296 17804 6330
rect 17704 6258 17804 6296
rect 17862 6330 17962 6346
rect 17862 6296 17878 6330
rect 17946 6296 17962 6330
rect 17862 6258 17962 6296
rect 18020 6330 18120 6346
rect 18020 6296 18036 6330
rect 18104 6296 18120 6330
rect 18020 6258 18120 6296
rect 18178 6330 18278 6346
rect 18178 6296 18194 6330
rect 18262 6296 18278 6330
rect 18178 6258 18278 6296
rect 18336 6330 18436 6346
rect 18336 6296 18352 6330
rect 18420 6296 18436 6330
rect 18336 6258 18436 6296
rect 18494 6330 18594 6346
rect 18494 6296 18510 6330
rect 18578 6296 18594 6330
rect 18494 6258 18594 6296
rect 18652 6330 18752 6346
rect 18652 6296 18668 6330
rect 18736 6296 18752 6330
rect 18652 6258 18752 6296
rect 18810 6330 18910 6346
rect 18810 6296 18826 6330
rect 18894 6296 18910 6330
rect 18810 6258 18910 6296
rect 14228 220 14328 258
rect 14228 186 14244 220
rect 14312 186 14328 220
rect 14228 170 14328 186
rect 14386 220 14486 258
rect 14386 186 14402 220
rect 14470 186 14486 220
rect 14386 170 14486 186
rect 14544 220 14644 258
rect 14544 186 14560 220
rect 14628 186 14644 220
rect 14544 170 14644 186
rect 14702 220 14802 258
rect 14702 186 14718 220
rect 14786 186 14802 220
rect 14702 170 14802 186
rect 14860 220 14960 258
rect 14860 186 14876 220
rect 14944 186 14960 220
rect 14860 170 14960 186
rect 15018 220 15118 258
rect 15018 186 15034 220
rect 15102 186 15118 220
rect 15018 170 15118 186
rect 15176 220 15276 258
rect 15176 186 15192 220
rect 15260 186 15276 220
rect 15176 170 15276 186
rect 15334 220 15434 258
rect 15334 186 15350 220
rect 15418 186 15434 220
rect 15334 170 15434 186
rect 15492 220 15592 258
rect 15492 186 15508 220
rect 15576 186 15592 220
rect 15492 170 15592 186
rect 15650 220 15750 258
rect 15650 186 15666 220
rect 15734 186 15750 220
rect 15650 170 15750 186
rect 15808 220 15908 258
rect 15808 186 15824 220
rect 15892 186 15908 220
rect 15808 170 15908 186
rect 15966 220 16066 258
rect 15966 186 15982 220
rect 16050 186 16066 220
rect 15966 170 16066 186
rect 16124 220 16224 258
rect 16124 186 16140 220
rect 16208 186 16224 220
rect 16124 170 16224 186
rect 16282 220 16382 258
rect 16282 186 16298 220
rect 16366 186 16382 220
rect 16282 170 16382 186
rect 16440 220 16540 258
rect 16440 186 16456 220
rect 16524 186 16540 220
rect 16440 170 16540 186
rect 16598 220 16698 258
rect 16598 186 16614 220
rect 16682 186 16698 220
rect 16598 170 16698 186
rect 16756 220 16856 258
rect 16756 186 16772 220
rect 16840 186 16856 220
rect 16756 170 16856 186
rect 16914 220 17014 258
rect 16914 186 16930 220
rect 16998 186 17014 220
rect 16914 170 17014 186
rect 17072 220 17172 258
rect 17072 186 17088 220
rect 17156 186 17172 220
rect 17072 170 17172 186
rect 17230 220 17330 258
rect 17230 186 17246 220
rect 17314 186 17330 220
rect 17230 170 17330 186
rect 17388 220 17488 258
rect 17388 186 17404 220
rect 17472 186 17488 220
rect 17388 170 17488 186
rect 17546 220 17646 258
rect 17546 186 17562 220
rect 17630 186 17646 220
rect 17546 170 17646 186
rect 17704 220 17804 258
rect 17704 186 17720 220
rect 17788 186 17804 220
rect 17704 170 17804 186
rect 17862 220 17962 258
rect 17862 186 17878 220
rect 17946 186 17962 220
rect 17862 170 17962 186
rect 18020 220 18120 258
rect 18020 186 18036 220
rect 18104 186 18120 220
rect 18020 170 18120 186
rect 18178 220 18278 258
rect 18178 186 18194 220
rect 18262 186 18278 220
rect 18178 170 18278 186
rect 18336 220 18436 258
rect 18336 186 18352 220
rect 18420 186 18436 220
rect 18336 170 18436 186
rect 18494 220 18594 258
rect 18494 186 18510 220
rect 18578 186 18594 220
rect 18494 170 18594 186
rect 18652 220 18752 258
rect 18652 186 18668 220
rect 18736 186 18752 220
rect 18652 170 18752 186
rect 18810 220 18910 258
rect 18810 186 18826 220
rect 18894 186 18910 220
rect 18810 170 18910 186
rect 21228 6330 21328 6346
rect 21228 6296 21244 6330
rect 21312 6296 21328 6330
rect 21228 6258 21328 6296
rect 21386 6330 21486 6346
rect 21386 6296 21402 6330
rect 21470 6296 21486 6330
rect 21386 6258 21486 6296
rect 21544 6330 21644 6346
rect 21544 6296 21560 6330
rect 21628 6296 21644 6330
rect 21544 6258 21644 6296
rect 21702 6330 21802 6346
rect 21702 6296 21718 6330
rect 21786 6296 21802 6330
rect 21702 6258 21802 6296
rect 21860 6330 21960 6346
rect 21860 6296 21876 6330
rect 21944 6296 21960 6330
rect 21860 6258 21960 6296
rect 22018 6330 22118 6346
rect 22018 6296 22034 6330
rect 22102 6296 22118 6330
rect 22018 6258 22118 6296
rect 22176 6330 22276 6346
rect 22176 6296 22192 6330
rect 22260 6296 22276 6330
rect 22176 6258 22276 6296
rect 22334 6330 22434 6346
rect 22334 6296 22350 6330
rect 22418 6296 22434 6330
rect 22334 6258 22434 6296
rect 22492 6330 22592 6346
rect 22492 6296 22508 6330
rect 22576 6296 22592 6330
rect 22492 6258 22592 6296
rect 22650 6330 22750 6346
rect 22650 6296 22666 6330
rect 22734 6296 22750 6330
rect 22650 6258 22750 6296
rect 22808 6330 22908 6346
rect 22808 6296 22824 6330
rect 22892 6296 22908 6330
rect 22808 6258 22908 6296
rect 22966 6330 23066 6346
rect 22966 6296 22982 6330
rect 23050 6296 23066 6330
rect 22966 6258 23066 6296
rect 23124 6330 23224 6346
rect 23124 6296 23140 6330
rect 23208 6296 23224 6330
rect 23124 6258 23224 6296
rect 23282 6330 23382 6346
rect 23282 6296 23298 6330
rect 23366 6296 23382 6330
rect 23282 6258 23382 6296
rect 23440 6330 23540 6346
rect 23440 6296 23456 6330
rect 23524 6296 23540 6330
rect 23440 6258 23540 6296
rect 23598 6330 23698 6346
rect 23598 6296 23614 6330
rect 23682 6296 23698 6330
rect 23598 6258 23698 6296
rect 23756 6330 23856 6346
rect 23756 6296 23772 6330
rect 23840 6296 23856 6330
rect 23756 6258 23856 6296
rect 23914 6330 24014 6346
rect 23914 6296 23930 6330
rect 23998 6296 24014 6330
rect 23914 6258 24014 6296
rect 24072 6330 24172 6346
rect 24072 6296 24088 6330
rect 24156 6296 24172 6330
rect 24072 6258 24172 6296
rect 24230 6330 24330 6346
rect 24230 6296 24246 6330
rect 24314 6296 24330 6330
rect 24230 6258 24330 6296
rect 24388 6330 24488 6346
rect 24388 6296 24404 6330
rect 24472 6296 24488 6330
rect 24388 6258 24488 6296
rect 24546 6330 24646 6346
rect 24546 6296 24562 6330
rect 24630 6296 24646 6330
rect 24546 6258 24646 6296
rect 24704 6330 24804 6346
rect 24704 6296 24720 6330
rect 24788 6296 24804 6330
rect 24704 6258 24804 6296
rect 24862 6330 24962 6346
rect 24862 6296 24878 6330
rect 24946 6296 24962 6330
rect 24862 6258 24962 6296
rect 25020 6330 25120 6346
rect 25020 6296 25036 6330
rect 25104 6296 25120 6330
rect 25020 6258 25120 6296
rect 25178 6330 25278 6346
rect 25178 6296 25194 6330
rect 25262 6296 25278 6330
rect 25178 6258 25278 6296
rect 25336 6330 25436 6346
rect 25336 6296 25352 6330
rect 25420 6296 25436 6330
rect 25336 6258 25436 6296
rect 25494 6330 25594 6346
rect 25494 6296 25510 6330
rect 25578 6296 25594 6330
rect 25494 6258 25594 6296
rect 25652 6330 25752 6346
rect 25652 6296 25668 6330
rect 25736 6296 25752 6330
rect 25652 6258 25752 6296
rect 25810 6330 25910 6346
rect 25810 6296 25826 6330
rect 25894 6296 25910 6330
rect 25810 6258 25910 6296
rect 21228 220 21328 258
rect 21228 186 21244 220
rect 21312 186 21328 220
rect 21228 170 21328 186
rect 21386 220 21486 258
rect 21386 186 21402 220
rect 21470 186 21486 220
rect 21386 170 21486 186
rect 21544 220 21644 258
rect 21544 186 21560 220
rect 21628 186 21644 220
rect 21544 170 21644 186
rect 21702 220 21802 258
rect 21702 186 21718 220
rect 21786 186 21802 220
rect 21702 170 21802 186
rect 21860 220 21960 258
rect 21860 186 21876 220
rect 21944 186 21960 220
rect 21860 170 21960 186
rect 22018 220 22118 258
rect 22018 186 22034 220
rect 22102 186 22118 220
rect 22018 170 22118 186
rect 22176 220 22276 258
rect 22176 186 22192 220
rect 22260 186 22276 220
rect 22176 170 22276 186
rect 22334 220 22434 258
rect 22334 186 22350 220
rect 22418 186 22434 220
rect 22334 170 22434 186
rect 22492 220 22592 258
rect 22492 186 22508 220
rect 22576 186 22592 220
rect 22492 170 22592 186
rect 22650 220 22750 258
rect 22650 186 22666 220
rect 22734 186 22750 220
rect 22650 170 22750 186
rect 22808 220 22908 258
rect 22808 186 22824 220
rect 22892 186 22908 220
rect 22808 170 22908 186
rect 22966 220 23066 258
rect 22966 186 22982 220
rect 23050 186 23066 220
rect 22966 170 23066 186
rect 23124 220 23224 258
rect 23124 186 23140 220
rect 23208 186 23224 220
rect 23124 170 23224 186
rect 23282 220 23382 258
rect 23282 186 23298 220
rect 23366 186 23382 220
rect 23282 170 23382 186
rect 23440 220 23540 258
rect 23440 186 23456 220
rect 23524 186 23540 220
rect 23440 170 23540 186
rect 23598 220 23698 258
rect 23598 186 23614 220
rect 23682 186 23698 220
rect 23598 170 23698 186
rect 23756 220 23856 258
rect 23756 186 23772 220
rect 23840 186 23856 220
rect 23756 170 23856 186
rect 23914 220 24014 258
rect 23914 186 23930 220
rect 23998 186 24014 220
rect 23914 170 24014 186
rect 24072 220 24172 258
rect 24072 186 24088 220
rect 24156 186 24172 220
rect 24072 170 24172 186
rect 24230 220 24330 258
rect 24230 186 24246 220
rect 24314 186 24330 220
rect 24230 170 24330 186
rect 24388 220 24488 258
rect 24388 186 24404 220
rect 24472 186 24488 220
rect 24388 170 24488 186
rect 24546 220 24646 258
rect 24546 186 24562 220
rect 24630 186 24646 220
rect 24546 170 24646 186
rect 24704 220 24804 258
rect 24704 186 24720 220
rect 24788 186 24804 220
rect 24704 170 24804 186
rect 24862 220 24962 258
rect 24862 186 24878 220
rect 24946 186 24962 220
rect 24862 170 24962 186
rect 25020 220 25120 258
rect 25020 186 25036 220
rect 25104 186 25120 220
rect 25020 170 25120 186
rect 25178 220 25278 258
rect 25178 186 25194 220
rect 25262 186 25278 220
rect 25178 170 25278 186
rect 25336 220 25436 258
rect 25336 186 25352 220
rect 25420 186 25436 220
rect 25336 170 25436 186
rect 25494 220 25594 258
rect 25494 186 25510 220
rect 25578 186 25594 220
rect 25494 170 25594 186
rect 25652 220 25752 258
rect 25652 186 25668 220
rect 25736 186 25752 220
rect 25652 170 25752 186
rect 25810 220 25910 258
rect 25810 186 25826 220
rect 25894 186 25910 220
rect 25810 170 25910 186
rect 228 -670 328 -654
rect 228 -704 244 -670
rect 312 -704 328 -670
rect 228 -742 328 -704
rect 386 -670 486 -654
rect 386 -704 402 -670
rect 470 -704 486 -670
rect 386 -742 486 -704
rect 544 -670 644 -654
rect 544 -704 560 -670
rect 628 -704 644 -670
rect 544 -742 644 -704
rect 702 -670 802 -654
rect 702 -704 718 -670
rect 786 -704 802 -670
rect 702 -742 802 -704
rect 860 -670 960 -654
rect 860 -704 876 -670
rect 944 -704 960 -670
rect 860 -742 960 -704
rect 1018 -670 1118 -654
rect 1018 -704 1034 -670
rect 1102 -704 1118 -670
rect 1018 -742 1118 -704
rect 1176 -670 1276 -654
rect 1176 -704 1192 -670
rect 1260 -704 1276 -670
rect 1176 -742 1276 -704
rect 1334 -670 1434 -654
rect 1334 -704 1350 -670
rect 1418 -704 1434 -670
rect 1334 -742 1434 -704
rect 1492 -670 1592 -654
rect 1492 -704 1508 -670
rect 1576 -704 1592 -670
rect 1492 -742 1592 -704
rect 1650 -670 1750 -654
rect 1650 -704 1666 -670
rect 1734 -704 1750 -670
rect 1650 -742 1750 -704
rect 1808 -670 1908 -654
rect 1808 -704 1824 -670
rect 1892 -704 1908 -670
rect 1808 -742 1908 -704
rect 1966 -670 2066 -654
rect 1966 -704 1982 -670
rect 2050 -704 2066 -670
rect 1966 -742 2066 -704
rect 2124 -670 2224 -654
rect 2124 -704 2140 -670
rect 2208 -704 2224 -670
rect 2124 -742 2224 -704
rect 2282 -670 2382 -654
rect 2282 -704 2298 -670
rect 2366 -704 2382 -670
rect 2282 -742 2382 -704
rect 2440 -670 2540 -654
rect 2440 -704 2456 -670
rect 2524 -704 2540 -670
rect 2440 -742 2540 -704
rect 2598 -670 2698 -654
rect 2598 -704 2614 -670
rect 2682 -704 2698 -670
rect 2598 -742 2698 -704
rect 2756 -670 2856 -654
rect 2756 -704 2772 -670
rect 2840 -704 2856 -670
rect 2756 -742 2856 -704
rect 2914 -670 3014 -654
rect 2914 -704 2930 -670
rect 2998 -704 3014 -670
rect 2914 -742 3014 -704
rect 3072 -670 3172 -654
rect 3072 -704 3088 -670
rect 3156 -704 3172 -670
rect 3072 -742 3172 -704
rect 3230 -670 3330 -654
rect 3230 -704 3246 -670
rect 3314 -704 3330 -670
rect 3230 -742 3330 -704
rect 3388 -670 3488 -654
rect 3388 -704 3404 -670
rect 3472 -704 3488 -670
rect 3388 -742 3488 -704
rect 3546 -670 3646 -654
rect 3546 -704 3562 -670
rect 3630 -704 3646 -670
rect 3546 -742 3646 -704
rect 3704 -670 3804 -654
rect 3704 -704 3720 -670
rect 3788 -704 3804 -670
rect 3704 -742 3804 -704
rect 3862 -670 3962 -654
rect 3862 -704 3878 -670
rect 3946 -704 3962 -670
rect 3862 -742 3962 -704
rect 4020 -670 4120 -654
rect 4020 -704 4036 -670
rect 4104 -704 4120 -670
rect 4020 -742 4120 -704
rect 4178 -670 4278 -654
rect 4178 -704 4194 -670
rect 4262 -704 4278 -670
rect 4178 -742 4278 -704
rect 4336 -670 4436 -654
rect 4336 -704 4352 -670
rect 4420 -704 4436 -670
rect 4336 -742 4436 -704
rect 4494 -670 4594 -654
rect 4494 -704 4510 -670
rect 4578 -704 4594 -670
rect 4494 -742 4594 -704
rect 4652 -670 4752 -654
rect 4652 -704 4668 -670
rect 4736 -704 4752 -670
rect 4652 -742 4752 -704
rect 4810 -670 4910 -654
rect 4810 -704 4826 -670
rect 4894 -704 4910 -670
rect 4810 -742 4910 -704
rect 228 -6780 328 -6742
rect 228 -6814 244 -6780
rect 312 -6814 328 -6780
rect 228 -6830 328 -6814
rect 386 -6780 486 -6742
rect 386 -6814 402 -6780
rect 470 -6814 486 -6780
rect 386 -6830 486 -6814
rect 544 -6780 644 -6742
rect 544 -6814 560 -6780
rect 628 -6814 644 -6780
rect 544 -6830 644 -6814
rect 702 -6780 802 -6742
rect 702 -6814 718 -6780
rect 786 -6814 802 -6780
rect 702 -6830 802 -6814
rect 860 -6780 960 -6742
rect 860 -6814 876 -6780
rect 944 -6814 960 -6780
rect 860 -6830 960 -6814
rect 1018 -6780 1118 -6742
rect 1018 -6814 1034 -6780
rect 1102 -6814 1118 -6780
rect 1018 -6830 1118 -6814
rect 1176 -6780 1276 -6742
rect 1176 -6814 1192 -6780
rect 1260 -6814 1276 -6780
rect 1176 -6830 1276 -6814
rect 1334 -6780 1434 -6742
rect 1334 -6814 1350 -6780
rect 1418 -6814 1434 -6780
rect 1334 -6830 1434 -6814
rect 1492 -6780 1592 -6742
rect 1492 -6814 1508 -6780
rect 1576 -6814 1592 -6780
rect 1492 -6830 1592 -6814
rect 1650 -6780 1750 -6742
rect 1650 -6814 1666 -6780
rect 1734 -6814 1750 -6780
rect 1650 -6830 1750 -6814
rect 1808 -6780 1908 -6742
rect 1808 -6814 1824 -6780
rect 1892 -6814 1908 -6780
rect 1808 -6830 1908 -6814
rect 1966 -6780 2066 -6742
rect 1966 -6814 1982 -6780
rect 2050 -6814 2066 -6780
rect 1966 -6830 2066 -6814
rect 2124 -6780 2224 -6742
rect 2124 -6814 2140 -6780
rect 2208 -6814 2224 -6780
rect 2124 -6830 2224 -6814
rect 2282 -6780 2382 -6742
rect 2282 -6814 2298 -6780
rect 2366 -6814 2382 -6780
rect 2282 -6830 2382 -6814
rect 2440 -6780 2540 -6742
rect 2440 -6814 2456 -6780
rect 2524 -6814 2540 -6780
rect 2440 -6830 2540 -6814
rect 2598 -6780 2698 -6742
rect 2598 -6814 2614 -6780
rect 2682 -6814 2698 -6780
rect 2598 -6830 2698 -6814
rect 2756 -6780 2856 -6742
rect 2756 -6814 2772 -6780
rect 2840 -6814 2856 -6780
rect 2756 -6830 2856 -6814
rect 2914 -6780 3014 -6742
rect 2914 -6814 2930 -6780
rect 2998 -6814 3014 -6780
rect 2914 -6830 3014 -6814
rect 3072 -6780 3172 -6742
rect 3072 -6814 3088 -6780
rect 3156 -6814 3172 -6780
rect 3072 -6830 3172 -6814
rect 3230 -6780 3330 -6742
rect 3230 -6814 3246 -6780
rect 3314 -6814 3330 -6780
rect 3230 -6830 3330 -6814
rect 3388 -6780 3488 -6742
rect 3388 -6814 3404 -6780
rect 3472 -6814 3488 -6780
rect 3388 -6830 3488 -6814
rect 3546 -6780 3646 -6742
rect 3546 -6814 3562 -6780
rect 3630 -6814 3646 -6780
rect 3546 -6830 3646 -6814
rect 3704 -6780 3804 -6742
rect 3704 -6814 3720 -6780
rect 3788 -6814 3804 -6780
rect 3704 -6830 3804 -6814
rect 3862 -6780 3962 -6742
rect 3862 -6814 3878 -6780
rect 3946 -6814 3962 -6780
rect 3862 -6830 3962 -6814
rect 4020 -6780 4120 -6742
rect 4020 -6814 4036 -6780
rect 4104 -6814 4120 -6780
rect 4020 -6830 4120 -6814
rect 4178 -6780 4278 -6742
rect 4178 -6814 4194 -6780
rect 4262 -6814 4278 -6780
rect 4178 -6830 4278 -6814
rect 4336 -6780 4436 -6742
rect 4336 -6814 4352 -6780
rect 4420 -6814 4436 -6780
rect 4336 -6830 4436 -6814
rect 4494 -6780 4594 -6742
rect 4494 -6814 4510 -6780
rect 4578 -6814 4594 -6780
rect 4494 -6830 4594 -6814
rect 4652 -6780 4752 -6742
rect 4652 -6814 4668 -6780
rect 4736 -6814 4752 -6780
rect 4652 -6830 4752 -6814
rect 4810 -6780 4910 -6742
rect 4810 -6814 4826 -6780
rect 4894 -6814 4910 -6780
rect 4810 -6830 4910 -6814
rect 7228 -670 7328 -654
rect 7228 -704 7244 -670
rect 7312 -704 7328 -670
rect 7228 -742 7328 -704
rect 7386 -670 7486 -654
rect 7386 -704 7402 -670
rect 7470 -704 7486 -670
rect 7386 -742 7486 -704
rect 7544 -670 7644 -654
rect 7544 -704 7560 -670
rect 7628 -704 7644 -670
rect 7544 -742 7644 -704
rect 7702 -670 7802 -654
rect 7702 -704 7718 -670
rect 7786 -704 7802 -670
rect 7702 -742 7802 -704
rect 7860 -670 7960 -654
rect 7860 -704 7876 -670
rect 7944 -704 7960 -670
rect 7860 -742 7960 -704
rect 8018 -670 8118 -654
rect 8018 -704 8034 -670
rect 8102 -704 8118 -670
rect 8018 -742 8118 -704
rect 8176 -670 8276 -654
rect 8176 -704 8192 -670
rect 8260 -704 8276 -670
rect 8176 -742 8276 -704
rect 8334 -670 8434 -654
rect 8334 -704 8350 -670
rect 8418 -704 8434 -670
rect 8334 -742 8434 -704
rect 8492 -670 8592 -654
rect 8492 -704 8508 -670
rect 8576 -704 8592 -670
rect 8492 -742 8592 -704
rect 8650 -670 8750 -654
rect 8650 -704 8666 -670
rect 8734 -704 8750 -670
rect 8650 -742 8750 -704
rect 8808 -670 8908 -654
rect 8808 -704 8824 -670
rect 8892 -704 8908 -670
rect 8808 -742 8908 -704
rect 8966 -670 9066 -654
rect 8966 -704 8982 -670
rect 9050 -704 9066 -670
rect 8966 -742 9066 -704
rect 9124 -670 9224 -654
rect 9124 -704 9140 -670
rect 9208 -704 9224 -670
rect 9124 -742 9224 -704
rect 9282 -670 9382 -654
rect 9282 -704 9298 -670
rect 9366 -704 9382 -670
rect 9282 -742 9382 -704
rect 9440 -670 9540 -654
rect 9440 -704 9456 -670
rect 9524 -704 9540 -670
rect 9440 -742 9540 -704
rect 9598 -670 9698 -654
rect 9598 -704 9614 -670
rect 9682 -704 9698 -670
rect 9598 -742 9698 -704
rect 9756 -670 9856 -654
rect 9756 -704 9772 -670
rect 9840 -704 9856 -670
rect 9756 -742 9856 -704
rect 9914 -670 10014 -654
rect 9914 -704 9930 -670
rect 9998 -704 10014 -670
rect 9914 -742 10014 -704
rect 10072 -670 10172 -654
rect 10072 -704 10088 -670
rect 10156 -704 10172 -670
rect 10072 -742 10172 -704
rect 10230 -670 10330 -654
rect 10230 -704 10246 -670
rect 10314 -704 10330 -670
rect 10230 -742 10330 -704
rect 10388 -670 10488 -654
rect 10388 -704 10404 -670
rect 10472 -704 10488 -670
rect 10388 -742 10488 -704
rect 10546 -670 10646 -654
rect 10546 -704 10562 -670
rect 10630 -704 10646 -670
rect 10546 -742 10646 -704
rect 10704 -670 10804 -654
rect 10704 -704 10720 -670
rect 10788 -704 10804 -670
rect 10704 -742 10804 -704
rect 10862 -670 10962 -654
rect 10862 -704 10878 -670
rect 10946 -704 10962 -670
rect 10862 -742 10962 -704
rect 11020 -670 11120 -654
rect 11020 -704 11036 -670
rect 11104 -704 11120 -670
rect 11020 -742 11120 -704
rect 11178 -670 11278 -654
rect 11178 -704 11194 -670
rect 11262 -704 11278 -670
rect 11178 -742 11278 -704
rect 11336 -670 11436 -654
rect 11336 -704 11352 -670
rect 11420 -704 11436 -670
rect 11336 -742 11436 -704
rect 11494 -670 11594 -654
rect 11494 -704 11510 -670
rect 11578 -704 11594 -670
rect 11494 -742 11594 -704
rect 11652 -670 11752 -654
rect 11652 -704 11668 -670
rect 11736 -704 11752 -670
rect 11652 -742 11752 -704
rect 11810 -670 11910 -654
rect 11810 -704 11826 -670
rect 11894 -704 11910 -670
rect 11810 -742 11910 -704
rect 7228 -6780 7328 -6742
rect 7228 -6814 7244 -6780
rect 7312 -6814 7328 -6780
rect 7228 -6830 7328 -6814
rect 7386 -6780 7486 -6742
rect 7386 -6814 7402 -6780
rect 7470 -6814 7486 -6780
rect 7386 -6830 7486 -6814
rect 7544 -6780 7644 -6742
rect 7544 -6814 7560 -6780
rect 7628 -6814 7644 -6780
rect 7544 -6830 7644 -6814
rect 7702 -6780 7802 -6742
rect 7702 -6814 7718 -6780
rect 7786 -6814 7802 -6780
rect 7702 -6830 7802 -6814
rect 7860 -6780 7960 -6742
rect 7860 -6814 7876 -6780
rect 7944 -6814 7960 -6780
rect 7860 -6830 7960 -6814
rect 8018 -6780 8118 -6742
rect 8018 -6814 8034 -6780
rect 8102 -6814 8118 -6780
rect 8018 -6830 8118 -6814
rect 8176 -6780 8276 -6742
rect 8176 -6814 8192 -6780
rect 8260 -6814 8276 -6780
rect 8176 -6830 8276 -6814
rect 8334 -6780 8434 -6742
rect 8334 -6814 8350 -6780
rect 8418 -6814 8434 -6780
rect 8334 -6830 8434 -6814
rect 8492 -6780 8592 -6742
rect 8492 -6814 8508 -6780
rect 8576 -6814 8592 -6780
rect 8492 -6830 8592 -6814
rect 8650 -6780 8750 -6742
rect 8650 -6814 8666 -6780
rect 8734 -6814 8750 -6780
rect 8650 -6830 8750 -6814
rect 8808 -6780 8908 -6742
rect 8808 -6814 8824 -6780
rect 8892 -6814 8908 -6780
rect 8808 -6830 8908 -6814
rect 8966 -6780 9066 -6742
rect 8966 -6814 8982 -6780
rect 9050 -6814 9066 -6780
rect 8966 -6830 9066 -6814
rect 9124 -6780 9224 -6742
rect 9124 -6814 9140 -6780
rect 9208 -6814 9224 -6780
rect 9124 -6830 9224 -6814
rect 9282 -6780 9382 -6742
rect 9282 -6814 9298 -6780
rect 9366 -6814 9382 -6780
rect 9282 -6830 9382 -6814
rect 9440 -6780 9540 -6742
rect 9440 -6814 9456 -6780
rect 9524 -6814 9540 -6780
rect 9440 -6830 9540 -6814
rect 9598 -6780 9698 -6742
rect 9598 -6814 9614 -6780
rect 9682 -6814 9698 -6780
rect 9598 -6830 9698 -6814
rect 9756 -6780 9856 -6742
rect 9756 -6814 9772 -6780
rect 9840 -6814 9856 -6780
rect 9756 -6830 9856 -6814
rect 9914 -6780 10014 -6742
rect 9914 -6814 9930 -6780
rect 9998 -6814 10014 -6780
rect 9914 -6830 10014 -6814
rect 10072 -6780 10172 -6742
rect 10072 -6814 10088 -6780
rect 10156 -6814 10172 -6780
rect 10072 -6830 10172 -6814
rect 10230 -6780 10330 -6742
rect 10230 -6814 10246 -6780
rect 10314 -6814 10330 -6780
rect 10230 -6830 10330 -6814
rect 10388 -6780 10488 -6742
rect 10388 -6814 10404 -6780
rect 10472 -6814 10488 -6780
rect 10388 -6830 10488 -6814
rect 10546 -6780 10646 -6742
rect 10546 -6814 10562 -6780
rect 10630 -6814 10646 -6780
rect 10546 -6830 10646 -6814
rect 10704 -6780 10804 -6742
rect 10704 -6814 10720 -6780
rect 10788 -6814 10804 -6780
rect 10704 -6830 10804 -6814
rect 10862 -6780 10962 -6742
rect 10862 -6814 10878 -6780
rect 10946 -6814 10962 -6780
rect 10862 -6830 10962 -6814
rect 11020 -6780 11120 -6742
rect 11020 -6814 11036 -6780
rect 11104 -6814 11120 -6780
rect 11020 -6830 11120 -6814
rect 11178 -6780 11278 -6742
rect 11178 -6814 11194 -6780
rect 11262 -6814 11278 -6780
rect 11178 -6830 11278 -6814
rect 11336 -6780 11436 -6742
rect 11336 -6814 11352 -6780
rect 11420 -6814 11436 -6780
rect 11336 -6830 11436 -6814
rect 11494 -6780 11594 -6742
rect 11494 -6814 11510 -6780
rect 11578 -6814 11594 -6780
rect 11494 -6830 11594 -6814
rect 11652 -6780 11752 -6742
rect 11652 -6814 11668 -6780
rect 11736 -6814 11752 -6780
rect 11652 -6830 11752 -6814
rect 11810 -6780 11910 -6742
rect 11810 -6814 11826 -6780
rect 11894 -6814 11910 -6780
rect 11810 -6830 11910 -6814
rect 14228 -670 14328 -654
rect 14228 -704 14244 -670
rect 14312 -704 14328 -670
rect 14228 -742 14328 -704
rect 14386 -670 14486 -654
rect 14386 -704 14402 -670
rect 14470 -704 14486 -670
rect 14386 -742 14486 -704
rect 14544 -670 14644 -654
rect 14544 -704 14560 -670
rect 14628 -704 14644 -670
rect 14544 -742 14644 -704
rect 14702 -670 14802 -654
rect 14702 -704 14718 -670
rect 14786 -704 14802 -670
rect 14702 -742 14802 -704
rect 14860 -670 14960 -654
rect 14860 -704 14876 -670
rect 14944 -704 14960 -670
rect 14860 -742 14960 -704
rect 15018 -670 15118 -654
rect 15018 -704 15034 -670
rect 15102 -704 15118 -670
rect 15018 -742 15118 -704
rect 15176 -670 15276 -654
rect 15176 -704 15192 -670
rect 15260 -704 15276 -670
rect 15176 -742 15276 -704
rect 15334 -670 15434 -654
rect 15334 -704 15350 -670
rect 15418 -704 15434 -670
rect 15334 -742 15434 -704
rect 15492 -670 15592 -654
rect 15492 -704 15508 -670
rect 15576 -704 15592 -670
rect 15492 -742 15592 -704
rect 15650 -670 15750 -654
rect 15650 -704 15666 -670
rect 15734 -704 15750 -670
rect 15650 -742 15750 -704
rect 15808 -670 15908 -654
rect 15808 -704 15824 -670
rect 15892 -704 15908 -670
rect 15808 -742 15908 -704
rect 15966 -670 16066 -654
rect 15966 -704 15982 -670
rect 16050 -704 16066 -670
rect 15966 -742 16066 -704
rect 16124 -670 16224 -654
rect 16124 -704 16140 -670
rect 16208 -704 16224 -670
rect 16124 -742 16224 -704
rect 16282 -670 16382 -654
rect 16282 -704 16298 -670
rect 16366 -704 16382 -670
rect 16282 -742 16382 -704
rect 16440 -670 16540 -654
rect 16440 -704 16456 -670
rect 16524 -704 16540 -670
rect 16440 -742 16540 -704
rect 16598 -670 16698 -654
rect 16598 -704 16614 -670
rect 16682 -704 16698 -670
rect 16598 -742 16698 -704
rect 16756 -670 16856 -654
rect 16756 -704 16772 -670
rect 16840 -704 16856 -670
rect 16756 -742 16856 -704
rect 16914 -670 17014 -654
rect 16914 -704 16930 -670
rect 16998 -704 17014 -670
rect 16914 -742 17014 -704
rect 17072 -670 17172 -654
rect 17072 -704 17088 -670
rect 17156 -704 17172 -670
rect 17072 -742 17172 -704
rect 17230 -670 17330 -654
rect 17230 -704 17246 -670
rect 17314 -704 17330 -670
rect 17230 -742 17330 -704
rect 17388 -670 17488 -654
rect 17388 -704 17404 -670
rect 17472 -704 17488 -670
rect 17388 -742 17488 -704
rect 17546 -670 17646 -654
rect 17546 -704 17562 -670
rect 17630 -704 17646 -670
rect 17546 -742 17646 -704
rect 17704 -670 17804 -654
rect 17704 -704 17720 -670
rect 17788 -704 17804 -670
rect 17704 -742 17804 -704
rect 17862 -670 17962 -654
rect 17862 -704 17878 -670
rect 17946 -704 17962 -670
rect 17862 -742 17962 -704
rect 18020 -670 18120 -654
rect 18020 -704 18036 -670
rect 18104 -704 18120 -670
rect 18020 -742 18120 -704
rect 18178 -670 18278 -654
rect 18178 -704 18194 -670
rect 18262 -704 18278 -670
rect 18178 -742 18278 -704
rect 18336 -670 18436 -654
rect 18336 -704 18352 -670
rect 18420 -704 18436 -670
rect 18336 -742 18436 -704
rect 18494 -670 18594 -654
rect 18494 -704 18510 -670
rect 18578 -704 18594 -670
rect 18494 -742 18594 -704
rect 18652 -670 18752 -654
rect 18652 -704 18668 -670
rect 18736 -704 18752 -670
rect 18652 -742 18752 -704
rect 18810 -670 18910 -654
rect 18810 -704 18826 -670
rect 18894 -704 18910 -670
rect 18810 -742 18910 -704
rect 14228 -6780 14328 -6742
rect 14228 -6814 14244 -6780
rect 14312 -6814 14328 -6780
rect 14228 -6830 14328 -6814
rect 14386 -6780 14486 -6742
rect 14386 -6814 14402 -6780
rect 14470 -6814 14486 -6780
rect 14386 -6830 14486 -6814
rect 14544 -6780 14644 -6742
rect 14544 -6814 14560 -6780
rect 14628 -6814 14644 -6780
rect 14544 -6830 14644 -6814
rect 14702 -6780 14802 -6742
rect 14702 -6814 14718 -6780
rect 14786 -6814 14802 -6780
rect 14702 -6830 14802 -6814
rect 14860 -6780 14960 -6742
rect 14860 -6814 14876 -6780
rect 14944 -6814 14960 -6780
rect 14860 -6830 14960 -6814
rect 15018 -6780 15118 -6742
rect 15018 -6814 15034 -6780
rect 15102 -6814 15118 -6780
rect 15018 -6830 15118 -6814
rect 15176 -6780 15276 -6742
rect 15176 -6814 15192 -6780
rect 15260 -6814 15276 -6780
rect 15176 -6830 15276 -6814
rect 15334 -6780 15434 -6742
rect 15334 -6814 15350 -6780
rect 15418 -6814 15434 -6780
rect 15334 -6830 15434 -6814
rect 15492 -6780 15592 -6742
rect 15492 -6814 15508 -6780
rect 15576 -6814 15592 -6780
rect 15492 -6830 15592 -6814
rect 15650 -6780 15750 -6742
rect 15650 -6814 15666 -6780
rect 15734 -6814 15750 -6780
rect 15650 -6830 15750 -6814
rect 15808 -6780 15908 -6742
rect 15808 -6814 15824 -6780
rect 15892 -6814 15908 -6780
rect 15808 -6830 15908 -6814
rect 15966 -6780 16066 -6742
rect 15966 -6814 15982 -6780
rect 16050 -6814 16066 -6780
rect 15966 -6830 16066 -6814
rect 16124 -6780 16224 -6742
rect 16124 -6814 16140 -6780
rect 16208 -6814 16224 -6780
rect 16124 -6830 16224 -6814
rect 16282 -6780 16382 -6742
rect 16282 -6814 16298 -6780
rect 16366 -6814 16382 -6780
rect 16282 -6830 16382 -6814
rect 16440 -6780 16540 -6742
rect 16440 -6814 16456 -6780
rect 16524 -6814 16540 -6780
rect 16440 -6830 16540 -6814
rect 16598 -6780 16698 -6742
rect 16598 -6814 16614 -6780
rect 16682 -6814 16698 -6780
rect 16598 -6830 16698 -6814
rect 16756 -6780 16856 -6742
rect 16756 -6814 16772 -6780
rect 16840 -6814 16856 -6780
rect 16756 -6830 16856 -6814
rect 16914 -6780 17014 -6742
rect 16914 -6814 16930 -6780
rect 16998 -6814 17014 -6780
rect 16914 -6830 17014 -6814
rect 17072 -6780 17172 -6742
rect 17072 -6814 17088 -6780
rect 17156 -6814 17172 -6780
rect 17072 -6830 17172 -6814
rect 17230 -6780 17330 -6742
rect 17230 -6814 17246 -6780
rect 17314 -6814 17330 -6780
rect 17230 -6830 17330 -6814
rect 17388 -6780 17488 -6742
rect 17388 -6814 17404 -6780
rect 17472 -6814 17488 -6780
rect 17388 -6830 17488 -6814
rect 17546 -6780 17646 -6742
rect 17546 -6814 17562 -6780
rect 17630 -6814 17646 -6780
rect 17546 -6830 17646 -6814
rect 17704 -6780 17804 -6742
rect 17704 -6814 17720 -6780
rect 17788 -6814 17804 -6780
rect 17704 -6830 17804 -6814
rect 17862 -6780 17962 -6742
rect 17862 -6814 17878 -6780
rect 17946 -6814 17962 -6780
rect 17862 -6830 17962 -6814
rect 18020 -6780 18120 -6742
rect 18020 -6814 18036 -6780
rect 18104 -6814 18120 -6780
rect 18020 -6830 18120 -6814
rect 18178 -6780 18278 -6742
rect 18178 -6814 18194 -6780
rect 18262 -6814 18278 -6780
rect 18178 -6830 18278 -6814
rect 18336 -6780 18436 -6742
rect 18336 -6814 18352 -6780
rect 18420 -6814 18436 -6780
rect 18336 -6830 18436 -6814
rect 18494 -6780 18594 -6742
rect 18494 -6814 18510 -6780
rect 18578 -6814 18594 -6780
rect 18494 -6830 18594 -6814
rect 18652 -6780 18752 -6742
rect 18652 -6814 18668 -6780
rect 18736 -6814 18752 -6780
rect 18652 -6830 18752 -6814
rect 18810 -6780 18910 -6742
rect 18810 -6814 18826 -6780
rect 18894 -6814 18910 -6780
rect 18810 -6830 18910 -6814
rect 21228 -670 21328 -654
rect 21228 -704 21244 -670
rect 21312 -704 21328 -670
rect 21228 -742 21328 -704
rect 21386 -670 21486 -654
rect 21386 -704 21402 -670
rect 21470 -704 21486 -670
rect 21386 -742 21486 -704
rect 21544 -670 21644 -654
rect 21544 -704 21560 -670
rect 21628 -704 21644 -670
rect 21544 -742 21644 -704
rect 21702 -670 21802 -654
rect 21702 -704 21718 -670
rect 21786 -704 21802 -670
rect 21702 -742 21802 -704
rect 21860 -670 21960 -654
rect 21860 -704 21876 -670
rect 21944 -704 21960 -670
rect 21860 -742 21960 -704
rect 22018 -670 22118 -654
rect 22018 -704 22034 -670
rect 22102 -704 22118 -670
rect 22018 -742 22118 -704
rect 22176 -670 22276 -654
rect 22176 -704 22192 -670
rect 22260 -704 22276 -670
rect 22176 -742 22276 -704
rect 22334 -670 22434 -654
rect 22334 -704 22350 -670
rect 22418 -704 22434 -670
rect 22334 -742 22434 -704
rect 22492 -670 22592 -654
rect 22492 -704 22508 -670
rect 22576 -704 22592 -670
rect 22492 -742 22592 -704
rect 22650 -670 22750 -654
rect 22650 -704 22666 -670
rect 22734 -704 22750 -670
rect 22650 -742 22750 -704
rect 22808 -670 22908 -654
rect 22808 -704 22824 -670
rect 22892 -704 22908 -670
rect 22808 -742 22908 -704
rect 22966 -670 23066 -654
rect 22966 -704 22982 -670
rect 23050 -704 23066 -670
rect 22966 -742 23066 -704
rect 23124 -670 23224 -654
rect 23124 -704 23140 -670
rect 23208 -704 23224 -670
rect 23124 -742 23224 -704
rect 23282 -670 23382 -654
rect 23282 -704 23298 -670
rect 23366 -704 23382 -670
rect 23282 -742 23382 -704
rect 23440 -670 23540 -654
rect 23440 -704 23456 -670
rect 23524 -704 23540 -670
rect 23440 -742 23540 -704
rect 23598 -670 23698 -654
rect 23598 -704 23614 -670
rect 23682 -704 23698 -670
rect 23598 -742 23698 -704
rect 23756 -670 23856 -654
rect 23756 -704 23772 -670
rect 23840 -704 23856 -670
rect 23756 -742 23856 -704
rect 23914 -670 24014 -654
rect 23914 -704 23930 -670
rect 23998 -704 24014 -670
rect 23914 -742 24014 -704
rect 24072 -670 24172 -654
rect 24072 -704 24088 -670
rect 24156 -704 24172 -670
rect 24072 -742 24172 -704
rect 24230 -670 24330 -654
rect 24230 -704 24246 -670
rect 24314 -704 24330 -670
rect 24230 -742 24330 -704
rect 24388 -670 24488 -654
rect 24388 -704 24404 -670
rect 24472 -704 24488 -670
rect 24388 -742 24488 -704
rect 24546 -670 24646 -654
rect 24546 -704 24562 -670
rect 24630 -704 24646 -670
rect 24546 -742 24646 -704
rect 24704 -670 24804 -654
rect 24704 -704 24720 -670
rect 24788 -704 24804 -670
rect 24704 -742 24804 -704
rect 24862 -670 24962 -654
rect 24862 -704 24878 -670
rect 24946 -704 24962 -670
rect 24862 -742 24962 -704
rect 25020 -670 25120 -654
rect 25020 -704 25036 -670
rect 25104 -704 25120 -670
rect 25020 -742 25120 -704
rect 25178 -670 25278 -654
rect 25178 -704 25194 -670
rect 25262 -704 25278 -670
rect 25178 -742 25278 -704
rect 25336 -670 25436 -654
rect 25336 -704 25352 -670
rect 25420 -704 25436 -670
rect 25336 -742 25436 -704
rect 25494 -670 25594 -654
rect 25494 -704 25510 -670
rect 25578 -704 25594 -670
rect 25494 -742 25594 -704
rect 25652 -670 25752 -654
rect 25652 -704 25668 -670
rect 25736 -704 25752 -670
rect 25652 -742 25752 -704
rect 25810 -670 25910 -654
rect 25810 -704 25826 -670
rect 25894 -704 25910 -670
rect 25810 -742 25910 -704
rect 21228 -6780 21328 -6742
rect 21228 -6814 21244 -6780
rect 21312 -6814 21328 -6780
rect 21228 -6830 21328 -6814
rect 21386 -6780 21486 -6742
rect 21386 -6814 21402 -6780
rect 21470 -6814 21486 -6780
rect 21386 -6830 21486 -6814
rect 21544 -6780 21644 -6742
rect 21544 -6814 21560 -6780
rect 21628 -6814 21644 -6780
rect 21544 -6830 21644 -6814
rect 21702 -6780 21802 -6742
rect 21702 -6814 21718 -6780
rect 21786 -6814 21802 -6780
rect 21702 -6830 21802 -6814
rect 21860 -6780 21960 -6742
rect 21860 -6814 21876 -6780
rect 21944 -6814 21960 -6780
rect 21860 -6830 21960 -6814
rect 22018 -6780 22118 -6742
rect 22018 -6814 22034 -6780
rect 22102 -6814 22118 -6780
rect 22018 -6830 22118 -6814
rect 22176 -6780 22276 -6742
rect 22176 -6814 22192 -6780
rect 22260 -6814 22276 -6780
rect 22176 -6830 22276 -6814
rect 22334 -6780 22434 -6742
rect 22334 -6814 22350 -6780
rect 22418 -6814 22434 -6780
rect 22334 -6830 22434 -6814
rect 22492 -6780 22592 -6742
rect 22492 -6814 22508 -6780
rect 22576 -6814 22592 -6780
rect 22492 -6830 22592 -6814
rect 22650 -6780 22750 -6742
rect 22650 -6814 22666 -6780
rect 22734 -6814 22750 -6780
rect 22650 -6830 22750 -6814
rect 22808 -6780 22908 -6742
rect 22808 -6814 22824 -6780
rect 22892 -6814 22908 -6780
rect 22808 -6830 22908 -6814
rect 22966 -6780 23066 -6742
rect 22966 -6814 22982 -6780
rect 23050 -6814 23066 -6780
rect 22966 -6830 23066 -6814
rect 23124 -6780 23224 -6742
rect 23124 -6814 23140 -6780
rect 23208 -6814 23224 -6780
rect 23124 -6830 23224 -6814
rect 23282 -6780 23382 -6742
rect 23282 -6814 23298 -6780
rect 23366 -6814 23382 -6780
rect 23282 -6830 23382 -6814
rect 23440 -6780 23540 -6742
rect 23440 -6814 23456 -6780
rect 23524 -6814 23540 -6780
rect 23440 -6830 23540 -6814
rect 23598 -6780 23698 -6742
rect 23598 -6814 23614 -6780
rect 23682 -6814 23698 -6780
rect 23598 -6830 23698 -6814
rect 23756 -6780 23856 -6742
rect 23756 -6814 23772 -6780
rect 23840 -6814 23856 -6780
rect 23756 -6830 23856 -6814
rect 23914 -6780 24014 -6742
rect 23914 -6814 23930 -6780
rect 23998 -6814 24014 -6780
rect 23914 -6830 24014 -6814
rect 24072 -6780 24172 -6742
rect 24072 -6814 24088 -6780
rect 24156 -6814 24172 -6780
rect 24072 -6830 24172 -6814
rect 24230 -6780 24330 -6742
rect 24230 -6814 24246 -6780
rect 24314 -6814 24330 -6780
rect 24230 -6830 24330 -6814
rect 24388 -6780 24488 -6742
rect 24388 -6814 24404 -6780
rect 24472 -6814 24488 -6780
rect 24388 -6830 24488 -6814
rect 24546 -6780 24646 -6742
rect 24546 -6814 24562 -6780
rect 24630 -6814 24646 -6780
rect 24546 -6830 24646 -6814
rect 24704 -6780 24804 -6742
rect 24704 -6814 24720 -6780
rect 24788 -6814 24804 -6780
rect 24704 -6830 24804 -6814
rect 24862 -6780 24962 -6742
rect 24862 -6814 24878 -6780
rect 24946 -6814 24962 -6780
rect 24862 -6830 24962 -6814
rect 25020 -6780 25120 -6742
rect 25020 -6814 25036 -6780
rect 25104 -6814 25120 -6780
rect 25020 -6830 25120 -6814
rect 25178 -6780 25278 -6742
rect 25178 -6814 25194 -6780
rect 25262 -6814 25278 -6780
rect 25178 -6830 25278 -6814
rect 25336 -6780 25436 -6742
rect 25336 -6814 25352 -6780
rect 25420 -6814 25436 -6780
rect 25336 -6830 25436 -6814
rect 25494 -6780 25594 -6742
rect 25494 -6814 25510 -6780
rect 25578 -6814 25594 -6780
rect 25494 -6830 25594 -6814
rect 25652 -6780 25752 -6742
rect 25652 -6814 25668 -6780
rect 25736 -6814 25752 -6780
rect 25652 -6830 25752 -6814
rect 25810 -6780 25910 -6742
rect 25810 -6814 25826 -6780
rect 25894 -6814 25910 -6780
rect 25810 -6830 25910 -6814
<< polycont >>
rect 244 6296 312 6330
rect 402 6296 470 6330
rect 560 6296 628 6330
rect 718 6296 786 6330
rect 876 6296 944 6330
rect 1034 6296 1102 6330
rect 1192 6296 1260 6330
rect 1350 6296 1418 6330
rect 1508 6296 1576 6330
rect 1666 6296 1734 6330
rect 1824 6296 1892 6330
rect 1982 6296 2050 6330
rect 2140 6296 2208 6330
rect 2298 6296 2366 6330
rect 2456 6296 2524 6330
rect 2614 6296 2682 6330
rect 2772 6296 2840 6330
rect 2930 6296 2998 6330
rect 3088 6296 3156 6330
rect 3246 6296 3314 6330
rect 3404 6296 3472 6330
rect 3562 6296 3630 6330
rect 3720 6296 3788 6330
rect 3878 6296 3946 6330
rect 4036 6296 4104 6330
rect 4194 6296 4262 6330
rect 4352 6296 4420 6330
rect 4510 6296 4578 6330
rect 4668 6296 4736 6330
rect 4826 6296 4894 6330
rect 244 186 312 220
rect 402 186 470 220
rect 560 186 628 220
rect 718 186 786 220
rect 876 186 944 220
rect 1034 186 1102 220
rect 1192 186 1260 220
rect 1350 186 1418 220
rect 1508 186 1576 220
rect 1666 186 1734 220
rect 1824 186 1892 220
rect 1982 186 2050 220
rect 2140 186 2208 220
rect 2298 186 2366 220
rect 2456 186 2524 220
rect 2614 186 2682 220
rect 2772 186 2840 220
rect 2930 186 2998 220
rect 3088 186 3156 220
rect 3246 186 3314 220
rect 3404 186 3472 220
rect 3562 186 3630 220
rect 3720 186 3788 220
rect 3878 186 3946 220
rect 4036 186 4104 220
rect 4194 186 4262 220
rect 4352 186 4420 220
rect 4510 186 4578 220
rect 4668 186 4736 220
rect 4826 186 4894 220
rect 7244 6296 7312 6330
rect 7402 6296 7470 6330
rect 7560 6296 7628 6330
rect 7718 6296 7786 6330
rect 7876 6296 7944 6330
rect 8034 6296 8102 6330
rect 8192 6296 8260 6330
rect 8350 6296 8418 6330
rect 8508 6296 8576 6330
rect 8666 6296 8734 6330
rect 8824 6296 8892 6330
rect 8982 6296 9050 6330
rect 9140 6296 9208 6330
rect 9298 6296 9366 6330
rect 9456 6296 9524 6330
rect 9614 6296 9682 6330
rect 9772 6296 9840 6330
rect 9930 6296 9998 6330
rect 10088 6296 10156 6330
rect 10246 6296 10314 6330
rect 10404 6296 10472 6330
rect 10562 6296 10630 6330
rect 10720 6296 10788 6330
rect 10878 6296 10946 6330
rect 11036 6296 11104 6330
rect 11194 6296 11262 6330
rect 11352 6296 11420 6330
rect 11510 6296 11578 6330
rect 11668 6296 11736 6330
rect 11826 6296 11894 6330
rect 7244 186 7312 220
rect 7402 186 7470 220
rect 7560 186 7628 220
rect 7718 186 7786 220
rect 7876 186 7944 220
rect 8034 186 8102 220
rect 8192 186 8260 220
rect 8350 186 8418 220
rect 8508 186 8576 220
rect 8666 186 8734 220
rect 8824 186 8892 220
rect 8982 186 9050 220
rect 9140 186 9208 220
rect 9298 186 9366 220
rect 9456 186 9524 220
rect 9614 186 9682 220
rect 9772 186 9840 220
rect 9930 186 9998 220
rect 10088 186 10156 220
rect 10246 186 10314 220
rect 10404 186 10472 220
rect 10562 186 10630 220
rect 10720 186 10788 220
rect 10878 186 10946 220
rect 11036 186 11104 220
rect 11194 186 11262 220
rect 11352 186 11420 220
rect 11510 186 11578 220
rect 11668 186 11736 220
rect 11826 186 11894 220
rect 14244 6296 14312 6330
rect 14402 6296 14470 6330
rect 14560 6296 14628 6330
rect 14718 6296 14786 6330
rect 14876 6296 14944 6330
rect 15034 6296 15102 6330
rect 15192 6296 15260 6330
rect 15350 6296 15418 6330
rect 15508 6296 15576 6330
rect 15666 6296 15734 6330
rect 15824 6296 15892 6330
rect 15982 6296 16050 6330
rect 16140 6296 16208 6330
rect 16298 6296 16366 6330
rect 16456 6296 16524 6330
rect 16614 6296 16682 6330
rect 16772 6296 16840 6330
rect 16930 6296 16998 6330
rect 17088 6296 17156 6330
rect 17246 6296 17314 6330
rect 17404 6296 17472 6330
rect 17562 6296 17630 6330
rect 17720 6296 17788 6330
rect 17878 6296 17946 6330
rect 18036 6296 18104 6330
rect 18194 6296 18262 6330
rect 18352 6296 18420 6330
rect 18510 6296 18578 6330
rect 18668 6296 18736 6330
rect 18826 6296 18894 6330
rect 14244 186 14312 220
rect 14402 186 14470 220
rect 14560 186 14628 220
rect 14718 186 14786 220
rect 14876 186 14944 220
rect 15034 186 15102 220
rect 15192 186 15260 220
rect 15350 186 15418 220
rect 15508 186 15576 220
rect 15666 186 15734 220
rect 15824 186 15892 220
rect 15982 186 16050 220
rect 16140 186 16208 220
rect 16298 186 16366 220
rect 16456 186 16524 220
rect 16614 186 16682 220
rect 16772 186 16840 220
rect 16930 186 16998 220
rect 17088 186 17156 220
rect 17246 186 17314 220
rect 17404 186 17472 220
rect 17562 186 17630 220
rect 17720 186 17788 220
rect 17878 186 17946 220
rect 18036 186 18104 220
rect 18194 186 18262 220
rect 18352 186 18420 220
rect 18510 186 18578 220
rect 18668 186 18736 220
rect 18826 186 18894 220
rect 21244 6296 21312 6330
rect 21402 6296 21470 6330
rect 21560 6296 21628 6330
rect 21718 6296 21786 6330
rect 21876 6296 21944 6330
rect 22034 6296 22102 6330
rect 22192 6296 22260 6330
rect 22350 6296 22418 6330
rect 22508 6296 22576 6330
rect 22666 6296 22734 6330
rect 22824 6296 22892 6330
rect 22982 6296 23050 6330
rect 23140 6296 23208 6330
rect 23298 6296 23366 6330
rect 23456 6296 23524 6330
rect 23614 6296 23682 6330
rect 23772 6296 23840 6330
rect 23930 6296 23998 6330
rect 24088 6296 24156 6330
rect 24246 6296 24314 6330
rect 24404 6296 24472 6330
rect 24562 6296 24630 6330
rect 24720 6296 24788 6330
rect 24878 6296 24946 6330
rect 25036 6296 25104 6330
rect 25194 6296 25262 6330
rect 25352 6296 25420 6330
rect 25510 6296 25578 6330
rect 25668 6296 25736 6330
rect 25826 6296 25894 6330
rect 21244 186 21312 220
rect 21402 186 21470 220
rect 21560 186 21628 220
rect 21718 186 21786 220
rect 21876 186 21944 220
rect 22034 186 22102 220
rect 22192 186 22260 220
rect 22350 186 22418 220
rect 22508 186 22576 220
rect 22666 186 22734 220
rect 22824 186 22892 220
rect 22982 186 23050 220
rect 23140 186 23208 220
rect 23298 186 23366 220
rect 23456 186 23524 220
rect 23614 186 23682 220
rect 23772 186 23840 220
rect 23930 186 23998 220
rect 24088 186 24156 220
rect 24246 186 24314 220
rect 24404 186 24472 220
rect 24562 186 24630 220
rect 24720 186 24788 220
rect 24878 186 24946 220
rect 25036 186 25104 220
rect 25194 186 25262 220
rect 25352 186 25420 220
rect 25510 186 25578 220
rect 25668 186 25736 220
rect 25826 186 25894 220
rect 244 -704 312 -670
rect 402 -704 470 -670
rect 560 -704 628 -670
rect 718 -704 786 -670
rect 876 -704 944 -670
rect 1034 -704 1102 -670
rect 1192 -704 1260 -670
rect 1350 -704 1418 -670
rect 1508 -704 1576 -670
rect 1666 -704 1734 -670
rect 1824 -704 1892 -670
rect 1982 -704 2050 -670
rect 2140 -704 2208 -670
rect 2298 -704 2366 -670
rect 2456 -704 2524 -670
rect 2614 -704 2682 -670
rect 2772 -704 2840 -670
rect 2930 -704 2998 -670
rect 3088 -704 3156 -670
rect 3246 -704 3314 -670
rect 3404 -704 3472 -670
rect 3562 -704 3630 -670
rect 3720 -704 3788 -670
rect 3878 -704 3946 -670
rect 4036 -704 4104 -670
rect 4194 -704 4262 -670
rect 4352 -704 4420 -670
rect 4510 -704 4578 -670
rect 4668 -704 4736 -670
rect 4826 -704 4894 -670
rect 244 -6814 312 -6780
rect 402 -6814 470 -6780
rect 560 -6814 628 -6780
rect 718 -6814 786 -6780
rect 876 -6814 944 -6780
rect 1034 -6814 1102 -6780
rect 1192 -6814 1260 -6780
rect 1350 -6814 1418 -6780
rect 1508 -6814 1576 -6780
rect 1666 -6814 1734 -6780
rect 1824 -6814 1892 -6780
rect 1982 -6814 2050 -6780
rect 2140 -6814 2208 -6780
rect 2298 -6814 2366 -6780
rect 2456 -6814 2524 -6780
rect 2614 -6814 2682 -6780
rect 2772 -6814 2840 -6780
rect 2930 -6814 2998 -6780
rect 3088 -6814 3156 -6780
rect 3246 -6814 3314 -6780
rect 3404 -6814 3472 -6780
rect 3562 -6814 3630 -6780
rect 3720 -6814 3788 -6780
rect 3878 -6814 3946 -6780
rect 4036 -6814 4104 -6780
rect 4194 -6814 4262 -6780
rect 4352 -6814 4420 -6780
rect 4510 -6814 4578 -6780
rect 4668 -6814 4736 -6780
rect 4826 -6814 4894 -6780
rect 7244 -704 7312 -670
rect 7402 -704 7470 -670
rect 7560 -704 7628 -670
rect 7718 -704 7786 -670
rect 7876 -704 7944 -670
rect 8034 -704 8102 -670
rect 8192 -704 8260 -670
rect 8350 -704 8418 -670
rect 8508 -704 8576 -670
rect 8666 -704 8734 -670
rect 8824 -704 8892 -670
rect 8982 -704 9050 -670
rect 9140 -704 9208 -670
rect 9298 -704 9366 -670
rect 9456 -704 9524 -670
rect 9614 -704 9682 -670
rect 9772 -704 9840 -670
rect 9930 -704 9998 -670
rect 10088 -704 10156 -670
rect 10246 -704 10314 -670
rect 10404 -704 10472 -670
rect 10562 -704 10630 -670
rect 10720 -704 10788 -670
rect 10878 -704 10946 -670
rect 11036 -704 11104 -670
rect 11194 -704 11262 -670
rect 11352 -704 11420 -670
rect 11510 -704 11578 -670
rect 11668 -704 11736 -670
rect 11826 -704 11894 -670
rect 7244 -6814 7312 -6780
rect 7402 -6814 7470 -6780
rect 7560 -6814 7628 -6780
rect 7718 -6814 7786 -6780
rect 7876 -6814 7944 -6780
rect 8034 -6814 8102 -6780
rect 8192 -6814 8260 -6780
rect 8350 -6814 8418 -6780
rect 8508 -6814 8576 -6780
rect 8666 -6814 8734 -6780
rect 8824 -6814 8892 -6780
rect 8982 -6814 9050 -6780
rect 9140 -6814 9208 -6780
rect 9298 -6814 9366 -6780
rect 9456 -6814 9524 -6780
rect 9614 -6814 9682 -6780
rect 9772 -6814 9840 -6780
rect 9930 -6814 9998 -6780
rect 10088 -6814 10156 -6780
rect 10246 -6814 10314 -6780
rect 10404 -6814 10472 -6780
rect 10562 -6814 10630 -6780
rect 10720 -6814 10788 -6780
rect 10878 -6814 10946 -6780
rect 11036 -6814 11104 -6780
rect 11194 -6814 11262 -6780
rect 11352 -6814 11420 -6780
rect 11510 -6814 11578 -6780
rect 11668 -6814 11736 -6780
rect 11826 -6814 11894 -6780
rect 14244 -704 14312 -670
rect 14402 -704 14470 -670
rect 14560 -704 14628 -670
rect 14718 -704 14786 -670
rect 14876 -704 14944 -670
rect 15034 -704 15102 -670
rect 15192 -704 15260 -670
rect 15350 -704 15418 -670
rect 15508 -704 15576 -670
rect 15666 -704 15734 -670
rect 15824 -704 15892 -670
rect 15982 -704 16050 -670
rect 16140 -704 16208 -670
rect 16298 -704 16366 -670
rect 16456 -704 16524 -670
rect 16614 -704 16682 -670
rect 16772 -704 16840 -670
rect 16930 -704 16998 -670
rect 17088 -704 17156 -670
rect 17246 -704 17314 -670
rect 17404 -704 17472 -670
rect 17562 -704 17630 -670
rect 17720 -704 17788 -670
rect 17878 -704 17946 -670
rect 18036 -704 18104 -670
rect 18194 -704 18262 -670
rect 18352 -704 18420 -670
rect 18510 -704 18578 -670
rect 18668 -704 18736 -670
rect 18826 -704 18894 -670
rect 14244 -6814 14312 -6780
rect 14402 -6814 14470 -6780
rect 14560 -6814 14628 -6780
rect 14718 -6814 14786 -6780
rect 14876 -6814 14944 -6780
rect 15034 -6814 15102 -6780
rect 15192 -6814 15260 -6780
rect 15350 -6814 15418 -6780
rect 15508 -6814 15576 -6780
rect 15666 -6814 15734 -6780
rect 15824 -6814 15892 -6780
rect 15982 -6814 16050 -6780
rect 16140 -6814 16208 -6780
rect 16298 -6814 16366 -6780
rect 16456 -6814 16524 -6780
rect 16614 -6814 16682 -6780
rect 16772 -6814 16840 -6780
rect 16930 -6814 16998 -6780
rect 17088 -6814 17156 -6780
rect 17246 -6814 17314 -6780
rect 17404 -6814 17472 -6780
rect 17562 -6814 17630 -6780
rect 17720 -6814 17788 -6780
rect 17878 -6814 17946 -6780
rect 18036 -6814 18104 -6780
rect 18194 -6814 18262 -6780
rect 18352 -6814 18420 -6780
rect 18510 -6814 18578 -6780
rect 18668 -6814 18736 -6780
rect 18826 -6814 18894 -6780
rect 21244 -704 21312 -670
rect 21402 -704 21470 -670
rect 21560 -704 21628 -670
rect 21718 -704 21786 -670
rect 21876 -704 21944 -670
rect 22034 -704 22102 -670
rect 22192 -704 22260 -670
rect 22350 -704 22418 -670
rect 22508 -704 22576 -670
rect 22666 -704 22734 -670
rect 22824 -704 22892 -670
rect 22982 -704 23050 -670
rect 23140 -704 23208 -670
rect 23298 -704 23366 -670
rect 23456 -704 23524 -670
rect 23614 -704 23682 -670
rect 23772 -704 23840 -670
rect 23930 -704 23998 -670
rect 24088 -704 24156 -670
rect 24246 -704 24314 -670
rect 24404 -704 24472 -670
rect 24562 -704 24630 -670
rect 24720 -704 24788 -670
rect 24878 -704 24946 -670
rect 25036 -704 25104 -670
rect 25194 -704 25262 -670
rect 25352 -704 25420 -670
rect 25510 -704 25578 -670
rect 25668 -704 25736 -670
rect 25826 -704 25894 -670
rect 21244 -6814 21312 -6780
rect 21402 -6814 21470 -6780
rect 21560 -6814 21628 -6780
rect 21718 -6814 21786 -6780
rect 21876 -6814 21944 -6780
rect 22034 -6814 22102 -6780
rect 22192 -6814 22260 -6780
rect 22350 -6814 22418 -6780
rect 22508 -6814 22576 -6780
rect 22666 -6814 22734 -6780
rect 22824 -6814 22892 -6780
rect 22982 -6814 23050 -6780
rect 23140 -6814 23208 -6780
rect 23298 -6814 23366 -6780
rect 23456 -6814 23524 -6780
rect 23614 -6814 23682 -6780
rect 23772 -6814 23840 -6780
rect 23930 -6814 23998 -6780
rect 24088 -6814 24156 -6780
rect 24246 -6814 24314 -6780
rect 24404 -6814 24472 -6780
rect 24562 -6814 24630 -6780
rect 24720 -6814 24788 -6780
rect 24878 -6814 24946 -6780
rect 25036 -6814 25104 -6780
rect 25194 -6814 25262 -6780
rect 25352 -6814 25420 -6780
rect 25510 -6814 25578 -6780
rect 25668 -6814 25736 -6780
rect 25826 -6814 25894 -6780
<< locali >>
rect 48 6434 144 6468
rect 4994 6434 5090 6468
rect 48 6372 82 6434
rect 5056 6372 5090 6434
rect 228 6296 244 6330
rect 312 6296 328 6330
rect 386 6296 402 6330
rect 470 6296 486 6330
rect 544 6296 560 6330
rect 628 6296 644 6330
rect 702 6296 718 6330
rect 786 6296 802 6330
rect 860 6296 876 6330
rect 944 6296 960 6330
rect 1018 6296 1034 6330
rect 1102 6296 1118 6330
rect 1176 6296 1192 6330
rect 1260 6296 1276 6330
rect 1334 6296 1350 6330
rect 1418 6296 1434 6330
rect 1492 6296 1508 6330
rect 1576 6296 1592 6330
rect 1650 6296 1666 6330
rect 1734 6296 1750 6330
rect 1808 6296 1824 6330
rect 1892 6296 1908 6330
rect 1966 6296 1982 6330
rect 2050 6296 2066 6330
rect 2124 6296 2140 6330
rect 2208 6296 2224 6330
rect 2282 6296 2298 6330
rect 2366 6296 2382 6330
rect 2440 6296 2456 6330
rect 2524 6296 2540 6330
rect 2598 6296 2614 6330
rect 2682 6296 2698 6330
rect 2756 6296 2772 6330
rect 2840 6296 2856 6330
rect 2914 6296 2930 6330
rect 2998 6296 3014 6330
rect 3072 6296 3088 6330
rect 3156 6296 3172 6330
rect 3230 6296 3246 6330
rect 3314 6296 3330 6330
rect 3388 6296 3404 6330
rect 3472 6296 3488 6330
rect 3546 6296 3562 6330
rect 3630 6296 3646 6330
rect 3704 6296 3720 6330
rect 3788 6296 3804 6330
rect 3862 6296 3878 6330
rect 3946 6296 3962 6330
rect 4020 6296 4036 6330
rect 4104 6296 4120 6330
rect 4178 6296 4194 6330
rect 4262 6296 4278 6330
rect 4336 6296 4352 6330
rect 4420 6296 4436 6330
rect 4494 6296 4510 6330
rect 4578 6296 4594 6330
rect 4652 6296 4668 6330
rect 4736 6296 4752 6330
rect 4810 6296 4826 6330
rect 4894 6296 4910 6330
rect 7048 6434 7144 6468
rect 11994 6434 12090 6468
rect 7048 6372 7082 6434
rect 12056 6372 12090 6434
rect 7228 6296 7244 6330
rect 7312 6296 7328 6330
rect 7386 6296 7402 6330
rect 7470 6296 7486 6330
rect 7544 6296 7560 6330
rect 7628 6296 7644 6330
rect 7702 6296 7718 6330
rect 7786 6296 7802 6330
rect 7860 6296 7876 6330
rect 7944 6296 7960 6330
rect 8018 6296 8034 6330
rect 8102 6296 8118 6330
rect 8176 6296 8192 6330
rect 8260 6296 8276 6330
rect 8334 6296 8350 6330
rect 8418 6296 8434 6330
rect 8492 6296 8508 6330
rect 8576 6296 8592 6330
rect 8650 6296 8666 6330
rect 8734 6296 8750 6330
rect 8808 6296 8824 6330
rect 8892 6296 8908 6330
rect 8966 6296 8982 6330
rect 9050 6296 9066 6330
rect 9124 6296 9140 6330
rect 9208 6296 9224 6330
rect 9282 6296 9298 6330
rect 9366 6296 9382 6330
rect 9440 6296 9456 6330
rect 9524 6296 9540 6330
rect 9598 6296 9614 6330
rect 9682 6296 9698 6330
rect 9756 6296 9772 6330
rect 9840 6296 9856 6330
rect 9914 6296 9930 6330
rect 9998 6296 10014 6330
rect 10072 6296 10088 6330
rect 10156 6296 10172 6330
rect 10230 6296 10246 6330
rect 10314 6296 10330 6330
rect 10388 6296 10404 6330
rect 10472 6296 10488 6330
rect 10546 6296 10562 6330
rect 10630 6296 10646 6330
rect 10704 6296 10720 6330
rect 10788 6296 10804 6330
rect 10862 6296 10878 6330
rect 10946 6296 10962 6330
rect 11020 6296 11036 6330
rect 11104 6296 11120 6330
rect 11178 6296 11194 6330
rect 11262 6296 11278 6330
rect 11336 6296 11352 6330
rect 11420 6296 11436 6330
rect 11494 6296 11510 6330
rect 11578 6296 11594 6330
rect 11652 6296 11668 6330
rect 11736 6296 11752 6330
rect 11810 6296 11826 6330
rect 11894 6296 11910 6330
rect 14048 6434 14144 6468
rect 18994 6434 19090 6468
rect 14048 6372 14082 6434
rect 19056 6372 19090 6434
rect 14228 6296 14244 6330
rect 14312 6296 14328 6330
rect 14386 6296 14402 6330
rect 14470 6296 14486 6330
rect 14544 6296 14560 6330
rect 14628 6296 14644 6330
rect 14702 6296 14718 6330
rect 14786 6296 14802 6330
rect 14860 6296 14876 6330
rect 14944 6296 14960 6330
rect 15018 6296 15034 6330
rect 15102 6296 15118 6330
rect 15176 6296 15192 6330
rect 15260 6296 15276 6330
rect 15334 6296 15350 6330
rect 15418 6296 15434 6330
rect 15492 6296 15508 6330
rect 15576 6296 15592 6330
rect 15650 6296 15666 6330
rect 15734 6296 15750 6330
rect 15808 6296 15824 6330
rect 15892 6296 15908 6330
rect 15966 6296 15982 6330
rect 16050 6296 16066 6330
rect 16124 6296 16140 6330
rect 16208 6296 16224 6330
rect 16282 6296 16298 6330
rect 16366 6296 16382 6330
rect 16440 6296 16456 6330
rect 16524 6296 16540 6330
rect 16598 6296 16614 6330
rect 16682 6296 16698 6330
rect 16756 6296 16772 6330
rect 16840 6296 16856 6330
rect 16914 6296 16930 6330
rect 16998 6296 17014 6330
rect 17072 6296 17088 6330
rect 17156 6296 17172 6330
rect 17230 6296 17246 6330
rect 17314 6296 17330 6330
rect 17388 6296 17404 6330
rect 17472 6296 17488 6330
rect 17546 6296 17562 6330
rect 17630 6296 17646 6330
rect 17704 6296 17720 6330
rect 17788 6296 17804 6330
rect 17862 6296 17878 6330
rect 17946 6296 17962 6330
rect 18020 6296 18036 6330
rect 18104 6296 18120 6330
rect 18178 6296 18194 6330
rect 18262 6296 18278 6330
rect 18336 6296 18352 6330
rect 18420 6296 18436 6330
rect 18494 6296 18510 6330
rect 18578 6296 18594 6330
rect 18652 6296 18668 6330
rect 18736 6296 18752 6330
rect 18810 6296 18826 6330
rect 18894 6296 18910 6330
rect 21048 6434 21144 6468
rect 25994 6434 26090 6468
rect 21048 6372 21082 6434
rect 26056 6372 26090 6434
rect 21228 6296 21244 6330
rect 21312 6296 21328 6330
rect 21386 6296 21402 6330
rect 21470 6296 21486 6330
rect 21544 6296 21560 6330
rect 21628 6296 21644 6330
rect 21702 6296 21718 6330
rect 21786 6296 21802 6330
rect 21860 6296 21876 6330
rect 21944 6296 21960 6330
rect 22018 6296 22034 6330
rect 22102 6296 22118 6330
rect 22176 6296 22192 6330
rect 22260 6296 22276 6330
rect 22334 6296 22350 6330
rect 22418 6296 22434 6330
rect 22492 6296 22508 6330
rect 22576 6296 22592 6330
rect 22650 6296 22666 6330
rect 22734 6296 22750 6330
rect 22808 6296 22824 6330
rect 22892 6296 22908 6330
rect 22966 6296 22982 6330
rect 23050 6296 23066 6330
rect 23124 6296 23140 6330
rect 23208 6296 23224 6330
rect 23282 6296 23298 6330
rect 23366 6296 23382 6330
rect 23440 6296 23456 6330
rect 23524 6296 23540 6330
rect 23598 6296 23614 6330
rect 23682 6296 23698 6330
rect 23756 6296 23772 6330
rect 23840 6296 23856 6330
rect 23914 6296 23930 6330
rect 23998 6296 24014 6330
rect 24072 6296 24088 6330
rect 24156 6296 24172 6330
rect 24230 6296 24246 6330
rect 24314 6296 24330 6330
rect 24388 6296 24404 6330
rect 24472 6296 24488 6330
rect 24546 6296 24562 6330
rect 24630 6296 24646 6330
rect 24704 6296 24720 6330
rect 24788 6296 24804 6330
rect 24862 6296 24878 6330
rect 24946 6296 24962 6330
rect 25020 6296 25036 6330
rect 25104 6296 25120 6330
rect 25178 6296 25194 6330
rect 25262 6296 25278 6330
rect 25336 6296 25352 6330
rect 25420 6296 25436 6330
rect 25494 6296 25510 6330
rect 25578 6296 25594 6330
rect 25652 6296 25668 6330
rect 25736 6296 25752 6330
rect 25810 6296 25826 6330
rect 25894 6296 25910 6330
rect 182 6246 216 6262
rect 182 254 216 270
rect 340 6246 374 6262
rect 340 254 374 270
rect 498 6246 532 6262
rect 498 254 532 270
rect 656 6246 690 6262
rect 656 254 690 270
rect 814 6246 848 6262
rect 814 254 848 270
rect 972 6246 1006 6262
rect 972 254 1006 270
rect 1130 6246 1164 6262
rect 1130 254 1164 270
rect 1288 6246 1322 6262
rect 1288 254 1322 270
rect 1446 6246 1480 6262
rect 1446 254 1480 270
rect 1604 6246 1638 6262
rect 1604 254 1638 270
rect 1762 6246 1796 6262
rect 1762 254 1796 270
rect 1920 6246 1954 6262
rect 1920 254 1954 270
rect 2078 6246 2112 6262
rect 2078 254 2112 270
rect 2236 6246 2270 6262
rect 2236 254 2270 270
rect 2394 6246 2428 6262
rect 2394 254 2428 270
rect 2552 6246 2586 6262
rect 2552 254 2586 270
rect 2710 6246 2744 6262
rect 2710 254 2744 270
rect 2868 6246 2902 6262
rect 2868 254 2902 270
rect 3026 6246 3060 6262
rect 3026 254 3060 270
rect 3184 6246 3218 6262
rect 3184 254 3218 270
rect 3342 6246 3376 6262
rect 3342 254 3376 270
rect 3500 6246 3534 6262
rect 3500 254 3534 270
rect 3658 6246 3692 6262
rect 3658 254 3692 270
rect 3816 6246 3850 6262
rect 3816 254 3850 270
rect 3974 6246 4008 6262
rect 3974 254 4008 270
rect 4132 6246 4166 6262
rect 4132 254 4166 270
rect 4290 6246 4324 6262
rect 4290 254 4324 270
rect 4448 6246 4482 6262
rect 4448 254 4482 270
rect 4606 6246 4640 6262
rect 4606 254 4640 270
rect 4764 6246 4798 6262
rect 4764 254 4798 270
rect 4922 6246 4956 6262
rect 4922 254 4956 270
rect 7182 6246 7216 6262
rect 7182 254 7216 270
rect 7340 6246 7374 6262
rect 7340 254 7374 270
rect 7498 6246 7532 6262
rect 7498 254 7532 270
rect 7656 6246 7690 6262
rect 7656 254 7690 270
rect 7814 6246 7848 6262
rect 7814 254 7848 270
rect 7972 6246 8006 6262
rect 7972 254 8006 270
rect 8130 6246 8164 6262
rect 8130 254 8164 270
rect 8288 6246 8322 6262
rect 8288 254 8322 270
rect 8446 6246 8480 6262
rect 8446 254 8480 270
rect 8604 6246 8638 6262
rect 8604 254 8638 270
rect 8762 6246 8796 6262
rect 8762 254 8796 270
rect 8920 6246 8954 6262
rect 8920 254 8954 270
rect 9078 6246 9112 6262
rect 9078 254 9112 270
rect 9236 6246 9270 6262
rect 9236 254 9270 270
rect 9394 6246 9428 6262
rect 9394 254 9428 270
rect 9552 6246 9586 6262
rect 9552 254 9586 270
rect 9710 6246 9744 6262
rect 9710 254 9744 270
rect 9868 6246 9902 6262
rect 9868 254 9902 270
rect 10026 6246 10060 6262
rect 10026 254 10060 270
rect 10184 6246 10218 6262
rect 10184 254 10218 270
rect 10342 6246 10376 6262
rect 10342 254 10376 270
rect 10500 6246 10534 6262
rect 10500 254 10534 270
rect 10658 6246 10692 6262
rect 10658 254 10692 270
rect 10816 6246 10850 6262
rect 10816 254 10850 270
rect 10974 6246 11008 6262
rect 10974 254 11008 270
rect 11132 6246 11166 6262
rect 11132 254 11166 270
rect 11290 6246 11324 6262
rect 11290 254 11324 270
rect 11448 6246 11482 6262
rect 11448 254 11482 270
rect 11606 6246 11640 6262
rect 11606 254 11640 270
rect 11764 6246 11798 6262
rect 11764 254 11798 270
rect 11922 6246 11956 6262
rect 11922 254 11956 270
rect 14182 6246 14216 6262
rect 14182 254 14216 270
rect 14340 6246 14374 6262
rect 14340 254 14374 270
rect 14498 6246 14532 6262
rect 14498 254 14532 270
rect 14656 6246 14690 6262
rect 14656 254 14690 270
rect 14814 6246 14848 6262
rect 14814 254 14848 270
rect 14972 6246 15006 6262
rect 14972 254 15006 270
rect 15130 6246 15164 6262
rect 15130 254 15164 270
rect 15288 6246 15322 6262
rect 15288 254 15322 270
rect 15446 6246 15480 6262
rect 15446 254 15480 270
rect 15604 6246 15638 6262
rect 15604 254 15638 270
rect 15762 6246 15796 6262
rect 15762 254 15796 270
rect 15920 6246 15954 6262
rect 15920 254 15954 270
rect 16078 6246 16112 6262
rect 16078 254 16112 270
rect 16236 6246 16270 6262
rect 16236 254 16270 270
rect 16394 6246 16428 6262
rect 16394 254 16428 270
rect 16552 6246 16586 6262
rect 16552 254 16586 270
rect 16710 6246 16744 6262
rect 16710 254 16744 270
rect 16868 6246 16902 6262
rect 16868 254 16902 270
rect 17026 6246 17060 6262
rect 17026 254 17060 270
rect 17184 6246 17218 6262
rect 17184 254 17218 270
rect 17342 6246 17376 6262
rect 17342 254 17376 270
rect 17500 6246 17534 6262
rect 17500 254 17534 270
rect 17658 6246 17692 6262
rect 17658 254 17692 270
rect 17816 6246 17850 6262
rect 17816 254 17850 270
rect 17974 6246 18008 6262
rect 17974 254 18008 270
rect 18132 6246 18166 6262
rect 18132 254 18166 270
rect 18290 6246 18324 6262
rect 18290 254 18324 270
rect 18448 6246 18482 6262
rect 18448 254 18482 270
rect 18606 6246 18640 6262
rect 18606 254 18640 270
rect 18764 6246 18798 6262
rect 18764 254 18798 270
rect 18922 6246 18956 6262
rect 18922 254 18956 270
rect 21182 6246 21216 6262
rect 21182 254 21216 270
rect 21340 6246 21374 6262
rect 21340 254 21374 270
rect 21498 6246 21532 6262
rect 21498 254 21532 270
rect 21656 6246 21690 6262
rect 21656 254 21690 270
rect 21814 6246 21848 6262
rect 21814 254 21848 270
rect 21972 6246 22006 6262
rect 21972 254 22006 270
rect 22130 6246 22164 6262
rect 22130 254 22164 270
rect 22288 6246 22322 6262
rect 22288 254 22322 270
rect 22446 6246 22480 6262
rect 22446 254 22480 270
rect 22604 6246 22638 6262
rect 22604 254 22638 270
rect 22762 6246 22796 6262
rect 22762 254 22796 270
rect 22920 6246 22954 6262
rect 22920 254 22954 270
rect 23078 6246 23112 6262
rect 23078 254 23112 270
rect 23236 6246 23270 6262
rect 23236 254 23270 270
rect 23394 6246 23428 6262
rect 23394 254 23428 270
rect 23552 6246 23586 6262
rect 23552 254 23586 270
rect 23710 6246 23744 6262
rect 23710 254 23744 270
rect 23868 6246 23902 6262
rect 23868 254 23902 270
rect 24026 6246 24060 6262
rect 24026 254 24060 270
rect 24184 6246 24218 6262
rect 24184 254 24218 270
rect 24342 6246 24376 6262
rect 24342 254 24376 270
rect 24500 6246 24534 6262
rect 24500 254 24534 270
rect 24658 6246 24692 6262
rect 24658 254 24692 270
rect 24816 6246 24850 6262
rect 24816 254 24850 270
rect 24974 6246 25008 6262
rect 24974 254 25008 270
rect 25132 6246 25166 6262
rect 25132 254 25166 270
rect 25290 6246 25324 6262
rect 25290 254 25324 270
rect 25448 6246 25482 6262
rect 25448 254 25482 270
rect 25606 6246 25640 6262
rect 25606 254 25640 270
rect 25764 6246 25798 6262
rect 25764 254 25798 270
rect 25922 6246 25956 6262
rect 25922 254 25956 270
rect 228 186 244 220
rect 312 186 328 220
rect 386 186 402 220
rect 470 186 486 220
rect 544 186 560 220
rect 628 186 644 220
rect 702 186 718 220
rect 786 186 802 220
rect 860 186 876 220
rect 944 186 960 220
rect 1018 186 1034 220
rect 1102 186 1118 220
rect 1176 186 1192 220
rect 1260 186 1276 220
rect 1334 186 1350 220
rect 1418 186 1434 220
rect 1492 186 1508 220
rect 1576 186 1592 220
rect 1650 186 1666 220
rect 1734 186 1750 220
rect 1808 186 1824 220
rect 1892 186 1908 220
rect 1966 186 1982 220
rect 2050 186 2066 220
rect 2124 186 2140 220
rect 2208 186 2224 220
rect 2282 186 2298 220
rect 2366 186 2382 220
rect 2440 186 2456 220
rect 2524 186 2540 220
rect 2598 186 2614 220
rect 2682 186 2698 220
rect 2756 186 2772 220
rect 2840 186 2856 220
rect 2914 186 2930 220
rect 2998 186 3014 220
rect 3072 186 3088 220
rect 3156 186 3172 220
rect 3230 186 3246 220
rect 3314 186 3330 220
rect 3388 186 3404 220
rect 3472 186 3488 220
rect 3546 186 3562 220
rect 3630 186 3646 220
rect 3704 186 3720 220
rect 3788 186 3804 220
rect 3862 186 3878 220
rect 3946 186 3962 220
rect 4020 186 4036 220
rect 4104 186 4120 220
rect 4178 186 4194 220
rect 4262 186 4278 220
rect 4336 186 4352 220
rect 4420 186 4436 220
rect 4494 186 4510 220
rect 4578 186 4594 220
rect 4652 186 4668 220
rect 4736 186 4752 220
rect 4810 186 4826 220
rect 4894 186 4910 220
rect 48 82 82 144
rect 5056 82 5090 144
rect 48 48 144 82
rect 4994 48 5090 82
rect 7228 186 7244 220
rect 7312 186 7328 220
rect 7386 186 7402 220
rect 7470 186 7486 220
rect 7544 186 7560 220
rect 7628 186 7644 220
rect 7702 186 7718 220
rect 7786 186 7802 220
rect 7860 186 7876 220
rect 7944 186 7960 220
rect 8018 186 8034 220
rect 8102 186 8118 220
rect 8176 186 8192 220
rect 8260 186 8276 220
rect 8334 186 8350 220
rect 8418 186 8434 220
rect 8492 186 8508 220
rect 8576 186 8592 220
rect 8650 186 8666 220
rect 8734 186 8750 220
rect 8808 186 8824 220
rect 8892 186 8908 220
rect 8966 186 8982 220
rect 9050 186 9066 220
rect 9124 186 9140 220
rect 9208 186 9224 220
rect 9282 186 9298 220
rect 9366 186 9382 220
rect 9440 186 9456 220
rect 9524 186 9540 220
rect 9598 186 9614 220
rect 9682 186 9698 220
rect 9756 186 9772 220
rect 9840 186 9856 220
rect 9914 186 9930 220
rect 9998 186 10014 220
rect 10072 186 10088 220
rect 10156 186 10172 220
rect 10230 186 10246 220
rect 10314 186 10330 220
rect 10388 186 10404 220
rect 10472 186 10488 220
rect 10546 186 10562 220
rect 10630 186 10646 220
rect 10704 186 10720 220
rect 10788 186 10804 220
rect 10862 186 10878 220
rect 10946 186 10962 220
rect 11020 186 11036 220
rect 11104 186 11120 220
rect 11178 186 11194 220
rect 11262 186 11278 220
rect 11336 186 11352 220
rect 11420 186 11436 220
rect 11494 186 11510 220
rect 11578 186 11594 220
rect 11652 186 11668 220
rect 11736 186 11752 220
rect 11810 186 11826 220
rect 11894 186 11910 220
rect 7048 82 7082 144
rect 12056 82 12090 144
rect 7048 48 7144 82
rect 11994 48 12090 82
rect 14228 186 14244 220
rect 14312 186 14328 220
rect 14386 186 14402 220
rect 14470 186 14486 220
rect 14544 186 14560 220
rect 14628 186 14644 220
rect 14702 186 14718 220
rect 14786 186 14802 220
rect 14860 186 14876 220
rect 14944 186 14960 220
rect 15018 186 15034 220
rect 15102 186 15118 220
rect 15176 186 15192 220
rect 15260 186 15276 220
rect 15334 186 15350 220
rect 15418 186 15434 220
rect 15492 186 15508 220
rect 15576 186 15592 220
rect 15650 186 15666 220
rect 15734 186 15750 220
rect 15808 186 15824 220
rect 15892 186 15908 220
rect 15966 186 15982 220
rect 16050 186 16066 220
rect 16124 186 16140 220
rect 16208 186 16224 220
rect 16282 186 16298 220
rect 16366 186 16382 220
rect 16440 186 16456 220
rect 16524 186 16540 220
rect 16598 186 16614 220
rect 16682 186 16698 220
rect 16756 186 16772 220
rect 16840 186 16856 220
rect 16914 186 16930 220
rect 16998 186 17014 220
rect 17072 186 17088 220
rect 17156 186 17172 220
rect 17230 186 17246 220
rect 17314 186 17330 220
rect 17388 186 17404 220
rect 17472 186 17488 220
rect 17546 186 17562 220
rect 17630 186 17646 220
rect 17704 186 17720 220
rect 17788 186 17804 220
rect 17862 186 17878 220
rect 17946 186 17962 220
rect 18020 186 18036 220
rect 18104 186 18120 220
rect 18178 186 18194 220
rect 18262 186 18278 220
rect 18336 186 18352 220
rect 18420 186 18436 220
rect 18494 186 18510 220
rect 18578 186 18594 220
rect 18652 186 18668 220
rect 18736 186 18752 220
rect 18810 186 18826 220
rect 18894 186 18910 220
rect 14048 82 14082 144
rect 19056 82 19090 144
rect 14048 48 14144 82
rect 18994 48 19090 82
rect 21228 186 21244 220
rect 21312 186 21328 220
rect 21386 186 21402 220
rect 21470 186 21486 220
rect 21544 186 21560 220
rect 21628 186 21644 220
rect 21702 186 21718 220
rect 21786 186 21802 220
rect 21860 186 21876 220
rect 21944 186 21960 220
rect 22018 186 22034 220
rect 22102 186 22118 220
rect 22176 186 22192 220
rect 22260 186 22276 220
rect 22334 186 22350 220
rect 22418 186 22434 220
rect 22492 186 22508 220
rect 22576 186 22592 220
rect 22650 186 22666 220
rect 22734 186 22750 220
rect 22808 186 22824 220
rect 22892 186 22908 220
rect 22966 186 22982 220
rect 23050 186 23066 220
rect 23124 186 23140 220
rect 23208 186 23224 220
rect 23282 186 23298 220
rect 23366 186 23382 220
rect 23440 186 23456 220
rect 23524 186 23540 220
rect 23598 186 23614 220
rect 23682 186 23698 220
rect 23756 186 23772 220
rect 23840 186 23856 220
rect 23914 186 23930 220
rect 23998 186 24014 220
rect 24072 186 24088 220
rect 24156 186 24172 220
rect 24230 186 24246 220
rect 24314 186 24330 220
rect 24388 186 24404 220
rect 24472 186 24488 220
rect 24546 186 24562 220
rect 24630 186 24646 220
rect 24704 186 24720 220
rect 24788 186 24804 220
rect 24862 186 24878 220
rect 24946 186 24962 220
rect 25020 186 25036 220
rect 25104 186 25120 220
rect 25178 186 25194 220
rect 25262 186 25278 220
rect 25336 186 25352 220
rect 25420 186 25436 220
rect 25494 186 25510 220
rect 25578 186 25594 220
rect 25652 186 25668 220
rect 25736 186 25752 220
rect 25810 186 25826 220
rect 25894 186 25910 220
rect 21048 82 21082 144
rect 26056 82 26090 144
rect 21048 48 21144 82
rect 25994 48 26090 82
rect 48 -566 144 -532
rect 4994 -566 5090 -532
rect 48 -628 82 -566
rect 5056 -628 5090 -566
rect 228 -704 244 -670
rect 312 -704 328 -670
rect 386 -704 402 -670
rect 470 -704 486 -670
rect 544 -704 560 -670
rect 628 -704 644 -670
rect 702 -704 718 -670
rect 786 -704 802 -670
rect 860 -704 876 -670
rect 944 -704 960 -670
rect 1018 -704 1034 -670
rect 1102 -704 1118 -670
rect 1176 -704 1192 -670
rect 1260 -704 1276 -670
rect 1334 -704 1350 -670
rect 1418 -704 1434 -670
rect 1492 -704 1508 -670
rect 1576 -704 1592 -670
rect 1650 -704 1666 -670
rect 1734 -704 1750 -670
rect 1808 -704 1824 -670
rect 1892 -704 1908 -670
rect 1966 -704 1982 -670
rect 2050 -704 2066 -670
rect 2124 -704 2140 -670
rect 2208 -704 2224 -670
rect 2282 -704 2298 -670
rect 2366 -704 2382 -670
rect 2440 -704 2456 -670
rect 2524 -704 2540 -670
rect 2598 -704 2614 -670
rect 2682 -704 2698 -670
rect 2756 -704 2772 -670
rect 2840 -704 2856 -670
rect 2914 -704 2930 -670
rect 2998 -704 3014 -670
rect 3072 -704 3088 -670
rect 3156 -704 3172 -670
rect 3230 -704 3246 -670
rect 3314 -704 3330 -670
rect 3388 -704 3404 -670
rect 3472 -704 3488 -670
rect 3546 -704 3562 -670
rect 3630 -704 3646 -670
rect 3704 -704 3720 -670
rect 3788 -704 3804 -670
rect 3862 -704 3878 -670
rect 3946 -704 3962 -670
rect 4020 -704 4036 -670
rect 4104 -704 4120 -670
rect 4178 -704 4194 -670
rect 4262 -704 4278 -670
rect 4336 -704 4352 -670
rect 4420 -704 4436 -670
rect 4494 -704 4510 -670
rect 4578 -704 4594 -670
rect 4652 -704 4668 -670
rect 4736 -704 4752 -670
rect 4810 -704 4826 -670
rect 4894 -704 4910 -670
rect 7048 -566 7144 -532
rect 11994 -566 12090 -532
rect 7048 -628 7082 -566
rect 12056 -628 12090 -566
rect 7228 -704 7244 -670
rect 7312 -704 7328 -670
rect 7386 -704 7402 -670
rect 7470 -704 7486 -670
rect 7544 -704 7560 -670
rect 7628 -704 7644 -670
rect 7702 -704 7718 -670
rect 7786 -704 7802 -670
rect 7860 -704 7876 -670
rect 7944 -704 7960 -670
rect 8018 -704 8034 -670
rect 8102 -704 8118 -670
rect 8176 -704 8192 -670
rect 8260 -704 8276 -670
rect 8334 -704 8350 -670
rect 8418 -704 8434 -670
rect 8492 -704 8508 -670
rect 8576 -704 8592 -670
rect 8650 -704 8666 -670
rect 8734 -704 8750 -670
rect 8808 -704 8824 -670
rect 8892 -704 8908 -670
rect 8966 -704 8982 -670
rect 9050 -704 9066 -670
rect 9124 -704 9140 -670
rect 9208 -704 9224 -670
rect 9282 -704 9298 -670
rect 9366 -704 9382 -670
rect 9440 -704 9456 -670
rect 9524 -704 9540 -670
rect 9598 -704 9614 -670
rect 9682 -704 9698 -670
rect 9756 -704 9772 -670
rect 9840 -704 9856 -670
rect 9914 -704 9930 -670
rect 9998 -704 10014 -670
rect 10072 -704 10088 -670
rect 10156 -704 10172 -670
rect 10230 -704 10246 -670
rect 10314 -704 10330 -670
rect 10388 -704 10404 -670
rect 10472 -704 10488 -670
rect 10546 -704 10562 -670
rect 10630 -704 10646 -670
rect 10704 -704 10720 -670
rect 10788 -704 10804 -670
rect 10862 -704 10878 -670
rect 10946 -704 10962 -670
rect 11020 -704 11036 -670
rect 11104 -704 11120 -670
rect 11178 -704 11194 -670
rect 11262 -704 11278 -670
rect 11336 -704 11352 -670
rect 11420 -704 11436 -670
rect 11494 -704 11510 -670
rect 11578 -704 11594 -670
rect 11652 -704 11668 -670
rect 11736 -704 11752 -670
rect 11810 -704 11826 -670
rect 11894 -704 11910 -670
rect 14048 -566 14144 -532
rect 18994 -566 19090 -532
rect 14048 -628 14082 -566
rect 19056 -628 19090 -566
rect 14228 -704 14244 -670
rect 14312 -704 14328 -670
rect 14386 -704 14402 -670
rect 14470 -704 14486 -670
rect 14544 -704 14560 -670
rect 14628 -704 14644 -670
rect 14702 -704 14718 -670
rect 14786 -704 14802 -670
rect 14860 -704 14876 -670
rect 14944 -704 14960 -670
rect 15018 -704 15034 -670
rect 15102 -704 15118 -670
rect 15176 -704 15192 -670
rect 15260 -704 15276 -670
rect 15334 -704 15350 -670
rect 15418 -704 15434 -670
rect 15492 -704 15508 -670
rect 15576 -704 15592 -670
rect 15650 -704 15666 -670
rect 15734 -704 15750 -670
rect 15808 -704 15824 -670
rect 15892 -704 15908 -670
rect 15966 -704 15982 -670
rect 16050 -704 16066 -670
rect 16124 -704 16140 -670
rect 16208 -704 16224 -670
rect 16282 -704 16298 -670
rect 16366 -704 16382 -670
rect 16440 -704 16456 -670
rect 16524 -704 16540 -670
rect 16598 -704 16614 -670
rect 16682 -704 16698 -670
rect 16756 -704 16772 -670
rect 16840 -704 16856 -670
rect 16914 -704 16930 -670
rect 16998 -704 17014 -670
rect 17072 -704 17088 -670
rect 17156 -704 17172 -670
rect 17230 -704 17246 -670
rect 17314 -704 17330 -670
rect 17388 -704 17404 -670
rect 17472 -704 17488 -670
rect 17546 -704 17562 -670
rect 17630 -704 17646 -670
rect 17704 -704 17720 -670
rect 17788 -704 17804 -670
rect 17862 -704 17878 -670
rect 17946 -704 17962 -670
rect 18020 -704 18036 -670
rect 18104 -704 18120 -670
rect 18178 -704 18194 -670
rect 18262 -704 18278 -670
rect 18336 -704 18352 -670
rect 18420 -704 18436 -670
rect 18494 -704 18510 -670
rect 18578 -704 18594 -670
rect 18652 -704 18668 -670
rect 18736 -704 18752 -670
rect 18810 -704 18826 -670
rect 18894 -704 18910 -670
rect 21048 -566 21144 -532
rect 25994 -566 26090 -532
rect 21048 -628 21082 -566
rect 26056 -628 26090 -566
rect 21228 -704 21244 -670
rect 21312 -704 21328 -670
rect 21386 -704 21402 -670
rect 21470 -704 21486 -670
rect 21544 -704 21560 -670
rect 21628 -704 21644 -670
rect 21702 -704 21718 -670
rect 21786 -704 21802 -670
rect 21860 -704 21876 -670
rect 21944 -704 21960 -670
rect 22018 -704 22034 -670
rect 22102 -704 22118 -670
rect 22176 -704 22192 -670
rect 22260 -704 22276 -670
rect 22334 -704 22350 -670
rect 22418 -704 22434 -670
rect 22492 -704 22508 -670
rect 22576 -704 22592 -670
rect 22650 -704 22666 -670
rect 22734 -704 22750 -670
rect 22808 -704 22824 -670
rect 22892 -704 22908 -670
rect 22966 -704 22982 -670
rect 23050 -704 23066 -670
rect 23124 -704 23140 -670
rect 23208 -704 23224 -670
rect 23282 -704 23298 -670
rect 23366 -704 23382 -670
rect 23440 -704 23456 -670
rect 23524 -704 23540 -670
rect 23598 -704 23614 -670
rect 23682 -704 23698 -670
rect 23756 -704 23772 -670
rect 23840 -704 23856 -670
rect 23914 -704 23930 -670
rect 23998 -704 24014 -670
rect 24072 -704 24088 -670
rect 24156 -704 24172 -670
rect 24230 -704 24246 -670
rect 24314 -704 24330 -670
rect 24388 -704 24404 -670
rect 24472 -704 24488 -670
rect 24546 -704 24562 -670
rect 24630 -704 24646 -670
rect 24704 -704 24720 -670
rect 24788 -704 24804 -670
rect 24862 -704 24878 -670
rect 24946 -704 24962 -670
rect 25020 -704 25036 -670
rect 25104 -704 25120 -670
rect 25178 -704 25194 -670
rect 25262 -704 25278 -670
rect 25336 -704 25352 -670
rect 25420 -704 25436 -670
rect 25494 -704 25510 -670
rect 25578 -704 25594 -670
rect 25652 -704 25668 -670
rect 25736 -704 25752 -670
rect 25810 -704 25826 -670
rect 25894 -704 25910 -670
rect 182 -754 216 -738
rect 182 -6746 216 -6730
rect 340 -754 374 -738
rect 340 -6746 374 -6730
rect 498 -754 532 -738
rect 498 -6746 532 -6730
rect 656 -754 690 -738
rect 656 -6746 690 -6730
rect 814 -754 848 -738
rect 814 -6746 848 -6730
rect 972 -754 1006 -738
rect 972 -6746 1006 -6730
rect 1130 -754 1164 -738
rect 1130 -6746 1164 -6730
rect 1288 -754 1322 -738
rect 1288 -6746 1322 -6730
rect 1446 -754 1480 -738
rect 1446 -6746 1480 -6730
rect 1604 -754 1638 -738
rect 1604 -6746 1638 -6730
rect 1762 -754 1796 -738
rect 1762 -6746 1796 -6730
rect 1920 -754 1954 -738
rect 1920 -6746 1954 -6730
rect 2078 -754 2112 -738
rect 2078 -6746 2112 -6730
rect 2236 -754 2270 -738
rect 2236 -6746 2270 -6730
rect 2394 -754 2428 -738
rect 2394 -6746 2428 -6730
rect 2552 -754 2586 -738
rect 2552 -6746 2586 -6730
rect 2710 -754 2744 -738
rect 2710 -6746 2744 -6730
rect 2868 -754 2902 -738
rect 2868 -6746 2902 -6730
rect 3026 -754 3060 -738
rect 3026 -6746 3060 -6730
rect 3184 -754 3218 -738
rect 3184 -6746 3218 -6730
rect 3342 -754 3376 -738
rect 3342 -6746 3376 -6730
rect 3500 -754 3534 -738
rect 3500 -6746 3534 -6730
rect 3658 -754 3692 -738
rect 3658 -6746 3692 -6730
rect 3816 -754 3850 -738
rect 3816 -6746 3850 -6730
rect 3974 -754 4008 -738
rect 3974 -6746 4008 -6730
rect 4132 -754 4166 -738
rect 4132 -6746 4166 -6730
rect 4290 -754 4324 -738
rect 4290 -6746 4324 -6730
rect 4448 -754 4482 -738
rect 4448 -6746 4482 -6730
rect 4606 -754 4640 -738
rect 4606 -6746 4640 -6730
rect 4764 -754 4798 -738
rect 4764 -6746 4798 -6730
rect 4922 -754 4956 -738
rect 4922 -6746 4956 -6730
rect 7182 -754 7216 -738
rect 7182 -6746 7216 -6730
rect 7340 -754 7374 -738
rect 7340 -6746 7374 -6730
rect 7498 -754 7532 -738
rect 7498 -6746 7532 -6730
rect 7656 -754 7690 -738
rect 7656 -6746 7690 -6730
rect 7814 -754 7848 -738
rect 7814 -6746 7848 -6730
rect 7972 -754 8006 -738
rect 7972 -6746 8006 -6730
rect 8130 -754 8164 -738
rect 8130 -6746 8164 -6730
rect 8288 -754 8322 -738
rect 8288 -6746 8322 -6730
rect 8446 -754 8480 -738
rect 8446 -6746 8480 -6730
rect 8604 -754 8638 -738
rect 8604 -6746 8638 -6730
rect 8762 -754 8796 -738
rect 8762 -6746 8796 -6730
rect 8920 -754 8954 -738
rect 8920 -6746 8954 -6730
rect 9078 -754 9112 -738
rect 9078 -6746 9112 -6730
rect 9236 -754 9270 -738
rect 9236 -6746 9270 -6730
rect 9394 -754 9428 -738
rect 9394 -6746 9428 -6730
rect 9552 -754 9586 -738
rect 9552 -6746 9586 -6730
rect 9710 -754 9744 -738
rect 9710 -6746 9744 -6730
rect 9868 -754 9902 -738
rect 9868 -6746 9902 -6730
rect 10026 -754 10060 -738
rect 10026 -6746 10060 -6730
rect 10184 -754 10218 -738
rect 10184 -6746 10218 -6730
rect 10342 -754 10376 -738
rect 10342 -6746 10376 -6730
rect 10500 -754 10534 -738
rect 10500 -6746 10534 -6730
rect 10658 -754 10692 -738
rect 10658 -6746 10692 -6730
rect 10816 -754 10850 -738
rect 10816 -6746 10850 -6730
rect 10974 -754 11008 -738
rect 10974 -6746 11008 -6730
rect 11132 -754 11166 -738
rect 11132 -6746 11166 -6730
rect 11290 -754 11324 -738
rect 11290 -6746 11324 -6730
rect 11448 -754 11482 -738
rect 11448 -6746 11482 -6730
rect 11606 -754 11640 -738
rect 11606 -6746 11640 -6730
rect 11764 -754 11798 -738
rect 11764 -6746 11798 -6730
rect 11922 -754 11956 -738
rect 11922 -6746 11956 -6730
rect 14182 -754 14216 -738
rect 14182 -6746 14216 -6730
rect 14340 -754 14374 -738
rect 14340 -6746 14374 -6730
rect 14498 -754 14532 -738
rect 14498 -6746 14532 -6730
rect 14656 -754 14690 -738
rect 14656 -6746 14690 -6730
rect 14814 -754 14848 -738
rect 14814 -6746 14848 -6730
rect 14972 -754 15006 -738
rect 14972 -6746 15006 -6730
rect 15130 -754 15164 -738
rect 15130 -6746 15164 -6730
rect 15288 -754 15322 -738
rect 15288 -6746 15322 -6730
rect 15446 -754 15480 -738
rect 15446 -6746 15480 -6730
rect 15604 -754 15638 -738
rect 15604 -6746 15638 -6730
rect 15762 -754 15796 -738
rect 15762 -6746 15796 -6730
rect 15920 -754 15954 -738
rect 15920 -6746 15954 -6730
rect 16078 -754 16112 -738
rect 16078 -6746 16112 -6730
rect 16236 -754 16270 -738
rect 16236 -6746 16270 -6730
rect 16394 -754 16428 -738
rect 16394 -6746 16428 -6730
rect 16552 -754 16586 -738
rect 16552 -6746 16586 -6730
rect 16710 -754 16744 -738
rect 16710 -6746 16744 -6730
rect 16868 -754 16902 -738
rect 16868 -6746 16902 -6730
rect 17026 -754 17060 -738
rect 17026 -6746 17060 -6730
rect 17184 -754 17218 -738
rect 17184 -6746 17218 -6730
rect 17342 -754 17376 -738
rect 17342 -6746 17376 -6730
rect 17500 -754 17534 -738
rect 17500 -6746 17534 -6730
rect 17658 -754 17692 -738
rect 17658 -6746 17692 -6730
rect 17816 -754 17850 -738
rect 17816 -6746 17850 -6730
rect 17974 -754 18008 -738
rect 17974 -6746 18008 -6730
rect 18132 -754 18166 -738
rect 18132 -6746 18166 -6730
rect 18290 -754 18324 -738
rect 18290 -6746 18324 -6730
rect 18448 -754 18482 -738
rect 18448 -6746 18482 -6730
rect 18606 -754 18640 -738
rect 18606 -6746 18640 -6730
rect 18764 -754 18798 -738
rect 18764 -6746 18798 -6730
rect 18922 -754 18956 -738
rect 18922 -6746 18956 -6730
rect 21182 -754 21216 -738
rect 21182 -6746 21216 -6730
rect 21340 -754 21374 -738
rect 21340 -6746 21374 -6730
rect 21498 -754 21532 -738
rect 21498 -6746 21532 -6730
rect 21656 -754 21690 -738
rect 21656 -6746 21690 -6730
rect 21814 -754 21848 -738
rect 21814 -6746 21848 -6730
rect 21972 -754 22006 -738
rect 21972 -6746 22006 -6730
rect 22130 -754 22164 -738
rect 22130 -6746 22164 -6730
rect 22288 -754 22322 -738
rect 22288 -6746 22322 -6730
rect 22446 -754 22480 -738
rect 22446 -6746 22480 -6730
rect 22604 -754 22638 -738
rect 22604 -6746 22638 -6730
rect 22762 -754 22796 -738
rect 22762 -6746 22796 -6730
rect 22920 -754 22954 -738
rect 22920 -6746 22954 -6730
rect 23078 -754 23112 -738
rect 23078 -6746 23112 -6730
rect 23236 -754 23270 -738
rect 23236 -6746 23270 -6730
rect 23394 -754 23428 -738
rect 23394 -6746 23428 -6730
rect 23552 -754 23586 -738
rect 23552 -6746 23586 -6730
rect 23710 -754 23744 -738
rect 23710 -6746 23744 -6730
rect 23868 -754 23902 -738
rect 23868 -6746 23902 -6730
rect 24026 -754 24060 -738
rect 24026 -6746 24060 -6730
rect 24184 -754 24218 -738
rect 24184 -6746 24218 -6730
rect 24342 -754 24376 -738
rect 24342 -6746 24376 -6730
rect 24500 -754 24534 -738
rect 24500 -6746 24534 -6730
rect 24658 -754 24692 -738
rect 24658 -6746 24692 -6730
rect 24816 -754 24850 -738
rect 24816 -6746 24850 -6730
rect 24974 -754 25008 -738
rect 24974 -6746 25008 -6730
rect 25132 -754 25166 -738
rect 25132 -6746 25166 -6730
rect 25290 -754 25324 -738
rect 25290 -6746 25324 -6730
rect 25448 -754 25482 -738
rect 25448 -6746 25482 -6730
rect 25606 -754 25640 -738
rect 25606 -6746 25640 -6730
rect 25764 -754 25798 -738
rect 25764 -6746 25798 -6730
rect 25922 -754 25956 -738
rect 25922 -6746 25956 -6730
rect 228 -6814 244 -6780
rect 312 -6814 328 -6780
rect 386 -6814 402 -6780
rect 470 -6814 486 -6780
rect 544 -6814 560 -6780
rect 628 -6814 644 -6780
rect 702 -6814 718 -6780
rect 786 -6814 802 -6780
rect 860 -6814 876 -6780
rect 944 -6814 960 -6780
rect 1018 -6814 1034 -6780
rect 1102 -6814 1118 -6780
rect 1176 -6814 1192 -6780
rect 1260 -6814 1276 -6780
rect 1334 -6814 1350 -6780
rect 1418 -6814 1434 -6780
rect 1492 -6814 1508 -6780
rect 1576 -6814 1592 -6780
rect 1650 -6814 1666 -6780
rect 1734 -6814 1750 -6780
rect 1808 -6814 1824 -6780
rect 1892 -6814 1908 -6780
rect 1966 -6814 1982 -6780
rect 2050 -6814 2066 -6780
rect 2124 -6814 2140 -6780
rect 2208 -6814 2224 -6780
rect 2282 -6814 2298 -6780
rect 2366 -6814 2382 -6780
rect 2440 -6814 2456 -6780
rect 2524 -6814 2540 -6780
rect 2598 -6814 2614 -6780
rect 2682 -6814 2698 -6780
rect 2756 -6814 2772 -6780
rect 2840 -6814 2856 -6780
rect 2914 -6814 2930 -6780
rect 2998 -6814 3014 -6780
rect 3072 -6814 3088 -6780
rect 3156 -6814 3172 -6780
rect 3230 -6814 3246 -6780
rect 3314 -6814 3330 -6780
rect 3388 -6814 3404 -6780
rect 3472 -6814 3488 -6780
rect 3546 -6814 3562 -6780
rect 3630 -6814 3646 -6780
rect 3704 -6814 3720 -6780
rect 3788 -6814 3804 -6780
rect 3862 -6814 3878 -6780
rect 3946 -6814 3962 -6780
rect 4020 -6814 4036 -6780
rect 4104 -6814 4120 -6780
rect 4178 -6814 4194 -6780
rect 4262 -6814 4278 -6780
rect 4336 -6814 4352 -6780
rect 4420 -6814 4436 -6780
rect 4494 -6814 4510 -6780
rect 4578 -6814 4594 -6780
rect 4652 -6814 4668 -6780
rect 4736 -6814 4752 -6780
rect 4810 -6814 4826 -6780
rect 4894 -6814 4910 -6780
rect 48 -6918 82 -6856
rect 5056 -6918 5090 -6856
rect 48 -6952 144 -6918
rect 4994 -6952 5090 -6918
rect 7228 -6814 7244 -6780
rect 7312 -6814 7328 -6780
rect 7386 -6814 7402 -6780
rect 7470 -6814 7486 -6780
rect 7544 -6814 7560 -6780
rect 7628 -6814 7644 -6780
rect 7702 -6814 7718 -6780
rect 7786 -6814 7802 -6780
rect 7860 -6814 7876 -6780
rect 7944 -6814 7960 -6780
rect 8018 -6814 8034 -6780
rect 8102 -6814 8118 -6780
rect 8176 -6814 8192 -6780
rect 8260 -6814 8276 -6780
rect 8334 -6814 8350 -6780
rect 8418 -6814 8434 -6780
rect 8492 -6814 8508 -6780
rect 8576 -6814 8592 -6780
rect 8650 -6814 8666 -6780
rect 8734 -6814 8750 -6780
rect 8808 -6814 8824 -6780
rect 8892 -6814 8908 -6780
rect 8966 -6814 8982 -6780
rect 9050 -6814 9066 -6780
rect 9124 -6814 9140 -6780
rect 9208 -6814 9224 -6780
rect 9282 -6814 9298 -6780
rect 9366 -6814 9382 -6780
rect 9440 -6814 9456 -6780
rect 9524 -6814 9540 -6780
rect 9598 -6814 9614 -6780
rect 9682 -6814 9698 -6780
rect 9756 -6814 9772 -6780
rect 9840 -6814 9856 -6780
rect 9914 -6814 9930 -6780
rect 9998 -6814 10014 -6780
rect 10072 -6814 10088 -6780
rect 10156 -6814 10172 -6780
rect 10230 -6814 10246 -6780
rect 10314 -6814 10330 -6780
rect 10388 -6814 10404 -6780
rect 10472 -6814 10488 -6780
rect 10546 -6814 10562 -6780
rect 10630 -6814 10646 -6780
rect 10704 -6814 10720 -6780
rect 10788 -6814 10804 -6780
rect 10862 -6814 10878 -6780
rect 10946 -6814 10962 -6780
rect 11020 -6814 11036 -6780
rect 11104 -6814 11120 -6780
rect 11178 -6814 11194 -6780
rect 11262 -6814 11278 -6780
rect 11336 -6814 11352 -6780
rect 11420 -6814 11436 -6780
rect 11494 -6814 11510 -6780
rect 11578 -6814 11594 -6780
rect 11652 -6814 11668 -6780
rect 11736 -6814 11752 -6780
rect 11810 -6814 11826 -6780
rect 11894 -6814 11910 -6780
rect 7048 -6918 7082 -6856
rect 12056 -6918 12090 -6856
rect 7048 -6952 7144 -6918
rect 11994 -6952 12090 -6918
rect 14228 -6814 14244 -6780
rect 14312 -6814 14328 -6780
rect 14386 -6814 14402 -6780
rect 14470 -6814 14486 -6780
rect 14544 -6814 14560 -6780
rect 14628 -6814 14644 -6780
rect 14702 -6814 14718 -6780
rect 14786 -6814 14802 -6780
rect 14860 -6814 14876 -6780
rect 14944 -6814 14960 -6780
rect 15018 -6814 15034 -6780
rect 15102 -6814 15118 -6780
rect 15176 -6814 15192 -6780
rect 15260 -6814 15276 -6780
rect 15334 -6814 15350 -6780
rect 15418 -6814 15434 -6780
rect 15492 -6814 15508 -6780
rect 15576 -6814 15592 -6780
rect 15650 -6814 15666 -6780
rect 15734 -6814 15750 -6780
rect 15808 -6814 15824 -6780
rect 15892 -6814 15908 -6780
rect 15966 -6814 15982 -6780
rect 16050 -6814 16066 -6780
rect 16124 -6814 16140 -6780
rect 16208 -6814 16224 -6780
rect 16282 -6814 16298 -6780
rect 16366 -6814 16382 -6780
rect 16440 -6814 16456 -6780
rect 16524 -6814 16540 -6780
rect 16598 -6814 16614 -6780
rect 16682 -6814 16698 -6780
rect 16756 -6814 16772 -6780
rect 16840 -6814 16856 -6780
rect 16914 -6814 16930 -6780
rect 16998 -6814 17014 -6780
rect 17072 -6814 17088 -6780
rect 17156 -6814 17172 -6780
rect 17230 -6814 17246 -6780
rect 17314 -6814 17330 -6780
rect 17388 -6814 17404 -6780
rect 17472 -6814 17488 -6780
rect 17546 -6814 17562 -6780
rect 17630 -6814 17646 -6780
rect 17704 -6814 17720 -6780
rect 17788 -6814 17804 -6780
rect 17862 -6814 17878 -6780
rect 17946 -6814 17962 -6780
rect 18020 -6814 18036 -6780
rect 18104 -6814 18120 -6780
rect 18178 -6814 18194 -6780
rect 18262 -6814 18278 -6780
rect 18336 -6814 18352 -6780
rect 18420 -6814 18436 -6780
rect 18494 -6814 18510 -6780
rect 18578 -6814 18594 -6780
rect 18652 -6814 18668 -6780
rect 18736 -6814 18752 -6780
rect 18810 -6814 18826 -6780
rect 18894 -6814 18910 -6780
rect 14048 -6918 14082 -6856
rect 19056 -6918 19090 -6856
rect 14048 -6952 14144 -6918
rect 18994 -6952 19090 -6918
rect 21228 -6814 21244 -6780
rect 21312 -6814 21328 -6780
rect 21386 -6814 21402 -6780
rect 21470 -6814 21486 -6780
rect 21544 -6814 21560 -6780
rect 21628 -6814 21644 -6780
rect 21702 -6814 21718 -6780
rect 21786 -6814 21802 -6780
rect 21860 -6814 21876 -6780
rect 21944 -6814 21960 -6780
rect 22018 -6814 22034 -6780
rect 22102 -6814 22118 -6780
rect 22176 -6814 22192 -6780
rect 22260 -6814 22276 -6780
rect 22334 -6814 22350 -6780
rect 22418 -6814 22434 -6780
rect 22492 -6814 22508 -6780
rect 22576 -6814 22592 -6780
rect 22650 -6814 22666 -6780
rect 22734 -6814 22750 -6780
rect 22808 -6814 22824 -6780
rect 22892 -6814 22908 -6780
rect 22966 -6814 22982 -6780
rect 23050 -6814 23066 -6780
rect 23124 -6814 23140 -6780
rect 23208 -6814 23224 -6780
rect 23282 -6814 23298 -6780
rect 23366 -6814 23382 -6780
rect 23440 -6814 23456 -6780
rect 23524 -6814 23540 -6780
rect 23598 -6814 23614 -6780
rect 23682 -6814 23698 -6780
rect 23756 -6814 23772 -6780
rect 23840 -6814 23856 -6780
rect 23914 -6814 23930 -6780
rect 23998 -6814 24014 -6780
rect 24072 -6814 24088 -6780
rect 24156 -6814 24172 -6780
rect 24230 -6814 24246 -6780
rect 24314 -6814 24330 -6780
rect 24388 -6814 24404 -6780
rect 24472 -6814 24488 -6780
rect 24546 -6814 24562 -6780
rect 24630 -6814 24646 -6780
rect 24704 -6814 24720 -6780
rect 24788 -6814 24804 -6780
rect 24862 -6814 24878 -6780
rect 24946 -6814 24962 -6780
rect 25020 -6814 25036 -6780
rect 25104 -6814 25120 -6780
rect 25178 -6814 25194 -6780
rect 25262 -6814 25278 -6780
rect 25336 -6814 25352 -6780
rect 25420 -6814 25436 -6780
rect 25494 -6814 25510 -6780
rect 25578 -6814 25594 -6780
rect 25652 -6814 25668 -6780
rect 25736 -6814 25752 -6780
rect 25810 -6814 25826 -6780
rect 25894 -6814 25910 -6780
rect 21048 -6918 21082 -6856
rect 26056 -6918 26090 -6856
rect 21048 -6952 21144 -6918
rect 25994 -6952 26090 -6918
<< viali >>
rect 236 6468 4959 6470
rect 7236 6468 11959 6470
rect 14236 6468 18959 6470
rect 21236 6468 25959 6470
rect 236 6434 4959 6468
rect 236 6432 4959 6434
rect 244 6296 312 6330
rect 402 6296 470 6330
rect 560 6296 628 6330
rect 718 6296 786 6330
rect 876 6296 944 6330
rect 1034 6296 1102 6330
rect 1192 6296 1260 6330
rect 1350 6296 1418 6330
rect 1508 6296 1576 6330
rect 1666 6296 1734 6330
rect 1824 6296 1892 6330
rect 1982 6296 2050 6330
rect 2140 6296 2208 6330
rect 2298 6296 2366 6330
rect 2456 6296 2524 6330
rect 2614 6296 2682 6330
rect 2772 6296 2840 6330
rect 2930 6296 2998 6330
rect 3088 6296 3156 6330
rect 3246 6296 3314 6330
rect 3404 6296 3472 6330
rect 3562 6296 3630 6330
rect 3720 6296 3788 6330
rect 3878 6296 3946 6330
rect 4036 6296 4104 6330
rect 4194 6296 4262 6330
rect 4352 6296 4420 6330
rect 4510 6296 4578 6330
rect 4668 6296 4736 6330
rect 4826 6296 4894 6330
rect 7236 6434 11959 6468
rect 7236 6432 11959 6434
rect 7244 6296 7312 6330
rect 7402 6296 7470 6330
rect 7560 6296 7628 6330
rect 7718 6296 7786 6330
rect 7876 6296 7944 6330
rect 8034 6296 8102 6330
rect 8192 6296 8260 6330
rect 8350 6296 8418 6330
rect 8508 6296 8576 6330
rect 8666 6296 8734 6330
rect 8824 6296 8892 6330
rect 8982 6296 9050 6330
rect 9140 6296 9208 6330
rect 9298 6296 9366 6330
rect 9456 6296 9524 6330
rect 9614 6296 9682 6330
rect 9772 6296 9840 6330
rect 9930 6296 9998 6330
rect 10088 6296 10156 6330
rect 10246 6296 10314 6330
rect 10404 6296 10472 6330
rect 10562 6296 10630 6330
rect 10720 6296 10788 6330
rect 10878 6296 10946 6330
rect 11036 6296 11104 6330
rect 11194 6296 11262 6330
rect 11352 6296 11420 6330
rect 11510 6296 11578 6330
rect 11668 6296 11736 6330
rect 11826 6296 11894 6330
rect 14236 6434 18959 6468
rect 14236 6432 18959 6434
rect 14244 6296 14312 6330
rect 14402 6296 14470 6330
rect 14560 6296 14628 6330
rect 14718 6296 14786 6330
rect 14876 6296 14944 6330
rect 15034 6296 15102 6330
rect 15192 6296 15260 6330
rect 15350 6296 15418 6330
rect 15508 6296 15576 6330
rect 15666 6296 15734 6330
rect 15824 6296 15892 6330
rect 15982 6296 16050 6330
rect 16140 6296 16208 6330
rect 16298 6296 16366 6330
rect 16456 6296 16524 6330
rect 16614 6296 16682 6330
rect 16772 6296 16840 6330
rect 16930 6296 16998 6330
rect 17088 6296 17156 6330
rect 17246 6296 17314 6330
rect 17404 6296 17472 6330
rect 17562 6296 17630 6330
rect 17720 6296 17788 6330
rect 17878 6296 17946 6330
rect 18036 6296 18104 6330
rect 18194 6296 18262 6330
rect 18352 6296 18420 6330
rect 18510 6296 18578 6330
rect 18668 6296 18736 6330
rect 18826 6296 18894 6330
rect 21236 6434 25959 6468
rect 21236 6432 25959 6434
rect 21244 6296 21312 6330
rect 21402 6296 21470 6330
rect 21560 6296 21628 6330
rect 21718 6296 21786 6330
rect 21876 6296 21944 6330
rect 22034 6296 22102 6330
rect 22192 6296 22260 6330
rect 22350 6296 22418 6330
rect 22508 6296 22576 6330
rect 22666 6296 22734 6330
rect 22824 6296 22892 6330
rect 22982 6296 23050 6330
rect 23140 6296 23208 6330
rect 23298 6296 23366 6330
rect 23456 6296 23524 6330
rect 23614 6296 23682 6330
rect 23772 6296 23840 6330
rect 23930 6296 23998 6330
rect 24088 6296 24156 6330
rect 24246 6296 24314 6330
rect 24404 6296 24472 6330
rect 24562 6296 24630 6330
rect 24720 6296 24788 6330
rect 24878 6296 24946 6330
rect 25036 6296 25104 6330
rect 25194 6296 25262 6330
rect 25352 6296 25420 6330
rect 25510 6296 25578 6330
rect 25668 6296 25736 6330
rect 25826 6296 25894 6330
rect 46 236 48 6280
rect 48 236 82 6280
rect 82 236 84 6280
rect 182 270 216 6246
rect 340 270 374 6246
rect 498 270 532 6246
rect 656 270 690 6246
rect 814 270 848 6246
rect 972 270 1006 6246
rect 1130 270 1164 6246
rect 1288 270 1322 6246
rect 1446 270 1480 6246
rect 1604 270 1638 6246
rect 1762 270 1796 6246
rect 1920 270 1954 6246
rect 2078 270 2112 6246
rect 2236 270 2270 6246
rect 2394 270 2428 6246
rect 2552 270 2586 6246
rect 2710 270 2744 6246
rect 2868 270 2902 6246
rect 3026 270 3060 6246
rect 3184 270 3218 6246
rect 3342 270 3376 6246
rect 3500 270 3534 6246
rect 3658 270 3692 6246
rect 3816 270 3850 6246
rect 3974 270 4008 6246
rect 4132 270 4166 6246
rect 4290 270 4324 6246
rect 4448 270 4482 6246
rect 4606 270 4640 6246
rect 4764 270 4798 6246
rect 4922 270 4956 6246
rect 5054 236 5056 6280
rect 5056 236 5090 6280
rect 5090 236 5092 6280
rect 7046 236 7048 6280
rect 7048 236 7082 6280
rect 7082 236 7084 6280
rect 7182 270 7216 6246
rect 7340 270 7374 6246
rect 7498 270 7532 6246
rect 7656 270 7690 6246
rect 7814 270 7848 6246
rect 7972 270 8006 6246
rect 8130 270 8164 6246
rect 8288 270 8322 6246
rect 8446 270 8480 6246
rect 8604 270 8638 6246
rect 8762 270 8796 6246
rect 8920 270 8954 6246
rect 9078 270 9112 6246
rect 9236 270 9270 6246
rect 9394 270 9428 6246
rect 9552 270 9586 6246
rect 9710 270 9744 6246
rect 9868 270 9902 6246
rect 10026 270 10060 6246
rect 10184 270 10218 6246
rect 10342 270 10376 6246
rect 10500 270 10534 6246
rect 10658 270 10692 6246
rect 10816 270 10850 6246
rect 10974 270 11008 6246
rect 11132 270 11166 6246
rect 11290 270 11324 6246
rect 11448 270 11482 6246
rect 11606 270 11640 6246
rect 11764 270 11798 6246
rect 11922 270 11956 6246
rect 12054 236 12056 6280
rect 12056 236 12090 6280
rect 12090 236 12092 6280
rect 14046 236 14048 6280
rect 14048 236 14082 6280
rect 14082 236 14084 6280
rect 14182 270 14216 6246
rect 14340 270 14374 6246
rect 14498 270 14532 6246
rect 14656 270 14690 6246
rect 14814 270 14848 6246
rect 14972 270 15006 6246
rect 15130 270 15164 6246
rect 15288 270 15322 6246
rect 15446 270 15480 6246
rect 15604 270 15638 6246
rect 15762 270 15796 6246
rect 15920 270 15954 6246
rect 16078 270 16112 6246
rect 16236 270 16270 6246
rect 16394 270 16428 6246
rect 16552 270 16586 6246
rect 16710 270 16744 6246
rect 16868 270 16902 6246
rect 17026 270 17060 6246
rect 17184 270 17218 6246
rect 17342 270 17376 6246
rect 17500 270 17534 6246
rect 17658 270 17692 6246
rect 17816 270 17850 6246
rect 17974 270 18008 6246
rect 18132 270 18166 6246
rect 18290 270 18324 6246
rect 18448 270 18482 6246
rect 18606 270 18640 6246
rect 18764 270 18798 6246
rect 18922 270 18956 6246
rect 19054 236 19056 6280
rect 19056 236 19090 6280
rect 19090 236 19092 6280
rect 21046 236 21048 6280
rect 21048 236 21082 6280
rect 21082 236 21084 6280
rect 21182 270 21216 6246
rect 21340 270 21374 6246
rect 21498 270 21532 6246
rect 21656 270 21690 6246
rect 21814 270 21848 6246
rect 21972 270 22006 6246
rect 22130 270 22164 6246
rect 22288 270 22322 6246
rect 22446 270 22480 6246
rect 22604 270 22638 6246
rect 22762 270 22796 6246
rect 22920 270 22954 6246
rect 23078 270 23112 6246
rect 23236 270 23270 6246
rect 23394 270 23428 6246
rect 23552 270 23586 6246
rect 23710 270 23744 6246
rect 23868 270 23902 6246
rect 24026 270 24060 6246
rect 24184 270 24218 6246
rect 24342 270 24376 6246
rect 24500 270 24534 6246
rect 24658 270 24692 6246
rect 24816 270 24850 6246
rect 24974 270 25008 6246
rect 25132 270 25166 6246
rect 25290 270 25324 6246
rect 25448 270 25482 6246
rect 25606 270 25640 6246
rect 25764 270 25798 6246
rect 25922 270 25956 6246
rect 26054 236 26056 6280
rect 26056 236 26090 6280
rect 26090 236 26092 6280
rect 244 186 312 220
rect 402 186 470 220
rect 560 186 628 220
rect 718 186 786 220
rect 876 186 944 220
rect 1034 186 1102 220
rect 1192 186 1260 220
rect 1350 186 1418 220
rect 1508 186 1576 220
rect 1666 186 1734 220
rect 1824 186 1892 220
rect 1982 186 2050 220
rect 2140 186 2208 220
rect 2298 186 2366 220
rect 2456 186 2524 220
rect 2614 186 2682 220
rect 2772 186 2840 220
rect 2930 186 2998 220
rect 3088 186 3156 220
rect 3246 186 3314 220
rect 3404 186 3472 220
rect 3562 186 3630 220
rect 3720 186 3788 220
rect 3878 186 3946 220
rect 4036 186 4104 220
rect 4194 186 4262 220
rect 4352 186 4420 220
rect 4510 186 4578 220
rect 4668 186 4736 220
rect 4826 186 4894 220
rect 236 82 4902 84
rect 236 48 4902 82
rect 7244 186 7312 220
rect 7402 186 7470 220
rect 7560 186 7628 220
rect 7718 186 7786 220
rect 7876 186 7944 220
rect 8034 186 8102 220
rect 8192 186 8260 220
rect 8350 186 8418 220
rect 8508 186 8576 220
rect 8666 186 8734 220
rect 8824 186 8892 220
rect 8982 186 9050 220
rect 9140 186 9208 220
rect 9298 186 9366 220
rect 9456 186 9524 220
rect 9614 186 9682 220
rect 9772 186 9840 220
rect 9930 186 9998 220
rect 10088 186 10156 220
rect 10246 186 10314 220
rect 10404 186 10472 220
rect 10562 186 10630 220
rect 10720 186 10788 220
rect 10878 186 10946 220
rect 11036 186 11104 220
rect 11194 186 11262 220
rect 11352 186 11420 220
rect 11510 186 11578 220
rect 11668 186 11736 220
rect 11826 186 11894 220
rect 7236 82 11902 84
rect 7236 48 11902 82
rect 14244 186 14312 220
rect 14402 186 14470 220
rect 14560 186 14628 220
rect 14718 186 14786 220
rect 14876 186 14944 220
rect 15034 186 15102 220
rect 15192 186 15260 220
rect 15350 186 15418 220
rect 15508 186 15576 220
rect 15666 186 15734 220
rect 15824 186 15892 220
rect 15982 186 16050 220
rect 16140 186 16208 220
rect 16298 186 16366 220
rect 16456 186 16524 220
rect 16614 186 16682 220
rect 16772 186 16840 220
rect 16930 186 16998 220
rect 17088 186 17156 220
rect 17246 186 17314 220
rect 17404 186 17472 220
rect 17562 186 17630 220
rect 17720 186 17788 220
rect 17878 186 17946 220
rect 18036 186 18104 220
rect 18194 186 18262 220
rect 18352 186 18420 220
rect 18510 186 18578 220
rect 18668 186 18736 220
rect 18826 186 18894 220
rect 14236 82 18902 84
rect 14236 48 18902 82
rect 21244 186 21312 220
rect 21402 186 21470 220
rect 21560 186 21628 220
rect 21718 186 21786 220
rect 21876 186 21944 220
rect 22034 186 22102 220
rect 22192 186 22260 220
rect 22350 186 22418 220
rect 22508 186 22576 220
rect 22666 186 22734 220
rect 22824 186 22892 220
rect 22982 186 23050 220
rect 23140 186 23208 220
rect 23298 186 23366 220
rect 23456 186 23524 220
rect 23614 186 23682 220
rect 23772 186 23840 220
rect 23930 186 23998 220
rect 24088 186 24156 220
rect 24246 186 24314 220
rect 24404 186 24472 220
rect 24562 186 24630 220
rect 24720 186 24788 220
rect 24878 186 24946 220
rect 25036 186 25104 220
rect 25194 186 25262 220
rect 25352 186 25420 220
rect 25510 186 25578 220
rect 25668 186 25736 220
rect 25826 186 25894 220
rect 21236 82 25902 84
rect 21236 48 25902 82
rect 236 46 4902 48
rect 7236 46 11902 48
rect 14236 46 18902 48
rect 21236 46 25902 48
rect 236 -532 4959 -530
rect 7236 -532 11959 -530
rect 14236 -532 18959 -530
rect 21236 -532 25959 -530
rect 236 -566 4959 -532
rect 236 -568 4959 -566
rect 244 -704 312 -670
rect 402 -704 470 -670
rect 560 -704 628 -670
rect 718 -704 786 -670
rect 876 -704 944 -670
rect 1034 -704 1102 -670
rect 1192 -704 1260 -670
rect 1350 -704 1418 -670
rect 1508 -704 1576 -670
rect 1666 -704 1734 -670
rect 1824 -704 1892 -670
rect 1982 -704 2050 -670
rect 2140 -704 2208 -670
rect 2298 -704 2366 -670
rect 2456 -704 2524 -670
rect 2614 -704 2682 -670
rect 2772 -704 2840 -670
rect 2930 -704 2998 -670
rect 3088 -704 3156 -670
rect 3246 -704 3314 -670
rect 3404 -704 3472 -670
rect 3562 -704 3630 -670
rect 3720 -704 3788 -670
rect 3878 -704 3946 -670
rect 4036 -704 4104 -670
rect 4194 -704 4262 -670
rect 4352 -704 4420 -670
rect 4510 -704 4578 -670
rect 4668 -704 4736 -670
rect 4826 -704 4894 -670
rect 7236 -566 11959 -532
rect 7236 -568 11959 -566
rect 7244 -704 7312 -670
rect 7402 -704 7470 -670
rect 7560 -704 7628 -670
rect 7718 -704 7786 -670
rect 7876 -704 7944 -670
rect 8034 -704 8102 -670
rect 8192 -704 8260 -670
rect 8350 -704 8418 -670
rect 8508 -704 8576 -670
rect 8666 -704 8734 -670
rect 8824 -704 8892 -670
rect 8982 -704 9050 -670
rect 9140 -704 9208 -670
rect 9298 -704 9366 -670
rect 9456 -704 9524 -670
rect 9614 -704 9682 -670
rect 9772 -704 9840 -670
rect 9930 -704 9998 -670
rect 10088 -704 10156 -670
rect 10246 -704 10314 -670
rect 10404 -704 10472 -670
rect 10562 -704 10630 -670
rect 10720 -704 10788 -670
rect 10878 -704 10946 -670
rect 11036 -704 11104 -670
rect 11194 -704 11262 -670
rect 11352 -704 11420 -670
rect 11510 -704 11578 -670
rect 11668 -704 11736 -670
rect 11826 -704 11894 -670
rect 14236 -566 18959 -532
rect 14236 -568 18959 -566
rect 14244 -704 14312 -670
rect 14402 -704 14470 -670
rect 14560 -704 14628 -670
rect 14718 -704 14786 -670
rect 14876 -704 14944 -670
rect 15034 -704 15102 -670
rect 15192 -704 15260 -670
rect 15350 -704 15418 -670
rect 15508 -704 15576 -670
rect 15666 -704 15734 -670
rect 15824 -704 15892 -670
rect 15982 -704 16050 -670
rect 16140 -704 16208 -670
rect 16298 -704 16366 -670
rect 16456 -704 16524 -670
rect 16614 -704 16682 -670
rect 16772 -704 16840 -670
rect 16930 -704 16998 -670
rect 17088 -704 17156 -670
rect 17246 -704 17314 -670
rect 17404 -704 17472 -670
rect 17562 -704 17630 -670
rect 17720 -704 17788 -670
rect 17878 -704 17946 -670
rect 18036 -704 18104 -670
rect 18194 -704 18262 -670
rect 18352 -704 18420 -670
rect 18510 -704 18578 -670
rect 18668 -704 18736 -670
rect 18826 -704 18894 -670
rect 21236 -566 25959 -532
rect 21236 -568 25959 -566
rect 21244 -704 21312 -670
rect 21402 -704 21470 -670
rect 21560 -704 21628 -670
rect 21718 -704 21786 -670
rect 21876 -704 21944 -670
rect 22034 -704 22102 -670
rect 22192 -704 22260 -670
rect 22350 -704 22418 -670
rect 22508 -704 22576 -670
rect 22666 -704 22734 -670
rect 22824 -704 22892 -670
rect 22982 -704 23050 -670
rect 23140 -704 23208 -670
rect 23298 -704 23366 -670
rect 23456 -704 23524 -670
rect 23614 -704 23682 -670
rect 23772 -704 23840 -670
rect 23930 -704 23998 -670
rect 24088 -704 24156 -670
rect 24246 -704 24314 -670
rect 24404 -704 24472 -670
rect 24562 -704 24630 -670
rect 24720 -704 24788 -670
rect 24878 -704 24946 -670
rect 25036 -704 25104 -670
rect 25194 -704 25262 -670
rect 25352 -704 25420 -670
rect 25510 -704 25578 -670
rect 25668 -704 25736 -670
rect 25826 -704 25894 -670
rect 46 -6764 48 -720
rect 48 -6764 82 -720
rect 82 -6764 84 -720
rect 182 -6730 216 -754
rect 340 -6730 374 -754
rect 498 -6730 532 -754
rect 656 -6730 690 -754
rect 814 -6730 848 -754
rect 972 -6730 1006 -754
rect 1130 -6730 1164 -754
rect 1288 -6730 1322 -754
rect 1446 -6730 1480 -754
rect 1604 -6730 1638 -754
rect 1762 -6730 1796 -754
rect 1920 -6730 1954 -754
rect 2078 -6730 2112 -754
rect 2236 -6730 2270 -754
rect 2394 -6730 2428 -754
rect 2552 -6730 2586 -754
rect 2710 -6730 2744 -754
rect 2868 -6730 2902 -754
rect 3026 -6730 3060 -754
rect 3184 -6730 3218 -754
rect 3342 -6730 3376 -754
rect 3500 -6730 3534 -754
rect 3658 -6730 3692 -754
rect 3816 -6730 3850 -754
rect 3974 -6730 4008 -754
rect 4132 -6730 4166 -754
rect 4290 -6730 4324 -754
rect 4448 -6730 4482 -754
rect 4606 -6730 4640 -754
rect 4764 -6730 4798 -754
rect 4922 -6730 4956 -754
rect 5054 -6764 5056 -720
rect 5056 -6764 5090 -720
rect 5090 -6764 5092 -720
rect 7046 -6764 7048 -720
rect 7048 -6764 7082 -720
rect 7082 -6764 7084 -720
rect 7182 -6730 7216 -754
rect 7340 -6730 7374 -754
rect 7498 -6730 7532 -754
rect 7656 -6730 7690 -754
rect 7814 -6730 7848 -754
rect 7972 -6730 8006 -754
rect 8130 -6730 8164 -754
rect 8288 -6730 8322 -754
rect 8446 -6730 8480 -754
rect 8604 -6730 8638 -754
rect 8762 -6730 8796 -754
rect 8920 -6730 8954 -754
rect 9078 -6730 9112 -754
rect 9236 -6730 9270 -754
rect 9394 -6730 9428 -754
rect 9552 -6730 9586 -754
rect 9710 -6730 9744 -754
rect 9868 -6730 9902 -754
rect 10026 -6730 10060 -754
rect 10184 -6730 10218 -754
rect 10342 -6730 10376 -754
rect 10500 -6730 10534 -754
rect 10658 -6730 10692 -754
rect 10816 -6730 10850 -754
rect 10974 -6730 11008 -754
rect 11132 -6730 11166 -754
rect 11290 -6730 11324 -754
rect 11448 -6730 11482 -754
rect 11606 -6730 11640 -754
rect 11764 -6730 11798 -754
rect 11922 -6730 11956 -754
rect 12054 -6764 12056 -720
rect 12056 -6764 12090 -720
rect 12090 -6764 12092 -720
rect 14046 -6764 14048 -720
rect 14048 -6764 14082 -720
rect 14082 -6764 14084 -720
rect 14182 -6730 14216 -754
rect 14340 -6730 14374 -754
rect 14498 -6730 14532 -754
rect 14656 -6730 14690 -754
rect 14814 -6730 14848 -754
rect 14972 -6730 15006 -754
rect 15130 -6730 15164 -754
rect 15288 -6730 15322 -754
rect 15446 -6730 15480 -754
rect 15604 -6730 15638 -754
rect 15762 -6730 15796 -754
rect 15920 -6730 15954 -754
rect 16078 -6730 16112 -754
rect 16236 -6730 16270 -754
rect 16394 -6730 16428 -754
rect 16552 -6730 16586 -754
rect 16710 -6730 16744 -754
rect 16868 -6730 16902 -754
rect 17026 -6730 17060 -754
rect 17184 -6730 17218 -754
rect 17342 -6730 17376 -754
rect 17500 -6730 17534 -754
rect 17658 -6730 17692 -754
rect 17816 -6730 17850 -754
rect 17974 -6730 18008 -754
rect 18132 -6730 18166 -754
rect 18290 -6730 18324 -754
rect 18448 -6730 18482 -754
rect 18606 -6730 18640 -754
rect 18764 -6730 18798 -754
rect 18922 -6730 18956 -754
rect 19054 -6764 19056 -720
rect 19056 -6764 19090 -720
rect 19090 -6764 19092 -720
rect 21046 -6764 21048 -720
rect 21048 -6764 21082 -720
rect 21082 -6764 21084 -720
rect 21182 -6730 21216 -754
rect 21340 -6730 21374 -754
rect 21498 -6730 21532 -754
rect 21656 -6730 21690 -754
rect 21814 -6730 21848 -754
rect 21972 -6730 22006 -754
rect 22130 -6730 22164 -754
rect 22288 -6730 22322 -754
rect 22446 -6730 22480 -754
rect 22604 -6730 22638 -754
rect 22762 -6730 22796 -754
rect 22920 -6730 22954 -754
rect 23078 -6730 23112 -754
rect 23236 -6730 23270 -754
rect 23394 -6730 23428 -754
rect 23552 -6730 23586 -754
rect 23710 -6730 23744 -754
rect 23868 -6730 23902 -754
rect 24026 -6730 24060 -754
rect 24184 -6730 24218 -754
rect 24342 -6730 24376 -754
rect 24500 -6730 24534 -754
rect 24658 -6730 24692 -754
rect 24816 -6730 24850 -754
rect 24974 -6730 25008 -754
rect 25132 -6730 25166 -754
rect 25290 -6730 25324 -754
rect 25448 -6730 25482 -754
rect 25606 -6730 25640 -754
rect 25764 -6730 25798 -754
rect 25922 -6730 25956 -754
rect 26054 -6764 26056 -720
rect 26056 -6764 26090 -720
rect 26090 -6764 26092 -720
rect 244 -6814 312 -6780
rect 402 -6814 470 -6780
rect 560 -6814 628 -6780
rect 718 -6814 786 -6780
rect 876 -6814 944 -6780
rect 1034 -6814 1102 -6780
rect 1192 -6814 1260 -6780
rect 1350 -6814 1418 -6780
rect 1508 -6814 1576 -6780
rect 1666 -6814 1734 -6780
rect 1824 -6814 1892 -6780
rect 1982 -6814 2050 -6780
rect 2140 -6814 2208 -6780
rect 2298 -6814 2366 -6780
rect 2456 -6814 2524 -6780
rect 2614 -6814 2682 -6780
rect 2772 -6814 2840 -6780
rect 2930 -6814 2998 -6780
rect 3088 -6814 3156 -6780
rect 3246 -6814 3314 -6780
rect 3404 -6814 3472 -6780
rect 3562 -6814 3630 -6780
rect 3720 -6814 3788 -6780
rect 3878 -6814 3946 -6780
rect 4036 -6814 4104 -6780
rect 4194 -6814 4262 -6780
rect 4352 -6814 4420 -6780
rect 4510 -6814 4578 -6780
rect 4668 -6814 4736 -6780
rect 4826 -6814 4894 -6780
rect 236 -6918 4902 -6916
rect 236 -6952 4902 -6918
rect 7244 -6814 7312 -6780
rect 7402 -6814 7470 -6780
rect 7560 -6814 7628 -6780
rect 7718 -6814 7786 -6780
rect 7876 -6814 7944 -6780
rect 8034 -6814 8102 -6780
rect 8192 -6814 8260 -6780
rect 8350 -6814 8418 -6780
rect 8508 -6814 8576 -6780
rect 8666 -6814 8734 -6780
rect 8824 -6814 8892 -6780
rect 8982 -6814 9050 -6780
rect 9140 -6814 9208 -6780
rect 9298 -6814 9366 -6780
rect 9456 -6814 9524 -6780
rect 9614 -6814 9682 -6780
rect 9772 -6814 9840 -6780
rect 9930 -6814 9998 -6780
rect 10088 -6814 10156 -6780
rect 10246 -6814 10314 -6780
rect 10404 -6814 10472 -6780
rect 10562 -6814 10630 -6780
rect 10720 -6814 10788 -6780
rect 10878 -6814 10946 -6780
rect 11036 -6814 11104 -6780
rect 11194 -6814 11262 -6780
rect 11352 -6814 11420 -6780
rect 11510 -6814 11578 -6780
rect 11668 -6814 11736 -6780
rect 11826 -6814 11894 -6780
rect 7236 -6918 11902 -6916
rect 7236 -6952 11902 -6918
rect 14244 -6814 14312 -6780
rect 14402 -6814 14470 -6780
rect 14560 -6814 14628 -6780
rect 14718 -6814 14786 -6780
rect 14876 -6814 14944 -6780
rect 15034 -6814 15102 -6780
rect 15192 -6814 15260 -6780
rect 15350 -6814 15418 -6780
rect 15508 -6814 15576 -6780
rect 15666 -6814 15734 -6780
rect 15824 -6814 15892 -6780
rect 15982 -6814 16050 -6780
rect 16140 -6814 16208 -6780
rect 16298 -6814 16366 -6780
rect 16456 -6814 16524 -6780
rect 16614 -6814 16682 -6780
rect 16772 -6814 16840 -6780
rect 16930 -6814 16998 -6780
rect 17088 -6814 17156 -6780
rect 17246 -6814 17314 -6780
rect 17404 -6814 17472 -6780
rect 17562 -6814 17630 -6780
rect 17720 -6814 17788 -6780
rect 17878 -6814 17946 -6780
rect 18036 -6814 18104 -6780
rect 18194 -6814 18262 -6780
rect 18352 -6814 18420 -6780
rect 18510 -6814 18578 -6780
rect 18668 -6814 18736 -6780
rect 18826 -6814 18894 -6780
rect 14236 -6918 18902 -6916
rect 14236 -6952 18902 -6918
rect 21244 -6814 21312 -6780
rect 21402 -6814 21470 -6780
rect 21560 -6814 21628 -6780
rect 21718 -6814 21786 -6780
rect 21876 -6814 21944 -6780
rect 22034 -6814 22102 -6780
rect 22192 -6814 22260 -6780
rect 22350 -6814 22418 -6780
rect 22508 -6814 22576 -6780
rect 22666 -6814 22734 -6780
rect 22824 -6814 22892 -6780
rect 22982 -6814 23050 -6780
rect 23140 -6814 23208 -6780
rect 23298 -6814 23366 -6780
rect 23456 -6814 23524 -6780
rect 23614 -6814 23682 -6780
rect 23772 -6814 23840 -6780
rect 23930 -6814 23998 -6780
rect 24088 -6814 24156 -6780
rect 24246 -6814 24314 -6780
rect 24404 -6814 24472 -6780
rect 24562 -6814 24630 -6780
rect 24720 -6814 24788 -6780
rect 24878 -6814 24946 -6780
rect 25036 -6814 25104 -6780
rect 25194 -6814 25262 -6780
rect 25352 -6814 25420 -6780
rect 25510 -6814 25578 -6780
rect 25668 -6814 25736 -6780
rect 25826 -6814 25894 -6780
rect 21236 -6918 25902 -6916
rect 21236 -6952 25902 -6918
rect 236 -6954 4902 -6952
rect 7236 -6954 11902 -6952
rect 14236 -6954 18902 -6952
rect 21236 -6954 25902 -6952
<< metal1 >>
rect 30 6470 5110 6480
rect 30 6432 236 6470
rect 4959 6432 5110 6470
rect 30 6422 5110 6432
rect 30 6420 100 6422
rect 5040 6420 5110 6422
rect 232 6330 252 6390
rect 4886 6330 4906 6390
rect 232 6296 244 6330
rect 4894 6296 4906 6330
rect 232 6290 252 6296
rect 4886 6290 4906 6296
rect 165 6246 231 6258
rect 165 6238 182 6246
rect 216 6238 231 6246
rect 165 270 182 278
rect 216 270 231 278
rect 165 258 231 270
rect 323 6246 389 6258
rect 323 6238 340 6246
rect 374 6238 389 6246
rect 323 270 340 278
rect 374 270 389 278
rect 323 258 389 270
rect 481 6246 547 6258
rect 481 6238 498 6246
rect 532 6238 547 6246
rect 481 270 498 278
rect 532 270 547 278
rect 481 258 547 270
rect 639 6246 705 6258
rect 639 6238 656 6246
rect 690 6238 705 6246
rect 639 270 656 278
rect 690 270 705 278
rect 639 258 705 270
rect 797 6246 863 6258
rect 797 6238 814 6246
rect 848 6238 863 6246
rect 797 270 814 278
rect 848 270 863 278
rect 797 258 863 270
rect 955 6246 1021 6258
rect 955 6238 972 6246
rect 1006 6238 1021 6246
rect 955 270 972 278
rect 1006 270 1021 278
rect 955 258 1021 270
rect 1113 6246 1179 6258
rect 1113 6238 1130 6246
rect 1164 6238 1179 6246
rect 1113 270 1130 278
rect 1164 270 1179 278
rect 1113 258 1179 270
rect 1271 6246 1337 6258
rect 1271 6238 1288 6246
rect 1322 6238 1337 6246
rect 1271 270 1288 278
rect 1322 270 1337 278
rect 1271 258 1337 270
rect 1429 6246 1495 6258
rect 1429 6238 1446 6246
rect 1480 6238 1495 6246
rect 1429 270 1446 278
rect 1480 270 1495 278
rect 1429 258 1495 270
rect 1587 6246 1653 6258
rect 1587 6238 1604 6246
rect 1638 6238 1653 6246
rect 1587 270 1604 278
rect 1638 270 1653 278
rect 1587 258 1653 270
rect 1745 6246 1811 6258
rect 1745 6238 1762 6246
rect 1796 6238 1811 6246
rect 1745 270 1762 278
rect 1796 270 1811 278
rect 1745 258 1811 270
rect 1903 6246 1969 6258
rect 1903 6238 1920 6246
rect 1954 6238 1969 6246
rect 1903 270 1920 278
rect 1954 270 1969 278
rect 1903 258 1969 270
rect 2061 6246 2127 6258
rect 2061 6238 2078 6246
rect 2112 6238 2127 6246
rect 2061 270 2078 278
rect 2112 270 2127 278
rect 2061 258 2127 270
rect 2219 6246 2285 6258
rect 2219 6238 2236 6246
rect 2270 6238 2285 6246
rect 2219 270 2236 278
rect 2270 270 2285 278
rect 2219 258 2285 270
rect 2377 6246 2443 6258
rect 2377 6238 2394 6246
rect 2428 6238 2443 6246
rect 2377 270 2394 278
rect 2428 270 2443 278
rect 2377 258 2443 270
rect 2535 6246 2601 6258
rect 2535 6238 2552 6246
rect 2586 6238 2601 6246
rect 2535 270 2552 278
rect 2586 270 2601 278
rect 2535 258 2601 270
rect 2693 6246 2759 6258
rect 2693 6238 2710 6246
rect 2744 6238 2759 6246
rect 2693 270 2710 278
rect 2744 270 2759 278
rect 2693 258 2759 270
rect 2851 6246 2917 6258
rect 2851 6238 2868 6246
rect 2902 6238 2917 6246
rect 2851 270 2868 278
rect 2902 270 2917 278
rect 2851 258 2917 270
rect 3009 6246 3075 6258
rect 3009 6238 3026 6246
rect 3060 6238 3075 6246
rect 3009 270 3026 278
rect 3060 270 3075 278
rect 3009 258 3075 270
rect 3167 6246 3233 6258
rect 3167 6238 3184 6246
rect 3218 6238 3233 6246
rect 3167 270 3184 278
rect 3218 270 3233 278
rect 3167 258 3233 270
rect 3325 6246 3391 6258
rect 3325 6238 3342 6246
rect 3376 6238 3391 6246
rect 3325 270 3342 278
rect 3376 270 3391 278
rect 3325 258 3391 270
rect 3483 6246 3549 6258
rect 3483 6238 3500 6246
rect 3534 6238 3549 6246
rect 3483 270 3500 278
rect 3534 270 3549 278
rect 3483 258 3549 270
rect 3641 6246 3707 6258
rect 3641 6238 3658 6246
rect 3692 6238 3707 6246
rect 3641 270 3658 278
rect 3692 270 3707 278
rect 3641 258 3707 270
rect 3799 6246 3865 6258
rect 3799 6238 3816 6246
rect 3850 6238 3865 6246
rect 3799 270 3816 278
rect 3850 270 3865 278
rect 3799 258 3865 270
rect 3957 6246 4023 6258
rect 3957 6238 3974 6246
rect 4008 6238 4023 6246
rect 3957 270 3974 278
rect 4008 270 4023 278
rect 3957 258 4023 270
rect 4115 6246 4181 6258
rect 4115 6238 4132 6246
rect 4166 6238 4181 6246
rect 4115 270 4132 278
rect 4166 270 4181 278
rect 4115 258 4181 270
rect 4273 6246 4339 6258
rect 4273 6238 4290 6246
rect 4324 6238 4339 6246
rect 4273 270 4290 278
rect 4324 270 4339 278
rect 4273 258 4339 270
rect 4431 6246 4497 6258
rect 4431 6238 4448 6246
rect 4482 6238 4497 6246
rect 4431 270 4448 278
rect 4482 270 4497 278
rect 4431 258 4497 270
rect 4589 6246 4655 6258
rect 4589 6238 4606 6246
rect 4640 6238 4655 6246
rect 4589 270 4606 278
rect 4640 270 4655 278
rect 4589 258 4655 270
rect 4747 6246 4813 6258
rect 4747 6238 4764 6246
rect 4798 6238 4813 6246
rect 4747 270 4764 278
rect 4798 270 4813 278
rect 4747 258 4813 270
rect 4905 6246 4971 6258
rect 4905 6238 4922 6246
rect 4956 6238 4971 6246
rect 4905 270 4922 278
rect 4956 270 4971 278
rect 4905 258 4971 270
rect 232 220 252 226
rect 4886 220 4906 226
rect 232 186 244 220
rect 4894 186 4906 220
rect 232 126 252 186
rect 4886 126 4906 186
rect 30 94 100 100
rect 5040 94 5110 100
rect 30 84 5110 94
rect 30 46 236 84
rect 4902 46 5110 84
rect 30 30 5110 46
rect 7030 6470 12110 6480
rect 7030 6432 7236 6470
rect 11959 6432 12110 6470
rect 7030 6422 12110 6432
rect 7030 6420 7100 6422
rect 12040 6420 12110 6422
rect 7232 6330 7252 6390
rect 11886 6330 11906 6390
rect 7232 6296 7244 6330
rect 11894 6296 11906 6330
rect 7232 6290 7252 6296
rect 11886 6290 11906 6296
rect 7165 6246 7231 6258
rect 7165 6238 7182 6246
rect 7216 6238 7231 6246
rect 7165 270 7182 278
rect 7216 270 7231 278
rect 7165 258 7231 270
rect 7323 6246 7389 6258
rect 7323 6238 7340 6246
rect 7374 6238 7389 6246
rect 7323 270 7340 278
rect 7374 270 7389 278
rect 7323 258 7389 270
rect 7481 6246 7547 6258
rect 7481 6238 7498 6246
rect 7532 6238 7547 6246
rect 7481 270 7498 278
rect 7532 270 7547 278
rect 7481 258 7547 270
rect 7639 6246 7705 6258
rect 7639 6238 7656 6246
rect 7690 6238 7705 6246
rect 7639 270 7656 278
rect 7690 270 7705 278
rect 7639 258 7705 270
rect 7797 6246 7863 6258
rect 7797 6238 7814 6246
rect 7848 6238 7863 6246
rect 7797 270 7814 278
rect 7848 270 7863 278
rect 7797 258 7863 270
rect 7955 6246 8021 6258
rect 7955 6238 7972 6246
rect 8006 6238 8021 6246
rect 7955 270 7972 278
rect 8006 270 8021 278
rect 7955 258 8021 270
rect 8113 6246 8179 6258
rect 8113 6238 8130 6246
rect 8164 6238 8179 6246
rect 8113 270 8130 278
rect 8164 270 8179 278
rect 8113 258 8179 270
rect 8271 6246 8337 6258
rect 8271 6238 8288 6246
rect 8322 6238 8337 6246
rect 8271 270 8288 278
rect 8322 270 8337 278
rect 8271 258 8337 270
rect 8429 6246 8495 6258
rect 8429 6238 8446 6246
rect 8480 6238 8495 6246
rect 8429 270 8446 278
rect 8480 270 8495 278
rect 8429 258 8495 270
rect 8587 6246 8653 6258
rect 8587 6238 8604 6246
rect 8638 6238 8653 6246
rect 8587 270 8604 278
rect 8638 270 8653 278
rect 8587 258 8653 270
rect 8745 6246 8811 6258
rect 8745 6238 8762 6246
rect 8796 6238 8811 6246
rect 8745 270 8762 278
rect 8796 270 8811 278
rect 8745 258 8811 270
rect 8903 6246 8969 6258
rect 8903 6238 8920 6246
rect 8954 6238 8969 6246
rect 8903 270 8920 278
rect 8954 270 8969 278
rect 8903 258 8969 270
rect 9061 6246 9127 6258
rect 9061 6238 9078 6246
rect 9112 6238 9127 6246
rect 9061 270 9078 278
rect 9112 270 9127 278
rect 9061 258 9127 270
rect 9219 6246 9285 6258
rect 9219 6238 9236 6246
rect 9270 6238 9285 6246
rect 9219 270 9236 278
rect 9270 270 9285 278
rect 9219 258 9285 270
rect 9377 6246 9443 6258
rect 9377 6238 9394 6246
rect 9428 6238 9443 6246
rect 9377 270 9394 278
rect 9428 270 9443 278
rect 9377 258 9443 270
rect 9535 6246 9601 6258
rect 9535 6238 9552 6246
rect 9586 6238 9601 6246
rect 9535 270 9552 278
rect 9586 270 9601 278
rect 9535 258 9601 270
rect 9693 6246 9759 6258
rect 9693 6238 9710 6246
rect 9744 6238 9759 6246
rect 9693 270 9710 278
rect 9744 270 9759 278
rect 9693 258 9759 270
rect 9851 6246 9917 6258
rect 9851 6238 9868 6246
rect 9902 6238 9917 6246
rect 9851 270 9868 278
rect 9902 270 9917 278
rect 9851 258 9917 270
rect 10009 6246 10075 6258
rect 10009 6238 10026 6246
rect 10060 6238 10075 6246
rect 10009 270 10026 278
rect 10060 270 10075 278
rect 10009 258 10075 270
rect 10167 6246 10233 6258
rect 10167 6238 10184 6246
rect 10218 6238 10233 6246
rect 10167 270 10184 278
rect 10218 270 10233 278
rect 10167 258 10233 270
rect 10325 6246 10391 6258
rect 10325 6238 10342 6246
rect 10376 6238 10391 6246
rect 10325 270 10342 278
rect 10376 270 10391 278
rect 10325 258 10391 270
rect 10483 6246 10549 6258
rect 10483 6238 10500 6246
rect 10534 6238 10549 6246
rect 10483 270 10500 278
rect 10534 270 10549 278
rect 10483 258 10549 270
rect 10641 6246 10707 6258
rect 10641 6238 10658 6246
rect 10692 6238 10707 6246
rect 10641 270 10658 278
rect 10692 270 10707 278
rect 10641 258 10707 270
rect 10799 6246 10865 6258
rect 10799 6238 10816 6246
rect 10850 6238 10865 6246
rect 10799 270 10816 278
rect 10850 270 10865 278
rect 10799 258 10865 270
rect 10957 6246 11023 6258
rect 10957 6238 10974 6246
rect 11008 6238 11023 6246
rect 10957 270 10974 278
rect 11008 270 11023 278
rect 10957 258 11023 270
rect 11115 6246 11181 6258
rect 11115 6238 11132 6246
rect 11166 6238 11181 6246
rect 11115 270 11132 278
rect 11166 270 11181 278
rect 11115 258 11181 270
rect 11273 6246 11339 6258
rect 11273 6238 11290 6246
rect 11324 6238 11339 6246
rect 11273 270 11290 278
rect 11324 270 11339 278
rect 11273 258 11339 270
rect 11431 6246 11497 6258
rect 11431 6238 11448 6246
rect 11482 6238 11497 6246
rect 11431 270 11448 278
rect 11482 270 11497 278
rect 11431 258 11497 270
rect 11589 6246 11655 6258
rect 11589 6238 11606 6246
rect 11640 6238 11655 6246
rect 11589 270 11606 278
rect 11640 270 11655 278
rect 11589 258 11655 270
rect 11747 6246 11813 6258
rect 11747 6238 11764 6246
rect 11798 6238 11813 6246
rect 11747 270 11764 278
rect 11798 270 11813 278
rect 11747 258 11813 270
rect 11905 6246 11971 6258
rect 11905 6238 11922 6246
rect 11956 6238 11971 6246
rect 11905 270 11922 278
rect 11956 270 11971 278
rect 11905 258 11971 270
rect 7232 220 7252 226
rect 11886 220 11906 226
rect 7232 186 7244 220
rect 11894 186 11906 220
rect 7232 126 7252 186
rect 11886 126 11906 186
rect 7030 94 7100 100
rect 12040 94 12110 100
rect 7030 84 12110 94
rect 7030 46 7236 84
rect 11902 46 12110 84
rect 7030 30 12110 46
rect 14030 6470 19110 6480
rect 14030 6432 14236 6470
rect 18959 6432 19110 6470
rect 14030 6422 19110 6432
rect 14030 6420 14100 6422
rect 19040 6420 19110 6422
rect 14232 6330 14252 6390
rect 18886 6330 18906 6390
rect 14232 6296 14244 6330
rect 18894 6296 18906 6330
rect 14232 6290 14252 6296
rect 18886 6290 18906 6296
rect 14165 6246 14231 6258
rect 14165 6238 14182 6246
rect 14216 6238 14231 6246
rect 14165 270 14182 278
rect 14216 270 14231 278
rect 14165 258 14231 270
rect 14323 6246 14389 6258
rect 14323 6238 14340 6246
rect 14374 6238 14389 6246
rect 14323 270 14340 278
rect 14374 270 14389 278
rect 14323 258 14389 270
rect 14481 6246 14547 6258
rect 14481 6238 14498 6246
rect 14532 6238 14547 6246
rect 14481 270 14498 278
rect 14532 270 14547 278
rect 14481 258 14547 270
rect 14639 6246 14705 6258
rect 14639 6238 14656 6246
rect 14690 6238 14705 6246
rect 14639 270 14656 278
rect 14690 270 14705 278
rect 14639 258 14705 270
rect 14797 6246 14863 6258
rect 14797 6238 14814 6246
rect 14848 6238 14863 6246
rect 14797 270 14814 278
rect 14848 270 14863 278
rect 14797 258 14863 270
rect 14955 6246 15021 6258
rect 14955 6238 14972 6246
rect 15006 6238 15021 6246
rect 14955 270 14972 278
rect 15006 270 15021 278
rect 14955 258 15021 270
rect 15113 6246 15179 6258
rect 15113 6238 15130 6246
rect 15164 6238 15179 6246
rect 15113 270 15130 278
rect 15164 270 15179 278
rect 15113 258 15179 270
rect 15271 6246 15337 6258
rect 15271 6238 15288 6246
rect 15322 6238 15337 6246
rect 15271 270 15288 278
rect 15322 270 15337 278
rect 15271 258 15337 270
rect 15429 6246 15495 6258
rect 15429 6238 15446 6246
rect 15480 6238 15495 6246
rect 15429 270 15446 278
rect 15480 270 15495 278
rect 15429 258 15495 270
rect 15587 6246 15653 6258
rect 15587 6238 15604 6246
rect 15638 6238 15653 6246
rect 15587 270 15604 278
rect 15638 270 15653 278
rect 15587 258 15653 270
rect 15745 6246 15811 6258
rect 15745 6238 15762 6246
rect 15796 6238 15811 6246
rect 15745 270 15762 278
rect 15796 270 15811 278
rect 15745 258 15811 270
rect 15903 6246 15969 6258
rect 15903 6238 15920 6246
rect 15954 6238 15969 6246
rect 15903 270 15920 278
rect 15954 270 15969 278
rect 15903 258 15969 270
rect 16061 6246 16127 6258
rect 16061 6238 16078 6246
rect 16112 6238 16127 6246
rect 16061 270 16078 278
rect 16112 270 16127 278
rect 16061 258 16127 270
rect 16219 6246 16285 6258
rect 16219 6238 16236 6246
rect 16270 6238 16285 6246
rect 16219 270 16236 278
rect 16270 270 16285 278
rect 16219 258 16285 270
rect 16377 6246 16443 6258
rect 16377 6238 16394 6246
rect 16428 6238 16443 6246
rect 16377 270 16394 278
rect 16428 270 16443 278
rect 16377 258 16443 270
rect 16535 6246 16601 6258
rect 16535 6238 16552 6246
rect 16586 6238 16601 6246
rect 16535 270 16552 278
rect 16586 270 16601 278
rect 16535 258 16601 270
rect 16693 6246 16759 6258
rect 16693 6238 16710 6246
rect 16744 6238 16759 6246
rect 16693 270 16710 278
rect 16744 270 16759 278
rect 16693 258 16759 270
rect 16851 6246 16917 6258
rect 16851 6238 16868 6246
rect 16902 6238 16917 6246
rect 16851 270 16868 278
rect 16902 270 16917 278
rect 16851 258 16917 270
rect 17009 6246 17075 6258
rect 17009 6238 17026 6246
rect 17060 6238 17075 6246
rect 17009 270 17026 278
rect 17060 270 17075 278
rect 17009 258 17075 270
rect 17167 6246 17233 6258
rect 17167 6238 17184 6246
rect 17218 6238 17233 6246
rect 17167 270 17184 278
rect 17218 270 17233 278
rect 17167 258 17233 270
rect 17325 6246 17391 6258
rect 17325 6238 17342 6246
rect 17376 6238 17391 6246
rect 17325 270 17342 278
rect 17376 270 17391 278
rect 17325 258 17391 270
rect 17483 6246 17549 6258
rect 17483 6238 17500 6246
rect 17534 6238 17549 6246
rect 17483 270 17500 278
rect 17534 270 17549 278
rect 17483 258 17549 270
rect 17641 6246 17707 6258
rect 17641 6238 17658 6246
rect 17692 6238 17707 6246
rect 17641 270 17658 278
rect 17692 270 17707 278
rect 17641 258 17707 270
rect 17799 6246 17865 6258
rect 17799 6238 17816 6246
rect 17850 6238 17865 6246
rect 17799 270 17816 278
rect 17850 270 17865 278
rect 17799 258 17865 270
rect 17957 6246 18023 6258
rect 17957 6238 17974 6246
rect 18008 6238 18023 6246
rect 17957 270 17974 278
rect 18008 270 18023 278
rect 17957 258 18023 270
rect 18115 6246 18181 6258
rect 18115 6238 18132 6246
rect 18166 6238 18181 6246
rect 18115 270 18132 278
rect 18166 270 18181 278
rect 18115 258 18181 270
rect 18273 6246 18339 6258
rect 18273 6238 18290 6246
rect 18324 6238 18339 6246
rect 18273 270 18290 278
rect 18324 270 18339 278
rect 18273 258 18339 270
rect 18431 6246 18497 6258
rect 18431 6238 18448 6246
rect 18482 6238 18497 6246
rect 18431 270 18448 278
rect 18482 270 18497 278
rect 18431 258 18497 270
rect 18589 6246 18655 6258
rect 18589 6238 18606 6246
rect 18640 6238 18655 6246
rect 18589 270 18606 278
rect 18640 270 18655 278
rect 18589 258 18655 270
rect 18747 6246 18813 6258
rect 18747 6238 18764 6246
rect 18798 6238 18813 6246
rect 18747 270 18764 278
rect 18798 270 18813 278
rect 18747 258 18813 270
rect 18905 6246 18971 6258
rect 18905 6238 18922 6246
rect 18956 6238 18971 6246
rect 18905 270 18922 278
rect 18956 270 18971 278
rect 18905 258 18971 270
rect 14232 220 14252 226
rect 18886 220 18906 226
rect 14232 186 14244 220
rect 18894 186 18906 220
rect 14232 126 14252 186
rect 18886 126 18906 186
rect 14030 94 14100 100
rect 19040 94 19110 100
rect 14030 84 19110 94
rect 14030 46 14236 84
rect 18902 46 19110 84
rect 14030 30 19110 46
rect 21030 6470 26110 6480
rect 21030 6432 21236 6470
rect 25959 6432 26110 6470
rect 21030 6422 26110 6432
rect 21030 6420 21100 6422
rect 26040 6420 26110 6422
rect 21232 6330 21252 6390
rect 25886 6330 25906 6390
rect 21232 6296 21244 6330
rect 25894 6296 25906 6330
rect 21232 6290 21252 6296
rect 25886 6290 25906 6296
rect 21165 6246 21231 6258
rect 21165 6238 21182 6246
rect 21216 6238 21231 6246
rect 21165 270 21182 278
rect 21216 270 21231 278
rect 21165 258 21231 270
rect 21323 6246 21389 6258
rect 21323 6238 21340 6246
rect 21374 6238 21389 6246
rect 21323 270 21340 278
rect 21374 270 21389 278
rect 21323 258 21389 270
rect 21481 6246 21547 6258
rect 21481 6238 21498 6246
rect 21532 6238 21547 6246
rect 21481 270 21498 278
rect 21532 270 21547 278
rect 21481 258 21547 270
rect 21639 6246 21705 6258
rect 21639 6238 21656 6246
rect 21690 6238 21705 6246
rect 21639 270 21656 278
rect 21690 270 21705 278
rect 21639 258 21705 270
rect 21797 6246 21863 6258
rect 21797 6238 21814 6246
rect 21848 6238 21863 6246
rect 21797 270 21814 278
rect 21848 270 21863 278
rect 21797 258 21863 270
rect 21955 6246 22021 6258
rect 21955 6238 21972 6246
rect 22006 6238 22021 6246
rect 21955 270 21972 278
rect 22006 270 22021 278
rect 21955 258 22021 270
rect 22113 6246 22179 6258
rect 22113 6238 22130 6246
rect 22164 6238 22179 6246
rect 22113 270 22130 278
rect 22164 270 22179 278
rect 22113 258 22179 270
rect 22271 6246 22337 6258
rect 22271 6238 22288 6246
rect 22322 6238 22337 6246
rect 22271 270 22288 278
rect 22322 270 22337 278
rect 22271 258 22337 270
rect 22429 6246 22495 6258
rect 22429 6238 22446 6246
rect 22480 6238 22495 6246
rect 22429 270 22446 278
rect 22480 270 22495 278
rect 22429 258 22495 270
rect 22587 6246 22653 6258
rect 22587 6238 22604 6246
rect 22638 6238 22653 6246
rect 22587 270 22604 278
rect 22638 270 22653 278
rect 22587 258 22653 270
rect 22745 6246 22811 6258
rect 22745 6238 22762 6246
rect 22796 6238 22811 6246
rect 22745 270 22762 278
rect 22796 270 22811 278
rect 22745 258 22811 270
rect 22903 6246 22969 6258
rect 22903 6238 22920 6246
rect 22954 6238 22969 6246
rect 22903 270 22920 278
rect 22954 270 22969 278
rect 22903 258 22969 270
rect 23061 6246 23127 6258
rect 23061 6238 23078 6246
rect 23112 6238 23127 6246
rect 23061 270 23078 278
rect 23112 270 23127 278
rect 23061 258 23127 270
rect 23219 6246 23285 6258
rect 23219 6238 23236 6246
rect 23270 6238 23285 6246
rect 23219 270 23236 278
rect 23270 270 23285 278
rect 23219 258 23285 270
rect 23377 6246 23443 6258
rect 23377 6238 23394 6246
rect 23428 6238 23443 6246
rect 23377 270 23394 278
rect 23428 270 23443 278
rect 23377 258 23443 270
rect 23535 6246 23601 6258
rect 23535 6238 23552 6246
rect 23586 6238 23601 6246
rect 23535 270 23552 278
rect 23586 270 23601 278
rect 23535 258 23601 270
rect 23693 6246 23759 6258
rect 23693 6238 23710 6246
rect 23744 6238 23759 6246
rect 23693 270 23710 278
rect 23744 270 23759 278
rect 23693 258 23759 270
rect 23851 6246 23917 6258
rect 23851 6238 23868 6246
rect 23902 6238 23917 6246
rect 23851 270 23868 278
rect 23902 270 23917 278
rect 23851 258 23917 270
rect 24009 6246 24075 6258
rect 24009 6238 24026 6246
rect 24060 6238 24075 6246
rect 24009 270 24026 278
rect 24060 270 24075 278
rect 24009 258 24075 270
rect 24167 6246 24233 6258
rect 24167 6238 24184 6246
rect 24218 6238 24233 6246
rect 24167 270 24184 278
rect 24218 270 24233 278
rect 24167 258 24233 270
rect 24325 6246 24391 6258
rect 24325 6238 24342 6246
rect 24376 6238 24391 6246
rect 24325 270 24342 278
rect 24376 270 24391 278
rect 24325 258 24391 270
rect 24483 6246 24549 6258
rect 24483 6238 24500 6246
rect 24534 6238 24549 6246
rect 24483 270 24500 278
rect 24534 270 24549 278
rect 24483 258 24549 270
rect 24641 6246 24707 6258
rect 24641 6238 24658 6246
rect 24692 6238 24707 6246
rect 24641 270 24658 278
rect 24692 270 24707 278
rect 24641 258 24707 270
rect 24799 6246 24865 6258
rect 24799 6238 24816 6246
rect 24850 6238 24865 6246
rect 24799 270 24816 278
rect 24850 270 24865 278
rect 24799 258 24865 270
rect 24957 6246 25023 6258
rect 24957 6238 24974 6246
rect 25008 6238 25023 6246
rect 24957 270 24974 278
rect 25008 270 25023 278
rect 24957 258 25023 270
rect 25115 6246 25181 6258
rect 25115 6238 25132 6246
rect 25166 6238 25181 6246
rect 25115 270 25132 278
rect 25166 270 25181 278
rect 25115 258 25181 270
rect 25273 6246 25339 6258
rect 25273 6238 25290 6246
rect 25324 6238 25339 6246
rect 25273 270 25290 278
rect 25324 270 25339 278
rect 25273 258 25339 270
rect 25431 6246 25497 6258
rect 25431 6238 25448 6246
rect 25482 6238 25497 6246
rect 25431 270 25448 278
rect 25482 270 25497 278
rect 25431 258 25497 270
rect 25589 6246 25655 6258
rect 25589 6238 25606 6246
rect 25640 6238 25655 6246
rect 25589 270 25606 278
rect 25640 270 25655 278
rect 25589 258 25655 270
rect 25747 6246 25813 6258
rect 25747 6238 25764 6246
rect 25798 6238 25813 6246
rect 25747 270 25764 278
rect 25798 270 25813 278
rect 25747 258 25813 270
rect 25905 6246 25971 6258
rect 25905 6238 25922 6246
rect 25956 6238 25971 6246
rect 25905 270 25922 278
rect 25956 270 25971 278
rect 25905 258 25971 270
rect 21232 220 21252 226
rect 25886 220 25906 226
rect 21232 186 21244 220
rect 25894 186 25906 220
rect 21232 126 21252 186
rect 25886 126 25906 186
rect 21030 94 21100 100
rect 26040 94 26110 100
rect 21030 84 26110 94
rect 21030 46 21236 84
rect 25902 46 26110 84
rect 21030 30 26110 46
rect 30 -530 5110 -520
rect 30 -568 236 -530
rect 4959 -568 5110 -530
rect 30 -578 5110 -568
rect 30 -580 100 -578
rect 5040 -580 5110 -578
rect 232 -670 252 -610
rect 4886 -670 4906 -610
rect 232 -704 244 -670
rect 4894 -704 4906 -670
rect 232 -710 252 -704
rect 4886 -710 4906 -704
rect 165 -754 231 -742
rect 165 -762 182 -754
rect 216 -762 231 -754
rect 165 -6730 182 -6722
rect 216 -6730 231 -6722
rect 165 -6742 231 -6730
rect 323 -754 389 -742
rect 323 -762 340 -754
rect 374 -762 389 -754
rect 323 -6730 340 -6722
rect 374 -6730 389 -6722
rect 323 -6742 389 -6730
rect 481 -754 547 -742
rect 481 -762 498 -754
rect 532 -762 547 -754
rect 481 -6730 498 -6722
rect 532 -6730 547 -6722
rect 481 -6742 547 -6730
rect 639 -754 705 -742
rect 639 -762 656 -754
rect 690 -762 705 -754
rect 639 -6730 656 -6722
rect 690 -6730 705 -6722
rect 639 -6742 705 -6730
rect 797 -754 863 -742
rect 797 -762 814 -754
rect 848 -762 863 -754
rect 797 -6730 814 -6722
rect 848 -6730 863 -6722
rect 797 -6742 863 -6730
rect 955 -754 1021 -742
rect 955 -762 972 -754
rect 1006 -762 1021 -754
rect 955 -6730 972 -6722
rect 1006 -6730 1021 -6722
rect 955 -6742 1021 -6730
rect 1113 -754 1179 -742
rect 1113 -762 1130 -754
rect 1164 -762 1179 -754
rect 1113 -6730 1130 -6722
rect 1164 -6730 1179 -6722
rect 1113 -6742 1179 -6730
rect 1271 -754 1337 -742
rect 1271 -762 1288 -754
rect 1322 -762 1337 -754
rect 1271 -6730 1288 -6722
rect 1322 -6730 1337 -6722
rect 1271 -6742 1337 -6730
rect 1429 -754 1495 -742
rect 1429 -762 1446 -754
rect 1480 -762 1495 -754
rect 1429 -6730 1446 -6722
rect 1480 -6730 1495 -6722
rect 1429 -6742 1495 -6730
rect 1587 -754 1653 -742
rect 1587 -762 1604 -754
rect 1638 -762 1653 -754
rect 1587 -6730 1604 -6722
rect 1638 -6730 1653 -6722
rect 1587 -6742 1653 -6730
rect 1745 -754 1811 -742
rect 1745 -762 1762 -754
rect 1796 -762 1811 -754
rect 1745 -6730 1762 -6722
rect 1796 -6730 1811 -6722
rect 1745 -6742 1811 -6730
rect 1903 -754 1969 -742
rect 1903 -762 1920 -754
rect 1954 -762 1969 -754
rect 1903 -6730 1920 -6722
rect 1954 -6730 1969 -6722
rect 1903 -6742 1969 -6730
rect 2061 -754 2127 -742
rect 2061 -762 2078 -754
rect 2112 -762 2127 -754
rect 2061 -6730 2078 -6722
rect 2112 -6730 2127 -6722
rect 2061 -6742 2127 -6730
rect 2219 -754 2285 -742
rect 2219 -762 2236 -754
rect 2270 -762 2285 -754
rect 2219 -6730 2236 -6722
rect 2270 -6730 2285 -6722
rect 2219 -6742 2285 -6730
rect 2377 -754 2443 -742
rect 2377 -762 2394 -754
rect 2428 -762 2443 -754
rect 2377 -6730 2394 -6722
rect 2428 -6730 2443 -6722
rect 2377 -6742 2443 -6730
rect 2535 -754 2601 -742
rect 2535 -762 2552 -754
rect 2586 -762 2601 -754
rect 2535 -6730 2552 -6722
rect 2586 -6730 2601 -6722
rect 2535 -6742 2601 -6730
rect 2693 -754 2759 -742
rect 2693 -762 2710 -754
rect 2744 -762 2759 -754
rect 2693 -6730 2710 -6722
rect 2744 -6730 2759 -6722
rect 2693 -6742 2759 -6730
rect 2851 -754 2917 -742
rect 2851 -762 2868 -754
rect 2902 -762 2917 -754
rect 2851 -6730 2868 -6722
rect 2902 -6730 2917 -6722
rect 2851 -6742 2917 -6730
rect 3009 -754 3075 -742
rect 3009 -762 3026 -754
rect 3060 -762 3075 -754
rect 3009 -6730 3026 -6722
rect 3060 -6730 3075 -6722
rect 3009 -6742 3075 -6730
rect 3167 -754 3233 -742
rect 3167 -762 3184 -754
rect 3218 -762 3233 -754
rect 3167 -6730 3184 -6722
rect 3218 -6730 3233 -6722
rect 3167 -6742 3233 -6730
rect 3325 -754 3391 -742
rect 3325 -762 3342 -754
rect 3376 -762 3391 -754
rect 3325 -6730 3342 -6722
rect 3376 -6730 3391 -6722
rect 3325 -6742 3391 -6730
rect 3483 -754 3549 -742
rect 3483 -762 3500 -754
rect 3534 -762 3549 -754
rect 3483 -6730 3500 -6722
rect 3534 -6730 3549 -6722
rect 3483 -6742 3549 -6730
rect 3641 -754 3707 -742
rect 3641 -762 3658 -754
rect 3692 -762 3707 -754
rect 3641 -6730 3658 -6722
rect 3692 -6730 3707 -6722
rect 3641 -6742 3707 -6730
rect 3799 -754 3865 -742
rect 3799 -762 3816 -754
rect 3850 -762 3865 -754
rect 3799 -6730 3816 -6722
rect 3850 -6730 3865 -6722
rect 3799 -6742 3865 -6730
rect 3957 -754 4023 -742
rect 3957 -762 3974 -754
rect 4008 -762 4023 -754
rect 3957 -6730 3974 -6722
rect 4008 -6730 4023 -6722
rect 3957 -6742 4023 -6730
rect 4115 -754 4181 -742
rect 4115 -762 4132 -754
rect 4166 -762 4181 -754
rect 4115 -6730 4132 -6722
rect 4166 -6730 4181 -6722
rect 4115 -6742 4181 -6730
rect 4273 -754 4339 -742
rect 4273 -762 4290 -754
rect 4324 -762 4339 -754
rect 4273 -6730 4290 -6722
rect 4324 -6730 4339 -6722
rect 4273 -6742 4339 -6730
rect 4431 -754 4497 -742
rect 4431 -762 4448 -754
rect 4482 -762 4497 -754
rect 4431 -6730 4448 -6722
rect 4482 -6730 4497 -6722
rect 4431 -6742 4497 -6730
rect 4589 -754 4655 -742
rect 4589 -762 4606 -754
rect 4640 -762 4655 -754
rect 4589 -6730 4606 -6722
rect 4640 -6730 4655 -6722
rect 4589 -6742 4655 -6730
rect 4747 -754 4813 -742
rect 4747 -762 4764 -754
rect 4798 -762 4813 -754
rect 4747 -6730 4764 -6722
rect 4798 -6730 4813 -6722
rect 4747 -6742 4813 -6730
rect 4905 -754 4971 -742
rect 4905 -762 4922 -754
rect 4956 -762 4971 -754
rect 4905 -6730 4922 -6722
rect 4956 -6730 4971 -6722
rect 4905 -6742 4971 -6730
rect 232 -6780 252 -6774
rect 4886 -6780 4906 -6774
rect 232 -6814 244 -6780
rect 4894 -6814 4906 -6780
rect 232 -6874 252 -6814
rect 4886 -6874 4906 -6814
rect 30 -6906 100 -6900
rect 5040 -6906 5110 -6900
rect 30 -6916 5110 -6906
rect 30 -6954 236 -6916
rect 4902 -6954 5110 -6916
rect 30 -6970 5110 -6954
rect 7030 -530 12110 -520
rect 7030 -568 7236 -530
rect 11959 -568 12110 -530
rect 7030 -578 12110 -568
rect 7030 -580 7100 -578
rect 12040 -580 12110 -578
rect 7232 -670 7252 -610
rect 11886 -670 11906 -610
rect 7232 -704 7244 -670
rect 11894 -704 11906 -670
rect 7232 -710 7252 -704
rect 11886 -710 11906 -704
rect 7165 -754 7231 -742
rect 7165 -762 7182 -754
rect 7216 -762 7231 -754
rect 7165 -6730 7182 -6722
rect 7216 -6730 7231 -6722
rect 7165 -6742 7231 -6730
rect 7323 -754 7389 -742
rect 7323 -762 7340 -754
rect 7374 -762 7389 -754
rect 7323 -6730 7340 -6722
rect 7374 -6730 7389 -6722
rect 7323 -6742 7389 -6730
rect 7481 -754 7547 -742
rect 7481 -762 7498 -754
rect 7532 -762 7547 -754
rect 7481 -6730 7498 -6722
rect 7532 -6730 7547 -6722
rect 7481 -6742 7547 -6730
rect 7639 -754 7705 -742
rect 7639 -762 7656 -754
rect 7690 -762 7705 -754
rect 7639 -6730 7656 -6722
rect 7690 -6730 7705 -6722
rect 7639 -6742 7705 -6730
rect 7797 -754 7863 -742
rect 7797 -762 7814 -754
rect 7848 -762 7863 -754
rect 7797 -6730 7814 -6722
rect 7848 -6730 7863 -6722
rect 7797 -6742 7863 -6730
rect 7955 -754 8021 -742
rect 7955 -762 7972 -754
rect 8006 -762 8021 -754
rect 7955 -6730 7972 -6722
rect 8006 -6730 8021 -6722
rect 7955 -6742 8021 -6730
rect 8113 -754 8179 -742
rect 8113 -762 8130 -754
rect 8164 -762 8179 -754
rect 8113 -6730 8130 -6722
rect 8164 -6730 8179 -6722
rect 8113 -6742 8179 -6730
rect 8271 -754 8337 -742
rect 8271 -762 8288 -754
rect 8322 -762 8337 -754
rect 8271 -6730 8288 -6722
rect 8322 -6730 8337 -6722
rect 8271 -6742 8337 -6730
rect 8429 -754 8495 -742
rect 8429 -762 8446 -754
rect 8480 -762 8495 -754
rect 8429 -6730 8446 -6722
rect 8480 -6730 8495 -6722
rect 8429 -6742 8495 -6730
rect 8587 -754 8653 -742
rect 8587 -762 8604 -754
rect 8638 -762 8653 -754
rect 8587 -6730 8604 -6722
rect 8638 -6730 8653 -6722
rect 8587 -6742 8653 -6730
rect 8745 -754 8811 -742
rect 8745 -762 8762 -754
rect 8796 -762 8811 -754
rect 8745 -6730 8762 -6722
rect 8796 -6730 8811 -6722
rect 8745 -6742 8811 -6730
rect 8903 -754 8969 -742
rect 8903 -762 8920 -754
rect 8954 -762 8969 -754
rect 8903 -6730 8920 -6722
rect 8954 -6730 8969 -6722
rect 8903 -6742 8969 -6730
rect 9061 -754 9127 -742
rect 9061 -762 9078 -754
rect 9112 -762 9127 -754
rect 9061 -6730 9078 -6722
rect 9112 -6730 9127 -6722
rect 9061 -6742 9127 -6730
rect 9219 -754 9285 -742
rect 9219 -762 9236 -754
rect 9270 -762 9285 -754
rect 9219 -6730 9236 -6722
rect 9270 -6730 9285 -6722
rect 9219 -6742 9285 -6730
rect 9377 -754 9443 -742
rect 9377 -762 9394 -754
rect 9428 -762 9443 -754
rect 9377 -6730 9394 -6722
rect 9428 -6730 9443 -6722
rect 9377 -6742 9443 -6730
rect 9535 -754 9601 -742
rect 9535 -762 9552 -754
rect 9586 -762 9601 -754
rect 9535 -6730 9552 -6722
rect 9586 -6730 9601 -6722
rect 9535 -6742 9601 -6730
rect 9693 -754 9759 -742
rect 9693 -762 9710 -754
rect 9744 -762 9759 -754
rect 9693 -6730 9710 -6722
rect 9744 -6730 9759 -6722
rect 9693 -6742 9759 -6730
rect 9851 -754 9917 -742
rect 9851 -762 9868 -754
rect 9902 -762 9917 -754
rect 9851 -6730 9868 -6722
rect 9902 -6730 9917 -6722
rect 9851 -6742 9917 -6730
rect 10009 -754 10075 -742
rect 10009 -762 10026 -754
rect 10060 -762 10075 -754
rect 10009 -6730 10026 -6722
rect 10060 -6730 10075 -6722
rect 10009 -6742 10075 -6730
rect 10167 -754 10233 -742
rect 10167 -762 10184 -754
rect 10218 -762 10233 -754
rect 10167 -6730 10184 -6722
rect 10218 -6730 10233 -6722
rect 10167 -6742 10233 -6730
rect 10325 -754 10391 -742
rect 10325 -762 10342 -754
rect 10376 -762 10391 -754
rect 10325 -6730 10342 -6722
rect 10376 -6730 10391 -6722
rect 10325 -6742 10391 -6730
rect 10483 -754 10549 -742
rect 10483 -762 10500 -754
rect 10534 -762 10549 -754
rect 10483 -6730 10500 -6722
rect 10534 -6730 10549 -6722
rect 10483 -6742 10549 -6730
rect 10641 -754 10707 -742
rect 10641 -762 10658 -754
rect 10692 -762 10707 -754
rect 10641 -6730 10658 -6722
rect 10692 -6730 10707 -6722
rect 10641 -6742 10707 -6730
rect 10799 -754 10865 -742
rect 10799 -762 10816 -754
rect 10850 -762 10865 -754
rect 10799 -6730 10816 -6722
rect 10850 -6730 10865 -6722
rect 10799 -6742 10865 -6730
rect 10957 -754 11023 -742
rect 10957 -762 10974 -754
rect 11008 -762 11023 -754
rect 10957 -6730 10974 -6722
rect 11008 -6730 11023 -6722
rect 10957 -6742 11023 -6730
rect 11115 -754 11181 -742
rect 11115 -762 11132 -754
rect 11166 -762 11181 -754
rect 11115 -6730 11132 -6722
rect 11166 -6730 11181 -6722
rect 11115 -6742 11181 -6730
rect 11273 -754 11339 -742
rect 11273 -762 11290 -754
rect 11324 -762 11339 -754
rect 11273 -6730 11290 -6722
rect 11324 -6730 11339 -6722
rect 11273 -6742 11339 -6730
rect 11431 -754 11497 -742
rect 11431 -762 11448 -754
rect 11482 -762 11497 -754
rect 11431 -6730 11448 -6722
rect 11482 -6730 11497 -6722
rect 11431 -6742 11497 -6730
rect 11589 -754 11655 -742
rect 11589 -762 11606 -754
rect 11640 -762 11655 -754
rect 11589 -6730 11606 -6722
rect 11640 -6730 11655 -6722
rect 11589 -6742 11655 -6730
rect 11747 -754 11813 -742
rect 11747 -762 11764 -754
rect 11798 -762 11813 -754
rect 11747 -6730 11764 -6722
rect 11798 -6730 11813 -6722
rect 11747 -6742 11813 -6730
rect 11905 -754 11971 -742
rect 11905 -762 11922 -754
rect 11956 -762 11971 -754
rect 11905 -6730 11922 -6722
rect 11956 -6730 11971 -6722
rect 11905 -6742 11971 -6730
rect 7232 -6780 7252 -6774
rect 11886 -6780 11906 -6774
rect 7232 -6814 7244 -6780
rect 11894 -6814 11906 -6780
rect 7232 -6874 7252 -6814
rect 11886 -6874 11906 -6814
rect 7030 -6906 7100 -6900
rect 12040 -6906 12110 -6900
rect 7030 -6916 12110 -6906
rect 7030 -6954 7236 -6916
rect 11902 -6954 12110 -6916
rect 7030 -6970 12110 -6954
rect 14030 -530 19110 -520
rect 14030 -568 14236 -530
rect 18959 -568 19110 -530
rect 14030 -578 19110 -568
rect 14030 -580 14100 -578
rect 19040 -580 19110 -578
rect 14232 -670 14252 -610
rect 18886 -670 18906 -610
rect 14232 -704 14244 -670
rect 18894 -704 18906 -670
rect 14232 -710 14252 -704
rect 18886 -710 18906 -704
rect 14165 -754 14231 -742
rect 14165 -762 14182 -754
rect 14216 -762 14231 -754
rect 14165 -6730 14182 -6722
rect 14216 -6730 14231 -6722
rect 14165 -6742 14231 -6730
rect 14323 -754 14389 -742
rect 14323 -762 14340 -754
rect 14374 -762 14389 -754
rect 14323 -6730 14340 -6722
rect 14374 -6730 14389 -6722
rect 14323 -6742 14389 -6730
rect 14481 -754 14547 -742
rect 14481 -762 14498 -754
rect 14532 -762 14547 -754
rect 14481 -6730 14498 -6722
rect 14532 -6730 14547 -6722
rect 14481 -6742 14547 -6730
rect 14639 -754 14705 -742
rect 14639 -762 14656 -754
rect 14690 -762 14705 -754
rect 14639 -6730 14656 -6722
rect 14690 -6730 14705 -6722
rect 14639 -6742 14705 -6730
rect 14797 -754 14863 -742
rect 14797 -762 14814 -754
rect 14848 -762 14863 -754
rect 14797 -6730 14814 -6722
rect 14848 -6730 14863 -6722
rect 14797 -6742 14863 -6730
rect 14955 -754 15021 -742
rect 14955 -762 14972 -754
rect 15006 -762 15021 -754
rect 14955 -6730 14972 -6722
rect 15006 -6730 15021 -6722
rect 14955 -6742 15021 -6730
rect 15113 -754 15179 -742
rect 15113 -762 15130 -754
rect 15164 -762 15179 -754
rect 15113 -6730 15130 -6722
rect 15164 -6730 15179 -6722
rect 15113 -6742 15179 -6730
rect 15271 -754 15337 -742
rect 15271 -762 15288 -754
rect 15322 -762 15337 -754
rect 15271 -6730 15288 -6722
rect 15322 -6730 15337 -6722
rect 15271 -6742 15337 -6730
rect 15429 -754 15495 -742
rect 15429 -762 15446 -754
rect 15480 -762 15495 -754
rect 15429 -6730 15446 -6722
rect 15480 -6730 15495 -6722
rect 15429 -6742 15495 -6730
rect 15587 -754 15653 -742
rect 15587 -762 15604 -754
rect 15638 -762 15653 -754
rect 15587 -6730 15604 -6722
rect 15638 -6730 15653 -6722
rect 15587 -6742 15653 -6730
rect 15745 -754 15811 -742
rect 15745 -762 15762 -754
rect 15796 -762 15811 -754
rect 15745 -6730 15762 -6722
rect 15796 -6730 15811 -6722
rect 15745 -6742 15811 -6730
rect 15903 -754 15969 -742
rect 15903 -762 15920 -754
rect 15954 -762 15969 -754
rect 15903 -6730 15920 -6722
rect 15954 -6730 15969 -6722
rect 15903 -6742 15969 -6730
rect 16061 -754 16127 -742
rect 16061 -762 16078 -754
rect 16112 -762 16127 -754
rect 16061 -6730 16078 -6722
rect 16112 -6730 16127 -6722
rect 16061 -6742 16127 -6730
rect 16219 -754 16285 -742
rect 16219 -762 16236 -754
rect 16270 -762 16285 -754
rect 16219 -6730 16236 -6722
rect 16270 -6730 16285 -6722
rect 16219 -6742 16285 -6730
rect 16377 -754 16443 -742
rect 16377 -762 16394 -754
rect 16428 -762 16443 -754
rect 16377 -6730 16394 -6722
rect 16428 -6730 16443 -6722
rect 16377 -6742 16443 -6730
rect 16535 -754 16601 -742
rect 16535 -762 16552 -754
rect 16586 -762 16601 -754
rect 16535 -6730 16552 -6722
rect 16586 -6730 16601 -6722
rect 16535 -6742 16601 -6730
rect 16693 -754 16759 -742
rect 16693 -762 16710 -754
rect 16744 -762 16759 -754
rect 16693 -6730 16710 -6722
rect 16744 -6730 16759 -6722
rect 16693 -6742 16759 -6730
rect 16851 -754 16917 -742
rect 16851 -762 16868 -754
rect 16902 -762 16917 -754
rect 16851 -6730 16868 -6722
rect 16902 -6730 16917 -6722
rect 16851 -6742 16917 -6730
rect 17009 -754 17075 -742
rect 17009 -762 17026 -754
rect 17060 -762 17075 -754
rect 17009 -6730 17026 -6722
rect 17060 -6730 17075 -6722
rect 17009 -6742 17075 -6730
rect 17167 -754 17233 -742
rect 17167 -762 17184 -754
rect 17218 -762 17233 -754
rect 17167 -6730 17184 -6722
rect 17218 -6730 17233 -6722
rect 17167 -6742 17233 -6730
rect 17325 -754 17391 -742
rect 17325 -762 17342 -754
rect 17376 -762 17391 -754
rect 17325 -6730 17342 -6722
rect 17376 -6730 17391 -6722
rect 17325 -6742 17391 -6730
rect 17483 -754 17549 -742
rect 17483 -762 17500 -754
rect 17534 -762 17549 -754
rect 17483 -6730 17500 -6722
rect 17534 -6730 17549 -6722
rect 17483 -6742 17549 -6730
rect 17641 -754 17707 -742
rect 17641 -762 17658 -754
rect 17692 -762 17707 -754
rect 17641 -6730 17658 -6722
rect 17692 -6730 17707 -6722
rect 17641 -6742 17707 -6730
rect 17799 -754 17865 -742
rect 17799 -762 17816 -754
rect 17850 -762 17865 -754
rect 17799 -6730 17816 -6722
rect 17850 -6730 17865 -6722
rect 17799 -6742 17865 -6730
rect 17957 -754 18023 -742
rect 17957 -762 17974 -754
rect 18008 -762 18023 -754
rect 17957 -6730 17974 -6722
rect 18008 -6730 18023 -6722
rect 17957 -6742 18023 -6730
rect 18115 -754 18181 -742
rect 18115 -762 18132 -754
rect 18166 -762 18181 -754
rect 18115 -6730 18132 -6722
rect 18166 -6730 18181 -6722
rect 18115 -6742 18181 -6730
rect 18273 -754 18339 -742
rect 18273 -762 18290 -754
rect 18324 -762 18339 -754
rect 18273 -6730 18290 -6722
rect 18324 -6730 18339 -6722
rect 18273 -6742 18339 -6730
rect 18431 -754 18497 -742
rect 18431 -762 18448 -754
rect 18482 -762 18497 -754
rect 18431 -6730 18448 -6722
rect 18482 -6730 18497 -6722
rect 18431 -6742 18497 -6730
rect 18589 -754 18655 -742
rect 18589 -762 18606 -754
rect 18640 -762 18655 -754
rect 18589 -6730 18606 -6722
rect 18640 -6730 18655 -6722
rect 18589 -6742 18655 -6730
rect 18747 -754 18813 -742
rect 18747 -762 18764 -754
rect 18798 -762 18813 -754
rect 18747 -6730 18764 -6722
rect 18798 -6730 18813 -6722
rect 18747 -6742 18813 -6730
rect 18905 -754 18971 -742
rect 18905 -762 18922 -754
rect 18956 -762 18971 -754
rect 18905 -6730 18922 -6722
rect 18956 -6730 18971 -6722
rect 18905 -6742 18971 -6730
rect 14232 -6780 14252 -6774
rect 18886 -6780 18906 -6774
rect 14232 -6814 14244 -6780
rect 18894 -6814 18906 -6780
rect 14232 -6874 14252 -6814
rect 18886 -6874 18906 -6814
rect 14030 -6906 14100 -6900
rect 19040 -6906 19110 -6900
rect 14030 -6916 19110 -6906
rect 14030 -6954 14236 -6916
rect 18902 -6954 19110 -6916
rect 14030 -6970 19110 -6954
rect 21030 -530 26110 -520
rect 21030 -568 21236 -530
rect 25959 -568 26110 -530
rect 21030 -578 26110 -568
rect 21030 -580 21100 -578
rect 26040 -580 26110 -578
rect 21232 -670 21252 -610
rect 25886 -670 25906 -610
rect 21232 -704 21244 -670
rect 25894 -704 25906 -670
rect 21232 -710 21252 -704
rect 25886 -710 25906 -704
rect 21165 -754 21231 -742
rect 21165 -762 21182 -754
rect 21216 -762 21231 -754
rect 21165 -6730 21182 -6722
rect 21216 -6730 21231 -6722
rect 21165 -6742 21231 -6730
rect 21323 -754 21389 -742
rect 21323 -762 21340 -754
rect 21374 -762 21389 -754
rect 21323 -6730 21340 -6722
rect 21374 -6730 21389 -6722
rect 21323 -6742 21389 -6730
rect 21481 -754 21547 -742
rect 21481 -762 21498 -754
rect 21532 -762 21547 -754
rect 21481 -6730 21498 -6722
rect 21532 -6730 21547 -6722
rect 21481 -6742 21547 -6730
rect 21639 -754 21705 -742
rect 21639 -762 21656 -754
rect 21690 -762 21705 -754
rect 21639 -6730 21656 -6722
rect 21690 -6730 21705 -6722
rect 21639 -6742 21705 -6730
rect 21797 -754 21863 -742
rect 21797 -762 21814 -754
rect 21848 -762 21863 -754
rect 21797 -6730 21814 -6722
rect 21848 -6730 21863 -6722
rect 21797 -6742 21863 -6730
rect 21955 -754 22021 -742
rect 21955 -762 21972 -754
rect 22006 -762 22021 -754
rect 21955 -6730 21972 -6722
rect 22006 -6730 22021 -6722
rect 21955 -6742 22021 -6730
rect 22113 -754 22179 -742
rect 22113 -762 22130 -754
rect 22164 -762 22179 -754
rect 22113 -6730 22130 -6722
rect 22164 -6730 22179 -6722
rect 22113 -6742 22179 -6730
rect 22271 -754 22337 -742
rect 22271 -762 22288 -754
rect 22322 -762 22337 -754
rect 22271 -6730 22288 -6722
rect 22322 -6730 22337 -6722
rect 22271 -6742 22337 -6730
rect 22429 -754 22495 -742
rect 22429 -762 22446 -754
rect 22480 -762 22495 -754
rect 22429 -6730 22446 -6722
rect 22480 -6730 22495 -6722
rect 22429 -6742 22495 -6730
rect 22587 -754 22653 -742
rect 22587 -762 22604 -754
rect 22638 -762 22653 -754
rect 22587 -6730 22604 -6722
rect 22638 -6730 22653 -6722
rect 22587 -6742 22653 -6730
rect 22745 -754 22811 -742
rect 22745 -762 22762 -754
rect 22796 -762 22811 -754
rect 22745 -6730 22762 -6722
rect 22796 -6730 22811 -6722
rect 22745 -6742 22811 -6730
rect 22903 -754 22969 -742
rect 22903 -762 22920 -754
rect 22954 -762 22969 -754
rect 22903 -6730 22920 -6722
rect 22954 -6730 22969 -6722
rect 22903 -6742 22969 -6730
rect 23061 -754 23127 -742
rect 23061 -762 23078 -754
rect 23112 -762 23127 -754
rect 23061 -6730 23078 -6722
rect 23112 -6730 23127 -6722
rect 23061 -6742 23127 -6730
rect 23219 -754 23285 -742
rect 23219 -762 23236 -754
rect 23270 -762 23285 -754
rect 23219 -6730 23236 -6722
rect 23270 -6730 23285 -6722
rect 23219 -6742 23285 -6730
rect 23377 -754 23443 -742
rect 23377 -762 23394 -754
rect 23428 -762 23443 -754
rect 23377 -6730 23394 -6722
rect 23428 -6730 23443 -6722
rect 23377 -6742 23443 -6730
rect 23535 -754 23601 -742
rect 23535 -762 23552 -754
rect 23586 -762 23601 -754
rect 23535 -6730 23552 -6722
rect 23586 -6730 23601 -6722
rect 23535 -6742 23601 -6730
rect 23693 -754 23759 -742
rect 23693 -762 23710 -754
rect 23744 -762 23759 -754
rect 23693 -6730 23710 -6722
rect 23744 -6730 23759 -6722
rect 23693 -6742 23759 -6730
rect 23851 -754 23917 -742
rect 23851 -762 23868 -754
rect 23902 -762 23917 -754
rect 23851 -6730 23868 -6722
rect 23902 -6730 23917 -6722
rect 23851 -6742 23917 -6730
rect 24009 -754 24075 -742
rect 24009 -762 24026 -754
rect 24060 -762 24075 -754
rect 24009 -6730 24026 -6722
rect 24060 -6730 24075 -6722
rect 24009 -6742 24075 -6730
rect 24167 -754 24233 -742
rect 24167 -762 24184 -754
rect 24218 -762 24233 -754
rect 24167 -6730 24184 -6722
rect 24218 -6730 24233 -6722
rect 24167 -6742 24233 -6730
rect 24325 -754 24391 -742
rect 24325 -762 24342 -754
rect 24376 -762 24391 -754
rect 24325 -6730 24342 -6722
rect 24376 -6730 24391 -6722
rect 24325 -6742 24391 -6730
rect 24483 -754 24549 -742
rect 24483 -762 24500 -754
rect 24534 -762 24549 -754
rect 24483 -6730 24500 -6722
rect 24534 -6730 24549 -6722
rect 24483 -6742 24549 -6730
rect 24641 -754 24707 -742
rect 24641 -762 24658 -754
rect 24692 -762 24707 -754
rect 24641 -6730 24658 -6722
rect 24692 -6730 24707 -6722
rect 24641 -6742 24707 -6730
rect 24799 -754 24865 -742
rect 24799 -762 24816 -754
rect 24850 -762 24865 -754
rect 24799 -6730 24816 -6722
rect 24850 -6730 24865 -6722
rect 24799 -6742 24865 -6730
rect 24957 -754 25023 -742
rect 24957 -762 24974 -754
rect 25008 -762 25023 -754
rect 24957 -6730 24974 -6722
rect 25008 -6730 25023 -6722
rect 24957 -6742 25023 -6730
rect 25115 -754 25181 -742
rect 25115 -762 25132 -754
rect 25166 -762 25181 -754
rect 25115 -6730 25132 -6722
rect 25166 -6730 25181 -6722
rect 25115 -6742 25181 -6730
rect 25273 -754 25339 -742
rect 25273 -762 25290 -754
rect 25324 -762 25339 -754
rect 25273 -6730 25290 -6722
rect 25324 -6730 25339 -6722
rect 25273 -6742 25339 -6730
rect 25431 -754 25497 -742
rect 25431 -762 25448 -754
rect 25482 -762 25497 -754
rect 25431 -6730 25448 -6722
rect 25482 -6730 25497 -6722
rect 25431 -6742 25497 -6730
rect 25589 -754 25655 -742
rect 25589 -762 25606 -754
rect 25640 -762 25655 -754
rect 25589 -6730 25606 -6722
rect 25640 -6730 25655 -6722
rect 25589 -6742 25655 -6730
rect 25747 -754 25813 -742
rect 25747 -762 25764 -754
rect 25798 -762 25813 -754
rect 25747 -6730 25764 -6722
rect 25798 -6730 25813 -6722
rect 25747 -6742 25813 -6730
rect 25905 -754 25971 -742
rect 25905 -762 25922 -754
rect 25956 -762 25971 -754
rect 25905 -6730 25922 -6722
rect 25956 -6730 25971 -6722
rect 25905 -6742 25971 -6730
rect 21232 -6780 21252 -6774
rect 25886 -6780 25906 -6774
rect 21232 -6814 21244 -6780
rect 25894 -6814 25906 -6780
rect 21232 -6874 21252 -6814
rect 25886 -6874 25906 -6814
rect 21030 -6906 21100 -6900
rect 26040 -6906 26110 -6900
rect 21030 -6916 26110 -6906
rect 21030 -6954 21236 -6916
rect 25902 -6954 26110 -6916
rect 21030 -6970 26110 -6954
<< via1 >>
rect 30 6280 100 6420
rect 252 6330 4886 6390
rect 252 6296 312 6330
rect 312 6296 402 6330
rect 402 6296 470 6330
rect 470 6296 560 6330
rect 560 6296 628 6330
rect 628 6296 718 6330
rect 718 6296 786 6330
rect 786 6296 876 6330
rect 876 6296 944 6330
rect 944 6296 1034 6330
rect 1034 6296 1102 6330
rect 1102 6296 1192 6330
rect 1192 6296 1260 6330
rect 1260 6296 1350 6330
rect 1350 6296 1418 6330
rect 1418 6296 1508 6330
rect 1508 6296 1576 6330
rect 1576 6296 1666 6330
rect 1666 6296 1734 6330
rect 1734 6296 1824 6330
rect 1824 6296 1892 6330
rect 1892 6296 1982 6330
rect 1982 6296 2050 6330
rect 2050 6296 2140 6330
rect 2140 6296 2208 6330
rect 2208 6296 2298 6330
rect 2298 6296 2366 6330
rect 2366 6296 2456 6330
rect 2456 6296 2524 6330
rect 2524 6296 2614 6330
rect 2614 6296 2682 6330
rect 2682 6296 2772 6330
rect 2772 6296 2840 6330
rect 2840 6296 2930 6330
rect 2930 6296 2998 6330
rect 2998 6296 3088 6330
rect 3088 6296 3156 6330
rect 3156 6296 3246 6330
rect 3246 6296 3314 6330
rect 3314 6296 3404 6330
rect 3404 6296 3472 6330
rect 3472 6296 3562 6330
rect 3562 6296 3630 6330
rect 3630 6296 3720 6330
rect 3720 6296 3788 6330
rect 3788 6296 3878 6330
rect 3878 6296 3946 6330
rect 3946 6296 4036 6330
rect 4036 6296 4104 6330
rect 4104 6296 4194 6330
rect 4194 6296 4262 6330
rect 4262 6296 4352 6330
rect 4352 6296 4420 6330
rect 4420 6296 4510 6330
rect 4510 6296 4578 6330
rect 4578 6296 4668 6330
rect 4668 6296 4736 6330
rect 4736 6296 4826 6330
rect 4826 6296 4886 6330
rect 252 6290 4886 6296
rect 30 236 46 6280
rect 46 236 84 6280
rect 84 236 100 6280
rect 5040 6280 5110 6420
rect 165 278 182 6238
rect 182 278 216 6238
rect 216 278 231 6238
rect 323 278 340 6238
rect 340 278 374 6238
rect 374 278 389 6238
rect 481 278 498 6238
rect 498 278 532 6238
rect 532 278 547 6238
rect 639 278 656 6238
rect 656 278 690 6238
rect 690 278 705 6238
rect 797 278 814 6238
rect 814 278 848 6238
rect 848 278 863 6238
rect 955 278 972 6238
rect 972 278 1006 6238
rect 1006 278 1021 6238
rect 1113 278 1130 6238
rect 1130 278 1164 6238
rect 1164 278 1179 6238
rect 1271 278 1288 6238
rect 1288 278 1322 6238
rect 1322 278 1337 6238
rect 1429 278 1446 6238
rect 1446 278 1480 6238
rect 1480 278 1495 6238
rect 1587 278 1604 6238
rect 1604 278 1638 6238
rect 1638 278 1653 6238
rect 1745 278 1762 6238
rect 1762 278 1796 6238
rect 1796 278 1811 6238
rect 1903 278 1920 6238
rect 1920 278 1954 6238
rect 1954 278 1969 6238
rect 2061 278 2078 6238
rect 2078 278 2112 6238
rect 2112 278 2127 6238
rect 2219 278 2236 6238
rect 2236 278 2270 6238
rect 2270 278 2285 6238
rect 2377 278 2394 6238
rect 2394 278 2428 6238
rect 2428 278 2443 6238
rect 2535 278 2552 6238
rect 2552 278 2586 6238
rect 2586 278 2601 6238
rect 2693 278 2710 6238
rect 2710 278 2744 6238
rect 2744 278 2759 6238
rect 2851 278 2868 6238
rect 2868 278 2902 6238
rect 2902 278 2917 6238
rect 3009 278 3026 6238
rect 3026 278 3060 6238
rect 3060 278 3075 6238
rect 3167 278 3184 6238
rect 3184 278 3218 6238
rect 3218 278 3233 6238
rect 3325 278 3342 6238
rect 3342 278 3376 6238
rect 3376 278 3391 6238
rect 3483 278 3500 6238
rect 3500 278 3534 6238
rect 3534 278 3549 6238
rect 3641 278 3658 6238
rect 3658 278 3692 6238
rect 3692 278 3707 6238
rect 3799 278 3816 6238
rect 3816 278 3850 6238
rect 3850 278 3865 6238
rect 3957 278 3974 6238
rect 3974 278 4008 6238
rect 4008 278 4023 6238
rect 4115 278 4132 6238
rect 4132 278 4166 6238
rect 4166 278 4181 6238
rect 4273 278 4290 6238
rect 4290 278 4324 6238
rect 4324 278 4339 6238
rect 4431 278 4448 6238
rect 4448 278 4482 6238
rect 4482 278 4497 6238
rect 4589 278 4606 6238
rect 4606 278 4640 6238
rect 4640 278 4655 6238
rect 4747 278 4764 6238
rect 4764 278 4798 6238
rect 4798 278 4813 6238
rect 4905 278 4922 6238
rect 4922 278 4956 6238
rect 4956 278 4971 6238
rect 30 100 100 236
rect 5040 236 5054 6280
rect 5054 236 5092 6280
rect 5092 236 5110 6280
rect 252 220 4886 226
rect 252 186 312 220
rect 312 186 402 220
rect 402 186 470 220
rect 470 186 560 220
rect 560 186 628 220
rect 628 186 718 220
rect 718 186 786 220
rect 786 186 876 220
rect 876 186 944 220
rect 944 186 1034 220
rect 1034 186 1102 220
rect 1102 186 1192 220
rect 1192 186 1260 220
rect 1260 186 1350 220
rect 1350 186 1418 220
rect 1418 186 1508 220
rect 1508 186 1576 220
rect 1576 186 1666 220
rect 1666 186 1734 220
rect 1734 186 1824 220
rect 1824 186 1892 220
rect 1892 186 1982 220
rect 1982 186 2050 220
rect 2050 186 2140 220
rect 2140 186 2208 220
rect 2208 186 2298 220
rect 2298 186 2366 220
rect 2366 186 2456 220
rect 2456 186 2524 220
rect 2524 186 2614 220
rect 2614 186 2682 220
rect 2682 186 2772 220
rect 2772 186 2840 220
rect 2840 186 2930 220
rect 2930 186 2998 220
rect 2998 186 3088 220
rect 3088 186 3156 220
rect 3156 186 3246 220
rect 3246 186 3314 220
rect 3314 186 3404 220
rect 3404 186 3472 220
rect 3472 186 3562 220
rect 3562 186 3630 220
rect 3630 186 3720 220
rect 3720 186 3788 220
rect 3788 186 3878 220
rect 3878 186 3946 220
rect 3946 186 4036 220
rect 4036 186 4104 220
rect 4104 186 4194 220
rect 4194 186 4262 220
rect 4262 186 4352 220
rect 4352 186 4420 220
rect 4420 186 4510 220
rect 4510 186 4578 220
rect 4578 186 4668 220
rect 4668 186 4736 220
rect 4736 186 4826 220
rect 4826 186 4886 220
rect 252 126 4886 186
rect 5040 100 5110 236
rect 7030 6280 7100 6420
rect 7252 6330 11886 6390
rect 7252 6296 7312 6330
rect 7312 6296 7402 6330
rect 7402 6296 7470 6330
rect 7470 6296 7560 6330
rect 7560 6296 7628 6330
rect 7628 6296 7718 6330
rect 7718 6296 7786 6330
rect 7786 6296 7876 6330
rect 7876 6296 7944 6330
rect 7944 6296 8034 6330
rect 8034 6296 8102 6330
rect 8102 6296 8192 6330
rect 8192 6296 8260 6330
rect 8260 6296 8350 6330
rect 8350 6296 8418 6330
rect 8418 6296 8508 6330
rect 8508 6296 8576 6330
rect 8576 6296 8666 6330
rect 8666 6296 8734 6330
rect 8734 6296 8824 6330
rect 8824 6296 8892 6330
rect 8892 6296 8982 6330
rect 8982 6296 9050 6330
rect 9050 6296 9140 6330
rect 9140 6296 9208 6330
rect 9208 6296 9298 6330
rect 9298 6296 9366 6330
rect 9366 6296 9456 6330
rect 9456 6296 9524 6330
rect 9524 6296 9614 6330
rect 9614 6296 9682 6330
rect 9682 6296 9772 6330
rect 9772 6296 9840 6330
rect 9840 6296 9930 6330
rect 9930 6296 9998 6330
rect 9998 6296 10088 6330
rect 10088 6296 10156 6330
rect 10156 6296 10246 6330
rect 10246 6296 10314 6330
rect 10314 6296 10404 6330
rect 10404 6296 10472 6330
rect 10472 6296 10562 6330
rect 10562 6296 10630 6330
rect 10630 6296 10720 6330
rect 10720 6296 10788 6330
rect 10788 6296 10878 6330
rect 10878 6296 10946 6330
rect 10946 6296 11036 6330
rect 11036 6296 11104 6330
rect 11104 6296 11194 6330
rect 11194 6296 11262 6330
rect 11262 6296 11352 6330
rect 11352 6296 11420 6330
rect 11420 6296 11510 6330
rect 11510 6296 11578 6330
rect 11578 6296 11668 6330
rect 11668 6296 11736 6330
rect 11736 6296 11826 6330
rect 11826 6296 11886 6330
rect 7252 6290 11886 6296
rect 7030 236 7046 6280
rect 7046 236 7084 6280
rect 7084 236 7100 6280
rect 12040 6280 12110 6420
rect 7165 278 7182 6238
rect 7182 278 7216 6238
rect 7216 278 7231 6238
rect 7323 278 7340 6238
rect 7340 278 7374 6238
rect 7374 278 7389 6238
rect 7481 278 7498 6238
rect 7498 278 7532 6238
rect 7532 278 7547 6238
rect 7639 278 7656 6238
rect 7656 278 7690 6238
rect 7690 278 7705 6238
rect 7797 278 7814 6238
rect 7814 278 7848 6238
rect 7848 278 7863 6238
rect 7955 278 7972 6238
rect 7972 278 8006 6238
rect 8006 278 8021 6238
rect 8113 278 8130 6238
rect 8130 278 8164 6238
rect 8164 278 8179 6238
rect 8271 278 8288 6238
rect 8288 278 8322 6238
rect 8322 278 8337 6238
rect 8429 278 8446 6238
rect 8446 278 8480 6238
rect 8480 278 8495 6238
rect 8587 278 8604 6238
rect 8604 278 8638 6238
rect 8638 278 8653 6238
rect 8745 278 8762 6238
rect 8762 278 8796 6238
rect 8796 278 8811 6238
rect 8903 278 8920 6238
rect 8920 278 8954 6238
rect 8954 278 8969 6238
rect 9061 278 9078 6238
rect 9078 278 9112 6238
rect 9112 278 9127 6238
rect 9219 278 9236 6238
rect 9236 278 9270 6238
rect 9270 278 9285 6238
rect 9377 278 9394 6238
rect 9394 278 9428 6238
rect 9428 278 9443 6238
rect 9535 278 9552 6238
rect 9552 278 9586 6238
rect 9586 278 9601 6238
rect 9693 278 9710 6238
rect 9710 278 9744 6238
rect 9744 278 9759 6238
rect 9851 278 9868 6238
rect 9868 278 9902 6238
rect 9902 278 9917 6238
rect 10009 278 10026 6238
rect 10026 278 10060 6238
rect 10060 278 10075 6238
rect 10167 278 10184 6238
rect 10184 278 10218 6238
rect 10218 278 10233 6238
rect 10325 278 10342 6238
rect 10342 278 10376 6238
rect 10376 278 10391 6238
rect 10483 278 10500 6238
rect 10500 278 10534 6238
rect 10534 278 10549 6238
rect 10641 278 10658 6238
rect 10658 278 10692 6238
rect 10692 278 10707 6238
rect 10799 278 10816 6238
rect 10816 278 10850 6238
rect 10850 278 10865 6238
rect 10957 278 10974 6238
rect 10974 278 11008 6238
rect 11008 278 11023 6238
rect 11115 278 11132 6238
rect 11132 278 11166 6238
rect 11166 278 11181 6238
rect 11273 278 11290 6238
rect 11290 278 11324 6238
rect 11324 278 11339 6238
rect 11431 278 11448 6238
rect 11448 278 11482 6238
rect 11482 278 11497 6238
rect 11589 278 11606 6238
rect 11606 278 11640 6238
rect 11640 278 11655 6238
rect 11747 278 11764 6238
rect 11764 278 11798 6238
rect 11798 278 11813 6238
rect 11905 278 11922 6238
rect 11922 278 11956 6238
rect 11956 278 11971 6238
rect 7030 100 7100 236
rect 12040 236 12054 6280
rect 12054 236 12092 6280
rect 12092 236 12110 6280
rect 7252 220 11886 226
rect 7252 186 7312 220
rect 7312 186 7402 220
rect 7402 186 7470 220
rect 7470 186 7560 220
rect 7560 186 7628 220
rect 7628 186 7718 220
rect 7718 186 7786 220
rect 7786 186 7876 220
rect 7876 186 7944 220
rect 7944 186 8034 220
rect 8034 186 8102 220
rect 8102 186 8192 220
rect 8192 186 8260 220
rect 8260 186 8350 220
rect 8350 186 8418 220
rect 8418 186 8508 220
rect 8508 186 8576 220
rect 8576 186 8666 220
rect 8666 186 8734 220
rect 8734 186 8824 220
rect 8824 186 8892 220
rect 8892 186 8982 220
rect 8982 186 9050 220
rect 9050 186 9140 220
rect 9140 186 9208 220
rect 9208 186 9298 220
rect 9298 186 9366 220
rect 9366 186 9456 220
rect 9456 186 9524 220
rect 9524 186 9614 220
rect 9614 186 9682 220
rect 9682 186 9772 220
rect 9772 186 9840 220
rect 9840 186 9930 220
rect 9930 186 9998 220
rect 9998 186 10088 220
rect 10088 186 10156 220
rect 10156 186 10246 220
rect 10246 186 10314 220
rect 10314 186 10404 220
rect 10404 186 10472 220
rect 10472 186 10562 220
rect 10562 186 10630 220
rect 10630 186 10720 220
rect 10720 186 10788 220
rect 10788 186 10878 220
rect 10878 186 10946 220
rect 10946 186 11036 220
rect 11036 186 11104 220
rect 11104 186 11194 220
rect 11194 186 11262 220
rect 11262 186 11352 220
rect 11352 186 11420 220
rect 11420 186 11510 220
rect 11510 186 11578 220
rect 11578 186 11668 220
rect 11668 186 11736 220
rect 11736 186 11826 220
rect 11826 186 11886 220
rect 7252 126 11886 186
rect 12040 100 12110 236
rect 14030 6280 14100 6420
rect 14252 6330 18886 6390
rect 14252 6296 14312 6330
rect 14312 6296 14402 6330
rect 14402 6296 14470 6330
rect 14470 6296 14560 6330
rect 14560 6296 14628 6330
rect 14628 6296 14718 6330
rect 14718 6296 14786 6330
rect 14786 6296 14876 6330
rect 14876 6296 14944 6330
rect 14944 6296 15034 6330
rect 15034 6296 15102 6330
rect 15102 6296 15192 6330
rect 15192 6296 15260 6330
rect 15260 6296 15350 6330
rect 15350 6296 15418 6330
rect 15418 6296 15508 6330
rect 15508 6296 15576 6330
rect 15576 6296 15666 6330
rect 15666 6296 15734 6330
rect 15734 6296 15824 6330
rect 15824 6296 15892 6330
rect 15892 6296 15982 6330
rect 15982 6296 16050 6330
rect 16050 6296 16140 6330
rect 16140 6296 16208 6330
rect 16208 6296 16298 6330
rect 16298 6296 16366 6330
rect 16366 6296 16456 6330
rect 16456 6296 16524 6330
rect 16524 6296 16614 6330
rect 16614 6296 16682 6330
rect 16682 6296 16772 6330
rect 16772 6296 16840 6330
rect 16840 6296 16930 6330
rect 16930 6296 16998 6330
rect 16998 6296 17088 6330
rect 17088 6296 17156 6330
rect 17156 6296 17246 6330
rect 17246 6296 17314 6330
rect 17314 6296 17404 6330
rect 17404 6296 17472 6330
rect 17472 6296 17562 6330
rect 17562 6296 17630 6330
rect 17630 6296 17720 6330
rect 17720 6296 17788 6330
rect 17788 6296 17878 6330
rect 17878 6296 17946 6330
rect 17946 6296 18036 6330
rect 18036 6296 18104 6330
rect 18104 6296 18194 6330
rect 18194 6296 18262 6330
rect 18262 6296 18352 6330
rect 18352 6296 18420 6330
rect 18420 6296 18510 6330
rect 18510 6296 18578 6330
rect 18578 6296 18668 6330
rect 18668 6296 18736 6330
rect 18736 6296 18826 6330
rect 18826 6296 18886 6330
rect 14252 6290 18886 6296
rect 14030 236 14046 6280
rect 14046 236 14084 6280
rect 14084 236 14100 6280
rect 19040 6280 19110 6420
rect 14165 278 14182 6238
rect 14182 278 14216 6238
rect 14216 278 14231 6238
rect 14323 278 14340 6238
rect 14340 278 14374 6238
rect 14374 278 14389 6238
rect 14481 278 14498 6238
rect 14498 278 14532 6238
rect 14532 278 14547 6238
rect 14639 278 14656 6238
rect 14656 278 14690 6238
rect 14690 278 14705 6238
rect 14797 278 14814 6238
rect 14814 278 14848 6238
rect 14848 278 14863 6238
rect 14955 278 14972 6238
rect 14972 278 15006 6238
rect 15006 278 15021 6238
rect 15113 278 15130 6238
rect 15130 278 15164 6238
rect 15164 278 15179 6238
rect 15271 278 15288 6238
rect 15288 278 15322 6238
rect 15322 278 15337 6238
rect 15429 278 15446 6238
rect 15446 278 15480 6238
rect 15480 278 15495 6238
rect 15587 278 15604 6238
rect 15604 278 15638 6238
rect 15638 278 15653 6238
rect 15745 278 15762 6238
rect 15762 278 15796 6238
rect 15796 278 15811 6238
rect 15903 278 15920 6238
rect 15920 278 15954 6238
rect 15954 278 15969 6238
rect 16061 278 16078 6238
rect 16078 278 16112 6238
rect 16112 278 16127 6238
rect 16219 278 16236 6238
rect 16236 278 16270 6238
rect 16270 278 16285 6238
rect 16377 278 16394 6238
rect 16394 278 16428 6238
rect 16428 278 16443 6238
rect 16535 278 16552 6238
rect 16552 278 16586 6238
rect 16586 278 16601 6238
rect 16693 278 16710 6238
rect 16710 278 16744 6238
rect 16744 278 16759 6238
rect 16851 278 16868 6238
rect 16868 278 16902 6238
rect 16902 278 16917 6238
rect 17009 278 17026 6238
rect 17026 278 17060 6238
rect 17060 278 17075 6238
rect 17167 278 17184 6238
rect 17184 278 17218 6238
rect 17218 278 17233 6238
rect 17325 278 17342 6238
rect 17342 278 17376 6238
rect 17376 278 17391 6238
rect 17483 278 17500 6238
rect 17500 278 17534 6238
rect 17534 278 17549 6238
rect 17641 278 17658 6238
rect 17658 278 17692 6238
rect 17692 278 17707 6238
rect 17799 278 17816 6238
rect 17816 278 17850 6238
rect 17850 278 17865 6238
rect 17957 278 17974 6238
rect 17974 278 18008 6238
rect 18008 278 18023 6238
rect 18115 278 18132 6238
rect 18132 278 18166 6238
rect 18166 278 18181 6238
rect 18273 278 18290 6238
rect 18290 278 18324 6238
rect 18324 278 18339 6238
rect 18431 278 18448 6238
rect 18448 278 18482 6238
rect 18482 278 18497 6238
rect 18589 278 18606 6238
rect 18606 278 18640 6238
rect 18640 278 18655 6238
rect 18747 278 18764 6238
rect 18764 278 18798 6238
rect 18798 278 18813 6238
rect 18905 278 18922 6238
rect 18922 278 18956 6238
rect 18956 278 18971 6238
rect 14030 100 14100 236
rect 19040 236 19054 6280
rect 19054 236 19092 6280
rect 19092 236 19110 6280
rect 14252 220 18886 226
rect 14252 186 14312 220
rect 14312 186 14402 220
rect 14402 186 14470 220
rect 14470 186 14560 220
rect 14560 186 14628 220
rect 14628 186 14718 220
rect 14718 186 14786 220
rect 14786 186 14876 220
rect 14876 186 14944 220
rect 14944 186 15034 220
rect 15034 186 15102 220
rect 15102 186 15192 220
rect 15192 186 15260 220
rect 15260 186 15350 220
rect 15350 186 15418 220
rect 15418 186 15508 220
rect 15508 186 15576 220
rect 15576 186 15666 220
rect 15666 186 15734 220
rect 15734 186 15824 220
rect 15824 186 15892 220
rect 15892 186 15982 220
rect 15982 186 16050 220
rect 16050 186 16140 220
rect 16140 186 16208 220
rect 16208 186 16298 220
rect 16298 186 16366 220
rect 16366 186 16456 220
rect 16456 186 16524 220
rect 16524 186 16614 220
rect 16614 186 16682 220
rect 16682 186 16772 220
rect 16772 186 16840 220
rect 16840 186 16930 220
rect 16930 186 16998 220
rect 16998 186 17088 220
rect 17088 186 17156 220
rect 17156 186 17246 220
rect 17246 186 17314 220
rect 17314 186 17404 220
rect 17404 186 17472 220
rect 17472 186 17562 220
rect 17562 186 17630 220
rect 17630 186 17720 220
rect 17720 186 17788 220
rect 17788 186 17878 220
rect 17878 186 17946 220
rect 17946 186 18036 220
rect 18036 186 18104 220
rect 18104 186 18194 220
rect 18194 186 18262 220
rect 18262 186 18352 220
rect 18352 186 18420 220
rect 18420 186 18510 220
rect 18510 186 18578 220
rect 18578 186 18668 220
rect 18668 186 18736 220
rect 18736 186 18826 220
rect 18826 186 18886 220
rect 14252 126 18886 186
rect 19040 100 19110 236
rect 21030 6280 21100 6420
rect 21252 6330 25886 6390
rect 21252 6296 21312 6330
rect 21312 6296 21402 6330
rect 21402 6296 21470 6330
rect 21470 6296 21560 6330
rect 21560 6296 21628 6330
rect 21628 6296 21718 6330
rect 21718 6296 21786 6330
rect 21786 6296 21876 6330
rect 21876 6296 21944 6330
rect 21944 6296 22034 6330
rect 22034 6296 22102 6330
rect 22102 6296 22192 6330
rect 22192 6296 22260 6330
rect 22260 6296 22350 6330
rect 22350 6296 22418 6330
rect 22418 6296 22508 6330
rect 22508 6296 22576 6330
rect 22576 6296 22666 6330
rect 22666 6296 22734 6330
rect 22734 6296 22824 6330
rect 22824 6296 22892 6330
rect 22892 6296 22982 6330
rect 22982 6296 23050 6330
rect 23050 6296 23140 6330
rect 23140 6296 23208 6330
rect 23208 6296 23298 6330
rect 23298 6296 23366 6330
rect 23366 6296 23456 6330
rect 23456 6296 23524 6330
rect 23524 6296 23614 6330
rect 23614 6296 23682 6330
rect 23682 6296 23772 6330
rect 23772 6296 23840 6330
rect 23840 6296 23930 6330
rect 23930 6296 23998 6330
rect 23998 6296 24088 6330
rect 24088 6296 24156 6330
rect 24156 6296 24246 6330
rect 24246 6296 24314 6330
rect 24314 6296 24404 6330
rect 24404 6296 24472 6330
rect 24472 6296 24562 6330
rect 24562 6296 24630 6330
rect 24630 6296 24720 6330
rect 24720 6296 24788 6330
rect 24788 6296 24878 6330
rect 24878 6296 24946 6330
rect 24946 6296 25036 6330
rect 25036 6296 25104 6330
rect 25104 6296 25194 6330
rect 25194 6296 25262 6330
rect 25262 6296 25352 6330
rect 25352 6296 25420 6330
rect 25420 6296 25510 6330
rect 25510 6296 25578 6330
rect 25578 6296 25668 6330
rect 25668 6296 25736 6330
rect 25736 6296 25826 6330
rect 25826 6296 25886 6330
rect 21252 6290 25886 6296
rect 21030 236 21046 6280
rect 21046 236 21084 6280
rect 21084 236 21100 6280
rect 26040 6280 26110 6420
rect 21165 278 21182 6238
rect 21182 278 21216 6238
rect 21216 278 21231 6238
rect 21323 278 21340 6238
rect 21340 278 21374 6238
rect 21374 278 21389 6238
rect 21481 278 21498 6238
rect 21498 278 21532 6238
rect 21532 278 21547 6238
rect 21639 278 21656 6238
rect 21656 278 21690 6238
rect 21690 278 21705 6238
rect 21797 278 21814 6238
rect 21814 278 21848 6238
rect 21848 278 21863 6238
rect 21955 278 21972 6238
rect 21972 278 22006 6238
rect 22006 278 22021 6238
rect 22113 278 22130 6238
rect 22130 278 22164 6238
rect 22164 278 22179 6238
rect 22271 278 22288 6238
rect 22288 278 22322 6238
rect 22322 278 22337 6238
rect 22429 278 22446 6238
rect 22446 278 22480 6238
rect 22480 278 22495 6238
rect 22587 278 22604 6238
rect 22604 278 22638 6238
rect 22638 278 22653 6238
rect 22745 278 22762 6238
rect 22762 278 22796 6238
rect 22796 278 22811 6238
rect 22903 278 22920 6238
rect 22920 278 22954 6238
rect 22954 278 22969 6238
rect 23061 278 23078 6238
rect 23078 278 23112 6238
rect 23112 278 23127 6238
rect 23219 278 23236 6238
rect 23236 278 23270 6238
rect 23270 278 23285 6238
rect 23377 278 23394 6238
rect 23394 278 23428 6238
rect 23428 278 23443 6238
rect 23535 278 23552 6238
rect 23552 278 23586 6238
rect 23586 278 23601 6238
rect 23693 278 23710 6238
rect 23710 278 23744 6238
rect 23744 278 23759 6238
rect 23851 278 23868 6238
rect 23868 278 23902 6238
rect 23902 278 23917 6238
rect 24009 278 24026 6238
rect 24026 278 24060 6238
rect 24060 278 24075 6238
rect 24167 278 24184 6238
rect 24184 278 24218 6238
rect 24218 278 24233 6238
rect 24325 278 24342 6238
rect 24342 278 24376 6238
rect 24376 278 24391 6238
rect 24483 278 24500 6238
rect 24500 278 24534 6238
rect 24534 278 24549 6238
rect 24641 278 24658 6238
rect 24658 278 24692 6238
rect 24692 278 24707 6238
rect 24799 278 24816 6238
rect 24816 278 24850 6238
rect 24850 278 24865 6238
rect 24957 278 24974 6238
rect 24974 278 25008 6238
rect 25008 278 25023 6238
rect 25115 278 25132 6238
rect 25132 278 25166 6238
rect 25166 278 25181 6238
rect 25273 278 25290 6238
rect 25290 278 25324 6238
rect 25324 278 25339 6238
rect 25431 278 25448 6238
rect 25448 278 25482 6238
rect 25482 278 25497 6238
rect 25589 278 25606 6238
rect 25606 278 25640 6238
rect 25640 278 25655 6238
rect 25747 278 25764 6238
rect 25764 278 25798 6238
rect 25798 278 25813 6238
rect 25905 278 25922 6238
rect 25922 278 25956 6238
rect 25956 278 25971 6238
rect 21030 100 21100 236
rect 26040 236 26054 6280
rect 26054 236 26092 6280
rect 26092 236 26110 6280
rect 21252 220 25886 226
rect 21252 186 21312 220
rect 21312 186 21402 220
rect 21402 186 21470 220
rect 21470 186 21560 220
rect 21560 186 21628 220
rect 21628 186 21718 220
rect 21718 186 21786 220
rect 21786 186 21876 220
rect 21876 186 21944 220
rect 21944 186 22034 220
rect 22034 186 22102 220
rect 22102 186 22192 220
rect 22192 186 22260 220
rect 22260 186 22350 220
rect 22350 186 22418 220
rect 22418 186 22508 220
rect 22508 186 22576 220
rect 22576 186 22666 220
rect 22666 186 22734 220
rect 22734 186 22824 220
rect 22824 186 22892 220
rect 22892 186 22982 220
rect 22982 186 23050 220
rect 23050 186 23140 220
rect 23140 186 23208 220
rect 23208 186 23298 220
rect 23298 186 23366 220
rect 23366 186 23456 220
rect 23456 186 23524 220
rect 23524 186 23614 220
rect 23614 186 23682 220
rect 23682 186 23772 220
rect 23772 186 23840 220
rect 23840 186 23930 220
rect 23930 186 23998 220
rect 23998 186 24088 220
rect 24088 186 24156 220
rect 24156 186 24246 220
rect 24246 186 24314 220
rect 24314 186 24404 220
rect 24404 186 24472 220
rect 24472 186 24562 220
rect 24562 186 24630 220
rect 24630 186 24720 220
rect 24720 186 24788 220
rect 24788 186 24878 220
rect 24878 186 24946 220
rect 24946 186 25036 220
rect 25036 186 25104 220
rect 25104 186 25194 220
rect 25194 186 25262 220
rect 25262 186 25352 220
rect 25352 186 25420 220
rect 25420 186 25510 220
rect 25510 186 25578 220
rect 25578 186 25668 220
rect 25668 186 25736 220
rect 25736 186 25826 220
rect 25826 186 25886 220
rect 21252 126 25886 186
rect 26040 100 26110 236
rect 30 -720 100 -580
rect 252 -670 4886 -610
rect 252 -704 312 -670
rect 312 -704 402 -670
rect 402 -704 470 -670
rect 470 -704 560 -670
rect 560 -704 628 -670
rect 628 -704 718 -670
rect 718 -704 786 -670
rect 786 -704 876 -670
rect 876 -704 944 -670
rect 944 -704 1034 -670
rect 1034 -704 1102 -670
rect 1102 -704 1192 -670
rect 1192 -704 1260 -670
rect 1260 -704 1350 -670
rect 1350 -704 1418 -670
rect 1418 -704 1508 -670
rect 1508 -704 1576 -670
rect 1576 -704 1666 -670
rect 1666 -704 1734 -670
rect 1734 -704 1824 -670
rect 1824 -704 1892 -670
rect 1892 -704 1982 -670
rect 1982 -704 2050 -670
rect 2050 -704 2140 -670
rect 2140 -704 2208 -670
rect 2208 -704 2298 -670
rect 2298 -704 2366 -670
rect 2366 -704 2456 -670
rect 2456 -704 2524 -670
rect 2524 -704 2614 -670
rect 2614 -704 2682 -670
rect 2682 -704 2772 -670
rect 2772 -704 2840 -670
rect 2840 -704 2930 -670
rect 2930 -704 2998 -670
rect 2998 -704 3088 -670
rect 3088 -704 3156 -670
rect 3156 -704 3246 -670
rect 3246 -704 3314 -670
rect 3314 -704 3404 -670
rect 3404 -704 3472 -670
rect 3472 -704 3562 -670
rect 3562 -704 3630 -670
rect 3630 -704 3720 -670
rect 3720 -704 3788 -670
rect 3788 -704 3878 -670
rect 3878 -704 3946 -670
rect 3946 -704 4036 -670
rect 4036 -704 4104 -670
rect 4104 -704 4194 -670
rect 4194 -704 4262 -670
rect 4262 -704 4352 -670
rect 4352 -704 4420 -670
rect 4420 -704 4510 -670
rect 4510 -704 4578 -670
rect 4578 -704 4668 -670
rect 4668 -704 4736 -670
rect 4736 -704 4826 -670
rect 4826 -704 4886 -670
rect 252 -710 4886 -704
rect 30 -6764 46 -720
rect 46 -6764 84 -720
rect 84 -6764 100 -720
rect 5040 -720 5110 -580
rect 165 -6722 182 -762
rect 182 -6722 216 -762
rect 216 -6722 231 -762
rect 323 -6722 340 -762
rect 340 -6722 374 -762
rect 374 -6722 389 -762
rect 481 -6722 498 -762
rect 498 -6722 532 -762
rect 532 -6722 547 -762
rect 639 -6722 656 -762
rect 656 -6722 690 -762
rect 690 -6722 705 -762
rect 797 -6722 814 -762
rect 814 -6722 848 -762
rect 848 -6722 863 -762
rect 955 -6722 972 -762
rect 972 -6722 1006 -762
rect 1006 -6722 1021 -762
rect 1113 -6722 1130 -762
rect 1130 -6722 1164 -762
rect 1164 -6722 1179 -762
rect 1271 -6722 1288 -762
rect 1288 -6722 1322 -762
rect 1322 -6722 1337 -762
rect 1429 -6722 1446 -762
rect 1446 -6722 1480 -762
rect 1480 -6722 1495 -762
rect 1587 -6722 1604 -762
rect 1604 -6722 1638 -762
rect 1638 -6722 1653 -762
rect 1745 -6722 1762 -762
rect 1762 -6722 1796 -762
rect 1796 -6722 1811 -762
rect 1903 -6722 1920 -762
rect 1920 -6722 1954 -762
rect 1954 -6722 1969 -762
rect 2061 -6722 2078 -762
rect 2078 -6722 2112 -762
rect 2112 -6722 2127 -762
rect 2219 -6722 2236 -762
rect 2236 -6722 2270 -762
rect 2270 -6722 2285 -762
rect 2377 -6722 2394 -762
rect 2394 -6722 2428 -762
rect 2428 -6722 2443 -762
rect 2535 -6722 2552 -762
rect 2552 -6722 2586 -762
rect 2586 -6722 2601 -762
rect 2693 -6722 2710 -762
rect 2710 -6722 2744 -762
rect 2744 -6722 2759 -762
rect 2851 -6722 2868 -762
rect 2868 -6722 2902 -762
rect 2902 -6722 2917 -762
rect 3009 -6722 3026 -762
rect 3026 -6722 3060 -762
rect 3060 -6722 3075 -762
rect 3167 -6722 3184 -762
rect 3184 -6722 3218 -762
rect 3218 -6722 3233 -762
rect 3325 -6722 3342 -762
rect 3342 -6722 3376 -762
rect 3376 -6722 3391 -762
rect 3483 -6722 3500 -762
rect 3500 -6722 3534 -762
rect 3534 -6722 3549 -762
rect 3641 -6722 3658 -762
rect 3658 -6722 3692 -762
rect 3692 -6722 3707 -762
rect 3799 -6722 3816 -762
rect 3816 -6722 3850 -762
rect 3850 -6722 3865 -762
rect 3957 -6722 3974 -762
rect 3974 -6722 4008 -762
rect 4008 -6722 4023 -762
rect 4115 -6722 4132 -762
rect 4132 -6722 4166 -762
rect 4166 -6722 4181 -762
rect 4273 -6722 4290 -762
rect 4290 -6722 4324 -762
rect 4324 -6722 4339 -762
rect 4431 -6722 4448 -762
rect 4448 -6722 4482 -762
rect 4482 -6722 4497 -762
rect 4589 -6722 4606 -762
rect 4606 -6722 4640 -762
rect 4640 -6722 4655 -762
rect 4747 -6722 4764 -762
rect 4764 -6722 4798 -762
rect 4798 -6722 4813 -762
rect 4905 -6722 4922 -762
rect 4922 -6722 4956 -762
rect 4956 -6722 4971 -762
rect 30 -6900 100 -6764
rect 5040 -6764 5054 -720
rect 5054 -6764 5092 -720
rect 5092 -6764 5110 -720
rect 252 -6780 4886 -6774
rect 252 -6814 312 -6780
rect 312 -6814 402 -6780
rect 402 -6814 470 -6780
rect 470 -6814 560 -6780
rect 560 -6814 628 -6780
rect 628 -6814 718 -6780
rect 718 -6814 786 -6780
rect 786 -6814 876 -6780
rect 876 -6814 944 -6780
rect 944 -6814 1034 -6780
rect 1034 -6814 1102 -6780
rect 1102 -6814 1192 -6780
rect 1192 -6814 1260 -6780
rect 1260 -6814 1350 -6780
rect 1350 -6814 1418 -6780
rect 1418 -6814 1508 -6780
rect 1508 -6814 1576 -6780
rect 1576 -6814 1666 -6780
rect 1666 -6814 1734 -6780
rect 1734 -6814 1824 -6780
rect 1824 -6814 1892 -6780
rect 1892 -6814 1982 -6780
rect 1982 -6814 2050 -6780
rect 2050 -6814 2140 -6780
rect 2140 -6814 2208 -6780
rect 2208 -6814 2298 -6780
rect 2298 -6814 2366 -6780
rect 2366 -6814 2456 -6780
rect 2456 -6814 2524 -6780
rect 2524 -6814 2614 -6780
rect 2614 -6814 2682 -6780
rect 2682 -6814 2772 -6780
rect 2772 -6814 2840 -6780
rect 2840 -6814 2930 -6780
rect 2930 -6814 2998 -6780
rect 2998 -6814 3088 -6780
rect 3088 -6814 3156 -6780
rect 3156 -6814 3246 -6780
rect 3246 -6814 3314 -6780
rect 3314 -6814 3404 -6780
rect 3404 -6814 3472 -6780
rect 3472 -6814 3562 -6780
rect 3562 -6814 3630 -6780
rect 3630 -6814 3720 -6780
rect 3720 -6814 3788 -6780
rect 3788 -6814 3878 -6780
rect 3878 -6814 3946 -6780
rect 3946 -6814 4036 -6780
rect 4036 -6814 4104 -6780
rect 4104 -6814 4194 -6780
rect 4194 -6814 4262 -6780
rect 4262 -6814 4352 -6780
rect 4352 -6814 4420 -6780
rect 4420 -6814 4510 -6780
rect 4510 -6814 4578 -6780
rect 4578 -6814 4668 -6780
rect 4668 -6814 4736 -6780
rect 4736 -6814 4826 -6780
rect 4826 -6814 4886 -6780
rect 252 -6874 4886 -6814
rect 5040 -6900 5110 -6764
rect 7030 -720 7100 -580
rect 7252 -670 11886 -610
rect 7252 -704 7312 -670
rect 7312 -704 7402 -670
rect 7402 -704 7470 -670
rect 7470 -704 7560 -670
rect 7560 -704 7628 -670
rect 7628 -704 7718 -670
rect 7718 -704 7786 -670
rect 7786 -704 7876 -670
rect 7876 -704 7944 -670
rect 7944 -704 8034 -670
rect 8034 -704 8102 -670
rect 8102 -704 8192 -670
rect 8192 -704 8260 -670
rect 8260 -704 8350 -670
rect 8350 -704 8418 -670
rect 8418 -704 8508 -670
rect 8508 -704 8576 -670
rect 8576 -704 8666 -670
rect 8666 -704 8734 -670
rect 8734 -704 8824 -670
rect 8824 -704 8892 -670
rect 8892 -704 8982 -670
rect 8982 -704 9050 -670
rect 9050 -704 9140 -670
rect 9140 -704 9208 -670
rect 9208 -704 9298 -670
rect 9298 -704 9366 -670
rect 9366 -704 9456 -670
rect 9456 -704 9524 -670
rect 9524 -704 9614 -670
rect 9614 -704 9682 -670
rect 9682 -704 9772 -670
rect 9772 -704 9840 -670
rect 9840 -704 9930 -670
rect 9930 -704 9998 -670
rect 9998 -704 10088 -670
rect 10088 -704 10156 -670
rect 10156 -704 10246 -670
rect 10246 -704 10314 -670
rect 10314 -704 10404 -670
rect 10404 -704 10472 -670
rect 10472 -704 10562 -670
rect 10562 -704 10630 -670
rect 10630 -704 10720 -670
rect 10720 -704 10788 -670
rect 10788 -704 10878 -670
rect 10878 -704 10946 -670
rect 10946 -704 11036 -670
rect 11036 -704 11104 -670
rect 11104 -704 11194 -670
rect 11194 -704 11262 -670
rect 11262 -704 11352 -670
rect 11352 -704 11420 -670
rect 11420 -704 11510 -670
rect 11510 -704 11578 -670
rect 11578 -704 11668 -670
rect 11668 -704 11736 -670
rect 11736 -704 11826 -670
rect 11826 -704 11886 -670
rect 7252 -710 11886 -704
rect 7030 -6764 7046 -720
rect 7046 -6764 7084 -720
rect 7084 -6764 7100 -720
rect 12040 -720 12110 -580
rect 7165 -6722 7182 -762
rect 7182 -6722 7216 -762
rect 7216 -6722 7231 -762
rect 7323 -6722 7340 -762
rect 7340 -6722 7374 -762
rect 7374 -6722 7389 -762
rect 7481 -6722 7498 -762
rect 7498 -6722 7532 -762
rect 7532 -6722 7547 -762
rect 7639 -6722 7656 -762
rect 7656 -6722 7690 -762
rect 7690 -6722 7705 -762
rect 7797 -6722 7814 -762
rect 7814 -6722 7848 -762
rect 7848 -6722 7863 -762
rect 7955 -6722 7972 -762
rect 7972 -6722 8006 -762
rect 8006 -6722 8021 -762
rect 8113 -6722 8130 -762
rect 8130 -6722 8164 -762
rect 8164 -6722 8179 -762
rect 8271 -6722 8288 -762
rect 8288 -6722 8322 -762
rect 8322 -6722 8337 -762
rect 8429 -6722 8446 -762
rect 8446 -6722 8480 -762
rect 8480 -6722 8495 -762
rect 8587 -6722 8604 -762
rect 8604 -6722 8638 -762
rect 8638 -6722 8653 -762
rect 8745 -6722 8762 -762
rect 8762 -6722 8796 -762
rect 8796 -6722 8811 -762
rect 8903 -6722 8920 -762
rect 8920 -6722 8954 -762
rect 8954 -6722 8969 -762
rect 9061 -6722 9078 -762
rect 9078 -6722 9112 -762
rect 9112 -6722 9127 -762
rect 9219 -6722 9236 -762
rect 9236 -6722 9270 -762
rect 9270 -6722 9285 -762
rect 9377 -6722 9394 -762
rect 9394 -6722 9428 -762
rect 9428 -6722 9443 -762
rect 9535 -6722 9552 -762
rect 9552 -6722 9586 -762
rect 9586 -6722 9601 -762
rect 9693 -6722 9710 -762
rect 9710 -6722 9744 -762
rect 9744 -6722 9759 -762
rect 9851 -6722 9868 -762
rect 9868 -6722 9902 -762
rect 9902 -6722 9917 -762
rect 10009 -6722 10026 -762
rect 10026 -6722 10060 -762
rect 10060 -6722 10075 -762
rect 10167 -6722 10184 -762
rect 10184 -6722 10218 -762
rect 10218 -6722 10233 -762
rect 10325 -6722 10342 -762
rect 10342 -6722 10376 -762
rect 10376 -6722 10391 -762
rect 10483 -6722 10500 -762
rect 10500 -6722 10534 -762
rect 10534 -6722 10549 -762
rect 10641 -6722 10658 -762
rect 10658 -6722 10692 -762
rect 10692 -6722 10707 -762
rect 10799 -6722 10816 -762
rect 10816 -6722 10850 -762
rect 10850 -6722 10865 -762
rect 10957 -6722 10974 -762
rect 10974 -6722 11008 -762
rect 11008 -6722 11023 -762
rect 11115 -6722 11132 -762
rect 11132 -6722 11166 -762
rect 11166 -6722 11181 -762
rect 11273 -6722 11290 -762
rect 11290 -6722 11324 -762
rect 11324 -6722 11339 -762
rect 11431 -6722 11448 -762
rect 11448 -6722 11482 -762
rect 11482 -6722 11497 -762
rect 11589 -6722 11606 -762
rect 11606 -6722 11640 -762
rect 11640 -6722 11655 -762
rect 11747 -6722 11764 -762
rect 11764 -6722 11798 -762
rect 11798 -6722 11813 -762
rect 11905 -6722 11922 -762
rect 11922 -6722 11956 -762
rect 11956 -6722 11971 -762
rect 7030 -6900 7100 -6764
rect 12040 -6764 12054 -720
rect 12054 -6764 12092 -720
rect 12092 -6764 12110 -720
rect 7252 -6780 11886 -6774
rect 7252 -6814 7312 -6780
rect 7312 -6814 7402 -6780
rect 7402 -6814 7470 -6780
rect 7470 -6814 7560 -6780
rect 7560 -6814 7628 -6780
rect 7628 -6814 7718 -6780
rect 7718 -6814 7786 -6780
rect 7786 -6814 7876 -6780
rect 7876 -6814 7944 -6780
rect 7944 -6814 8034 -6780
rect 8034 -6814 8102 -6780
rect 8102 -6814 8192 -6780
rect 8192 -6814 8260 -6780
rect 8260 -6814 8350 -6780
rect 8350 -6814 8418 -6780
rect 8418 -6814 8508 -6780
rect 8508 -6814 8576 -6780
rect 8576 -6814 8666 -6780
rect 8666 -6814 8734 -6780
rect 8734 -6814 8824 -6780
rect 8824 -6814 8892 -6780
rect 8892 -6814 8982 -6780
rect 8982 -6814 9050 -6780
rect 9050 -6814 9140 -6780
rect 9140 -6814 9208 -6780
rect 9208 -6814 9298 -6780
rect 9298 -6814 9366 -6780
rect 9366 -6814 9456 -6780
rect 9456 -6814 9524 -6780
rect 9524 -6814 9614 -6780
rect 9614 -6814 9682 -6780
rect 9682 -6814 9772 -6780
rect 9772 -6814 9840 -6780
rect 9840 -6814 9930 -6780
rect 9930 -6814 9998 -6780
rect 9998 -6814 10088 -6780
rect 10088 -6814 10156 -6780
rect 10156 -6814 10246 -6780
rect 10246 -6814 10314 -6780
rect 10314 -6814 10404 -6780
rect 10404 -6814 10472 -6780
rect 10472 -6814 10562 -6780
rect 10562 -6814 10630 -6780
rect 10630 -6814 10720 -6780
rect 10720 -6814 10788 -6780
rect 10788 -6814 10878 -6780
rect 10878 -6814 10946 -6780
rect 10946 -6814 11036 -6780
rect 11036 -6814 11104 -6780
rect 11104 -6814 11194 -6780
rect 11194 -6814 11262 -6780
rect 11262 -6814 11352 -6780
rect 11352 -6814 11420 -6780
rect 11420 -6814 11510 -6780
rect 11510 -6814 11578 -6780
rect 11578 -6814 11668 -6780
rect 11668 -6814 11736 -6780
rect 11736 -6814 11826 -6780
rect 11826 -6814 11886 -6780
rect 7252 -6874 11886 -6814
rect 12040 -6900 12110 -6764
rect 14030 -720 14100 -580
rect 14252 -670 18886 -610
rect 14252 -704 14312 -670
rect 14312 -704 14402 -670
rect 14402 -704 14470 -670
rect 14470 -704 14560 -670
rect 14560 -704 14628 -670
rect 14628 -704 14718 -670
rect 14718 -704 14786 -670
rect 14786 -704 14876 -670
rect 14876 -704 14944 -670
rect 14944 -704 15034 -670
rect 15034 -704 15102 -670
rect 15102 -704 15192 -670
rect 15192 -704 15260 -670
rect 15260 -704 15350 -670
rect 15350 -704 15418 -670
rect 15418 -704 15508 -670
rect 15508 -704 15576 -670
rect 15576 -704 15666 -670
rect 15666 -704 15734 -670
rect 15734 -704 15824 -670
rect 15824 -704 15892 -670
rect 15892 -704 15982 -670
rect 15982 -704 16050 -670
rect 16050 -704 16140 -670
rect 16140 -704 16208 -670
rect 16208 -704 16298 -670
rect 16298 -704 16366 -670
rect 16366 -704 16456 -670
rect 16456 -704 16524 -670
rect 16524 -704 16614 -670
rect 16614 -704 16682 -670
rect 16682 -704 16772 -670
rect 16772 -704 16840 -670
rect 16840 -704 16930 -670
rect 16930 -704 16998 -670
rect 16998 -704 17088 -670
rect 17088 -704 17156 -670
rect 17156 -704 17246 -670
rect 17246 -704 17314 -670
rect 17314 -704 17404 -670
rect 17404 -704 17472 -670
rect 17472 -704 17562 -670
rect 17562 -704 17630 -670
rect 17630 -704 17720 -670
rect 17720 -704 17788 -670
rect 17788 -704 17878 -670
rect 17878 -704 17946 -670
rect 17946 -704 18036 -670
rect 18036 -704 18104 -670
rect 18104 -704 18194 -670
rect 18194 -704 18262 -670
rect 18262 -704 18352 -670
rect 18352 -704 18420 -670
rect 18420 -704 18510 -670
rect 18510 -704 18578 -670
rect 18578 -704 18668 -670
rect 18668 -704 18736 -670
rect 18736 -704 18826 -670
rect 18826 -704 18886 -670
rect 14252 -710 18886 -704
rect 14030 -6764 14046 -720
rect 14046 -6764 14084 -720
rect 14084 -6764 14100 -720
rect 19040 -720 19110 -580
rect 14165 -6722 14182 -762
rect 14182 -6722 14216 -762
rect 14216 -6722 14231 -762
rect 14323 -6722 14340 -762
rect 14340 -6722 14374 -762
rect 14374 -6722 14389 -762
rect 14481 -6722 14498 -762
rect 14498 -6722 14532 -762
rect 14532 -6722 14547 -762
rect 14639 -6722 14656 -762
rect 14656 -6722 14690 -762
rect 14690 -6722 14705 -762
rect 14797 -6722 14814 -762
rect 14814 -6722 14848 -762
rect 14848 -6722 14863 -762
rect 14955 -6722 14972 -762
rect 14972 -6722 15006 -762
rect 15006 -6722 15021 -762
rect 15113 -6722 15130 -762
rect 15130 -6722 15164 -762
rect 15164 -6722 15179 -762
rect 15271 -6722 15288 -762
rect 15288 -6722 15322 -762
rect 15322 -6722 15337 -762
rect 15429 -6722 15446 -762
rect 15446 -6722 15480 -762
rect 15480 -6722 15495 -762
rect 15587 -6722 15604 -762
rect 15604 -6722 15638 -762
rect 15638 -6722 15653 -762
rect 15745 -6722 15762 -762
rect 15762 -6722 15796 -762
rect 15796 -6722 15811 -762
rect 15903 -6722 15920 -762
rect 15920 -6722 15954 -762
rect 15954 -6722 15969 -762
rect 16061 -6722 16078 -762
rect 16078 -6722 16112 -762
rect 16112 -6722 16127 -762
rect 16219 -6722 16236 -762
rect 16236 -6722 16270 -762
rect 16270 -6722 16285 -762
rect 16377 -6722 16394 -762
rect 16394 -6722 16428 -762
rect 16428 -6722 16443 -762
rect 16535 -6722 16552 -762
rect 16552 -6722 16586 -762
rect 16586 -6722 16601 -762
rect 16693 -6722 16710 -762
rect 16710 -6722 16744 -762
rect 16744 -6722 16759 -762
rect 16851 -6722 16868 -762
rect 16868 -6722 16902 -762
rect 16902 -6722 16917 -762
rect 17009 -6722 17026 -762
rect 17026 -6722 17060 -762
rect 17060 -6722 17075 -762
rect 17167 -6722 17184 -762
rect 17184 -6722 17218 -762
rect 17218 -6722 17233 -762
rect 17325 -6722 17342 -762
rect 17342 -6722 17376 -762
rect 17376 -6722 17391 -762
rect 17483 -6722 17500 -762
rect 17500 -6722 17534 -762
rect 17534 -6722 17549 -762
rect 17641 -6722 17658 -762
rect 17658 -6722 17692 -762
rect 17692 -6722 17707 -762
rect 17799 -6722 17816 -762
rect 17816 -6722 17850 -762
rect 17850 -6722 17865 -762
rect 17957 -6722 17974 -762
rect 17974 -6722 18008 -762
rect 18008 -6722 18023 -762
rect 18115 -6722 18132 -762
rect 18132 -6722 18166 -762
rect 18166 -6722 18181 -762
rect 18273 -6722 18290 -762
rect 18290 -6722 18324 -762
rect 18324 -6722 18339 -762
rect 18431 -6722 18448 -762
rect 18448 -6722 18482 -762
rect 18482 -6722 18497 -762
rect 18589 -6722 18606 -762
rect 18606 -6722 18640 -762
rect 18640 -6722 18655 -762
rect 18747 -6722 18764 -762
rect 18764 -6722 18798 -762
rect 18798 -6722 18813 -762
rect 18905 -6722 18922 -762
rect 18922 -6722 18956 -762
rect 18956 -6722 18971 -762
rect 14030 -6900 14100 -6764
rect 19040 -6764 19054 -720
rect 19054 -6764 19092 -720
rect 19092 -6764 19110 -720
rect 14252 -6780 18886 -6774
rect 14252 -6814 14312 -6780
rect 14312 -6814 14402 -6780
rect 14402 -6814 14470 -6780
rect 14470 -6814 14560 -6780
rect 14560 -6814 14628 -6780
rect 14628 -6814 14718 -6780
rect 14718 -6814 14786 -6780
rect 14786 -6814 14876 -6780
rect 14876 -6814 14944 -6780
rect 14944 -6814 15034 -6780
rect 15034 -6814 15102 -6780
rect 15102 -6814 15192 -6780
rect 15192 -6814 15260 -6780
rect 15260 -6814 15350 -6780
rect 15350 -6814 15418 -6780
rect 15418 -6814 15508 -6780
rect 15508 -6814 15576 -6780
rect 15576 -6814 15666 -6780
rect 15666 -6814 15734 -6780
rect 15734 -6814 15824 -6780
rect 15824 -6814 15892 -6780
rect 15892 -6814 15982 -6780
rect 15982 -6814 16050 -6780
rect 16050 -6814 16140 -6780
rect 16140 -6814 16208 -6780
rect 16208 -6814 16298 -6780
rect 16298 -6814 16366 -6780
rect 16366 -6814 16456 -6780
rect 16456 -6814 16524 -6780
rect 16524 -6814 16614 -6780
rect 16614 -6814 16682 -6780
rect 16682 -6814 16772 -6780
rect 16772 -6814 16840 -6780
rect 16840 -6814 16930 -6780
rect 16930 -6814 16998 -6780
rect 16998 -6814 17088 -6780
rect 17088 -6814 17156 -6780
rect 17156 -6814 17246 -6780
rect 17246 -6814 17314 -6780
rect 17314 -6814 17404 -6780
rect 17404 -6814 17472 -6780
rect 17472 -6814 17562 -6780
rect 17562 -6814 17630 -6780
rect 17630 -6814 17720 -6780
rect 17720 -6814 17788 -6780
rect 17788 -6814 17878 -6780
rect 17878 -6814 17946 -6780
rect 17946 -6814 18036 -6780
rect 18036 -6814 18104 -6780
rect 18104 -6814 18194 -6780
rect 18194 -6814 18262 -6780
rect 18262 -6814 18352 -6780
rect 18352 -6814 18420 -6780
rect 18420 -6814 18510 -6780
rect 18510 -6814 18578 -6780
rect 18578 -6814 18668 -6780
rect 18668 -6814 18736 -6780
rect 18736 -6814 18826 -6780
rect 18826 -6814 18886 -6780
rect 14252 -6874 18886 -6814
rect 19040 -6900 19110 -6764
rect 21030 -720 21100 -580
rect 21252 -670 25886 -610
rect 21252 -704 21312 -670
rect 21312 -704 21402 -670
rect 21402 -704 21470 -670
rect 21470 -704 21560 -670
rect 21560 -704 21628 -670
rect 21628 -704 21718 -670
rect 21718 -704 21786 -670
rect 21786 -704 21876 -670
rect 21876 -704 21944 -670
rect 21944 -704 22034 -670
rect 22034 -704 22102 -670
rect 22102 -704 22192 -670
rect 22192 -704 22260 -670
rect 22260 -704 22350 -670
rect 22350 -704 22418 -670
rect 22418 -704 22508 -670
rect 22508 -704 22576 -670
rect 22576 -704 22666 -670
rect 22666 -704 22734 -670
rect 22734 -704 22824 -670
rect 22824 -704 22892 -670
rect 22892 -704 22982 -670
rect 22982 -704 23050 -670
rect 23050 -704 23140 -670
rect 23140 -704 23208 -670
rect 23208 -704 23298 -670
rect 23298 -704 23366 -670
rect 23366 -704 23456 -670
rect 23456 -704 23524 -670
rect 23524 -704 23614 -670
rect 23614 -704 23682 -670
rect 23682 -704 23772 -670
rect 23772 -704 23840 -670
rect 23840 -704 23930 -670
rect 23930 -704 23998 -670
rect 23998 -704 24088 -670
rect 24088 -704 24156 -670
rect 24156 -704 24246 -670
rect 24246 -704 24314 -670
rect 24314 -704 24404 -670
rect 24404 -704 24472 -670
rect 24472 -704 24562 -670
rect 24562 -704 24630 -670
rect 24630 -704 24720 -670
rect 24720 -704 24788 -670
rect 24788 -704 24878 -670
rect 24878 -704 24946 -670
rect 24946 -704 25036 -670
rect 25036 -704 25104 -670
rect 25104 -704 25194 -670
rect 25194 -704 25262 -670
rect 25262 -704 25352 -670
rect 25352 -704 25420 -670
rect 25420 -704 25510 -670
rect 25510 -704 25578 -670
rect 25578 -704 25668 -670
rect 25668 -704 25736 -670
rect 25736 -704 25826 -670
rect 25826 -704 25886 -670
rect 21252 -710 25886 -704
rect 21030 -6764 21046 -720
rect 21046 -6764 21084 -720
rect 21084 -6764 21100 -720
rect 26040 -720 26110 -580
rect 21165 -6722 21182 -762
rect 21182 -6722 21216 -762
rect 21216 -6722 21231 -762
rect 21323 -6722 21340 -762
rect 21340 -6722 21374 -762
rect 21374 -6722 21389 -762
rect 21481 -6722 21498 -762
rect 21498 -6722 21532 -762
rect 21532 -6722 21547 -762
rect 21639 -6722 21656 -762
rect 21656 -6722 21690 -762
rect 21690 -6722 21705 -762
rect 21797 -6722 21814 -762
rect 21814 -6722 21848 -762
rect 21848 -6722 21863 -762
rect 21955 -6722 21972 -762
rect 21972 -6722 22006 -762
rect 22006 -6722 22021 -762
rect 22113 -6722 22130 -762
rect 22130 -6722 22164 -762
rect 22164 -6722 22179 -762
rect 22271 -6722 22288 -762
rect 22288 -6722 22322 -762
rect 22322 -6722 22337 -762
rect 22429 -6722 22446 -762
rect 22446 -6722 22480 -762
rect 22480 -6722 22495 -762
rect 22587 -6722 22604 -762
rect 22604 -6722 22638 -762
rect 22638 -6722 22653 -762
rect 22745 -6722 22762 -762
rect 22762 -6722 22796 -762
rect 22796 -6722 22811 -762
rect 22903 -6722 22920 -762
rect 22920 -6722 22954 -762
rect 22954 -6722 22969 -762
rect 23061 -6722 23078 -762
rect 23078 -6722 23112 -762
rect 23112 -6722 23127 -762
rect 23219 -6722 23236 -762
rect 23236 -6722 23270 -762
rect 23270 -6722 23285 -762
rect 23377 -6722 23394 -762
rect 23394 -6722 23428 -762
rect 23428 -6722 23443 -762
rect 23535 -6722 23552 -762
rect 23552 -6722 23586 -762
rect 23586 -6722 23601 -762
rect 23693 -6722 23710 -762
rect 23710 -6722 23744 -762
rect 23744 -6722 23759 -762
rect 23851 -6722 23868 -762
rect 23868 -6722 23902 -762
rect 23902 -6722 23917 -762
rect 24009 -6722 24026 -762
rect 24026 -6722 24060 -762
rect 24060 -6722 24075 -762
rect 24167 -6722 24184 -762
rect 24184 -6722 24218 -762
rect 24218 -6722 24233 -762
rect 24325 -6722 24342 -762
rect 24342 -6722 24376 -762
rect 24376 -6722 24391 -762
rect 24483 -6722 24500 -762
rect 24500 -6722 24534 -762
rect 24534 -6722 24549 -762
rect 24641 -6722 24658 -762
rect 24658 -6722 24692 -762
rect 24692 -6722 24707 -762
rect 24799 -6722 24816 -762
rect 24816 -6722 24850 -762
rect 24850 -6722 24865 -762
rect 24957 -6722 24974 -762
rect 24974 -6722 25008 -762
rect 25008 -6722 25023 -762
rect 25115 -6722 25132 -762
rect 25132 -6722 25166 -762
rect 25166 -6722 25181 -762
rect 25273 -6722 25290 -762
rect 25290 -6722 25324 -762
rect 25324 -6722 25339 -762
rect 25431 -6722 25448 -762
rect 25448 -6722 25482 -762
rect 25482 -6722 25497 -762
rect 25589 -6722 25606 -762
rect 25606 -6722 25640 -762
rect 25640 -6722 25655 -762
rect 25747 -6722 25764 -762
rect 25764 -6722 25798 -762
rect 25798 -6722 25813 -762
rect 25905 -6722 25922 -762
rect 25922 -6722 25956 -762
rect 25956 -6722 25971 -762
rect 21030 -6900 21100 -6764
rect 26040 -6764 26054 -720
rect 26054 -6764 26092 -720
rect 26092 -6764 26110 -720
rect 21252 -6780 25886 -6774
rect 21252 -6814 21312 -6780
rect 21312 -6814 21402 -6780
rect 21402 -6814 21470 -6780
rect 21470 -6814 21560 -6780
rect 21560 -6814 21628 -6780
rect 21628 -6814 21718 -6780
rect 21718 -6814 21786 -6780
rect 21786 -6814 21876 -6780
rect 21876 -6814 21944 -6780
rect 21944 -6814 22034 -6780
rect 22034 -6814 22102 -6780
rect 22102 -6814 22192 -6780
rect 22192 -6814 22260 -6780
rect 22260 -6814 22350 -6780
rect 22350 -6814 22418 -6780
rect 22418 -6814 22508 -6780
rect 22508 -6814 22576 -6780
rect 22576 -6814 22666 -6780
rect 22666 -6814 22734 -6780
rect 22734 -6814 22824 -6780
rect 22824 -6814 22892 -6780
rect 22892 -6814 22982 -6780
rect 22982 -6814 23050 -6780
rect 23050 -6814 23140 -6780
rect 23140 -6814 23208 -6780
rect 23208 -6814 23298 -6780
rect 23298 -6814 23366 -6780
rect 23366 -6814 23456 -6780
rect 23456 -6814 23524 -6780
rect 23524 -6814 23614 -6780
rect 23614 -6814 23682 -6780
rect 23682 -6814 23772 -6780
rect 23772 -6814 23840 -6780
rect 23840 -6814 23930 -6780
rect 23930 -6814 23998 -6780
rect 23998 -6814 24088 -6780
rect 24088 -6814 24156 -6780
rect 24156 -6814 24246 -6780
rect 24246 -6814 24314 -6780
rect 24314 -6814 24404 -6780
rect 24404 -6814 24472 -6780
rect 24472 -6814 24562 -6780
rect 24562 -6814 24630 -6780
rect 24630 -6814 24720 -6780
rect 24720 -6814 24788 -6780
rect 24788 -6814 24878 -6780
rect 24878 -6814 24946 -6780
rect 24946 -6814 25036 -6780
rect 25036 -6814 25104 -6780
rect 25104 -6814 25194 -6780
rect 25194 -6814 25262 -6780
rect 25262 -6814 25352 -6780
rect 25352 -6814 25420 -6780
rect 25420 -6814 25510 -6780
rect 25510 -6814 25578 -6780
rect 25578 -6814 25668 -6780
rect 25668 -6814 25736 -6780
rect 25736 -6814 25826 -6780
rect 25826 -6814 25886 -6780
rect 21252 -6874 25886 -6814
rect 26040 -6900 26110 -6764
<< metal2 >>
rect 12600 11700 13600 11900
rect 12600 6500 13000 11700
rect 13200 6500 13600 11700
rect 5100 6480 7100 6500
rect 12100 6480 14100 6500
rect 19100 6480 21100 6500
rect 30 6420 100 6480
rect 5040 6420 7100 6480
rect 232 6380 252 6390
rect 4886 6380 4906 6390
rect 232 6310 240 6380
rect 4900 6310 4906 6380
rect 232 6290 252 6310
rect 4886 6290 4906 6310
rect 165 6238 231 6258
rect 165 258 231 278
rect 323 6238 389 6258
rect 323 258 389 278
rect 481 6238 547 6258
rect 481 258 547 278
rect 639 6238 705 6258
rect 639 258 705 278
rect 797 6238 863 6258
rect 797 258 863 278
rect 955 6238 1021 6258
rect 955 258 1021 278
rect 1113 6238 1179 6258
rect 1113 258 1179 278
rect 1271 6238 1337 6258
rect 1271 258 1337 278
rect 1429 6238 1495 6258
rect 1429 258 1495 278
rect 1587 6238 1653 6258
rect 1587 258 1653 278
rect 1745 6238 1811 6258
rect 1745 258 1811 278
rect 1903 6238 1969 6258
rect 1903 258 1969 278
rect 2061 6238 2127 6258
rect 2061 258 2127 278
rect 2219 6238 2285 6258
rect 2219 258 2285 278
rect 2377 6238 2443 6258
rect 2377 258 2443 278
rect 2535 6238 2601 6258
rect 2535 258 2601 278
rect 2693 6238 2759 6258
rect 2693 258 2759 278
rect 2851 6238 2917 6258
rect 2851 258 2917 278
rect 3009 6238 3075 6258
rect 3009 258 3075 278
rect 3167 6238 3233 6258
rect 3167 258 3233 278
rect 3325 6238 3391 6258
rect 3325 258 3391 278
rect 3483 6238 3549 6258
rect 3483 258 3549 278
rect 3641 6238 3707 6258
rect 3641 258 3707 278
rect 3799 6238 3865 6258
rect 3799 258 3865 278
rect 3957 6238 4023 6258
rect 3957 258 4023 278
rect 4115 6238 4181 6258
rect 4115 258 4181 278
rect 4273 6238 4339 6258
rect 4273 258 4339 278
rect 4431 6238 4497 6258
rect 4431 258 4497 278
rect 4589 6238 4655 6258
rect 4589 258 4655 278
rect 4747 6238 4813 6258
rect 4747 258 4813 278
rect 4905 6238 4971 6258
rect 4905 258 4971 278
rect 232 210 252 226
rect 4886 210 4906 226
rect 232 140 240 210
rect 4890 140 4906 210
rect 232 126 252 140
rect 4886 126 4906 140
rect 30 30 100 100
rect 5110 6300 7030 6420
rect 5300 5800 5700 6300
rect 5900 5800 6300 6300
rect 6500 5800 6900 6300
rect 5110 5600 7030 5800
rect 5110 100 7030 200
rect 12040 6420 14100 6480
rect 7232 6380 7252 6390
rect 11886 6380 11906 6390
rect 7232 6310 7240 6380
rect 11900 6310 11906 6380
rect 7232 6290 7252 6310
rect 11886 6290 11906 6310
rect 7165 6238 7231 6258
rect 7165 258 7231 278
rect 7323 6238 7389 6258
rect 7323 258 7389 278
rect 7481 6238 7547 6258
rect 7481 258 7547 278
rect 7639 6238 7705 6258
rect 7639 258 7705 278
rect 7797 6238 7863 6258
rect 7797 258 7863 278
rect 7955 6238 8021 6258
rect 7955 258 8021 278
rect 8113 6238 8179 6258
rect 8113 258 8179 278
rect 8271 6238 8337 6258
rect 8271 258 8337 278
rect 8429 6238 8495 6258
rect 8429 258 8495 278
rect 8587 6238 8653 6258
rect 8587 258 8653 278
rect 8745 6238 8811 6258
rect 8745 258 8811 278
rect 8903 6238 8969 6258
rect 8903 258 8969 278
rect 9061 6238 9127 6258
rect 9061 258 9127 278
rect 9219 6238 9285 6258
rect 9219 258 9285 278
rect 9377 6238 9443 6258
rect 9377 258 9443 278
rect 9535 6238 9601 6258
rect 9535 258 9601 278
rect 9693 6238 9759 6258
rect 9693 258 9759 278
rect 9851 6238 9917 6258
rect 9851 258 9917 278
rect 10009 6238 10075 6258
rect 10009 258 10075 278
rect 10167 6238 10233 6258
rect 10167 258 10233 278
rect 10325 6238 10391 6258
rect 10325 258 10391 278
rect 10483 6238 10549 6258
rect 10483 258 10549 278
rect 10641 6238 10707 6258
rect 10641 258 10707 278
rect 10799 6238 10865 6258
rect 10799 258 10865 278
rect 10957 6238 11023 6258
rect 10957 258 11023 278
rect 11115 6238 11181 6258
rect 11115 258 11181 278
rect 11273 6238 11339 6258
rect 11273 258 11339 278
rect 11431 6238 11497 6258
rect 11431 258 11497 278
rect 11589 6238 11655 6258
rect 11589 258 11655 278
rect 11747 6238 11813 6258
rect 11747 258 11813 278
rect 11905 6238 11971 6258
rect 11905 258 11971 278
rect 7232 210 7252 226
rect 11886 210 11906 226
rect 7232 140 7240 210
rect 11890 140 11906 210
rect 7232 126 7252 140
rect 11886 126 11906 140
rect 5040 30 7100 100
rect 12110 6300 14030 6420
rect 12300 5800 12700 6300
rect 12900 5800 13300 6300
rect 13500 5800 13900 6300
rect 12110 5600 14030 5800
rect 12600 200 13000 5600
rect 13200 200 13600 5600
rect 12110 100 14030 200
rect 19040 6420 21100 6480
rect 14232 6380 14252 6390
rect 18886 6380 18906 6390
rect 14232 6310 14240 6380
rect 18900 6310 18906 6380
rect 14232 6290 14252 6310
rect 18886 6290 18906 6310
rect 14165 6238 14231 6258
rect 14165 258 14231 278
rect 14323 6238 14389 6258
rect 14323 258 14389 278
rect 14481 6238 14547 6258
rect 14481 258 14547 278
rect 14639 6238 14705 6258
rect 14639 258 14705 278
rect 14797 6238 14863 6258
rect 14797 258 14863 278
rect 14955 6238 15021 6258
rect 14955 258 15021 278
rect 15113 6238 15179 6258
rect 15113 258 15179 278
rect 15271 6238 15337 6258
rect 15271 258 15337 278
rect 15429 6238 15495 6258
rect 15429 258 15495 278
rect 15587 6238 15653 6258
rect 15587 258 15653 278
rect 15745 6238 15811 6258
rect 15745 258 15811 278
rect 15903 6238 15969 6258
rect 15903 258 15969 278
rect 16061 6238 16127 6258
rect 16061 258 16127 278
rect 16219 6238 16285 6258
rect 16219 258 16285 278
rect 16377 6238 16443 6258
rect 16377 258 16443 278
rect 16535 6238 16601 6258
rect 16535 258 16601 278
rect 16693 6238 16759 6258
rect 16693 258 16759 278
rect 16851 6238 16917 6258
rect 16851 258 16917 278
rect 17009 6238 17075 6258
rect 17009 258 17075 278
rect 17167 6238 17233 6258
rect 17167 258 17233 278
rect 17325 6238 17391 6258
rect 17325 258 17391 278
rect 17483 6238 17549 6258
rect 17483 258 17549 278
rect 17641 6238 17707 6258
rect 17641 258 17707 278
rect 17799 6238 17865 6258
rect 17799 258 17865 278
rect 17957 6238 18023 6258
rect 17957 258 18023 278
rect 18115 6238 18181 6258
rect 18115 258 18181 278
rect 18273 6238 18339 6258
rect 18273 258 18339 278
rect 18431 6238 18497 6258
rect 18431 258 18497 278
rect 18589 6238 18655 6258
rect 18589 258 18655 278
rect 18747 6238 18813 6258
rect 18747 258 18813 278
rect 18905 6238 18971 6258
rect 18905 258 18971 278
rect 14232 210 14252 226
rect 18886 210 18906 226
rect 14232 140 14240 210
rect 18890 140 18906 210
rect 14232 126 14252 140
rect 18886 126 18906 140
rect 12040 30 14100 100
rect 19110 6300 21030 6420
rect 19300 5800 19700 6300
rect 19900 5800 20300 6300
rect 20500 5800 20900 6300
rect 19110 5600 21030 5800
rect 19110 100 21030 200
rect 26040 6420 26110 6480
rect 21232 6380 21252 6390
rect 25886 6380 25906 6390
rect 21232 6310 21240 6380
rect 25900 6310 25906 6380
rect 21232 6290 21252 6310
rect 25886 6290 25906 6310
rect 21165 6238 21231 6258
rect 21165 258 21231 278
rect 21323 6238 21389 6258
rect 21323 258 21389 278
rect 21481 6238 21547 6258
rect 21481 258 21547 278
rect 21639 6238 21705 6258
rect 21639 258 21705 278
rect 21797 6238 21863 6258
rect 21797 258 21863 278
rect 21955 6238 22021 6258
rect 21955 258 22021 278
rect 22113 6238 22179 6258
rect 22113 258 22179 278
rect 22271 6238 22337 6258
rect 22271 258 22337 278
rect 22429 6238 22495 6258
rect 22429 258 22495 278
rect 22587 6238 22653 6258
rect 22587 258 22653 278
rect 22745 6238 22811 6258
rect 22745 258 22811 278
rect 22903 6238 22969 6258
rect 22903 258 22969 278
rect 23061 6238 23127 6258
rect 23061 258 23127 278
rect 23219 6238 23285 6258
rect 23219 258 23285 278
rect 23377 6238 23443 6258
rect 23377 258 23443 278
rect 23535 6238 23601 6258
rect 23535 258 23601 278
rect 23693 6238 23759 6258
rect 23693 258 23759 278
rect 23851 6238 23917 6258
rect 23851 258 23917 278
rect 24009 6238 24075 6258
rect 24009 258 24075 278
rect 24167 6238 24233 6258
rect 24167 258 24233 278
rect 24325 6238 24391 6258
rect 24325 258 24391 278
rect 24483 6238 24549 6258
rect 24483 258 24549 278
rect 24641 6238 24707 6258
rect 24641 258 24707 278
rect 24799 6238 24865 6258
rect 24799 258 24865 278
rect 24957 6238 25023 6258
rect 24957 258 25023 278
rect 25115 6238 25181 6258
rect 25115 258 25181 278
rect 25273 6238 25339 6258
rect 25273 258 25339 278
rect 25431 6238 25497 6258
rect 25431 258 25497 278
rect 25589 6238 25655 6258
rect 25589 258 25655 278
rect 25747 6238 25813 6258
rect 25747 258 25813 278
rect 25905 6238 25971 6258
rect 25905 258 25971 278
rect 21232 210 21252 226
rect 25886 210 25906 226
rect 21232 140 21240 210
rect 25890 140 25906 210
rect 21232 126 21252 140
rect 25886 126 25906 140
rect 19040 30 21100 100
rect 26040 30 26110 100
rect 5100 0 7100 30
rect 12100 0 14100 30
rect 19100 0 21100 30
rect 5300 -500 5700 0
rect 5900 -500 6300 0
rect 6500 -500 6900 0
rect 12300 -500 12700 0
rect 12900 -500 13300 0
rect 13500 -500 13900 0
rect 19300 -500 19700 0
rect 19900 -500 20300 0
rect 20500 -500 20900 0
rect 5100 -520 7100 -500
rect 12100 -520 14100 -500
rect 19100 -520 21100 -500
rect 30 -580 100 -520
rect 5040 -580 7100 -520
rect 232 -620 252 -610
rect 4886 -620 4906 -610
rect 232 -690 240 -620
rect 4900 -690 4906 -620
rect 232 -710 252 -690
rect 4886 -710 4906 -690
rect 165 -762 231 -742
rect 165 -6742 231 -6722
rect 323 -762 389 -742
rect 323 -6742 389 -6722
rect 481 -762 547 -742
rect 481 -6742 547 -6722
rect 639 -762 705 -742
rect 639 -6742 705 -6722
rect 797 -762 863 -742
rect 797 -6742 863 -6722
rect 955 -762 1021 -742
rect 955 -6742 1021 -6722
rect 1113 -762 1179 -742
rect 1113 -6742 1179 -6722
rect 1271 -762 1337 -742
rect 1271 -6742 1337 -6722
rect 1429 -762 1495 -742
rect 1429 -6742 1495 -6722
rect 1587 -762 1653 -742
rect 1587 -6742 1653 -6722
rect 1745 -762 1811 -742
rect 1745 -6742 1811 -6722
rect 1903 -762 1969 -742
rect 1903 -6742 1969 -6722
rect 2061 -762 2127 -742
rect 2061 -6742 2127 -6722
rect 2219 -762 2285 -742
rect 2219 -6742 2285 -6722
rect 2377 -762 2443 -742
rect 2377 -6742 2443 -6722
rect 2535 -762 2601 -742
rect 2535 -6742 2601 -6722
rect 2693 -762 2759 -742
rect 2693 -6742 2759 -6722
rect 2851 -762 2917 -742
rect 2851 -6742 2917 -6722
rect 3009 -762 3075 -742
rect 3009 -6742 3075 -6722
rect 3167 -762 3233 -742
rect 3167 -6742 3233 -6722
rect 3325 -762 3391 -742
rect 3325 -6742 3391 -6722
rect 3483 -762 3549 -742
rect 3483 -6742 3549 -6722
rect 3641 -762 3707 -742
rect 3641 -6742 3707 -6722
rect 3799 -762 3865 -742
rect 3799 -6742 3865 -6722
rect 3957 -762 4023 -742
rect 3957 -6742 4023 -6722
rect 4115 -762 4181 -742
rect 4115 -6742 4181 -6722
rect 4273 -762 4339 -742
rect 4273 -6742 4339 -6722
rect 4431 -762 4497 -742
rect 4431 -6742 4497 -6722
rect 4589 -762 4655 -742
rect 4589 -6742 4655 -6722
rect 4747 -762 4813 -742
rect 4747 -6742 4813 -6722
rect 4905 -762 4971 -742
rect 4905 -6742 4971 -6722
rect 232 -6790 252 -6774
rect 4886 -6790 4906 -6774
rect 232 -6860 240 -6790
rect 4890 -6860 4906 -6790
rect 232 -6874 252 -6860
rect 4886 -6874 4906 -6860
rect 30 -6970 100 -6900
rect 5110 -700 7030 -580
rect 5110 -6200 7030 -6000
rect 5300 -6700 5700 -6200
rect 5900 -6700 6300 -6200
rect 6500 -6700 6900 -6200
rect 5110 -6900 7030 -6700
rect 12040 -580 14100 -520
rect 7232 -620 7252 -610
rect 11886 -620 11906 -610
rect 7232 -690 7240 -620
rect 11900 -690 11906 -620
rect 7232 -710 7252 -690
rect 11886 -710 11906 -690
rect 7165 -762 7231 -742
rect 7165 -6742 7231 -6722
rect 7323 -762 7389 -742
rect 7323 -6742 7389 -6722
rect 7481 -762 7547 -742
rect 7481 -6742 7547 -6722
rect 7639 -762 7705 -742
rect 7639 -6742 7705 -6722
rect 7797 -762 7863 -742
rect 7797 -6742 7863 -6722
rect 7955 -762 8021 -742
rect 7955 -6742 8021 -6722
rect 8113 -762 8179 -742
rect 8113 -6742 8179 -6722
rect 8271 -762 8337 -742
rect 8271 -6742 8337 -6722
rect 8429 -762 8495 -742
rect 8429 -6742 8495 -6722
rect 8587 -762 8653 -742
rect 8587 -6742 8653 -6722
rect 8745 -762 8811 -742
rect 8745 -6742 8811 -6722
rect 8903 -762 8969 -742
rect 8903 -6742 8969 -6722
rect 9061 -762 9127 -742
rect 9061 -6742 9127 -6722
rect 9219 -762 9285 -742
rect 9219 -6742 9285 -6722
rect 9377 -762 9443 -742
rect 9377 -6742 9443 -6722
rect 9535 -762 9601 -742
rect 9535 -6742 9601 -6722
rect 9693 -762 9759 -742
rect 9693 -6742 9759 -6722
rect 9851 -762 9917 -742
rect 9851 -6742 9917 -6722
rect 10009 -762 10075 -742
rect 10009 -6742 10075 -6722
rect 10167 -762 10233 -742
rect 10167 -6742 10233 -6722
rect 10325 -762 10391 -742
rect 10325 -6742 10391 -6722
rect 10483 -762 10549 -742
rect 10483 -6742 10549 -6722
rect 10641 -762 10707 -742
rect 10641 -6742 10707 -6722
rect 10799 -762 10865 -742
rect 10799 -6742 10865 -6722
rect 10957 -762 11023 -742
rect 10957 -6742 11023 -6722
rect 11115 -762 11181 -742
rect 11115 -6742 11181 -6722
rect 11273 -762 11339 -742
rect 11273 -6742 11339 -6722
rect 11431 -762 11497 -742
rect 11431 -6742 11497 -6722
rect 11589 -762 11655 -742
rect 11589 -6742 11655 -6722
rect 11747 -762 11813 -742
rect 11747 -6742 11813 -6722
rect 11905 -762 11971 -742
rect 11905 -6742 11971 -6722
rect 7232 -6790 7252 -6774
rect 11886 -6790 11906 -6774
rect 7232 -6860 7240 -6790
rect 11890 -6860 11906 -6790
rect 7232 -6874 7252 -6860
rect 11886 -6874 11906 -6860
rect 5040 -6970 5110 -6900
rect 7030 -6970 7100 -6900
rect 12110 -700 14030 -580
rect 12600 -6000 13000 -700
rect 13200 -6000 13600 -700
rect 12110 -6200 14030 -6000
rect 12300 -6700 12700 -6200
rect 12900 -6700 13300 -6200
rect 13500 -6700 13900 -6200
rect 12110 -6900 14030 -6700
rect 19040 -580 21100 -520
rect 14232 -620 14252 -610
rect 18886 -620 18906 -610
rect 14232 -690 14240 -620
rect 18900 -690 18906 -620
rect 14232 -710 14252 -690
rect 18886 -710 18906 -690
rect 14165 -762 14231 -742
rect 14165 -6742 14231 -6722
rect 14323 -762 14389 -742
rect 14323 -6742 14389 -6722
rect 14481 -762 14547 -742
rect 14481 -6742 14547 -6722
rect 14639 -762 14705 -742
rect 14639 -6742 14705 -6722
rect 14797 -762 14863 -742
rect 14797 -6742 14863 -6722
rect 14955 -762 15021 -742
rect 14955 -6742 15021 -6722
rect 15113 -762 15179 -742
rect 15113 -6742 15179 -6722
rect 15271 -762 15337 -742
rect 15271 -6742 15337 -6722
rect 15429 -762 15495 -742
rect 15429 -6742 15495 -6722
rect 15587 -762 15653 -742
rect 15587 -6742 15653 -6722
rect 15745 -762 15811 -742
rect 15745 -6742 15811 -6722
rect 15903 -762 15969 -742
rect 15903 -6742 15969 -6722
rect 16061 -762 16127 -742
rect 16061 -6742 16127 -6722
rect 16219 -762 16285 -742
rect 16219 -6742 16285 -6722
rect 16377 -762 16443 -742
rect 16377 -6742 16443 -6722
rect 16535 -762 16601 -742
rect 16535 -6742 16601 -6722
rect 16693 -762 16759 -742
rect 16693 -6742 16759 -6722
rect 16851 -762 16917 -742
rect 16851 -6742 16917 -6722
rect 17009 -762 17075 -742
rect 17009 -6742 17075 -6722
rect 17167 -762 17233 -742
rect 17167 -6742 17233 -6722
rect 17325 -762 17391 -742
rect 17325 -6742 17391 -6722
rect 17483 -762 17549 -742
rect 17483 -6742 17549 -6722
rect 17641 -762 17707 -742
rect 17641 -6742 17707 -6722
rect 17799 -762 17865 -742
rect 17799 -6742 17865 -6722
rect 17957 -762 18023 -742
rect 17957 -6742 18023 -6722
rect 18115 -762 18181 -742
rect 18115 -6742 18181 -6722
rect 18273 -762 18339 -742
rect 18273 -6742 18339 -6722
rect 18431 -762 18497 -742
rect 18431 -6742 18497 -6722
rect 18589 -762 18655 -742
rect 18589 -6742 18655 -6722
rect 18747 -762 18813 -742
rect 18747 -6742 18813 -6722
rect 18905 -762 18971 -742
rect 18905 -6742 18971 -6722
rect 14232 -6790 14252 -6774
rect 18886 -6790 18906 -6774
rect 14232 -6860 14240 -6790
rect 18890 -6860 18906 -6790
rect 14232 -6874 14252 -6860
rect 18886 -6874 18906 -6860
rect 12040 -6970 12110 -6900
rect 12600 -12100 13000 -6900
rect 13200 -12100 13600 -6900
rect 14030 -6970 14100 -6900
rect 19110 -700 21030 -580
rect 19110 -6200 21030 -6000
rect 19300 -6700 19700 -6200
rect 19900 -6700 20300 -6200
rect 20500 -6700 20900 -6200
rect 19110 -6900 21030 -6700
rect 26040 -580 26110 -520
rect 21232 -620 21252 -610
rect 25886 -620 25906 -610
rect 21232 -690 21240 -620
rect 25900 -690 25906 -620
rect 21232 -710 21252 -690
rect 25886 -710 25906 -690
rect 21165 -762 21231 -742
rect 21165 -6742 21231 -6722
rect 21323 -762 21389 -742
rect 21323 -6742 21389 -6722
rect 21481 -762 21547 -742
rect 21481 -6742 21547 -6722
rect 21639 -762 21705 -742
rect 21639 -6742 21705 -6722
rect 21797 -762 21863 -742
rect 21797 -6742 21863 -6722
rect 21955 -762 22021 -742
rect 21955 -6742 22021 -6722
rect 22113 -762 22179 -742
rect 22113 -6742 22179 -6722
rect 22271 -762 22337 -742
rect 22271 -6742 22337 -6722
rect 22429 -762 22495 -742
rect 22429 -6742 22495 -6722
rect 22587 -762 22653 -742
rect 22587 -6742 22653 -6722
rect 22745 -762 22811 -742
rect 22745 -6742 22811 -6722
rect 22903 -762 22969 -742
rect 22903 -6742 22969 -6722
rect 23061 -762 23127 -742
rect 23061 -6742 23127 -6722
rect 23219 -762 23285 -742
rect 23219 -6742 23285 -6722
rect 23377 -762 23443 -742
rect 23377 -6742 23443 -6722
rect 23535 -762 23601 -742
rect 23535 -6742 23601 -6722
rect 23693 -762 23759 -742
rect 23693 -6742 23759 -6722
rect 23851 -762 23917 -742
rect 23851 -6742 23917 -6722
rect 24009 -762 24075 -742
rect 24009 -6742 24075 -6722
rect 24167 -762 24233 -742
rect 24167 -6742 24233 -6722
rect 24325 -762 24391 -742
rect 24325 -6742 24391 -6722
rect 24483 -762 24549 -742
rect 24483 -6742 24549 -6722
rect 24641 -762 24707 -742
rect 24641 -6742 24707 -6722
rect 24799 -762 24865 -742
rect 24799 -6742 24865 -6722
rect 24957 -762 25023 -742
rect 24957 -6742 25023 -6722
rect 25115 -762 25181 -742
rect 25115 -6742 25181 -6722
rect 25273 -762 25339 -742
rect 25273 -6742 25339 -6722
rect 25431 -762 25497 -742
rect 25431 -6742 25497 -6722
rect 25589 -762 25655 -742
rect 25589 -6742 25655 -6722
rect 25747 -762 25813 -742
rect 25747 -6742 25813 -6722
rect 25905 -762 25971 -742
rect 25905 -6742 25971 -6722
rect 21232 -6790 21252 -6774
rect 25886 -6790 25906 -6774
rect 21232 -6860 21240 -6790
rect 25890 -6860 25906 -6790
rect 21232 -6874 21252 -6860
rect 25886 -6874 25906 -6860
rect 19040 -6970 19110 -6900
rect 21030 -6970 21100 -6900
rect 26040 -6970 26110 -6900
rect 12600 -12300 13600 -12100
<< via2 >>
rect 240 6310 252 6380
rect 252 6310 4886 6380
rect 4886 6310 4900 6380
rect 165 885 231 2645
rect 323 3885 389 5645
rect 481 885 547 2645
rect 639 3885 705 5645
rect 797 885 863 2645
rect 955 3885 1021 5645
rect 1113 885 1179 2645
rect 1271 3885 1337 5645
rect 1429 885 1495 2645
rect 1587 3885 1653 5645
rect 1745 885 1811 2645
rect 1903 3885 1969 5645
rect 2061 885 2127 2645
rect 2219 3885 2285 5645
rect 2377 885 2443 2645
rect 2535 3885 2601 5645
rect 2693 885 2759 2645
rect 2851 3885 2917 5645
rect 3009 885 3075 2645
rect 3167 3885 3233 5645
rect 3325 885 3391 2645
rect 3483 3885 3549 5645
rect 3641 885 3707 2645
rect 3799 3885 3865 5645
rect 3957 885 4023 2645
rect 4115 3885 4181 5645
rect 4273 885 4339 2645
rect 4431 3885 4497 5645
rect 4589 885 4655 2645
rect 4747 3885 4813 5645
rect 4905 885 4971 2645
rect 240 140 252 210
rect 252 140 4886 210
rect 4886 140 4890 210
rect 7240 6310 7252 6380
rect 7252 6310 11886 6380
rect 11886 6310 11900 6380
rect 7165 885 7231 2645
rect 7323 3885 7389 5645
rect 7481 885 7547 2645
rect 7639 3885 7705 5645
rect 7797 885 7863 2645
rect 7955 3885 8021 5645
rect 8113 885 8179 2645
rect 8271 3885 8337 5645
rect 8429 885 8495 2645
rect 8587 3885 8653 5645
rect 8745 885 8811 2645
rect 8903 3885 8969 5645
rect 9061 885 9127 2645
rect 9219 3885 9285 5645
rect 9377 885 9443 2645
rect 9535 3885 9601 5645
rect 9693 885 9759 2645
rect 9851 3885 9917 5645
rect 10009 885 10075 2645
rect 10167 3885 10233 5645
rect 10325 885 10391 2645
rect 10483 3885 10549 5645
rect 10641 885 10707 2645
rect 10799 3885 10865 5645
rect 10957 885 11023 2645
rect 11115 3885 11181 5645
rect 11273 885 11339 2645
rect 11431 3885 11497 5645
rect 11589 885 11655 2645
rect 11747 3885 11813 5645
rect 11905 885 11971 2645
rect 7240 140 7252 210
rect 7252 140 11886 210
rect 11886 140 11890 210
rect 14240 6310 14252 6380
rect 14252 6310 18886 6380
rect 18886 6310 18900 6380
rect 14165 885 14231 2645
rect 14323 3885 14389 5645
rect 14481 885 14547 2645
rect 14639 3885 14705 5645
rect 14797 885 14863 2645
rect 14955 3885 15021 5645
rect 15113 885 15179 2645
rect 15271 3885 15337 5645
rect 15429 885 15495 2645
rect 15587 3885 15653 5645
rect 15745 885 15811 2645
rect 15903 3885 15969 5645
rect 16061 885 16127 2645
rect 16219 3885 16285 5645
rect 16377 885 16443 2645
rect 16535 3885 16601 5645
rect 16693 885 16759 2645
rect 16851 3885 16917 5645
rect 17009 885 17075 2645
rect 17167 3885 17233 5645
rect 17325 885 17391 2645
rect 17483 3885 17549 5645
rect 17641 885 17707 2645
rect 17799 3885 17865 5645
rect 17957 885 18023 2645
rect 18115 3885 18181 5645
rect 18273 885 18339 2645
rect 18431 3885 18497 5645
rect 18589 885 18655 2645
rect 18747 3885 18813 5645
rect 18905 885 18971 2645
rect 14240 140 14252 210
rect 14252 140 18886 210
rect 18886 140 18890 210
rect 21240 6310 21252 6380
rect 21252 6310 25886 6380
rect 25886 6310 25900 6380
rect 21165 885 21231 2645
rect 21323 3885 21389 5645
rect 21481 885 21547 2645
rect 21639 3885 21705 5645
rect 21797 885 21863 2645
rect 21955 3885 22021 5645
rect 22113 885 22179 2645
rect 22271 3885 22337 5645
rect 22429 885 22495 2645
rect 22587 3885 22653 5645
rect 22745 885 22811 2645
rect 22903 3885 22969 5645
rect 23061 885 23127 2645
rect 23219 3885 23285 5645
rect 23377 885 23443 2645
rect 23535 3885 23601 5645
rect 23693 885 23759 2645
rect 23851 3885 23917 5645
rect 24009 885 24075 2645
rect 24167 3885 24233 5645
rect 24325 885 24391 2645
rect 24483 3885 24549 5645
rect 24641 885 24707 2645
rect 24799 3885 24865 5645
rect 24957 885 25023 2645
rect 25115 3885 25181 5645
rect 25273 885 25339 2645
rect 25431 3885 25497 5645
rect 25589 885 25655 2645
rect 25747 3885 25813 5645
rect 25905 885 25971 2645
rect 21240 140 21252 210
rect 21252 140 25886 210
rect 25886 140 25890 210
rect 240 -690 252 -620
rect 252 -690 4886 -620
rect 4886 -690 4900 -620
rect 165 -6115 231 -4355
rect 323 -3115 389 -1355
rect 481 -6115 547 -4355
rect 639 -3115 705 -1355
rect 797 -6115 863 -4355
rect 955 -3115 1021 -1355
rect 1113 -6115 1179 -4355
rect 1271 -3115 1337 -1355
rect 1429 -6115 1495 -4355
rect 1587 -3115 1653 -1355
rect 1745 -6115 1811 -4355
rect 1903 -3115 1969 -1355
rect 2061 -6115 2127 -4355
rect 2219 -3115 2285 -1355
rect 2377 -6115 2443 -4355
rect 2535 -3115 2601 -1355
rect 2693 -6115 2759 -4355
rect 2851 -3115 2917 -1355
rect 3009 -6115 3075 -4355
rect 3167 -3115 3233 -1355
rect 3325 -6115 3391 -4355
rect 3483 -3115 3549 -1355
rect 3641 -6115 3707 -4355
rect 3799 -3115 3865 -1355
rect 3957 -6115 4023 -4355
rect 4115 -3115 4181 -1355
rect 4273 -6115 4339 -4355
rect 4431 -3115 4497 -1355
rect 4589 -6115 4655 -4355
rect 4747 -3115 4813 -1355
rect 4905 -6115 4971 -4355
rect 240 -6860 252 -6790
rect 252 -6860 4886 -6790
rect 4886 -6860 4890 -6790
rect 7240 -690 7252 -620
rect 7252 -690 11886 -620
rect 11886 -690 11900 -620
rect 7165 -6115 7231 -4355
rect 7323 -3115 7389 -1355
rect 7481 -6115 7547 -4355
rect 7639 -3115 7705 -1355
rect 7797 -6115 7863 -4355
rect 7955 -3115 8021 -1355
rect 8113 -6115 8179 -4355
rect 8271 -3115 8337 -1355
rect 8429 -6115 8495 -4355
rect 8587 -3115 8653 -1355
rect 8745 -6115 8811 -4355
rect 8903 -3115 8969 -1355
rect 9061 -6115 9127 -4355
rect 9219 -3115 9285 -1355
rect 9377 -6115 9443 -4355
rect 9535 -3115 9601 -1355
rect 9693 -6115 9759 -4355
rect 9851 -3115 9917 -1355
rect 10009 -6115 10075 -4355
rect 10167 -3115 10233 -1355
rect 10325 -6115 10391 -4355
rect 10483 -3115 10549 -1355
rect 10641 -6115 10707 -4355
rect 10799 -3115 10865 -1355
rect 10957 -6115 11023 -4355
rect 11115 -3115 11181 -1355
rect 11273 -6115 11339 -4355
rect 11431 -3115 11497 -1355
rect 11589 -6115 11655 -4355
rect 11747 -3115 11813 -1355
rect 11905 -6115 11971 -4355
rect 7240 -6860 7252 -6790
rect 7252 -6860 11886 -6790
rect 11886 -6860 11890 -6790
rect 14240 -690 14252 -620
rect 14252 -690 18886 -620
rect 18886 -690 18900 -620
rect 14165 -6115 14231 -4355
rect 14323 -3115 14389 -1355
rect 14481 -6115 14547 -4355
rect 14639 -3115 14705 -1355
rect 14797 -6115 14863 -4355
rect 14955 -3115 15021 -1355
rect 15113 -6115 15179 -4355
rect 15271 -3115 15337 -1355
rect 15429 -6115 15495 -4355
rect 15587 -3115 15653 -1355
rect 15745 -6115 15811 -4355
rect 15903 -3115 15969 -1355
rect 16061 -6115 16127 -4355
rect 16219 -3115 16285 -1355
rect 16377 -6115 16443 -4355
rect 16535 -3115 16601 -1355
rect 16693 -6115 16759 -4355
rect 16851 -3115 16917 -1355
rect 17009 -6115 17075 -4355
rect 17167 -3115 17233 -1355
rect 17325 -6115 17391 -4355
rect 17483 -3115 17549 -1355
rect 17641 -6115 17707 -4355
rect 17799 -3115 17865 -1355
rect 17957 -6115 18023 -4355
rect 18115 -3115 18181 -1355
rect 18273 -6115 18339 -4355
rect 18431 -3115 18497 -1355
rect 18589 -6115 18655 -4355
rect 18747 -3115 18813 -1355
rect 18905 -6115 18971 -4355
rect 14240 -6860 14252 -6790
rect 14252 -6860 18886 -6790
rect 18886 -6860 18890 -6790
rect 21240 -690 21252 -620
rect 21252 -690 25886 -620
rect 25886 -690 25900 -620
rect 21165 -6115 21231 -4355
rect 21323 -3115 21389 -1355
rect 21481 -6115 21547 -4355
rect 21639 -3115 21705 -1355
rect 21797 -6115 21863 -4355
rect 21955 -3115 22021 -1355
rect 22113 -6115 22179 -4355
rect 22271 -3115 22337 -1355
rect 22429 -6115 22495 -4355
rect 22587 -3115 22653 -1355
rect 22745 -6115 22811 -4355
rect 22903 -3115 22969 -1355
rect 23061 -6115 23127 -4355
rect 23219 -3115 23285 -1355
rect 23377 -6115 23443 -4355
rect 23535 -3115 23601 -1355
rect 23693 -6115 23759 -4355
rect 23851 -3115 23917 -1355
rect 24009 -6115 24075 -4355
rect 24167 -3115 24233 -1355
rect 24325 -6115 24391 -4355
rect 24483 -3115 24549 -1355
rect 24641 -6115 24707 -4355
rect 24799 -3115 24865 -1355
rect 24957 -6115 25023 -4355
rect 25115 -3115 25181 -1355
rect 25273 -6115 25339 -4355
rect 25431 -3115 25497 -1355
rect 25589 -6115 25655 -4355
rect 25747 -3115 25813 -1355
rect 25905 -6115 25971 -4355
rect 21240 -6860 21252 -6790
rect 21252 -6860 25886 -6790
rect 25886 -6860 25890 -6790
<< metal3 >>
rect 100 6380 5100 6500
rect 100 6310 240 6380
rect 4900 6310 5100 6380
rect 100 6300 5100 6310
rect 7100 6380 12100 6500
rect 7100 6310 7240 6380
rect 11900 6310 12100 6380
rect 7100 6300 12100 6310
rect 14100 6380 19100 6500
rect 14100 6310 14240 6380
rect 18900 6310 19100 6380
rect 14100 6300 19100 6310
rect 21100 6380 26100 6500
rect 21100 6310 21240 6380
rect 25900 6310 26100 6380
rect 21100 6300 26100 6310
rect 30 5645 5110 5800
rect 30 5600 323 5645
rect 389 5600 639 5645
rect 705 5600 955 5645
rect 1021 5600 1271 5645
rect 1337 5600 1587 5645
rect 30 4000 200 5600
rect 1400 4000 1587 5600
rect 30 3885 323 4000
rect 389 3885 639 4000
rect 705 3885 955 4000
rect 1021 3885 1271 4000
rect 1337 3885 1587 4000
rect 1653 3885 1903 5645
rect 1969 3885 2219 5645
rect 2285 3885 2535 5645
rect 2601 3885 2851 5645
rect 2917 3885 3167 5645
rect 3233 3885 3483 5645
rect 3549 3885 3799 5645
rect 3865 3885 4115 5645
rect 4181 3885 4431 5645
rect 4497 3885 4747 5645
rect 4813 3885 5110 5645
rect 30 3800 5110 3885
rect 7030 5645 12110 5800
rect 7030 5600 7323 5645
rect 7389 5600 7639 5645
rect 7705 5600 7955 5645
rect 8021 5600 8271 5645
rect 8337 5600 8587 5645
rect 7030 4000 7200 5600
rect 8400 4000 8587 5600
rect 7030 3885 7323 4000
rect 7389 3885 7639 4000
rect 7705 3885 7955 4000
rect 8021 3885 8271 4000
rect 8337 3885 8587 4000
rect 8653 3885 8903 5645
rect 8969 3885 9219 5645
rect 9285 3885 9535 5645
rect 9601 3885 9851 5645
rect 9917 3885 10167 5645
rect 10233 3885 10483 5645
rect 10549 3885 10799 5645
rect 10865 3885 11115 5645
rect 11181 3885 11431 5645
rect 11497 3885 11747 5645
rect 11813 3885 12110 5645
rect 7030 3800 12110 3885
rect 14030 5645 19110 5800
rect 14030 5600 14323 5645
rect 14389 5600 14639 5645
rect 14705 5600 14955 5645
rect 15021 5600 15271 5645
rect 15337 5600 15587 5645
rect 14030 4000 14200 5600
rect 15400 4000 15587 5600
rect 14030 3885 14323 4000
rect 14389 3885 14639 4000
rect 14705 3885 14955 4000
rect 15021 3885 15271 4000
rect 15337 3885 15587 4000
rect 15653 3885 15903 5645
rect 15969 3885 16219 5645
rect 16285 3885 16535 5645
rect 16601 3885 16851 5645
rect 16917 3885 17167 5645
rect 17233 3885 17483 5645
rect 17549 3885 17799 5645
rect 17865 3885 18115 5645
rect 18181 3885 18431 5645
rect 18497 3885 18747 5645
rect 18813 3885 19110 5645
rect 14030 3800 19110 3885
rect 21030 5645 26110 5800
rect 21030 5600 21323 5645
rect 21389 5600 21639 5645
rect 21705 5600 21955 5645
rect 22021 5600 22271 5645
rect 22337 5600 22587 5645
rect 21030 4000 21200 5600
rect 22400 4000 22587 5600
rect 21030 3885 21323 4000
rect 21389 3885 21639 4000
rect 21705 3885 21955 4000
rect 22021 3885 22271 4000
rect 22337 3885 22587 4000
rect 22653 3885 22903 5645
rect 22969 3885 23219 5645
rect 23285 3885 23535 5645
rect 23601 3885 23851 5645
rect 23917 3885 24167 5645
rect 24233 3885 24483 5645
rect 24549 3885 24799 5645
rect 24865 3885 25115 5645
rect 25181 3885 25431 5645
rect 25497 3885 25747 5645
rect 25813 3885 26110 5645
rect 21030 3800 26110 3885
rect 30 2645 5110 2800
rect 30 885 165 2645
rect 231 2600 481 2645
rect 547 2600 797 2645
rect 863 2600 1113 2645
rect 1179 2600 1429 2645
rect 1400 1000 1429 2600
rect 231 885 481 1000
rect 547 885 797 1000
rect 863 885 1113 1000
rect 1179 885 1429 1000
rect 1495 885 1745 2645
rect 1811 885 2061 2645
rect 2127 885 2377 2645
rect 2443 885 2693 2645
rect 2759 885 3009 2645
rect 3075 885 3325 2645
rect 3391 885 3641 2645
rect 3707 885 3957 2645
rect 4023 885 4273 2645
rect 4339 885 4589 2645
rect 4655 885 4905 2645
rect 4971 885 5110 2645
rect 30 800 5110 885
rect 7030 2645 12110 2800
rect 7030 885 7165 2645
rect 7231 2600 7481 2645
rect 7547 2600 7797 2645
rect 7863 2600 8113 2645
rect 8179 2600 8429 2645
rect 8400 1000 8429 2600
rect 7231 885 7481 1000
rect 7547 885 7797 1000
rect 7863 885 8113 1000
rect 8179 885 8429 1000
rect 8495 885 8745 2645
rect 8811 885 9061 2645
rect 9127 885 9377 2645
rect 9443 885 9693 2645
rect 9759 885 10009 2645
rect 10075 885 10325 2645
rect 10391 885 10641 2645
rect 10707 885 10957 2645
rect 11023 885 11273 2645
rect 11339 885 11589 2645
rect 11655 885 11905 2645
rect 11971 885 12110 2645
rect 7030 800 12110 885
rect 14030 2645 19110 2800
rect 14030 885 14165 2645
rect 14231 2600 14481 2645
rect 14547 2600 14797 2645
rect 14863 2600 15113 2645
rect 15179 2600 15429 2645
rect 15400 1000 15429 2600
rect 14231 885 14481 1000
rect 14547 885 14797 1000
rect 14863 885 15113 1000
rect 15179 885 15429 1000
rect 15495 885 15745 2645
rect 15811 885 16061 2645
rect 16127 885 16377 2645
rect 16443 885 16693 2645
rect 16759 885 17009 2645
rect 17075 885 17325 2645
rect 17391 885 17641 2645
rect 17707 885 17957 2645
rect 18023 885 18273 2645
rect 18339 885 18589 2645
rect 18655 885 18905 2645
rect 18971 885 19110 2645
rect 14030 800 19110 885
rect 21030 2645 26110 2800
rect 21030 885 21165 2645
rect 21231 2600 21481 2645
rect 21547 2600 21797 2645
rect 21863 2600 22113 2645
rect 22179 2600 22429 2645
rect 22400 1000 22429 2600
rect 21231 885 21481 1000
rect 21547 885 21797 1000
rect 21863 885 22113 1000
rect 22179 885 22429 1000
rect 22495 885 22745 2645
rect 22811 885 23061 2645
rect 23127 885 23377 2645
rect 23443 885 23693 2645
rect 23759 885 24009 2645
rect 24075 885 24325 2645
rect 24391 885 24641 2645
rect 24707 885 24957 2645
rect 25023 885 25273 2645
rect 25339 885 25589 2645
rect 25655 885 25905 2645
rect 25971 885 26110 2645
rect 21030 800 26110 885
rect 1900 300 4100 400
rect 15900 300 18100 400
rect 1700 230 2000 300
rect 100 210 2000 230
rect 4000 230 4300 300
rect 8700 230 11300 300
rect 15700 230 16000 300
rect 4000 210 5100 230
rect 100 140 240 210
rect 4890 200 5100 210
rect 7100 210 12100 230
rect 7100 200 7240 210
rect 4890 180 6700 200
rect 4890 140 6320 180
rect 100 100 2000 140
rect 4000 100 6320 140
rect 100 30 6320 100
rect 1700 -100 4300 30
rect 4500 20 6320 30
rect 6680 20 6700 180
rect 4500 0 6700 20
rect 6900 140 7240 200
rect 11890 200 12100 210
rect 14100 210 16000 230
rect 18000 230 18300 300
rect 22700 230 25300 300
rect 18000 210 19100 230
rect 14100 200 14240 210
rect 11890 180 13700 200
rect 11890 140 13320 180
rect 6900 20 13320 140
rect 13680 20 13700 180
rect 6900 0 13700 20
rect 13900 140 14240 200
rect 18890 200 19100 210
rect 21100 210 26100 230
rect 21100 200 21240 210
rect 18890 180 20700 200
rect 18890 140 20320 180
rect 13900 100 16000 140
rect 18000 100 20320 140
rect 13900 30 20320 100
rect 13900 20 14220 30
rect 15700 20 20320 30
rect 20680 20 20700 180
rect 13900 0 14200 20
rect 15700 0 20700 20
rect 20900 140 21240 200
rect 25890 140 26100 210
rect 20900 30 26100 140
rect 6900 -200 7100 0
rect 8700 -100 11300 0
rect 13900 -100 14100 0
rect 15700 -100 18300 0
rect 20900 -100 21200 30
rect 22700 -100 25300 30
rect 5900 -400 7100 -200
rect 12900 -300 14100 -100
rect 19900 -300 21200 -100
rect 1700 -500 4300 -400
rect 5900 -500 6100 -400
rect 8700 -500 11300 -400
rect 12900 -500 13100 -300
rect 15700 -500 18300 -400
rect 19900 -500 20100 -300
rect 22700 -500 25300 -400
rect 100 -620 2000 -500
rect 4000 -620 6100 -500
rect 100 -690 240 -620
rect 4900 -690 6100 -620
rect 100 -700 2000 -690
rect 4000 -700 6100 -690
rect 6300 -520 13100 -500
rect 6300 -680 6320 -520
rect 6680 -620 13100 -520
rect 6680 -680 7240 -620
rect 6300 -690 7240 -680
rect 11900 -690 13100 -620
rect 6300 -700 13100 -690
rect 13300 -520 16000 -500
rect 13300 -680 13320 -520
rect 13680 -620 16000 -520
rect 18000 -620 20100 -500
rect 13680 -680 14240 -620
rect 13300 -690 14240 -680
rect 18900 -690 20100 -620
rect 13300 -700 16000 -690
rect 18000 -700 20100 -690
rect 20300 -520 26100 -500
rect 20300 -680 20320 -520
rect 20680 -620 26100 -520
rect 20680 -680 21240 -620
rect 20300 -690 21240 -680
rect 25900 -690 26100 -620
rect 20300 -700 26100 -690
rect 1700 -800 4300 -700
rect 8700 -800 11300 -700
rect 15700 -800 18300 -700
rect 22700 -800 25300 -700
rect 30 -1355 5110 -1200
rect 30 -3115 323 -1355
rect 389 -3115 639 -1355
rect 705 -3115 955 -1355
rect 1021 -3115 1271 -1355
rect 1337 -3115 1587 -1355
rect 1653 -3115 1903 -1355
rect 1969 -3115 2219 -1355
rect 2285 -1400 2535 -1355
rect 2601 -1400 2851 -1355
rect 2917 -1400 3167 -1355
rect 3233 -1400 3483 -1355
rect 3549 -1400 3799 -1355
rect 2285 -3000 2400 -1400
rect 3600 -3000 3799 -1400
rect 2285 -3115 2535 -3000
rect 2601 -3115 2851 -3000
rect 2917 -3115 3167 -3000
rect 3233 -3115 3483 -3000
rect 3549 -3115 3799 -3000
rect 3865 -3115 4115 -1355
rect 4181 -3115 4431 -1355
rect 4497 -3115 4747 -1355
rect 4813 -3115 5110 -1355
rect 30 -3200 5110 -3115
rect 7030 -1355 12110 -1200
rect 7030 -3115 7323 -1355
rect 7389 -3115 7639 -1355
rect 7705 -3115 7955 -1355
rect 8021 -3115 8271 -1355
rect 8337 -3115 8587 -1355
rect 8653 -3115 8903 -1355
rect 8969 -3115 9219 -1355
rect 9285 -1400 9535 -1355
rect 9601 -1400 9851 -1355
rect 9917 -1400 10167 -1355
rect 10233 -1400 10483 -1355
rect 10549 -1400 10799 -1355
rect 9285 -3000 9400 -1400
rect 10600 -3000 10799 -1400
rect 9285 -3115 9535 -3000
rect 9601 -3115 9851 -3000
rect 9917 -3115 10167 -3000
rect 10233 -3115 10483 -3000
rect 10549 -3115 10799 -3000
rect 10865 -3115 11115 -1355
rect 11181 -3115 11431 -1355
rect 11497 -3115 11747 -1355
rect 11813 -3115 12110 -1355
rect 7030 -3200 12110 -3115
rect 14030 -1355 19110 -1200
rect 14030 -3115 14323 -1355
rect 14389 -3115 14639 -1355
rect 14705 -3115 14955 -1355
rect 15021 -3115 15271 -1355
rect 15337 -3115 15587 -1355
rect 15653 -3115 15903 -1355
rect 15969 -3115 16219 -1355
rect 16285 -1400 16535 -1355
rect 16601 -1400 16851 -1355
rect 16917 -1400 17167 -1355
rect 17233 -1400 17483 -1355
rect 17549 -1400 17799 -1355
rect 16285 -3000 16400 -1400
rect 17600 -3000 17799 -1400
rect 16285 -3115 16535 -3000
rect 16601 -3115 16851 -3000
rect 16917 -3115 17167 -3000
rect 17233 -3115 17483 -3000
rect 17549 -3115 17799 -3000
rect 17865 -3115 18115 -1355
rect 18181 -3115 18431 -1355
rect 18497 -3115 18747 -1355
rect 18813 -3115 19110 -1355
rect 14030 -3200 19110 -3115
rect 21030 -1355 26110 -1200
rect 21030 -3115 21323 -1355
rect 21389 -3115 21639 -1355
rect 21705 -3115 21955 -1355
rect 22021 -3115 22271 -1355
rect 22337 -3115 22587 -1355
rect 22653 -3115 22903 -1355
rect 22969 -3115 23219 -1355
rect 23285 -1400 23535 -1355
rect 23601 -1400 23851 -1355
rect 23917 -1400 24167 -1355
rect 24233 -1400 24483 -1355
rect 24549 -1400 24799 -1355
rect 23285 -3000 23400 -1400
rect 24600 -3000 24799 -1400
rect 23285 -3115 23535 -3000
rect 23601 -3115 23851 -3000
rect 23917 -3115 24167 -3000
rect 24233 -3115 24483 -3000
rect 24549 -3115 24799 -3000
rect 24865 -3115 25115 -1355
rect 25181 -3115 25431 -1355
rect 25497 -3115 25747 -1355
rect 25813 -3115 26110 -1355
rect 21030 -3200 26110 -3115
rect 30 -4355 6200 -4200
rect 30 -6115 165 -4355
rect 231 -6115 481 -4355
rect 547 -6115 797 -4355
rect 863 -6115 1113 -4355
rect 1179 -6115 1429 -4355
rect 1495 -6115 1745 -4355
rect 1811 -6115 2061 -4355
rect 2127 -6115 2377 -4355
rect 2443 -6115 2693 -4355
rect 2759 -6115 3009 -4355
rect 3075 -6115 3325 -4355
rect 3391 -6115 3641 -4355
rect 3707 -6115 3957 -4355
rect 4023 -6115 4273 -4355
rect 4339 -6115 4589 -4355
rect 4655 -4400 4905 -4355
rect 4971 -4400 6200 -4355
rect 5800 -6000 6200 -4400
rect 4655 -6115 4905 -6000
rect 4971 -6115 6200 -6000
rect 30 -6200 6200 -6115
rect 7030 -4355 13200 -4200
rect 7030 -6115 7165 -4355
rect 7231 -6115 7481 -4355
rect 7547 -6115 7797 -4355
rect 7863 -6115 8113 -4355
rect 8179 -6115 8429 -4355
rect 8495 -6115 8745 -4355
rect 8811 -6115 9061 -4355
rect 9127 -6115 9377 -4355
rect 9443 -6115 9693 -4355
rect 9759 -6115 10009 -4355
rect 10075 -6115 10325 -4355
rect 10391 -6115 10641 -4355
rect 10707 -6115 10957 -4355
rect 11023 -6115 11273 -4355
rect 11339 -6115 11589 -4355
rect 11655 -4400 11905 -4355
rect 11971 -4400 13200 -4355
rect 12800 -6000 13200 -4400
rect 11655 -6115 11905 -6000
rect 11971 -6115 13200 -6000
rect 7030 -6200 13200 -6115
rect 14030 -4355 20200 -4200
rect 14030 -6115 14165 -4355
rect 14231 -6115 14481 -4355
rect 14547 -6115 14797 -4355
rect 14863 -6115 15113 -4355
rect 15179 -6115 15429 -4355
rect 15495 -6115 15745 -4355
rect 15811 -6115 16061 -4355
rect 16127 -6115 16377 -4355
rect 16443 -6115 16693 -4355
rect 16759 -6115 17009 -4355
rect 17075 -6115 17325 -4355
rect 17391 -6115 17641 -4355
rect 17707 -6115 17957 -4355
rect 18023 -6115 18273 -4355
rect 18339 -6115 18589 -4355
rect 18655 -4400 18905 -4355
rect 18971 -4400 20200 -4355
rect 19800 -6000 20200 -4400
rect 18655 -6115 18905 -6000
rect 18971 -6115 20200 -6000
rect 14030 -6200 20200 -6115
rect 21030 -4355 27200 -4200
rect 21030 -6115 21165 -4355
rect 21231 -6115 21481 -4355
rect 21547 -6115 21797 -4355
rect 21863 -6115 22113 -4355
rect 22179 -6115 22429 -4355
rect 22495 -6115 22745 -4355
rect 22811 -6115 23061 -4355
rect 23127 -6115 23377 -4355
rect 23443 -6115 23693 -4355
rect 23759 -6115 24009 -4355
rect 24075 -6115 24325 -4355
rect 24391 -6115 24641 -4355
rect 24707 -6115 24957 -4355
rect 25023 -6115 25273 -4355
rect 25339 -6115 25589 -4355
rect 25655 -4400 25905 -4355
rect 25971 -4400 27200 -4355
rect 26800 -6000 27200 -4400
rect 25655 -6115 25905 -6000
rect 25971 -6115 27200 -6000
rect 21030 -6200 27200 -6115
rect 100 -6790 5100 -6770
rect 100 -6860 240 -6790
rect 4890 -6860 5100 -6790
rect 100 -6970 5100 -6860
rect 7100 -6790 12100 -6770
rect 7100 -6860 7240 -6790
rect 11890 -6860 12100 -6790
rect 7100 -6970 12100 -6860
rect 14100 -6790 19100 -6770
rect 14100 -6860 14240 -6790
rect 18890 -6860 19100 -6790
rect 14100 -6970 19100 -6860
rect 21100 -6790 26100 -6770
rect 21100 -6860 21240 -6790
rect 25890 -6860 26100 -6790
rect 21100 -6970 26100 -6860
<< via3 >>
rect 200 4000 323 5600
rect 323 4000 389 5600
rect 389 4000 639 5600
rect 639 4000 705 5600
rect 705 4000 955 5600
rect 955 4000 1021 5600
rect 1021 4000 1271 5600
rect 1271 4000 1337 5600
rect 1337 4000 1400 5600
rect 7200 4000 7323 5600
rect 7323 4000 7389 5600
rect 7389 4000 7639 5600
rect 7639 4000 7705 5600
rect 7705 4000 7955 5600
rect 7955 4000 8021 5600
rect 8021 4000 8271 5600
rect 8271 4000 8337 5600
rect 8337 4000 8400 5600
rect 14200 4000 14323 5600
rect 14323 4000 14389 5600
rect 14389 4000 14639 5600
rect 14639 4000 14705 5600
rect 14705 4000 14955 5600
rect 14955 4000 15021 5600
rect 15021 4000 15271 5600
rect 15271 4000 15337 5600
rect 15337 4000 15400 5600
rect 21200 4000 21323 5600
rect 21323 4000 21389 5600
rect 21389 4000 21639 5600
rect 21639 4000 21705 5600
rect 21705 4000 21955 5600
rect 21955 4000 22021 5600
rect 22021 4000 22271 5600
rect 22271 4000 22337 5600
rect 22337 4000 22400 5600
rect 200 1000 231 2600
rect 231 1000 481 2600
rect 481 1000 547 2600
rect 547 1000 797 2600
rect 797 1000 863 2600
rect 863 1000 1113 2600
rect 1113 1000 1179 2600
rect 1179 1000 1400 2600
rect 7200 1000 7231 2600
rect 7231 1000 7481 2600
rect 7481 1000 7547 2600
rect 7547 1000 7797 2600
rect 7797 1000 7863 2600
rect 7863 1000 8113 2600
rect 8113 1000 8179 2600
rect 8179 1000 8400 2600
rect 14200 1000 14231 2600
rect 14231 1000 14481 2600
rect 14481 1000 14547 2600
rect 14547 1000 14797 2600
rect 14797 1000 14863 2600
rect 14863 1000 15113 2600
rect 15113 1000 15179 2600
rect 15179 1000 15400 2600
rect 21200 1000 21231 2600
rect 21231 1000 21481 2600
rect 21481 1000 21547 2600
rect 21547 1000 21797 2600
rect 21797 1000 21863 2600
rect 21863 1000 22113 2600
rect 22113 1000 22179 2600
rect 22179 1000 22400 2600
rect 2000 210 4000 300
rect 2000 140 4000 210
rect 2000 100 4000 140
rect 6320 20 6680 180
rect 16000 210 18000 300
rect 13320 20 13680 180
rect 16000 140 18000 210
rect 16000 100 18000 140
rect 20320 20 20680 180
rect 2000 -620 4000 -500
rect 2000 -690 4000 -620
rect 2000 -700 4000 -690
rect 6320 -680 6680 -520
rect 13320 -680 13680 -520
rect 16000 -620 18000 -500
rect 16000 -690 18000 -620
rect 16000 -700 18000 -690
rect 20320 -680 20680 -520
rect 2400 -3000 2535 -1400
rect 2535 -3000 2601 -1400
rect 2601 -3000 2851 -1400
rect 2851 -3000 2917 -1400
rect 2917 -3000 3167 -1400
rect 3167 -3000 3233 -1400
rect 3233 -3000 3483 -1400
rect 3483 -3000 3549 -1400
rect 3549 -3000 3600 -1400
rect 9400 -3000 9535 -1400
rect 9535 -3000 9601 -1400
rect 9601 -3000 9851 -1400
rect 9851 -3000 9917 -1400
rect 9917 -3000 10167 -1400
rect 10167 -3000 10233 -1400
rect 10233 -3000 10483 -1400
rect 10483 -3000 10549 -1400
rect 10549 -3000 10600 -1400
rect 16400 -3000 16535 -1400
rect 16535 -3000 16601 -1400
rect 16601 -3000 16851 -1400
rect 16851 -3000 16917 -1400
rect 16917 -3000 17167 -1400
rect 17167 -3000 17233 -1400
rect 17233 -3000 17483 -1400
rect 17483 -3000 17549 -1400
rect 17549 -3000 17600 -1400
rect 23400 -3000 23535 -1400
rect 23535 -3000 23601 -1400
rect 23601 -3000 23851 -1400
rect 23851 -3000 23917 -1400
rect 23917 -3000 24167 -1400
rect 24167 -3000 24233 -1400
rect 24233 -3000 24483 -1400
rect 24483 -3000 24549 -1400
rect 24549 -3000 24600 -1400
rect 4600 -6000 4655 -4400
rect 4655 -6000 4905 -4400
rect 4905 -6000 4971 -4400
rect 4971 -6000 5800 -4400
rect 11600 -6000 11655 -4400
rect 11655 -6000 11905 -4400
rect 11905 -6000 11971 -4400
rect 11971 -6000 12800 -4400
rect 18600 -6000 18655 -4400
rect 18655 -6000 18905 -4400
rect 18905 -6000 18971 -4400
rect 18971 -6000 19800 -4400
rect 25600 -6000 25655 -4400
rect 25655 -6000 25905 -4400
rect 25905 -6000 25971 -4400
rect 25971 -6000 26800 -4400
<< metal4 >>
rect 4400 11000 6000 11200
rect 4400 9600 4600 11000
rect 5800 9600 6000 11000
rect 0 8000 1600 8200
rect 0 6600 200 8000
rect 1400 6600 1600 8000
rect 0 5600 1600 6600
rect 0 4000 200 5600
rect 1400 4000 1600 5600
rect 0 3800 1600 4000
rect 0 2600 1600 2800
rect 0 1000 200 2600
rect 1400 1000 1600 2600
rect 0 -10000 1600 1000
rect 1900 400 4100 500
rect 1900 100 2000 400
rect 4000 100 4100 400
rect 1900 0 4100 100
rect 1900 -500 4100 -400
rect 1900 -800 2000 -500
rect 4000 -800 4100 -500
rect 1900 -900 4100 -800
rect 2200 -1400 3800 -1200
rect 2200 -3000 2400 -1400
rect 3600 -3000 3800 -1400
rect 2200 -7000 3800 -3000
rect 4400 -4400 6000 9600
rect 11400 11000 13000 11200
rect 11400 9600 11600 11000
rect 12800 9600 13000 11000
rect 7000 8000 8600 8200
rect 7000 6600 7200 8000
rect 8400 6600 8600 8000
rect 7000 5600 8600 6600
rect 7000 4000 7200 5600
rect 8400 4000 8600 5600
rect 7000 3800 8600 4000
rect 7000 2600 8600 2800
rect 7000 1000 7200 2600
rect 8400 1000 8600 2600
rect 6300 180 6700 200
rect 6300 20 6320 180
rect 6680 20 6700 180
rect 6300 -520 6700 20
rect 6300 -680 6320 -520
rect 6680 -680 6700 -520
rect 6300 -700 6700 -680
rect 4400 -6000 4600 -4400
rect 5800 -6000 6000 -4400
rect 4400 -6200 6000 -6000
rect 2200 -8400 2400 -7000
rect 3600 -8400 3800 -7000
rect 2200 -8600 3800 -8400
rect 0 -11400 200 -10000
rect 1400 -11400 1600 -10000
rect 0 -11600 1600 -11400
rect 7000 -10000 8600 1000
rect 9200 -1400 10800 -1200
rect 9200 -3000 9400 -1400
rect 10600 -3000 10800 -1400
rect 9200 -7000 10800 -3000
rect 11400 -4400 13000 9600
rect 18400 11000 20000 11200
rect 18400 9600 18600 11000
rect 19800 9600 20000 11000
rect 14000 8000 15600 8200
rect 14000 6600 14200 8000
rect 15400 6600 15600 8000
rect 14000 5600 15600 6600
rect 14000 4000 14200 5600
rect 15400 4000 15600 5600
rect 14000 3800 15600 4000
rect 14000 2600 15600 2800
rect 14000 1000 14200 2600
rect 15400 1000 15600 2600
rect 13300 180 13700 200
rect 13300 20 13320 180
rect 13680 20 13700 180
rect 13300 -520 13700 20
rect 13300 -680 13320 -520
rect 13680 -680 13700 -520
rect 13300 -700 13700 -680
rect 11400 -6000 11600 -4400
rect 12800 -6000 13000 -4400
rect 11400 -6200 13000 -6000
rect 9200 -8400 9400 -7000
rect 10600 -8400 10800 -7000
rect 9200 -8600 10800 -8400
rect 7000 -11400 7200 -10000
rect 8400 -11400 8600 -10000
rect 7000 -11600 8600 -11400
rect 14000 -10000 15600 1000
rect 15900 400 18100 500
rect 15900 100 16000 400
rect 18000 100 18100 400
rect 15900 0 18100 100
rect 15900 -500 18100 -400
rect 15900 -800 16000 -500
rect 18000 -800 18100 -500
rect 15900 -900 18100 -800
rect 16200 -1400 17800 -1200
rect 16200 -3000 16400 -1400
rect 17600 -3000 17800 -1400
rect 16200 -7000 17800 -3000
rect 18400 -4400 20000 9600
rect 25400 11000 27000 11200
rect 25400 9600 25600 11000
rect 26800 9600 27000 11000
rect 21000 8000 22600 8200
rect 21000 6600 21200 8000
rect 22400 6600 22600 8000
rect 21000 5600 22600 6600
rect 21000 4000 21200 5600
rect 22400 4000 22600 5600
rect 21000 3800 22600 4000
rect 21000 2600 22600 2800
rect 21000 1000 21200 2600
rect 22400 1000 22600 2600
rect 20300 180 20700 200
rect 20300 20 20320 180
rect 20680 20 20700 180
rect 20300 -520 20700 20
rect 20300 -680 20320 -520
rect 20680 -680 20700 -520
rect 20300 -700 20700 -680
rect 18400 -6000 18600 -4400
rect 19800 -6000 20000 -4400
rect 18400 -6200 20000 -6000
rect 16200 -8400 16400 -7000
rect 17600 -8400 17800 -7000
rect 16200 -8600 17800 -8400
rect 14000 -11400 14200 -10000
rect 15400 -11400 15600 -10000
rect 14000 -11600 15600 -11400
rect 21000 -10000 22600 1000
rect 23200 -1400 24800 -1200
rect 23200 -3000 23400 -1400
rect 24600 -3000 24800 -1400
rect 23200 -7000 24800 -3000
rect 25400 -4400 27000 9600
rect 25400 -6000 25600 -4400
rect 26800 -6000 27000 -4400
rect 25400 -6200 27000 -6000
rect 23200 -8400 23400 -7000
rect 24600 -8400 24800 -7000
rect 23200 -8600 24800 -8400
rect 21000 -11400 21200 -10000
rect 22400 -11400 22600 -10000
rect 21000 -11600 22600 -11400
<< via4 >>
rect 4600 9600 5800 11000
rect 200 6600 1400 8000
rect 2000 300 4000 400
rect 2000 100 4000 300
rect 2000 -700 4000 -500
rect 2000 -800 4000 -700
rect 11600 9600 12800 11000
rect 7200 6600 8400 8000
rect 2400 -8400 3600 -7000
rect 200 -11400 1400 -10000
rect 18600 9600 19800 11000
rect 14200 6600 15400 8000
rect 9400 -8400 10600 -7000
rect 7200 -11400 8400 -10000
rect 16000 300 18000 400
rect 16000 100 18000 300
rect 16000 -700 18000 -500
rect 16000 -800 18000 -700
rect 25600 9600 26800 11000
rect 21200 6600 22400 8000
rect 16400 -8400 17600 -7000
rect 14200 -11400 15400 -10000
rect 23400 -8400 24600 -7000
rect 21200 -11400 22400 -10000
<< metal5 >>
rect 0 8200 2800 11400
rect 24200 11200 27000 11400
rect 4400 11000 27000 11200
rect 4400 9600 4600 11000
rect 5800 9600 11600 11000
rect 12800 9600 18600 11000
rect 19800 9600 25600 11000
rect 26800 9600 27000 11000
rect 4400 9400 27000 9600
rect 0 8000 22600 8200
rect 0 6600 200 8000
rect 1400 6600 7200 8000
rect 8400 6600 14200 8000
rect 15400 6600 21200 8000
rect 22400 6600 22600 8000
rect 0 6400 22600 6600
rect -100 400 27000 500
rect -100 100 2000 400
rect 4000 100 16000 400
rect 18000 100 27000 400
rect -100 0 27000 100
rect -100 -500 27000 -400
rect -100 -800 2000 -500
rect 4000 -800 16000 -500
rect 18000 -800 27000 -500
rect -100 -900 27000 -800
rect 2200 -7000 27000 -6800
rect 2200 -8400 2400 -7000
rect 3600 -8400 9400 -7000
rect 10600 -8400 16400 -7000
rect 17600 -8400 23400 -7000
rect 24600 -8400 27000 -7000
rect 2200 -8600 27000 -8400
rect 0 -10000 22600 -9800
rect 0 -11400 200 -10000
rect 1400 -11400 7200 -10000
rect 8400 -11400 14200 -10000
rect 15400 -11400 21200 -10000
rect 22400 -11400 22600 -10000
rect 0 -11600 22600 -11400
rect 0 -11800 2800 -11600
rect 24200 -11800 27000 -8600
<< labels >>
rlabel metal5 24200 11200 27000 11400 1 SD1R
rlabel metal5 0 11200 2800 11400 1 SD1L
rlabel metal5 0 -11800 2800 -11600 1 SD2L
rlabel metal5 24200 -11800 27000 -11600 1 SD2R
rlabel metal5 -100 0 0 500 1 GL
rlabel metal5 -100 -900 0 -400 1 GR
rlabel metal2 14030 5720 14100 5780 1 SUB
rlabel metal2 7030 5720 7100 5780 1 SUB
rlabel metal2 21030 5720 21100 5780 1 SUB
rlabel metal2 7030 -6780 7100 -6720 1 SUB
rlabel metal2 14030 -6780 14100 -6720 1 SUB
rlabel metal2 21030 -6780 21100 -6720 1 SUB
rlabel metal2 12600 -12300 13600 -12100 1 SUB
<< end >>
