magic
tech sky130B
timestamp 1659057364
<< metal4 >>
rect 2400 2250 3200 2300
rect 2400 1650 2450 2250
rect 3150 1650 3200 2250
rect 2400 -400 3200 1650
<< via4 >>
rect 2450 1650 3150 2250
<< metal5 >>
rect 0 9500 10000 10000
rect 0 0 500 9500
rect 800 8700 9200 9200
rect 800 500 1300 8700
rect 1600 7900 8400 8400
rect 1600 1300 2100 7900
rect 2400 2250 3200 2300
rect 2400 1650 2450 2250
rect 3150 2200 3250 2250
rect 3150 2150 3300 2200
rect 3150 2100 3350 2150
rect 7900 2100 8400 7900
rect 3150 1650 8400 2100
rect 2400 1600 8400 1650
rect 8700 1300 9200 8700
rect 1600 800 9200 1300
rect 9500 500 10000 9500
rect 800 0 10000 500
<< labels >>
rlabel metal4 2400 -400 3200 -100 1 B
rlabel metal5 0 0 500 250 1 A
<< end >>
