magic
tech sky130B
timestamp 1662008789
<< metal3 >>
rect 8097 81150 10597 82000
rect 34097 81150 36597 82000
rect 60097 81150 62597 82000
rect 82797 81150 85297 82000
rect 85447 81150 86547 82000
rect 86697 81150 87797 82000
rect 87947 81150 90447 82000
rect 108647 81150 111147 82000
rect 111297 81150 112397 82000
rect 112547 81150 113647 82000
rect 113797 81150 116297 82000
rect 159497 81150 161997 82000
rect 162147 81150 163247 82000
rect 163397 81150 164497 82000
rect 164647 81150 167147 82000
rect 206697 81150 209197 82000
rect 232697 81150 235197 82000
rect 255297 81170 257697 82000
rect 260297 81170 262697 82000
rect 283297 81150 285797 82000
rect 0 70121 850 72621
rect 291150 68992 292000 71492
rect 0 51921 830 54321
rect 291170 49892 292000 52292
rect 0 46921 830 49321
rect 291170 44892 292000 47292
rect 291760 24736 292400 24792
rect 291760 24145 292400 24201
rect 291760 23554 292400 23610
rect 291760 22963 292400 23019
rect 291760 22372 292400 22428
rect 291760 21781 292400 21837
rect 0 9721 830 12121
rect 0 4721 830 7121
rect 291170 5281 292000 7681
rect 291170 281 292000 2681
rect 10000 0 10056 200
rect 13100 0 13156 200
rect 16200 0 16256 200
rect 19300 0 19356 200
rect 22400 0 22456 200
rect 25500 0 25556 200
rect 28600 0 28656 200
rect 31700 0 31756 200
rect 34800 0 34856 200
rect 37900 0 37956 200
rect 41000 0 41056 200
rect 44100 0 44156 200
rect 47200 0 47256 200
rect 50300 0 50356 200
rect 53400 0 53456 200
rect 56500 0 56556 200
rect 59600 0 59656 200
rect 62700 0 62756 200
rect 65800 0 65856 200
rect 68900 0 68956 200
rect 72000 0 72056 200
rect 75100 0 75156 200
rect 78200 0 78256 200
rect 81300 0 81356 200
rect 84400 0 84456 200
rect 87500 0 87556 200
rect 90600 0 90656 200
rect 93700 0 93756 200
rect 96800 0 96856 200
rect 99900 0 99956 200
rect 103000 0 103056 200
rect 106100 0 106156 200
rect 109200 0 109256 200
rect 112300 0 112356 200
rect 115400 0 115456 200
rect 118500 0 118556 200
rect 121600 0 121656 200
rect 124700 0 124756 200
rect 127800 0 127856 200
rect 130900 0 130956 200
rect 134000 0 134056 200
rect 137100 0 137156 200
rect 140200 0 140256 200
rect 143300 0 143356 200
rect 146400 0 146456 200
rect 149500 0 149556 200
rect 152600 0 152656 200
rect 155700 0 155756 200
rect 158800 0 158856 200
rect 161900 0 161956 200
rect 165000 0 165056 200
rect 168100 0 168156 200
rect 171200 0 171256 200
rect 174300 0 174356 200
rect 177400 0 177456 200
rect 180500 0 180556 200
rect 183600 0 183656 200
rect 186700 0 186756 200
rect 189800 0 189856 200
rect 192900 0 192956 200
<< metal4 >>
rect 3049 0 6899 400
rect 7229 0 11079 400
rect 282049 0 285899 400
rect 286229 0 290079 400
<< labels >>
rlabel metal3 s 10000 0 10056 200 0 analog_la_out[0]
port 1 nsew
rlabel metal3 s 13100 0 13156 200 0 analog_la_out[1]
port 2 nsew
rlabel metal3 s 16200 0 16256 200 0 analog_la_out[2]
port 3 nsew
rlabel metal3 s 19300 0 19356 200 0 analog_la_out[3]
port 4 nsew
rlabel metal3 s 22400 0 22456 200 0 analog_la_out[4]
port 5 nsew
rlabel metal3 s 25500 0 25556 200 0 analog_la_out[5]
port 6 nsew
rlabel metal3 s 28600 0 28656 200 0 analog_la_out[6]
port 7 nsew
rlabel metal3 s 31700 0 31756 200 0 analog_la_out[7]
port 8 nsew
rlabel metal3 s 34800 0 34856 200 0 analog_la_out[8]
port 9 nsew
rlabel metal3 s 37900 0 37956 200 0 analog_la_out[9]
port 10 nsew
rlabel metal3 s 41000 0 41056 200 0 analog_la_out[10]
port 11 nsew
rlabel metal3 s 44100 0 44156 200 0 analog_la_out[11]
port 12 nsew
rlabel metal3 s 47200 0 47256 200 0 analog_la_out[12]
port 13 nsew
rlabel metal3 s 50300 0 50356 200 0 analog_la_out[13]
port 14 nsew
rlabel metal3 s 53400 0 53456 200 0 analog_la_out[14]
port 15 nsew
rlabel metal3 s 56500 0 56556 200 0 analog_la_out[15]
port 16 nsew
rlabel metal3 s 59600 0 59656 200 0 analog_la_out[16]
port 17 nsew
rlabel metal3 s 62700 0 62756 200 0 analog_la_out[17]
port 18 nsew
rlabel metal3 s 65800 0 65856 200 0 analog_la_out[18]
port 19 nsew
rlabel metal3 s 68900 0 68956 200 0 analog_la_out[19]
port 20 nsew
rlabel metal3 s 72000 0 72056 200 0 analog_la_out[20]
port 21 nsew
rlabel metal3 s 75100 0 75156 200 0 analog_la_out[21]
port 22 nsew
rlabel metal3 s 78200 0 78256 200 0 analog_la_out[22]
port 23 nsew
rlabel metal3 s 81300 0 81356 200 0 analog_la_out[23]
port 24 nsew
rlabel metal3 s 84400 0 84456 200 0 analog_la_out[24]
port 25 nsew
rlabel metal3 s 87500 0 87556 200 0 analog_la_out[25]
port 26 nsew
rlabel metal3 s 90600 0 90656 200 0 analog_la_out[26]
port 27 nsew
rlabel metal3 s 93700 0 93756 200 0 analog_la_out[27]
port 28 nsew
rlabel metal3 s 96800 0 96856 200 0 analog_la_out[28]
port 29 nsew
rlabel metal3 s 99900 0 99956 200 0 analog_la_out[29]
port 30 nsew
rlabel metal3 s 103000 0 103056 200 0 analog_la_in[0]
port 31 nsew
rlabel metal3 s 106100 0 106156 200 0 analog_la_in[1]
port 32 nsew
rlabel metal3 s 109200 0 109256 200 0 analog_la_in[2]
port 33 nsew
rlabel metal3 s 112300 0 112356 200 0 analog_la_in[3]
port 34 nsew
rlabel metal3 s 115400 0 115456 200 0 analog_la_in[4]
port 35 nsew
rlabel metal3 s 118500 0 118556 200 0 analog_la_in[5]
port 36 nsew
rlabel metal3 s 121600 0 121656 200 0 analog_la_in[6]
port 37 nsew
rlabel metal3 s 124700 0 124756 200 0 analog_la_in[7]
port 38 nsew
rlabel metal3 s 127800 0 127856 200 0 analog_la_in[8]
port 39 nsew
rlabel metal3 s 130900 0 130956 200 0 analog_la_in[9]
port 40 nsew
rlabel metal3 s 134000 0 134056 200 0 analog_la_in[10]
port 41 nsew
rlabel metal3 s 137100 0 137156 200 0 analog_la_in[11]
port 42 nsew
rlabel metal3 s 140200 0 140256 200 0 analog_la_in[12]
port 43 nsew
rlabel metal3 s 143300 0 143356 200 0 analog_la_in[13]
port 44 nsew
rlabel metal3 s 146400 0 146456 200 0 analog_la_in[14]
port 45 nsew
rlabel metal3 s 149500 0 149556 200 0 analog_la_in[15]
port 46 nsew
rlabel metal3 s 152600 0 152656 200 0 analog_la_in[16]
port 47 nsew
rlabel metal3 s 155700 0 155756 200 0 analog_la_in[17]
port 48 nsew
rlabel metal3 s 158800 0 158856 200 0 analog_la_in[18]
port 49 nsew
rlabel metal3 s 161900 0 161956 200 0 analog_la_in[19]
port 50 nsew
rlabel metal3 s 165000 0 165056 200 0 analog_la_in[20]
port 51 nsew
rlabel metal3 s 168100 0 168156 200 0 analog_la_in[21]
port 52 nsew
rlabel metal3 s 171200 0 171256 200 0 analog_la_in[22]
port 53 nsew
rlabel metal3 s 174300 0 174356 200 0 analog_la_in[23]
port 54 nsew
rlabel metal3 s 177400 0 177456 200 0 analog_la_in[24]
port 55 nsew
rlabel metal3 s 180500 0 180556 200 0 analog_la_in[25]
port 56 nsew
rlabel metal3 s 183600 0 183656 200 0 analog_la_in[26]
port 57 nsew
rlabel metal3 s 186700 0 186756 200 0 analog_la_in[27]
port 58 nsew
rlabel metal3 s 189800 0 189856 200 0 analog_la_in[28]
port 59 nsew
rlabel metal3 s 192900 0 192956 200 0 analog_la_in[29]
port 60 nsew
rlabel metal3 s 291760 21781 292400 21837 0 gpio_analog[6]
port 61 nsew
rlabel metal3 s 291760 22372 292400 22428 0 gpio_noesd[6]
port 62 nsew
rlabel metal3 s 291150 68992 292000 71492 0 io_analog[0]
port 63 nsew
rlabel metal3 s 0 70121 850 72621 0 io_analog[10]
port 64 nsew
rlabel metal3 s 283297 81150 285797 82000 0 io_analog[1]
port 65 nsew
rlabel metal3 s 232697 81150 235197 82000 0 io_analog[2]
port 66 nsew
rlabel metal3 s 206697 81150 209197 82000 0 io_analog[3]
port 67 nsew
rlabel metal3 s 159497 81150 161997 82000 0 io_analog[4]
port 68 nsew
rlabel metal3 s 108647 81150 111147 82000 0 io_analog[5]
port 69 nsew
rlabel metal3 s 82797 81150 85297 82000 0 io_analog[6]
port 70 nsew
rlabel metal3 s 60097 81150 62597 82000 0 io_analog[7]
port 71 nsew
rlabel metal3 s 34097 81150 36597 82000 0 io_analog[8]
port 72 nsew
rlabel metal3 s 8097 81150 10597 82000 0 io_analog[9]
port 73 nsew
rlabel metal3 s 163397 81150 164497 82000 0 io_clamp_high[0]
port 74 nsew
rlabel metal3 s 112547 81150 113647 82000 0 io_clamp_high[1]
port 75 nsew
rlabel metal3 s 86697 81150 87797 82000 0 io_clamp_high[2]
port 76 nsew
rlabel metal3 s 162147 81150 163247 82000 0 io_clamp_low[0]
port 77 nsew
rlabel metal3 s 111297 81150 112397 82000 0 io_clamp_low[1]
port 78 nsew
rlabel metal3 s 85447 81150 86547 82000 0 io_clamp_low[2]
port 79 nsew
rlabel metal3 s 291760 23554 292400 23610 0 io_in[13]
port 80 nsew
rlabel metal3 s 291760 22963 292400 23019 0 io_in_3v3[13]
port 81 nsew
rlabel metal3 s 291760 24736 292400 24792 0 io_oeb[13]
port 82 nsew
rlabel metal3 s 291760 24145 292400 24201 0 io_out[13]
port 83 nsew
rlabel metal3 s 291170 44892 292000 47292 0 vccd1
port 84 nsew
rlabel metal3 s 0 46921 830 49321 0 vccd2
port 85 nsew
rlabel metal3 s 291170 5281 292000 7681 0 vdda1
port 86 nsew
rlabel metal3 s 255297 81170 257697 82000 0 vssa1
port 87 nsew
rlabel metal3 s 0 4721 830 7121 0 vssa2
port 88 nsew
rlabel metal4 s 282049 0 285899 400 0 vdda1
port 86 nsew
rlabel metal4 s 286229 0 290079 400 0 vssa1
port 87 nsew
rlabel metal4 s 3049 0 6899 400 0 vdda2
port 89 nsew
rlabel metal4 s 7229 0 11079 400 0 vssd2
port 90 nsew
<< properties >>
string FIXED_BBOX 0 0 292000 82000
string path 1929.280 0.000 1929.280 2.000 
<< end >>
