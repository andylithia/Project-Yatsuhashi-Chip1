magic
tech sky130A
timestamp 1664680375
<< metal4 >>
rect -6700 25850 -5950 25900
rect -6700 25250 -6650 25850
rect -6000 25250 -5950 25850
rect -6700 24250 -5950 25250
rect -2600 25850 -1850 25900
rect -2600 25250 -2550 25850
rect -1900 25250 -1850 25850
rect -4800 24950 -4050 25000
rect -4800 24350 -4750 24950
rect -4100 24350 -4050 24950
rect -4800 24200 -4050 24350
rect -3550 24950 -2800 25000
rect -3550 24350 -3500 24950
rect -2850 24350 -2800 24950
rect -3550 24200 -2800 24350
rect -2600 24300 -1850 25250
rect -400 25850 350 25900
rect -400 25250 -350 25850
rect 300 25250 350 25850
rect -400 24300 350 25250
rect 3700 25850 4450 25900
rect 3700 25250 3750 25850
rect 4400 25250 4450 25850
rect 1500 24950 2250 25000
rect 1500 24350 1550 24950
rect 2200 24350 2250 24950
rect 1500 24200 2250 24350
rect 2750 24950 3500 25000
rect 2750 24350 2800 24950
rect 3450 24350 3500 24950
rect 2750 24200 3500 24350
rect 3700 24250 4450 25250
rect -6700 18500 -5950 18550
rect -6700 17950 -6650 18500
rect -6000 17950 -5950 18500
rect -6700 17000 -5950 17950
rect -5750 17600 -5000 18600
rect -3550 18500 -2800 18950
rect -3550 17950 -3500 18500
rect -2850 17950 -2800 18500
rect -3550 17900 -2800 17950
rect -2600 18500 -1850 18550
rect -2600 17950 -2550 18500
rect -1900 17950 -1850 18500
rect -5750 17050 -5700 17600
rect -5050 17050 -5000 17600
rect -5750 17000 -5000 17050
rect -4800 17600 -4050 17650
rect -4800 17050 -4750 17600
rect -4100 17050 -4050 17600
rect -4800 17000 -4050 17050
rect -3550 17600 -2800 17650
rect -3550 17050 -3500 17600
rect -2850 17050 -2800 17600
rect -3550 17000 -2800 17050
rect -2600 17000 -1850 17950
rect -1650 17600 -900 18600
rect -1650 17050 -1600 17600
rect -950 17050 -900 17600
rect -1650 17000 -900 17050
rect -400 18500 350 18550
rect -400 17950 -350 18500
rect 300 17950 350 18500
rect 2750 18500 3500 18600
rect -400 17000 350 17950
rect 550 17600 1300 18400
rect 2750 17950 2800 18500
rect 3450 17950 3500 18500
rect 2750 17900 3500 17950
rect 3700 18500 4450 18550
rect 3700 17950 3750 18500
rect 4400 17950 4450 18500
rect 550 17050 600 17600
rect 1250 17050 1300 17600
rect 550 17000 1300 17050
rect 1500 17600 2250 17650
rect 1500 17050 1550 17600
rect 2200 17050 2250 17600
rect 1500 16650 2250 17050
rect 2750 17600 3500 17650
rect 2750 17050 2800 17600
rect 3450 17050 3500 17600
rect 2750 16650 3500 17050
rect 3700 16650 4450 17950
rect 4650 17600 5400 18550
rect 4650 17050 4700 17600
rect 5350 17050 5400 17600
rect 4650 17000 5400 17050
rect -6700 10850 -5950 10900
rect -6700 10300 -6650 10850
rect -6000 10300 -5950 10850
rect -6700 9350 -5950 10300
rect -5750 9950 -5000 10950
rect -3550 10850 -2800 11300
rect -3550 10300 -3500 10850
rect -2850 10300 -2800 10850
rect -3550 10250 -2800 10300
rect -2600 10850 -1850 10900
rect -2600 10300 -2550 10850
rect -1900 10300 -1850 10850
rect -5750 9400 -5700 9950
rect -5050 9400 -5000 9950
rect -5750 9350 -5000 9400
rect -4800 9950 -4050 10000
rect -4800 9400 -4750 9950
rect -4100 9400 -4050 9950
rect -4800 9350 -4050 9400
rect -3550 9950 -2800 10000
rect -3550 9400 -3500 9950
rect -2850 9400 -2800 9950
rect -3550 9350 -2800 9400
rect -2600 9350 -1850 10300
rect -1650 9950 -900 10950
rect -1650 9400 -1600 9950
rect -950 9400 -900 9950
rect -1650 9350 -900 9400
rect -400 10850 350 10900
rect -400 10300 -350 10850
rect 300 10300 350 10850
rect 2750 10850 3500 10950
rect -400 9350 350 10300
rect 550 9950 1300 10750
rect 2750 10300 2800 10850
rect 3450 10300 3500 10850
rect 2750 10250 3500 10300
rect 3700 10850 4450 10900
rect 3700 10300 3750 10850
rect 4400 10300 4450 10850
rect 550 9400 600 9950
rect 1250 9400 1300 9950
rect 550 9350 1300 9400
rect 1500 9950 2250 10000
rect 1500 9400 1550 9950
rect 2200 9400 2250 9950
rect 1500 9000 2250 9400
rect 2750 9950 3500 10000
rect 2750 9400 2800 9950
rect 3450 9400 3500 9950
rect 2750 9000 3500 9400
rect 3700 9000 4450 10300
rect 4650 9950 5400 10900
rect 4650 9400 4700 9950
rect 5350 9400 5400 9950
rect 4650 9350 5400 9400
rect -5750 2700 -5000 3650
rect -5750 2100 -5700 2700
rect -5050 2100 -5000 2700
rect -5750 2050 -5000 2100
rect -1650 2700 -900 3650
rect -1650 2100 -1600 2700
rect -950 2100 -900 2700
rect -1650 2050 -900 2100
rect 550 2700 1300 3650
rect 550 2100 600 2700
rect 1250 2100 1300 2700
rect 550 2050 1300 2100
rect 4650 2700 5400 3650
rect 4650 2100 4700 2700
rect 5350 2100 5400 2700
rect 4650 2050 5400 2100
<< via4 >>
rect -6650 25250 -6000 25850
rect -2550 25250 -1900 25850
rect -4750 24350 -4100 24950
rect -3500 24350 -2850 24950
rect -350 25250 300 25850
rect 3750 25250 4400 25850
rect 1550 24350 2200 24950
rect 2800 24350 3450 24950
rect -6650 17950 -6000 18500
rect -3500 17950 -2850 18500
rect -2550 17950 -1900 18500
rect -5700 17050 -5050 17600
rect -4750 17050 -4100 17600
rect -3500 17050 -2850 17600
rect -1600 17050 -950 17600
rect -350 17950 300 18500
rect 2800 17950 3450 18500
rect 3750 17950 4400 18500
rect 600 17050 1250 17600
rect 1550 17050 2200 17600
rect 2800 17050 3450 17600
rect 4700 17050 5350 17600
rect -6650 10300 -6000 10850
rect -3500 10300 -2850 10850
rect -2550 10300 -1900 10850
rect -5700 9400 -5050 9950
rect -4750 9400 -4100 9950
rect -3500 9400 -2850 9950
rect -1600 9400 -950 9950
rect -350 10300 300 10850
rect 2800 10300 3450 10850
rect 3750 10300 4400 10850
rect 600 9400 1250 9950
rect 1550 9400 2200 9950
rect 2800 9400 3450 9950
rect 4700 9400 5350 9950
rect -6650 3000 -6000 3600
rect -3500 3000 -2850 3600
rect -5700 2100 -5050 2700
rect -350 3000 300 3600
rect -1600 2100 -950 2700
rect 2800 3000 3450 3600
rect 600 2100 1250 2700
rect 4700 2100 5350 2700
<< metal5 >>
rect -6700 25900 -5950 26100
rect -6700 25850 4450 25900
rect -6700 25250 -6650 25850
rect -6000 25250 -2550 25850
rect -1900 25250 -350 25850
rect 300 25250 3750 25850
rect 4400 25250 4450 25850
rect -6700 25200 4450 25250
rect 4650 25000 5400 26100
rect -4800 24950 5400 25000
rect -4800 24350 -4750 24950
rect -4100 24350 -3500 24950
rect -2850 24350 1550 24950
rect 2200 24350 2800 24950
rect 3450 24350 5400 24950
rect -4800 24300 5400 24350
rect -6750 21700 -6700 21950
rect -6750 21250 -6700 21500
rect -6700 18500 5400 18550
rect -6700 17950 -6650 18500
rect -6000 17950 -3500 18500
rect -2850 17950 -2550 18500
rect -1900 17950 -350 18500
rect 300 17950 2800 18500
rect 3450 17950 3750 18500
rect 4400 17950 5400 18500
rect -6700 17900 5400 17950
rect -6700 17600 5400 17650
rect -6700 17050 -5700 17600
rect -5050 17050 -4750 17600
rect -4100 17050 -3500 17600
rect -2850 17050 -1600 17600
rect -950 17050 600 17600
rect 1250 17050 1550 17600
rect 2200 17050 2800 17600
rect 3450 17050 4700 17600
rect 5350 17050 5400 17600
rect -6700 17000 5400 17050
rect -6750 14050 -6700 14300
rect -6750 13600 -6700 13850
rect -6700 10850 5400 10900
rect -6700 10300 -6650 10850
rect -6000 10300 -3500 10850
rect -2850 10300 -2550 10850
rect -1900 10300 -350 10850
rect 300 10300 2800 10850
rect 3450 10300 3750 10850
rect 4400 10300 5400 10850
rect -6700 10250 5400 10300
rect -6700 9950 5400 10000
rect -6700 9400 -5700 9950
rect -5050 9400 -4750 9950
rect -4100 9400 -3500 9950
rect -2850 9400 -1600 9950
rect -950 9400 600 9950
rect 1250 9400 1550 9950
rect 2200 9400 2800 9950
rect 3450 9400 4700 9950
rect 5350 9400 5400 9950
rect -6700 9350 5400 9400
rect -6750 6400 -6700 6650
rect -6750 5950 -6700 6200
rect -6700 3600 3500 3650
rect -6700 3000 -6650 3600
rect -6000 3000 -3500 3600
rect -2850 3000 -350 3600
rect 300 3000 2800 3600
rect 3450 3000 3500 3600
rect -6700 2950 3500 3000
rect -6700 1850 -5950 2950
rect -5750 2700 5400 2750
rect -5750 2100 -5700 2700
rect -5050 2100 -1600 2700
rect -950 2100 600 2700
rect 1250 2100 4700 2700
rect 5350 2100 5400 2700
rect -5750 2050 5400 2100
rect 4650 1850 5400 2050
<< comment >>
rect -7250 24900 -7200 24950
rect -7300 24800 -7250 24900
rect -7200 24800 -7150 24850
rect -7300 24750 -7150 24800
rect -7200 24700 -7150 24750
rect -7350 17550 -7200 17600
rect -7250 17500 -7200 17550
rect -7300 17450 -7200 17500
rect -7250 17400 -7200 17450
rect -7350 17350 -7200 17400
rect -7300 9650 -7150 9700
rect -7200 9600 -7150 9650
rect -7250 9550 -7150 9600
rect -7300 9500 -7250 9550
rect -7300 9450 -7150 9500
rect -7150 2250 -7100 2300
rect -7200 2200 -7100 2250
rect -7150 2100 -7100 2200
rect -7200 2050 -7050 2100
use NMOS_30_0p5_30_diff4x_2s  NMOS_30_0p5_30_diff4x_2s_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/CLASSE
timestamp 1664504783
transform 1 0 -7400 0 1 6400
box 650 -3650 12800 3500
use NMOS_30_0p5_30_diff4x_2s  NMOS_30_0p5_30_diff4x_2s_1
timestamp 1664504783
transform 1 0 -7400 0 1 14050
box 650 -3650 12800 3500
use NMOS_30_0p5_30_diff4x_2s  NMOS_30_0p5_30_diff4x_2s_2
timestamp 1664504783
transform 1 0 -7400 0 1 21700
box 650 -3650 12800 3500
<< labels >>
rlabel metal5 -6700 1850 -5950 2050 1 SD1L
rlabel metal5 4650 1850 5400 2050 1 SD1R
rlabel metal5 -6700 25900 -5950 26100 1 SD4L
rlabel metal5 4650 25900 5400 26100 1 SD4R
rlabel metal5 -6750 6400 -6700 6650 1 G12L
rlabel metal5 -6750 5950 -6700 6200 1 G12R
rlabel metal5 -6750 13600 -6700 13850 1 G23R
rlabel metal5 -6750 14050 -6700 14300 1 G23L
rlabel metal5 -6750 21250 -6700 21500 1 G34R
rlabel metal5 -6750 21700 -6700 21950 1 G34L
rlabel metal4 -6700 17850 -6550 18550 1 SD3L
rlabel space -6700 16950 -6550 17650 1 SD3R
rlabel metal4 -6700 10200 -6550 10900 1 SD3L
rlabel space -6700 9300 -6550 10000 1 SD3R
<< end >>
