magic
tech sky130B
timestamp 0
<< end >>
