magic
tech sky130B
timestamp 1664070670
<< metal2 >>
rect 6300 5850 6800 5950
rect 6300 3250 6500 5850
rect 6600 3250 6800 5850
rect 2550 3150 3550 3250
rect 6050 3150 7050 3250
rect 9550 3150 10550 3250
rect 2650 2900 2850 3150
rect 2950 2900 3150 3150
rect 3250 2900 3450 3150
rect 6150 2900 6350 3150
rect 6450 2900 6650 3150
rect 6750 2900 6950 3150
rect 9650 2900 9850 3150
rect 9950 2900 10150 3150
rect 10250 2900 10450 3150
rect 2550 2800 3550 2900
rect 6050 2800 7050 2900
rect 9550 2800 10550 2900
rect 6300 100 6500 2800
rect 6600 100 6800 2800
rect 2550 0 3550 100
rect 6050 0 7050 100
rect 9550 0 10550 100
rect 2650 -250 2850 0
rect 2950 -250 3150 0
rect 3250 -250 3450 0
rect 6150 -250 6350 0
rect 6450 -250 6650 0
rect 6750 -250 6950 0
rect 9650 -250 9850 0
rect 9950 -250 10150 0
rect 10250 -250 10450 0
rect 2550 -350 3550 -250
rect 6050 -350 7050 -250
rect 9550 -350 10550 -250
rect 6300 -3000 6500 -350
rect 6600 -3000 6800 -350
rect 2550 -3100 3550 -3000
rect 6050 -3100 7050 -3000
rect 9550 -3100 10550 -3000
rect 2650 -3350 2850 -3100
rect 2950 -3350 3150 -3100
rect 3250 -3350 3450 -3100
rect 6150 -3350 6350 -3100
rect 6450 -3350 6650 -3100
rect 6750 -3350 6950 -3100
rect 9650 -3350 9850 -3100
rect 9950 -3350 10150 -3100
rect 10250 -3350 10450 -3100
rect 2550 -3450 3550 -3350
rect 6050 -3450 7050 -3350
rect 9550 -3450 10550 -3350
rect 6300 -6050 6500 -3450
rect 6600 -6050 6800 -3450
rect 6300 -6150 6800 -6050
<< metal3 >>
rect 950 150 2050 200
rect 7950 150 9050 200
rect 850 50 1000 150
rect 2000 50 2150 150
rect 4350 100 5650 150
rect 850 -50 2150 50
rect 2250 90 3350 100
rect 2250 10 3160 90
rect 3340 10 3350 90
rect 2250 0 3350 10
rect 3450 90 6850 100
rect 3450 10 6660 90
rect 6840 10 6850 90
rect 3450 0 6850 10
rect 6950 10 7110 100
rect 7850 50 8000 150
rect 9000 100 9150 150
rect 9000 90 10350 100
rect 9000 50 10160 90
rect 7850 10 10160 50
rect 10340 10 10350 90
rect 6950 0 7100 10
rect 7850 0 10350 10
rect 3450 -100 3550 0
rect 4350 -50 5650 0
rect 6950 -50 7050 0
rect 7850 -50 9150 0
rect 10450 -50 10600 100
rect 11350 -50 12650 150
rect 2950 -200 3550 -100
rect 6450 -150 7050 -50
rect 9950 -150 10600 -50
rect 850 -250 2150 -200
rect 2950 -250 3050 -200
rect 850 -350 1000 -250
rect 2000 -350 3050 -250
rect 3150 -260 3700 -250
rect 3150 -340 3160 -260
rect 3340 -340 3700 -260
rect 3150 -350 3700 -340
rect 850 -400 2150 -350
rect 4350 -400 5650 -200
rect 6450 -250 6550 -150
rect 7850 -250 9150 -200
rect 9950 -250 10050 -150
rect 6040 -350 6550 -250
rect 6650 -260 7570 -250
rect 6650 -340 6660 -260
rect 6840 -340 7570 -260
rect 6650 -350 7570 -340
rect 7850 -350 8000 -250
rect 9000 -350 9150 -250
rect 9300 -350 10050 -250
rect 10150 -260 10650 -250
rect 10150 -340 10160 -260
rect 10340 -340 10650 -260
rect 10150 -350 10650 -340
rect 7850 -400 9150 -350
rect 11350 -400 12650 -200
rect 100 -2200 3100 -2100
rect 100 -3000 2300 -2200
rect 2900 -3000 3100 -2200
rect 100 -3100 3100 -3000
rect 3600 -2200 6600 -2100
rect 3600 -3000 5800 -2200
rect 6400 -3000 6600 -2200
rect 3600 -3100 6600 -3000
rect 7100 -2200 10100 -2100
rect 7100 -3000 9300 -2200
rect 9900 -3000 10100 -2200
rect 7100 -3100 10100 -3000
rect 10600 -2200 13600 -2100
rect 10600 -3000 12800 -2200
rect 13400 -3000 13600 -2200
rect 10600 -3100 13600 -3000
<< via3 >>
rect 100 2000 700 2800
rect 3600 2000 4200 2800
rect 7100 2000 7700 2800
rect 10600 2000 11200 2800
rect 100 500 700 1300
rect 3600 500 4200 1300
rect 7100 500 7700 1300
rect 10600 500 11200 1300
rect 1000 50 2000 150
rect 3160 10 3340 90
rect 6660 10 6840 90
rect 8000 50 9000 150
rect 10160 10 10340 90
rect 1000 -350 2000 -250
rect 3160 -340 3340 -260
rect 6660 -340 6840 -260
rect 8000 -350 9000 -250
rect 10160 -340 10340 -260
rect 1200 -1500 1800 -700
rect 4700 -1500 5300 -700
rect 8200 -1500 8800 -700
rect 11700 -1500 12300 -700
rect 2300 -3000 2900 -2200
rect 5800 -3000 6400 -2200
rect 9300 -3000 9900 -2200
rect 12800 -3000 13400 -2200
<< metal4 >>
rect 2200 5500 3000 5600
rect 2200 4800 2300 5500
rect 2900 4800 3000 5500
rect 0 4000 800 4100
rect 0 3300 100 4000
rect 700 3300 800 4000
rect 0 2800 800 3300
rect 0 2000 100 2800
rect 700 2000 800 2800
rect 0 1900 800 2000
rect 0 1300 800 1400
rect 0 500 100 1300
rect 700 500 800 1300
rect 0 -5000 800 500
rect 950 200 2050 250
rect 950 50 1000 200
rect 2000 50 2050 200
rect 950 0 2050 50
rect 950 -250 2050 -200
rect 950 -400 1000 -250
rect 2000 -400 2050 -250
rect 950 -450 2050 -400
rect 1100 -700 1900 -600
rect 1100 -1500 1200 -700
rect 1800 -1500 1900 -700
rect 1100 -3500 1900 -1500
rect 2200 -2200 3000 4800
rect 5700 5500 6500 5600
rect 5700 4800 5800 5500
rect 6400 4800 6500 5500
rect 3500 4000 4300 4100
rect 3500 3300 3600 4000
rect 4200 3300 4300 4000
rect 3500 2800 4300 3300
rect 3500 2000 3600 2800
rect 4200 2000 4300 2800
rect 3500 1900 4300 2000
rect 3500 1300 4300 1400
rect 3500 500 3600 1300
rect 4200 500 4300 1300
rect 3150 90 3350 100
rect 3150 10 3160 90
rect 3340 10 3350 90
rect 3150 -260 3350 10
rect 3150 -340 3160 -260
rect 3340 -340 3350 -260
rect 3150 -350 3350 -340
rect 2200 -3000 2300 -2200
rect 2900 -3000 3000 -2200
rect 2200 -3100 3000 -3000
rect 1100 -4200 1200 -3500
rect 1800 -4200 1900 -3500
rect 1100 -4300 1900 -4200
rect 0 -5700 100 -5000
rect 700 -5700 800 -5000
rect 0 -5800 800 -5700
rect 3500 -5000 4300 500
rect 4600 -700 5400 -600
rect 4600 -1500 4700 -700
rect 5300 -1500 5400 -700
rect 4600 -3500 5400 -1500
rect 5700 -2200 6500 4800
rect 9200 5500 10000 5600
rect 9200 4800 9300 5500
rect 9900 4800 10000 5500
rect 7000 4000 7800 4100
rect 7000 3300 7100 4000
rect 7700 3300 7800 4000
rect 7000 2800 7800 3300
rect 7000 2000 7100 2800
rect 7700 2000 7800 2800
rect 7000 1900 7800 2000
rect 7000 1300 7800 1400
rect 7000 500 7100 1300
rect 7700 500 7800 1300
rect 6650 90 6850 100
rect 6650 10 6660 90
rect 6840 10 6850 90
rect 6650 -260 6850 10
rect 6650 -340 6660 -260
rect 6840 -340 6850 -260
rect 6650 -350 6850 -340
rect 5700 -3000 5800 -2200
rect 6400 -3000 6500 -2200
rect 5700 -3100 6500 -3000
rect 4600 -4200 4700 -3500
rect 5300 -4200 5400 -3500
rect 4600 -4300 5400 -4200
rect 3500 -5700 3600 -5000
rect 4200 -5700 4300 -5000
rect 3500 -5800 4300 -5700
rect 7000 -5000 7800 500
rect 7950 200 9050 250
rect 7950 50 8000 200
rect 9000 50 9050 200
rect 7950 0 9050 50
rect 7950 -250 9050 -200
rect 7950 -400 8000 -250
rect 9000 -400 9050 -250
rect 7950 -450 9050 -400
rect 8100 -700 8900 -600
rect 8100 -1500 8200 -700
rect 8800 -1500 8900 -700
rect 8100 -3500 8900 -1500
rect 9200 -2200 10000 4800
rect 12700 5500 13500 5600
rect 12700 4800 12800 5500
rect 13400 4800 13500 5500
rect 10500 4000 11300 4100
rect 10500 3300 10600 4000
rect 11200 3300 11300 4000
rect 10500 2800 11300 3300
rect 10500 2000 10600 2800
rect 11200 2000 11300 2800
rect 10500 1900 11300 2000
rect 10500 1300 11300 1400
rect 10500 500 10600 1300
rect 11200 500 11300 1300
rect 10150 90 10350 100
rect 10150 10 10160 90
rect 10340 10 10350 90
rect 10150 -260 10350 10
rect 10150 -340 10160 -260
rect 10340 -340 10350 -260
rect 10150 -350 10350 -340
rect 9200 -3000 9300 -2200
rect 9900 -3000 10000 -2200
rect 9200 -3100 10000 -3000
rect 8100 -4200 8200 -3500
rect 8800 -4200 8900 -3500
rect 8100 -4300 8900 -4200
rect 7000 -5700 7100 -5000
rect 7700 -5700 7800 -5000
rect 7000 -5800 7800 -5700
rect 10500 -5000 11300 500
rect 11600 -700 12400 -600
rect 11600 -1500 11700 -700
rect 12300 -1500 12400 -700
rect 11600 -3500 12400 -1500
rect 12700 -2200 13500 4800
rect 12700 -3000 12800 -2200
rect 13400 -3000 13500 -2200
rect 12700 -3100 13500 -3000
rect 11600 -4200 11700 -3500
rect 12300 -4200 12400 -3500
rect 11600 -4300 12400 -4200
rect 10500 -5700 10600 -5000
rect 11200 -5700 11300 -5000
rect 10500 -5800 11300 -5700
<< via4 >>
rect 2300 4800 2900 5500
rect 100 3300 700 4000
rect 1000 150 2000 200
rect 1000 50 2000 150
rect 1000 -350 2000 -250
rect 1000 -400 2000 -350
rect 5800 4800 6400 5500
rect 3600 3300 4200 4000
rect 1200 -4200 1800 -3500
rect 100 -5700 700 -5000
rect 9300 4800 9900 5500
rect 7100 3300 7700 4000
rect 4700 -4200 5300 -3500
rect 3600 -5700 4200 -5000
rect 8000 150 9000 200
rect 8000 50 9000 150
rect 8000 -350 9000 -250
rect 8000 -400 9000 -350
rect 12800 4800 13400 5500
rect 10600 3300 11200 4000
rect 8200 -4200 8800 -3500
rect 7100 -5700 7700 -5000
rect 11700 -4200 12300 -3500
rect 10600 -5700 11200 -5000
<< metal5 >>
rect 0 4100 1400 5700
rect 12100 5600 13500 5700
rect 2200 5500 13500 5600
rect 2200 4800 2300 5500
rect 2900 4800 5800 5500
rect 6400 4800 9300 5500
rect 9900 4800 12800 5500
rect 13400 4800 13500 5500
rect 2200 4700 13500 4800
rect 0 4000 11300 4100
rect 0 3300 100 4000
rect 700 3300 3600 4000
rect 4200 3300 7100 4000
rect 7700 3300 10600 4000
rect 11200 3300 11300 4000
rect 0 3200 11300 3300
rect -50 200 13500 250
rect -50 50 1000 200
rect 2000 50 8000 200
rect 9000 50 13500 200
rect -50 0 13500 50
rect -50 -250 13500 -200
rect -50 -400 1000 -250
rect 2000 -400 8000 -250
rect 9000 -400 13500 -250
rect -50 -450 13500 -400
rect 1100 -3500 13500 -3400
rect 1100 -4200 1200 -3500
rect 1800 -4200 4700 -3500
rect 5300 -4200 8200 -3500
rect 8800 -4200 11700 -3500
rect 12300 -4200 13500 -3500
rect 1100 -4300 13500 -4200
rect 0 -5000 11300 -4900
rect 0 -5700 100 -5000
rect 700 -5700 3600 -5000
rect 4200 -5700 7100 -5000
rect 7700 -5700 10600 -5000
rect 11200 -5700 11300 -5000
rect 0 -5800 11300 -5700
rect 0 -5900 1400 -5800
rect 12100 -5900 13500 -4300
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_0
timestamp 1663721312
transform 1 0 0 0 1 0
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_1
timestamp 1663721312
transform 1 0 3500 0 1 0
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_2
timestamp 1663721312
transform 1 0 7000 0 1 0
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_3
timestamp 1663721312
transform 1 0 10500 0 1 0
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_4
timestamp 1663721312
transform 1 0 10500 0 1 -3500
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_5
timestamp 1663721312
transform 1 0 7000 0 1 -3500
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_6
timestamp 1663721312
transform 1 0 3500 0 1 -3500
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_7
timestamp 1663721312
transform 1 0 0 0 1 -3500
box 0 0 2569 3258
<< labels >>
rlabel metal5 12100 5600 13500 5700 1 SD1R
rlabel metal5 0 5600 1400 5700 1 SD1L
rlabel metal5 0 -5900 1400 -5800 1 SD2L
rlabel metal5 12100 -5900 13500 -5800 1 SD2R
rlabel metal5 -50 0 0 250 1 GL
rlabel metal5 -50 -450 0 -200 1 GR
rlabel metal2 7015 2860 7050 2890 1 SUB
rlabel metal2 3515 2860 3550 2890 1 SUB
rlabel metal2 10515 2860 10550 2890 1 SUB
rlabel metal2 3515 -3390 3550 -3360 1 SUB
rlabel metal2 7015 -3390 7050 -3360 1 SUB
rlabel metal2 10515 -3390 10550 -3360 1 SUB
rlabel metal2 6300 -6150 6800 -6050 1 SUB
<< end >>
