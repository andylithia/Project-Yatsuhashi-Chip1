magic
tech sky130A
timestamp 1660789662
use hash_m1m2_W2p5L2p5  hash_m1m2_W2p5L2p5_0
timestamp 1660275339
transform 1 0 -50 0 1 -50
box 50 -550 300 -300
use hash_m1m2_W2p5L2p5  hash_m1m2_W2p5L2p5_1
timestamp 1660275339
transform 1 0 200 0 1 -50
box 50 -550 300 -300
use hash_m1m2_W2p5L2p5  hash_m1m2_W2p5L2p5_2
timestamp 1660275339
transform 1 0 -50 0 1 -300
box 50 -550 300 -300
use hash_m1m2_W2p5L2p5  hash_m1m2_W2p5L2p5_3
timestamp 1660275339
transform 1 0 200 0 1 -300
box 50 -550 300 -300
<< end >>
