magic
tech sky130A
magscale 1 2
timestamp 1664327147
<< pwell >>
rect 1400 400 6538 6916
rect 7700 400 12838 6916
rect 14000 400 19138 6916
rect 20300 400 25438 6916
rect 1400 -7200 6538 -684
rect 7700 -7200 12838 -684
rect 14000 -7200 19138 -684
rect 20300 -7200 25438 -684
<< mvnmos >>
rect 1628 658 1728 6658
rect 1786 658 1886 6658
rect 1944 658 2044 6658
rect 2102 658 2202 6658
rect 2260 658 2360 6658
rect 2418 658 2518 6658
rect 2576 658 2676 6658
rect 2734 658 2834 6658
rect 2892 658 2992 6658
rect 3050 658 3150 6658
rect 3208 658 3308 6658
rect 3366 658 3466 6658
rect 3524 658 3624 6658
rect 3682 658 3782 6658
rect 3840 658 3940 6658
rect 3998 658 4098 6658
rect 4156 658 4256 6658
rect 4314 658 4414 6658
rect 4472 658 4572 6658
rect 4630 658 4730 6658
rect 4788 658 4888 6658
rect 4946 658 5046 6658
rect 5104 658 5204 6658
rect 5262 658 5362 6658
rect 5420 658 5520 6658
rect 5578 658 5678 6658
rect 5736 658 5836 6658
rect 5894 658 5994 6658
rect 6052 658 6152 6658
rect 6210 658 6310 6658
rect 7928 658 8028 6658
rect 8086 658 8186 6658
rect 8244 658 8344 6658
rect 8402 658 8502 6658
rect 8560 658 8660 6658
rect 8718 658 8818 6658
rect 8876 658 8976 6658
rect 9034 658 9134 6658
rect 9192 658 9292 6658
rect 9350 658 9450 6658
rect 9508 658 9608 6658
rect 9666 658 9766 6658
rect 9824 658 9924 6658
rect 9982 658 10082 6658
rect 10140 658 10240 6658
rect 10298 658 10398 6658
rect 10456 658 10556 6658
rect 10614 658 10714 6658
rect 10772 658 10872 6658
rect 10930 658 11030 6658
rect 11088 658 11188 6658
rect 11246 658 11346 6658
rect 11404 658 11504 6658
rect 11562 658 11662 6658
rect 11720 658 11820 6658
rect 11878 658 11978 6658
rect 12036 658 12136 6658
rect 12194 658 12294 6658
rect 12352 658 12452 6658
rect 12510 658 12610 6658
rect 14228 658 14328 6658
rect 14386 658 14486 6658
rect 14544 658 14644 6658
rect 14702 658 14802 6658
rect 14860 658 14960 6658
rect 15018 658 15118 6658
rect 15176 658 15276 6658
rect 15334 658 15434 6658
rect 15492 658 15592 6658
rect 15650 658 15750 6658
rect 15808 658 15908 6658
rect 15966 658 16066 6658
rect 16124 658 16224 6658
rect 16282 658 16382 6658
rect 16440 658 16540 6658
rect 16598 658 16698 6658
rect 16756 658 16856 6658
rect 16914 658 17014 6658
rect 17072 658 17172 6658
rect 17230 658 17330 6658
rect 17388 658 17488 6658
rect 17546 658 17646 6658
rect 17704 658 17804 6658
rect 17862 658 17962 6658
rect 18020 658 18120 6658
rect 18178 658 18278 6658
rect 18336 658 18436 6658
rect 18494 658 18594 6658
rect 18652 658 18752 6658
rect 18810 658 18910 6658
rect 20528 658 20628 6658
rect 20686 658 20786 6658
rect 20844 658 20944 6658
rect 21002 658 21102 6658
rect 21160 658 21260 6658
rect 21318 658 21418 6658
rect 21476 658 21576 6658
rect 21634 658 21734 6658
rect 21792 658 21892 6658
rect 21950 658 22050 6658
rect 22108 658 22208 6658
rect 22266 658 22366 6658
rect 22424 658 22524 6658
rect 22582 658 22682 6658
rect 22740 658 22840 6658
rect 22898 658 22998 6658
rect 23056 658 23156 6658
rect 23214 658 23314 6658
rect 23372 658 23472 6658
rect 23530 658 23630 6658
rect 23688 658 23788 6658
rect 23846 658 23946 6658
rect 24004 658 24104 6658
rect 24162 658 24262 6658
rect 24320 658 24420 6658
rect 24478 658 24578 6658
rect 24636 658 24736 6658
rect 24794 658 24894 6658
rect 24952 658 25052 6658
rect 25110 658 25210 6658
rect 1628 -6942 1728 -942
rect 1786 -6942 1886 -942
rect 1944 -6942 2044 -942
rect 2102 -6942 2202 -942
rect 2260 -6942 2360 -942
rect 2418 -6942 2518 -942
rect 2576 -6942 2676 -942
rect 2734 -6942 2834 -942
rect 2892 -6942 2992 -942
rect 3050 -6942 3150 -942
rect 3208 -6942 3308 -942
rect 3366 -6942 3466 -942
rect 3524 -6942 3624 -942
rect 3682 -6942 3782 -942
rect 3840 -6942 3940 -942
rect 3998 -6942 4098 -942
rect 4156 -6942 4256 -942
rect 4314 -6942 4414 -942
rect 4472 -6942 4572 -942
rect 4630 -6942 4730 -942
rect 4788 -6942 4888 -942
rect 4946 -6942 5046 -942
rect 5104 -6942 5204 -942
rect 5262 -6942 5362 -942
rect 5420 -6942 5520 -942
rect 5578 -6942 5678 -942
rect 5736 -6942 5836 -942
rect 5894 -6942 5994 -942
rect 6052 -6942 6152 -942
rect 6210 -6942 6310 -942
rect 7928 -6942 8028 -942
rect 8086 -6942 8186 -942
rect 8244 -6942 8344 -942
rect 8402 -6942 8502 -942
rect 8560 -6942 8660 -942
rect 8718 -6942 8818 -942
rect 8876 -6942 8976 -942
rect 9034 -6942 9134 -942
rect 9192 -6942 9292 -942
rect 9350 -6942 9450 -942
rect 9508 -6942 9608 -942
rect 9666 -6942 9766 -942
rect 9824 -6942 9924 -942
rect 9982 -6942 10082 -942
rect 10140 -6942 10240 -942
rect 10298 -6942 10398 -942
rect 10456 -6942 10556 -942
rect 10614 -6942 10714 -942
rect 10772 -6942 10872 -942
rect 10930 -6942 11030 -942
rect 11088 -6942 11188 -942
rect 11246 -6942 11346 -942
rect 11404 -6942 11504 -942
rect 11562 -6942 11662 -942
rect 11720 -6942 11820 -942
rect 11878 -6942 11978 -942
rect 12036 -6942 12136 -942
rect 12194 -6942 12294 -942
rect 12352 -6942 12452 -942
rect 12510 -6942 12610 -942
rect 14228 -6942 14328 -942
rect 14386 -6942 14486 -942
rect 14544 -6942 14644 -942
rect 14702 -6942 14802 -942
rect 14860 -6942 14960 -942
rect 15018 -6942 15118 -942
rect 15176 -6942 15276 -942
rect 15334 -6942 15434 -942
rect 15492 -6942 15592 -942
rect 15650 -6942 15750 -942
rect 15808 -6942 15908 -942
rect 15966 -6942 16066 -942
rect 16124 -6942 16224 -942
rect 16282 -6942 16382 -942
rect 16440 -6942 16540 -942
rect 16598 -6942 16698 -942
rect 16756 -6942 16856 -942
rect 16914 -6942 17014 -942
rect 17072 -6942 17172 -942
rect 17230 -6942 17330 -942
rect 17388 -6942 17488 -942
rect 17546 -6942 17646 -942
rect 17704 -6942 17804 -942
rect 17862 -6942 17962 -942
rect 18020 -6942 18120 -942
rect 18178 -6942 18278 -942
rect 18336 -6942 18436 -942
rect 18494 -6942 18594 -942
rect 18652 -6942 18752 -942
rect 18810 -6942 18910 -942
rect 20528 -6942 20628 -942
rect 20686 -6942 20786 -942
rect 20844 -6942 20944 -942
rect 21002 -6942 21102 -942
rect 21160 -6942 21260 -942
rect 21318 -6942 21418 -942
rect 21476 -6942 21576 -942
rect 21634 -6942 21734 -942
rect 21792 -6942 21892 -942
rect 21950 -6942 22050 -942
rect 22108 -6942 22208 -942
rect 22266 -6942 22366 -942
rect 22424 -6942 22524 -942
rect 22582 -6942 22682 -942
rect 22740 -6942 22840 -942
rect 22898 -6942 22998 -942
rect 23056 -6942 23156 -942
rect 23214 -6942 23314 -942
rect 23372 -6942 23472 -942
rect 23530 -6942 23630 -942
rect 23688 -6942 23788 -942
rect 23846 -6942 23946 -942
rect 24004 -6942 24104 -942
rect 24162 -6942 24262 -942
rect 24320 -6942 24420 -942
rect 24478 -6942 24578 -942
rect 24636 -6942 24736 -942
rect 24794 -6942 24894 -942
rect 24952 -6942 25052 -942
rect 25110 -6942 25210 -942
<< mvndiff >>
rect 1570 6646 1628 6658
rect 1570 670 1582 6646
rect 1616 670 1628 6646
rect 1570 658 1628 670
rect 1728 6646 1786 6658
rect 1728 670 1740 6646
rect 1774 670 1786 6646
rect 1728 658 1786 670
rect 1886 6646 1944 6658
rect 1886 670 1898 6646
rect 1932 670 1944 6646
rect 1886 658 1944 670
rect 2044 6646 2102 6658
rect 2044 670 2056 6646
rect 2090 670 2102 6646
rect 2044 658 2102 670
rect 2202 6646 2260 6658
rect 2202 670 2214 6646
rect 2248 670 2260 6646
rect 2202 658 2260 670
rect 2360 6646 2418 6658
rect 2360 670 2372 6646
rect 2406 670 2418 6646
rect 2360 658 2418 670
rect 2518 6646 2576 6658
rect 2518 670 2530 6646
rect 2564 670 2576 6646
rect 2518 658 2576 670
rect 2676 6646 2734 6658
rect 2676 670 2688 6646
rect 2722 670 2734 6646
rect 2676 658 2734 670
rect 2834 6646 2892 6658
rect 2834 670 2846 6646
rect 2880 670 2892 6646
rect 2834 658 2892 670
rect 2992 6646 3050 6658
rect 2992 670 3004 6646
rect 3038 670 3050 6646
rect 2992 658 3050 670
rect 3150 6646 3208 6658
rect 3150 670 3162 6646
rect 3196 670 3208 6646
rect 3150 658 3208 670
rect 3308 6646 3366 6658
rect 3308 670 3320 6646
rect 3354 670 3366 6646
rect 3308 658 3366 670
rect 3466 6646 3524 6658
rect 3466 670 3478 6646
rect 3512 670 3524 6646
rect 3466 658 3524 670
rect 3624 6646 3682 6658
rect 3624 670 3636 6646
rect 3670 670 3682 6646
rect 3624 658 3682 670
rect 3782 6646 3840 6658
rect 3782 670 3794 6646
rect 3828 670 3840 6646
rect 3782 658 3840 670
rect 3940 6646 3998 6658
rect 3940 670 3952 6646
rect 3986 670 3998 6646
rect 3940 658 3998 670
rect 4098 6646 4156 6658
rect 4098 670 4110 6646
rect 4144 670 4156 6646
rect 4098 658 4156 670
rect 4256 6646 4314 6658
rect 4256 670 4268 6646
rect 4302 670 4314 6646
rect 4256 658 4314 670
rect 4414 6646 4472 6658
rect 4414 670 4426 6646
rect 4460 670 4472 6646
rect 4414 658 4472 670
rect 4572 6646 4630 6658
rect 4572 670 4584 6646
rect 4618 670 4630 6646
rect 4572 658 4630 670
rect 4730 6646 4788 6658
rect 4730 670 4742 6646
rect 4776 670 4788 6646
rect 4730 658 4788 670
rect 4888 6646 4946 6658
rect 4888 670 4900 6646
rect 4934 670 4946 6646
rect 4888 658 4946 670
rect 5046 6646 5104 6658
rect 5046 670 5058 6646
rect 5092 670 5104 6646
rect 5046 658 5104 670
rect 5204 6646 5262 6658
rect 5204 670 5216 6646
rect 5250 670 5262 6646
rect 5204 658 5262 670
rect 5362 6646 5420 6658
rect 5362 670 5374 6646
rect 5408 670 5420 6646
rect 5362 658 5420 670
rect 5520 6646 5578 6658
rect 5520 670 5532 6646
rect 5566 670 5578 6646
rect 5520 658 5578 670
rect 5678 6646 5736 6658
rect 5678 670 5690 6646
rect 5724 670 5736 6646
rect 5678 658 5736 670
rect 5836 6646 5894 6658
rect 5836 670 5848 6646
rect 5882 670 5894 6646
rect 5836 658 5894 670
rect 5994 6646 6052 6658
rect 5994 670 6006 6646
rect 6040 670 6052 6646
rect 5994 658 6052 670
rect 6152 6646 6210 6658
rect 6152 670 6164 6646
rect 6198 670 6210 6646
rect 6152 658 6210 670
rect 6310 6646 6368 6658
rect 6310 670 6322 6646
rect 6356 670 6368 6646
rect 6310 658 6368 670
rect 7870 6646 7928 6658
rect 7870 670 7882 6646
rect 7916 670 7928 6646
rect 7870 658 7928 670
rect 8028 6646 8086 6658
rect 8028 670 8040 6646
rect 8074 670 8086 6646
rect 8028 658 8086 670
rect 8186 6646 8244 6658
rect 8186 670 8198 6646
rect 8232 670 8244 6646
rect 8186 658 8244 670
rect 8344 6646 8402 6658
rect 8344 670 8356 6646
rect 8390 670 8402 6646
rect 8344 658 8402 670
rect 8502 6646 8560 6658
rect 8502 670 8514 6646
rect 8548 670 8560 6646
rect 8502 658 8560 670
rect 8660 6646 8718 6658
rect 8660 670 8672 6646
rect 8706 670 8718 6646
rect 8660 658 8718 670
rect 8818 6646 8876 6658
rect 8818 670 8830 6646
rect 8864 670 8876 6646
rect 8818 658 8876 670
rect 8976 6646 9034 6658
rect 8976 670 8988 6646
rect 9022 670 9034 6646
rect 8976 658 9034 670
rect 9134 6646 9192 6658
rect 9134 670 9146 6646
rect 9180 670 9192 6646
rect 9134 658 9192 670
rect 9292 6646 9350 6658
rect 9292 670 9304 6646
rect 9338 670 9350 6646
rect 9292 658 9350 670
rect 9450 6646 9508 6658
rect 9450 670 9462 6646
rect 9496 670 9508 6646
rect 9450 658 9508 670
rect 9608 6646 9666 6658
rect 9608 670 9620 6646
rect 9654 670 9666 6646
rect 9608 658 9666 670
rect 9766 6646 9824 6658
rect 9766 670 9778 6646
rect 9812 670 9824 6646
rect 9766 658 9824 670
rect 9924 6646 9982 6658
rect 9924 670 9936 6646
rect 9970 670 9982 6646
rect 9924 658 9982 670
rect 10082 6646 10140 6658
rect 10082 670 10094 6646
rect 10128 670 10140 6646
rect 10082 658 10140 670
rect 10240 6646 10298 6658
rect 10240 670 10252 6646
rect 10286 670 10298 6646
rect 10240 658 10298 670
rect 10398 6646 10456 6658
rect 10398 670 10410 6646
rect 10444 670 10456 6646
rect 10398 658 10456 670
rect 10556 6646 10614 6658
rect 10556 670 10568 6646
rect 10602 670 10614 6646
rect 10556 658 10614 670
rect 10714 6646 10772 6658
rect 10714 670 10726 6646
rect 10760 670 10772 6646
rect 10714 658 10772 670
rect 10872 6646 10930 6658
rect 10872 670 10884 6646
rect 10918 670 10930 6646
rect 10872 658 10930 670
rect 11030 6646 11088 6658
rect 11030 670 11042 6646
rect 11076 670 11088 6646
rect 11030 658 11088 670
rect 11188 6646 11246 6658
rect 11188 670 11200 6646
rect 11234 670 11246 6646
rect 11188 658 11246 670
rect 11346 6646 11404 6658
rect 11346 670 11358 6646
rect 11392 670 11404 6646
rect 11346 658 11404 670
rect 11504 6646 11562 6658
rect 11504 670 11516 6646
rect 11550 670 11562 6646
rect 11504 658 11562 670
rect 11662 6646 11720 6658
rect 11662 670 11674 6646
rect 11708 670 11720 6646
rect 11662 658 11720 670
rect 11820 6646 11878 6658
rect 11820 670 11832 6646
rect 11866 670 11878 6646
rect 11820 658 11878 670
rect 11978 6646 12036 6658
rect 11978 670 11990 6646
rect 12024 670 12036 6646
rect 11978 658 12036 670
rect 12136 6646 12194 6658
rect 12136 670 12148 6646
rect 12182 670 12194 6646
rect 12136 658 12194 670
rect 12294 6646 12352 6658
rect 12294 670 12306 6646
rect 12340 670 12352 6646
rect 12294 658 12352 670
rect 12452 6646 12510 6658
rect 12452 670 12464 6646
rect 12498 670 12510 6646
rect 12452 658 12510 670
rect 12610 6646 12668 6658
rect 12610 670 12622 6646
rect 12656 670 12668 6646
rect 12610 658 12668 670
rect 14170 6646 14228 6658
rect 14170 670 14182 6646
rect 14216 670 14228 6646
rect 14170 658 14228 670
rect 14328 6646 14386 6658
rect 14328 670 14340 6646
rect 14374 670 14386 6646
rect 14328 658 14386 670
rect 14486 6646 14544 6658
rect 14486 670 14498 6646
rect 14532 670 14544 6646
rect 14486 658 14544 670
rect 14644 6646 14702 6658
rect 14644 670 14656 6646
rect 14690 670 14702 6646
rect 14644 658 14702 670
rect 14802 6646 14860 6658
rect 14802 670 14814 6646
rect 14848 670 14860 6646
rect 14802 658 14860 670
rect 14960 6646 15018 6658
rect 14960 670 14972 6646
rect 15006 670 15018 6646
rect 14960 658 15018 670
rect 15118 6646 15176 6658
rect 15118 670 15130 6646
rect 15164 670 15176 6646
rect 15118 658 15176 670
rect 15276 6646 15334 6658
rect 15276 670 15288 6646
rect 15322 670 15334 6646
rect 15276 658 15334 670
rect 15434 6646 15492 6658
rect 15434 670 15446 6646
rect 15480 670 15492 6646
rect 15434 658 15492 670
rect 15592 6646 15650 6658
rect 15592 670 15604 6646
rect 15638 670 15650 6646
rect 15592 658 15650 670
rect 15750 6646 15808 6658
rect 15750 670 15762 6646
rect 15796 670 15808 6646
rect 15750 658 15808 670
rect 15908 6646 15966 6658
rect 15908 670 15920 6646
rect 15954 670 15966 6646
rect 15908 658 15966 670
rect 16066 6646 16124 6658
rect 16066 670 16078 6646
rect 16112 670 16124 6646
rect 16066 658 16124 670
rect 16224 6646 16282 6658
rect 16224 670 16236 6646
rect 16270 670 16282 6646
rect 16224 658 16282 670
rect 16382 6646 16440 6658
rect 16382 670 16394 6646
rect 16428 670 16440 6646
rect 16382 658 16440 670
rect 16540 6646 16598 6658
rect 16540 670 16552 6646
rect 16586 670 16598 6646
rect 16540 658 16598 670
rect 16698 6646 16756 6658
rect 16698 670 16710 6646
rect 16744 670 16756 6646
rect 16698 658 16756 670
rect 16856 6646 16914 6658
rect 16856 670 16868 6646
rect 16902 670 16914 6646
rect 16856 658 16914 670
rect 17014 6646 17072 6658
rect 17014 670 17026 6646
rect 17060 670 17072 6646
rect 17014 658 17072 670
rect 17172 6646 17230 6658
rect 17172 670 17184 6646
rect 17218 670 17230 6646
rect 17172 658 17230 670
rect 17330 6646 17388 6658
rect 17330 670 17342 6646
rect 17376 670 17388 6646
rect 17330 658 17388 670
rect 17488 6646 17546 6658
rect 17488 670 17500 6646
rect 17534 670 17546 6646
rect 17488 658 17546 670
rect 17646 6646 17704 6658
rect 17646 670 17658 6646
rect 17692 670 17704 6646
rect 17646 658 17704 670
rect 17804 6646 17862 6658
rect 17804 670 17816 6646
rect 17850 670 17862 6646
rect 17804 658 17862 670
rect 17962 6646 18020 6658
rect 17962 670 17974 6646
rect 18008 670 18020 6646
rect 17962 658 18020 670
rect 18120 6646 18178 6658
rect 18120 670 18132 6646
rect 18166 670 18178 6646
rect 18120 658 18178 670
rect 18278 6646 18336 6658
rect 18278 670 18290 6646
rect 18324 670 18336 6646
rect 18278 658 18336 670
rect 18436 6646 18494 6658
rect 18436 670 18448 6646
rect 18482 670 18494 6646
rect 18436 658 18494 670
rect 18594 6646 18652 6658
rect 18594 670 18606 6646
rect 18640 670 18652 6646
rect 18594 658 18652 670
rect 18752 6646 18810 6658
rect 18752 670 18764 6646
rect 18798 670 18810 6646
rect 18752 658 18810 670
rect 18910 6646 18968 6658
rect 18910 670 18922 6646
rect 18956 670 18968 6646
rect 18910 658 18968 670
rect 20470 6646 20528 6658
rect 20470 670 20482 6646
rect 20516 670 20528 6646
rect 20470 658 20528 670
rect 20628 6646 20686 6658
rect 20628 670 20640 6646
rect 20674 670 20686 6646
rect 20628 658 20686 670
rect 20786 6646 20844 6658
rect 20786 670 20798 6646
rect 20832 670 20844 6646
rect 20786 658 20844 670
rect 20944 6646 21002 6658
rect 20944 670 20956 6646
rect 20990 670 21002 6646
rect 20944 658 21002 670
rect 21102 6646 21160 6658
rect 21102 670 21114 6646
rect 21148 670 21160 6646
rect 21102 658 21160 670
rect 21260 6646 21318 6658
rect 21260 670 21272 6646
rect 21306 670 21318 6646
rect 21260 658 21318 670
rect 21418 6646 21476 6658
rect 21418 670 21430 6646
rect 21464 670 21476 6646
rect 21418 658 21476 670
rect 21576 6646 21634 6658
rect 21576 670 21588 6646
rect 21622 670 21634 6646
rect 21576 658 21634 670
rect 21734 6646 21792 6658
rect 21734 670 21746 6646
rect 21780 670 21792 6646
rect 21734 658 21792 670
rect 21892 6646 21950 6658
rect 21892 670 21904 6646
rect 21938 670 21950 6646
rect 21892 658 21950 670
rect 22050 6646 22108 6658
rect 22050 670 22062 6646
rect 22096 670 22108 6646
rect 22050 658 22108 670
rect 22208 6646 22266 6658
rect 22208 670 22220 6646
rect 22254 670 22266 6646
rect 22208 658 22266 670
rect 22366 6646 22424 6658
rect 22366 670 22378 6646
rect 22412 670 22424 6646
rect 22366 658 22424 670
rect 22524 6646 22582 6658
rect 22524 670 22536 6646
rect 22570 670 22582 6646
rect 22524 658 22582 670
rect 22682 6646 22740 6658
rect 22682 670 22694 6646
rect 22728 670 22740 6646
rect 22682 658 22740 670
rect 22840 6646 22898 6658
rect 22840 670 22852 6646
rect 22886 670 22898 6646
rect 22840 658 22898 670
rect 22998 6646 23056 6658
rect 22998 670 23010 6646
rect 23044 670 23056 6646
rect 22998 658 23056 670
rect 23156 6646 23214 6658
rect 23156 670 23168 6646
rect 23202 670 23214 6646
rect 23156 658 23214 670
rect 23314 6646 23372 6658
rect 23314 670 23326 6646
rect 23360 670 23372 6646
rect 23314 658 23372 670
rect 23472 6646 23530 6658
rect 23472 670 23484 6646
rect 23518 670 23530 6646
rect 23472 658 23530 670
rect 23630 6646 23688 6658
rect 23630 670 23642 6646
rect 23676 670 23688 6646
rect 23630 658 23688 670
rect 23788 6646 23846 6658
rect 23788 670 23800 6646
rect 23834 670 23846 6646
rect 23788 658 23846 670
rect 23946 6646 24004 6658
rect 23946 670 23958 6646
rect 23992 670 24004 6646
rect 23946 658 24004 670
rect 24104 6646 24162 6658
rect 24104 670 24116 6646
rect 24150 670 24162 6646
rect 24104 658 24162 670
rect 24262 6646 24320 6658
rect 24262 670 24274 6646
rect 24308 670 24320 6646
rect 24262 658 24320 670
rect 24420 6646 24478 6658
rect 24420 670 24432 6646
rect 24466 670 24478 6646
rect 24420 658 24478 670
rect 24578 6646 24636 6658
rect 24578 670 24590 6646
rect 24624 670 24636 6646
rect 24578 658 24636 670
rect 24736 6646 24794 6658
rect 24736 670 24748 6646
rect 24782 670 24794 6646
rect 24736 658 24794 670
rect 24894 6646 24952 6658
rect 24894 670 24906 6646
rect 24940 670 24952 6646
rect 24894 658 24952 670
rect 25052 6646 25110 6658
rect 25052 670 25064 6646
rect 25098 670 25110 6646
rect 25052 658 25110 670
rect 25210 6646 25268 6658
rect 25210 670 25222 6646
rect 25256 670 25268 6646
rect 25210 658 25268 670
rect 1570 -954 1628 -942
rect 1570 -6930 1582 -954
rect 1616 -6930 1628 -954
rect 1570 -6942 1628 -6930
rect 1728 -954 1786 -942
rect 1728 -6930 1740 -954
rect 1774 -6930 1786 -954
rect 1728 -6942 1786 -6930
rect 1886 -954 1944 -942
rect 1886 -6930 1898 -954
rect 1932 -6930 1944 -954
rect 1886 -6942 1944 -6930
rect 2044 -954 2102 -942
rect 2044 -6930 2056 -954
rect 2090 -6930 2102 -954
rect 2044 -6942 2102 -6930
rect 2202 -954 2260 -942
rect 2202 -6930 2214 -954
rect 2248 -6930 2260 -954
rect 2202 -6942 2260 -6930
rect 2360 -954 2418 -942
rect 2360 -6930 2372 -954
rect 2406 -6930 2418 -954
rect 2360 -6942 2418 -6930
rect 2518 -954 2576 -942
rect 2518 -6930 2530 -954
rect 2564 -6930 2576 -954
rect 2518 -6942 2576 -6930
rect 2676 -954 2734 -942
rect 2676 -6930 2688 -954
rect 2722 -6930 2734 -954
rect 2676 -6942 2734 -6930
rect 2834 -954 2892 -942
rect 2834 -6930 2846 -954
rect 2880 -6930 2892 -954
rect 2834 -6942 2892 -6930
rect 2992 -954 3050 -942
rect 2992 -6930 3004 -954
rect 3038 -6930 3050 -954
rect 2992 -6942 3050 -6930
rect 3150 -954 3208 -942
rect 3150 -6930 3162 -954
rect 3196 -6930 3208 -954
rect 3150 -6942 3208 -6930
rect 3308 -954 3366 -942
rect 3308 -6930 3320 -954
rect 3354 -6930 3366 -954
rect 3308 -6942 3366 -6930
rect 3466 -954 3524 -942
rect 3466 -6930 3478 -954
rect 3512 -6930 3524 -954
rect 3466 -6942 3524 -6930
rect 3624 -954 3682 -942
rect 3624 -6930 3636 -954
rect 3670 -6930 3682 -954
rect 3624 -6942 3682 -6930
rect 3782 -954 3840 -942
rect 3782 -6930 3794 -954
rect 3828 -6930 3840 -954
rect 3782 -6942 3840 -6930
rect 3940 -954 3998 -942
rect 3940 -6930 3952 -954
rect 3986 -6930 3998 -954
rect 3940 -6942 3998 -6930
rect 4098 -954 4156 -942
rect 4098 -6930 4110 -954
rect 4144 -6930 4156 -954
rect 4098 -6942 4156 -6930
rect 4256 -954 4314 -942
rect 4256 -6930 4268 -954
rect 4302 -6930 4314 -954
rect 4256 -6942 4314 -6930
rect 4414 -954 4472 -942
rect 4414 -6930 4426 -954
rect 4460 -6930 4472 -954
rect 4414 -6942 4472 -6930
rect 4572 -954 4630 -942
rect 4572 -6930 4584 -954
rect 4618 -6930 4630 -954
rect 4572 -6942 4630 -6930
rect 4730 -954 4788 -942
rect 4730 -6930 4742 -954
rect 4776 -6930 4788 -954
rect 4730 -6942 4788 -6930
rect 4888 -954 4946 -942
rect 4888 -6930 4900 -954
rect 4934 -6930 4946 -954
rect 4888 -6942 4946 -6930
rect 5046 -954 5104 -942
rect 5046 -6930 5058 -954
rect 5092 -6930 5104 -954
rect 5046 -6942 5104 -6930
rect 5204 -954 5262 -942
rect 5204 -6930 5216 -954
rect 5250 -6930 5262 -954
rect 5204 -6942 5262 -6930
rect 5362 -954 5420 -942
rect 5362 -6930 5374 -954
rect 5408 -6930 5420 -954
rect 5362 -6942 5420 -6930
rect 5520 -954 5578 -942
rect 5520 -6930 5532 -954
rect 5566 -6930 5578 -954
rect 5520 -6942 5578 -6930
rect 5678 -954 5736 -942
rect 5678 -6930 5690 -954
rect 5724 -6930 5736 -954
rect 5678 -6942 5736 -6930
rect 5836 -954 5894 -942
rect 5836 -6930 5848 -954
rect 5882 -6930 5894 -954
rect 5836 -6942 5894 -6930
rect 5994 -954 6052 -942
rect 5994 -6930 6006 -954
rect 6040 -6930 6052 -954
rect 5994 -6942 6052 -6930
rect 6152 -954 6210 -942
rect 6152 -6930 6164 -954
rect 6198 -6930 6210 -954
rect 6152 -6942 6210 -6930
rect 6310 -954 6368 -942
rect 6310 -6930 6322 -954
rect 6356 -6930 6368 -954
rect 6310 -6942 6368 -6930
rect 7870 -954 7928 -942
rect 7870 -6930 7882 -954
rect 7916 -6930 7928 -954
rect 7870 -6942 7928 -6930
rect 8028 -954 8086 -942
rect 8028 -6930 8040 -954
rect 8074 -6930 8086 -954
rect 8028 -6942 8086 -6930
rect 8186 -954 8244 -942
rect 8186 -6930 8198 -954
rect 8232 -6930 8244 -954
rect 8186 -6942 8244 -6930
rect 8344 -954 8402 -942
rect 8344 -6930 8356 -954
rect 8390 -6930 8402 -954
rect 8344 -6942 8402 -6930
rect 8502 -954 8560 -942
rect 8502 -6930 8514 -954
rect 8548 -6930 8560 -954
rect 8502 -6942 8560 -6930
rect 8660 -954 8718 -942
rect 8660 -6930 8672 -954
rect 8706 -6930 8718 -954
rect 8660 -6942 8718 -6930
rect 8818 -954 8876 -942
rect 8818 -6930 8830 -954
rect 8864 -6930 8876 -954
rect 8818 -6942 8876 -6930
rect 8976 -954 9034 -942
rect 8976 -6930 8988 -954
rect 9022 -6930 9034 -954
rect 8976 -6942 9034 -6930
rect 9134 -954 9192 -942
rect 9134 -6930 9146 -954
rect 9180 -6930 9192 -954
rect 9134 -6942 9192 -6930
rect 9292 -954 9350 -942
rect 9292 -6930 9304 -954
rect 9338 -6930 9350 -954
rect 9292 -6942 9350 -6930
rect 9450 -954 9508 -942
rect 9450 -6930 9462 -954
rect 9496 -6930 9508 -954
rect 9450 -6942 9508 -6930
rect 9608 -954 9666 -942
rect 9608 -6930 9620 -954
rect 9654 -6930 9666 -954
rect 9608 -6942 9666 -6930
rect 9766 -954 9824 -942
rect 9766 -6930 9778 -954
rect 9812 -6930 9824 -954
rect 9766 -6942 9824 -6930
rect 9924 -954 9982 -942
rect 9924 -6930 9936 -954
rect 9970 -6930 9982 -954
rect 9924 -6942 9982 -6930
rect 10082 -954 10140 -942
rect 10082 -6930 10094 -954
rect 10128 -6930 10140 -954
rect 10082 -6942 10140 -6930
rect 10240 -954 10298 -942
rect 10240 -6930 10252 -954
rect 10286 -6930 10298 -954
rect 10240 -6942 10298 -6930
rect 10398 -954 10456 -942
rect 10398 -6930 10410 -954
rect 10444 -6930 10456 -954
rect 10398 -6942 10456 -6930
rect 10556 -954 10614 -942
rect 10556 -6930 10568 -954
rect 10602 -6930 10614 -954
rect 10556 -6942 10614 -6930
rect 10714 -954 10772 -942
rect 10714 -6930 10726 -954
rect 10760 -6930 10772 -954
rect 10714 -6942 10772 -6930
rect 10872 -954 10930 -942
rect 10872 -6930 10884 -954
rect 10918 -6930 10930 -954
rect 10872 -6942 10930 -6930
rect 11030 -954 11088 -942
rect 11030 -6930 11042 -954
rect 11076 -6930 11088 -954
rect 11030 -6942 11088 -6930
rect 11188 -954 11246 -942
rect 11188 -6930 11200 -954
rect 11234 -6930 11246 -954
rect 11188 -6942 11246 -6930
rect 11346 -954 11404 -942
rect 11346 -6930 11358 -954
rect 11392 -6930 11404 -954
rect 11346 -6942 11404 -6930
rect 11504 -954 11562 -942
rect 11504 -6930 11516 -954
rect 11550 -6930 11562 -954
rect 11504 -6942 11562 -6930
rect 11662 -954 11720 -942
rect 11662 -6930 11674 -954
rect 11708 -6930 11720 -954
rect 11662 -6942 11720 -6930
rect 11820 -954 11878 -942
rect 11820 -6930 11832 -954
rect 11866 -6930 11878 -954
rect 11820 -6942 11878 -6930
rect 11978 -954 12036 -942
rect 11978 -6930 11990 -954
rect 12024 -6930 12036 -954
rect 11978 -6942 12036 -6930
rect 12136 -954 12194 -942
rect 12136 -6930 12148 -954
rect 12182 -6930 12194 -954
rect 12136 -6942 12194 -6930
rect 12294 -954 12352 -942
rect 12294 -6930 12306 -954
rect 12340 -6930 12352 -954
rect 12294 -6942 12352 -6930
rect 12452 -954 12510 -942
rect 12452 -6930 12464 -954
rect 12498 -6930 12510 -954
rect 12452 -6942 12510 -6930
rect 12610 -954 12668 -942
rect 12610 -6930 12622 -954
rect 12656 -6930 12668 -954
rect 12610 -6942 12668 -6930
rect 14170 -954 14228 -942
rect 14170 -6930 14182 -954
rect 14216 -6930 14228 -954
rect 14170 -6942 14228 -6930
rect 14328 -954 14386 -942
rect 14328 -6930 14340 -954
rect 14374 -6930 14386 -954
rect 14328 -6942 14386 -6930
rect 14486 -954 14544 -942
rect 14486 -6930 14498 -954
rect 14532 -6930 14544 -954
rect 14486 -6942 14544 -6930
rect 14644 -954 14702 -942
rect 14644 -6930 14656 -954
rect 14690 -6930 14702 -954
rect 14644 -6942 14702 -6930
rect 14802 -954 14860 -942
rect 14802 -6930 14814 -954
rect 14848 -6930 14860 -954
rect 14802 -6942 14860 -6930
rect 14960 -954 15018 -942
rect 14960 -6930 14972 -954
rect 15006 -6930 15018 -954
rect 14960 -6942 15018 -6930
rect 15118 -954 15176 -942
rect 15118 -6930 15130 -954
rect 15164 -6930 15176 -954
rect 15118 -6942 15176 -6930
rect 15276 -954 15334 -942
rect 15276 -6930 15288 -954
rect 15322 -6930 15334 -954
rect 15276 -6942 15334 -6930
rect 15434 -954 15492 -942
rect 15434 -6930 15446 -954
rect 15480 -6930 15492 -954
rect 15434 -6942 15492 -6930
rect 15592 -954 15650 -942
rect 15592 -6930 15604 -954
rect 15638 -6930 15650 -954
rect 15592 -6942 15650 -6930
rect 15750 -954 15808 -942
rect 15750 -6930 15762 -954
rect 15796 -6930 15808 -954
rect 15750 -6942 15808 -6930
rect 15908 -954 15966 -942
rect 15908 -6930 15920 -954
rect 15954 -6930 15966 -954
rect 15908 -6942 15966 -6930
rect 16066 -954 16124 -942
rect 16066 -6930 16078 -954
rect 16112 -6930 16124 -954
rect 16066 -6942 16124 -6930
rect 16224 -954 16282 -942
rect 16224 -6930 16236 -954
rect 16270 -6930 16282 -954
rect 16224 -6942 16282 -6930
rect 16382 -954 16440 -942
rect 16382 -6930 16394 -954
rect 16428 -6930 16440 -954
rect 16382 -6942 16440 -6930
rect 16540 -954 16598 -942
rect 16540 -6930 16552 -954
rect 16586 -6930 16598 -954
rect 16540 -6942 16598 -6930
rect 16698 -954 16756 -942
rect 16698 -6930 16710 -954
rect 16744 -6930 16756 -954
rect 16698 -6942 16756 -6930
rect 16856 -954 16914 -942
rect 16856 -6930 16868 -954
rect 16902 -6930 16914 -954
rect 16856 -6942 16914 -6930
rect 17014 -954 17072 -942
rect 17014 -6930 17026 -954
rect 17060 -6930 17072 -954
rect 17014 -6942 17072 -6930
rect 17172 -954 17230 -942
rect 17172 -6930 17184 -954
rect 17218 -6930 17230 -954
rect 17172 -6942 17230 -6930
rect 17330 -954 17388 -942
rect 17330 -6930 17342 -954
rect 17376 -6930 17388 -954
rect 17330 -6942 17388 -6930
rect 17488 -954 17546 -942
rect 17488 -6930 17500 -954
rect 17534 -6930 17546 -954
rect 17488 -6942 17546 -6930
rect 17646 -954 17704 -942
rect 17646 -6930 17658 -954
rect 17692 -6930 17704 -954
rect 17646 -6942 17704 -6930
rect 17804 -954 17862 -942
rect 17804 -6930 17816 -954
rect 17850 -6930 17862 -954
rect 17804 -6942 17862 -6930
rect 17962 -954 18020 -942
rect 17962 -6930 17974 -954
rect 18008 -6930 18020 -954
rect 17962 -6942 18020 -6930
rect 18120 -954 18178 -942
rect 18120 -6930 18132 -954
rect 18166 -6930 18178 -954
rect 18120 -6942 18178 -6930
rect 18278 -954 18336 -942
rect 18278 -6930 18290 -954
rect 18324 -6930 18336 -954
rect 18278 -6942 18336 -6930
rect 18436 -954 18494 -942
rect 18436 -6930 18448 -954
rect 18482 -6930 18494 -954
rect 18436 -6942 18494 -6930
rect 18594 -954 18652 -942
rect 18594 -6930 18606 -954
rect 18640 -6930 18652 -954
rect 18594 -6942 18652 -6930
rect 18752 -954 18810 -942
rect 18752 -6930 18764 -954
rect 18798 -6930 18810 -954
rect 18752 -6942 18810 -6930
rect 18910 -954 18968 -942
rect 18910 -6930 18922 -954
rect 18956 -6930 18968 -954
rect 18910 -6942 18968 -6930
rect 20470 -954 20528 -942
rect 20470 -6930 20482 -954
rect 20516 -6930 20528 -954
rect 20470 -6942 20528 -6930
rect 20628 -954 20686 -942
rect 20628 -6930 20640 -954
rect 20674 -6930 20686 -954
rect 20628 -6942 20686 -6930
rect 20786 -954 20844 -942
rect 20786 -6930 20798 -954
rect 20832 -6930 20844 -954
rect 20786 -6942 20844 -6930
rect 20944 -954 21002 -942
rect 20944 -6930 20956 -954
rect 20990 -6930 21002 -954
rect 20944 -6942 21002 -6930
rect 21102 -954 21160 -942
rect 21102 -6930 21114 -954
rect 21148 -6930 21160 -954
rect 21102 -6942 21160 -6930
rect 21260 -954 21318 -942
rect 21260 -6930 21272 -954
rect 21306 -6930 21318 -954
rect 21260 -6942 21318 -6930
rect 21418 -954 21476 -942
rect 21418 -6930 21430 -954
rect 21464 -6930 21476 -954
rect 21418 -6942 21476 -6930
rect 21576 -954 21634 -942
rect 21576 -6930 21588 -954
rect 21622 -6930 21634 -954
rect 21576 -6942 21634 -6930
rect 21734 -954 21792 -942
rect 21734 -6930 21746 -954
rect 21780 -6930 21792 -954
rect 21734 -6942 21792 -6930
rect 21892 -954 21950 -942
rect 21892 -6930 21904 -954
rect 21938 -6930 21950 -954
rect 21892 -6942 21950 -6930
rect 22050 -954 22108 -942
rect 22050 -6930 22062 -954
rect 22096 -6930 22108 -954
rect 22050 -6942 22108 -6930
rect 22208 -954 22266 -942
rect 22208 -6930 22220 -954
rect 22254 -6930 22266 -954
rect 22208 -6942 22266 -6930
rect 22366 -954 22424 -942
rect 22366 -6930 22378 -954
rect 22412 -6930 22424 -954
rect 22366 -6942 22424 -6930
rect 22524 -954 22582 -942
rect 22524 -6930 22536 -954
rect 22570 -6930 22582 -954
rect 22524 -6942 22582 -6930
rect 22682 -954 22740 -942
rect 22682 -6930 22694 -954
rect 22728 -6930 22740 -954
rect 22682 -6942 22740 -6930
rect 22840 -954 22898 -942
rect 22840 -6930 22852 -954
rect 22886 -6930 22898 -954
rect 22840 -6942 22898 -6930
rect 22998 -954 23056 -942
rect 22998 -6930 23010 -954
rect 23044 -6930 23056 -954
rect 22998 -6942 23056 -6930
rect 23156 -954 23214 -942
rect 23156 -6930 23168 -954
rect 23202 -6930 23214 -954
rect 23156 -6942 23214 -6930
rect 23314 -954 23372 -942
rect 23314 -6930 23326 -954
rect 23360 -6930 23372 -954
rect 23314 -6942 23372 -6930
rect 23472 -954 23530 -942
rect 23472 -6930 23484 -954
rect 23518 -6930 23530 -954
rect 23472 -6942 23530 -6930
rect 23630 -954 23688 -942
rect 23630 -6930 23642 -954
rect 23676 -6930 23688 -954
rect 23630 -6942 23688 -6930
rect 23788 -954 23846 -942
rect 23788 -6930 23800 -954
rect 23834 -6930 23846 -954
rect 23788 -6942 23846 -6930
rect 23946 -954 24004 -942
rect 23946 -6930 23958 -954
rect 23992 -6930 24004 -954
rect 23946 -6942 24004 -6930
rect 24104 -954 24162 -942
rect 24104 -6930 24116 -954
rect 24150 -6930 24162 -954
rect 24104 -6942 24162 -6930
rect 24262 -954 24320 -942
rect 24262 -6930 24274 -954
rect 24308 -6930 24320 -954
rect 24262 -6942 24320 -6930
rect 24420 -954 24478 -942
rect 24420 -6930 24432 -954
rect 24466 -6930 24478 -954
rect 24420 -6942 24478 -6930
rect 24578 -954 24636 -942
rect 24578 -6930 24590 -954
rect 24624 -6930 24636 -954
rect 24578 -6942 24636 -6930
rect 24736 -954 24794 -942
rect 24736 -6930 24748 -954
rect 24782 -6930 24794 -954
rect 24736 -6942 24794 -6930
rect 24894 -954 24952 -942
rect 24894 -6930 24906 -954
rect 24940 -6930 24952 -954
rect 24894 -6942 24952 -6930
rect 25052 -954 25110 -942
rect 25052 -6930 25064 -954
rect 25098 -6930 25110 -954
rect 25052 -6942 25110 -6930
rect 25210 -954 25268 -942
rect 25210 -6930 25222 -954
rect 25256 -6930 25268 -954
rect 25210 -6942 25268 -6930
<< mvndiffc >>
rect 1582 670 1616 6646
rect 1740 670 1774 6646
rect 1898 670 1932 6646
rect 2056 670 2090 6646
rect 2214 670 2248 6646
rect 2372 670 2406 6646
rect 2530 670 2564 6646
rect 2688 670 2722 6646
rect 2846 670 2880 6646
rect 3004 670 3038 6646
rect 3162 670 3196 6646
rect 3320 670 3354 6646
rect 3478 670 3512 6646
rect 3636 670 3670 6646
rect 3794 670 3828 6646
rect 3952 670 3986 6646
rect 4110 670 4144 6646
rect 4268 670 4302 6646
rect 4426 670 4460 6646
rect 4584 670 4618 6646
rect 4742 670 4776 6646
rect 4900 670 4934 6646
rect 5058 670 5092 6646
rect 5216 670 5250 6646
rect 5374 670 5408 6646
rect 5532 670 5566 6646
rect 5690 670 5724 6646
rect 5848 670 5882 6646
rect 6006 670 6040 6646
rect 6164 670 6198 6646
rect 6322 670 6356 6646
rect 7882 670 7916 6646
rect 8040 670 8074 6646
rect 8198 670 8232 6646
rect 8356 670 8390 6646
rect 8514 670 8548 6646
rect 8672 670 8706 6646
rect 8830 670 8864 6646
rect 8988 670 9022 6646
rect 9146 670 9180 6646
rect 9304 670 9338 6646
rect 9462 670 9496 6646
rect 9620 670 9654 6646
rect 9778 670 9812 6646
rect 9936 670 9970 6646
rect 10094 670 10128 6646
rect 10252 670 10286 6646
rect 10410 670 10444 6646
rect 10568 670 10602 6646
rect 10726 670 10760 6646
rect 10884 670 10918 6646
rect 11042 670 11076 6646
rect 11200 670 11234 6646
rect 11358 670 11392 6646
rect 11516 670 11550 6646
rect 11674 670 11708 6646
rect 11832 670 11866 6646
rect 11990 670 12024 6646
rect 12148 670 12182 6646
rect 12306 670 12340 6646
rect 12464 670 12498 6646
rect 12622 670 12656 6646
rect 14182 670 14216 6646
rect 14340 670 14374 6646
rect 14498 670 14532 6646
rect 14656 670 14690 6646
rect 14814 670 14848 6646
rect 14972 670 15006 6646
rect 15130 670 15164 6646
rect 15288 670 15322 6646
rect 15446 670 15480 6646
rect 15604 670 15638 6646
rect 15762 670 15796 6646
rect 15920 670 15954 6646
rect 16078 670 16112 6646
rect 16236 670 16270 6646
rect 16394 670 16428 6646
rect 16552 670 16586 6646
rect 16710 670 16744 6646
rect 16868 670 16902 6646
rect 17026 670 17060 6646
rect 17184 670 17218 6646
rect 17342 670 17376 6646
rect 17500 670 17534 6646
rect 17658 670 17692 6646
rect 17816 670 17850 6646
rect 17974 670 18008 6646
rect 18132 670 18166 6646
rect 18290 670 18324 6646
rect 18448 670 18482 6646
rect 18606 670 18640 6646
rect 18764 670 18798 6646
rect 18922 670 18956 6646
rect 20482 670 20516 6646
rect 20640 670 20674 6646
rect 20798 670 20832 6646
rect 20956 670 20990 6646
rect 21114 670 21148 6646
rect 21272 670 21306 6646
rect 21430 670 21464 6646
rect 21588 670 21622 6646
rect 21746 670 21780 6646
rect 21904 670 21938 6646
rect 22062 670 22096 6646
rect 22220 670 22254 6646
rect 22378 670 22412 6646
rect 22536 670 22570 6646
rect 22694 670 22728 6646
rect 22852 670 22886 6646
rect 23010 670 23044 6646
rect 23168 670 23202 6646
rect 23326 670 23360 6646
rect 23484 670 23518 6646
rect 23642 670 23676 6646
rect 23800 670 23834 6646
rect 23958 670 23992 6646
rect 24116 670 24150 6646
rect 24274 670 24308 6646
rect 24432 670 24466 6646
rect 24590 670 24624 6646
rect 24748 670 24782 6646
rect 24906 670 24940 6646
rect 25064 670 25098 6646
rect 25222 670 25256 6646
rect 1582 -6930 1616 -954
rect 1740 -6930 1774 -954
rect 1898 -6930 1932 -954
rect 2056 -6930 2090 -954
rect 2214 -6930 2248 -954
rect 2372 -6930 2406 -954
rect 2530 -6930 2564 -954
rect 2688 -6930 2722 -954
rect 2846 -6930 2880 -954
rect 3004 -6930 3038 -954
rect 3162 -6930 3196 -954
rect 3320 -6930 3354 -954
rect 3478 -6930 3512 -954
rect 3636 -6930 3670 -954
rect 3794 -6930 3828 -954
rect 3952 -6930 3986 -954
rect 4110 -6930 4144 -954
rect 4268 -6930 4302 -954
rect 4426 -6930 4460 -954
rect 4584 -6930 4618 -954
rect 4742 -6930 4776 -954
rect 4900 -6930 4934 -954
rect 5058 -6930 5092 -954
rect 5216 -6930 5250 -954
rect 5374 -6930 5408 -954
rect 5532 -6930 5566 -954
rect 5690 -6930 5724 -954
rect 5848 -6930 5882 -954
rect 6006 -6930 6040 -954
rect 6164 -6930 6198 -954
rect 6322 -6930 6356 -954
rect 7882 -6930 7916 -954
rect 8040 -6930 8074 -954
rect 8198 -6930 8232 -954
rect 8356 -6930 8390 -954
rect 8514 -6930 8548 -954
rect 8672 -6930 8706 -954
rect 8830 -6930 8864 -954
rect 8988 -6930 9022 -954
rect 9146 -6930 9180 -954
rect 9304 -6930 9338 -954
rect 9462 -6930 9496 -954
rect 9620 -6930 9654 -954
rect 9778 -6930 9812 -954
rect 9936 -6930 9970 -954
rect 10094 -6930 10128 -954
rect 10252 -6930 10286 -954
rect 10410 -6930 10444 -954
rect 10568 -6930 10602 -954
rect 10726 -6930 10760 -954
rect 10884 -6930 10918 -954
rect 11042 -6930 11076 -954
rect 11200 -6930 11234 -954
rect 11358 -6930 11392 -954
rect 11516 -6930 11550 -954
rect 11674 -6930 11708 -954
rect 11832 -6930 11866 -954
rect 11990 -6930 12024 -954
rect 12148 -6930 12182 -954
rect 12306 -6930 12340 -954
rect 12464 -6930 12498 -954
rect 12622 -6930 12656 -954
rect 14182 -6930 14216 -954
rect 14340 -6930 14374 -954
rect 14498 -6930 14532 -954
rect 14656 -6930 14690 -954
rect 14814 -6930 14848 -954
rect 14972 -6930 15006 -954
rect 15130 -6930 15164 -954
rect 15288 -6930 15322 -954
rect 15446 -6930 15480 -954
rect 15604 -6930 15638 -954
rect 15762 -6930 15796 -954
rect 15920 -6930 15954 -954
rect 16078 -6930 16112 -954
rect 16236 -6930 16270 -954
rect 16394 -6930 16428 -954
rect 16552 -6930 16586 -954
rect 16710 -6930 16744 -954
rect 16868 -6930 16902 -954
rect 17026 -6930 17060 -954
rect 17184 -6930 17218 -954
rect 17342 -6930 17376 -954
rect 17500 -6930 17534 -954
rect 17658 -6930 17692 -954
rect 17816 -6930 17850 -954
rect 17974 -6930 18008 -954
rect 18132 -6930 18166 -954
rect 18290 -6930 18324 -954
rect 18448 -6930 18482 -954
rect 18606 -6930 18640 -954
rect 18764 -6930 18798 -954
rect 18922 -6930 18956 -954
rect 20482 -6930 20516 -954
rect 20640 -6930 20674 -954
rect 20798 -6930 20832 -954
rect 20956 -6930 20990 -954
rect 21114 -6930 21148 -954
rect 21272 -6930 21306 -954
rect 21430 -6930 21464 -954
rect 21588 -6930 21622 -954
rect 21746 -6930 21780 -954
rect 21904 -6930 21938 -954
rect 22062 -6930 22096 -954
rect 22220 -6930 22254 -954
rect 22378 -6930 22412 -954
rect 22536 -6930 22570 -954
rect 22694 -6930 22728 -954
rect 22852 -6930 22886 -954
rect 23010 -6930 23044 -954
rect 23168 -6930 23202 -954
rect 23326 -6930 23360 -954
rect 23484 -6930 23518 -954
rect 23642 -6930 23676 -954
rect 23800 -6930 23834 -954
rect 23958 -6930 23992 -954
rect 24116 -6930 24150 -954
rect 24274 -6930 24308 -954
rect 24432 -6930 24466 -954
rect 24590 -6930 24624 -954
rect 24748 -6930 24782 -954
rect 24906 -6930 24940 -954
rect 25064 -6930 25098 -954
rect 25222 -6930 25256 -954
<< mvpsubdiff >>
rect 1436 6868 6502 6880
rect 1436 6834 1544 6868
rect 6394 6834 6502 6868
rect 1436 6822 6502 6834
rect 1436 6772 1494 6822
rect 1436 544 1448 6772
rect 1482 544 1494 6772
rect 6444 6772 6502 6822
rect 1436 494 1494 544
rect 6444 544 6456 6772
rect 6490 544 6502 6772
rect 6444 494 6502 544
rect 1436 482 6502 494
rect 1436 448 1544 482
rect 6394 448 6502 482
rect 1436 436 6502 448
rect 7736 6868 12802 6880
rect 7736 6834 7844 6868
rect 12694 6834 12802 6868
rect 7736 6822 12802 6834
rect 7736 6772 7794 6822
rect 7736 544 7748 6772
rect 7782 544 7794 6772
rect 12744 6772 12802 6822
rect 7736 494 7794 544
rect 12744 544 12756 6772
rect 12790 544 12802 6772
rect 12744 494 12802 544
rect 7736 482 12802 494
rect 7736 448 7844 482
rect 12694 448 12802 482
rect 7736 436 12802 448
rect 14036 6868 19102 6880
rect 14036 6834 14144 6868
rect 18994 6834 19102 6868
rect 14036 6822 19102 6834
rect 14036 6772 14094 6822
rect 14036 544 14048 6772
rect 14082 544 14094 6772
rect 19044 6772 19102 6822
rect 14036 494 14094 544
rect 19044 544 19056 6772
rect 19090 544 19102 6772
rect 19044 494 19102 544
rect 14036 482 19102 494
rect 14036 448 14144 482
rect 18994 448 19102 482
rect 14036 436 19102 448
rect 20336 6868 25402 6880
rect 20336 6834 20444 6868
rect 25294 6834 25402 6868
rect 20336 6822 25402 6834
rect 20336 6772 20394 6822
rect 20336 544 20348 6772
rect 20382 544 20394 6772
rect 25344 6772 25402 6822
rect 20336 494 20394 544
rect 25344 544 25356 6772
rect 25390 544 25402 6772
rect 25344 494 25402 544
rect 20336 482 25402 494
rect 20336 448 20444 482
rect 25294 448 25402 482
rect 20336 436 25402 448
rect 1436 -732 6502 -720
rect 1436 -766 1544 -732
rect 6394 -766 6502 -732
rect 1436 -778 6502 -766
rect 1436 -828 1494 -778
rect 1436 -7056 1448 -828
rect 1482 -7056 1494 -828
rect 6444 -828 6502 -778
rect 1436 -7106 1494 -7056
rect 6444 -7056 6456 -828
rect 6490 -7056 6502 -828
rect 6444 -7106 6502 -7056
rect 1436 -7118 6502 -7106
rect 1436 -7152 1544 -7118
rect 6394 -7152 6502 -7118
rect 1436 -7164 6502 -7152
rect 7736 -732 12802 -720
rect 7736 -766 7844 -732
rect 12694 -766 12802 -732
rect 7736 -778 12802 -766
rect 7736 -828 7794 -778
rect 7736 -7056 7748 -828
rect 7782 -7056 7794 -828
rect 12744 -828 12802 -778
rect 7736 -7106 7794 -7056
rect 12744 -7056 12756 -828
rect 12790 -7056 12802 -828
rect 12744 -7106 12802 -7056
rect 7736 -7118 12802 -7106
rect 7736 -7152 7844 -7118
rect 12694 -7152 12802 -7118
rect 7736 -7164 12802 -7152
rect 14036 -732 19102 -720
rect 14036 -766 14144 -732
rect 18994 -766 19102 -732
rect 14036 -778 19102 -766
rect 14036 -828 14094 -778
rect 14036 -7056 14048 -828
rect 14082 -7056 14094 -828
rect 19044 -828 19102 -778
rect 14036 -7106 14094 -7056
rect 19044 -7056 19056 -828
rect 19090 -7056 19102 -828
rect 19044 -7106 19102 -7056
rect 14036 -7118 19102 -7106
rect 14036 -7152 14144 -7118
rect 18994 -7152 19102 -7118
rect 14036 -7164 19102 -7152
rect 20336 -732 25402 -720
rect 20336 -766 20444 -732
rect 25294 -766 25402 -732
rect 20336 -778 25402 -766
rect 20336 -828 20394 -778
rect 20336 -7056 20348 -828
rect 20382 -7056 20394 -828
rect 25344 -828 25402 -778
rect 20336 -7106 20394 -7056
rect 25344 -7056 25356 -828
rect 25390 -7056 25402 -828
rect 25344 -7106 25402 -7056
rect 20336 -7118 25402 -7106
rect 20336 -7152 20444 -7118
rect 25294 -7152 25402 -7118
rect 20336 -7164 25402 -7152
<< mvpsubdiffcont >>
rect 1544 6834 6394 6868
rect 1448 544 1482 6772
rect 6456 544 6490 6772
rect 1544 448 6394 482
rect 7844 6834 12694 6868
rect 7748 544 7782 6772
rect 12756 544 12790 6772
rect 7844 448 12694 482
rect 14144 6834 18994 6868
rect 14048 544 14082 6772
rect 19056 544 19090 6772
rect 14144 448 18994 482
rect 20444 6834 25294 6868
rect 20348 544 20382 6772
rect 25356 544 25390 6772
rect 20444 448 25294 482
rect 1544 -766 6394 -732
rect 1448 -7056 1482 -828
rect 6456 -7056 6490 -828
rect 1544 -7152 6394 -7118
rect 7844 -766 12694 -732
rect 7748 -7056 7782 -828
rect 12756 -7056 12790 -828
rect 7844 -7152 12694 -7118
rect 14144 -766 18994 -732
rect 14048 -7056 14082 -828
rect 19056 -7056 19090 -828
rect 14144 -7152 18994 -7118
rect 20444 -766 25294 -732
rect 20348 -7056 20382 -828
rect 25356 -7056 25390 -828
rect 20444 -7152 25294 -7118
<< poly >>
rect 1628 6730 1728 6746
rect 1628 6696 1644 6730
rect 1712 6696 1728 6730
rect 1628 6658 1728 6696
rect 1786 6730 1886 6746
rect 1786 6696 1802 6730
rect 1870 6696 1886 6730
rect 1786 6658 1886 6696
rect 1944 6730 2044 6746
rect 1944 6696 1960 6730
rect 2028 6696 2044 6730
rect 1944 6658 2044 6696
rect 2102 6730 2202 6746
rect 2102 6696 2118 6730
rect 2186 6696 2202 6730
rect 2102 6658 2202 6696
rect 2260 6730 2360 6746
rect 2260 6696 2276 6730
rect 2344 6696 2360 6730
rect 2260 6658 2360 6696
rect 2418 6730 2518 6746
rect 2418 6696 2434 6730
rect 2502 6696 2518 6730
rect 2418 6658 2518 6696
rect 2576 6730 2676 6746
rect 2576 6696 2592 6730
rect 2660 6696 2676 6730
rect 2576 6658 2676 6696
rect 2734 6730 2834 6746
rect 2734 6696 2750 6730
rect 2818 6696 2834 6730
rect 2734 6658 2834 6696
rect 2892 6730 2992 6746
rect 2892 6696 2908 6730
rect 2976 6696 2992 6730
rect 2892 6658 2992 6696
rect 3050 6730 3150 6746
rect 3050 6696 3066 6730
rect 3134 6696 3150 6730
rect 3050 6658 3150 6696
rect 3208 6730 3308 6746
rect 3208 6696 3224 6730
rect 3292 6696 3308 6730
rect 3208 6658 3308 6696
rect 3366 6730 3466 6746
rect 3366 6696 3382 6730
rect 3450 6696 3466 6730
rect 3366 6658 3466 6696
rect 3524 6730 3624 6746
rect 3524 6696 3540 6730
rect 3608 6696 3624 6730
rect 3524 6658 3624 6696
rect 3682 6730 3782 6746
rect 3682 6696 3698 6730
rect 3766 6696 3782 6730
rect 3682 6658 3782 6696
rect 3840 6730 3940 6746
rect 3840 6696 3856 6730
rect 3924 6696 3940 6730
rect 3840 6658 3940 6696
rect 3998 6730 4098 6746
rect 3998 6696 4014 6730
rect 4082 6696 4098 6730
rect 3998 6658 4098 6696
rect 4156 6730 4256 6746
rect 4156 6696 4172 6730
rect 4240 6696 4256 6730
rect 4156 6658 4256 6696
rect 4314 6730 4414 6746
rect 4314 6696 4330 6730
rect 4398 6696 4414 6730
rect 4314 6658 4414 6696
rect 4472 6730 4572 6746
rect 4472 6696 4488 6730
rect 4556 6696 4572 6730
rect 4472 6658 4572 6696
rect 4630 6730 4730 6746
rect 4630 6696 4646 6730
rect 4714 6696 4730 6730
rect 4630 6658 4730 6696
rect 4788 6730 4888 6746
rect 4788 6696 4804 6730
rect 4872 6696 4888 6730
rect 4788 6658 4888 6696
rect 4946 6730 5046 6746
rect 4946 6696 4962 6730
rect 5030 6696 5046 6730
rect 4946 6658 5046 6696
rect 5104 6730 5204 6746
rect 5104 6696 5120 6730
rect 5188 6696 5204 6730
rect 5104 6658 5204 6696
rect 5262 6730 5362 6746
rect 5262 6696 5278 6730
rect 5346 6696 5362 6730
rect 5262 6658 5362 6696
rect 5420 6730 5520 6746
rect 5420 6696 5436 6730
rect 5504 6696 5520 6730
rect 5420 6658 5520 6696
rect 5578 6730 5678 6746
rect 5578 6696 5594 6730
rect 5662 6696 5678 6730
rect 5578 6658 5678 6696
rect 5736 6730 5836 6746
rect 5736 6696 5752 6730
rect 5820 6696 5836 6730
rect 5736 6658 5836 6696
rect 5894 6730 5994 6746
rect 5894 6696 5910 6730
rect 5978 6696 5994 6730
rect 5894 6658 5994 6696
rect 6052 6730 6152 6746
rect 6052 6696 6068 6730
rect 6136 6696 6152 6730
rect 6052 6658 6152 6696
rect 6210 6730 6310 6746
rect 6210 6696 6226 6730
rect 6294 6696 6310 6730
rect 6210 6658 6310 6696
rect 1628 620 1728 658
rect 1628 586 1644 620
rect 1712 586 1728 620
rect 1628 570 1728 586
rect 1786 620 1886 658
rect 1786 586 1802 620
rect 1870 586 1886 620
rect 1786 570 1886 586
rect 1944 620 2044 658
rect 1944 586 1960 620
rect 2028 586 2044 620
rect 1944 570 2044 586
rect 2102 620 2202 658
rect 2102 586 2118 620
rect 2186 586 2202 620
rect 2102 570 2202 586
rect 2260 620 2360 658
rect 2260 586 2276 620
rect 2344 586 2360 620
rect 2260 570 2360 586
rect 2418 620 2518 658
rect 2418 586 2434 620
rect 2502 586 2518 620
rect 2418 570 2518 586
rect 2576 620 2676 658
rect 2576 586 2592 620
rect 2660 586 2676 620
rect 2576 570 2676 586
rect 2734 620 2834 658
rect 2734 586 2750 620
rect 2818 586 2834 620
rect 2734 570 2834 586
rect 2892 620 2992 658
rect 2892 586 2908 620
rect 2976 586 2992 620
rect 2892 570 2992 586
rect 3050 620 3150 658
rect 3050 586 3066 620
rect 3134 586 3150 620
rect 3050 570 3150 586
rect 3208 620 3308 658
rect 3208 586 3224 620
rect 3292 586 3308 620
rect 3208 570 3308 586
rect 3366 620 3466 658
rect 3366 586 3382 620
rect 3450 586 3466 620
rect 3366 570 3466 586
rect 3524 620 3624 658
rect 3524 586 3540 620
rect 3608 586 3624 620
rect 3524 570 3624 586
rect 3682 620 3782 658
rect 3682 586 3698 620
rect 3766 586 3782 620
rect 3682 570 3782 586
rect 3840 620 3940 658
rect 3840 586 3856 620
rect 3924 586 3940 620
rect 3840 570 3940 586
rect 3998 620 4098 658
rect 3998 586 4014 620
rect 4082 586 4098 620
rect 3998 570 4098 586
rect 4156 620 4256 658
rect 4156 586 4172 620
rect 4240 586 4256 620
rect 4156 570 4256 586
rect 4314 620 4414 658
rect 4314 586 4330 620
rect 4398 586 4414 620
rect 4314 570 4414 586
rect 4472 620 4572 658
rect 4472 586 4488 620
rect 4556 586 4572 620
rect 4472 570 4572 586
rect 4630 620 4730 658
rect 4630 586 4646 620
rect 4714 586 4730 620
rect 4630 570 4730 586
rect 4788 620 4888 658
rect 4788 586 4804 620
rect 4872 586 4888 620
rect 4788 570 4888 586
rect 4946 620 5046 658
rect 4946 586 4962 620
rect 5030 586 5046 620
rect 4946 570 5046 586
rect 5104 620 5204 658
rect 5104 586 5120 620
rect 5188 586 5204 620
rect 5104 570 5204 586
rect 5262 620 5362 658
rect 5262 586 5278 620
rect 5346 586 5362 620
rect 5262 570 5362 586
rect 5420 620 5520 658
rect 5420 586 5436 620
rect 5504 586 5520 620
rect 5420 570 5520 586
rect 5578 620 5678 658
rect 5578 586 5594 620
rect 5662 586 5678 620
rect 5578 570 5678 586
rect 5736 620 5836 658
rect 5736 586 5752 620
rect 5820 586 5836 620
rect 5736 570 5836 586
rect 5894 620 5994 658
rect 5894 586 5910 620
rect 5978 586 5994 620
rect 5894 570 5994 586
rect 6052 620 6152 658
rect 6052 586 6068 620
rect 6136 586 6152 620
rect 6052 570 6152 586
rect 6210 620 6310 658
rect 6210 586 6226 620
rect 6294 586 6310 620
rect 6210 570 6310 586
rect 7928 6730 8028 6746
rect 7928 6696 7944 6730
rect 8012 6696 8028 6730
rect 7928 6658 8028 6696
rect 8086 6730 8186 6746
rect 8086 6696 8102 6730
rect 8170 6696 8186 6730
rect 8086 6658 8186 6696
rect 8244 6730 8344 6746
rect 8244 6696 8260 6730
rect 8328 6696 8344 6730
rect 8244 6658 8344 6696
rect 8402 6730 8502 6746
rect 8402 6696 8418 6730
rect 8486 6696 8502 6730
rect 8402 6658 8502 6696
rect 8560 6730 8660 6746
rect 8560 6696 8576 6730
rect 8644 6696 8660 6730
rect 8560 6658 8660 6696
rect 8718 6730 8818 6746
rect 8718 6696 8734 6730
rect 8802 6696 8818 6730
rect 8718 6658 8818 6696
rect 8876 6730 8976 6746
rect 8876 6696 8892 6730
rect 8960 6696 8976 6730
rect 8876 6658 8976 6696
rect 9034 6730 9134 6746
rect 9034 6696 9050 6730
rect 9118 6696 9134 6730
rect 9034 6658 9134 6696
rect 9192 6730 9292 6746
rect 9192 6696 9208 6730
rect 9276 6696 9292 6730
rect 9192 6658 9292 6696
rect 9350 6730 9450 6746
rect 9350 6696 9366 6730
rect 9434 6696 9450 6730
rect 9350 6658 9450 6696
rect 9508 6730 9608 6746
rect 9508 6696 9524 6730
rect 9592 6696 9608 6730
rect 9508 6658 9608 6696
rect 9666 6730 9766 6746
rect 9666 6696 9682 6730
rect 9750 6696 9766 6730
rect 9666 6658 9766 6696
rect 9824 6730 9924 6746
rect 9824 6696 9840 6730
rect 9908 6696 9924 6730
rect 9824 6658 9924 6696
rect 9982 6730 10082 6746
rect 9982 6696 9998 6730
rect 10066 6696 10082 6730
rect 9982 6658 10082 6696
rect 10140 6730 10240 6746
rect 10140 6696 10156 6730
rect 10224 6696 10240 6730
rect 10140 6658 10240 6696
rect 10298 6730 10398 6746
rect 10298 6696 10314 6730
rect 10382 6696 10398 6730
rect 10298 6658 10398 6696
rect 10456 6730 10556 6746
rect 10456 6696 10472 6730
rect 10540 6696 10556 6730
rect 10456 6658 10556 6696
rect 10614 6730 10714 6746
rect 10614 6696 10630 6730
rect 10698 6696 10714 6730
rect 10614 6658 10714 6696
rect 10772 6730 10872 6746
rect 10772 6696 10788 6730
rect 10856 6696 10872 6730
rect 10772 6658 10872 6696
rect 10930 6730 11030 6746
rect 10930 6696 10946 6730
rect 11014 6696 11030 6730
rect 10930 6658 11030 6696
rect 11088 6730 11188 6746
rect 11088 6696 11104 6730
rect 11172 6696 11188 6730
rect 11088 6658 11188 6696
rect 11246 6730 11346 6746
rect 11246 6696 11262 6730
rect 11330 6696 11346 6730
rect 11246 6658 11346 6696
rect 11404 6730 11504 6746
rect 11404 6696 11420 6730
rect 11488 6696 11504 6730
rect 11404 6658 11504 6696
rect 11562 6730 11662 6746
rect 11562 6696 11578 6730
rect 11646 6696 11662 6730
rect 11562 6658 11662 6696
rect 11720 6730 11820 6746
rect 11720 6696 11736 6730
rect 11804 6696 11820 6730
rect 11720 6658 11820 6696
rect 11878 6730 11978 6746
rect 11878 6696 11894 6730
rect 11962 6696 11978 6730
rect 11878 6658 11978 6696
rect 12036 6730 12136 6746
rect 12036 6696 12052 6730
rect 12120 6696 12136 6730
rect 12036 6658 12136 6696
rect 12194 6730 12294 6746
rect 12194 6696 12210 6730
rect 12278 6696 12294 6730
rect 12194 6658 12294 6696
rect 12352 6730 12452 6746
rect 12352 6696 12368 6730
rect 12436 6696 12452 6730
rect 12352 6658 12452 6696
rect 12510 6730 12610 6746
rect 12510 6696 12526 6730
rect 12594 6696 12610 6730
rect 12510 6658 12610 6696
rect 7928 620 8028 658
rect 7928 586 7944 620
rect 8012 586 8028 620
rect 7928 570 8028 586
rect 8086 620 8186 658
rect 8086 586 8102 620
rect 8170 586 8186 620
rect 8086 570 8186 586
rect 8244 620 8344 658
rect 8244 586 8260 620
rect 8328 586 8344 620
rect 8244 570 8344 586
rect 8402 620 8502 658
rect 8402 586 8418 620
rect 8486 586 8502 620
rect 8402 570 8502 586
rect 8560 620 8660 658
rect 8560 586 8576 620
rect 8644 586 8660 620
rect 8560 570 8660 586
rect 8718 620 8818 658
rect 8718 586 8734 620
rect 8802 586 8818 620
rect 8718 570 8818 586
rect 8876 620 8976 658
rect 8876 586 8892 620
rect 8960 586 8976 620
rect 8876 570 8976 586
rect 9034 620 9134 658
rect 9034 586 9050 620
rect 9118 586 9134 620
rect 9034 570 9134 586
rect 9192 620 9292 658
rect 9192 586 9208 620
rect 9276 586 9292 620
rect 9192 570 9292 586
rect 9350 620 9450 658
rect 9350 586 9366 620
rect 9434 586 9450 620
rect 9350 570 9450 586
rect 9508 620 9608 658
rect 9508 586 9524 620
rect 9592 586 9608 620
rect 9508 570 9608 586
rect 9666 620 9766 658
rect 9666 586 9682 620
rect 9750 586 9766 620
rect 9666 570 9766 586
rect 9824 620 9924 658
rect 9824 586 9840 620
rect 9908 586 9924 620
rect 9824 570 9924 586
rect 9982 620 10082 658
rect 9982 586 9998 620
rect 10066 586 10082 620
rect 9982 570 10082 586
rect 10140 620 10240 658
rect 10140 586 10156 620
rect 10224 586 10240 620
rect 10140 570 10240 586
rect 10298 620 10398 658
rect 10298 586 10314 620
rect 10382 586 10398 620
rect 10298 570 10398 586
rect 10456 620 10556 658
rect 10456 586 10472 620
rect 10540 586 10556 620
rect 10456 570 10556 586
rect 10614 620 10714 658
rect 10614 586 10630 620
rect 10698 586 10714 620
rect 10614 570 10714 586
rect 10772 620 10872 658
rect 10772 586 10788 620
rect 10856 586 10872 620
rect 10772 570 10872 586
rect 10930 620 11030 658
rect 10930 586 10946 620
rect 11014 586 11030 620
rect 10930 570 11030 586
rect 11088 620 11188 658
rect 11088 586 11104 620
rect 11172 586 11188 620
rect 11088 570 11188 586
rect 11246 620 11346 658
rect 11246 586 11262 620
rect 11330 586 11346 620
rect 11246 570 11346 586
rect 11404 620 11504 658
rect 11404 586 11420 620
rect 11488 586 11504 620
rect 11404 570 11504 586
rect 11562 620 11662 658
rect 11562 586 11578 620
rect 11646 586 11662 620
rect 11562 570 11662 586
rect 11720 620 11820 658
rect 11720 586 11736 620
rect 11804 586 11820 620
rect 11720 570 11820 586
rect 11878 620 11978 658
rect 11878 586 11894 620
rect 11962 586 11978 620
rect 11878 570 11978 586
rect 12036 620 12136 658
rect 12036 586 12052 620
rect 12120 586 12136 620
rect 12036 570 12136 586
rect 12194 620 12294 658
rect 12194 586 12210 620
rect 12278 586 12294 620
rect 12194 570 12294 586
rect 12352 620 12452 658
rect 12352 586 12368 620
rect 12436 586 12452 620
rect 12352 570 12452 586
rect 12510 620 12610 658
rect 12510 586 12526 620
rect 12594 586 12610 620
rect 12510 570 12610 586
rect 14228 6730 14328 6746
rect 14228 6696 14244 6730
rect 14312 6696 14328 6730
rect 14228 6658 14328 6696
rect 14386 6730 14486 6746
rect 14386 6696 14402 6730
rect 14470 6696 14486 6730
rect 14386 6658 14486 6696
rect 14544 6730 14644 6746
rect 14544 6696 14560 6730
rect 14628 6696 14644 6730
rect 14544 6658 14644 6696
rect 14702 6730 14802 6746
rect 14702 6696 14718 6730
rect 14786 6696 14802 6730
rect 14702 6658 14802 6696
rect 14860 6730 14960 6746
rect 14860 6696 14876 6730
rect 14944 6696 14960 6730
rect 14860 6658 14960 6696
rect 15018 6730 15118 6746
rect 15018 6696 15034 6730
rect 15102 6696 15118 6730
rect 15018 6658 15118 6696
rect 15176 6730 15276 6746
rect 15176 6696 15192 6730
rect 15260 6696 15276 6730
rect 15176 6658 15276 6696
rect 15334 6730 15434 6746
rect 15334 6696 15350 6730
rect 15418 6696 15434 6730
rect 15334 6658 15434 6696
rect 15492 6730 15592 6746
rect 15492 6696 15508 6730
rect 15576 6696 15592 6730
rect 15492 6658 15592 6696
rect 15650 6730 15750 6746
rect 15650 6696 15666 6730
rect 15734 6696 15750 6730
rect 15650 6658 15750 6696
rect 15808 6730 15908 6746
rect 15808 6696 15824 6730
rect 15892 6696 15908 6730
rect 15808 6658 15908 6696
rect 15966 6730 16066 6746
rect 15966 6696 15982 6730
rect 16050 6696 16066 6730
rect 15966 6658 16066 6696
rect 16124 6730 16224 6746
rect 16124 6696 16140 6730
rect 16208 6696 16224 6730
rect 16124 6658 16224 6696
rect 16282 6730 16382 6746
rect 16282 6696 16298 6730
rect 16366 6696 16382 6730
rect 16282 6658 16382 6696
rect 16440 6730 16540 6746
rect 16440 6696 16456 6730
rect 16524 6696 16540 6730
rect 16440 6658 16540 6696
rect 16598 6730 16698 6746
rect 16598 6696 16614 6730
rect 16682 6696 16698 6730
rect 16598 6658 16698 6696
rect 16756 6730 16856 6746
rect 16756 6696 16772 6730
rect 16840 6696 16856 6730
rect 16756 6658 16856 6696
rect 16914 6730 17014 6746
rect 16914 6696 16930 6730
rect 16998 6696 17014 6730
rect 16914 6658 17014 6696
rect 17072 6730 17172 6746
rect 17072 6696 17088 6730
rect 17156 6696 17172 6730
rect 17072 6658 17172 6696
rect 17230 6730 17330 6746
rect 17230 6696 17246 6730
rect 17314 6696 17330 6730
rect 17230 6658 17330 6696
rect 17388 6730 17488 6746
rect 17388 6696 17404 6730
rect 17472 6696 17488 6730
rect 17388 6658 17488 6696
rect 17546 6730 17646 6746
rect 17546 6696 17562 6730
rect 17630 6696 17646 6730
rect 17546 6658 17646 6696
rect 17704 6730 17804 6746
rect 17704 6696 17720 6730
rect 17788 6696 17804 6730
rect 17704 6658 17804 6696
rect 17862 6730 17962 6746
rect 17862 6696 17878 6730
rect 17946 6696 17962 6730
rect 17862 6658 17962 6696
rect 18020 6730 18120 6746
rect 18020 6696 18036 6730
rect 18104 6696 18120 6730
rect 18020 6658 18120 6696
rect 18178 6730 18278 6746
rect 18178 6696 18194 6730
rect 18262 6696 18278 6730
rect 18178 6658 18278 6696
rect 18336 6730 18436 6746
rect 18336 6696 18352 6730
rect 18420 6696 18436 6730
rect 18336 6658 18436 6696
rect 18494 6730 18594 6746
rect 18494 6696 18510 6730
rect 18578 6696 18594 6730
rect 18494 6658 18594 6696
rect 18652 6730 18752 6746
rect 18652 6696 18668 6730
rect 18736 6696 18752 6730
rect 18652 6658 18752 6696
rect 18810 6730 18910 6746
rect 18810 6696 18826 6730
rect 18894 6696 18910 6730
rect 18810 6658 18910 6696
rect 14228 620 14328 658
rect 14228 586 14244 620
rect 14312 586 14328 620
rect 14228 570 14328 586
rect 14386 620 14486 658
rect 14386 586 14402 620
rect 14470 586 14486 620
rect 14386 570 14486 586
rect 14544 620 14644 658
rect 14544 586 14560 620
rect 14628 586 14644 620
rect 14544 570 14644 586
rect 14702 620 14802 658
rect 14702 586 14718 620
rect 14786 586 14802 620
rect 14702 570 14802 586
rect 14860 620 14960 658
rect 14860 586 14876 620
rect 14944 586 14960 620
rect 14860 570 14960 586
rect 15018 620 15118 658
rect 15018 586 15034 620
rect 15102 586 15118 620
rect 15018 570 15118 586
rect 15176 620 15276 658
rect 15176 586 15192 620
rect 15260 586 15276 620
rect 15176 570 15276 586
rect 15334 620 15434 658
rect 15334 586 15350 620
rect 15418 586 15434 620
rect 15334 570 15434 586
rect 15492 620 15592 658
rect 15492 586 15508 620
rect 15576 586 15592 620
rect 15492 570 15592 586
rect 15650 620 15750 658
rect 15650 586 15666 620
rect 15734 586 15750 620
rect 15650 570 15750 586
rect 15808 620 15908 658
rect 15808 586 15824 620
rect 15892 586 15908 620
rect 15808 570 15908 586
rect 15966 620 16066 658
rect 15966 586 15982 620
rect 16050 586 16066 620
rect 15966 570 16066 586
rect 16124 620 16224 658
rect 16124 586 16140 620
rect 16208 586 16224 620
rect 16124 570 16224 586
rect 16282 620 16382 658
rect 16282 586 16298 620
rect 16366 586 16382 620
rect 16282 570 16382 586
rect 16440 620 16540 658
rect 16440 586 16456 620
rect 16524 586 16540 620
rect 16440 570 16540 586
rect 16598 620 16698 658
rect 16598 586 16614 620
rect 16682 586 16698 620
rect 16598 570 16698 586
rect 16756 620 16856 658
rect 16756 586 16772 620
rect 16840 586 16856 620
rect 16756 570 16856 586
rect 16914 620 17014 658
rect 16914 586 16930 620
rect 16998 586 17014 620
rect 16914 570 17014 586
rect 17072 620 17172 658
rect 17072 586 17088 620
rect 17156 586 17172 620
rect 17072 570 17172 586
rect 17230 620 17330 658
rect 17230 586 17246 620
rect 17314 586 17330 620
rect 17230 570 17330 586
rect 17388 620 17488 658
rect 17388 586 17404 620
rect 17472 586 17488 620
rect 17388 570 17488 586
rect 17546 620 17646 658
rect 17546 586 17562 620
rect 17630 586 17646 620
rect 17546 570 17646 586
rect 17704 620 17804 658
rect 17704 586 17720 620
rect 17788 586 17804 620
rect 17704 570 17804 586
rect 17862 620 17962 658
rect 17862 586 17878 620
rect 17946 586 17962 620
rect 17862 570 17962 586
rect 18020 620 18120 658
rect 18020 586 18036 620
rect 18104 586 18120 620
rect 18020 570 18120 586
rect 18178 620 18278 658
rect 18178 586 18194 620
rect 18262 586 18278 620
rect 18178 570 18278 586
rect 18336 620 18436 658
rect 18336 586 18352 620
rect 18420 586 18436 620
rect 18336 570 18436 586
rect 18494 620 18594 658
rect 18494 586 18510 620
rect 18578 586 18594 620
rect 18494 570 18594 586
rect 18652 620 18752 658
rect 18652 586 18668 620
rect 18736 586 18752 620
rect 18652 570 18752 586
rect 18810 620 18910 658
rect 18810 586 18826 620
rect 18894 586 18910 620
rect 18810 570 18910 586
rect 20528 6730 20628 6746
rect 20528 6696 20544 6730
rect 20612 6696 20628 6730
rect 20528 6658 20628 6696
rect 20686 6730 20786 6746
rect 20686 6696 20702 6730
rect 20770 6696 20786 6730
rect 20686 6658 20786 6696
rect 20844 6730 20944 6746
rect 20844 6696 20860 6730
rect 20928 6696 20944 6730
rect 20844 6658 20944 6696
rect 21002 6730 21102 6746
rect 21002 6696 21018 6730
rect 21086 6696 21102 6730
rect 21002 6658 21102 6696
rect 21160 6730 21260 6746
rect 21160 6696 21176 6730
rect 21244 6696 21260 6730
rect 21160 6658 21260 6696
rect 21318 6730 21418 6746
rect 21318 6696 21334 6730
rect 21402 6696 21418 6730
rect 21318 6658 21418 6696
rect 21476 6730 21576 6746
rect 21476 6696 21492 6730
rect 21560 6696 21576 6730
rect 21476 6658 21576 6696
rect 21634 6730 21734 6746
rect 21634 6696 21650 6730
rect 21718 6696 21734 6730
rect 21634 6658 21734 6696
rect 21792 6730 21892 6746
rect 21792 6696 21808 6730
rect 21876 6696 21892 6730
rect 21792 6658 21892 6696
rect 21950 6730 22050 6746
rect 21950 6696 21966 6730
rect 22034 6696 22050 6730
rect 21950 6658 22050 6696
rect 22108 6730 22208 6746
rect 22108 6696 22124 6730
rect 22192 6696 22208 6730
rect 22108 6658 22208 6696
rect 22266 6730 22366 6746
rect 22266 6696 22282 6730
rect 22350 6696 22366 6730
rect 22266 6658 22366 6696
rect 22424 6730 22524 6746
rect 22424 6696 22440 6730
rect 22508 6696 22524 6730
rect 22424 6658 22524 6696
rect 22582 6730 22682 6746
rect 22582 6696 22598 6730
rect 22666 6696 22682 6730
rect 22582 6658 22682 6696
rect 22740 6730 22840 6746
rect 22740 6696 22756 6730
rect 22824 6696 22840 6730
rect 22740 6658 22840 6696
rect 22898 6730 22998 6746
rect 22898 6696 22914 6730
rect 22982 6696 22998 6730
rect 22898 6658 22998 6696
rect 23056 6730 23156 6746
rect 23056 6696 23072 6730
rect 23140 6696 23156 6730
rect 23056 6658 23156 6696
rect 23214 6730 23314 6746
rect 23214 6696 23230 6730
rect 23298 6696 23314 6730
rect 23214 6658 23314 6696
rect 23372 6730 23472 6746
rect 23372 6696 23388 6730
rect 23456 6696 23472 6730
rect 23372 6658 23472 6696
rect 23530 6730 23630 6746
rect 23530 6696 23546 6730
rect 23614 6696 23630 6730
rect 23530 6658 23630 6696
rect 23688 6730 23788 6746
rect 23688 6696 23704 6730
rect 23772 6696 23788 6730
rect 23688 6658 23788 6696
rect 23846 6730 23946 6746
rect 23846 6696 23862 6730
rect 23930 6696 23946 6730
rect 23846 6658 23946 6696
rect 24004 6730 24104 6746
rect 24004 6696 24020 6730
rect 24088 6696 24104 6730
rect 24004 6658 24104 6696
rect 24162 6730 24262 6746
rect 24162 6696 24178 6730
rect 24246 6696 24262 6730
rect 24162 6658 24262 6696
rect 24320 6730 24420 6746
rect 24320 6696 24336 6730
rect 24404 6696 24420 6730
rect 24320 6658 24420 6696
rect 24478 6730 24578 6746
rect 24478 6696 24494 6730
rect 24562 6696 24578 6730
rect 24478 6658 24578 6696
rect 24636 6730 24736 6746
rect 24636 6696 24652 6730
rect 24720 6696 24736 6730
rect 24636 6658 24736 6696
rect 24794 6730 24894 6746
rect 24794 6696 24810 6730
rect 24878 6696 24894 6730
rect 24794 6658 24894 6696
rect 24952 6730 25052 6746
rect 24952 6696 24968 6730
rect 25036 6696 25052 6730
rect 24952 6658 25052 6696
rect 25110 6730 25210 6746
rect 25110 6696 25126 6730
rect 25194 6696 25210 6730
rect 25110 6658 25210 6696
rect 20528 620 20628 658
rect 20528 586 20544 620
rect 20612 586 20628 620
rect 20528 570 20628 586
rect 20686 620 20786 658
rect 20686 586 20702 620
rect 20770 586 20786 620
rect 20686 570 20786 586
rect 20844 620 20944 658
rect 20844 586 20860 620
rect 20928 586 20944 620
rect 20844 570 20944 586
rect 21002 620 21102 658
rect 21002 586 21018 620
rect 21086 586 21102 620
rect 21002 570 21102 586
rect 21160 620 21260 658
rect 21160 586 21176 620
rect 21244 586 21260 620
rect 21160 570 21260 586
rect 21318 620 21418 658
rect 21318 586 21334 620
rect 21402 586 21418 620
rect 21318 570 21418 586
rect 21476 620 21576 658
rect 21476 586 21492 620
rect 21560 586 21576 620
rect 21476 570 21576 586
rect 21634 620 21734 658
rect 21634 586 21650 620
rect 21718 586 21734 620
rect 21634 570 21734 586
rect 21792 620 21892 658
rect 21792 586 21808 620
rect 21876 586 21892 620
rect 21792 570 21892 586
rect 21950 620 22050 658
rect 21950 586 21966 620
rect 22034 586 22050 620
rect 21950 570 22050 586
rect 22108 620 22208 658
rect 22108 586 22124 620
rect 22192 586 22208 620
rect 22108 570 22208 586
rect 22266 620 22366 658
rect 22266 586 22282 620
rect 22350 586 22366 620
rect 22266 570 22366 586
rect 22424 620 22524 658
rect 22424 586 22440 620
rect 22508 586 22524 620
rect 22424 570 22524 586
rect 22582 620 22682 658
rect 22582 586 22598 620
rect 22666 586 22682 620
rect 22582 570 22682 586
rect 22740 620 22840 658
rect 22740 586 22756 620
rect 22824 586 22840 620
rect 22740 570 22840 586
rect 22898 620 22998 658
rect 22898 586 22914 620
rect 22982 586 22998 620
rect 22898 570 22998 586
rect 23056 620 23156 658
rect 23056 586 23072 620
rect 23140 586 23156 620
rect 23056 570 23156 586
rect 23214 620 23314 658
rect 23214 586 23230 620
rect 23298 586 23314 620
rect 23214 570 23314 586
rect 23372 620 23472 658
rect 23372 586 23388 620
rect 23456 586 23472 620
rect 23372 570 23472 586
rect 23530 620 23630 658
rect 23530 586 23546 620
rect 23614 586 23630 620
rect 23530 570 23630 586
rect 23688 620 23788 658
rect 23688 586 23704 620
rect 23772 586 23788 620
rect 23688 570 23788 586
rect 23846 620 23946 658
rect 23846 586 23862 620
rect 23930 586 23946 620
rect 23846 570 23946 586
rect 24004 620 24104 658
rect 24004 586 24020 620
rect 24088 586 24104 620
rect 24004 570 24104 586
rect 24162 620 24262 658
rect 24162 586 24178 620
rect 24246 586 24262 620
rect 24162 570 24262 586
rect 24320 620 24420 658
rect 24320 586 24336 620
rect 24404 586 24420 620
rect 24320 570 24420 586
rect 24478 620 24578 658
rect 24478 586 24494 620
rect 24562 586 24578 620
rect 24478 570 24578 586
rect 24636 620 24736 658
rect 24636 586 24652 620
rect 24720 586 24736 620
rect 24636 570 24736 586
rect 24794 620 24894 658
rect 24794 586 24810 620
rect 24878 586 24894 620
rect 24794 570 24894 586
rect 24952 620 25052 658
rect 24952 586 24968 620
rect 25036 586 25052 620
rect 24952 570 25052 586
rect 25110 620 25210 658
rect 25110 586 25126 620
rect 25194 586 25210 620
rect 25110 570 25210 586
rect 1628 -870 1728 -854
rect 1628 -904 1644 -870
rect 1712 -904 1728 -870
rect 1628 -942 1728 -904
rect 1786 -870 1886 -854
rect 1786 -904 1802 -870
rect 1870 -904 1886 -870
rect 1786 -942 1886 -904
rect 1944 -870 2044 -854
rect 1944 -904 1960 -870
rect 2028 -904 2044 -870
rect 1944 -942 2044 -904
rect 2102 -870 2202 -854
rect 2102 -904 2118 -870
rect 2186 -904 2202 -870
rect 2102 -942 2202 -904
rect 2260 -870 2360 -854
rect 2260 -904 2276 -870
rect 2344 -904 2360 -870
rect 2260 -942 2360 -904
rect 2418 -870 2518 -854
rect 2418 -904 2434 -870
rect 2502 -904 2518 -870
rect 2418 -942 2518 -904
rect 2576 -870 2676 -854
rect 2576 -904 2592 -870
rect 2660 -904 2676 -870
rect 2576 -942 2676 -904
rect 2734 -870 2834 -854
rect 2734 -904 2750 -870
rect 2818 -904 2834 -870
rect 2734 -942 2834 -904
rect 2892 -870 2992 -854
rect 2892 -904 2908 -870
rect 2976 -904 2992 -870
rect 2892 -942 2992 -904
rect 3050 -870 3150 -854
rect 3050 -904 3066 -870
rect 3134 -904 3150 -870
rect 3050 -942 3150 -904
rect 3208 -870 3308 -854
rect 3208 -904 3224 -870
rect 3292 -904 3308 -870
rect 3208 -942 3308 -904
rect 3366 -870 3466 -854
rect 3366 -904 3382 -870
rect 3450 -904 3466 -870
rect 3366 -942 3466 -904
rect 3524 -870 3624 -854
rect 3524 -904 3540 -870
rect 3608 -904 3624 -870
rect 3524 -942 3624 -904
rect 3682 -870 3782 -854
rect 3682 -904 3698 -870
rect 3766 -904 3782 -870
rect 3682 -942 3782 -904
rect 3840 -870 3940 -854
rect 3840 -904 3856 -870
rect 3924 -904 3940 -870
rect 3840 -942 3940 -904
rect 3998 -870 4098 -854
rect 3998 -904 4014 -870
rect 4082 -904 4098 -870
rect 3998 -942 4098 -904
rect 4156 -870 4256 -854
rect 4156 -904 4172 -870
rect 4240 -904 4256 -870
rect 4156 -942 4256 -904
rect 4314 -870 4414 -854
rect 4314 -904 4330 -870
rect 4398 -904 4414 -870
rect 4314 -942 4414 -904
rect 4472 -870 4572 -854
rect 4472 -904 4488 -870
rect 4556 -904 4572 -870
rect 4472 -942 4572 -904
rect 4630 -870 4730 -854
rect 4630 -904 4646 -870
rect 4714 -904 4730 -870
rect 4630 -942 4730 -904
rect 4788 -870 4888 -854
rect 4788 -904 4804 -870
rect 4872 -904 4888 -870
rect 4788 -942 4888 -904
rect 4946 -870 5046 -854
rect 4946 -904 4962 -870
rect 5030 -904 5046 -870
rect 4946 -942 5046 -904
rect 5104 -870 5204 -854
rect 5104 -904 5120 -870
rect 5188 -904 5204 -870
rect 5104 -942 5204 -904
rect 5262 -870 5362 -854
rect 5262 -904 5278 -870
rect 5346 -904 5362 -870
rect 5262 -942 5362 -904
rect 5420 -870 5520 -854
rect 5420 -904 5436 -870
rect 5504 -904 5520 -870
rect 5420 -942 5520 -904
rect 5578 -870 5678 -854
rect 5578 -904 5594 -870
rect 5662 -904 5678 -870
rect 5578 -942 5678 -904
rect 5736 -870 5836 -854
rect 5736 -904 5752 -870
rect 5820 -904 5836 -870
rect 5736 -942 5836 -904
rect 5894 -870 5994 -854
rect 5894 -904 5910 -870
rect 5978 -904 5994 -870
rect 5894 -942 5994 -904
rect 6052 -870 6152 -854
rect 6052 -904 6068 -870
rect 6136 -904 6152 -870
rect 6052 -942 6152 -904
rect 6210 -870 6310 -854
rect 6210 -904 6226 -870
rect 6294 -904 6310 -870
rect 6210 -942 6310 -904
rect 1628 -6980 1728 -6942
rect 1628 -7014 1644 -6980
rect 1712 -7014 1728 -6980
rect 1628 -7030 1728 -7014
rect 1786 -6980 1886 -6942
rect 1786 -7014 1802 -6980
rect 1870 -7014 1886 -6980
rect 1786 -7030 1886 -7014
rect 1944 -6980 2044 -6942
rect 1944 -7014 1960 -6980
rect 2028 -7014 2044 -6980
rect 1944 -7030 2044 -7014
rect 2102 -6980 2202 -6942
rect 2102 -7014 2118 -6980
rect 2186 -7014 2202 -6980
rect 2102 -7030 2202 -7014
rect 2260 -6980 2360 -6942
rect 2260 -7014 2276 -6980
rect 2344 -7014 2360 -6980
rect 2260 -7030 2360 -7014
rect 2418 -6980 2518 -6942
rect 2418 -7014 2434 -6980
rect 2502 -7014 2518 -6980
rect 2418 -7030 2518 -7014
rect 2576 -6980 2676 -6942
rect 2576 -7014 2592 -6980
rect 2660 -7014 2676 -6980
rect 2576 -7030 2676 -7014
rect 2734 -6980 2834 -6942
rect 2734 -7014 2750 -6980
rect 2818 -7014 2834 -6980
rect 2734 -7030 2834 -7014
rect 2892 -6980 2992 -6942
rect 2892 -7014 2908 -6980
rect 2976 -7014 2992 -6980
rect 2892 -7030 2992 -7014
rect 3050 -6980 3150 -6942
rect 3050 -7014 3066 -6980
rect 3134 -7014 3150 -6980
rect 3050 -7030 3150 -7014
rect 3208 -6980 3308 -6942
rect 3208 -7014 3224 -6980
rect 3292 -7014 3308 -6980
rect 3208 -7030 3308 -7014
rect 3366 -6980 3466 -6942
rect 3366 -7014 3382 -6980
rect 3450 -7014 3466 -6980
rect 3366 -7030 3466 -7014
rect 3524 -6980 3624 -6942
rect 3524 -7014 3540 -6980
rect 3608 -7014 3624 -6980
rect 3524 -7030 3624 -7014
rect 3682 -6980 3782 -6942
rect 3682 -7014 3698 -6980
rect 3766 -7014 3782 -6980
rect 3682 -7030 3782 -7014
rect 3840 -6980 3940 -6942
rect 3840 -7014 3856 -6980
rect 3924 -7014 3940 -6980
rect 3840 -7030 3940 -7014
rect 3998 -6980 4098 -6942
rect 3998 -7014 4014 -6980
rect 4082 -7014 4098 -6980
rect 3998 -7030 4098 -7014
rect 4156 -6980 4256 -6942
rect 4156 -7014 4172 -6980
rect 4240 -7014 4256 -6980
rect 4156 -7030 4256 -7014
rect 4314 -6980 4414 -6942
rect 4314 -7014 4330 -6980
rect 4398 -7014 4414 -6980
rect 4314 -7030 4414 -7014
rect 4472 -6980 4572 -6942
rect 4472 -7014 4488 -6980
rect 4556 -7014 4572 -6980
rect 4472 -7030 4572 -7014
rect 4630 -6980 4730 -6942
rect 4630 -7014 4646 -6980
rect 4714 -7014 4730 -6980
rect 4630 -7030 4730 -7014
rect 4788 -6980 4888 -6942
rect 4788 -7014 4804 -6980
rect 4872 -7014 4888 -6980
rect 4788 -7030 4888 -7014
rect 4946 -6980 5046 -6942
rect 4946 -7014 4962 -6980
rect 5030 -7014 5046 -6980
rect 4946 -7030 5046 -7014
rect 5104 -6980 5204 -6942
rect 5104 -7014 5120 -6980
rect 5188 -7014 5204 -6980
rect 5104 -7030 5204 -7014
rect 5262 -6980 5362 -6942
rect 5262 -7014 5278 -6980
rect 5346 -7014 5362 -6980
rect 5262 -7030 5362 -7014
rect 5420 -6980 5520 -6942
rect 5420 -7014 5436 -6980
rect 5504 -7014 5520 -6980
rect 5420 -7030 5520 -7014
rect 5578 -6980 5678 -6942
rect 5578 -7014 5594 -6980
rect 5662 -7014 5678 -6980
rect 5578 -7030 5678 -7014
rect 5736 -6980 5836 -6942
rect 5736 -7014 5752 -6980
rect 5820 -7014 5836 -6980
rect 5736 -7030 5836 -7014
rect 5894 -6980 5994 -6942
rect 5894 -7014 5910 -6980
rect 5978 -7014 5994 -6980
rect 5894 -7030 5994 -7014
rect 6052 -6980 6152 -6942
rect 6052 -7014 6068 -6980
rect 6136 -7014 6152 -6980
rect 6052 -7030 6152 -7014
rect 6210 -6980 6310 -6942
rect 6210 -7014 6226 -6980
rect 6294 -7014 6310 -6980
rect 6210 -7030 6310 -7014
rect 7928 -870 8028 -854
rect 7928 -904 7944 -870
rect 8012 -904 8028 -870
rect 7928 -942 8028 -904
rect 8086 -870 8186 -854
rect 8086 -904 8102 -870
rect 8170 -904 8186 -870
rect 8086 -942 8186 -904
rect 8244 -870 8344 -854
rect 8244 -904 8260 -870
rect 8328 -904 8344 -870
rect 8244 -942 8344 -904
rect 8402 -870 8502 -854
rect 8402 -904 8418 -870
rect 8486 -904 8502 -870
rect 8402 -942 8502 -904
rect 8560 -870 8660 -854
rect 8560 -904 8576 -870
rect 8644 -904 8660 -870
rect 8560 -942 8660 -904
rect 8718 -870 8818 -854
rect 8718 -904 8734 -870
rect 8802 -904 8818 -870
rect 8718 -942 8818 -904
rect 8876 -870 8976 -854
rect 8876 -904 8892 -870
rect 8960 -904 8976 -870
rect 8876 -942 8976 -904
rect 9034 -870 9134 -854
rect 9034 -904 9050 -870
rect 9118 -904 9134 -870
rect 9034 -942 9134 -904
rect 9192 -870 9292 -854
rect 9192 -904 9208 -870
rect 9276 -904 9292 -870
rect 9192 -942 9292 -904
rect 9350 -870 9450 -854
rect 9350 -904 9366 -870
rect 9434 -904 9450 -870
rect 9350 -942 9450 -904
rect 9508 -870 9608 -854
rect 9508 -904 9524 -870
rect 9592 -904 9608 -870
rect 9508 -942 9608 -904
rect 9666 -870 9766 -854
rect 9666 -904 9682 -870
rect 9750 -904 9766 -870
rect 9666 -942 9766 -904
rect 9824 -870 9924 -854
rect 9824 -904 9840 -870
rect 9908 -904 9924 -870
rect 9824 -942 9924 -904
rect 9982 -870 10082 -854
rect 9982 -904 9998 -870
rect 10066 -904 10082 -870
rect 9982 -942 10082 -904
rect 10140 -870 10240 -854
rect 10140 -904 10156 -870
rect 10224 -904 10240 -870
rect 10140 -942 10240 -904
rect 10298 -870 10398 -854
rect 10298 -904 10314 -870
rect 10382 -904 10398 -870
rect 10298 -942 10398 -904
rect 10456 -870 10556 -854
rect 10456 -904 10472 -870
rect 10540 -904 10556 -870
rect 10456 -942 10556 -904
rect 10614 -870 10714 -854
rect 10614 -904 10630 -870
rect 10698 -904 10714 -870
rect 10614 -942 10714 -904
rect 10772 -870 10872 -854
rect 10772 -904 10788 -870
rect 10856 -904 10872 -870
rect 10772 -942 10872 -904
rect 10930 -870 11030 -854
rect 10930 -904 10946 -870
rect 11014 -904 11030 -870
rect 10930 -942 11030 -904
rect 11088 -870 11188 -854
rect 11088 -904 11104 -870
rect 11172 -904 11188 -870
rect 11088 -942 11188 -904
rect 11246 -870 11346 -854
rect 11246 -904 11262 -870
rect 11330 -904 11346 -870
rect 11246 -942 11346 -904
rect 11404 -870 11504 -854
rect 11404 -904 11420 -870
rect 11488 -904 11504 -870
rect 11404 -942 11504 -904
rect 11562 -870 11662 -854
rect 11562 -904 11578 -870
rect 11646 -904 11662 -870
rect 11562 -942 11662 -904
rect 11720 -870 11820 -854
rect 11720 -904 11736 -870
rect 11804 -904 11820 -870
rect 11720 -942 11820 -904
rect 11878 -870 11978 -854
rect 11878 -904 11894 -870
rect 11962 -904 11978 -870
rect 11878 -942 11978 -904
rect 12036 -870 12136 -854
rect 12036 -904 12052 -870
rect 12120 -904 12136 -870
rect 12036 -942 12136 -904
rect 12194 -870 12294 -854
rect 12194 -904 12210 -870
rect 12278 -904 12294 -870
rect 12194 -942 12294 -904
rect 12352 -870 12452 -854
rect 12352 -904 12368 -870
rect 12436 -904 12452 -870
rect 12352 -942 12452 -904
rect 12510 -870 12610 -854
rect 12510 -904 12526 -870
rect 12594 -904 12610 -870
rect 12510 -942 12610 -904
rect 7928 -6980 8028 -6942
rect 7928 -7014 7944 -6980
rect 8012 -7014 8028 -6980
rect 7928 -7030 8028 -7014
rect 8086 -6980 8186 -6942
rect 8086 -7014 8102 -6980
rect 8170 -7014 8186 -6980
rect 8086 -7030 8186 -7014
rect 8244 -6980 8344 -6942
rect 8244 -7014 8260 -6980
rect 8328 -7014 8344 -6980
rect 8244 -7030 8344 -7014
rect 8402 -6980 8502 -6942
rect 8402 -7014 8418 -6980
rect 8486 -7014 8502 -6980
rect 8402 -7030 8502 -7014
rect 8560 -6980 8660 -6942
rect 8560 -7014 8576 -6980
rect 8644 -7014 8660 -6980
rect 8560 -7030 8660 -7014
rect 8718 -6980 8818 -6942
rect 8718 -7014 8734 -6980
rect 8802 -7014 8818 -6980
rect 8718 -7030 8818 -7014
rect 8876 -6980 8976 -6942
rect 8876 -7014 8892 -6980
rect 8960 -7014 8976 -6980
rect 8876 -7030 8976 -7014
rect 9034 -6980 9134 -6942
rect 9034 -7014 9050 -6980
rect 9118 -7014 9134 -6980
rect 9034 -7030 9134 -7014
rect 9192 -6980 9292 -6942
rect 9192 -7014 9208 -6980
rect 9276 -7014 9292 -6980
rect 9192 -7030 9292 -7014
rect 9350 -6980 9450 -6942
rect 9350 -7014 9366 -6980
rect 9434 -7014 9450 -6980
rect 9350 -7030 9450 -7014
rect 9508 -6980 9608 -6942
rect 9508 -7014 9524 -6980
rect 9592 -7014 9608 -6980
rect 9508 -7030 9608 -7014
rect 9666 -6980 9766 -6942
rect 9666 -7014 9682 -6980
rect 9750 -7014 9766 -6980
rect 9666 -7030 9766 -7014
rect 9824 -6980 9924 -6942
rect 9824 -7014 9840 -6980
rect 9908 -7014 9924 -6980
rect 9824 -7030 9924 -7014
rect 9982 -6980 10082 -6942
rect 9982 -7014 9998 -6980
rect 10066 -7014 10082 -6980
rect 9982 -7030 10082 -7014
rect 10140 -6980 10240 -6942
rect 10140 -7014 10156 -6980
rect 10224 -7014 10240 -6980
rect 10140 -7030 10240 -7014
rect 10298 -6980 10398 -6942
rect 10298 -7014 10314 -6980
rect 10382 -7014 10398 -6980
rect 10298 -7030 10398 -7014
rect 10456 -6980 10556 -6942
rect 10456 -7014 10472 -6980
rect 10540 -7014 10556 -6980
rect 10456 -7030 10556 -7014
rect 10614 -6980 10714 -6942
rect 10614 -7014 10630 -6980
rect 10698 -7014 10714 -6980
rect 10614 -7030 10714 -7014
rect 10772 -6980 10872 -6942
rect 10772 -7014 10788 -6980
rect 10856 -7014 10872 -6980
rect 10772 -7030 10872 -7014
rect 10930 -6980 11030 -6942
rect 10930 -7014 10946 -6980
rect 11014 -7014 11030 -6980
rect 10930 -7030 11030 -7014
rect 11088 -6980 11188 -6942
rect 11088 -7014 11104 -6980
rect 11172 -7014 11188 -6980
rect 11088 -7030 11188 -7014
rect 11246 -6980 11346 -6942
rect 11246 -7014 11262 -6980
rect 11330 -7014 11346 -6980
rect 11246 -7030 11346 -7014
rect 11404 -6980 11504 -6942
rect 11404 -7014 11420 -6980
rect 11488 -7014 11504 -6980
rect 11404 -7030 11504 -7014
rect 11562 -6980 11662 -6942
rect 11562 -7014 11578 -6980
rect 11646 -7014 11662 -6980
rect 11562 -7030 11662 -7014
rect 11720 -6980 11820 -6942
rect 11720 -7014 11736 -6980
rect 11804 -7014 11820 -6980
rect 11720 -7030 11820 -7014
rect 11878 -6980 11978 -6942
rect 11878 -7014 11894 -6980
rect 11962 -7014 11978 -6980
rect 11878 -7030 11978 -7014
rect 12036 -6980 12136 -6942
rect 12036 -7014 12052 -6980
rect 12120 -7014 12136 -6980
rect 12036 -7030 12136 -7014
rect 12194 -6980 12294 -6942
rect 12194 -7014 12210 -6980
rect 12278 -7014 12294 -6980
rect 12194 -7030 12294 -7014
rect 12352 -6980 12452 -6942
rect 12352 -7014 12368 -6980
rect 12436 -7014 12452 -6980
rect 12352 -7030 12452 -7014
rect 12510 -6980 12610 -6942
rect 12510 -7014 12526 -6980
rect 12594 -7014 12610 -6980
rect 12510 -7030 12610 -7014
rect 14228 -870 14328 -854
rect 14228 -904 14244 -870
rect 14312 -904 14328 -870
rect 14228 -942 14328 -904
rect 14386 -870 14486 -854
rect 14386 -904 14402 -870
rect 14470 -904 14486 -870
rect 14386 -942 14486 -904
rect 14544 -870 14644 -854
rect 14544 -904 14560 -870
rect 14628 -904 14644 -870
rect 14544 -942 14644 -904
rect 14702 -870 14802 -854
rect 14702 -904 14718 -870
rect 14786 -904 14802 -870
rect 14702 -942 14802 -904
rect 14860 -870 14960 -854
rect 14860 -904 14876 -870
rect 14944 -904 14960 -870
rect 14860 -942 14960 -904
rect 15018 -870 15118 -854
rect 15018 -904 15034 -870
rect 15102 -904 15118 -870
rect 15018 -942 15118 -904
rect 15176 -870 15276 -854
rect 15176 -904 15192 -870
rect 15260 -904 15276 -870
rect 15176 -942 15276 -904
rect 15334 -870 15434 -854
rect 15334 -904 15350 -870
rect 15418 -904 15434 -870
rect 15334 -942 15434 -904
rect 15492 -870 15592 -854
rect 15492 -904 15508 -870
rect 15576 -904 15592 -870
rect 15492 -942 15592 -904
rect 15650 -870 15750 -854
rect 15650 -904 15666 -870
rect 15734 -904 15750 -870
rect 15650 -942 15750 -904
rect 15808 -870 15908 -854
rect 15808 -904 15824 -870
rect 15892 -904 15908 -870
rect 15808 -942 15908 -904
rect 15966 -870 16066 -854
rect 15966 -904 15982 -870
rect 16050 -904 16066 -870
rect 15966 -942 16066 -904
rect 16124 -870 16224 -854
rect 16124 -904 16140 -870
rect 16208 -904 16224 -870
rect 16124 -942 16224 -904
rect 16282 -870 16382 -854
rect 16282 -904 16298 -870
rect 16366 -904 16382 -870
rect 16282 -942 16382 -904
rect 16440 -870 16540 -854
rect 16440 -904 16456 -870
rect 16524 -904 16540 -870
rect 16440 -942 16540 -904
rect 16598 -870 16698 -854
rect 16598 -904 16614 -870
rect 16682 -904 16698 -870
rect 16598 -942 16698 -904
rect 16756 -870 16856 -854
rect 16756 -904 16772 -870
rect 16840 -904 16856 -870
rect 16756 -942 16856 -904
rect 16914 -870 17014 -854
rect 16914 -904 16930 -870
rect 16998 -904 17014 -870
rect 16914 -942 17014 -904
rect 17072 -870 17172 -854
rect 17072 -904 17088 -870
rect 17156 -904 17172 -870
rect 17072 -942 17172 -904
rect 17230 -870 17330 -854
rect 17230 -904 17246 -870
rect 17314 -904 17330 -870
rect 17230 -942 17330 -904
rect 17388 -870 17488 -854
rect 17388 -904 17404 -870
rect 17472 -904 17488 -870
rect 17388 -942 17488 -904
rect 17546 -870 17646 -854
rect 17546 -904 17562 -870
rect 17630 -904 17646 -870
rect 17546 -942 17646 -904
rect 17704 -870 17804 -854
rect 17704 -904 17720 -870
rect 17788 -904 17804 -870
rect 17704 -942 17804 -904
rect 17862 -870 17962 -854
rect 17862 -904 17878 -870
rect 17946 -904 17962 -870
rect 17862 -942 17962 -904
rect 18020 -870 18120 -854
rect 18020 -904 18036 -870
rect 18104 -904 18120 -870
rect 18020 -942 18120 -904
rect 18178 -870 18278 -854
rect 18178 -904 18194 -870
rect 18262 -904 18278 -870
rect 18178 -942 18278 -904
rect 18336 -870 18436 -854
rect 18336 -904 18352 -870
rect 18420 -904 18436 -870
rect 18336 -942 18436 -904
rect 18494 -870 18594 -854
rect 18494 -904 18510 -870
rect 18578 -904 18594 -870
rect 18494 -942 18594 -904
rect 18652 -870 18752 -854
rect 18652 -904 18668 -870
rect 18736 -904 18752 -870
rect 18652 -942 18752 -904
rect 18810 -870 18910 -854
rect 18810 -904 18826 -870
rect 18894 -904 18910 -870
rect 18810 -942 18910 -904
rect 14228 -6980 14328 -6942
rect 14228 -7014 14244 -6980
rect 14312 -7014 14328 -6980
rect 14228 -7030 14328 -7014
rect 14386 -6980 14486 -6942
rect 14386 -7014 14402 -6980
rect 14470 -7014 14486 -6980
rect 14386 -7030 14486 -7014
rect 14544 -6980 14644 -6942
rect 14544 -7014 14560 -6980
rect 14628 -7014 14644 -6980
rect 14544 -7030 14644 -7014
rect 14702 -6980 14802 -6942
rect 14702 -7014 14718 -6980
rect 14786 -7014 14802 -6980
rect 14702 -7030 14802 -7014
rect 14860 -6980 14960 -6942
rect 14860 -7014 14876 -6980
rect 14944 -7014 14960 -6980
rect 14860 -7030 14960 -7014
rect 15018 -6980 15118 -6942
rect 15018 -7014 15034 -6980
rect 15102 -7014 15118 -6980
rect 15018 -7030 15118 -7014
rect 15176 -6980 15276 -6942
rect 15176 -7014 15192 -6980
rect 15260 -7014 15276 -6980
rect 15176 -7030 15276 -7014
rect 15334 -6980 15434 -6942
rect 15334 -7014 15350 -6980
rect 15418 -7014 15434 -6980
rect 15334 -7030 15434 -7014
rect 15492 -6980 15592 -6942
rect 15492 -7014 15508 -6980
rect 15576 -7014 15592 -6980
rect 15492 -7030 15592 -7014
rect 15650 -6980 15750 -6942
rect 15650 -7014 15666 -6980
rect 15734 -7014 15750 -6980
rect 15650 -7030 15750 -7014
rect 15808 -6980 15908 -6942
rect 15808 -7014 15824 -6980
rect 15892 -7014 15908 -6980
rect 15808 -7030 15908 -7014
rect 15966 -6980 16066 -6942
rect 15966 -7014 15982 -6980
rect 16050 -7014 16066 -6980
rect 15966 -7030 16066 -7014
rect 16124 -6980 16224 -6942
rect 16124 -7014 16140 -6980
rect 16208 -7014 16224 -6980
rect 16124 -7030 16224 -7014
rect 16282 -6980 16382 -6942
rect 16282 -7014 16298 -6980
rect 16366 -7014 16382 -6980
rect 16282 -7030 16382 -7014
rect 16440 -6980 16540 -6942
rect 16440 -7014 16456 -6980
rect 16524 -7014 16540 -6980
rect 16440 -7030 16540 -7014
rect 16598 -6980 16698 -6942
rect 16598 -7014 16614 -6980
rect 16682 -7014 16698 -6980
rect 16598 -7030 16698 -7014
rect 16756 -6980 16856 -6942
rect 16756 -7014 16772 -6980
rect 16840 -7014 16856 -6980
rect 16756 -7030 16856 -7014
rect 16914 -6980 17014 -6942
rect 16914 -7014 16930 -6980
rect 16998 -7014 17014 -6980
rect 16914 -7030 17014 -7014
rect 17072 -6980 17172 -6942
rect 17072 -7014 17088 -6980
rect 17156 -7014 17172 -6980
rect 17072 -7030 17172 -7014
rect 17230 -6980 17330 -6942
rect 17230 -7014 17246 -6980
rect 17314 -7014 17330 -6980
rect 17230 -7030 17330 -7014
rect 17388 -6980 17488 -6942
rect 17388 -7014 17404 -6980
rect 17472 -7014 17488 -6980
rect 17388 -7030 17488 -7014
rect 17546 -6980 17646 -6942
rect 17546 -7014 17562 -6980
rect 17630 -7014 17646 -6980
rect 17546 -7030 17646 -7014
rect 17704 -6980 17804 -6942
rect 17704 -7014 17720 -6980
rect 17788 -7014 17804 -6980
rect 17704 -7030 17804 -7014
rect 17862 -6980 17962 -6942
rect 17862 -7014 17878 -6980
rect 17946 -7014 17962 -6980
rect 17862 -7030 17962 -7014
rect 18020 -6980 18120 -6942
rect 18020 -7014 18036 -6980
rect 18104 -7014 18120 -6980
rect 18020 -7030 18120 -7014
rect 18178 -6980 18278 -6942
rect 18178 -7014 18194 -6980
rect 18262 -7014 18278 -6980
rect 18178 -7030 18278 -7014
rect 18336 -6980 18436 -6942
rect 18336 -7014 18352 -6980
rect 18420 -7014 18436 -6980
rect 18336 -7030 18436 -7014
rect 18494 -6980 18594 -6942
rect 18494 -7014 18510 -6980
rect 18578 -7014 18594 -6980
rect 18494 -7030 18594 -7014
rect 18652 -6980 18752 -6942
rect 18652 -7014 18668 -6980
rect 18736 -7014 18752 -6980
rect 18652 -7030 18752 -7014
rect 18810 -6980 18910 -6942
rect 18810 -7014 18826 -6980
rect 18894 -7014 18910 -6980
rect 18810 -7030 18910 -7014
rect 20528 -870 20628 -854
rect 20528 -904 20544 -870
rect 20612 -904 20628 -870
rect 20528 -942 20628 -904
rect 20686 -870 20786 -854
rect 20686 -904 20702 -870
rect 20770 -904 20786 -870
rect 20686 -942 20786 -904
rect 20844 -870 20944 -854
rect 20844 -904 20860 -870
rect 20928 -904 20944 -870
rect 20844 -942 20944 -904
rect 21002 -870 21102 -854
rect 21002 -904 21018 -870
rect 21086 -904 21102 -870
rect 21002 -942 21102 -904
rect 21160 -870 21260 -854
rect 21160 -904 21176 -870
rect 21244 -904 21260 -870
rect 21160 -942 21260 -904
rect 21318 -870 21418 -854
rect 21318 -904 21334 -870
rect 21402 -904 21418 -870
rect 21318 -942 21418 -904
rect 21476 -870 21576 -854
rect 21476 -904 21492 -870
rect 21560 -904 21576 -870
rect 21476 -942 21576 -904
rect 21634 -870 21734 -854
rect 21634 -904 21650 -870
rect 21718 -904 21734 -870
rect 21634 -942 21734 -904
rect 21792 -870 21892 -854
rect 21792 -904 21808 -870
rect 21876 -904 21892 -870
rect 21792 -942 21892 -904
rect 21950 -870 22050 -854
rect 21950 -904 21966 -870
rect 22034 -904 22050 -870
rect 21950 -942 22050 -904
rect 22108 -870 22208 -854
rect 22108 -904 22124 -870
rect 22192 -904 22208 -870
rect 22108 -942 22208 -904
rect 22266 -870 22366 -854
rect 22266 -904 22282 -870
rect 22350 -904 22366 -870
rect 22266 -942 22366 -904
rect 22424 -870 22524 -854
rect 22424 -904 22440 -870
rect 22508 -904 22524 -870
rect 22424 -942 22524 -904
rect 22582 -870 22682 -854
rect 22582 -904 22598 -870
rect 22666 -904 22682 -870
rect 22582 -942 22682 -904
rect 22740 -870 22840 -854
rect 22740 -904 22756 -870
rect 22824 -904 22840 -870
rect 22740 -942 22840 -904
rect 22898 -870 22998 -854
rect 22898 -904 22914 -870
rect 22982 -904 22998 -870
rect 22898 -942 22998 -904
rect 23056 -870 23156 -854
rect 23056 -904 23072 -870
rect 23140 -904 23156 -870
rect 23056 -942 23156 -904
rect 23214 -870 23314 -854
rect 23214 -904 23230 -870
rect 23298 -904 23314 -870
rect 23214 -942 23314 -904
rect 23372 -870 23472 -854
rect 23372 -904 23388 -870
rect 23456 -904 23472 -870
rect 23372 -942 23472 -904
rect 23530 -870 23630 -854
rect 23530 -904 23546 -870
rect 23614 -904 23630 -870
rect 23530 -942 23630 -904
rect 23688 -870 23788 -854
rect 23688 -904 23704 -870
rect 23772 -904 23788 -870
rect 23688 -942 23788 -904
rect 23846 -870 23946 -854
rect 23846 -904 23862 -870
rect 23930 -904 23946 -870
rect 23846 -942 23946 -904
rect 24004 -870 24104 -854
rect 24004 -904 24020 -870
rect 24088 -904 24104 -870
rect 24004 -942 24104 -904
rect 24162 -870 24262 -854
rect 24162 -904 24178 -870
rect 24246 -904 24262 -870
rect 24162 -942 24262 -904
rect 24320 -870 24420 -854
rect 24320 -904 24336 -870
rect 24404 -904 24420 -870
rect 24320 -942 24420 -904
rect 24478 -870 24578 -854
rect 24478 -904 24494 -870
rect 24562 -904 24578 -870
rect 24478 -942 24578 -904
rect 24636 -870 24736 -854
rect 24636 -904 24652 -870
rect 24720 -904 24736 -870
rect 24636 -942 24736 -904
rect 24794 -870 24894 -854
rect 24794 -904 24810 -870
rect 24878 -904 24894 -870
rect 24794 -942 24894 -904
rect 24952 -870 25052 -854
rect 24952 -904 24968 -870
rect 25036 -904 25052 -870
rect 24952 -942 25052 -904
rect 25110 -870 25210 -854
rect 25110 -904 25126 -870
rect 25194 -904 25210 -870
rect 25110 -942 25210 -904
rect 20528 -6980 20628 -6942
rect 20528 -7014 20544 -6980
rect 20612 -7014 20628 -6980
rect 20528 -7030 20628 -7014
rect 20686 -6980 20786 -6942
rect 20686 -7014 20702 -6980
rect 20770 -7014 20786 -6980
rect 20686 -7030 20786 -7014
rect 20844 -6980 20944 -6942
rect 20844 -7014 20860 -6980
rect 20928 -7014 20944 -6980
rect 20844 -7030 20944 -7014
rect 21002 -6980 21102 -6942
rect 21002 -7014 21018 -6980
rect 21086 -7014 21102 -6980
rect 21002 -7030 21102 -7014
rect 21160 -6980 21260 -6942
rect 21160 -7014 21176 -6980
rect 21244 -7014 21260 -6980
rect 21160 -7030 21260 -7014
rect 21318 -6980 21418 -6942
rect 21318 -7014 21334 -6980
rect 21402 -7014 21418 -6980
rect 21318 -7030 21418 -7014
rect 21476 -6980 21576 -6942
rect 21476 -7014 21492 -6980
rect 21560 -7014 21576 -6980
rect 21476 -7030 21576 -7014
rect 21634 -6980 21734 -6942
rect 21634 -7014 21650 -6980
rect 21718 -7014 21734 -6980
rect 21634 -7030 21734 -7014
rect 21792 -6980 21892 -6942
rect 21792 -7014 21808 -6980
rect 21876 -7014 21892 -6980
rect 21792 -7030 21892 -7014
rect 21950 -6980 22050 -6942
rect 21950 -7014 21966 -6980
rect 22034 -7014 22050 -6980
rect 21950 -7030 22050 -7014
rect 22108 -6980 22208 -6942
rect 22108 -7014 22124 -6980
rect 22192 -7014 22208 -6980
rect 22108 -7030 22208 -7014
rect 22266 -6980 22366 -6942
rect 22266 -7014 22282 -6980
rect 22350 -7014 22366 -6980
rect 22266 -7030 22366 -7014
rect 22424 -6980 22524 -6942
rect 22424 -7014 22440 -6980
rect 22508 -7014 22524 -6980
rect 22424 -7030 22524 -7014
rect 22582 -6980 22682 -6942
rect 22582 -7014 22598 -6980
rect 22666 -7014 22682 -6980
rect 22582 -7030 22682 -7014
rect 22740 -6980 22840 -6942
rect 22740 -7014 22756 -6980
rect 22824 -7014 22840 -6980
rect 22740 -7030 22840 -7014
rect 22898 -6980 22998 -6942
rect 22898 -7014 22914 -6980
rect 22982 -7014 22998 -6980
rect 22898 -7030 22998 -7014
rect 23056 -6980 23156 -6942
rect 23056 -7014 23072 -6980
rect 23140 -7014 23156 -6980
rect 23056 -7030 23156 -7014
rect 23214 -6980 23314 -6942
rect 23214 -7014 23230 -6980
rect 23298 -7014 23314 -6980
rect 23214 -7030 23314 -7014
rect 23372 -6980 23472 -6942
rect 23372 -7014 23388 -6980
rect 23456 -7014 23472 -6980
rect 23372 -7030 23472 -7014
rect 23530 -6980 23630 -6942
rect 23530 -7014 23546 -6980
rect 23614 -7014 23630 -6980
rect 23530 -7030 23630 -7014
rect 23688 -6980 23788 -6942
rect 23688 -7014 23704 -6980
rect 23772 -7014 23788 -6980
rect 23688 -7030 23788 -7014
rect 23846 -6980 23946 -6942
rect 23846 -7014 23862 -6980
rect 23930 -7014 23946 -6980
rect 23846 -7030 23946 -7014
rect 24004 -6980 24104 -6942
rect 24004 -7014 24020 -6980
rect 24088 -7014 24104 -6980
rect 24004 -7030 24104 -7014
rect 24162 -6980 24262 -6942
rect 24162 -7014 24178 -6980
rect 24246 -7014 24262 -6980
rect 24162 -7030 24262 -7014
rect 24320 -6980 24420 -6942
rect 24320 -7014 24336 -6980
rect 24404 -7014 24420 -6980
rect 24320 -7030 24420 -7014
rect 24478 -6980 24578 -6942
rect 24478 -7014 24494 -6980
rect 24562 -7014 24578 -6980
rect 24478 -7030 24578 -7014
rect 24636 -6980 24736 -6942
rect 24636 -7014 24652 -6980
rect 24720 -7014 24736 -6980
rect 24636 -7030 24736 -7014
rect 24794 -6980 24894 -6942
rect 24794 -7014 24810 -6980
rect 24878 -7014 24894 -6980
rect 24794 -7030 24894 -7014
rect 24952 -6980 25052 -6942
rect 24952 -7014 24968 -6980
rect 25036 -7014 25052 -6980
rect 24952 -7030 25052 -7014
rect 25110 -6980 25210 -6942
rect 25110 -7014 25126 -6980
rect 25194 -7014 25210 -6980
rect 25110 -7030 25210 -7014
<< polycont >>
rect 1644 6696 1712 6730
rect 1802 6696 1870 6730
rect 1960 6696 2028 6730
rect 2118 6696 2186 6730
rect 2276 6696 2344 6730
rect 2434 6696 2502 6730
rect 2592 6696 2660 6730
rect 2750 6696 2818 6730
rect 2908 6696 2976 6730
rect 3066 6696 3134 6730
rect 3224 6696 3292 6730
rect 3382 6696 3450 6730
rect 3540 6696 3608 6730
rect 3698 6696 3766 6730
rect 3856 6696 3924 6730
rect 4014 6696 4082 6730
rect 4172 6696 4240 6730
rect 4330 6696 4398 6730
rect 4488 6696 4556 6730
rect 4646 6696 4714 6730
rect 4804 6696 4872 6730
rect 4962 6696 5030 6730
rect 5120 6696 5188 6730
rect 5278 6696 5346 6730
rect 5436 6696 5504 6730
rect 5594 6696 5662 6730
rect 5752 6696 5820 6730
rect 5910 6696 5978 6730
rect 6068 6696 6136 6730
rect 6226 6696 6294 6730
rect 1644 586 1712 620
rect 1802 586 1870 620
rect 1960 586 2028 620
rect 2118 586 2186 620
rect 2276 586 2344 620
rect 2434 586 2502 620
rect 2592 586 2660 620
rect 2750 586 2818 620
rect 2908 586 2976 620
rect 3066 586 3134 620
rect 3224 586 3292 620
rect 3382 586 3450 620
rect 3540 586 3608 620
rect 3698 586 3766 620
rect 3856 586 3924 620
rect 4014 586 4082 620
rect 4172 586 4240 620
rect 4330 586 4398 620
rect 4488 586 4556 620
rect 4646 586 4714 620
rect 4804 586 4872 620
rect 4962 586 5030 620
rect 5120 586 5188 620
rect 5278 586 5346 620
rect 5436 586 5504 620
rect 5594 586 5662 620
rect 5752 586 5820 620
rect 5910 586 5978 620
rect 6068 586 6136 620
rect 6226 586 6294 620
rect 7944 6696 8012 6730
rect 8102 6696 8170 6730
rect 8260 6696 8328 6730
rect 8418 6696 8486 6730
rect 8576 6696 8644 6730
rect 8734 6696 8802 6730
rect 8892 6696 8960 6730
rect 9050 6696 9118 6730
rect 9208 6696 9276 6730
rect 9366 6696 9434 6730
rect 9524 6696 9592 6730
rect 9682 6696 9750 6730
rect 9840 6696 9908 6730
rect 9998 6696 10066 6730
rect 10156 6696 10224 6730
rect 10314 6696 10382 6730
rect 10472 6696 10540 6730
rect 10630 6696 10698 6730
rect 10788 6696 10856 6730
rect 10946 6696 11014 6730
rect 11104 6696 11172 6730
rect 11262 6696 11330 6730
rect 11420 6696 11488 6730
rect 11578 6696 11646 6730
rect 11736 6696 11804 6730
rect 11894 6696 11962 6730
rect 12052 6696 12120 6730
rect 12210 6696 12278 6730
rect 12368 6696 12436 6730
rect 12526 6696 12594 6730
rect 7944 586 8012 620
rect 8102 586 8170 620
rect 8260 586 8328 620
rect 8418 586 8486 620
rect 8576 586 8644 620
rect 8734 586 8802 620
rect 8892 586 8960 620
rect 9050 586 9118 620
rect 9208 586 9276 620
rect 9366 586 9434 620
rect 9524 586 9592 620
rect 9682 586 9750 620
rect 9840 586 9908 620
rect 9998 586 10066 620
rect 10156 586 10224 620
rect 10314 586 10382 620
rect 10472 586 10540 620
rect 10630 586 10698 620
rect 10788 586 10856 620
rect 10946 586 11014 620
rect 11104 586 11172 620
rect 11262 586 11330 620
rect 11420 586 11488 620
rect 11578 586 11646 620
rect 11736 586 11804 620
rect 11894 586 11962 620
rect 12052 586 12120 620
rect 12210 586 12278 620
rect 12368 586 12436 620
rect 12526 586 12594 620
rect 14244 6696 14312 6730
rect 14402 6696 14470 6730
rect 14560 6696 14628 6730
rect 14718 6696 14786 6730
rect 14876 6696 14944 6730
rect 15034 6696 15102 6730
rect 15192 6696 15260 6730
rect 15350 6696 15418 6730
rect 15508 6696 15576 6730
rect 15666 6696 15734 6730
rect 15824 6696 15892 6730
rect 15982 6696 16050 6730
rect 16140 6696 16208 6730
rect 16298 6696 16366 6730
rect 16456 6696 16524 6730
rect 16614 6696 16682 6730
rect 16772 6696 16840 6730
rect 16930 6696 16998 6730
rect 17088 6696 17156 6730
rect 17246 6696 17314 6730
rect 17404 6696 17472 6730
rect 17562 6696 17630 6730
rect 17720 6696 17788 6730
rect 17878 6696 17946 6730
rect 18036 6696 18104 6730
rect 18194 6696 18262 6730
rect 18352 6696 18420 6730
rect 18510 6696 18578 6730
rect 18668 6696 18736 6730
rect 18826 6696 18894 6730
rect 14244 586 14312 620
rect 14402 586 14470 620
rect 14560 586 14628 620
rect 14718 586 14786 620
rect 14876 586 14944 620
rect 15034 586 15102 620
rect 15192 586 15260 620
rect 15350 586 15418 620
rect 15508 586 15576 620
rect 15666 586 15734 620
rect 15824 586 15892 620
rect 15982 586 16050 620
rect 16140 586 16208 620
rect 16298 586 16366 620
rect 16456 586 16524 620
rect 16614 586 16682 620
rect 16772 586 16840 620
rect 16930 586 16998 620
rect 17088 586 17156 620
rect 17246 586 17314 620
rect 17404 586 17472 620
rect 17562 586 17630 620
rect 17720 586 17788 620
rect 17878 586 17946 620
rect 18036 586 18104 620
rect 18194 586 18262 620
rect 18352 586 18420 620
rect 18510 586 18578 620
rect 18668 586 18736 620
rect 18826 586 18894 620
rect 20544 6696 20612 6730
rect 20702 6696 20770 6730
rect 20860 6696 20928 6730
rect 21018 6696 21086 6730
rect 21176 6696 21244 6730
rect 21334 6696 21402 6730
rect 21492 6696 21560 6730
rect 21650 6696 21718 6730
rect 21808 6696 21876 6730
rect 21966 6696 22034 6730
rect 22124 6696 22192 6730
rect 22282 6696 22350 6730
rect 22440 6696 22508 6730
rect 22598 6696 22666 6730
rect 22756 6696 22824 6730
rect 22914 6696 22982 6730
rect 23072 6696 23140 6730
rect 23230 6696 23298 6730
rect 23388 6696 23456 6730
rect 23546 6696 23614 6730
rect 23704 6696 23772 6730
rect 23862 6696 23930 6730
rect 24020 6696 24088 6730
rect 24178 6696 24246 6730
rect 24336 6696 24404 6730
rect 24494 6696 24562 6730
rect 24652 6696 24720 6730
rect 24810 6696 24878 6730
rect 24968 6696 25036 6730
rect 25126 6696 25194 6730
rect 20544 586 20612 620
rect 20702 586 20770 620
rect 20860 586 20928 620
rect 21018 586 21086 620
rect 21176 586 21244 620
rect 21334 586 21402 620
rect 21492 586 21560 620
rect 21650 586 21718 620
rect 21808 586 21876 620
rect 21966 586 22034 620
rect 22124 586 22192 620
rect 22282 586 22350 620
rect 22440 586 22508 620
rect 22598 586 22666 620
rect 22756 586 22824 620
rect 22914 586 22982 620
rect 23072 586 23140 620
rect 23230 586 23298 620
rect 23388 586 23456 620
rect 23546 586 23614 620
rect 23704 586 23772 620
rect 23862 586 23930 620
rect 24020 586 24088 620
rect 24178 586 24246 620
rect 24336 586 24404 620
rect 24494 586 24562 620
rect 24652 586 24720 620
rect 24810 586 24878 620
rect 24968 586 25036 620
rect 25126 586 25194 620
rect 1644 -904 1712 -870
rect 1802 -904 1870 -870
rect 1960 -904 2028 -870
rect 2118 -904 2186 -870
rect 2276 -904 2344 -870
rect 2434 -904 2502 -870
rect 2592 -904 2660 -870
rect 2750 -904 2818 -870
rect 2908 -904 2976 -870
rect 3066 -904 3134 -870
rect 3224 -904 3292 -870
rect 3382 -904 3450 -870
rect 3540 -904 3608 -870
rect 3698 -904 3766 -870
rect 3856 -904 3924 -870
rect 4014 -904 4082 -870
rect 4172 -904 4240 -870
rect 4330 -904 4398 -870
rect 4488 -904 4556 -870
rect 4646 -904 4714 -870
rect 4804 -904 4872 -870
rect 4962 -904 5030 -870
rect 5120 -904 5188 -870
rect 5278 -904 5346 -870
rect 5436 -904 5504 -870
rect 5594 -904 5662 -870
rect 5752 -904 5820 -870
rect 5910 -904 5978 -870
rect 6068 -904 6136 -870
rect 6226 -904 6294 -870
rect 1644 -7014 1712 -6980
rect 1802 -7014 1870 -6980
rect 1960 -7014 2028 -6980
rect 2118 -7014 2186 -6980
rect 2276 -7014 2344 -6980
rect 2434 -7014 2502 -6980
rect 2592 -7014 2660 -6980
rect 2750 -7014 2818 -6980
rect 2908 -7014 2976 -6980
rect 3066 -7014 3134 -6980
rect 3224 -7014 3292 -6980
rect 3382 -7014 3450 -6980
rect 3540 -7014 3608 -6980
rect 3698 -7014 3766 -6980
rect 3856 -7014 3924 -6980
rect 4014 -7014 4082 -6980
rect 4172 -7014 4240 -6980
rect 4330 -7014 4398 -6980
rect 4488 -7014 4556 -6980
rect 4646 -7014 4714 -6980
rect 4804 -7014 4872 -6980
rect 4962 -7014 5030 -6980
rect 5120 -7014 5188 -6980
rect 5278 -7014 5346 -6980
rect 5436 -7014 5504 -6980
rect 5594 -7014 5662 -6980
rect 5752 -7014 5820 -6980
rect 5910 -7014 5978 -6980
rect 6068 -7014 6136 -6980
rect 6226 -7014 6294 -6980
rect 7944 -904 8012 -870
rect 8102 -904 8170 -870
rect 8260 -904 8328 -870
rect 8418 -904 8486 -870
rect 8576 -904 8644 -870
rect 8734 -904 8802 -870
rect 8892 -904 8960 -870
rect 9050 -904 9118 -870
rect 9208 -904 9276 -870
rect 9366 -904 9434 -870
rect 9524 -904 9592 -870
rect 9682 -904 9750 -870
rect 9840 -904 9908 -870
rect 9998 -904 10066 -870
rect 10156 -904 10224 -870
rect 10314 -904 10382 -870
rect 10472 -904 10540 -870
rect 10630 -904 10698 -870
rect 10788 -904 10856 -870
rect 10946 -904 11014 -870
rect 11104 -904 11172 -870
rect 11262 -904 11330 -870
rect 11420 -904 11488 -870
rect 11578 -904 11646 -870
rect 11736 -904 11804 -870
rect 11894 -904 11962 -870
rect 12052 -904 12120 -870
rect 12210 -904 12278 -870
rect 12368 -904 12436 -870
rect 12526 -904 12594 -870
rect 7944 -7014 8012 -6980
rect 8102 -7014 8170 -6980
rect 8260 -7014 8328 -6980
rect 8418 -7014 8486 -6980
rect 8576 -7014 8644 -6980
rect 8734 -7014 8802 -6980
rect 8892 -7014 8960 -6980
rect 9050 -7014 9118 -6980
rect 9208 -7014 9276 -6980
rect 9366 -7014 9434 -6980
rect 9524 -7014 9592 -6980
rect 9682 -7014 9750 -6980
rect 9840 -7014 9908 -6980
rect 9998 -7014 10066 -6980
rect 10156 -7014 10224 -6980
rect 10314 -7014 10382 -6980
rect 10472 -7014 10540 -6980
rect 10630 -7014 10698 -6980
rect 10788 -7014 10856 -6980
rect 10946 -7014 11014 -6980
rect 11104 -7014 11172 -6980
rect 11262 -7014 11330 -6980
rect 11420 -7014 11488 -6980
rect 11578 -7014 11646 -6980
rect 11736 -7014 11804 -6980
rect 11894 -7014 11962 -6980
rect 12052 -7014 12120 -6980
rect 12210 -7014 12278 -6980
rect 12368 -7014 12436 -6980
rect 12526 -7014 12594 -6980
rect 14244 -904 14312 -870
rect 14402 -904 14470 -870
rect 14560 -904 14628 -870
rect 14718 -904 14786 -870
rect 14876 -904 14944 -870
rect 15034 -904 15102 -870
rect 15192 -904 15260 -870
rect 15350 -904 15418 -870
rect 15508 -904 15576 -870
rect 15666 -904 15734 -870
rect 15824 -904 15892 -870
rect 15982 -904 16050 -870
rect 16140 -904 16208 -870
rect 16298 -904 16366 -870
rect 16456 -904 16524 -870
rect 16614 -904 16682 -870
rect 16772 -904 16840 -870
rect 16930 -904 16998 -870
rect 17088 -904 17156 -870
rect 17246 -904 17314 -870
rect 17404 -904 17472 -870
rect 17562 -904 17630 -870
rect 17720 -904 17788 -870
rect 17878 -904 17946 -870
rect 18036 -904 18104 -870
rect 18194 -904 18262 -870
rect 18352 -904 18420 -870
rect 18510 -904 18578 -870
rect 18668 -904 18736 -870
rect 18826 -904 18894 -870
rect 14244 -7014 14312 -6980
rect 14402 -7014 14470 -6980
rect 14560 -7014 14628 -6980
rect 14718 -7014 14786 -6980
rect 14876 -7014 14944 -6980
rect 15034 -7014 15102 -6980
rect 15192 -7014 15260 -6980
rect 15350 -7014 15418 -6980
rect 15508 -7014 15576 -6980
rect 15666 -7014 15734 -6980
rect 15824 -7014 15892 -6980
rect 15982 -7014 16050 -6980
rect 16140 -7014 16208 -6980
rect 16298 -7014 16366 -6980
rect 16456 -7014 16524 -6980
rect 16614 -7014 16682 -6980
rect 16772 -7014 16840 -6980
rect 16930 -7014 16998 -6980
rect 17088 -7014 17156 -6980
rect 17246 -7014 17314 -6980
rect 17404 -7014 17472 -6980
rect 17562 -7014 17630 -6980
rect 17720 -7014 17788 -6980
rect 17878 -7014 17946 -6980
rect 18036 -7014 18104 -6980
rect 18194 -7014 18262 -6980
rect 18352 -7014 18420 -6980
rect 18510 -7014 18578 -6980
rect 18668 -7014 18736 -6980
rect 18826 -7014 18894 -6980
rect 20544 -904 20612 -870
rect 20702 -904 20770 -870
rect 20860 -904 20928 -870
rect 21018 -904 21086 -870
rect 21176 -904 21244 -870
rect 21334 -904 21402 -870
rect 21492 -904 21560 -870
rect 21650 -904 21718 -870
rect 21808 -904 21876 -870
rect 21966 -904 22034 -870
rect 22124 -904 22192 -870
rect 22282 -904 22350 -870
rect 22440 -904 22508 -870
rect 22598 -904 22666 -870
rect 22756 -904 22824 -870
rect 22914 -904 22982 -870
rect 23072 -904 23140 -870
rect 23230 -904 23298 -870
rect 23388 -904 23456 -870
rect 23546 -904 23614 -870
rect 23704 -904 23772 -870
rect 23862 -904 23930 -870
rect 24020 -904 24088 -870
rect 24178 -904 24246 -870
rect 24336 -904 24404 -870
rect 24494 -904 24562 -870
rect 24652 -904 24720 -870
rect 24810 -904 24878 -870
rect 24968 -904 25036 -870
rect 25126 -904 25194 -870
rect 20544 -7014 20612 -6980
rect 20702 -7014 20770 -6980
rect 20860 -7014 20928 -6980
rect 21018 -7014 21086 -6980
rect 21176 -7014 21244 -6980
rect 21334 -7014 21402 -6980
rect 21492 -7014 21560 -6980
rect 21650 -7014 21718 -6980
rect 21808 -7014 21876 -6980
rect 21966 -7014 22034 -6980
rect 22124 -7014 22192 -6980
rect 22282 -7014 22350 -6980
rect 22440 -7014 22508 -6980
rect 22598 -7014 22666 -6980
rect 22756 -7014 22824 -6980
rect 22914 -7014 22982 -6980
rect 23072 -7014 23140 -6980
rect 23230 -7014 23298 -6980
rect 23388 -7014 23456 -6980
rect 23546 -7014 23614 -6980
rect 23704 -7014 23772 -6980
rect 23862 -7014 23930 -6980
rect 24020 -7014 24088 -6980
rect 24178 -7014 24246 -6980
rect 24336 -7014 24404 -6980
rect 24494 -7014 24562 -6980
rect 24652 -7014 24720 -6980
rect 24810 -7014 24878 -6980
rect 24968 -7014 25036 -6980
rect 25126 -7014 25194 -6980
<< locali >>
rect 1448 6834 1544 6868
rect 6394 6834 6490 6868
rect 1448 6772 1482 6834
rect 6456 6772 6490 6834
rect 1628 6696 1644 6730
rect 1712 6696 1728 6730
rect 1786 6696 1802 6730
rect 1870 6696 1886 6730
rect 1944 6696 1960 6730
rect 2028 6696 2044 6730
rect 2102 6696 2118 6730
rect 2186 6696 2202 6730
rect 2260 6696 2276 6730
rect 2344 6696 2360 6730
rect 2418 6696 2434 6730
rect 2502 6696 2518 6730
rect 2576 6696 2592 6730
rect 2660 6696 2676 6730
rect 2734 6696 2750 6730
rect 2818 6696 2834 6730
rect 2892 6696 2908 6730
rect 2976 6696 2992 6730
rect 3050 6696 3066 6730
rect 3134 6696 3150 6730
rect 3208 6696 3224 6730
rect 3292 6696 3308 6730
rect 3366 6696 3382 6730
rect 3450 6696 3466 6730
rect 3524 6696 3540 6730
rect 3608 6696 3624 6730
rect 3682 6696 3698 6730
rect 3766 6696 3782 6730
rect 3840 6696 3856 6730
rect 3924 6696 3940 6730
rect 3998 6696 4014 6730
rect 4082 6696 4098 6730
rect 4156 6696 4172 6730
rect 4240 6696 4256 6730
rect 4314 6696 4330 6730
rect 4398 6696 4414 6730
rect 4472 6696 4488 6730
rect 4556 6696 4572 6730
rect 4630 6696 4646 6730
rect 4714 6696 4730 6730
rect 4788 6696 4804 6730
rect 4872 6696 4888 6730
rect 4946 6696 4962 6730
rect 5030 6696 5046 6730
rect 5104 6696 5120 6730
rect 5188 6696 5204 6730
rect 5262 6696 5278 6730
rect 5346 6696 5362 6730
rect 5420 6696 5436 6730
rect 5504 6696 5520 6730
rect 5578 6696 5594 6730
rect 5662 6696 5678 6730
rect 5736 6696 5752 6730
rect 5820 6696 5836 6730
rect 5894 6696 5910 6730
rect 5978 6696 5994 6730
rect 6052 6696 6068 6730
rect 6136 6696 6152 6730
rect 6210 6696 6226 6730
rect 6294 6696 6310 6730
rect 7748 6834 7844 6868
rect 12694 6834 12790 6868
rect 7748 6772 7782 6834
rect 12756 6772 12790 6834
rect 7928 6696 7944 6730
rect 8012 6696 8028 6730
rect 8086 6696 8102 6730
rect 8170 6696 8186 6730
rect 8244 6696 8260 6730
rect 8328 6696 8344 6730
rect 8402 6696 8418 6730
rect 8486 6696 8502 6730
rect 8560 6696 8576 6730
rect 8644 6696 8660 6730
rect 8718 6696 8734 6730
rect 8802 6696 8818 6730
rect 8876 6696 8892 6730
rect 8960 6696 8976 6730
rect 9034 6696 9050 6730
rect 9118 6696 9134 6730
rect 9192 6696 9208 6730
rect 9276 6696 9292 6730
rect 9350 6696 9366 6730
rect 9434 6696 9450 6730
rect 9508 6696 9524 6730
rect 9592 6696 9608 6730
rect 9666 6696 9682 6730
rect 9750 6696 9766 6730
rect 9824 6696 9840 6730
rect 9908 6696 9924 6730
rect 9982 6696 9998 6730
rect 10066 6696 10082 6730
rect 10140 6696 10156 6730
rect 10224 6696 10240 6730
rect 10298 6696 10314 6730
rect 10382 6696 10398 6730
rect 10456 6696 10472 6730
rect 10540 6696 10556 6730
rect 10614 6696 10630 6730
rect 10698 6696 10714 6730
rect 10772 6696 10788 6730
rect 10856 6696 10872 6730
rect 10930 6696 10946 6730
rect 11014 6696 11030 6730
rect 11088 6696 11104 6730
rect 11172 6696 11188 6730
rect 11246 6696 11262 6730
rect 11330 6696 11346 6730
rect 11404 6696 11420 6730
rect 11488 6696 11504 6730
rect 11562 6696 11578 6730
rect 11646 6696 11662 6730
rect 11720 6696 11736 6730
rect 11804 6696 11820 6730
rect 11878 6696 11894 6730
rect 11962 6696 11978 6730
rect 12036 6696 12052 6730
rect 12120 6696 12136 6730
rect 12194 6696 12210 6730
rect 12278 6696 12294 6730
rect 12352 6696 12368 6730
rect 12436 6696 12452 6730
rect 12510 6696 12526 6730
rect 12594 6696 12610 6730
rect 14048 6834 14144 6868
rect 18994 6834 19090 6868
rect 14048 6772 14082 6834
rect 19056 6772 19090 6834
rect 14228 6696 14244 6730
rect 14312 6696 14328 6730
rect 14386 6696 14402 6730
rect 14470 6696 14486 6730
rect 14544 6696 14560 6730
rect 14628 6696 14644 6730
rect 14702 6696 14718 6730
rect 14786 6696 14802 6730
rect 14860 6696 14876 6730
rect 14944 6696 14960 6730
rect 15018 6696 15034 6730
rect 15102 6696 15118 6730
rect 15176 6696 15192 6730
rect 15260 6696 15276 6730
rect 15334 6696 15350 6730
rect 15418 6696 15434 6730
rect 15492 6696 15508 6730
rect 15576 6696 15592 6730
rect 15650 6696 15666 6730
rect 15734 6696 15750 6730
rect 15808 6696 15824 6730
rect 15892 6696 15908 6730
rect 15966 6696 15982 6730
rect 16050 6696 16066 6730
rect 16124 6696 16140 6730
rect 16208 6696 16224 6730
rect 16282 6696 16298 6730
rect 16366 6696 16382 6730
rect 16440 6696 16456 6730
rect 16524 6696 16540 6730
rect 16598 6696 16614 6730
rect 16682 6696 16698 6730
rect 16756 6696 16772 6730
rect 16840 6696 16856 6730
rect 16914 6696 16930 6730
rect 16998 6696 17014 6730
rect 17072 6696 17088 6730
rect 17156 6696 17172 6730
rect 17230 6696 17246 6730
rect 17314 6696 17330 6730
rect 17388 6696 17404 6730
rect 17472 6696 17488 6730
rect 17546 6696 17562 6730
rect 17630 6696 17646 6730
rect 17704 6696 17720 6730
rect 17788 6696 17804 6730
rect 17862 6696 17878 6730
rect 17946 6696 17962 6730
rect 18020 6696 18036 6730
rect 18104 6696 18120 6730
rect 18178 6696 18194 6730
rect 18262 6696 18278 6730
rect 18336 6696 18352 6730
rect 18420 6696 18436 6730
rect 18494 6696 18510 6730
rect 18578 6696 18594 6730
rect 18652 6696 18668 6730
rect 18736 6696 18752 6730
rect 18810 6696 18826 6730
rect 18894 6696 18910 6730
rect 20348 6834 20444 6868
rect 25294 6834 25390 6868
rect 20348 6772 20382 6834
rect 25356 6772 25390 6834
rect 20528 6696 20544 6730
rect 20612 6696 20628 6730
rect 20686 6696 20702 6730
rect 20770 6696 20786 6730
rect 20844 6696 20860 6730
rect 20928 6696 20944 6730
rect 21002 6696 21018 6730
rect 21086 6696 21102 6730
rect 21160 6696 21176 6730
rect 21244 6696 21260 6730
rect 21318 6696 21334 6730
rect 21402 6696 21418 6730
rect 21476 6696 21492 6730
rect 21560 6696 21576 6730
rect 21634 6696 21650 6730
rect 21718 6696 21734 6730
rect 21792 6696 21808 6730
rect 21876 6696 21892 6730
rect 21950 6696 21966 6730
rect 22034 6696 22050 6730
rect 22108 6696 22124 6730
rect 22192 6696 22208 6730
rect 22266 6696 22282 6730
rect 22350 6696 22366 6730
rect 22424 6696 22440 6730
rect 22508 6696 22524 6730
rect 22582 6696 22598 6730
rect 22666 6696 22682 6730
rect 22740 6696 22756 6730
rect 22824 6696 22840 6730
rect 22898 6696 22914 6730
rect 22982 6696 22998 6730
rect 23056 6696 23072 6730
rect 23140 6696 23156 6730
rect 23214 6696 23230 6730
rect 23298 6696 23314 6730
rect 23372 6696 23388 6730
rect 23456 6696 23472 6730
rect 23530 6696 23546 6730
rect 23614 6696 23630 6730
rect 23688 6696 23704 6730
rect 23772 6696 23788 6730
rect 23846 6696 23862 6730
rect 23930 6696 23946 6730
rect 24004 6696 24020 6730
rect 24088 6696 24104 6730
rect 24162 6696 24178 6730
rect 24246 6696 24262 6730
rect 24320 6696 24336 6730
rect 24404 6696 24420 6730
rect 24478 6696 24494 6730
rect 24562 6696 24578 6730
rect 24636 6696 24652 6730
rect 24720 6696 24736 6730
rect 24794 6696 24810 6730
rect 24878 6696 24894 6730
rect 24952 6696 24968 6730
rect 25036 6696 25052 6730
rect 25110 6696 25126 6730
rect 25194 6696 25210 6730
rect 1582 6646 1616 6662
rect 1582 654 1616 670
rect 1740 6646 1774 6662
rect 1740 654 1774 670
rect 1898 6646 1932 6662
rect 1898 654 1932 670
rect 2056 6646 2090 6662
rect 2056 654 2090 670
rect 2214 6646 2248 6662
rect 2214 654 2248 670
rect 2372 6646 2406 6662
rect 2372 654 2406 670
rect 2530 6646 2564 6662
rect 2530 654 2564 670
rect 2688 6646 2722 6662
rect 2688 654 2722 670
rect 2846 6646 2880 6662
rect 2846 654 2880 670
rect 3004 6646 3038 6662
rect 3004 654 3038 670
rect 3162 6646 3196 6662
rect 3162 654 3196 670
rect 3320 6646 3354 6662
rect 3320 654 3354 670
rect 3478 6646 3512 6662
rect 3478 654 3512 670
rect 3636 6646 3670 6662
rect 3636 654 3670 670
rect 3794 6646 3828 6662
rect 3794 654 3828 670
rect 3952 6646 3986 6662
rect 3952 654 3986 670
rect 4110 6646 4144 6662
rect 4110 654 4144 670
rect 4268 6646 4302 6662
rect 4268 654 4302 670
rect 4426 6646 4460 6662
rect 4426 654 4460 670
rect 4584 6646 4618 6662
rect 4584 654 4618 670
rect 4742 6646 4776 6662
rect 4742 654 4776 670
rect 4900 6646 4934 6662
rect 4900 654 4934 670
rect 5058 6646 5092 6662
rect 5058 654 5092 670
rect 5216 6646 5250 6662
rect 5216 654 5250 670
rect 5374 6646 5408 6662
rect 5374 654 5408 670
rect 5532 6646 5566 6662
rect 5532 654 5566 670
rect 5690 6646 5724 6662
rect 5690 654 5724 670
rect 5848 6646 5882 6662
rect 5848 654 5882 670
rect 6006 6646 6040 6662
rect 6006 654 6040 670
rect 6164 6646 6198 6662
rect 6164 654 6198 670
rect 6322 6646 6356 6662
rect 6322 654 6356 670
rect 7882 6646 7916 6662
rect 7882 654 7916 670
rect 8040 6646 8074 6662
rect 8040 654 8074 670
rect 8198 6646 8232 6662
rect 8198 654 8232 670
rect 8356 6646 8390 6662
rect 8356 654 8390 670
rect 8514 6646 8548 6662
rect 8514 654 8548 670
rect 8672 6646 8706 6662
rect 8672 654 8706 670
rect 8830 6646 8864 6662
rect 8830 654 8864 670
rect 8988 6646 9022 6662
rect 8988 654 9022 670
rect 9146 6646 9180 6662
rect 9146 654 9180 670
rect 9304 6646 9338 6662
rect 9304 654 9338 670
rect 9462 6646 9496 6662
rect 9462 654 9496 670
rect 9620 6646 9654 6662
rect 9620 654 9654 670
rect 9778 6646 9812 6662
rect 9778 654 9812 670
rect 9936 6646 9970 6662
rect 9936 654 9970 670
rect 10094 6646 10128 6662
rect 10094 654 10128 670
rect 10252 6646 10286 6662
rect 10252 654 10286 670
rect 10410 6646 10444 6662
rect 10410 654 10444 670
rect 10568 6646 10602 6662
rect 10568 654 10602 670
rect 10726 6646 10760 6662
rect 10726 654 10760 670
rect 10884 6646 10918 6662
rect 10884 654 10918 670
rect 11042 6646 11076 6662
rect 11042 654 11076 670
rect 11200 6646 11234 6662
rect 11200 654 11234 670
rect 11358 6646 11392 6662
rect 11358 654 11392 670
rect 11516 6646 11550 6662
rect 11516 654 11550 670
rect 11674 6646 11708 6662
rect 11674 654 11708 670
rect 11832 6646 11866 6662
rect 11832 654 11866 670
rect 11990 6646 12024 6662
rect 11990 654 12024 670
rect 12148 6646 12182 6662
rect 12148 654 12182 670
rect 12306 6646 12340 6662
rect 12306 654 12340 670
rect 12464 6646 12498 6662
rect 12464 654 12498 670
rect 12622 6646 12656 6662
rect 12622 654 12656 670
rect 14182 6646 14216 6662
rect 14182 654 14216 670
rect 14340 6646 14374 6662
rect 14340 654 14374 670
rect 14498 6646 14532 6662
rect 14498 654 14532 670
rect 14656 6646 14690 6662
rect 14656 654 14690 670
rect 14814 6646 14848 6662
rect 14814 654 14848 670
rect 14972 6646 15006 6662
rect 14972 654 15006 670
rect 15130 6646 15164 6662
rect 15130 654 15164 670
rect 15288 6646 15322 6662
rect 15288 654 15322 670
rect 15446 6646 15480 6662
rect 15446 654 15480 670
rect 15604 6646 15638 6662
rect 15604 654 15638 670
rect 15762 6646 15796 6662
rect 15762 654 15796 670
rect 15920 6646 15954 6662
rect 15920 654 15954 670
rect 16078 6646 16112 6662
rect 16078 654 16112 670
rect 16236 6646 16270 6662
rect 16236 654 16270 670
rect 16394 6646 16428 6662
rect 16394 654 16428 670
rect 16552 6646 16586 6662
rect 16552 654 16586 670
rect 16710 6646 16744 6662
rect 16710 654 16744 670
rect 16868 6646 16902 6662
rect 16868 654 16902 670
rect 17026 6646 17060 6662
rect 17026 654 17060 670
rect 17184 6646 17218 6662
rect 17184 654 17218 670
rect 17342 6646 17376 6662
rect 17342 654 17376 670
rect 17500 6646 17534 6662
rect 17500 654 17534 670
rect 17658 6646 17692 6662
rect 17658 654 17692 670
rect 17816 6646 17850 6662
rect 17816 654 17850 670
rect 17974 6646 18008 6662
rect 17974 654 18008 670
rect 18132 6646 18166 6662
rect 18132 654 18166 670
rect 18290 6646 18324 6662
rect 18290 654 18324 670
rect 18448 6646 18482 6662
rect 18448 654 18482 670
rect 18606 6646 18640 6662
rect 18606 654 18640 670
rect 18764 6646 18798 6662
rect 18764 654 18798 670
rect 18922 6646 18956 6662
rect 18922 654 18956 670
rect 20482 6646 20516 6662
rect 20482 654 20516 670
rect 20640 6646 20674 6662
rect 20640 654 20674 670
rect 20798 6646 20832 6662
rect 20798 654 20832 670
rect 20956 6646 20990 6662
rect 20956 654 20990 670
rect 21114 6646 21148 6662
rect 21114 654 21148 670
rect 21272 6646 21306 6662
rect 21272 654 21306 670
rect 21430 6646 21464 6662
rect 21430 654 21464 670
rect 21588 6646 21622 6662
rect 21588 654 21622 670
rect 21746 6646 21780 6662
rect 21746 654 21780 670
rect 21904 6646 21938 6662
rect 21904 654 21938 670
rect 22062 6646 22096 6662
rect 22062 654 22096 670
rect 22220 6646 22254 6662
rect 22220 654 22254 670
rect 22378 6646 22412 6662
rect 22378 654 22412 670
rect 22536 6646 22570 6662
rect 22536 654 22570 670
rect 22694 6646 22728 6662
rect 22694 654 22728 670
rect 22852 6646 22886 6662
rect 22852 654 22886 670
rect 23010 6646 23044 6662
rect 23010 654 23044 670
rect 23168 6646 23202 6662
rect 23168 654 23202 670
rect 23326 6646 23360 6662
rect 23326 654 23360 670
rect 23484 6646 23518 6662
rect 23484 654 23518 670
rect 23642 6646 23676 6662
rect 23642 654 23676 670
rect 23800 6646 23834 6662
rect 23800 654 23834 670
rect 23958 6646 23992 6662
rect 23958 654 23992 670
rect 24116 6646 24150 6662
rect 24116 654 24150 670
rect 24274 6646 24308 6662
rect 24274 654 24308 670
rect 24432 6646 24466 6662
rect 24432 654 24466 670
rect 24590 6646 24624 6662
rect 24590 654 24624 670
rect 24748 6646 24782 6662
rect 24748 654 24782 670
rect 24906 6646 24940 6662
rect 24906 654 24940 670
rect 25064 6646 25098 6662
rect 25064 654 25098 670
rect 25222 6646 25256 6662
rect 25222 654 25256 670
rect 1628 586 1644 620
rect 1712 586 1728 620
rect 1786 586 1802 620
rect 1870 586 1886 620
rect 1944 586 1960 620
rect 2028 586 2044 620
rect 2102 586 2118 620
rect 2186 586 2202 620
rect 2260 586 2276 620
rect 2344 586 2360 620
rect 2418 586 2434 620
rect 2502 586 2518 620
rect 2576 586 2592 620
rect 2660 586 2676 620
rect 2734 586 2750 620
rect 2818 586 2834 620
rect 2892 586 2908 620
rect 2976 586 2992 620
rect 3050 586 3066 620
rect 3134 586 3150 620
rect 3208 586 3224 620
rect 3292 586 3308 620
rect 3366 586 3382 620
rect 3450 586 3466 620
rect 3524 586 3540 620
rect 3608 586 3624 620
rect 3682 586 3698 620
rect 3766 586 3782 620
rect 3840 586 3856 620
rect 3924 586 3940 620
rect 3998 586 4014 620
rect 4082 586 4098 620
rect 4156 586 4172 620
rect 4240 586 4256 620
rect 4314 586 4330 620
rect 4398 586 4414 620
rect 4472 586 4488 620
rect 4556 586 4572 620
rect 4630 586 4646 620
rect 4714 586 4730 620
rect 4788 586 4804 620
rect 4872 586 4888 620
rect 4946 586 4962 620
rect 5030 586 5046 620
rect 5104 586 5120 620
rect 5188 586 5204 620
rect 5262 586 5278 620
rect 5346 586 5362 620
rect 5420 586 5436 620
rect 5504 586 5520 620
rect 5578 586 5594 620
rect 5662 586 5678 620
rect 5736 586 5752 620
rect 5820 586 5836 620
rect 5894 586 5910 620
rect 5978 586 5994 620
rect 6052 586 6068 620
rect 6136 586 6152 620
rect 6210 586 6226 620
rect 6294 586 6310 620
rect 1448 482 1482 544
rect 6456 482 6490 544
rect 1448 448 1544 482
rect 6394 448 6490 482
rect 7928 586 7944 620
rect 8012 586 8028 620
rect 8086 586 8102 620
rect 8170 586 8186 620
rect 8244 586 8260 620
rect 8328 586 8344 620
rect 8402 586 8418 620
rect 8486 586 8502 620
rect 8560 586 8576 620
rect 8644 586 8660 620
rect 8718 586 8734 620
rect 8802 586 8818 620
rect 8876 586 8892 620
rect 8960 586 8976 620
rect 9034 586 9050 620
rect 9118 586 9134 620
rect 9192 586 9208 620
rect 9276 586 9292 620
rect 9350 586 9366 620
rect 9434 586 9450 620
rect 9508 586 9524 620
rect 9592 586 9608 620
rect 9666 586 9682 620
rect 9750 586 9766 620
rect 9824 586 9840 620
rect 9908 586 9924 620
rect 9982 586 9998 620
rect 10066 586 10082 620
rect 10140 586 10156 620
rect 10224 586 10240 620
rect 10298 586 10314 620
rect 10382 586 10398 620
rect 10456 586 10472 620
rect 10540 586 10556 620
rect 10614 586 10630 620
rect 10698 586 10714 620
rect 10772 586 10788 620
rect 10856 586 10872 620
rect 10930 586 10946 620
rect 11014 586 11030 620
rect 11088 586 11104 620
rect 11172 586 11188 620
rect 11246 586 11262 620
rect 11330 586 11346 620
rect 11404 586 11420 620
rect 11488 586 11504 620
rect 11562 586 11578 620
rect 11646 586 11662 620
rect 11720 586 11736 620
rect 11804 586 11820 620
rect 11878 586 11894 620
rect 11962 586 11978 620
rect 12036 586 12052 620
rect 12120 586 12136 620
rect 12194 586 12210 620
rect 12278 586 12294 620
rect 12352 586 12368 620
rect 12436 586 12452 620
rect 12510 586 12526 620
rect 12594 586 12610 620
rect 7748 482 7782 544
rect 12756 482 12790 544
rect 7748 448 7844 482
rect 12694 448 12790 482
rect 14228 586 14244 620
rect 14312 586 14328 620
rect 14386 586 14402 620
rect 14470 586 14486 620
rect 14544 586 14560 620
rect 14628 586 14644 620
rect 14702 586 14718 620
rect 14786 586 14802 620
rect 14860 586 14876 620
rect 14944 586 14960 620
rect 15018 586 15034 620
rect 15102 586 15118 620
rect 15176 586 15192 620
rect 15260 586 15276 620
rect 15334 586 15350 620
rect 15418 586 15434 620
rect 15492 586 15508 620
rect 15576 586 15592 620
rect 15650 586 15666 620
rect 15734 586 15750 620
rect 15808 586 15824 620
rect 15892 586 15908 620
rect 15966 586 15982 620
rect 16050 586 16066 620
rect 16124 586 16140 620
rect 16208 586 16224 620
rect 16282 586 16298 620
rect 16366 586 16382 620
rect 16440 586 16456 620
rect 16524 586 16540 620
rect 16598 586 16614 620
rect 16682 586 16698 620
rect 16756 586 16772 620
rect 16840 586 16856 620
rect 16914 586 16930 620
rect 16998 586 17014 620
rect 17072 586 17088 620
rect 17156 586 17172 620
rect 17230 586 17246 620
rect 17314 586 17330 620
rect 17388 586 17404 620
rect 17472 586 17488 620
rect 17546 586 17562 620
rect 17630 586 17646 620
rect 17704 586 17720 620
rect 17788 586 17804 620
rect 17862 586 17878 620
rect 17946 586 17962 620
rect 18020 586 18036 620
rect 18104 586 18120 620
rect 18178 586 18194 620
rect 18262 586 18278 620
rect 18336 586 18352 620
rect 18420 586 18436 620
rect 18494 586 18510 620
rect 18578 586 18594 620
rect 18652 586 18668 620
rect 18736 586 18752 620
rect 18810 586 18826 620
rect 18894 586 18910 620
rect 14048 482 14082 544
rect 19056 482 19090 544
rect 14048 448 14144 482
rect 18994 448 19090 482
rect 20528 586 20544 620
rect 20612 586 20628 620
rect 20686 586 20702 620
rect 20770 586 20786 620
rect 20844 586 20860 620
rect 20928 586 20944 620
rect 21002 586 21018 620
rect 21086 586 21102 620
rect 21160 586 21176 620
rect 21244 586 21260 620
rect 21318 586 21334 620
rect 21402 586 21418 620
rect 21476 586 21492 620
rect 21560 586 21576 620
rect 21634 586 21650 620
rect 21718 586 21734 620
rect 21792 586 21808 620
rect 21876 586 21892 620
rect 21950 586 21966 620
rect 22034 586 22050 620
rect 22108 586 22124 620
rect 22192 586 22208 620
rect 22266 586 22282 620
rect 22350 586 22366 620
rect 22424 586 22440 620
rect 22508 586 22524 620
rect 22582 586 22598 620
rect 22666 586 22682 620
rect 22740 586 22756 620
rect 22824 586 22840 620
rect 22898 586 22914 620
rect 22982 586 22998 620
rect 23056 586 23072 620
rect 23140 586 23156 620
rect 23214 586 23230 620
rect 23298 586 23314 620
rect 23372 586 23388 620
rect 23456 586 23472 620
rect 23530 586 23546 620
rect 23614 586 23630 620
rect 23688 586 23704 620
rect 23772 586 23788 620
rect 23846 586 23862 620
rect 23930 586 23946 620
rect 24004 586 24020 620
rect 24088 586 24104 620
rect 24162 586 24178 620
rect 24246 586 24262 620
rect 24320 586 24336 620
rect 24404 586 24420 620
rect 24478 586 24494 620
rect 24562 586 24578 620
rect 24636 586 24652 620
rect 24720 586 24736 620
rect 24794 586 24810 620
rect 24878 586 24894 620
rect 24952 586 24968 620
rect 25036 586 25052 620
rect 25110 586 25126 620
rect 25194 586 25210 620
rect 20348 482 20382 544
rect 25356 482 25390 544
rect 20348 448 20444 482
rect 25294 448 25390 482
rect 1448 -766 1544 -732
rect 6394 -766 6490 -732
rect 1448 -828 1482 -766
rect 6456 -828 6490 -766
rect 1628 -904 1644 -870
rect 1712 -904 1728 -870
rect 1786 -904 1802 -870
rect 1870 -904 1886 -870
rect 1944 -904 1960 -870
rect 2028 -904 2044 -870
rect 2102 -904 2118 -870
rect 2186 -904 2202 -870
rect 2260 -904 2276 -870
rect 2344 -904 2360 -870
rect 2418 -904 2434 -870
rect 2502 -904 2518 -870
rect 2576 -904 2592 -870
rect 2660 -904 2676 -870
rect 2734 -904 2750 -870
rect 2818 -904 2834 -870
rect 2892 -904 2908 -870
rect 2976 -904 2992 -870
rect 3050 -904 3066 -870
rect 3134 -904 3150 -870
rect 3208 -904 3224 -870
rect 3292 -904 3308 -870
rect 3366 -904 3382 -870
rect 3450 -904 3466 -870
rect 3524 -904 3540 -870
rect 3608 -904 3624 -870
rect 3682 -904 3698 -870
rect 3766 -904 3782 -870
rect 3840 -904 3856 -870
rect 3924 -904 3940 -870
rect 3998 -904 4014 -870
rect 4082 -904 4098 -870
rect 4156 -904 4172 -870
rect 4240 -904 4256 -870
rect 4314 -904 4330 -870
rect 4398 -904 4414 -870
rect 4472 -904 4488 -870
rect 4556 -904 4572 -870
rect 4630 -904 4646 -870
rect 4714 -904 4730 -870
rect 4788 -904 4804 -870
rect 4872 -904 4888 -870
rect 4946 -904 4962 -870
rect 5030 -904 5046 -870
rect 5104 -904 5120 -870
rect 5188 -904 5204 -870
rect 5262 -904 5278 -870
rect 5346 -904 5362 -870
rect 5420 -904 5436 -870
rect 5504 -904 5520 -870
rect 5578 -904 5594 -870
rect 5662 -904 5678 -870
rect 5736 -904 5752 -870
rect 5820 -904 5836 -870
rect 5894 -904 5910 -870
rect 5978 -904 5994 -870
rect 6052 -904 6068 -870
rect 6136 -904 6152 -870
rect 6210 -904 6226 -870
rect 6294 -904 6310 -870
rect 7748 -766 7844 -732
rect 12694 -766 12790 -732
rect 7748 -828 7782 -766
rect 12756 -828 12790 -766
rect 7928 -904 7944 -870
rect 8012 -904 8028 -870
rect 8086 -904 8102 -870
rect 8170 -904 8186 -870
rect 8244 -904 8260 -870
rect 8328 -904 8344 -870
rect 8402 -904 8418 -870
rect 8486 -904 8502 -870
rect 8560 -904 8576 -870
rect 8644 -904 8660 -870
rect 8718 -904 8734 -870
rect 8802 -904 8818 -870
rect 8876 -904 8892 -870
rect 8960 -904 8976 -870
rect 9034 -904 9050 -870
rect 9118 -904 9134 -870
rect 9192 -904 9208 -870
rect 9276 -904 9292 -870
rect 9350 -904 9366 -870
rect 9434 -904 9450 -870
rect 9508 -904 9524 -870
rect 9592 -904 9608 -870
rect 9666 -904 9682 -870
rect 9750 -904 9766 -870
rect 9824 -904 9840 -870
rect 9908 -904 9924 -870
rect 9982 -904 9998 -870
rect 10066 -904 10082 -870
rect 10140 -904 10156 -870
rect 10224 -904 10240 -870
rect 10298 -904 10314 -870
rect 10382 -904 10398 -870
rect 10456 -904 10472 -870
rect 10540 -904 10556 -870
rect 10614 -904 10630 -870
rect 10698 -904 10714 -870
rect 10772 -904 10788 -870
rect 10856 -904 10872 -870
rect 10930 -904 10946 -870
rect 11014 -904 11030 -870
rect 11088 -904 11104 -870
rect 11172 -904 11188 -870
rect 11246 -904 11262 -870
rect 11330 -904 11346 -870
rect 11404 -904 11420 -870
rect 11488 -904 11504 -870
rect 11562 -904 11578 -870
rect 11646 -904 11662 -870
rect 11720 -904 11736 -870
rect 11804 -904 11820 -870
rect 11878 -904 11894 -870
rect 11962 -904 11978 -870
rect 12036 -904 12052 -870
rect 12120 -904 12136 -870
rect 12194 -904 12210 -870
rect 12278 -904 12294 -870
rect 12352 -904 12368 -870
rect 12436 -904 12452 -870
rect 12510 -904 12526 -870
rect 12594 -904 12610 -870
rect 14048 -766 14144 -732
rect 18994 -766 19090 -732
rect 14048 -828 14082 -766
rect 19056 -828 19090 -766
rect 14228 -904 14244 -870
rect 14312 -904 14328 -870
rect 14386 -904 14402 -870
rect 14470 -904 14486 -870
rect 14544 -904 14560 -870
rect 14628 -904 14644 -870
rect 14702 -904 14718 -870
rect 14786 -904 14802 -870
rect 14860 -904 14876 -870
rect 14944 -904 14960 -870
rect 15018 -904 15034 -870
rect 15102 -904 15118 -870
rect 15176 -904 15192 -870
rect 15260 -904 15276 -870
rect 15334 -904 15350 -870
rect 15418 -904 15434 -870
rect 15492 -904 15508 -870
rect 15576 -904 15592 -870
rect 15650 -904 15666 -870
rect 15734 -904 15750 -870
rect 15808 -904 15824 -870
rect 15892 -904 15908 -870
rect 15966 -904 15982 -870
rect 16050 -904 16066 -870
rect 16124 -904 16140 -870
rect 16208 -904 16224 -870
rect 16282 -904 16298 -870
rect 16366 -904 16382 -870
rect 16440 -904 16456 -870
rect 16524 -904 16540 -870
rect 16598 -904 16614 -870
rect 16682 -904 16698 -870
rect 16756 -904 16772 -870
rect 16840 -904 16856 -870
rect 16914 -904 16930 -870
rect 16998 -904 17014 -870
rect 17072 -904 17088 -870
rect 17156 -904 17172 -870
rect 17230 -904 17246 -870
rect 17314 -904 17330 -870
rect 17388 -904 17404 -870
rect 17472 -904 17488 -870
rect 17546 -904 17562 -870
rect 17630 -904 17646 -870
rect 17704 -904 17720 -870
rect 17788 -904 17804 -870
rect 17862 -904 17878 -870
rect 17946 -904 17962 -870
rect 18020 -904 18036 -870
rect 18104 -904 18120 -870
rect 18178 -904 18194 -870
rect 18262 -904 18278 -870
rect 18336 -904 18352 -870
rect 18420 -904 18436 -870
rect 18494 -904 18510 -870
rect 18578 -904 18594 -870
rect 18652 -904 18668 -870
rect 18736 -904 18752 -870
rect 18810 -904 18826 -870
rect 18894 -904 18910 -870
rect 20348 -766 20444 -732
rect 25294 -766 25390 -732
rect 20348 -828 20382 -766
rect 25356 -828 25390 -766
rect 20528 -904 20544 -870
rect 20612 -904 20628 -870
rect 20686 -904 20702 -870
rect 20770 -904 20786 -870
rect 20844 -904 20860 -870
rect 20928 -904 20944 -870
rect 21002 -904 21018 -870
rect 21086 -904 21102 -870
rect 21160 -904 21176 -870
rect 21244 -904 21260 -870
rect 21318 -904 21334 -870
rect 21402 -904 21418 -870
rect 21476 -904 21492 -870
rect 21560 -904 21576 -870
rect 21634 -904 21650 -870
rect 21718 -904 21734 -870
rect 21792 -904 21808 -870
rect 21876 -904 21892 -870
rect 21950 -904 21966 -870
rect 22034 -904 22050 -870
rect 22108 -904 22124 -870
rect 22192 -904 22208 -870
rect 22266 -904 22282 -870
rect 22350 -904 22366 -870
rect 22424 -904 22440 -870
rect 22508 -904 22524 -870
rect 22582 -904 22598 -870
rect 22666 -904 22682 -870
rect 22740 -904 22756 -870
rect 22824 -904 22840 -870
rect 22898 -904 22914 -870
rect 22982 -904 22998 -870
rect 23056 -904 23072 -870
rect 23140 -904 23156 -870
rect 23214 -904 23230 -870
rect 23298 -904 23314 -870
rect 23372 -904 23388 -870
rect 23456 -904 23472 -870
rect 23530 -904 23546 -870
rect 23614 -904 23630 -870
rect 23688 -904 23704 -870
rect 23772 -904 23788 -870
rect 23846 -904 23862 -870
rect 23930 -904 23946 -870
rect 24004 -904 24020 -870
rect 24088 -904 24104 -870
rect 24162 -904 24178 -870
rect 24246 -904 24262 -870
rect 24320 -904 24336 -870
rect 24404 -904 24420 -870
rect 24478 -904 24494 -870
rect 24562 -904 24578 -870
rect 24636 -904 24652 -870
rect 24720 -904 24736 -870
rect 24794 -904 24810 -870
rect 24878 -904 24894 -870
rect 24952 -904 24968 -870
rect 25036 -904 25052 -870
rect 25110 -904 25126 -870
rect 25194 -904 25210 -870
rect 1582 -954 1616 -938
rect 1582 -6946 1616 -6930
rect 1740 -954 1774 -938
rect 1740 -6946 1774 -6930
rect 1898 -954 1932 -938
rect 1898 -6946 1932 -6930
rect 2056 -954 2090 -938
rect 2056 -6946 2090 -6930
rect 2214 -954 2248 -938
rect 2214 -6946 2248 -6930
rect 2372 -954 2406 -938
rect 2372 -6946 2406 -6930
rect 2530 -954 2564 -938
rect 2530 -6946 2564 -6930
rect 2688 -954 2722 -938
rect 2688 -6946 2722 -6930
rect 2846 -954 2880 -938
rect 2846 -6946 2880 -6930
rect 3004 -954 3038 -938
rect 3004 -6946 3038 -6930
rect 3162 -954 3196 -938
rect 3162 -6946 3196 -6930
rect 3320 -954 3354 -938
rect 3320 -6946 3354 -6930
rect 3478 -954 3512 -938
rect 3478 -6946 3512 -6930
rect 3636 -954 3670 -938
rect 3636 -6946 3670 -6930
rect 3794 -954 3828 -938
rect 3794 -6946 3828 -6930
rect 3952 -954 3986 -938
rect 3952 -6946 3986 -6930
rect 4110 -954 4144 -938
rect 4110 -6946 4144 -6930
rect 4268 -954 4302 -938
rect 4268 -6946 4302 -6930
rect 4426 -954 4460 -938
rect 4426 -6946 4460 -6930
rect 4584 -954 4618 -938
rect 4584 -6946 4618 -6930
rect 4742 -954 4776 -938
rect 4742 -6946 4776 -6930
rect 4900 -954 4934 -938
rect 4900 -6946 4934 -6930
rect 5058 -954 5092 -938
rect 5058 -6946 5092 -6930
rect 5216 -954 5250 -938
rect 5216 -6946 5250 -6930
rect 5374 -954 5408 -938
rect 5374 -6946 5408 -6930
rect 5532 -954 5566 -938
rect 5532 -6946 5566 -6930
rect 5690 -954 5724 -938
rect 5690 -6946 5724 -6930
rect 5848 -954 5882 -938
rect 5848 -6946 5882 -6930
rect 6006 -954 6040 -938
rect 6006 -6946 6040 -6930
rect 6164 -954 6198 -938
rect 6164 -6946 6198 -6930
rect 6322 -954 6356 -938
rect 6322 -6946 6356 -6930
rect 7882 -954 7916 -938
rect 7882 -6946 7916 -6930
rect 8040 -954 8074 -938
rect 8040 -6946 8074 -6930
rect 8198 -954 8232 -938
rect 8198 -6946 8232 -6930
rect 8356 -954 8390 -938
rect 8356 -6946 8390 -6930
rect 8514 -954 8548 -938
rect 8514 -6946 8548 -6930
rect 8672 -954 8706 -938
rect 8672 -6946 8706 -6930
rect 8830 -954 8864 -938
rect 8830 -6946 8864 -6930
rect 8988 -954 9022 -938
rect 8988 -6946 9022 -6930
rect 9146 -954 9180 -938
rect 9146 -6946 9180 -6930
rect 9304 -954 9338 -938
rect 9304 -6946 9338 -6930
rect 9462 -954 9496 -938
rect 9462 -6946 9496 -6930
rect 9620 -954 9654 -938
rect 9620 -6946 9654 -6930
rect 9778 -954 9812 -938
rect 9778 -6946 9812 -6930
rect 9936 -954 9970 -938
rect 9936 -6946 9970 -6930
rect 10094 -954 10128 -938
rect 10094 -6946 10128 -6930
rect 10252 -954 10286 -938
rect 10252 -6946 10286 -6930
rect 10410 -954 10444 -938
rect 10410 -6946 10444 -6930
rect 10568 -954 10602 -938
rect 10568 -6946 10602 -6930
rect 10726 -954 10760 -938
rect 10726 -6946 10760 -6930
rect 10884 -954 10918 -938
rect 10884 -6946 10918 -6930
rect 11042 -954 11076 -938
rect 11042 -6946 11076 -6930
rect 11200 -954 11234 -938
rect 11200 -6946 11234 -6930
rect 11358 -954 11392 -938
rect 11358 -6946 11392 -6930
rect 11516 -954 11550 -938
rect 11516 -6946 11550 -6930
rect 11674 -954 11708 -938
rect 11674 -6946 11708 -6930
rect 11832 -954 11866 -938
rect 11832 -6946 11866 -6930
rect 11990 -954 12024 -938
rect 11990 -6946 12024 -6930
rect 12148 -954 12182 -938
rect 12148 -6946 12182 -6930
rect 12306 -954 12340 -938
rect 12306 -6946 12340 -6930
rect 12464 -954 12498 -938
rect 12464 -6946 12498 -6930
rect 12622 -954 12656 -938
rect 12622 -6946 12656 -6930
rect 14182 -954 14216 -938
rect 14182 -6946 14216 -6930
rect 14340 -954 14374 -938
rect 14340 -6946 14374 -6930
rect 14498 -954 14532 -938
rect 14498 -6946 14532 -6930
rect 14656 -954 14690 -938
rect 14656 -6946 14690 -6930
rect 14814 -954 14848 -938
rect 14814 -6946 14848 -6930
rect 14972 -954 15006 -938
rect 14972 -6946 15006 -6930
rect 15130 -954 15164 -938
rect 15130 -6946 15164 -6930
rect 15288 -954 15322 -938
rect 15288 -6946 15322 -6930
rect 15446 -954 15480 -938
rect 15446 -6946 15480 -6930
rect 15604 -954 15638 -938
rect 15604 -6946 15638 -6930
rect 15762 -954 15796 -938
rect 15762 -6946 15796 -6930
rect 15920 -954 15954 -938
rect 15920 -6946 15954 -6930
rect 16078 -954 16112 -938
rect 16078 -6946 16112 -6930
rect 16236 -954 16270 -938
rect 16236 -6946 16270 -6930
rect 16394 -954 16428 -938
rect 16394 -6946 16428 -6930
rect 16552 -954 16586 -938
rect 16552 -6946 16586 -6930
rect 16710 -954 16744 -938
rect 16710 -6946 16744 -6930
rect 16868 -954 16902 -938
rect 16868 -6946 16902 -6930
rect 17026 -954 17060 -938
rect 17026 -6946 17060 -6930
rect 17184 -954 17218 -938
rect 17184 -6946 17218 -6930
rect 17342 -954 17376 -938
rect 17342 -6946 17376 -6930
rect 17500 -954 17534 -938
rect 17500 -6946 17534 -6930
rect 17658 -954 17692 -938
rect 17658 -6946 17692 -6930
rect 17816 -954 17850 -938
rect 17816 -6946 17850 -6930
rect 17974 -954 18008 -938
rect 17974 -6946 18008 -6930
rect 18132 -954 18166 -938
rect 18132 -6946 18166 -6930
rect 18290 -954 18324 -938
rect 18290 -6946 18324 -6930
rect 18448 -954 18482 -938
rect 18448 -6946 18482 -6930
rect 18606 -954 18640 -938
rect 18606 -6946 18640 -6930
rect 18764 -954 18798 -938
rect 18764 -6946 18798 -6930
rect 18922 -954 18956 -938
rect 18922 -6946 18956 -6930
rect 20482 -954 20516 -938
rect 20482 -6946 20516 -6930
rect 20640 -954 20674 -938
rect 20640 -6946 20674 -6930
rect 20798 -954 20832 -938
rect 20798 -6946 20832 -6930
rect 20956 -954 20990 -938
rect 20956 -6946 20990 -6930
rect 21114 -954 21148 -938
rect 21114 -6946 21148 -6930
rect 21272 -954 21306 -938
rect 21272 -6946 21306 -6930
rect 21430 -954 21464 -938
rect 21430 -6946 21464 -6930
rect 21588 -954 21622 -938
rect 21588 -6946 21622 -6930
rect 21746 -954 21780 -938
rect 21746 -6946 21780 -6930
rect 21904 -954 21938 -938
rect 21904 -6946 21938 -6930
rect 22062 -954 22096 -938
rect 22062 -6946 22096 -6930
rect 22220 -954 22254 -938
rect 22220 -6946 22254 -6930
rect 22378 -954 22412 -938
rect 22378 -6946 22412 -6930
rect 22536 -954 22570 -938
rect 22536 -6946 22570 -6930
rect 22694 -954 22728 -938
rect 22694 -6946 22728 -6930
rect 22852 -954 22886 -938
rect 22852 -6946 22886 -6930
rect 23010 -954 23044 -938
rect 23010 -6946 23044 -6930
rect 23168 -954 23202 -938
rect 23168 -6946 23202 -6930
rect 23326 -954 23360 -938
rect 23326 -6946 23360 -6930
rect 23484 -954 23518 -938
rect 23484 -6946 23518 -6930
rect 23642 -954 23676 -938
rect 23642 -6946 23676 -6930
rect 23800 -954 23834 -938
rect 23800 -6946 23834 -6930
rect 23958 -954 23992 -938
rect 23958 -6946 23992 -6930
rect 24116 -954 24150 -938
rect 24116 -6946 24150 -6930
rect 24274 -954 24308 -938
rect 24274 -6946 24308 -6930
rect 24432 -954 24466 -938
rect 24432 -6946 24466 -6930
rect 24590 -954 24624 -938
rect 24590 -6946 24624 -6930
rect 24748 -954 24782 -938
rect 24748 -6946 24782 -6930
rect 24906 -954 24940 -938
rect 24906 -6946 24940 -6930
rect 25064 -954 25098 -938
rect 25064 -6946 25098 -6930
rect 25222 -954 25256 -938
rect 25222 -6946 25256 -6930
rect 1628 -7014 1644 -6980
rect 1712 -7014 1728 -6980
rect 1786 -7014 1802 -6980
rect 1870 -7014 1886 -6980
rect 1944 -7014 1960 -6980
rect 2028 -7014 2044 -6980
rect 2102 -7014 2118 -6980
rect 2186 -7014 2202 -6980
rect 2260 -7014 2276 -6980
rect 2344 -7014 2360 -6980
rect 2418 -7014 2434 -6980
rect 2502 -7014 2518 -6980
rect 2576 -7014 2592 -6980
rect 2660 -7014 2676 -6980
rect 2734 -7014 2750 -6980
rect 2818 -7014 2834 -6980
rect 2892 -7014 2908 -6980
rect 2976 -7014 2992 -6980
rect 3050 -7014 3066 -6980
rect 3134 -7014 3150 -6980
rect 3208 -7014 3224 -6980
rect 3292 -7014 3308 -6980
rect 3366 -7014 3382 -6980
rect 3450 -7014 3466 -6980
rect 3524 -7014 3540 -6980
rect 3608 -7014 3624 -6980
rect 3682 -7014 3698 -6980
rect 3766 -7014 3782 -6980
rect 3840 -7014 3856 -6980
rect 3924 -7014 3940 -6980
rect 3998 -7014 4014 -6980
rect 4082 -7014 4098 -6980
rect 4156 -7014 4172 -6980
rect 4240 -7014 4256 -6980
rect 4314 -7014 4330 -6980
rect 4398 -7014 4414 -6980
rect 4472 -7014 4488 -6980
rect 4556 -7014 4572 -6980
rect 4630 -7014 4646 -6980
rect 4714 -7014 4730 -6980
rect 4788 -7014 4804 -6980
rect 4872 -7014 4888 -6980
rect 4946 -7014 4962 -6980
rect 5030 -7014 5046 -6980
rect 5104 -7014 5120 -6980
rect 5188 -7014 5204 -6980
rect 5262 -7014 5278 -6980
rect 5346 -7014 5362 -6980
rect 5420 -7014 5436 -6980
rect 5504 -7014 5520 -6980
rect 5578 -7014 5594 -6980
rect 5662 -7014 5678 -6980
rect 5736 -7014 5752 -6980
rect 5820 -7014 5836 -6980
rect 5894 -7014 5910 -6980
rect 5978 -7014 5994 -6980
rect 6052 -7014 6068 -6980
rect 6136 -7014 6152 -6980
rect 6210 -7014 6226 -6980
rect 6294 -7014 6310 -6980
rect 1448 -7118 1482 -7056
rect 6456 -7118 6490 -7056
rect 1448 -7152 1544 -7118
rect 6394 -7152 6490 -7118
rect 7928 -7014 7944 -6980
rect 8012 -7014 8028 -6980
rect 8086 -7014 8102 -6980
rect 8170 -7014 8186 -6980
rect 8244 -7014 8260 -6980
rect 8328 -7014 8344 -6980
rect 8402 -7014 8418 -6980
rect 8486 -7014 8502 -6980
rect 8560 -7014 8576 -6980
rect 8644 -7014 8660 -6980
rect 8718 -7014 8734 -6980
rect 8802 -7014 8818 -6980
rect 8876 -7014 8892 -6980
rect 8960 -7014 8976 -6980
rect 9034 -7014 9050 -6980
rect 9118 -7014 9134 -6980
rect 9192 -7014 9208 -6980
rect 9276 -7014 9292 -6980
rect 9350 -7014 9366 -6980
rect 9434 -7014 9450 -6980
rect 9508 -7014 9524 -6980
rect 9592 -7014 9608 -6980
rect 9666 -7014 9682 -6980
rect 9750 -7014 9766 -6980
rect 9824 -7014 9840 -6980
rect 9908 -7014 9924 -6980
rect 9982 -7014 9998 -6980
rect 10066 -7014 10082 -6980
rect 10140 -7014 10156 -6980
rect 10224 -7014 10240 -6980
rect 10298 -7014 10314 -6980
rect 10382 -7014 10398 -6980
rect 10456 -7014 10472 -6980
rect 10540 -7014 10556 -6980
rect 10614 -7014 10630 -6980
rect 10698 -7014 10714 -6980
rect 10772 -7014 10788 -6980
rect 10856 -7014 10872 -6980
rect 10930 -7014 10946 -6980
rect 11014 -7014 11030 -6980
rect 11088 -7014 11104 -6980
rect 11172 -7014 11188 -6980
rect 11246 -7014 11262 -6980
rect 11330 -7014 11346 -6980
rect 11404 -7014 11420 -6980
rect 11488 -7014 11504 -6980
rect 11562 -7014 11578 -6980
rect 11646 -7014 11662 -6980
rect 11720 -7014 11736 -6980
rect 11804 -7014 11820 -6980
rect 11878 -7014 11894 -6980
rect 11962 -7014 11978 -6980
rect 12036 -7014 12052 -6980
rect 12120 -7014 12136 -6980
rect 12194 -7014 12210 -6980
rect 12278 -7014 12294 -6980
rect 12352 -7014 12368 -6980
rect 12436 -7014 12452 -6980
rect 12510 -7014 12526 -6980
rect 12594 -7014 12610 -6980
rect 7748 -7118 7782 -7056
rect 12756 -7118 12790 -7056
rect 7748 -7152 7844 -7118
rect 12694 -7152 12790 -7118
rect 14228 -7014 14244 -6980
rect 14312 -7014 14328 -6980
rect 14386 -7014 14402 -6980
rect 14470 -7014 14486 -6980
rect 14544 -7014 14560 -6980
rect 14628 -7014 14644 -6980
rect 14702 -7014 14718 -6980
rect 14786 -7014 14802 -6980
rect 14860 -7014 14876 -6980
rect 14944 -7014 14960 -6980
rect 15018 -7014 15034 -6980
rect 15102 -7014 15118 -6980
rect 15176 -7014 15192 -6980
rect 15260 -7014 15276 -6980
rect 15334 -7014 15350 -6980
rect 15418 -7014 15434 -6980
rect 15492 -7014 15508 -6980
rect 15576 -7014 15592 -6980
rect 15650 -7014 15666 -6980
rect 15734 -7014 15750 -6980
rect 15808 -7014 15824 -6980
rect 15892 -7014 15908 -6980
rect 15966 -7014 15982 -6980
rect 16050 -7014 16066 -6980
rect 16124 -7014 16140 -6980
rect 16208 -7014 16224 -6980
rect 16282 -7014 16298 -6980
rect 16366 -7014 16382 -6980
rect 16440 -7014 16456 -6980
rect 16524 -7014 16540 -6980
rect 16598 -7014 16614 -6980
rect 16682 -7014 16698 -6980
rect 16756 -7014 16772 -6980
rect 16840 -7014 16856 -6980
rect 16914 -7014 16930 -6980
rect 16998 -7014 17014 -6980
rect 17072 -7014 17088 -6980
rect 17156 -7014 17172 -6980
rect 17230 -7014 17246 -6980
rect 17314 -7014 17330 -6980
rect 17388 -7014 17404 -6980
rect 17472 -7014 17488 -6980
rect 17546 -7014 17562 -6980
rect 17630 -7014 17646 -6980
rect 17704 -7014 17720 -6980
rect 17788 -7014 17804 -6980
rect 17862 -7014 17878 -6980
rect 17946 -7014 17962 -6980
rect 18020 -7014 18036 -6980
rect 18104 -7014 18120 -6980
rect 18178 -7014 18194 -6980
rect 18262 -7014 18278 -6980
rect 18336 -7014 18352 -6980
rect 18420 -7014 18436 -6980
rect 18494 -7014 18510 -6980
rect 18578 -7014 18594 -6980
rect 18652 -7014 18668 -6980
rect 18736 -7014 18752 -6980
rect 18810 -7014 18826 -6980
rect 18894 -7014 18910 -6980
rect 14048 -7118 14082 -7056
rect 19056 -7118 19090 -7056
rect 14048 -7152 14144 -7118
rect 18994 -7152 19090 -7118
rect 20528 -7014 20544 -6980
rect 20612 -7014 20628 -6980
rect 20686 -7014 20702 -6980
rect 20770 -7014 20786 -6980
rect 20844 -7014 20860 -6980
rect 20928 -7014 20944 -6980
rect 21002 -7014 21018 -6980
rect 21086 -7014 21102 -6980
rect 21160 -7014 21176 -6980
rect 21244 -7014 21260 -6980
rect 21318 -7014 21334 -6980
rect 21402 -7014 21418 -6980
rect 21476 -7014 21492 -6980
rect 21560 -7014 21576 -6980
rect 21634 -7014 21650 -6980
rect 21718 -7014 21734 -6980
rect 21792 -7014 21808 -6980
rect 21876 -7014 21892 -6980
rect 21950 -7014 21966 -6980
rect 22034 -7014 22050 -6980
rect 22108 -7014 22124 -6980
rect 22192 -7014 22208 -6980
rect 22266 -7014 22282 -6980
rect 22350 -7014 22366 -6980
rect 22424 -7014 22440 -6980
rect 22508 -7014 22524 -6980
rect 22582 -7014 22598 -6980
rect 22666 -7014 22682 -6980
rect 22740 -7014 22756 -6980
rect 22824 -7014 22840 -6980
rect 22898 -7014 22914 -6980
rect 22982 -7014 22998 -6980
rect 23056 -7014 23072 -6980
rect 23140 -7014 23156 -6980
rect 23214 -7014 23230 -6980
rect 23298 -7014 23314 -6980
rect 23372 -7014 23388 -6980
rect 23456 -7014 23472 -6980
rect 23530 -7014 23546 -6980
rect 23614 -7014 23630 -6980
rect 23688 -7014 23704 -6980
rect 23772 -7014 23788 -6980
rect 23846 -7014 23862 -6980
rect 23930 -7014 23946 -6980
rect 24004 -7014 24020 -6980
rect 24088 -7014 24104 -6980
rect 24162 -7014 24178 -6980
rect 24246 -7014 24262 -6980
rect 24320 -7014 24336 -6980
rect 24404 -7014 24420 -6980
rect 24478 -7014 24494 -6980
rect 24562 -7014 24578 -6980
rect 24636 -7014 24652 -6980
rect 24720 -7014 24736 -6980
rect 24794 -7014 24810 -6980
rect 24878 -7014 24894 -6980
rect 24952 -7014 24968 -6980
rect 25036 -7014 25052 -6980
rect 25110 -7014 25126 -6980
rect 25194 -7014 25210 -6980
rect 20348 -7118 20382 -7056
rect 25356 -7118 25390 -7056
rect 20348 -7152 20444 -7118
rect 25294 -7152 25390 -7118
<< viali >>
rect 1636 6868 6359 6870
rect 7936 6868 12659 6870
rect 14236 6868 18959 6870
rect 20536 6868 25259 6870
rect 1636 6834 6359 6868
rect 1636 6832 6359 6834
rect 1644 6696 1712 6730
rect 1802 6696 1870 6730
rect 1960 6696 2028 6730
rect 2118 6696 2186 6730
rect 2276 6696 2344 6730
rect 2434 6696 2502 6730
rect 2592 6696 2660 6730
rect 2750 6696 2818 6730
rect 2908 6696 2976 6730
rect 3066 6696 3134 6730
rect 3224 6696 3292 6730
rect 3382 6696 3450 6730
rect 3540 6696 3608 6730
rect 3698 6696 3766 6730
rect 3856 6696 3924 6730
rect 4014 6696 4082 6730
rect 4172 6696 4240 6730
rect 4330 6696 4398 6730
rect 4488 6696 4556 6730
rect 4646 6696 4714 6730
rect 4804 6696 4872 6730
rect 4962 6696 5030 6730
rect 5120 6696 5188 6730
rect 5278 6696 5346 6730
rect 5436 6696 5504 6730
rect 5594 6696 5662 6730
rect 5752 6696 5820 6730
rect 5910 6696 5978 6730
rect 6068 6696 6136 6730
rect 6226 6696 6294 6730
rect 7936 6834 12659 6868
rect 7936 6832 12659 6834
rect 7944 6696 8012 6730
rect 8102 6696 8170 6730
rect 8260 6696 8328 6730
rect 8418 6696 8486 6730
rect 8576 6696 8644 6730
rect 8734 6696 8802 6730
rect 8892 6696 8960 6730
rect 9050 6696 9118 6730
rect 9208 6696 9276 6730
rect 9366 6696 9434 6730
rect 9524 6696 9592 6730
rect 9682 6696 9750 6730
rect 9840 6696 9908 6730
rect 9998 6696 10066 6730
rect 10156 6696 10224 6730
rect 10314 6696 10382 6730
rect 10472 6696 10540 6730
rect 10630 6696 10698 6730
rect 10788 6696 10856 6730
rect 10946 6696 11014 6730
rect 11104 6696 11172 6730
rect 11262 6696 11330 6730
rect 11420 6696 11488 6730
rect 11578 6696 11646 6730
rect 11736 6696 11804 6730
rect 11894 6696 11962 6730
rect 12052 6696 12120 6730
rect 12210 6696 12278 6730
rect 12368 6696 12436 6730
rect 12526 6696 12594 6730
rect 14236 6834 18959 6868
rect 14236 6832 18959 6834
rect 14244 6696 14312 6730
rect 14402 6696 14470 6730
rect 14560 6696 14628 6730
rect 14718 6696 14786 6730
rect 14876 6696 14944 6730
rect 15034 6696 15102 6730
rect 15192 6696 15260 6730
rect 15350 6696 15418 6730
rect 15508 6696 15576 6730
rect 15666 6696 15734 6730
rect 15824 6696 15892 6730
rect 15982 6696 16050 6730
rect 16140 6696 16208 6730
rect 16298 6696 16366 6730
rect 16456 6696 16524 6730
rect 16614 6696 16682 6730
rect 16772 6696 16840 6730
rect 16930 6696 16998 6730
rect 17088 6696 17156 6730
rect 17246 6696 17314 6730
rect 17404 6696 17472 6730
rect 17562 6696 17630 6730
rect 17720 6696 17788 6730
rect 17878 6696 17946 6730
rect 18036 6696 18104 6730
rect 18194 6696 18262 6730
rect 18352 6696 18420 6730
rect 18510 6696 18578 6730
rect 18668 6696 18736 6730
rect 18826 6696 18894 6730
rect 20536 6834 25259 6868
rect 20536 6832 25259 6834
rect 20544 6696 20612 6730
rect 20702 6696 20770 6730
rect 20860 6696 20928 6730
rect 21018 6696 21086 6730
rect 21176 6696 21244 6730
rect 21334 6696 21402 6730
rect 21492 6696 21560 6730
rect 21650 6696 21718 6730
rect 21808 6696 21876 6730
rect 21966 6696 22034 6730
rect 22124 6696 22192 6730
rect 22282 6696 22350 6730
rect 22440 6696 22508 6730
rect 22598 6696 22666 6730
rect 22756 6696 22824 6730
rect 22914 6696 22982 6730
rect 23072 6696 23140 6730
rect 23230 6696 23298 6730
rect 23388 6696 23456 6730
rect 23546 6696 23614 6730
rect 23704 6696 23772 6730
rect 23862 6696 23930 6730
rect 24020 6696 24088 6730
rect 24178 6696 24246 6730
rect 24336 6696 24404 6730
rect 24494 6696 24562 6730
rect 24652 6696 24720 6730
rect 24810 6696 24878 6730
rect 24968 6696 25036 6730
rect 25126 6696 25194 6730
rect 1446 636 1448 6680
rect 1448 636 1482 6680
rect 1482 636 1484 6680
rect 1582 670 1616 6646
rect 1740 670 1774 6646
rect 1898 670 1932 6646
rect 2056 670 2090 6646
rect 2214 670 2248 6646
rect 2372 670 2406 6646
rect 2530 670 2564 6646
rect 2688 670 2722 6646
rect 2846 670 2880 6646
rect 3004 670 3038 6646
rect 3162 670 3196 6646
rect 3320 670 3354 6646
rect 3478 670 3512 6646
rect 3636 670 3670 6646
rect 3794 670 3828 6646
rect 3952 670 3986 6646
rect 4110 670 4144 6646
rect 4268 670 4302 6646
rect 4426 670 4460 6646
rect 4584 670 4618 6646
rect 4742 670 4776 6646
rect 4900 670 4934 6646
rect 5058 670 5092 6646
rect 5216 670 5250 6646
rect 5374 670 5408 6646
rect 5532 670 5566 6646
rect 5690 670 5724 6646
rect 5848 670 5882 6646
rect 6006 670 6040 6646
rect 6164 670 6198 6646
rect 6322 670 6356 6646
rect 6454 636 6456 6680
rect 6456 636 6490 6680
rect 6490 636 6492 6680
rect 7746 636 7748 6680
rect 7748 636 7782 6680
rect 7782 636 7784 6680
rect 7882 670 7916 6646
rect 8040 670 8074 6646
rect 8198 670 8232 6646
rect 8356 670 8390 6646
rect 8514 670 8548 6646
rect 8672 670 8706 6646
rect 8830 670 8864 6646
rect 8988 670 9022 6646
rect 9146 670 9180 6646
rect 9304 670 9338 6646
rect 9462 670 9496 6646
rect 9620 670 9654 6646
rect 9778 670 9812 6646
rect 9936 670 9970 6646
rect 10094 670 10128 6646
rect 10252 670 10286 6646
rect 10410 670 10444 6646
rect 10568 670 10602 6646
rect 10726 670 10760 6646
rect 10884 670 10918 6646
rect 11042 670 11076 6646
rect 11200 670 11234 6646
rect 11358 670 11392 6646
rect 11516 670 11550 6646
rect 11674 670 11708 6646
rect 11832 670 11866 6646
rect 11990 670 12024 6646
rect 12148 670 12182 6646
rect 12306 670 12340 6646
rect 12464 670 12498 6646
rect 12622 670 12656 6646
rect 12754 636 12756 6680
rect 12756 636 12790 6680
rect 12790 636 12792 6680
rect 14046 636 14048 6680
rect 14048 636 14082 6680
rect 14082 636 14084 6680
rect 14182 670 14216 6646
rect 14340 670 14374 6646
rect 14498 670 14532 6646
rect 14656 670 14690 6646
rect 14814 670 14848 6646
rect 14972 670 15006 6646
rect 15130 670 15164 6646
rect 15288 670 15322 6646
rect 15446 670 15480 6646
rect 15604 670 15638 6646
rect 15762 670 15796 6646
rect 15920 670 15954 6646
rect 16078 670 16112 6646
rect 16236 670 16270 6646
rect 16394 670 16428 6646
rect 16552 670 16586 6646
rect 16710 670 16744 6646
rect 16868 670 16902 6646
rect 17026 670 17060 6646
rect 17184 670 17218 6646
rect 17342 670 17376 6646
rect 17500 670 17534 6646
rect 17658 670 17692 6646
rect 17816 670 17850 6646
rect 17974 670 18008 6646
rect 18132 670 18166 6646
rect 18290 670 18324 6646
rect 18448 670 18482 6646
rect 18606 670 18640 6646
rect 18764 670 18798 6646
rect 18922 670 18956 6646
rect 19054 636 19056 6680
rect 19056 636 19090 6680
rect 19090 636 19092 6680
rect 20346 636 20348 6680
rect 20348 636 20382 6680
rect 20382 636 20384 6680
rect 20482 670 20516 6646
rect 20640 670 20674 6646
rect 20798 670 20832 6646
rect 20956 670 20990 6646
rect 21114 670 21148 6646
rect 21272 670 21306 6646
rect 21430 670 21464 6646
rect 21588 670 21622 6646
rect 21746 670 21780 6646
rect 21904 670 21938 6646
rect 22062 670 22096 6646
rect 22220 670 22254 6646
rect 22378 670 22412 6646
rect 22536 670 22570 6646
rect 22694 670 22728 6646
rect 22852 670 22886 6646
rect 23010 670 23044 6646
rect 23168 670 23202 6646
rect 23326 670 23360 6646
rect 23484 670 23518 6646
rect 23642 670 23676 6646
rect 23800 670 23834 6646
rect 23958 670 23992 6646
rect 24116 670 24150 6646
rect 24274 670 24308 6646
rect 24432 670 24466 6646
rect 24590 670 24624 6646
rect 24748 670 24782 6646
rect 24906 670 24940 6646
rect 25064 670 25098 6646
rect 25222 670 25256 6646
rect 25354 636 25356 6680
rect 25356 636 25390 6680
rect 25390 636 25392 6680
rect 1644 586 1712 620
rect 1802 586 1870 620
rect 1960 586 2028 620
rect 2118 586 2186 620
rect 2276 586 2344 620
rect 2434 586 2502 620
rect 2592 586 2660 620
rect 2750 586 2818 620
rect 2908 586 2976 620
rect 3066 586 3134 620
rect 3224 586 3292 620
rect 3382 586 3450 620
rect 3540 586 3608 620
rect 3698 586 3766 620
rect 3856 586 3924 620
rect 4014 586 4082 620
rect 4172 586 4240 620
rect 4330 586 4398 620
rect 4488 586 4556 620
rect 4646 586 4714 620
rect 4804 586 4872 620
rect 4962 586 5030 620
rect 5120 586 5188 620
rect 5278 586 5346 620
rect 5436 586 5504 620
rect 5594 586 5662 620
rect 5752 586 5820 620
rect 5910 586 5978 620
rect 6068 586 6136 620
rect 6226 586 6294 620
rect 1636 482 6302 484
rect 1636 448 6302 482
rect 7944 586 8012 620
rect 8102 586 8170 620
rect 8260 586 8328 620
rect 8418 586 8486 620
rect 8576 586 8644 620
rect 8734 586 8802 620
rect 8892 586 8960 620
rect 9050 586 9118 620
rect 9208 586 9276 620
rect 9366 586 9434 620
rect 9524 586 9592 620
rect 9682 586 9750 620
rect 9840 586 9908 620
rect 9998 586 10066 620
rect 10156 586 10224 620
rect 10314 586 10382 620
rect 10472 586 10540 620
rect 10630 586 10698 620
rect 10788 586 10856 620
rect 10946 586 11014 620
rect 11104 586 11172 620
rect 11262 586 11330 620
rect 11420 586 11488 620
rect 11578 586 11646 620
rect 11736 586 11804 620
rect 11894 586 11962 620
rect 12052 586 12120 620
rect 12210 586 12278 620
rect 12368 586 12436 620
rect 12526 586 12594 620
rect 7936 482 12602 484
rect 7936 448 12602 482
rect 14244 586 14312 620
rect 14402 586 14470 620
rect 14560 586 14628 620
rect 14718 586 14786 620
rect 14876 586 14944 620
rect 15034 586 15102 620
rect 15192 586 15260 620
rect 15350 586 15418 620
rect 15508 586 15576 620
rect 15666 586 15734 620
rect 15824 586 15892 620
rect 15982 586 16050 620
rect 16140 586 16208 620
rect 16298 586 16366 620
rect 16456 586 16524 620
rect 16614 586 16682 620
rect 16772 586 16840 620
rect 16930 586 16998 620
rect 17088 586 17156 620
rect 17246 586 17314 620
rect 17404 586 17472 620
rect 17562 586 17630 620
rect 17720 586 17788 620
rect 17878 586 17946 620
rect 18036 586 18104 620
rect 18194 586 18262 620
rect 18352 586 18420 620
rect 18510 586 18578 620
rect 18668 586 18736 620
rect 18826 586 18894 620
rect 14236 482 18902 484
rect 14236 448 18902 482
rect 20544 586 20612 620
rect 20702 586 20770 620
rect 20860 586 20928 620
rect 21018 586 21086 620
rect 21176 586 21244 620
rect 21334 586 21402 620
rect 21492 586 21560 620
rect 21650 586 21718 620
rect 21808 586 21876 620
rect 21966 586 22034 620
rect 22124 586 22192 620
rect 22282 586 22350 620
rect 22440 586 22508 620
rect 22598 586 22666 620
rect 22756 586 22824 620
rect 22914 586 22982 620
rect 23072 586 23140 620
rect 23230 586 23298 620
rect 23388 586 23456 620
rect 23546 586 23614 620
rect 23704 586 23772 620
rect 23862 586 23930 620
rect 24020 586 24088 620
rect 24178 586 24246 620
rect 24336 586 24404 620
rect 24494 586 24562 620
rect 24652 586 24720 620
rect 24810 586 24878 620
rect 24968 586 25036 620
rect 25126 586 25194 620
rect 20536 482 25202 484
rect 20536 448 25202 482
rect 1636 446 6302 448
rect 7936 446 12602 448
rect 14236 446 18902 448
rect 20536 446 25202 448
rect 1636 -732 6359 -730
rect 7936 -732 12659 -730
rect 14236 -732 18959 -730
rect 20536 -732 25259 -730
rect 1636 -766 6359 -732
rect 1636 -768 6359 -766
rect 1644 -904 1712 -870
rect 1802 -904 1870 -870
rect 1960 -904 2028 -870
rect 2118 -904 2186 -870
rect 2276 -904 2344 -870
rect 2434 -904 2502 -870
rect 2592 -904 2660 -870
rect 2750 -904 2818 -870
rect 2908 -904 2976 -870
rect 3066 -904 3134 -870
rect 3224 -904 3292 -870
rect 3382 -904 3450 -870
rect 3540 -904 3608 -870
rect 3698 -904 3766 -870
rect 3856 -904 3924 -870
rect 4014 -904 4082 -870
rect 4172 -904 4240 -870
rect 4330 -904 4398 -870
rect 4488 -904 4556 -870
rect 4646 -904 4714 -870
rect 4804 -904 4872 -870
rect 4962 -904 5030 -870
rect 5120 -904 5188 -870
rect 5278 -904 5346 -870
rect 5436 -904 5504 -870
rect 5594 -904 5662 -870
rect 5752 -904 5820 -870
rect 5910 -904 5978 -870
rect 6068 -904 6136 -870
rect 6226 -904 6294 -870
rect 7936 -766 12659 -732
rect 7936 -768 12659 -766
rect 7944 -904 8012 -870
rect 8102 -904 8170 -870
rect 8260 -904 8328 -870
rect 8418 -904 8486 -870
rect 8576 -904 8644 -870
rect 8734 -904 8802 -870
rect 8892 -904 8960 -870
rect 9050 -904 9118 -870
rect 9208 -904 9276 -870
rect 9366 -904 9434 -870
rect 9524 -904 9592 -870
rect 9682 -904 9750 -870
rect 9840 -904 9908 -870
rect 9998 -904 10066 -870
rect 10156 -904 10224 -870
rect 10314 -904 10382 -870
rect 10472 -904 10540 -870
rect 10630 -904 10698 -870
rect 10788 -904 10856 -870
rect 10946 -904 11014 -870
rect 11104 -904 11172 -870
rect 11262 -904 11330 -870
rect 11420 -904 11488 -870
rect 11578 -904 11646 -870
rect 11736 -904 11804 -870
rect 11894 -904 11962 -870
rect 12052 -904 12120 -870
rect 12210 -904 12278 -870
rect 12368 -904 12436 -870
rect 12526 -904 12594 -870
rect 14236 -766 18959 -732
rect 14236 -768 18959 -766
rect 14244 -904 14312 -870
rect 14402 -904 14470 -870
rect 14560 -904 14628 -870
rect 14718 -904 14786 -870
rect 14876 -904 14944 -870
rect 15034 -904 15102 -870
rect 15192 -904 15260 -870
rect 15350 -904 15418 -870
rect 15508 -904 15576 -870
rect 15666 -904 15734 -870
rect 15824 -904 15892 -870
rect 15982 -904 16050 -870
rect 16140 -904 16208 -870
rect 16298 -904 16366 -870
rect 16456 -904 16524 -870
rect 16614 -904 16682 -870
rect 16772 -904 16840 -870
rect 16930 -904 16998 -870
rect 17088 -904 17156 -870
rect 17246 -904 17314 -870
rect 17404 -904 17472 -870
rect 17562 -904 17630 -870
rect 17720 -904 17788 -870
rect 17878 -904 17946 -870
rect 18036 -904 18104 -870
rect 18194 -904 18262 -870
rect 18352 -904 18420 -870
rect 18510 -904 18578 -870
rect 18668 -904 18736 -870
rect 18826 -904 18894 -870
rect 20536 -766 25259 -732
rect 20536 -768 25259 -766
rect 20544 -904 20612 -870
rect 20702 -904 20770 -870
rect 20860 -904 20928 -870
rect 21018 -904 21086 -870
rect 21176 -904 21244 -870
rect 21334 -904 21402 -870
rect 21492 -904 21560 -870
rect 21650 -904 21718 -870
rect 21808 -904 21876 -870
rect 21966 -904 22034 -870
rect 22124 -904 22192 -870
rect 22282 -904 22350 -870
rect 22440 -904 22508 -870
rect 22598 -904 22666 -870
rect 22756 -904 22824 -870
rect 22914 -904 22982 -870
rect 23072 -904 23140 -870
rect 23230 -904 23298 -870
rect 23388 -904 23456 -870
rect 23546 -904 23614 -870
rect 23704 -904 23772 -870
rect 23862 -904 23930 -870
rect 24020 -904 24088 -870
rect 24178 -904 24246 -870
rect 24336 -904 24404 -870
rect 24494 -904 24562 -870
rect 24652 -904 24720 -870
rect 24810 -904 24878 -870
rect 24968 -904 25036 -870
rect 25126 -904 25194 -870
rect 1446 -6964 1448 -920
rect 1448 -6964 1482 -920
rect 1482 -6964 1484 -920
rect 1582 -6930 1616 -954
rect 1740 -6930 1774 -954
rect 1898 -6930 1932 -954
rect 2056 -6930 2090 -954
rect 2214 -6930 2248 -954
rect 2372 -6930 2406 -954
rect 2530 -6930 2564 -954
rect 2688 -6930 2722 -954
rect 2846 -6930 2880 -954
rect 3004 -6930 3038 -954
rect 3162 -6930 3196 -954
rect 3320 -6930 3354 -954
rect 3478 -6930 3512 -954
rect 3636 -6930 3670 -954
rect 3794 -6930 3828 -954
rect 3952 -6930 3986 -954
rect 4110 -6930 4144 -954
rect 4268 -6930 4302 -954
rect 4426 -6930 4460 -954
rect 4584 -6930 4618 -954
rect 4742 -6930 4776 -954
rect 4900 -6930 4934 -954
rect 5058 -6930 5092 -954
rect 5216 -6930 5250 -954
rect 5374 -6930 5408 -954
rect 5532 -6930 5566 -954
rect 5690 -6930 5724 -954
rect 5848 -6930 5882 -954
rect 6006 -6930 6040 -954
rect 6164 -6930 6198 -954
rect 6322 -6930 6356 -954
rect 6454 -6964 6456 -920
rect 6456 -6964 6490 -920
rect 6490 -6964 6492 -920
rect 7746 -6964 7748 -920
rect 7748 -6964 7782 -920
rect 7782 -6964 7784 -920
rect 7882 -6930 7916 -954
rect 8040 -6930 8074 -954
rect 8198 -6930 8232 -954
rect 8356 -6930 8390 -954
rect 8514 -6930 8548 -954
rect 8672 -6930 8706 -954
rect 8830 -6930 8864 -954
rect 8988 -6930 9022 -954
rect 9146 -6930 9180 -954
rect 9304 -6930 9338 -954
rect 9462 -6930 9496 -954
rect 9620 -6930 9654 -954
rect 9778 -6930 9812 -954
rect 9936 -6930 9970 -954
rect 10094 -6930 10128 -954
rect 10252 -6930 10286 -954
rect 10410 -6930 10444 -954
rect 10568 -6930 10602 -954
rect 10726 -6930 10760 -954
rect 10884 -6930 10918 -954
rect 11042 -6930 11076 -954
rect 11200 -6930 11234 -954
rect 11358 -6930 11392 -954
rect 11516 -6930 11550 -954
rect 11674 -6930 11708 -954
rect 11832 -6930 11866 -954
rect 11990 -6930 12024 -954
rect 12148 -6930 12182 -954
rect 12306 -6930 12340 -954
rect 12464 -6930 12498 -954
rect 12622 -6930 12656 -954
rect 12754 -6964 12756 -920
rect 12756 -6964 12790 -920
rect 12790 -6964 12792 -920
rect 14046 -6964 14048 -920
rect 14048 -6964 14082 -920
rect 14082 -6964 14084 -920
rect 14182 -6930 14216 -954
rect 14340 -6930 14374 -954
rect 14498 -6930 14532 -954
rect 14656 -6930 14690 -954
rect 14814 -6930 14848 -954
rect 14972 -6930 15006 -954
rect 15130 -6930 15164 -954
rect 15288 -6930 15322 -954
rect 15446 -6930 15480 -954
rect 15604 -6930 15638 -954
rect 15762 -6930 15796 -954
rect 15920 -6930 15954 -954
rect 16078 -6930 16112 -954
rect 16236 -6930 16270 -954
rect 16394 -6930 16428 -954
rect 16552 -6930 16586 -954
rect 16710 -6930 16744 -954
rect 16868 -6930 16902 -954
rect 17026 -6930 17060 -954
rect 17184 -6930 17218 -954
rect 17342 -6930 17376 -954
rect 17500 -6930 17534 -954
rect 17658 -6930 17692 -954
rect 17816 -6930 17850 -954
rect 17974 -6930 18008 -954
rect 18132 -6930 18166 -954
rect 18290 -6930 18324 -954
rect 18448 -6930 18482 -954
rect 18606 -6930 18640 -954
rect 18764 -6930 18798 -954
rect 18922 -6930 18956 -954
rect 19054 -6964 19056 -920
rect 19056 -6964 19090 -920
rect 19090 -6964 19092 -920
rect 20346 -6964 20348 -920
rect 20348 -6964 20382 -920
rect 20382 -6964 20384 -920
rect 20482 -6930 20516 -954
rect 20640 -6930 20674 -954
rect 20798 -6930 20832 -954
rect 20956 -6930 20990 -954
rect 21114 -6930 21148 -954
rect 21272 -6930 21306 -954
rect 21430 -6930 21464 -954
rect 21588 -6930 21622 -954
rect 21746 -6930 21780 -954
rect 21904 -6930 21938 -954
rect 22062 -6930 22096 -954
rect 22220 -6930 22254 -954
rect 22378 -6930 22412 -954
rect 22536 -6930 22570 -954
rect 22694 -6930 22728 -954
rect 22852 -6930 22886 -954
rect 23010 -6930 23044 -954
rect 23168 -6930 23202 -954
rect 23326 -6930 23360 -954
rect 23484 -6930 23518 -954
rect 23642 -6930 23676 -954
rect 23800 -6930 23834 -954
rect 23958 -6930 23992 -954
rect 24116 -6930 24150 -954
rect 24274 -6930 24308 -954
rect 24432 -6930 24466 -954
rect 24590 -6930 24624 -954
rect 24748 -6930 24782 -954
rect 24906 -6930 24940 -954
rect 25064 -6930 25098 -954
rect 25222 -6930 25256 -954
rect 25354 -6964 25356 -920
rect 25356 -6964 25390 -920
rect 25390 -6964 25392 -920
rect 1644 -7014 1712 -6980
rect 1802 -7014 1870 -6980
rect 1960 -7014 2028 -6980
rect 2118 -7014 2186 -6980
rect 2276 -7014 2344 -6980
rect 2434 -7014 2502 -6980
rect 2592 -7014 2660 -6980
rect 2750 -7014 2818 -6980
rect 2908 -7014 2976 -6980
rect 3066 -7014 3134 -6980
rect 3224 -7014 3292 -6980
rect 3382 -7014 3450 -6980
rect 3540 -7014 3608 -6980
rect 3698 -7014 3766 -6980
rect 3856 -7014 3924 -6980
rect 4014 -7014 4082 -6980
rect 4172 -7014 4240 -6980
rect 4330 -7014 4398 -6980
rect 4488 -7014 4556 -6980
rect 4646 -7014 4714 -6980
rect 4804 -7014 4872 -6980
rect 4962 -7014 5030 -6980
rect 5120 -7014 5188 -6980
rect 5278 -7014 5346 -6980
rect 5436 -7014 5504 -6980
rect 5594 -7014 5662 -6980
rect 5752 -7014 5820 -6980
rect 5910 -7014 5978 -6980
rect 6068 -7014 6136 -6980
rect 6226 -7014 6294 -6980
rect 1636 -7118 6302 -7116
rect 1636 -7152 6302 -7118
rect 7944 -7014 8012 -6980
rect 8102 -7014 8170 -6980
rect 8260 -7014 8328 -6980
rect 8418 -7014 8486 -6980
rect 8576 -7014 8644 -6980
rect 8734 -7014 8802 -6980
rect 8892 -7014 8960 -6980
rect 9050 -7014 9118 -6980
rect 9208 -7014 9276 -6980
rect 9366 -7014 9434 -6980
rect 9524 -7014 9592 -6980
rect 9682 -7014 9750 -6980
rect 9840 -7014 9908 -6980
rect 9998 -7014 10066 -6980
rect 10156 -7014 10224 -6980
rect 10314 -7014 10382 -6980
rect 10472 -7014 10540 -6980
rect 10630 -7014 10698 -6980
rect 10788 -7014 10856 -6980
rect 10946 -7014 11014 -6980
rect 11104 -7014 11172 -6980
rect 11262 -7014 11330 -6980
rect 11420 -7014 11488 -6980
rect 11578 -7014 11646 -6980
rect 11736 -7014 11804 -6980
rect 11894 -7014 11962 -6980
rect 12052 -7014 12120 -6980
rect 12210 -7014 12278 -6980
rect 12368 -7014 12436 -6980
rect 12526 -7014 12594 -6980
rect 7936 -7118 12602 -7116
rect 7936 -7152 12602 -7118
rect 14244 -7014 14312 -6980
rect 14402 -7014 14470 -6980
rect 14560 -7014 14628 -6980
rect 14718 -7014 14786 -6980
rect 14876 -7014 14944 -6980
rect 15034 -7014 15102 -6980
rect 15192 -7014 15260 -6980
rect 15350 -7014 15418 -6980
rect 15508 -7014 15576 -6980
rect 15666 -7014 15734 -6980
rect 15824 -7014 15892 -6980
rect 15982 -7014 16050 -6980
rect 16140 -7014 16208 -6980
rect 16298 -7014 16366 -6980
rect 16456 -7014 16524 -6980
rect 16614 -7014 16682 -6980
rect 16772 -7014 16840 -6980
rect 16930 -7014 16998 -6980
rect 17088 -7014 17156 -6980
rect 17246 -7014 17314 -6980
rect 17404 -7014 17472 -6980
rect 17562 -7014 17630 -6980
rect 17720 -7014 17788 -6980
rect 17878 -7014 17946 -6980
rect 18036 -7014 18104 -6980
rect 18194 -7014 18262 -6980
rect 18352 -7014 18420 -6980
rect 18510 -7014 18578 -6980
rect 18668 -7014 18736 -6980
rect 18826 -7014 18894 -6980
rect 14236 -7118 18902 -7116
rect 14236 -7152 18902 -7118
rect 20544 -7014 20612 -6980
rect 20702 -7014 20770 -6980
rect 20860 -7014 20928 -6980
rect 21018 -7014 21086 -6980
rect 21176 -7014 21244 -6980
rect 21334 -7014 21402 -6980
rect 21492 -7014 21560 -6980
rect 21650 -7014 21718 -6980
rect 21808 -7014 21876 -6980
rect 21966 -7014 22034 -6980
rect 22124 -7014 22192 -6980
rect 22282 -7014 22350 -6980
rect 22440 -7014 22508 -6980
rect 22598 -7014 22666 -6980
rect 22756 -7014 22824 -6980
rect 22914 -7014 22982 -6980
rect 23072 -7014 23140 -6980
rect 23230 -7014 23298 -6980
rect 23388 -7014 23456 -6980
rect 23546 -7014 23614 -6980
rect 23704 -7014 23772 -6980
rect 23862 -7014 23930 -6980
rect 24020 -7014 24088 -6980
rect 24178 -7014 24246 -6980
rect 24336 -7014 24404 -6980
rect 24494 -7014 24562 -6980
rect 24652 -7014 24720 -6980
rect 24810 -7014 24878 -6980
rect 24968 -7014 25036 -6980
rect 25126 -7014 25194 -6980
rect 20536 -7118 25202 -7116
rect 20536 -7152 25202 -7118
rect 1636 -7154 6302 -7152
rect 7936 -7154 12602 -7152
rect 14236 -7154 18902 -7152
rect 20536 -7154 25202 -7152
<< metal1 >>
rect 1430 6870 6510 6880
rect 1430 6832 1636 6870
rect 6359 6832 6510 6870
rect 1430 6822 6510 6832
rect 1430 6820 1500 6822
rect 6440 6820 6510 6822
rect 1632 6730 1652 6790
rect 6286 6730 6306 6790
rect 1632 6696 1644 6730
rect 6294 6696 6306 6730
rect 1632 6690 1652 6696
rect 6286 6690 6306 6696
rect 1565 6646 1635 6658
rect 1565 6638 1582 6646
rect 1616 6638 1635 6646
rect 1565 670 1582 678
rect 1616 670 1635 678
rect 1565 658 1635 670
rect 1723 6646 1793 6658
rect 1723 6638 1740 6646
rect 1774 6638 1793 6646
rect 1723 670 1740 678
rect 1774 670 1793 678
rect 1723 658 1793 670
rect 1881 6646 1951 6658
rect 1881 6638 1898 6646
rect 1932 6638 1951 6646
rect 1881 670 1898 678
rect 1932 670 1951 678
rect 1881 658 1951 670
rect 2039 6646 2109 6658
rect 2039 6638 2056 6646
rect 2090 6638 2109 6646
rect 2039 670 2056 678
rect 2090 670 2109 678
rect 2039 658 2109 670
rect 2197 6646 2267 6658
rect 2197 6638 2214 6646
rect 2248 6638 2267 6646
rect 2197 670 2214 678
rect 2248 670 2267 678
rect 2197 658 2267 670
rect 2355 6646 2425 6658
rect 2355 6638 2372 6646
rect 2406 6638 2425 6646
rect 2355 670 2372 678
rect 2406 670 2425 678
rect 2355 658 2425 670
rect 2513 6646 2583 6658
rect 2513 6638 2530 6646
rect 2564 6638 2583 6646
rect 2513 670 2530 678
rect 2564 670 2583 678
rect 2513 658 2583 670
rect 2671 6646 2741 6658
rect 2671 6638 2688 6646
rect 2722 6638 2741 6646
rect 2671 670 2688 678
rect 2722 670 2741 678
rect 2671 658 2741 670
rect 2829 6646 2899 6658
rect 2829 6638 2846 6646
rect 2880 6638 2899 6646
rect 2829 670 2846 678
rect 2880 670 2899 678
rect 2829 658 2899 670
rect 2987 6646 3057 6658
rect 2987 6638 3004 6646
rect 3038 6638 3057 6646
rect 2987 670 3004 678
rect 3038 670 3057 678
rect 2987 658 3057 670
rect 3145 6646 3215 6658
rect 3145 6638 3162 6646
rect 3196 6638 3215 6646
rect 3145 670 3162 678
rect 3196 670 3215 678
rect 3145 658 3215 670
rect 3303 6646 3373 6658
rect 3303 6638 3320 6646
rect 3354 6638 3373 6646
rect 3303 670 3320 678
rect 3354 670 3373 678
rect 3303 658 3373 670
rect 3461 6646 3531 6658
rect 3461 6638 3478 6646
rect 3512 6638 3531 6646
rect 3461 670 3478 678
rect 3512 670 3531 678
rect 3461 658 3531 670
rect 3619 6646 3689 6658
rect 3619 6638 3636 6646
rect 3670 6638 3689 6646
rect 3619 670 3636 678
rect 3670 670 3689 678
rect 3619 658 3689 670
rect 3777 6646 3847 6658
rect 3777 6638 3794 6646
rect 3828 6638 3847 6646
rect 3777 670 3794 678
rect 3828 670 3847 678
rect 3777 658 3847 670
rect 3935 6646 4005 6658
rect 3935 6638 3952 6646
rect 3986 6638 4005 6646
rect 3935 670 3952 678
rect 3986 670 4005 678
rect 3935 658 4005 670
rect 4093 6646 4163 6658
rect 4093 6638 4110 6646
rect 4144 6638 4163 6646
rect 4093 670 4110 678
rect 4144 670 4163 678
rect 4093 658 4163 670
rect 4251 6646 4321 6658
rect 4251 6638 4268 6646
rect 4302 6638 4321 6646
rect 4251 670 4268 678
rect 4302 670 4321 678
rect 4251 658 4321 670
rect 4409 6646 4479 6658
rect 4409 6638 4426 6646
rect 4460 6638 4479 6646
rect 4409 670 4426 678
rect 4460 670 4479 678
rect 4409 658 4479 670
rect 4567 6646 4637 6658
rect 4567 6638 4584 6646
rect 4618 6638 4637 6646
rect 4567 670 4584 678
rect 4618 670 4637 678
rect 4567 658 4637 670
rect 4725 6646 4795 6658
rect 4725 6638 4742 6646
rect 4776 6638 4795 6646
rect 4725 670 4742 678
rect 4776 670 4795 678
rect 4725 658 4795 670
rect 4883 6646 4953 6658
rect 4883 6638 4900 6646
rect 4934 6638 4953 6646
rect 4883 670 4900 678
rect 4934 670 4953 678
rect 4883 658 4953 670
rect 5041 6646 5111 6658
rect 5041 6638 5058 6646
rect 5092 6638 5111 6646
rect 5041 670 5058 678
rect 5092 670 5111 678
rect 5041 658 5111 670
rect 5199 6646 5269 6658
rect 5199 6638 5216 6646
rect 5250 6638 5269 6646
rect 5199 670 5216 678
rect 5250 670 5269 678
rect 5199 658 5269 670
rect 5357 6646 5427 6658
rect 5357 6638 5374 6646
rect 5408 6638 5427 6646
rect 5357 670 5374 678
rect 5408 670 5427 678
rect 5357 658 5427 670
rect 5515 6646 5585 6658
rect 5515 6638 5532 6646
rect 5566 6638 5585 6646
rect 5515 670 5532 678
rect 5566 670 5585 678
rect 5515 658 5585 670
rect 5673 6646 5743 6658
rect 5673 6638 5690 6646
rect 5724 6638 5743 6646
rect 5673 670 5690 678
rect 5724 670 5743 678
rect 5673 658 5743 670
rect 5831 6646 5901 6658
rect 5831 6638 5848 6646
rect 5882 6638 5901 6646
rect 5831 670 5848 678
rect 5882 670 5901 678
rect 5831 658 5901 670
rect 5989 6646 6059 6658
rect 5989 6638 6006 6646
rect 6040 6638 6059 6646
rect 5989 670 6006 678
rect 6040 670 6059 678
rect 5989 658 6059 670
rect 6147 6646 6217 6658
rect 6147 6638 6164 6646
rect 6198 6638 6217 6646
rect 6147 670 6164 678
rect 6198 670 6217 678
rect 6147 658 6217 670
rect 6305 6646 6375 6658
rect 6305 6638 6322 6646
rect 6356 6638 6375 6646
rect 6305 670 6322 678
rect 6356 670 6375 678
rect 6305 658 6375 670
rect 1632 620 1652 626
rect 6286 620 6306 626
rect 1632 586 1644 620
rect 6294 586 6306 620
rect 1632 526 1652 586
rect 6286 526 6306 586
rect 1430 494 1500 500
rect 6440 494 6510 500
rect 1430 484 6510 494
rect 1430 446 1636 484
rect 6302 446 6510 484
rect 1430 430 6510 446
rect 7730 6870 12810 6880
rect 7730 6832 7936 6870
rect 12659 6832 12810 6870
rect 7730 6822 12810 6832
rect 7730 6820 7800 6822
rect 12740 6820 12810 6822
rect 7932 6730 7952 6790
rect 12586 6730 12606 6790
rect 7932 6696 7944 6730
rect 12594 6696 12606 6730
rect 7932 6690 7952 6696
rect 12586 6690 12606 6696
rect 7865 6646 7935 6658
rect 7865 6638 7882 6646
rect 7916 6638 7935 6646
rect 7865 670 7882 678
rect 7916 670 7935 678
rect 7865 658 7935 670
rect 8023 6646 8093 6658
rect 8023 6638 8040 6646
rect 8074 6638 8093 6646
rect 8023 670 8040 678
rect 8074 670 8093 678
rect 8023 658 8093 670
rect 8181 6646 8251 6658
rect 8181 6638 8198 6646
rect 8232 6638 8251 6646
rect 8181 670 8198 678
rect 8232 670 8251 678
rect 8181 658 8251 670
rect 8339 6646 8409 6658
rect 8339 6638 8356 6646
rect 8390 6638 8409 6646
rect 8339 670 8356 678
rect 8390 670 8409 678
rect 8339 658 8409 670
rect 8497 6646 8567 6658
rect 8497 6638 8514 6646
rect 8548 6638 8567 6646
rect 8497 670 8514 678
rect 8548 670 8567 678
rect 8497 658 8567 670
rect 8655 6646 8725 6658
rect 8655 6638 8672 6646
rect 8706 6638 8725 6646
rect 8655 670 8672 678
rect 8706 670 8725 678
rect 8655 658 8725 670
rect 8813 6646 8883 6658
rect 8813 6638 8830 6646
rect 8864 6638 8883 6646
rect 8813 670 8830 678
rect 8864 670 8883 678
rect 8813 658 8883 670
rect 8971 6646 9041 6658
rect 8971 6638 8988 6646
rect 9022 6638 9041 6646
rect 8971 670 8988 678
rect 9022 670 9041 678
rect 8971 658 9041 670
rect 9129 6646 9199 6658
rect 9129 6638 9146 6646
rect 9180 6638 9199 6646
rect 9129 670 9146 678
rect 9180 670 9199 678
rect 9129 658 9199 670
rect 9287 6646 9357 6658
rect 9287 6638 9304 6646
rect 9338 6638 9357 6646
rect 9287 670 9304 678
rect 9338 670 9357 678
rect 9287 658 9357 670
rect 9445 6646 9515 6658
rect 9445 6638 9462 6646
rect 9496 6638 9515 6646
rect 9445 670 9462 678
rect 9496 670 9515 678
rect 9445 658 9515 670
rect 9603 6646 9673 6658
rect 9603 6638 9620 6646
rect 9654 6638 9673 6646
rect 9603 670 9620 678
rect 9654 670 9673 678
rect 9603 658 9673 670
rect 9761 6646 9831 6658
rect 9761 6638 9778 6646
rect 9812 6638 9831 6646
rect 9761 670 9778 678
rect 9812 670 9831 678
rect 9761 658 9831 670
rect 9919 6646 9989 6658
rect 9919 6638 9936 6646
rect 9970 6638 9989 6646
rect 9919 670 9936 678
rect 9970 670 9989 678
rect 9919 658 9989 670
rect 10077 6646 10147 6658
rect 10077 6638 10094 6646
rect 10128 6638 10147 6646
rect 10077 670 10094 678
rect 10128 670 10147 678
rect 10077 658 10147 670
rect 10235 6646 10305 6658
rect 10235 6638 10252 6646
rect 10286 6638 10305 6646
rect 10235 670 10252 678
rect 10286 670 10305 678
rect 10235 658 10305 670
rect 10393 6646 10463 6658
rect 10393 6638 10410 6646
rect 10444 6638 10463 6646
rect 10393 670 10410 678
rect 10444 670 10463 678
rect 10393 658 10463 670
rect 10551 6646 10621 6658
rect 10551 6638 10568 6646
rect 10602 6638 10621 6646
rect 10551 670 10568 678
rect 10602 670 10621 678
rect 10551 658 10621 670
rect 10709 6646 10779 6658
rect 10709 6638 10726 6646
rect 10760 6638 10779 6646
rect 10709 670 10726 678
rect 10760 670 10779 678
rect 10709 658 10779 670
rect 10867 6646 10937 6658
rect 10867 6638 10884 6646
rect 10918 6638 10937 6646
rect 10867 670 10884 678
rect 10918 670 10937 678
rect 10867 658 10937 670
rect 11025 6646 11095 6658
rect 11025 6638 11042 6646
rect 11076 6638 11095 6646
rect 11025 670 11042 678
rect 11076 670 11095 678
rect 11025 658 11095 670
rect 11183 6646 11253 6658
rect 11183 6638 11200 6646
rect 11234 6638 11253 6646
rect 11183 670 11200 678
rect 11234 670 11253 678
rect 11183 658 11253 670
rect 11341 6646 11411 6658
rect 11341 6638 11358 6646
rect 11392 6638 11411 6646
rect 11341 670 11358 678
rect 11392 670 11411 678
rect 11341 658 11411 670
rect 11499 6646 11569 6658
rect 11499 6638 11516 6646
rect 11550 6638 11569 6646
rect 11499 670 11516 678
rect 11550 670 11569 678
rect 11499 658 11569 670
rect 11657 6646 11727 6658
rect 11657 6638 11674 6646
rect 11708 6638 11727 6646
rect 11657 670 11674 678
rect 11708 670 11727 678
rect 11657 658 11727 670
rect 11815 6646 11885 6658
rect 11815 6638 11832 6646
rect 11866 6638 11885 6646
rect 11815 670 11832 678
rect 11866 670 11885 678
rect 11815 658 11885 670
rect 11973 6646 12043 6658
rect 11973 6638 11990 6646
rect 12024 6638 12043 6646
rect 11973 670 11990 678
rect 12024 670 12043 678
rect 11973 658 12043 670
rect 12131 6646 12201 6658
rect 12131 6638 12148 6646
rect 12182 6638 12201 6646
rect 12131 670 12148 678
rect 12182 670 12201 678
rect 12131 658 12201 670
rect 12289 6646 12359 6658
rect 12289 6638 12306 6646
rect 12340 6638 12359 6646
rect 12289 670 12306 678
rect 12340 670 12359 678
rect 12289 658 12359 670
rect 12447 6646 12517 6658
rect 12447 6638 12464 6646
rect 12498 6638 12517 6646
rect 12447 670 12464 678
rect 12498 670 12517 678
rect 12447 658 12517 670
rect 12605 6646 12675 6658
rect 12605 6638 12622 6646
rect 12656 6638 12675 6646
rect 12605 670 12622 678
rect 12656 670 12675 678
rect 12605 658 12675 670
rect 7932 620 7952 626
rect 12586 620 12606 626
rect 7932 586 7944 620
rect 12594 586 12606 620
rect 7932 526 7952 586
rect 12586 526 12606 586
rect 7730 494 7800 500
rect 12740 494 12810 500
rect 7730 484 12810 494
rect 7730 446 7936 484
rect 12602 446 12810 484
rect 7730 430 12810 446
rect 14030 6870 19110 6880
rect 14030 6832 14236 6870
rect 18959 6832 19110 6870
rect 14030 6822 19110 6832
rect 14030 6820 14100 6822
rect 19040 6820 19110 6822
rect 14232 6730 14252 6790
rect 18886 6730 18906 6790
rect 14232 6696 14244 6730
rect 18894 6696 18906 6730
rect 14232 6690 14252 6696
rect 18886 6690 18906 6696
rect 14165 6646 14235 6658
rect 14165 6638 14182 6646
rect 14216 6638 14235 6646
rect 14165 670 14182 678
rect 14216 670 14235 678
rect 14165 658 14235 670
rect 14323 6646 14393 6658
rect 14323 6638 14340 6646
rect 14374 6638 14393 6646
rect 14323 670 14340 678
rect 14374 670 14393 678
rect 14323 658 14393 670
rect 14481 6646 14551 6658
rect 14481 6638 14498 6646
rect 14532 6638 14551 6646
rect 14481 670 14498 678
rect 14532 670 14551 678
rect 14481 658 14551 670
rect 14639 6646 14709 6658
rect 14639 6638 14656 6646
rect 14690 6638 14709 6646
rect 14639 670 14656 678
rect 14690 670 14709 678
rect 14639 658 14709 670
rect 14797 6646 14867 6658
rect 14797 6638 14814 6646
rect 14848 6638 14867 6646
rect 14797 670 14814 678
rect 14848 670 14867 678
rect 14797 658 14867 670
rect 14955 6646 15025 6658
rect 14955 6638 14972 6646
rect 15006 6638 15025 6646
rect 14955 670 14972 678
rect 15006 670 15025 678
rect 14955 658 15025 670
rect 15113 6646 15183 6658
rect 15113 6638 15130 6646
rect 15164 6638 15183 6646
rect 15113 670 15130 678
rect 15164 670 15183 678
rect 15113 658 15183 670
rect 15271 6646 15341 6658
rect 15271 6638 15288 6646
rect 15322 6638 15341 6646
rect 15271 670 15288 678
rect 15322 670 15341 678
rect 15271 658 15341 670
rect 15429 6646 15499 6658
rect 15429 6638 15446 6646
rect 15480 6638 15499 6646
rect 15429 670 15446 678
rect 15480 670 15499 678
rect 15429 658 15499 670
rect 15587 6646 15657 6658
rect 15587 6638 15604 6646
rect 15638 6638 15657 6646
rect 15587 670 15604 678
rect 15638 670 15657 678
rect 15587 658 15657 670
rect 15745 6646 15815 6658
rect 15745 6638 15762 6646
rect 15796 6638 15815 6646
rect 15745 670 15762 678
rect 15796 670 15815 678
rect 15745 658 15815 670
rect 15903 6646 15973 6658
rect 15903 6638 15920 6646
rect 15954 6638 15973 6646
rect 15903 670 15920 678
rect 15954 670 15973 678
rect 15903 658 15973 670
rect 16061 6646 16131 6658
rect 16061 6638 16078 6646
rect 16112 6638 16131 6646
rect 16061 670 16078 678
rect 16112 670 16131 678
rect 16061 658 16131 670
rect 16219 6646 16289 6658
rect 16219 6638 16236 6646
rect 16270 6638 16289 6646
rect 16219 670 16236 678
rect 16270 670 16289 678
rect 16219 658 16289 670
rect 16377 6646 16447 6658
rect 16377 6638 16394 6646
rect 16428 6638 16447 6646
rect 16377 670 16394 678
rect 16428 670 16447 678
rect 16377 658 16447 670
rect 16535 6646 16605 6658
rect 16535 6638 16552 6646
rect 16586 6638 16605 6646
rect 16535 670 16552 678
rect 16586 670 16605 678
rect 16535 658 16605 670
rect 16693 6646 16763 6658
rect 16693 6638 16710 6646
rect 16744 6638 16763 6646
rect 16693 670 16710 678
rect 16744 670 16763 678
rect 16693 658 16763 670
rect 16851 6646 16921 6658
rect 16851 6638 16868 6646
rect 16902 6638 16921 6646
rect 16851 670 16868 678
rect 16902 670 16921 678
rect 16851 658 16921 670
rect 17009 6646 17079 6658
rect 17009 6638 17026 6646
rect 17060 6638 17079 6646
rect 17009 670 17026 678
rect 17060 670 17079 678
rect 17009 658 17079 670
rect 17167 6646 17237 6658
rect 17167 6638 17184 6646
rect 17218 6638 17237 6646
rect 17167 670 17184 678
rect 17218 670 17237 678
rect 17167 658 17237 670
rect 17325 6646 17395 6658
rect 17325 6638 17342 6646
rect 17376 6638 17395 6646
rect 17325 670 17342 678
rect 17376 670 17395 678
rect 17325 658 17395 670
rect 17483 6646 17553 6658
rect 17483 6638 17500 6646
rect 17534 6638 17553 6646
rect 17483 670 17500 678
rect 17534 670 17553 678
rect 17483 658 17553 670
rect 17641 6646 17711 6658
rect 17641 6638 17658 6646
rect 17692 6638 17711 6646
rect 17641 670 17658 678
rect 17692 670 17711 678
rect 17641 658 17711 670
rect 17799 6646 17869 6658
rect 17799 6638 17816 6646
rect 17850 6638 17869 6646
rect 17799 670 17816 678
rect 17850 670 17869 678
rect 17799 658 17869 670
rect 17957 6646 18027 6658
rect 17957 6638 17974 6646
rect 18008 6638 18027 6646
rect 17957 670 17974 678
rect 18008 670 18027 678
rect 17957 658 18027 670
rect 18115 6646 18185 6658
rect 18115 6638 18132 6646
rect 18166 6638 18185 6646
rect 18115 670 18132 678
rect 18166 670 18185 678
rect 18115 658 18185 670
rect 18273 6646 18343 6658
rect 18273 6638 18290 6646
rect 18324 6638 18343 6646
rect 18273 670 18290 678
rect 18324 670 18343 678
rect 18273 658 18343 670
rect 18431 6646 18501 6658
rect 18431 6638 18448 6646
rect 18482 6638 18501 6646
rect 18431 670 18448 678
rect 18482 670 18501 678
rect 18431 658 18501 670
rect 18589 6646 18659 6658
rect 18589 6638 18606 6646
rect 18640 6638 18659 6646
rect 18589 670 18606 678
rect 18640 670 18659 678
rect 18589 658 18659 670
rect 18747 6646 18817 6658
rect 18747 6638 18764 6646
rect 18798 6638 18817 6646
rect 18747 670 18764 678
rect 18798 670 18817 678
rect 18747 658 18817 670
rect 18905 6646 18975 6658
rect 18905 6638 18922 6646
rect 18956 6638 18975 6646
rect 18905 670 18922 678
rect 18956 670 18975 678
rect 18905 658 18975 670
rect 14232 620 14252 626
rect 18886 620 18906 626
rect 14232 586 14244 620
rect 18894 586 18906 620
rect 14232 526 14252 586
rect 18886 526 18906 586
rect 14030 494 14100 500
rect 19040 494 19110 500
rect 14030 484 19110 494
rect 14030 446 14236 484
rect 18902 446 19110 484
rect 14030 430 19110 446
rect 20330 6870 25410 6880
rect 20330 6832 20536 6870
rect 25259 6832 25410 6870
rect 20330 6822 25410 6832
rect 20330 6820 20400 6822
rect 25340 6820 25410 6822
rect 20532 6730 20552 6790
rect 25186 6730 25206 6790
rect 20532 6696 20544 6730
rect 25194 6696 25206 6730
rect 20532 6690 20552 6696
rect 25186 6690 25206 6696
rect 20465 6646 20535 6658
rect 20465 6638 20482 6646
rect 20516 6638 20535 6646
rect 20465 670 20482 678
rect 20516 670 20535 678
rect 20465 658 20535 670
rect 20623 6646 20693 6658
rect 20623 6638 20640 6646
rect 20674 6638 20693 6646
rect 20623 670 20640 678
rect 20674 670 20693 678
rect 20623 658 20693 670
rect 20781 6646 20851 6658
rect 20781 6638 20798 6646
rect 20832 6638 20851 6646
rect 20781 670 20798 678
rect 20832 670 20851 678
rect 20781 658 20851 670
rect 20939 6646 21009 6658
rect 20939 6638 20956 6646
rect 20990 6638 21009 6646
rect 20939 670 20956 678
rect 20990 670 21009 678
rect 20939 658 21009 670
rect 21097 6646 21167 6658
rect 21097 6638 21114 6646
rect 21148 6638 21167 6646
rect 21097 670 21114 678
rect 21148 670 21167 678
rect 21097 658 21167 670
rect 21255 6646 21325 6658
rect 21255 6638 21272 6646
rect 21306 6638 21325 6646
rect 21255 670 21272 678
rect 21306 670 21325 678
rect 21255 658 21325 670
rect 21413 6646 21483 6658
rect 21413 6638 21430 6646
rect 21464 6638 21483 6646
rect 21413 670 21430 678
rect 21464 670 21483 678
rect 21413 658 21483 670
rect 21571 6646 21641 6658
rect 21571 6638 21588 6646
rect 21622 6638 21641 6646
rect 21571 670 21588 678
rect 21622 670 21641 678
rect 21571 658 21641 670
rect 21729 6646 21799 6658
rect 21729 6638 21746 6646
rect 21780 6638 21799 6646
rect 21729 670 21746 678
rect 21780 670 21799 678
rect 21729 658 21799 670
rect 21887 6646 21957 6658
rect 21887 6638 21904 6646
rect 21938 6638 21957 6646
rect 21887 670 21904 678
rect 21938 670 21957 678
rect 21887 658 21957 670
rect 22045 6646 22115 6658
rect 22045 6638 22062 6646
rect 22096 6638 22115 6646
rect 22045 670 22062 678
rect 22096 670 22115 678
rect 22045 658 22115 670
rect 22203 6646 22273 6658
rect 22203 6638 22220 6646
rect 22254 6638 22273 6646
rect 22203 670 22220 678
rect 22254 670 22273 678
rect 22203 658 22273 670
rect 22361 6646 22431 6658
rect 22361 6638 22378 6646
rect 22412 6638 22431 6646
rect 22361 670 22378 678
rect 22412 670 22431 678
rect 22361 658 22431 670
rect 22519 6646 22589 6658
rect 22519 6638 22536 6646
rect 22570 6638 22589 6646
rect 22519 670 22536 678
rect 22570 670 22589 678
rect 22519 658 22589 670
rect 22677 6646 22747 6658
rect 22677 6638 22694 6646
rect 22728 6638 22747 6646
rect 22677 670 22694 678
rect 22728 670 22747 678
rect 22677 658 22747 670
rect 22835 6646 22905 6658
rect 22835 6638 22852 6646
rect 22886 6638 22905 6646
rect 22835 670 22852 678
rect 22886 670 22905 678
rect 22835 658 22905 670
rect 22993 6646 23063 6658
rect 22993 6638 23010 6646
rect 23044 6638 23063 6646
rect 22993 670 23010 678
rect 23044 670 23063 678
rect 22993 658 23063 670
rect 23151 6646 23221 6658
rect 23151 6638 23168 6646
rect 23202 6638 23221 6646
rect 23151 670 23168 678
rect 23202 670 23221 678
rect 23151 658 23221 670
rect 23309 6646 23379 6658
rect 23309 6638 23326 6646
rect 23360 6638 23379 6646
rect 23309 670 23326 678
rect 23360 670 23379 678
rect 23309 658 23379 670
rect 23467 6646 23537 6658
rect 23467 6638 23484 6646
rect 23518 6638 23537 6646
rect 23467 670 23484 678
rect 23518 670 23537 678
rect 23467 658 23537 670
rect 23625 6646 23695 6658
rect 23625 6638 23642 6646
rect 23676 6638 23695 6646
rect 23625 670 23642 678
rect 23676 670 23695 678
rect 23625 658 23695 670
rect 23783 6646 23853 6658
rect 23783 6638 23800 6646
rect 23834 6638 23853 6646
rect 23783 670 23800 678
rect 23834 670 23853 678
rect 23783 658 23853 670
rect 23941 6646 24011 6658
rect 23941 6638 23958 6646
rect 23992 6638 24011 6646
rect 23941 670 23958 678
rect 23992 670 24011 678
rect 23941 658 24011 670
rect 24099 6646 24169 6658
rect 24099 6638 24116 6646
rect 24150 6638 24169 6646
rect 24099 670 24116 678
rect 24150 670 24169 678
rect 24099 658 24169 670
rect 24257 6646 24327 6658
rect 24257 6638 24274 6646
rect 24308 6638 24327 6646
rect 24257 670 24274 678
rect 24308 670 24327 678
rect 24257 658 24327 670
rect 24415 6646 24485 6658
rect 24415 6638 24432 6646
rect 24466 6638 24485 6646
rect 24415 670 24432 678
rect 24466 670 24485 678
rect 24415 658 24485 670
rect 24573 6646 24643 6658
rect 24573 6638 24590 6646
rect 24624 6638 24643 6646
rect 24573 670 24590 678
rect 24624 670 24643 678
rect 24573 658 24643 670
rect 24731 6646 24801 6658
rect 24731 6638 24748 6646
rect 24782 6638 24801 6646
rect 24731 670 24748 678
rect 24782 670 24801 678
rect 24731 658 24801 670
rect 24889 6646 24959 6658
rect 24889 6638 24906 6646
rect 24940 6638 24959 6646
rect 24889 670 24906 678
rect 24940 670 24959 678
rect 24889 658 24959 670
rect 25047 6646 25117 6658
rect 25047 6638 25064 6646
rect 25098 6638 25117 6646
rect 25047 670 25064 678
rect 25098 670 25117 678
rect 25047 658 25117 670
rect 25205 6646 25275 6658
rect 25205 6638 25222 6646
rect 25256 6638 25275 6646
rect 25205 670 25222 678
rect 25256 670 25275 678
rect 25205 658 25275 670
rect 20532 620 20552 626
rect 25186 620 25206 626
rect 20532 586 20544 620
rect 25194 586 25206 620
rect 20532 526 20552 586
rect 25186 526 25206 586
rect 20330 494 20400 500
rect 25340 494 25410 500
rect 20330 484 25410 494
rect 20330 446 20536 484
rect 25202 446 25410 484
rect 20330 430 25410 446
rect 1430 -730 6510 -720
rect 1430 -768 1636 -730
rect 6359 -768 6510 -730
rect 1430 -778 6510 -768
rect 1430 -780 1500 -778
rect 6440 -780 6510 -778
rect 1632 -870 1652 -810
rect 6286 -870 6306 -810
rect 1632 -904 1644 -870
rect 6294 -904 6306 -870
rect 1632 -910 1652 -904
rect 6286 -910 6306 -904
rect 1565 -954 1635 -942
rect 1565 -962 1582 -954
rect 1616 -962 1635 -954
rect 1565 -6930 1582 -6922
rect 1616 -6930 1635 -6922
rect 1565 -6942 1635 -6930
rect 1723 -954 1793 -942
rect 1723 -962 1740 -954
rect 1774 -962 1793 -954
rect 1723 -6930 1740 -6922
rect 1774 -6930 1793 -6922
rect 1723 -6942 1793 -6930
rect 1881 -954 1951 -942
rect 1881 -962 1898 -954
rect 1932 -962 1951 -954
rect 1881 -6930 1898 -6922
rect 1932 -6930 1951 -6922
rect 1881 -6942 1951 -6930
rect 2039 -954 2109 -942
rect 2039 -962 2056 -954
rect 2090 -962 2109 -954
rect 2039 -6930 2056 -6922
rect 2090 -6930 2109 -6922
rect 2039 -6942 2109 -6930
rect 2197 -954 2267 -942
rect 2197 -962 2214 -954
rect 2248 -962 2267 -954
rect 2197 -6930 2214 -6922
rect 2248 -6930 2267 -6922
rect 2197 -6942 2267 -6930
rect 2355 -954 2425 -942
rect 2355 -962 2372 -954
rect 2406 -962 2425 -954
rect 2355 -6930 2372 -6922
rect 2406 -6930 2425 -6922
rect 2355 -6942 2425 -6930
rect 2513 -954 2583 -942
rect 2513 -962 2530 -954
rect 2564 -962 2583 -954
rect 2513 -6930 2530 -6922
rect 2564 -6930 2583 -6922
rect 2513 -6942 2583 -6930
rect 2671 -954 2741 -942
rect 2671 -962 2688 -954
rect 2722 -962 2741 -954
rect 2671 -6930 2688 -6922
rect 2722 -6930 2741 -6922
rect 2671 -6942 2741 -6930
rect 2829 -954 2899 -942
rect 2829 -962 2846 -954
rect 2880 -962 2899 -954
rect 2829 -6930 2846 -6922
rect 2880 -6930 2899 -6922
rect 2829 -6942 2899 -6930
rect 2987 -954 3057 -942
rect 2987 -962 3004 -954
rect 3038 -962 3057 -954
rect 2987 -6930 3004 -6922
rect 3038 -6930 3057 -6922
rect 2987 -6942 3057 -6930
rect 3145 -954 3215 -942
rect 3145 -962 3162 -954
rect 3196 -962 3215 -954
rect 3145 -6930 3162 -6922
rect 3196 -6930 3215 -6922
rect 3145 -6942 3215 -6930
rect 3303 -954 3373 -942
rect 3303 -962 3320 -954
rect 3354 -962 3373 -954
rect 3303 -6930 3320 -6922
rect 3354 -6930 3373 -6922
rect 3303 -6942 3373 -6930
rect 3461 -954 3531 -942
rect 3461 -962 3478 -954
rect 3512 -962 3531 -954
rect 3461 -6930 3478 -6922
rect 3512 -6930 3531 -6922
rect 3461 -6942 3531 -6930
rect 3619 -954 3689 -942
rect 3619 -962 3636 -954
rect 3670 -962 3689 -954
rect 3619 -6930 3636 -6922
rect 3670 -6930 3689 -6922
rect 3619 -6942 3689 -6930
rect 3777 -954 3847 -942
rect 3777 -962 3794 -954
rect 3828 -962 3847 -954
rect 3777 -6930 3794 -6922
rect 3828 -6930 3847 -6922
rect 3777 -6942 3847 -6930
rect 3935 -954 4005 -942
rect 3935 -962 3952 -954
rect 3986 -962 4005 -954
rect 3935 -6930 3952 -6922
rect 3986 -6930 4005 -6922
rect 3935 -6942 4005 -6930
rect 4093 -954 4163 -942
rect 4093 -962 4110 -954
rect 4144 -962 4163 -954
rect 4093 -6930 4110 -6922
rect 4144 -6930 4163 -6922
rect 4093 -6942 4163 -6930
rect 4251 -954 4321 -942
rect 4251 -962 4268 -954
rect 4302 -962 4321 -954
rect 4251 -6930 4268 -6922
rect 4302 -6930 4321 -6922
rect 4251 -6942 4321 -6930
rect 4409 -954 4479 -942
rect 4409 -962 4426 -954
rect 4460 -962 4479 -954
rect 4409 -6930 4426 -6922
rect 4460 -6930 4479 -6922
rect 4409 -6942 4479 -6930
rect 4567 -954 4637 -942
rect 4567 -962 4584 -954
rect 4618 -962 4637 -954
rect 4567 -6930 4584 -6922
rect 4618 -6930 4637 -6922
rect 4567 -6942 4637 -6930
rect 4725 -954 4795 -942
rect 4725 -962 4742 -954
rect 4776 -962 4795 -954
rect 4725 -6930 4742 -6922
rect 4776 -6930 4795 -6922
rect 4725 -6942 4795 -6930
rect 4883 -954 4953 -942
rect 4883 -962 4900 -954
rect 4934 -962 4953 -954
rect 4883 -6930 4900 -6922
rect 4934 -6930 4953 -6922
rect 4883 -6942 4953 -6930
rect 5041 -954 5111 -942
rect 5041 -962 5058 -954
rect 5092 -962 5111 -954
rect 5041 -6930 5058 -6922
rect 5092 -6930 5111 -6922
rect 5041 -6942 5111 -6930
rect 5199 -954 5269 -942
rect 5199 -962 5216 -954
rect 5250 -962 5269 -954
rect 5199 -6930 5216 -6922
rect 5250 -6930 5269 -6922
rect 5199 -6942 5269 -6930
rect 5357 -954 5427 -942
rect 5357 -962 5374 -954
rect 5408 -962 5427 -954
rect 5357 -6930 5374 -6922
rect 5408 -6930 5427 -6922
rect 5357 -6942 5427 -6930
rect 5515 -954 5585 -942
rect 5515 -962 5532 -954
rect 5566 -962 5585 -954
rect 5515 -6930 5532 -6922
rect 5566 -6930 5585 -6922
rect 5515 -6942 5585 -6930
rect 5673 -954 5743 -942
rect 5673 -962 5690 -954
rect 5724 -962 5743 -954
rect 5673 -6930 5690 -6922
rect 5724 -6930 5743 -6922
rect 5673 -6942 5743 -6930
rect 5831 -954 5901 -942
rect 5831 -962 5848 -954
rect 5882 -962 5901 -954
rect 5831 -6930 5848 -6922
rect 5882 -6930 5901 -6922
rect 5831 -6942 5901 -6930
rect 5989 -954 6059 -942
rect 5989 -962 6006 -954
rect 6040 -962 6059 -954
rect 5989 -6930 6006 -6922
rect 6040 -6930 6059 -6922
rect 5989 -6942 6059 -6930
rect 6147 -954 6217 -942
rect 6147 -962 6164 -954
rect 6198 -962 6217 -954
rect 6147 -6930 6164 -6922
rect 6198 -6930 6217 -6922
rect 6147 -6942 6217 -6930
rect 6305 -954 6375 -942
rect 6305 -962 6322 -954
rect 6356 -962 6375 -954
rect 6305 -6930 6322 -6922
rect 6356 -6930 6375 -6922
rect 6305 -6942 6375 -6930
rect 1632 -6980 1652 -6974
rect 6286 -6980 6306 -6974
rect 1632 -7014 1644 -6980
rect 6294 -7014 6306 -6980
rect 1632 -7074 1652 -7014
rect 6286 -7074 6306 -7014
rect 1430 -7106 1500 -7100
rect 6440 -7106 6510 -7100
rect 1430 -7116 6510 -7106
rect 1430 -7154 1636 -7116
rect 6302 -7154 6510 -7116
rect 1430 -7170 6510 -7154
rect 7730 -730 12810 -720
rect 7730 -768 7936 -730
rect 12659 -768 12810 -730
rect 7730 -778 12810 -768
rect 7730 -780 7800 -778
rect 12740 -780 12810 -778
rect 7932 -870 7952 -810
rect 12586 -870 12606 -810
rect 7932 -904 7944 -870
rect 12594 -904 12606 -870
rect 7932 -910 7952 -904
rect 12586 -910 12606 -904
rect 7865 -954 7935 -942
rect 7865 -962 7882 -954
rect 7916 -962 7935 -954
rect 7865 -6930 7882 -6922
rect 7916 -6930 7935 -6922
rect 7865 -6942 7935 -6930
rect 8023 -954 8093 -942
rect 8023 -962 8040 -954
rect 8074 -962 8093 -954
rect 8023 -6930 8040 -6922
rect 8074 -6930 8093 -6922
rect 8023 -6942 8093 -6930
rect 8181 -954 8251 -942
rect 8181 -962 8198 -954
rect 8232 -962 8251 -954
rect 8181 -6930 8198 -6922
rect 8232 -6930 8251 -6922
rect 8181 -6942 8251 -6930
rect 8339 -954 8409 -942
rect 8339 -962 8356 -954
rect 8390 -962 8409 -954
rect 8339 -6930 8356 -6922
rect 8390 -6930 8409 -6922
rect 8339 -6942 8409 -6930
rect 8497 -954 8567 -942
rect 8497 -962 8514 -954
rect 8548 -962 8567 -954
rect 8497 -6930 8514 -6922
rect 8548 -6930 8567 -6922
rect 8497 -6942 8567 -6930
rect 8655 -954 8725 -942
rect 8655 -962 8672 -954
rect 8706 -962 8725 -954
rect 8655 -6930 8672 -6922
rect 8706 -6930 8725 -6922
rect 8655 -6942 8725 -6930
rect 8813 -954 8883 -942
rect 8813 -962 8830 -954
rect 8864 -962 8883 -954
rect 8813 -6930 8830 -6922
rect 8864 -6930 8883 -6922
rect 8813 -6942 8883 -6930
rect 8971 -954 9041 -942
rect 8971 -962 8988 -954
rect 9022 -962 9041 -954
rect 8971 -6930 8988 -6922
rect 9022 -6930 9041 -6922
rect 8971 -6942 9041 -6930
rect 9129 -954 9199 -942
rect 9129 -962 9146 -954
rect 9180 -962 9199 -954
rect 9129 -6930 9146 -6922
rect 9180 -6930 9199 -6922
rect 9129 -6942 9199 -6930
rect 9287 -954 9357 -942
rect 9287 -962 9304 -954
rect 9338 -962 9357 -954
rect 9287 -6930 9304 -6922
rect 9338 -6930 9357 -6922
rect 9287 -6942 9357 -6930
rect 9445 -954 9515 -942
rect 9445 -962 9462 -954
rect 9496 -962 9515 -954
rect 9445 -6930 9462 -6922
rect 9496 -6930 9515 -6922
rect 9445 -6942 9515 -6930
rect 9603 -954 9673 -942
rect 9603 -962 9620 -954
rect 9654 -962 9673 -954
rect 9603 -6930 9620 -6922
rect 9654 -6930 9673 -6922
rect 9603 -6942 9673 -6930
rect 9761 -954 9831 -942
rect 9761 -962 9778 -954
rect 9812 -962 9831 -954
rect 9761 -6930 9778 -6922
rect 9812 -6930 9831 -6922
rect 9761 -6942 9831 -6930
rect 9919 -954 9989 -942
rect 9919 -962 9936 -954
rect 9970 -962 9989 -954
rect 9919 -6930 9936 -6922
rect 9970 -6930 9989 -6922
rect 9919 -6942 9989 -6930
rect 10077 -954 10147 -942
rect 10077 -962 10094 -954
rect 10128 -962 10147 -954
rect 10077 -6930 10094 -6922
rect 10128 -6930 10147 -6922
rect 10077 -6942 10147 -6930
rect 10235 -954 10305 -942
rect 10235 -962 10252 -954
rect 10286 -962 10305 -954
rect 10235 -6930 10252 -6922
rect 10286 -6930 10305 -6922
rect 10235 -6942 10305 -6930
rect 10393 -954 10463 -942
rect 10393 -962 10410 -954
rect 10444 -962 10463 -954
rect 10393 -6930 10410 -6922
rect 10444 -6930 10463 -6922
rect 10393 -6942 10463 -6930
rect 10551 -954 10621 -942
rect 10551 -962 10568 -954
rect 10602 -962 10621 -954
rect 10551 -6930 10568 -6922
rect 10602 -6930 10621 -6922
rect 10551 -6942 10621 -6930
rect 10709 -954 10779 -942
rect 10709 -962 10726 -954
rect 10760 -962 10779 -954
rect 10709 -6930 10726 -6922
rect 10760 -6930 10779 -6922
rect 10709 -6942 10779 -6930
rect 10867 -954 10937 -942
rect 10867 -962 10884 -954
rect 10918 -962 10937 -954
rect 10867 -6930 10884 -6922
rect 10918 -6930 10937 -6922
rect 10867 -6942 10937 -6930
rect 11025 -954 11095 -942
rect 11025 -962 11042 -954
rect 11076 -962 11095 -954
rect 11025 -6930 11042 -6922
rect 11076 -6930 11095 -6922
rect 11025 -6942 11095 -6930
rect 11183 -954 11253 -942
rect 11183 -962 11200 -954
rect 11234 -962 11253 -954
rect 11183 -6930 11200 -6922
rect 11234 -6930 11253 -6922
rect 11183 -6942 11253 -6930
rect 11341 -954 11411 -942
rect 11341 -962 11358 -954
rect 11392 -962 11411 -954
rect 11341 -6930 11358 -6922
rect 11392 -6930 11411 -6922
rect 11341 -6942 11411 -6930
rect 11499 -954 11569 -942
rect 11499 -962 11516 -954
rect 11550 -962 11569 -954
rect 11499 -6930 11516 -6922
rect 11550 -6930 11569 -6922
rect 11499 -6942 11569 -6930
rect 11657 -954 11727 -942
rect 11657 -962 11674 -954
rect 11708 -962 11727 -954
rect 11657 -6930 11674 -6922
rect 11708 -6930 11727 -6922
rect 11657 -6942 11727 -6930
rect 11815 -954 11885 -942
rect 11815 -962 11832 -954
rect 11866 -962 11885 -954
rect 11815 -6930 11832 -6922
rect 11866 -6930 11885 -6922
rect 11815 -6942 11885 -6930
rect 11973 -954 12043 -942
rect 11973 -962 11990 -954
rect 12024 -962 12043 -954
rect 11973 -6930 11990 -6922
rect 12024 -6930 12043 -6922
rect 11973 -6942 12043 -6930
rect 12131 -954 12201 -942
rect 12131 -962 12148 -954
rect 12182 -962 12201 -954
rect 12131 -6930 12148 -6922
rect 12182 -6930 12201 -6922
rect 12131 -6942 12201 -6930
rect 12289 -954 12359 -942
rect 12289 -962 12306 -954
rect 12340 -962 12359 -954
rect 12289 -6930 12306 -6922
rect 12340 -6930 12359 -6922
rect 12289 -6942 12359 -6930
rect 12447 -954 12517 -942
rect 12447 -962 12464 -954
rect 12498 -962 12517 -954
rect 12447 -6930 12464 -6922
rect 12498 -6930 12517 -6922
rect 12447 -6942 12517 -6930
rect 12605 -954 12675 -942
rect 12605 -962 12622 -954
rect 12656 -962 12675 -954
rect 12605 -6930 12622 -6922
rect 12656 -6930 12675 -6922
rect 12605 -6942 12675 -6930
rect 7932 -6980 7952 -6974
rect 12586 -6980 12606 -6974
rect 7932 -7014 7944 -6980
rect 12594 -7014 12606 -6980
rect 7932 -7074 7952 -7014
rect 12586 -7074 12606 -7014
rect 7730 -7106 7800 -7100
rect 12740 -7106 12810 -7100
rect 7730 -7116 12810 -7106
rect 7730 -7154 7936 -7116
rect 12602 -7154 12810 -7116
rect 7730 -7170 12810 -7154
rect 14030 -730 19110 -720
rect 14030 -768 14236 -730
rect 18959 -768 19110 -730
rect 14030 -778 19110 -768
rect 14030 -780 14100 -778
rect 19040 -780 19110 -778
rect 14232 -870 14252 -810
rect 18886 -870 18906 -810
rect 14232 -904 14244 -870
rect 18894 -904 18906 -870
rect 14232 -910 14252 -904
rect 18886 -910 18906 -904
rect 14165 -954 14235 -942
rect 14165 -962 14182 -954
rect 14216 -962 14235 -954
rect 14165 -6930 14182 -6922
rect 14216 -6930 14235 -6922
rect 14165 -6942 14235 -6930
rect 14323 -954 14393 -942
rect 14323 -962 14340 -954
rect 14374 -962 14393 -954
rect 14323 -6930 14340 -6922
rect 14374 -6930 14393 -6922
rect 14323 -6942 14393 -6930
rect 14481 -954 14551 -942
rect 14481 -962 14498 -954
rect 14532 -962 14551 -954
rect 14481 -6930 14498 -6922
rect 14532 -6930 14551 -6922
rect 14481 -6942 14551 -6930
rect 14639 -954 14709 -942
rect 14639 -962 14656 -954
rect 14690 -962 14709 -954
rect 14639 -6930 14656 -6922
rect 14690 -6930 14709 -6922
rect 14639 -6942 14709 -6930
rect 14797 -954 14867 -942
rect 14797 -962 14814 -954
rect 14848 -962 14867 -954
rect 14797 -6930 14814 -6922
rect 14848 -6930 14867 -6922
rect 14797 -6942 14867 -6930
rect 14955 -954 15025 -942
rect 14955 -962 14972 -954
rect 15006 -962 15025 -954
rect 14955 -6930 14972 -6922
rect 15006 -6930 15025 -6922
rect 14955 -6942 15025 -6930
rect 15113 -954 15183 -942
rect 15113 -962 15130 -954
rect 15164 -962 15183 -954
rect 15113 -6930 15130 -6922
rect 15164 -6930 15183 -6922
rect 15113 -6942 15183 -6930
rect 15271 -954 15341 -942
rect 15271 -962 15288 -954
rect 15322 -962 15341 -954
rect 15271 -6930 15288 -6922
rect 15322 -6930 15341 -6922
rect 15271 -6942 15341 -6930
rect 15429 -954 15499 -942
rect 15429 -962 15446 -954
rect 15480 -962 15499 -954
rect 15429 -6930 15446 -6922
rect 15480 -6930 15499 -6922
rect 15429 -6942 15499 -6930
rect 15587 -954 15657 -942
rect 15587 -962 15604 -954
rect 15638 -962 15657 -954
rect 15587 -6930 15604 -6922
rect 15638 -6930 15657 -6922
rect 15587 -6942 15657 -6930
rect 15745 -954 15815 -942
rect 15745 -962 15762 -954
rect 15796 -962 15815 -954
rect 15745 -6930 15762 -6922
rect 15796 -6930 15815 -6922
rect 15745 -6942 15815 -6930
rect 15903 -954 15973 -942
rect 15903 -962 15920 -954
rect 15954 -962 15973 -954
rect 15903 -6930 15920 -6922
rect 15954 -6930 15973 -6922
rect 15903 -6942 15973 -6930
rect 16061 -954 16131 -942
rect 16061 -962 16078 -954
rect 16112 -962 16131 -954
rect 16061 -6930 16078 -6922
rect 16112 -6930 16131 -6922
rect 16061 -6942 16131 -6930
rect 16219 -954 16289 -942
rect 16219 -962 16236 -954
rect 16270 -962 16289 -954
rect 16219 -6930 16236 -6922
rect 16270 -6930 16289 -6922
rect 16219 -6942 16289 -6930
rect 16377 -954 16447 -942
rect 16377 -962 16394 -954
rect 16428 -962 16447 -954
rect 16377 -6930 16394 -6922
rect 16428 -6930 16447 -6922
rect 16377 -6942 16447 -6930
rect 16535 -954 16605 -942
rect 16535 -962 16552 -954
rect 16586 -962 16605 -954
rect 16535 -6930 16552 -6922
rect 16586 -6930 16605 -6922
rect 16535 -6942 16605 -6930
rect 16693 -954 16763 -942
rect 16693 -962 16710 -954
rect 16744 -962 16763 -954
rect 16693 -6930 16710 -6922
rect 16744 -6930 16763 -6922
rect 16693 -6942 16763 -6930
rect 16851 -954 16921 -942
rect 16851 -962 16868 -954
rect 16902 -962 16921 -954
rect 16851 -6930 16868 -6922
rect 16902 -6930 16921 -6922
rect 16851 -6942 16921 -6930
rect 17009 -954 17079 -942
rect 17009 -962 17026 -954
rect 17060 -962 17079 -954
rect 17009 -6930 17026 -6922
rect 17060 -6930 17079 -6922
rect 17009 -6942 17079 -6930
rect 17167 -954 17237 -942
rect 17167 -962 17184 -954
rect 17218 -962 17237 -954
rect 17167 -6930 17184 -6922
rect 17218 -6930 17237 -6922
rect 17167 -6942 17237 -6930
rect 17325 -954 17395 -942
rect 17325 -962 17342 -954
rect 17376 -962 17395 -954
rect 17325 -6930 17342 -6922
rect 17376 -6930 17395 -6922
rect 17325 -6942 17395 -6930
rect 17483 -954 17553 -942
rect 17483 -962 17500 -954
rect 17534 -962 17553 -954
rect 17483 -6930 17500 -6922
rect 17534 -6930 17553 -6922
rect 17483 -6942 17553 -6930
rect 17641 -954 17711 -942
rect 17641 -962 17658 -954
rect 17692 -962 17711 -954
rect 17641 -6930 17658 -6922
rect 17692 -6930 17711 -6922
rect 17641 -6942 17711 -6930
rect 17799 -954 17869 -942
rect 17799 -962 17816 -954
rect 17850 -962 17869 -954
rect 17799 -6930 17816 -6922
rect 17850 -6930 17869 -6922
rect 17799 -6942 17869 -6930
rect 17957 -954 18027 -942
rect 17957 -962 17974 -954
rect 18008 -962 18027 -954
rect 17957 -6930 17974 -6922
rect 18008 -6930 18027 -6922
rect 17957 -6942 18027 -6930
rect 18115 -954 18185 -942
rect 18115 -962 18132 -954
rect 18166 -962 18185 -954
rect 18115 -6930 18132 -6922
rect 18166 -6930 18185 -6922
rect 18115 -6942 18185 -6930
rect 18273 -954 18343 -942
rect 18273 -962 18290 -954
rect 18324 -962 18343 -954
rect 18273 -6930 18290 -6922
rect 18324 -6930 18343 -6922
rect 18273 -6942 18343 -6930
rect 18431 -954 18501 -942
rect 18431 -962 18448 -954
rect 18482 -962 18501 -954
rect 18431 -6930 18448 -6922
rect 18482 -6930 18501 -6922
rect 18431 -6942 18501 -6930
rect 18589 -954 18659 -942
rect 18589 -962 18606 -954
rect 18640 -962 18659 -954
rect 18589 -6930 18606 -6922
rect 18640 -6930 18659 -6922
rect 18589 -6942 18659 -6930
rect 18747 -954 18817 -942
rect 18747 -962 18764 -954
rect 18798 -962 18817 -954
rect 18747 -6930 18764 -6922
rect 18798 -6930 18817 -6922
rect 18747 -6942 18817 -6930
rect 18905 -954 18975 -942
rect 18905 -962 18922 -954
rect 18956 -962 18975 -954
rect 18905 -6930 18922 -6922
rect 18956 -6930 18975 -6922
rect 18905 -6942 18975 -6930
rect 14232 -6980 14252 -6974
rect 18886 -6980 18906 -6974
rect 14232 -7014 14244 -6980
rect 18894 -7014 18906 -6980
rect 14232 -7074 14252 -7014
rect 18886 -7074 18906 -7014
rect 14030 -7106 14100 -7100
rect 19040 -7106 19110 -7100
rect 14030 -7116 19110 -7106
rect 14030 -7154 14236 -7116
rect 18902 -7154 19110 -7116
rect 14030 -7170 19110 -7154
rect 20330 -730 25410 -720
rect 20330 -768 20536 -730
rect 25259 -768 25410 -730
rect 20330 -778 25410 -768
rect 20330 -780 20400 -778
rect 25340 -780 25410 -778
rect 20532 -870 20552 -810
rect 25186 -870 25206 -810
rect 20532 -904 20544 -870
rect 25194 -904 25206 -870
rect 20532 -910 20552 -904
rect 25186 -910 25206 -904
rect 20465 -954 20535 -942
rect 20465 -962 20482 -954
rect 20516 -962 20535 -954
rect 20465 -6930 20482 -6922
rect 20516 -6930 20535 -6922
rect 20465 -6942 20535 -6930
rect 20623 -954 20693 -942
rect 20623 -962 20640 -954
rect 20674 -962 20693 -954
rect 20623 -6930 20640 -6922
rect 20674 -6930 20693 -6922
rect 20623 -6942 20693 -6930
rect 20781 -954 20851 -942
rect 20781 -962 20798 -954
rect 20832 -962 20851 -954
rect 20781 -6930 20798 -6922
rect 20832 -6930 20851 -6922
rect 20781 -6942 20851 -6930
rect 20939 -954 21009 -942
rect 20939 -962 20956 -954
rect 20990 -962 21009 -954
rect 20939 -6930 20956 -6922
rect 20990 -6930 21009 -6922
rect 20939 -6942 21009 -6930
rect 21097 -954 21167 -942
rect 21097 -962 21114 -954
rect 21148 -962 21167 -954
rect 21097 -6930 21114 -6922
rect 21148 -6930 21167 -6922
rect 21097 -6942 21167 -6930
rect 21255 -954 21325 -942
rect 21255 -962 21272 -954
rect 21306 -962 21325 -954
rect 21255 -6930 21272 -6922
rect 21306 -6930 21325 -6922
rect 21255 -6942 21325 -6930
rect 21413 -954 21483 -942
rect 21413 -962 21430 -954
rect 21464 -962 21483 -954
rect 21413 -6930 21430 -6922
rect 21464 -6930 21483 -6922
rect 21413 -6942 21483 -6930
rect 21571 -954 21641 -942
rect 21571 -962 21588 -954
rect 21622 -962 21641 -954
rect 21571 -6930 21588 -6922
rect 21622 -6930 21641 -6922
rect 21571 -6942 21641 -6930
rect 21729 -954 21799 -942
rect 21729 -962 21746 -954
rect 21780 -962 21799 -954
rect 21729 -6930 21746 -6922
rect 21780 -6930 21799 -6922
rect 21729 -6942 21799 -6930
rect 21887 -954 21957 -942
rect 21887 -962 21904 -954
rect 21938 -962 21957 -954
rect 21887 -6930 21904 -6922
rect 21938 -6930 21957 -6922
rect 21887 -6942 21957 -6930
rect 22045 -954 22115 -942
rect 22045 -962 22062 -954
rect 22096 -962 22115 -954
rect 22045 -6930 22062 -6922
rect 22096 -6930 22115 -6922
rect 22045 -6942 22115 -6930
rect 22203 -954 22273 -942
rect 22203 -962 22220 -954
rect 22254 -962 22273 -954
rect 22203 -6930 22220 -6922
rect 22254 -6930 22273 -6922
rect 22203 -6942 22273 -6930
rect 22361 -954 22431 -942
rect 22361 -962 22378 -954
rect 22412 -962 22431 -954
rect 22361 -6930 22378 -6922
rect 22412 -6930 22431 -6922
rect 22361 -6942 22431 -6930
rect 22519 -954 22589 -942
rect 22519 -962 22536 -954
rect 22570 -962 22589 -954
rect 22519 -6930 22536 -6922
rect 22570 -6930 22589 -6922
rect 22519 -6942 22589 -6930
rect 22677 -954 22747 -942
rect 22677 -962 22694 -954
rect 22728 -962 22747 -954
rect 22677 -6930 22694 -6922
rect 22728 -6930 22747 -6922
rect 22677 -6942 22747 -6930
rect 22835 -954 22905 -942
rect 22835 -962 22852 -954
rect 22886 -962 22905 -954
rect 22835 -6930 22852 -6922
rect 22886 -6930 22905 -6922
rect 22835 -6942 22905 -6930
rect 22993 -954 23063 -942
rect 22993 -962 23010 -954
rect 23044 -962 23063 -954
rect 22993 -6930 23010 -6922
rect 23044 -6930 23063 -6922
rect 22993 -6942 23063 -6930
rect 23151 -954 23221 -942
rect 23151 -962 23168 -954
rect 23202 -962 23221 -954
rect 23151 -6930 23168 -6922
rect 23202 -6930 23221 -6922
rect 23151 -6942 23221 -6930
rect 23309 -954 23379 -942
rect 23309 -962 23326 -954
rect 23360 -962 23379 -954
rect 23309 -6930 23326 -6922
rect 23360 -6930 23379 -6922
rect 23309 -6942 23379 -6930
rect 23467 -954 23537 -942
rect 23467 -962 23484 -954
rect 23518 -962 23537 -954
rect 23467 -6930 23484 -6922
rect 23518 -6930 23537 -6922
rect 23467 -6942 23537 -6930
rect 23625 -954 23695 -942
rect 23625 -962 23642 -954
rect 23676 -962 23695 -954
rect 23625 -6930 23642 -6922
rect 23676 -6930 23695 -6922
rect 23625 -6942 23695 -6930
rect 23783 -954 23853 -942
rect 23783 -962 23800 -954
rect 23834 -962 23853 -954
rect 23783 -6930 23800 -6922
rect 23834 -6930 23853 -6922
rect 23783 -6942 23853 -6930
rect 23941 -954 24011 -942
rect 23941 -962 23958 -954
rect 23992 -962 24011 -954
rect 23941 -6930 23958 -6922
rect 23992 -6930 24011 -6922
rect 23941 -6942 24011 -6930
rect 24099 -954 24169 -942
rect 24099 -962 24116 -954
rect 24150 -962 24169 -954
rect 24099 -6930 24116 -6922
rect 24150 -6930 24169 -6922
rect 24099 -6942 24169 -6930
rect 24257 -954 24327 -942
rect 24257 -962 24274 -954
rect 24308 -962 24327 -954
rect 24257 -6930 24274 -6922
rect 24308 -6930 24327 -6922
rect 24257 -6942 24327 -6930
rect 24415 -954 24485 -942
rect 24415 -962 24432 -954
rect 24466 -962 24485 -954
rect 24415 -6930 24432 -6922
rect 24466 -6930 24485 -6922
rect 24415 -6942 24485 -6930
rect 24573 -954 24643 -942
rect 24573 -962 24590 -954
rect 24624 -962 24643 -954
rect 24573 -6930 24590 -6922
rect 24624 -6930 24643 -6922
rect 24573 -6942 24643 -6930
rect 24731 -954 24801 -942
rect 24731 -962 24748 -954
rect 24782 -962 24801 -954
rect 24731 -6930 24748 -6922
rect 24782 -6930 24801 -6922
rect 24731 -6942 24801 -6930
rect 24889 -954 24959 -942
rect 24889 -962 24906 -954
rect 24940 -962 24959 -954
rect 24889 -6930 24906 -6922
rect 24940 -6930 24959 -6922
rect 24889 -6942 24959 -6930
rect 25047 -954 25117 -942
rect 25047 -962 25064 -954
rect 25098 -962 25117 -954
rect 25047 -6930 25064 -6922
rect 25098 -6930 25117 -6922
rect 25047 -6942 25117 -6930
rect 25205 -954 25275 -942
rect 25205 -962 25222 -954
rect 25256 -962 25275 -954
rect 25205 -6930 25222 -6922
rect 25256 -6930 25275 -6922
rect 25205 -6942 25275 -6930
rect 20532 -6980 20552 -6974
rect 25186 -6980 25206 -6974
rect 20532 -7014 20544 -6980
rect 25194 -7014 25206 -6980
rect 20532 -7074 20552 -7014
rect 25186 -7074 25206 -7014
rect 20330 -7106 20400 -7100
rect 25340 -7106 25410 -7100
rect 20330 -7116 25410 -7106
rect 20330 -7154 20536 -7116
rect 25202 -7154 25410 -7116
rect 20330 -7170 25410 -7154
<< via1 >>
rect 1430 6680 1500 6820
rect 1652 6730 6286 6790
rect 1652 6696 1712 6730
rect 1712 6696 1802 6730
rect 1802 6696 1870 6730
rect 1870 6696 1960 6730
rect 1960 6696 2028 6730
rect 2028 6696 2118 6730
rect 2118 6696 2186 6730
rect 2186 6696 2276 6730
rect 2276 6696 2344 6730
rect 2344 6696 2434 6730
rect 2434 6696 2502 6730
rect 2502 6696 2592 6730
rect 2592 6696 2660 6730
rect 2660 6696 2750 6730
rect 2750 6696 2818 6730
rect 2818 6696 2908 6730
rect 2908 6696 2976 6730
rect 2976 6696 3066 6730
rect 3066 6696 3134 6730
rect 3134 6696 3224 6730
rect 3224 6696 3292 6730
rect 3292 6696 3382 6730
rect 3382 6696 3450 6730
rect 3450 6696 3540 6730
rect 3540 6696 3608 6730
rect 3608 6696 3698 6730
rect 3698 6696 3766 6730
rect 3766 6696 3856 6730
rect 3856 6696 3924 6730
rect 3924 6696 4014 6730
rect 4014 6696 4082 6730
rect 4082 6696 4172 6730
rect 4172 6696 4240 6730
rect 4240 6696 4330 6730
rect 4330 6696 4398 6730
rect 4398 6696 4488 6730
rect 4488 6696 4556 6730
rect 4556 6696 4646 6730
rect 4646 6696 4714 6730
rect 4714 6696 4804 6730
rect 4804 6696 4872 6730
rect 4872 6696 4962 6730
rect 4962 6696 5030 6730
rect 5030 6696 5120 6730
rect 5120 6696 5188 6730
rect 5188 6696 5278 6730
rect 5278 6696 5346 6730
rect 5346 6696 5436 6730
rect 5436 6696 5504 6730
rect 5504 6696 5594 6730
rect 5594 6696 5662 6730
rect 5662 6696 5752 6730
rect 5752 6696 5820 6730
rect 5820 6696 5910 6730
rect 5910 6696 5978 6730
rect 5978 6696 6068 6730
rect 6068 6696 6136 6730
rect 6136 6696 6226 6730
rect 6226 6696 6286 6730
rect 1652 6690 6286 6696
rect 1430 636 1446 6680
rect 1446 636 1484 6680
rect 1484 636 1500 6680
rect 6440 6680 6510 6820
rect 1565 678 1582 6638
rect 1582 678 1616 6638
rect 1616 678 1635 6638
rect 1723 678 1740 6638
rect 1740 678 1774 6638
rect 1774 678 1793 6638
rect 1881 678 1898 6638
rect 1898 678 1932 6638
rect 1932 678 1951 6638
rect 2039 678 2056 6638
rect 2056 678 2090 6638
rect 2090 678 2109 6638
rect 2197 678 2214 6638
rect 2214 678 2248 6638
rect 2248 678 2267 6638
rect 2355 678 2372 6638
rect 2372 678 2406 6638
rect 2406 678 2425 6638
rect 2513 678 2530 6638
rect 2530 678 2564 6638
rect 2564 678 2583 6638
rect 2671 678 2688 6638
rect 2688 678 2722 6638
rect 2722 678 2741 6638
rect 2829 678 2846 6638
rect 2846 678 2880 6638
rect 2880 678 2899 6638
rect 2987 678 3004 6638
rect 3004 678 3038 6638
rect 3038 678 3057 6638
rect 3145 678 3162 6638
rect 3162 678 3196 6638
rect 3196 678 3215 6638
rect 3303 678 3320 6638
rect 3320 678 3354 6638
rect 3354 678 3373 6638
rect 3461 678 3478 6638
rect 3478 678 3512 6638
rect 3512 678 3531 6638
rect 3619 678 3636 6638
rect 3636 678 3670 6638
rect 3670 678 3689 6638
rect 3777 678 3794 6638
rect 3794 678 3828 6638
rect 3828 678 3847 6638
rect 3935 678 3952 6638
rect 3952 678 3986 6638
rect 3986 678 4005 6638
rect 4093 678 4110 6638
rect 4110 678 4144 6638
rect 4144 678 4163 6638
rect 4251 678 4268 6638
rect 4268 678 4302 6638
rect 4302 678 4321 6638
rect 4409 678 4426 6638
rect 4426 678 4460 6638
rect 4460 678 4479 6638
rect 4567 678 4584 6638
rect 4584 678 4618 6638
rect 4618 678 4637 6638
rect 4725 678 4742 6638
rect 4742 678 4776 6638
rect 4776 678 4795 6638
rect 4883 678 4900 6638
rect 4900 678 4934 6638
rect 4934 678 4953 6638
rect 5041 678 5058 6638
rect 5058 678 5092 6638
rect 5092 678 5111 6638
rect 5199 678 5216 6638
rect 5216 678 5250 6638
rect 5250 678 5269 6638
rect 5357 678 5374 6638
rect 5374 678 5408 6638
rect 5408 678 5427 6638
rect 5515 678 5532 6638
rect 5532 678 5566 6638
rect 5566 678 5585 6638
rect 5673 678 5690 6638
rect 5690 678 5724 6638
rect 5724 678 5743 6638
rect 5831 678 5848 6638
rect 5848 678 5882 6638
rect 5882 678 5901 6638
rect 5989 678 6006 6638
rect 6006 678 6040 6638
rect 6040 678 6059 6638
rect 6147 678 6164 6638
rect 6164 678 6198 6638
rect 6198 678 6217 6638
rect 6305 678 6322 6638
rect 6322 678 6356 6638
rect 6356 678 6375 6638
rect 1430 500 1500 636
rect 6440 636 6454 6680
rect 6454 636 6492 6680
rect 6492 636 6510 6680
rect 1652 620 6286 626
rect 1652 586 1712 620
rect 1712 586 1802 620
rect 1802 586 1870 620
rect 1870 586 1960 620
rect 1960 586 2028 620
rect 2028 586 2118 620
rect 2118 586 2186 620
rect 2186 586 2276 620
rect 2276 586 2344 620
rect 2344 586 2434 620
rect 2434 586 2502 620
rect 2502 586 2592 620
rect 2592 586 2660 620
rect 2660 586 2750 620
rect 2750 586 2818 620
rect 2818 586 2908 620
rect 2908 586 2976 620
rect 2976 586 3066 620
rect 3066 586 3134 620
rect 3134 586 3224 620
rect 3224 586 3292 620
rect 3292 586 3382 620
rect 3382 586 3450 620
rect 3450 586 3540 620
rect 3540 586 3608 620
rect 3608 586 3698 620
rect 3698 586 3766 620
rect 3766 586 3856 620
rect 3856 586 3924 620
rect 3924 586 4014 620
rect 4014 586 4082 620
rect 4082 586 4172 620
rect 4172 586 4240 620
rect 4240 586 4330 620
rect 4330 586 4398 620
rect 4398 586 4488 620
rect 4488 586 4556 620
rect 4556 586 4646 620
rect 4646 586 4714 620
rect 4714 586 4804 620
rect 4804 586 4872 620
rect 4872 586 4962 620
rect 4962 586 5030 620
rect 5030 586 5120 620
rect 5120 586 5188 620
rect 5188 586 5278 620
rect 5278 586 5346 620
rect 5346 586 5436 620
rect 5436 586 5504 620
rect 5504 586 5594 620
rect 5594 586 5662 620
rect 5662 586 5752 620
rect 5752 586 5820 620
rect 5820 586 5910 620
rect 5910 586 5978 620
rect 5978 586 6068 620
rect 6068 586 6136 620
rect 6136 586 6226 620
rect 6226 586 6286 620
rect 1652 526 6286 586
rect 6440 500 6510 636
rect 7730 6680 7800 6820
rect 7952 6730 12586 6790
rect 7952 6696 8012 6730
rect 8012 6696 8102 6730
rect 8102 6696 8170 6730
rect 8170 6696 8260 6730
rect 8260 6696 8328 6730
rect 8328 6696 8418 6730
rect 8418 6696 8486 6730
rect 8486 6696 8576 6730
rect 8576 6696 8644 6730
rect 8644 6696 8734 6730
rect 8734 6696 8802 6730
rect 8802 6696 8892 6730
rect 8892 6696 8960 6730
rect 8960 6696 9050 6730
rect 9050 6696 9118 6730
rect 9118 6696 9208 6730
rect 9208 6696 9276 6730
rect 9276 6696 9366 6730
rect 9366 6696 9434 6730
rect 9434 6696 9524 6730
rect 9524 6696 9592 6730
rect 9592 6696 9682 6730
rect 9682 6696 9750 6730
rect 9750 6696 9840 6730
rect 9840 6696 9908 6730
rect 9908 6696 9998 6730
rect 9998 6696 10066 6730
rect 10066 6696 10156 6730
rect 10156 6696 10224 6730
rect 10224 6696 10314 6730
rect 10314 6696 10382 6730
rect 10382 6696 10472 6730
rect 10472 6696 10540 6730
rect 10540 6696 10630 6730
rect 10630 6696 10698 6730
rect 10698 6696 10788 6730
rect 10788 6696 10856 6730
rect 10856 6696 10946 6730
rect 10946 6696 11014 6730
rect 11014 6696 11104 6730
rect 11104 6696 11172 6730
rect 11172 6696 11262 6730
rect 11262 6696 11330 6730
rect 11330 6696 11420 6730
rect 11420 6696 11488 6730
rect 11488 6696 11578 6730
rect 11578 6696 11646 6730
rect 11646 6696 11736 6730
rect 11736 6696 11804 6730
rect 11804 6696 11894 6730
rect 11894 6696 11962 6730
rect 11962 6696 12052 6730
rect 12052 6696 12120 6730
rect 12120 6696 12210 6730
rect 12210 6696 12278 6730
rect 12278 6696 12368 6730
rect 12368 6696 12436 6730
rect 12436 6696 12526 6730
rect 12526 6696 12586 6730
rect 7952 6690 12586 6696
rect 7730 636 7746 6680
rect 7746 636 7784 6680
rect 7784 636 7800 6680
rect 12740 6680 12810 6820
rect 7865 678 7882 6638
rect 7882 678 7916 6638
rect 7916 678 7935 6638
rect 8023 678 8040 6638
rect 8040 678 8074 6638
rect 8074 678 8093 6638
rect 8181 678 8198 6638
rect 8198 678 8232 6638
rect 8232 678 8251 6638
rect 8339 678 8356 6638
rect 8356 678 8390 6638
rect 8390 678 8409 6638
rect 8497 678 8514 6638
rect 8514 678 8548 6638
rect 8548 678 8567 6638
rect 8655 678 8672 6638
rect 8672 678 8706 6638
rect 8706 678 8725 6638
rect 8813 678 8830 6638
rect 8830 678 8864 6638
rect 8864 678 8883 6638
rect 8971 678 8988 6638
rect 8988 678 9022 6638
rect 9022 678 9041 6638
rect 9129 678 9146 6638
rect 9146 678 9180 6638
rect 9180 678 9199 6638
rect 9287 678 9304 6638
rect 9304 678 9338 6638
rect 9338 678 9357 6638
rect 9445 678 9462 6638
rect 9462 678 9496 6638
rect 9496 678 9515 6638
rect 9603 678 9620 6638
rect 9620 678 9654 6638
rect 9654 678 9673 6638
rect 9761 678 9778 6638
rect 9778 678 9812 6638
rect 9812 678 9831 6638
rect 9919 678 9936 6638
rect 9936 678 9970 6638
rect 9970 678 9989 6638
rect 10077 678 10094 6638
rect 10094 678 10128 6638
rect 10128 678 10147 6638
rect 10235 678 10252 6638
rect 10252 678 10286 6638
rect 10286 678 10305 6638
rect 10393 678 10410 6638
rect 10410 678 10444 6638
rect 10444 678 10463 6638
rect 10551 678 10568 6638
rect 10568 678 10602 6638
rect 10602 678 10621 6638
rect 10709 678 10726 6638
rect 10726 678 10760 6638
rect 10760 678 10779 6638
rect 10867 678 10884 6638
rect 10884 678 10918 6638
rect 10918 678 10937 6638
rect 11025 678 11042 6638
rect 11042 678 11076 6638
rect 11076 678 11095 6638
rect 11183 678 11200 6638
rect 11200 678 11234 6638
rect 11234 678 11253 6638
rect 11341 678 11358 6638
rect 11358 678 11392 6638
rect 11392 678 11411 6638
rect 11499 678 11516 6638
rect 11516 678 11550 6638
rect 11550 678 11569 6638
rect 11657 678 11674 6638
rect 11674 678 11708 6638
rect 11708 678 11727 6638
rect 11815 678 11832 6638
rect 11832 678 11866 6638
rect 11866 678 11885 6638
rect 11973 678 11990 6638
rect 11990 678 12024 6638
rect 12024 678 12043 6638
rect 12131 678 12148 6638
rect 12148 678 12182 6638
rect 12182 678 12201 6638
rect 12289 678 12306 6638
rect 12306 678 12340 6638
rect 12340 678 12359 6638
rect 12447 678 12464 6638
rect 12464 678 12498 6638
rect 12498 678 12517 6638
rect 12605 678 12622 6638
rect 12622 678 12656 6638
rect 12656 678 12675 6638
rect 7730 500 7800 636
rect 12740 636 12754 6680
rect 12754 636 12792 6680
rect 12792 636 12810 6680
rect 7952 620 12586 626
rect 7952 586 8012 620
rect 8012 586 8102 620
rect 8102 586 8170 620
rect 8170 586 8260 620
rect 8260 586 8328 620
rect 8328 586 8418 620
rect 8418 586 8486 620
rect 8486 586 8576 620
rect 8576 586 8644 620
rect 8644 586 8734 620
rect 8734 586 8802 620
rect 8802 586 8892 620
rect 8892 586 8960 620
rect 8960 586 9050 620
rect 9050 586 9118 620
rect 9118 586 9208 620
rect 9208 586 9276 620
rect 9276 586 9366 620
rect 9366 586 9434 620
rect 9434 586 9524 620
rect 9524 586 9592 620
rect 9592 586 9682 620
rect 9682 586 9750 620
rect 9750 586 9840 620
rect 9840 586 9908 620
rect 9908 586 9998 620
rect 9998 586 10066 620
rect 10066 586 10156 620
rect 10156 586 10224 620
rect 10224 586 10314 620
rect 10314 586 10382 620
rect 10382 586 10472 620
rect 10472 586 10540 620
rect 10540 586 10630 620
rect 10630 586 10698 620
rect 10698 586 10788 620
rect 10788 586 10856 620
rect 10856 586 10946 620
rect 10946 586 11014 620
rect 11014 586 11104 620
rect 11104 586 11172 620
rect 11172 586 11262 620
rect 11262 586 11330 620
rect 11330 586 11420 620
rect 11420 586 11488 620
rect 11488 586 11578 620
rect 11578 586 11646 620
rect 11646 586 11736 620
rect 11736 586 11804 620
rect 11804 586 11894 620
rect 11894 586 11962 620
rect 11962 586 12052 620
rect 12052 586 12120 620
rect 12120 586 12210 620
rect 12210 586 12278 620
rect 12278 586 12368 620
rect 12368 586 12436 620
rect 12436 586 12526 620
rect 12526 586 12586 620
rect 7952 526 12586 586
rect 12740 500 12810 636
rect 14030 6680 14100 6820
rect 14252 6730 18886 6790
rect 14252 6696 14312 6730
rect 14312 6696 14402 6730
rect 14402 6696 14470 6730
rect 14470 6696 14560 6730
rect 14560 6696 14628 6730
rect 14628 6696 14718 6730
rect 14718 6696 14786 6730
rect 14786 6696 14876 6730
rect 14876 6696 14944 6730
rect 14944 6696 15034 6730
rect 15034 6696 15102 6730
rect 15102 6696 15192 6730
rect 15192 6696 15260 6730
rect 15260 6696 15350 6730
rect 15350 6696 15418 6730
rect 15418 6696 15508 6730
rect 15508 6696 15576 6730
rect 15576 6696 15666 6730
rect 15666 6696 15734 6730
rect 15734 6696 15824 6730
rect 15824 6696 15892 6730
rect 15892 6696 15982 6730
rect 15982 6696 16050 6730
rect 16050 6696 16140 6730
rect 16140 6696 16208 6730
rect 16208 6696 16298 6730
rect 16298 6696 16366 6730
rect 16366 6696 16456 6730
rect 16456 6696 16524 6730
rect 16524 6696 16614 6730
rect 16614 6696 16682 6730
rect 16682 6696 16772 6730
rect 16772 6696 16840 6730
rect 16840 6696 16930 6730
rect 16930 6696 16998 6730
rect 16998 6696 17088 6730
rect 17088 6696 17156 6730
rect 17156 6696 17246 6730
rect 17246 6696 17314 6730
rect 17314 6696 17404 6730
rect 17404 6696 17472 6730
rect 17472 6696 17562 6730
rect 17562 6696 17630 6730
rect 17630 6696 17720 6730
rect 17720 6696 17788 6730
rect 17788 6696 17878 6730
rect 17878 6696 17946 6730
rect 17946 6696 18036 6730
rect 18036 6696 18104 6730
rect 18104 6696 18194 6730
rect 18194 6696 18262 6730
rect 18262 6696 18352 6730
rect 18352 6696 18420 6730
rect 18420 6696 18510 6730
rect 18510 6696 18578 6730
rect 18578 6696 18668 6730
rect 18668 6696 18736 6730
rect 18736 6696 18826 6730
rect 18826 6696 18886 6730
rect 14252 6690 18886 6696
rect 14030 636 14046 6680
rect 14046 636 14084 6680
rect 14084 636 14100 6680
rect 19040 6680 19110 6820
rect 14165 678 14182 6638
rect 14182 678 14216 6638
rect 14216 678 14235 6638
rect 14323 678 14340 6638
rect 14340 678 14374 6638
rect 14374 678 14393 6638
rect 14481 678 14498 6638
rect 14498 678 14532 6638
rect 14532 678 14551 6638
rect 14639 678 14656 6638
rect 14656 678 14690 6638
rect 14690 678 14709 6638
rect 14797 678 14814 6638
rect 14814 678 14848 6638
rect 14848 678 14867 6638
rect 14955 678 14972 6638
rect 14972 678 15006 6638
rect 15006 678 15025 6638
rect 15113 678 15130 6638
rect 15130 678 15164 6638
rect 15164 678 15183 6638
rect 15271 678 15288 6638
rect 15288 678 15322 6638
rect 15322 678 15341 6638
rect 15429 678 15446 6638
rect 15446 678 15480 6638
rect 15480 678 15499 6638
rect 15587 678 15604 6638
rect 15604 678 15638 6638
rect 15638 678 15657 6638
rect 15745 678 15762 6638
rect 15762 678 15796 6638
rect 15796 678 15815 6638
rect 15903 678 15920 6638
rect 15920 678 15954 6638
rect 15954 678 15973 6638
rect 16061 678 16078 6638
rect 16078 678 16112 6638
rect 16112 678 16131 6638
rect 16219 678 16236 6638
rect 16236 678 16270 6638
rect 16270 678 16289 6638
rect 16377 678 16394 6638
rect 16394 678 16428 6638
rect 16428 678 16447 6638
rect 16535 678 16552 6638
rect 16552 678 16586 6638
rect 16586 678 16605 6638
rect 16693 678 16710 6638
rect 16710 678 16744 6638
rect 16744 678 16763 6638
rect 16851 678 16868 6638
rect 16868 678 16902 6638
rect 16902 678 16921 6638
rect 17009 678 17026 6638
rect 17026 678 17060 6638
rect 17060 678 17079 6638
rect 17167 678 17184 6638
rect 17184 678 17218 6638
rect 17218 678 17237 6638
rect 17325 678 17342 6638
rect 17342 678 17376 6638
rect 17376 678 17395 6638
rect 17483 678 17500 6638
rect 17500 678 17534 6638
rect 17534 678 17553 6638
rect 17641 678 17658 6638
rect 17658 678 17692 6638
rect 17692 678 17711 6638
rect 17799 678 17816 6638
rect 17816 678 17850 6638
rect 17850 678 17869 6638
rect 17957 678 17974 6638
rect 17974 678 18008 6638
rect 18008 678 18027 6638
rect 18115 678 18132 6638
rect 18132 678 18166 6638
rect 18166 678 18185 6638
rect 18273 678 18290 6638
rect 18290 678 18324 6638
rect 18324 678 18343 6638
rect 18431 678 18448 6638
rect 18448 678 18482 6638
rect 18482 678 18501 6638
rect 18589 678 18606 6638
rect 18606 678 18640 6638
rect 18640 678 18659 6638
rect 18747 678 18764 6638
rect 18764 678 18798 6638
rect 18798 678 18817 6638
rect 18905 678 18922 6638
rect 18922 678 18956 6638
rect 18956 678 18975 6638
rect 14030 500 14100 636
rect 19040 636 19054 6680
rect 19054 636 19092 6680
rect 19092 636 19110 6680
rect 14252 620 18886 626
rect 14252 586 14312 620
rect 14312 586 14402 620
rect 14402 586 14470 620
rect 14470 586 14560 620
rect 14560 586 14628 620
rect 14628 586 14718 620
rect 14718 586 14786 620
rect 14786 586 14876 620
rect 14876 586 14944 620
rect 14944 586 15034 620
rect 15034 586 15102 620
rect 15102 586 15192 620
rect 15192 586 15260 620
rect 15260 586 15350 620
rect 15350 586 15418 620
rect 15418 586 15508 620
rect 15508 586 15576 620
rect 15576 586 15666 620
rect 15666 586 15734 620
rect 15734 586 15824 620
rect 15824 586 15892 620
rect 15892 586 15982 620
rect 15982 586 16050 620
rect 16050 586 16140 620
rect 16140 586 16208 620
rect 16208 586 16298 620
rect 16298 586 16366 620
rect 16366 586 16456 620
rect 16456 586 16524 620
rect 16524 586 16614 620
rect 16614 586 16682 620
rect 16682 586 16772 620
rect 16772 586 16840 620
rect 16840 586 16930 620
rect 16930 586 16998 620
rect 16998 586 17088 620
rect 17088 586 17156 620
rect 17156 586 17246 620
rect 17246 586 17314 620
rect 17314 586 17404 620
rect 17404 586 17472 620
rect 17472 586 17562 620
rect 17562 586 17630 620
rect 17630 586 17720 620
rect 17720 586 17788 620
rect 17788 586 17878 620
rect 17878 586 17946 620
rect 17946 586 18036 620
rect 18036 586 18104 620
rect 18104 586 18194 620
rect 18194 586 18262 620
rect 18262 586 18352 620
rect 18352 586 18420 620
rect 18420 586 18510 620
rect 18510 586 18578 620
rect 18578 586 18668 620
rect 18668 586 18736 620
rect 18736 586 18826 620
rect 18826 586 18886 620
rect 14252 526 18886 586
rect 19040 500 19110 636
rect 20330 6680 20400 6820
rect 20552 6730 25186 6790
rect 20552 6696 20612 6730
rect 20612 6696 20702 6730
rect 20702 6696 20770 6730
rect 20770 6696 20860 6730
rect 20860 6696 20928 6730
rect 20928 6696 21018 6730
rect 21018 6696 21086 6730
rect 21086 6696 21176 6730
rect 21176 6696 21244 6730
rect 21244 6696 21334 6730
rect 21334 6696 21402 6730
rect 21402 6696 21492 6730
rect 21492 6696 21560 6730
rect 21560 6696 21650 6730
rect 21650 6696 21718 6730
rect 21718 6696 21808 6730
rect 21808 6696 21876 6730
rect 21876 6696 21966 6730
rect 21966 6696 22034 6730
rect 22034 6696 22124 6730
rect 22124 6696 22192 6730
rect 22192 6696 22282 6730
rect 22282 6696 22350 6730
rect 22350 6696 22440 6730
rect 22440 6696 22508 6730
rect 22508 6696 22598 6730
rect 22598 6696 22666 6730
rect 22666 6696 22756 6730
rect 22756 6696 22824 6730
rect 22824 6696 22914 6730
rect 22914 6696 22982 6730
rect 22982 6696 23072 6730
rect 23072 6696 23140 6730
rect 23140 6696 23230 6730
rect 23230 6696 23298 6730
rect 23298 6696 23388 6730
rect 23388 6696 23456 6730
rect 23456 6696 23546 6730
rect 23546 6696 23614 6730
rect 23614 6696 23704 6730
rect 23704 6696 23772 6730
rect 23772 6696 23862 6730
rect 23862 6696 23930 6730
rect 23930 6696 24020 6730
rect 24020 6696 24088 6730
rect 24088 6696 24178 6730
rect 24178 6696 24246 6730
rect 24246 6696 24336 6730
rect 24336 6696 24404 6730
rect 24404 6696 24494 6730
rect 24494 6696 24562 6730
rect 24562 6696 24652 6730
rect 24652 6696 24720 6730
rect 24720 6696 24810 6730
rect 24810 6696 24878 6730
rect 24878 6696 24968 6730
rect 24968 6696 25036 6730
rect 25036 6696 25126 6730
rect 25126 6696 25186 6730
rect 20552 6690 25186 6696
rect 20330 636 20346 6680
rect 20346 636 20384 6680
rect 20384 636 20400 6680
rect 25340 6680 25410 6820
rect 20465 678 20482 6638
rect 20482 678 20516 6638
rect 20516 678 20535 6638
rect 20623 678 20640 6638
rect 20640 678 20674 6638
rect 20674 678 20693 6638
rect 20781 678 20798 6638
rect 20798 678 20832 6638
rect 20832 678 20851 6638
rect 20939 678 20956 6638
rect 20956 678 20990 6638
rect 20990 678 21009 6638
rect 21097 678 21114 6638
rect 21114 678 21148 6638
rect 21148 678 21167 6638
rect 21255 678 21272 6638
rect 21272 678 21306 6638
rect 21306 678 21325 6638
rect 21413 678 21430 6638
rect 21430 678 21464 6638
rect 21464 678 21483 6638
rect 21571 678 21588 6638
rect 21588 678 21622 6638
rect 21622 678 21641 6638
rect 21729 678 21746 6638
rect 21746 678 21780 6638
rect 21780 678 21799 6638
rect 21887 678 21904 6638
rect 21904 678 21938 6638
rect 21938 678 21957 6638
rect 22045 678 22062 6638
rect 22062 678 22096 6638
rect 22096 678 22115 6638
rect 22203 678 22220 6638
rect 22220 678 22254 6638
rect 22254 678 22273 6638
rect 22361 678 22378 6638
rect 22378 678 22412 6638
rect 22412 678 22431 6638
rect 22519 678 22536 6638
rect 22536 678 22570 6638
rect 22570 678 22589 6638
rect 22677 678 22694 6638
rect 22694 678 22728 6638
rect 22728 678 22747 6638
rect 22835 678 22852 6638
rect 22852 678 22886 6638
rect 22886 678 22905 6638
rect 22993 678 23010 6638
rect 23010 678 23044 6638
rect 23044 678 23063 6638
rect 23151 678 23168 6638
rect 23168 678 23202 6638
rect 23202 678 23221 6638
rect 23309 678 23326 6638
rect 23326 678 23360 6638
rect 23360 678 23379 6638
rect 23467 678 23484 6638
rect 23484 678 23518 6638
rect 23518 678 23537 6638
rect 23625 678 23642 6638
rect 23642 678 23676 6638
rect 23676 678 23695 6638
rect 23783 678 23800 6638
rect 23800 678 23834 6638
rect 23834 678 23853 6638
rect 23941 678 23958 6638
rect 23958 678 23992 6638
rect 23992 678 24011 6638
rect 24099 678 24116 6638
rect 24116 678 24150 6638
rect 24150 678 24169 6638
rect 24257 678 24274 6638
rect 24274 678 24308 6638
rect 24308 678 24327 6638
rect 24415 678 24432 6638
rect 24432 678 24466 6638
rect 24466 678 24485 6638
rect 24573 678 24590 6638
rect 24590 678 24624 6638
rect 24624 678 24643 6638
rect 24731 678 24748 6638
rect 24748 678 24782 6638
rect 24782 678 24801 6638
rect 24889 678 24906 6638
rect 24906 678 24940 6638
rect 24940 678 24959 6638
rect 25047 678 25064 6638
rect 25064 678 25098 6638
rect 25098 678 25117 6638
rect 25205 678 25222 6638
rect 25222 678 25256 6638
rect 25256 678 25275 6638
rect 20330 500 20400 636
rect 25340 636 25354 6680
rect 25354 636 25392 6680
rect 25392 636 25410 6680
rect 20552 620 25186 626
rect 20552 586 20612 620
rect 20612 586 20702 620
rect 20702 586 20770 620
rect 20770 586 20860 620
rect 20860 586 20928 620
rect 20928 586 21018 620
rect 21018 586 21086 620
rect 21086 586 21176 620
rect 21176 586 21244 620
rect 21244 586 21334 620
rect 21334 586 21402 620
rect 21402 586 21492 620
rect 21492 586 21560 620
rect 21560 586 21650 620
rect 21650 586 21718 620
rect 21718 586 21808 620
rect 21808 586 21876 620
rect 21876 586 21966 620
rect 21966 586 22034 620
rect 22034 586 22124 620
rect 22124 586 22192 620
rect 22192 586 22282 620
rect 22282 586 22350 620
rect 22350 586 22440 620
rect 22440 586 22508 620
rect 22508 586 22598 620
rect 22598 586 22666 620
rect 22666 586 22756 620
rect 22756 586 22824 620
rect 22824 586 22914 620
rect 22914 586 22982 620
rect 22982 586 23072 620
rect 23072 586 23140 620
rect 23140 586 23230 620
rect 23230 586 23298 620
rect 23298 586 23388 620
rect 23388 586 23456 620
rect 23456 586 23546 620
rect 23546 586 23614 620
rect 23614 586 23704 620
rect 23704 586 23772 620
rect 23772 586 23862 620
rect 23862 586 23930 620
rect 23930 586 24020 620
rect 24020 586 24088 620
rect 24088 586 24178 620
rect 24178 586 24246 620
rect 24246 586 24336 620
rect 24336 586 24404 620
rect 24404 586 24494 620
rect 24494 586 24562 620
rect 24562 586 24652 620
rect 24652 586 24720 620
rect 24720 586 24810 620
rect 24810 586 24878 620
rect 24878 586 24968 620
rect 24968 586 25036 620
rect 25036 586 25126 620
rect 25126 586 25186 620
rect 20552 526 25186 586
rect 25340 500 25410 636
rect 1430 -920 1500 -780
rect 1652 -870 6286 -810
rect 1652 -904 1712 -870
rect 1712 -904 1802 -870
rect 1802 -904 1870 -870
rect 1870 -904 1960 -870
rect 1960 -904 2028 -870
rect 2028 -904 2118 -870
rect 2118 -904 2186 -870
rect 2186 -904 2276 -870
rect 2276 -904 2344 -870
rect 2344 -904 2434 -870
rect 2434 -904 2502 -870
rect 2502 -904 2592 -870
rect 2592 -904 2660 -870
rect 2660 -904 2750 -870
rect 2750 -904 2818 -870
rect 2818 -904 2908 -870
rect 2908 -904 2976 -870
rect 2976 -904 3066 -870
rect 3066 -904 3134 -870
rect 3134 -904 3224 -870
rect 3224 -904 3292 -870
rect 3292 -904 3382 -870
rect 3382 -904 3450 -870
rect 3450 -904 3540 -870
rect 3540 -904 3608 -870
rect 3608 -904 3698 -870
rect 3698 -904 3766 -870
rect 3766 -904 3856 -870
rect 3856 -904 3924 -870
rect 3924 -904 4014 -870
rect 4014 -904 4082 -870
rect 4082 -904 4172 -870
rect 4172 -904 4240 -870
rect 4240 -904 4330 -870
rect 4330 -904 4398 -870
rect 4398 -904 4488 -870
rect 4488 -904 4556 -870
rect 4556 -904 4646 -870
rect 4646 -904 4714 -870
rect 4714 -904 4804 -870
rect 4804 -904 4872 -870
rect 4872 -904 4962 -870
rect 4962 -904 5030 -870
rect 5030 -904 5120 -870
rect 5120 -904 5188 -870
rect 5188 -904 5278 -870
rect 5278 -904 5346 -870
rect 5346 -904 5436 -870
rect 5436 -904 5504 -870
rect 5504 -904 5594 -870
rect 5594 -904 5662 -870
rect 5662 -904 5752 -870
rect 5752 -904 5820 -870
rect 5820 -904 5910 -870
rect 5910 -904 5978 -870
rect 5978 -904 6068 -870
rect 6068 -904 6136 -870
rect 6136 -904 6226 -870
rect 6226 -904 6286 -870
rect 1652 -910 6286 -904
rect 1430 -6964 1446 -920
rect 1446 -6964 1484 -920
rect 1484 -6964 1500 -920
rect 6440 -920 6510 -780
rect 1565 -6922 1582 -962
rect 1582 -6922 1616 -962
rect 1616 -6922 1635 -962
rect 1723 -6922 1740 -962
rect 1740 -6922 1774 -962
rect 1774 -6922 1793 -962
rect 1881 -6922 1898 -962
rect 1898 -6922 1932 -962
rect 1932 -6922 1951 -962
rect 2039 -6922 2056 -962
rect 2056 -6922 2090 -962
rect 2090 -6922 2109 -962
rect 2197 -6922 2214 -962
rect 2214 -6922 2248 -962
rect 2248 -6922 2267 -962
rect 2355 -6922 2372 -962
rect 2372 -6922 2406 -962
rect 2406 -6922 2425 -962
rect 2513 -6922 2530 -962
rect 2530 -6922 2564 -962
rect 2564 -6922 2583 -962
rect 2671 -6922 2688 -962
rect 2688 -6922 2722 -962
rect 2722 -6922 2741 -962
rect 2829 -6922 2846 -962
rect 2846 -6922 2880 -962
rect 2880 -6922 2899 -962
rect 2987 -6922 3004 -962
rect 3004 -6922 3038 -962
rect 3038 -6922 3057 -962
rect 3145 -6922 3162 -962
rect 3162 -6922 3196 -962
rect 3196 -6922 3215 -962
rect 3303 -6922 3320 -962
rect 3320 -6922 3354 -962
rect 3354 -6922 3373 -962
rect 3461 -6922 3478 -962
rect 3478 -6922 3512 -962
rect 3512 -6922 3531 -962
rect 3619 -6922 3636 -962
rect 3636 -6922 3670 -962
rect 3670 -6922 3689 -962
rect 3777 -6922 3794 -962
rect 3794 -6922 3828 -962
rect 3828 -6922 3847 -962
rect 3935 -6922 3952 -962
rect 3952 -6922 3986 -962
rect 3986 -6922 4005 -962
rect 4093 -6922 4110 -962
rect 4110 -6922 4144 -962
rect 4144 -6922 4163 -962
rect 4251 -6922 4268 -962
rect 4268 -6922 4302 -962
rect 4302 -6922 4321 -962
rect 4409 -6922 4426 -962
rect 4426 -6922 4460 -962
rect 4460 -6922 4479 -962
rect 4567 -6922 4584 -962
rect 4584 -6922 4618 -962
rect 4618 -6922 4637 -962
rect 4725 -6922 4742 -962
rect 4742 -6922 4776 -962
rect 4776 -6922 4795 -962
rect 4883 -6922 4900 -962
rect 4900 -6922 4934 -962
rect 4934 -6922 4953 -962
rect 5041 -6922 5058 -962
rect 5058 -6922 5092 -962
rect 5092 -6922 5111 -962
rect 5199 -6922 5216 -962
rect 5216 -6922 5250 -962
rect 5250 -6922 5269 -962
rect 5357 -6922 5374 -962
rect 5374 -6922 5408 -962
rect 5408 -6922 5427 -962
rect 5515 -6922 5532 -962
rect 5532 -6922 5566 -962
rect 5566 -6922 5585 -962
rect 5673 -6922 5690 -962
rect 5690 -6922 5724 -962
rect 5724 -6922 5743 -962
rect 5831 -6922 5848 -962
rect 5848 -6922 5882 -962
rect 5882 -6922 5901 -962
rect 5989 -6922 6006 -962
rect 6006 -6922 6040 -962
rect 6040 -6922 6059 -962
rect 6147 -6922 6164 -962
rect 6164 -6922 6198 -962
rect 6198 -6922 6217 -962
rect 6305 -6922 6322 -962
rect 6322 -6922 6356 -962
rect 6356 -6922 6375 -962
rect 1430 -7100 1500 -6964
rect 6440 -6964 6454 -920
rect 6454 -6964 6492 -920
rect 6492 -6964 6510 -920
rect 1652 -6980 6286 -6974
rect 1652 -7014 1712 -6980
rect 1712 -7014 1802 -6980
rect 1802 -7014 1870 -6980
rect 1870 -7014 1960 -6980
rect 1960 -7014 2028 -6980
rect 2028 -7014 2118 -6980
rect 2118 -7014 2186 -6980
rect 2186 -7014 2276 -6980
rect 2276 -7014 2344 -6980
rect 2344 -7014 2434 -6980
rect 2434 -7014 2502 -6980
rect 2502 -7014 2592 -6980
rect 2592 -7014 2660 -6980
rect 2660 -7014 2750 -6980
rect 2750 -7014 2818 -6980
rect 2818 -7014 2908 -6980
rect 2908 -7014 2976 -6980
rect 2976 -7014 3066 -6980
rect 3066 -7014 3134 -6980
rect 3134 -7014 3224 -6980
rect 3224 -7014 3292 -6980
rect 3292 -7014 3382 -6980
rect 3382 -7014 3450 -6980
rect 3450 -7014 3540 -6980
rect 3540 -7014 3608 -6980
rect 3608 -7014 3698 -6980
rect 3698 -7014 3766 -6980
rect 3766 -7014 3856 -6980
rect 3856 -7014 3924 -6980
rect 3924 -7014 4014 -6980
rect 4014 -7014 4082 -6980
rect 4082 -7014 4172 -6980
rect 4172 -7014 4240 -6980
rect 4240 -7014 4330 -6980
rect 4330 -7014 4398 -6980
rect 4398 -7014 4488 -6980
rect 4488 -7014 4556 -6980
rect 4556 -7014 4646 -6980
rect 4646 -7014 4714 -6980
rect 4714 -7014 4804 -6980
rect 4804 -7014 4872 -6980
rect 4872 -7014 4962 -6980
rect 4962 -7014 5030 -6980
rect 5030 -7014 5120 -6980
rect 5120 -7014 5188 -6980
rect 5188 -7014 5278 -6980
rect 5278 -7014 5346 -6980
rect 5346 -7014 5436 -6980
rect 5436 -7014 5504 -6980
rect 5504 -7014 5594 -6980
rect 5594 -7014 5662 -6980
rect 5662 -7014 5752 -6980
rect 5752 -7014 5820 -6980
rect 5820 -7014 5910 -6980
rect 5910 -7014 5978 -6980
rect 5978 -7014 6068 -6980
rect 6068 -7014 6136 -6980
rect 6136 -7014 6226 -6980
rect 6226 -7014 6286 -6980
rect 1652 -7074 6286 -7014
rect 6440 -7100 6510 -6964
rect 7730 -920 7800 -780
rect 7952 -870 12586 -810
rect 7952 -904 8012 -870
rect 8012 -904 8102 -870
rect 8102 -904 8170 -870
rect 8170 -904 8260 -870
rect 8260 -904 8328 -870
rect 8328 -904 8418 -870
rect 8418 -904 8486 -870
rect 8486 -904 8576 -870
rect 8576 -904 8644 -870
rect 8644 -904 8734 -870
rect 8734 -904 8802 -870
rect 8802 -904 8892 -870
rect 8892 -904 8960 -870
rect 8960 -904 9050 -870
rect 9050 -904 9118 -870
rect 9118 -904 9208 -870
rect 9208 -904 9276 -870
rect 9276 -904 9366 -870
rect 9366 -904 9434 -870
rect 9434 -904 9524 -870
rect 9524 -904 9592 -870
rect 9592 -904 9682 -870
rect 9682 -904 9750 -870
rect 9750 -904 9840 -870
rect 9840 -904 9908 -870
rect 9908 -904 9998 -870
rect 9998 -904 10066 -870
rect 10066 -904 10156 -870
rect 10156 -904 10224 -870
rect 10224 -904 10314 -870
rect 10314 -904 10382 -870
rect 10382 -904 10472 -870
rect 10472 -904 10540 -870
rect 10540 -904 10630 -870
rect 10630 -904 10698 -870
rect 10698 -904 10788 -870
rect 10788 -904 10856 -870
rect 10856 -904 10946 -870
rect 10946 -904 11014 -870
rect 11014 -904 11104 -870
rect 11104 -904 11172 -870
rect 11172 -904 11262 -870
rect 11262 -904 11330 -870
rect 11330 -904 11420 -870
rect 11420 -904 11488 -870
rect 11488 -904 11578 -870
rect 11578 -904 11646 -870
rect 11646 -904 11736 -870
rect 11736 -904 11804 -870
rect 11804 -904 11894 -870
rect 11894 -904 11962 -870
rect 11962 -904 12052 -870
rect 12052 -904 12120 -870
rect 12120 -904 12210 -870
rect 12210 -904 12278 -870
rect 12278 -904 12368 -870
rect 12368 -904 12436 -870
rect 12436 -904 12526 -870
rect 12526 -904 12586 -870
rect 7952 -910 12586 -904
rect 7730 -6964 7746 -920
rect 7746 -6964 7784 -920
rect 7784 -6964 7800 -920
rect 12740 -920 12810 -780
rect 7865 -6922 7882 -962
rect 7882 -6922 7916 -962
rect 7916 -6922 7935 -962
rect 8023 -6922 8040 -962
rect 8040 -6922 8074 -962
rect 8074 -6922 8093 -962
rect 8181 -6922 8198 -962
rect 8198 -6922 8232 -962
rect 8232 -6922 8251 -962
rect 8339 -6922 8356 -962
rect 8356 -6922 8390 -962
rect 8390 -6922 8409 -962
rect 8497 -6922 8514 -962
rect 8514 -6922 8548 -962
rect 8548 -6922 8567 -962
rect 8655 -6922 8672 -962
rect 8672 -6922 8706 -962
rect 8706 -6922 8725 -962
rect 8813 -6922 8830 -962
rect 8830 -6922 8864 -962
rect 8864 -6922 8883 -962
rect 8971 -6922 8988 -962
rect 8988 -6922 9022 -962
rect 9022 -6922 9041 -962
rect 9129 -6922 9146 -962
rect 9146 -6922 9180 -962
rect 9180 -6922 9199 -962
rect 9287 -6922 9304 -962
rect 9304 -6922 9338 -962
rect 9338 -6922 9357 -962
rect 9445 -6922 9462 -962
rect 9462 -6922 9496 -962
rect 9496 -6922 9515 -962
rect 9603 -6922 9620 -962
rect 9620 -6922 9654 -962
rect 9654 -6922 9673 -962
rect 9761 -6922 9778 -962
rect 9778 -6922 9812 -962
rect 9812 -6922 9831 -962
rect 9919 -6922 9936 -962
rect 9936 -6922 9970 -962
rect 9970 -6922 9989 -962
rect 10077 -6922 10094 -962
rect 10094 -6922 10128 -962
rect 10128 -6922 10147 -962
rect 10235 -6922 10252 -962
rect 10252 -6922 10286 -962
rect 10286 -6922 10305 -962
rect 10393 -6922 10410 -962
rect 10410 -6922 10444 -962
rect 10444 -6922 10463 -962
rect 10551 -6922 10568 -962
rect 10568 -6922 10602 -962
rect 10602 -6922 10621 -962
rect 10709 -6922 10726 -962
rect 10726 -6922 10760 -962
rect 10760 -6922 10779 -962
rect 10867 -6922 10884 -962
rect 10884 -6922 10918 -962
rect 10918 -6922 10937 -962
rect 11025 -6922 11042 -962
rect 11042 -6922 11076 -962
rect 11076 -6922 11095 -962
rect 11183 -6922 11200 -962
rect 11200 -6922 11234 -962
rect 11234 -6922 11253 -962
rect 11341 -6922 11358 -962
rect 11358 -6922 11392 -962
rect 11392 -6922 11411 -962
rect 11499 -6922 11516 -962
rect 11516 -6922 11550 -962
rect 11550 -6922 11569 -962
rect 11657 -6922 11674 -962
rect 11674 -6922 11708 -962
rect 11708 -6922 11727 -962
rect 11815 -6922 11832 -962
rect 11832 -6922 11866 -962
rect 11866 -6922 11885 -962
rect 11973 -6922 11990 -962
rect 11990 -6922 12024 -962
rect 12024 -6922 12043 -962
rect 12131 -6922 12148 -962
rect 12148 -6922 12182 -962
rect 12182 -6922 12201 -962
rect 12289 -6922 12306 -962
rect 12306 -6922 12340 -962
rect 12340 -6922 12359 -962
rect 12447 -6922 12464 -962
rect 12464 -6922 12498 -962
rect 12498 -6922 12517 -962
rect 12605 -6922 12622 -962
rect 12622 -6922 12656 -962
rect 12656 -6922 12675 -962
rect 7730 -7100 7800 -6964
rect 12740 -6964 12754 -920
rect 12754 -6964 12792 -920
rect 12792 -6964 12810 -920
rect 7952 -6980 12586 -6974
rect 7952 -7014 8012 -6980
rect 8012 -7014 8102 -6980
rect 8102 -7014 8170 -6980
rect 8170 -7014 8260 -6980
rect 8260 -7014 8328 -6980
rect 8328 -7014 8418 -6980
rect 8418 -7014 8486 -6980
rect 8486 -7014 8576 -6980
rect 8576 -7014 8644 -6980
rect 8644 -7014 8734 -6980
rect 8734 -7014 8802 -6980
rect 8802 -7014 8892 -6980
rect 8892 -7014 8960 -6980
rect 8960 -7014 9050 -6980
rect 9050 -7014 9118 -6980
rect 9118 -7014 9208 -6980
rect 9208 -7014 9276 -6980
rect 9276 -7014 9366 -6980
rect 9366 -7014 9434 -6980
rect 9434 -7014 9524 -6980
rect 9524 -7014 9592 -6980
rect 9592 -7014 9682 -6980
rect 9682 -7014 9750 -6980
rect 9750 -7014 9840 -6980
rect 9840 -7014 9908 -6980
rect 9908 -7014 9998 -6980
rect 9998 -7014 10066 -6980
rect 10066 -7014 10156 -6980
rect 10156 -7014 10224 -6980
rect 10224 -7014 10314 -6980
rect 10314 -7014 10382 -6980
rect 10382 -7014 10472 -6980
rect 10472 -7014 10540 -6980
rect 10540 -7014 10630 -6980
rect 10630 -7014 10698 -6980
rect 10698 -7014 10788 -6980
rect 10788 -7014 10856 -6980
rect 10856 -7014 10946 -6980
rect 10946 -7014 11014 -6980
rect 11014 -7014 11104 -6980
rect 11104 -7014 11172 -6980
rect 11172 -7014 11262 -6980
rect 11262 -7014 11330 -6980
rect 11330 -7014 11420 -6980
rect 11420 -7014 11488 -6980
rect 11488 -7014 11578 -6980
rect 11578 -7014 11646 -6980
rect 11646 -7014 11736 -6980
rect 11736 -7014 11804 -6980
rect 11804 -7014 11894 -6980
rect 11894 -7014 11962 -6980
rect 11962 -7014 12052 -6980
rect 12052 -7014 12120 -6980
rect 12120 -7014 12210 -6980
rect 12210 -7014 12278 -6980
rect 12278 -7014 12368 -6980
rect 12368 -7014 12436 -6980
rect 12436 -7014 12526 -6980
rect 12526 -7014 12586 -6980
rect 7952 -7074 12586 -7014
rect 12740 -7100 12810 -6964
rect 14030 -920 14100 -780
rect 14252 -870 18886 -810
rect 14252 -904 14312 -870
rect 14312 -904 14402 -870
rect 14402 -904 14470 -870
rect 14470 -904 14560 -870
rect 14560 -904 14628 -870
rect 14628 -904 14718 -870
rect 14718 -904 14786 -870
rect 14786 -904 14876 -870
rect 14876 -904 14944 -870
rect 14944 -904 15034 -870
rect 15034 -904 15102 -870
rect 15102 -904 15192 -870
rect 15192 -904 15260 -870
rect 15260 -904 15350 -870
rect 15350 -904 15418 -870
rect 15418 -904 15508 -870
rect 15508 -904 15576 -870
rect 15576 -904 15666 -870
rect 15666 -904 15734 -870
rect 15734 -904 15824 -870
rect 15824 -904 15892 -870
rect 15892 -904 15982 -870
rect 15982 -904 16050 -870
rect 16050 -904 16140 -870
rect 16140 -904 16208 -870
rect 16208 -904 16298 -870
rect 16298 -904 16366 -870
rect 16366 -904 16456 -870
rect 16456 -904 16524 -870
rect 16524 -904 16614 -870
rect 16614 -904 16682 -870
rect 16682 -904 16772 -870
rect 16772 -904 16840 -870
rect 16840 -904 16930 -870
rect 16930 -904 16998 -870
rect 16998 -904 17088 -870
rect 17088 -904 17156 -870
rect 17156 -904 17246 -870
rect 17246 -904 17314 -870
rect 17314 -904 17404 -870
rect 17404 -904 17472 -870
rect 17472 -904 17562 -870
rect 17562 -904 17630 -870
rect 17630 -904 17720 -870
rect 17720 -904 17788 -870
rect 17788 -904 17878 -870
rect 17878 -904 17946 -870
rect 17946 -904 18036 -870
rect 18036 -904 18104 -870
rect 18104 -904 18194 -870
rect 18194 -904 18262 -870
rect 18262 -904 18352 -870
rect 18352 -904 18420 -870
rect 18420 -904 18510 -870
rect 18510 -904 18578 -870
rect 18578 -904 18668 -870
rect 18668 -904 18736 -870
rect 18736 -904 18826 -870
rect 18826 -904 18886 -870
rect 14252 -910 18886 -904
rect 14030 -6964 14046 -920
rect 14046 -6964 14084 -920
rect 14084 -6964 14100 -920
rect 19040 -920 19110 -780
rect 14165 -6922 14182 -962
rect 14182 -6922 14216 -962
rect 14216 -6922 14235 -962
rect 14323 -6922 14340 -962
rect 14340 -6922 14374 -962
rect 14374 -6922 14393 -962
rect 14481 -6922 14498 -962
rect 14498 -6922 14532 -962
rect 14532 -6922 14551 -962
rect 14639 -6922 14656 -962
rect 14656 -6922 14690 -962
rect 14690 -6922 14709 -962
rect 14797 -6922 14814 -962
rect 14814 -6922 14848 -962
rect 14848 -6922 14867 -962
rect 14955 -6922 14972 -962
rect 14972 -6922 15006 -962
rect 15006 -6922 15025 -962
rect 15113 -6922 15130 -962
rect 15130 -6922 15164 -962
rect 15164 -6922 15183 -962
rect 15271 -6922 15288 -962
rect 15288 -6922 15322 -962
rect 15322 -6922 15341 -962
rect 15429 -6922 15446 -962
rect 15446 -6922 15480 -962
rect 15480 -6922 15499 -962
rect 15587 -6922 15604 -962
rect 15604 -6922 15638 -962
rect 15638 -6922 15657 -962
rect 15745 -6922 15762 -962
rect 15762 -6922 15796 -962
rect 15796 -6922 15815 -962
rect 15903 -6922 15920 -962
rect 15920 -6922 15954 -962
rect 15954 -6922 15973 -962
rect 16061 -6922 16078 -962
rect 16078 -6922 16112 -962
rect 16112 -6922 16131 -962
rect 16219 -6922 16236 -962
rect 16236 -6922 16270 -962
rect 16270 -6922 16289 -962
rect 16377 -6922 16394 -962
rect 16394 -6922 16428 -962
rect 16428 -6922 16447 -962
rect 16535 -6922 16552 -962
rect 16552 -6922 16586 -962
rect 16586 -6922 16605 -962
rect 16693 -6922 16710 -962
rect 16710 -6922 16744 -962
rect 16744 -6922 16763 -962
rect 16851 -6922 16868 -962
rect 16868 -6922 16902 -962
rect 16902 -6922 16921 -962
rect 17009 -6922 17026 -962
rect 17026 -6922 17060 -962
rect 17060 -6922 17079 -962
rect 17167 -6922 17184 -962
rect 17184 -6922 17218 -962
rect 17218 -6922 17237 -962
rect 17325 -6922 17342 -962
rect 17342 -6922 17376 -962
rect 17376 -6922 17395 -962
rect 17483 -6922 17500 -962
rect 17500 -6922 17534 -962
rect 17534 -6922 17553 -962
rect 17641 -6922 17658 -962
rect 17658 -6922 17692 -962
rect 17692 -6922 17711 -962
rect 17799 -6922 17816 -962
rect 17816 -6922 17850 -962
rect 17850 -6922 17869 -962
rect 17957 -6922 17974 -962
rect 17974 -6922 18008 -962
rect 18008 -6922 18027 -962
rect 18115 -6922 18132 -962
rect 18132 -6922 18166 -962
rect 18166 -6922 18185 -962
rect 18273 -6922 18290 -962
rect 18290 -6922 18324 -962
rect 18324 -6922 18343 -962
rect 18431 -6922 18448 -962
rect 18448 -6922 18482 -962
rect 18482 -6922 18501 -962
rect 18589 -6922 18606 -962
rect 18606 -6922 18640 -962
rect 18640 -6922 18659 -962
rect 18747 -6922 18764 -962
rect 18764 -6922 18798 -962
rect 18798 -6922 18817 -962
rect 18905 -6922 18922 -962
rect 18922 -6922 18956 -962
rect 18956 -6922 18975 -962
rect 14030 -7100 14100 -6964
rect 19040 -6964 19054 -920
rect 19054 -6964 19092 -920
rect 19092 -6964 19110 -920
rect 14252 -6980 18886 -6974
rect 14252 -7014 14312 -6980
rect 14312 -7014 14402 -6980
rect 14402 -7014 14470 -6980
rect 14470 -7014 14560 -6980
rect 14560 -7014 14628 -6980
rect 14628 -7014 14718 -6980
rect 14718 -7014 14786 -6980
rect 14786 -7014 14876 -6980
rect 14876 -7014 14944 -6980
rect 14944 -7014 15034 -6980
rect 15034 -7014 15102 -6980
rect 15102 -7014 15192 -6980
rect 15192 -7014 15260 -6980
rect 15260 -7014 15350 -6980
rect 15350 -7014 15418 -6980
rect 15418 -7014 15508 -6980
rect 15508 -7014 15576 -6980
rect 15576 -7014 15666 -6980
rect 15666 -7014 15734 -6980
rect 15734 -7014 15824 -6980
rect 15824 -7014 15892 -6980
rect 15892 -7014 15982 -6980
rect 15982 -7014 16050 -6980
rect 16050 -7014 16140 -6980
rect 16140 -7014 16208 -6980
rect 16208 -7014 16298 -6980
rect 16298 -7014 16366 -6980
rect 16366 -7014 16456 -6980
rect 16456 -7014 16524 -6980
rect 16524 -7014 16614 -6980
rect 16614 -7014 16682 -6980
rect 16682 -7014 16772 -6980
rect 16772 -7014 16840 -6980
rect 16840 -7014 16930 -6980
rect 16930 -7014 16998 -6980
rect 16998 -7014 17088 -6980
rect 17088 -7014 17156 -6980
rect 17156 -7014 17246 -6980
rect 17246 -7014 17314 -6980
rect 17314 -7014 17404 -6980
rect 17404 -7014 17472 -6980
rect 17472 -7014 17562 -6980
rect 17562 -7014 17630 -6980
rect 17630 -7014 17720 -6980
rect 17720 -7014 17788 -6980
rect 17788 -7014 17878 -6980
rect 17878 -7014 17946 -6980
rect 17946 -7014 18036 -6980
rect 18036 -7014 18104 -6980
rect 18104 -7014 18194 -6980
rect 18194 -7014 18262 -6980
rect 18262 -7014 18352 -6980
rect 18352 -7014 18420 -6980
rect 18420 -7014 18510 -6980
rect 18510 -7014 18578 -6980
rect 18578 -7014 18668 -6980
rect 18668 -7014 18736 -6980
rect 18736 -7014 18826 -6980
rect 18826 -7014 18886 -6980
rect 14252 -7074 18886 -7014
rect 19040 -7100 19110 -6964
rect 20330 -920 20400 -780
rect 20552 -870 25186 -810
rect 20552 -904 20612 -870
rect 20612 -904 20702 -870
rect 20702 -904 20770 -870
rect 20770 -904 20860 -870
rect 20860 -904 20928 -870
rect 20928 -904 21018 -870
rect 21018 -904 21086 -870
rect 21086 -904 21176 -870
rect 21176 -904 21244 -870
rect 21244 -904 21334 -870
rect 21334 -904 21402 -870
rect 21402 -904 21492 -870
rect 21492 -904 21560 -870
rect 21560 -904 21650 -870
rect 21650 -904 21718 -870
rect 21718 -904 21808 -870
rect 21808 -904 21876 -870
rect 21876 -904 21966 -870
rect 21966 -904 22034 -870
rect 22034 -904 22124 -870
rect 22124 -904 22192 -870
rect 22192 -904 22282 -870
rect 22282 -904 22350 -870
rect 22350 -904 22440 -870
rect 22440 -904 22508 -870
rect 22508 -904 22598 -870
rect 22598 -904 22666 -870
rect 22666 -904 22756 -870
rect 22756 -904 22824 -870
rect 22824 -904 22914 -870
rect 22914 -904 22982 -870
rect 22982 -904 23072 -870
rect 23072 -904 23140 -870
rect 23140 -904 23230 -870
rect 23230 -904 23298 -870
rect 23298 -904 23388 -870
rect 23388 -904 23456 -870
rect 23456 -904 23546 -870
rect 23546 -904 23614 -870
rect 23614 -904 23704 -870
rect 23704 -904 23772 -870
rect 23772 -904 23862 -870
rect 23862 -904 23930 -870
rect 23930 -904 24020 -870
rect 24020 -904 24088 -870
rect 24088 -904 24178 -870
rect 24178 -904 24246 -870
rect 24246 -904 24336 -870
rect 24336 -904 24404 -870
rect 24404 -904 24494 -870
rect 24494 -904 24562 -870
rect 24562 -904 24652 -870
rect 24652 -904 24720 -870
rect 24720 -904 24810 -870
rect 24810 -904 24878 -870
rect 24878 -904 24968 -870
rect 24968 -904 25036 -870
rect 25036 -904 25126 -870
rect 25126 -904 25186 -870
rect 20552 -910 25186 -904
rect 20330 -6964 20346 -920
rect 20346 -6964 20384 -920
rect 20384 -6964 20400 -920
rect 25340 -920 25410 -780
rect 20465 -6922 20482 -962
rect 20482 -6922 20516 -962
rect 20516 -6922 20535 -962
rect 20623 -6922 20640 -962
rect 20640 -6922 20674 -962
rect 20674 -6922 20693 -962
rect 20781 -6922 20798 -962
rect 20798 -6922 20832 -962
rect 20832 -6922 20851 -962
rect 20939 -6922 20956 -962
rect 20956 -6922 20990 -962
rect 20990 -6922 21009 -962
rect 21097 -6922 21114 -962
rect 21114 -6922 21148 -962
rect 21148 -6922 21167 -962
rect 21255 -6922 21272 -962
rect 21272 -6922 21306 -962
rect 21306 -6922 21325 -962
rect 21413 -6922 21430 -962
rect 21430 -6922 21464 -962
rect 21464 -6922 21483 -962
rect 21571 -6922 21588 -962
rect 21588 -6922 21622 -962
rect 21622 -6922 21641 -962
rect 21729 -6922 21746 -962
rect 21746 -6922 21780 -962
rect 21780 -6922 21799 -962
rect 21887 -6922 21904 -962
rect 21904 -6922 21938 -962
rect 21938 -6922 21957 -962
rect 22045 -6922 22062 -962
rect 22062 -6922 22096 -962
rect 22096 -6922 22115 -962
rect 22203 -6922 22220 -962
rect 22220 -6922 22254 -962
rect 22254 -6922 22273 -962
rect 22361 -6922 22378 -962
rect 22378 -6922 22412 -962
rect 22412 -6922 22431 -962
rect 22519 -6922 22536 -962
rect 22536 -6922 22570 -962
rect 22570 -6922 22589 -962
rect 22677 -6922 22694 -962
rect 22694 -6922 22728 -962
rect 22728 -6922 22747 -962
rect 22835 -6922 22852 -962
rect 22852 -6922 22886 -962
rect 22886 -6922 22905 -962
rect 22993 -6922 23010 -962
rect 23010 -6922 23044 -962
rect 23044 -6922 23063 -962
rect 23151 -6922 23168 -962
rect 23168 -6922 23202 -962
rect 23202 -6922 23221 -962
rect 23309 -6922 23326 -962
rect 23326 -6922 23360 -962
rect 23360 -6922 23379 -962
rect 23467 -6922 23484 -962
rect 23484 -6922 23518 -962
rect 23518 -6922 23537 -962
rect 23625 -6922 23642 -962
rect 23642 -6922 23676 -962
rect 23676 -6922 23695 -962
rect 23783 -6922 23800 -962
rect 23800 -6922 23834 -962
rect 23834 -6922 23853 -962
rect 23941 -6922 23958 -962
rect 23958 -6922 23992 -962
rect 23992 -6922 24011 -962
rect 24099 -6922 24116 -962
rect 24116 -6922 24150 -962
rect 24150 -6922 24169 -962
rect 24257 -6922 24274 -962
rect 24274 -6922 24308 -962
rect 24308 -6922 24327 -962
rect 24415 -6922 24432 -962
rect 24432 -6922 24466 -962
rect 24466 -6922 24485 -962
rect 24573 -6922 24590 -962
rect 24590 -6922 24624 -962
rect 24624 -6922 24643 -962
rect 24731 -6922 24748 -962
rect 24748 -6922 24782 -962
rect 24782 -6922 24801 -962
rect 24889 -6922 24906 -962
rect 24906 -6922 24940 -962
rect 24940 -6922 24959 -962
rect 25047 -6922 25064 -962
rect 25064 -6922 25098 -962
rect 25098 -6922 25117 -962
rect 25205 -6922 25222 -962
rect 25222 -6922 25256 -962
rect 25256 -6922 25275 -962
rect 20330 -7100 20400 -6964
rect 25340 -6964 25354 -920
rect 25354 -6964 25392 -920
rect 25392 -6964 25410 -920
rect 20552 -6980 25186 -6974
rect 20552 -7014 20612 -6980
rect 20612 -7014 20702 -6980
rect 20702 -7014 20770 -6980
rect 20770 -7014 20860 -6980
rect 20860 -7014 20928 -6980
rect 20928 -7014 21018 -6980
rect 21018 -7014 21086 -6980
rect 21086 -7014 21176 -6980
rect 21176 -7014 21244 -6980
rect 21244 -7014 21334 -6980
rect 21334 -7014 21402 -6980
rect 21402 -7014 21492 -6980
rect 21492 -7014 21560 -6980
rect 21560 -7014 21650 -6980
rect 21650 -7014 21718 -6980
rect 21718 -7014 21808 -6980
rect 21808 -7014 21876 -6980
rect 21876 -7014 21966 -6980
rect 21966 -7014 22034 -6980
rect 22034 -7014 22124 -6980
rect 22124 -7014 22192 -6980
rect 22192 -7014 22282 -6980
rect 22282 -7014 22350 -6980
rect 22350 -7014 22440 -6980
rect 22440 -7014 22508 -6980
rect 22508 -7014 22598 -6980
rect 22598 -7014 22666 -6980
rect 22666 -7014 22756 -6980
rect 22756 -7014 22824 -6980
rect 22824 -7014 22914 -6980
rect 22914 -7014 22982 -6980
rect 22982 -7014 23072 -6980
rect 23072 -7014 23140 -6980
rect 23140 -7014 23230 -6980
rect 23230 -7014 23298 -6980
rect 23298 -7014 23388 -6980
rect 23388 -7014 23456 -6980
rect 23456 -7014 23546 -6980
rect 23546 -7014 23614 -6980
rect 23614 -7014 23704 -6980
rect 23704 -7014 23772 -6980
rect 23772 -7014 23862 -6980
rect 23862 -7014 23930 -6980
rect 23930 -7014 24020 -6980
rect 24020 -7014 24088 -6980
rect 24088 -7014 24178 -6980
rect 24178 -7014 24246 -6980
rect 24246 -7014 24336 -6980
rect 24336 -7014 24404 -6980
rect 24404 -7014 24494 -6980
rect 24494 -7014 24562 -6980
rect 24562 -7014 24652 -6980
rect 24652 -7014 24720 -6980
rect 24720 -7014 24810 -6980
rect 24810 -7014 24878 -6980
rect 24878 -7014 24968 -6980
rect 24968 -7014 25036 -6980
rect 25036 -7014 25126 -6980
rect 25126 -7014 25186 -6980
rect 20552 -7074 25186 -7014
rect 25340 -7100 25410 -6964
<< metal2 >>
rect 1430 6820 1500 6880
rect 6440 6820 6510 6880
rect 1632 6780 1652 6790
rect 6286 6780 6306 6790
rect 1632 6710 1640 6780
rect 6300 6710 6306 6780
rect 1632 6690 1652 6710
rect 6286 6690 6306 6710
rect 1565 6638 1635 6658
rect 1565 658 1635 678
rect 1723 6638 1793 6658
rect 1723 658 1793 678
rect 1881 6638 1951 6658
rect 1881 658 1951 678
rect 2039 6638 2109 6658
rect 2039 658 2109 678
rect 2197 6638 2267 6658
rect 2197 658 2267 678
rect 2355 6638 2425 6658
rect 2355 658 2425 678
rect 2513 6638 2583 6658
rect 2513 658 2583 678
rect 2671 6638 2741 6658
rect 2671 658 2741 678
rect 2829 6638 2899 6658
rect 2829 658 2899 678
rect 2987 6638 3057 6658
rect 2987 658 3057 678
rect 3145 6638 3215 6658
rect 3145 658 3215 678
rect 3303 6638 3373 6658
rect 3303 658 3373 678
rect 3461 6638 3531 6658
rect 3461 658 3531 678
rect 3619 6638 3689 6658
rect 3619 658 3689 678
rect 3777 6638 3847 6658
rect 3777 658 3847 678
rect 3935 6638 4005 6658
rect 3935 658 4005 678
rect 4093 6638 4163 6658
rect 4093 658 4163 678
rect 4251 6638 4321 6658
rect 4251 658 4321 678
rect 4409 6638 4479 6658
rect 4409 658 4479 678
rect 4567 6638 4637 6658
rect 4567 658 4637 678
rect 4725 6638 4795 6658
rect 4725 658 4795 678
rect 4883 6638 4953 6658
rect 4883 658 4953 678
rect 5041 6638 5111 6658
rect 5041 658 5111 678
rect 5199 6638 5269 6658
rect 5199 658 5269 678
rect 5357 6638 5427 6658
rect 5357 658 5427 678
rect 5515 6638 5585 6658
rect 5515 658 5585 678
rect 5673 6638 5743 6658
rect 5673 658 5743 678
rect 5831 6638 5901 6658
rect 5831 658 5901 678
rect 5989 6638 6059 6658
rect 5989 658 6059 678
rect 6147 6638 6217 6658
rect 6147 658 6217 678
rect 6305 6638 6375 6658
rect 6305 658 6375 678
rect 1632 610 1652 626
rect 6286 610 6306 626
rect 1632 540 1640 610
rect 6290 540 6306 610
rect 1632 526 1652 540
rect 6286 526 6306 540
rect 1430 430 1500 500
rect 7730 6820 7800 6880
rect 6510 6100 7730 6500
rect 6510 5500 7730 5900
rect 6510 4900 7730 5300
rect 6510 4300 7730 4700
rect 6510 3700 7730 4100
rect 6510 3100 7730 3500
rect 6510 2500 7730 2900
rect 6510 1900 7730 2300
rect 6510 1300 7730 1700
rect 6510 700 7730 1100
rect 12740 6820 12810 6880
rect 7932 6780 7952 6790
rect 12586 6780 12606 6790
rect 7932 6710 7940 6780
rect 12600 6710 12606 6780
rect 7932 6690 7952 6710
rect 12586 6690 12606 6710
rect 7865 6638 7935 6658
rect 7865 658 7935 678
rect 8023 6638 8093 6658
rect 8023 658 8093 678
rect 8181 6638 8251 6658
rect 8181 658 8251 678
rect 8339 6638 8409 6658
rect 8339 658 8409 678
rect 8497 6638 8567 6658
rect 8497 658 8567 678
rect 8655 6638 8725 6658
rect 8655 658 8725 678
rect 8813 6638 8883 6658
rect 8813 658 8883 678
rect 8971 6638 9041 6658
rect 8971 658 9041 678
rect 9129 6638 9199 6658
rect 9129 658 9199 678
rect 9287 6638 9357 6658
rect 9287 658 9357 678
rect 9445 6638 9515 6658
rect 9445 658 9515 678
rect 9603 6638 9673 6658
rect 9603 658 9673 678
rect 9761 6638 9831 6658
rect 9761 658 9831 678
rect 9919 6638 9989 6658
rect 9919 658 9989 678
rect 10077 6638 10147 6658
rect 10077 658 10147 678
rect 10235 6638 10305 6658
rect 10235 658 10305 678
rect 10393 6638 10463 6658
rect 10393 658 10463 678
rect 10551 6638 10621 6658
rect 10551 658 10621 678
rect 10709 6638 10779 6658
rect 10709 658 10779 678
rect 10867 6638 10937 6658
rect 10867 658 10937 678
rect 11025 6638 11095 6658
rect 11025 658 11095 678
rect 11183 6638 11253 6658
rect 11183 658 11253 678
rect 11341 6638 11411 6658
rect 11341 658 11411 678
rect 11499 6638 11569 6658
rect 11499 658 11569 678
rect 11657 6638 11727 6658
rect 11657 658 11727 678
rect 11815 6638 11885 6658
rect 11815 658 11885 678
rect 11973 6638 12043 6658
rect 11973 658 12043 678
rect 12131 6638 12201 6658
rect 12131 658 12201 678
rect 12289 6638 12359 6658
rect 12289 658 12359 678
rect 12447 6638 12517 6658
rect 12447 658 12517 678
rect 12605 6638 12675 6658
rect 12605 658 12675 678
rect 7932 610 7952 626
rect 12586 610 12606 626
rect 7932 540 7940 610
rect 12590 540 12606 610
rect 7932 526 7952 540
rect 12586 526 12606 540
rect 6440 430 7800 500
rect 14030 6820 14100 6880
rect 12810 6100 14030 6500
rect 12810 5500 14030 5900
rect 12810 4900 14030 5300
rect 12810 4300 14030 4700
rect 12810 3700 14030 4100
rect 12810 3100 14030 3500
rect 12810 2500 14030 2900
rect 12810 1900 14030 2300
rect 12810 1300 14030 1700
rect 12810 700 14030 1100
rect 19040 6820 19110 6880
rect 14232 6780 14252 6790
rect 18886 6780 18906 6790
rect 14232 6710 14240 6780
rect 18900 6710 18906 6780
rect 14232 6690 14252 6710
rect 18886 6690 18906 6710
rect 14165 6638 14235 6658
rect 14165 658 14235 678
rect 14323 6638 14393 6658
rect 14323 658 14393 678
rect 14481 6638 14551 6658
rect 14481 658 14551 678
rect 14639 6638 14709 6658
rect 14639 658 14709 678
rect 14797 6638 14867 6658
rect 14797 658 14867 678
rect 14955 6638 15025 6658
rect 14955 658 15025 678
rect 15113 6638 15183 6658
rect 15113 658 15183 678
rect 15271 6638 15341 6658
rect 15271 658 15341 678
rect 15429 6638 15499 6658
rect 15429 658 15499 678
rect 15587 6638 15657 6658
rect 15587 658 15657 678
rect 15745 6638 15815 6658
rect 15745 658 15815 678
rect 15903 6638 15973 6658
rect 15903 658 15973 678
rect 16061 6638 16131 6658
rect 16061 658 16131 678
rect 16219 6638 16289 6658
rect 16219 658 16289 678
rect 16377 6638 16447 6658
rect 16377 658 16447 678
rect 16535 6638 16605 6658
rect 16535 658 16605 678
rect 16693 6638 16763 6658
rect 16693 658 16763 678
rect 16851 6638 16921 6658
rect 16851 658 16921 678
rect 17009 6638 17079 6658
rect 17009 658 17079 678
rect 17167 6638 17237 6658
rect 17167 658 17237 678
rect 17325 6638 17395 6658
rect 17325 658 17395 678
rect 17483 6638 17553 6658
rect 17483 658 17553 678
rect 17641 6638 17711 6658
rect 17641 658 17711 678
rect 17799 6638 17869 6658
rect 17799 658 17869 678
rect 17957 6638 18027 6658
rect 17957 658 18027 678
rect 18115 6638 18185 6658
rect 18115 658 18185 678
rect 18273 6638 18343 6658
rect 18273 658 18343 678
rect 18431 6638 18501 6658
rect 18431 658 18501 678
rect 18589 6638 18659 6658
rect 18589 658 18659 678
rect 18747 6638 18817 6658
rect 18747 658 18817 678
rect 18905 6638 18975 6658
rect 18905 658 18975 678
rect 14232 610 14252 626
rect 18886 610 18906 626
rect 14232 540 14240 610
rect 18890 540 18906 610
rect 14232 526 14252 540
rect 18886 526 18906 540
rect 12740 430 14100 500
rect 20330 6820 20400 6880
rect 19110 6100 20330 6500
rect 19110 5500 20330 5900
rect 19110 4900 20330 5300
rect 19110 4300 20330 4700
rect 19110 3700 20330 4100
rect 19110 3100 20330 3500
rect 19110 2500 20330 2900
rect 19110 1900 20330 2300
rect 19110 1300 20330 1700
rect 19110 700 20330 1100
rect 25340 6820 25410 6880
rect 20532 6780 20552 6790
rect 25186 6780 25206 6790
rect 20532 6710 20540 6780
rect 25200 6710 25206 6780
rect 20532 6690 20552 6710
rect 25186 6690 25206 6710
rect 20465 6638 20535 6658
rect 20465 658 20535 678
rect 20623 6638 20693 6658
rect 20623 658 20693 678
rect 20781 6638 20851 6658
rect 20781 658 20851 678
rect 20939 6638 21009 6658
rect 20939 658 21009 678
rect 21097 6638 21167 6658
rect 21097 658 21167 678
rect 21255 6638 21325 6658
rect 21255 658 21325 678
rect 21413 6638 21483 6658
rect 21413 658 21483 678
rect 21571 6638 21641 6658
rect 21571 658 21641 678
rect 21729 6638 21799 6658
rect 21729 658 21799 678
rect 21887 6638 21957 6658
rect 21887 658 21957 678
rect 22045 6638 22115 6658
rect 22045 658 22115 678
rect 22203 6638 22273 6658
rect 22203 658 22273 678
rect 22361 6638 22431 6658
rect 22361 658 22431 678
rect 22519 6638 22589 6658
rect 22519 658 22589 678
rect 22677 6638 22747 6658
rect 22677 658 22747 678
rect 22835 6638 22905 6658
rect 22835 658 22905 678
rect 22993 6638 23063 6658
rect 22993 658 23063 678
rect 23151 6638 23221 6658
rect 23151 658 23221 678
rect 23309 6638 23379 6658
rect 23309 658 23379 678
rect 23467 6638 23537 6658
rect 23467 658 23537 678
rect 23625 6638 23695 6658
rect 23625 658 23695 678
rect 23783 6638 23853 6658
rect 23783 658 23853 678
rect 23941 6638 24011 6658
rect 23941 658 24011 678
rect 24099 6638 24169 6658
rect 24099 658 24169 678
rect 24257 6638 24327 6658
rect 24257 658 24327 678
rect 24415 6638 24485 6658
rect 24415 658 24485 678
rect 24573 6638 24643 6658
rect 24573 658 24643 678
rect 24731 6638 24801 6658
rect 24731 658 24801 678
rect 24889 6638 24959 6658
rect 24889 658 24959 678
rect 25047 6638 25117 6658
rect 25047 658 25117 678
rect 25205 6638 25275 6658
rect 25205 658 25275 678
rect 20532 610 20552 626
rect 25186 610 25206 626
rect 20532 540 20540 610
rect 25190 540 25206 610
rect 20532 526 20552 540
rect 25186 526 25206 540
rect 19040 430 20400 500
rect 25340 430 25410 500
rect 6500 100 7800 430
rect 12800 100 14100 430
rect 19100 100 20400 430
rect 6900 -500 7400 100
rect 13200 -500 13700 100
rect 19500 -500 20000 100
rect 6500 -720 7800 -500
rect 12800 -720 14100 -500
rect 19100 -720 20400 -500
rect 1430 -780 1500 -720
rect 6440 -780 7800 -720
rect 1632 -820 1652 -810
rect 6286 -820 6306 -810
rect 1632 -890 1640 -820
rect 6300 -890 6306 -820
rect 1632 -910 1652 -890
rect 6286 -910 6306 -890
rect 1565 -962 1635 -942
rect 1565 -6942 1635 -6922
rect 1723 -962 1793 -942
rect 1723 -6942 1793 -6922
rect 1881 -962 1951 -942
rect 1881 -6942 1951 -6922
rect 2039 -962 2109 -942
rect 2039 -6942 2109 -6922
rect 2197 -962 2267 -942
rect 2197 -6942 2267 -6922
rect 2355 -962 2425 -942
rect 2355 -6942 2425 -6922
rect 2513 -962 2583 -942
rect 2513 -6942 2583 -6922
rect 2671 -962 2741 -942
rect 2671 -6942 2741 -6922
rect 2829 -962 2899 -942
rect 2829 -6942 2899 -6922
rect 2987 -962 3057 -942
rect 2987 -6942 3057 -6922
rect 3145 -962 3215 -942
rect 3145 -6942 3215 -6922
rect 3303 -962 3373 -942
rect 3303 -6942 3373 -6922
rect 3461 -962 3531 -942
rect 3461 -6942 3531 -6922
rect 3619 -962 3689 -942
rect 3619 -6942 3689 -6922
rect 3777 -962 3847 -942
rect 3777 -6942 3847 -6922
rect 3935 -962 4005 -942
rect 3935 -6942 4005 -6922
rect 4093 -962 4163 -942
rect 4093 -6942 4163 -6922
rect 4251 -962 4321 -942
rect 4251 -6942 4321 -6922
rect 4409 -962 4479 -942
rect 4409 -6942 4479 -6922
rect 4567 -962 4637 -942
rect 4567 -6942 4637 -6922
rect 4725 -962 4795 -942
rect 4725 -6942 4795 -6922
rect 4883 -962 4953 -942
rect 4883 -6942 4953 -6922
rect 5041 -962 5111 -942
rect 5041 -6942 5111 -6922
rect 5199 -962 5269 -942
rect 5199 -6942 5269 -6922
rect 5357 -962 5427 -942
rect 5357 -6942 5427 -6922
rect 5515 -962 5585 -942
rect 5515 -6942 5585 -6922
rect 5673 -962 5743 -942
rect 5673 -6942 5743 -6922
rect 5831 -962 5901 -942
rect 5831 -6942 5901 -6922
rect 5989 -962 6059 -942
rect 5989 -6942 6059 -6922
rect 6147 -962 6217 -942
rect 6147 -6942 6217 -6922
rect 6305 -962 6375 -942
rect 6305 -6942 6375 -6922
rect 1632 -6990 1652 -6974
rect 6286 -6990 6306 -6974
rect 1632 -7060 1640 -6990
rect 6290 -7060 6306 -6990
rect 1632 -7074 1652 -7060
rect 6286 -7074 6306 -7060
rect 1430 -7170 1500 -7100
rect 6510 -900 7730 -780
rect 6510 -1500 7730 -1100
rect 6510 -2100 7730 -1700
rect 6510 -2700 7730 -2300
rect 6510 -3300 7730 -2900
rect 6510 -3900 7730 -3500
rect 6510 -4500 7730 -4100
rect 6510 -5100 7730 -4700
rect 6510 -5700 7730 -5300
rect 6510 -6300 7730 -5900
rect 6510 -6900 7730 -6500
rect 6440 -7170 6510 -7100
rect 12740 -780 14100 -720
rect 7932 -820 7952 -810
rect 12586 -820 12606 -810
rect 7932 -890 7940 -820
rect 12600 -890 12606 -820
rect 7932 -910 7952 -890
rect 12586 -910 12606 -890
rect 7865 -962 7935 -942
rect 7865 -6942 7935 -6922
rect 8023 -962 8093 -942
rect 8023 -6942 8093 -6922
rect 8181 -962 8251 -942
rect 8181 -6942 8251 -6922
rect 8339 -962 8409 -942
rect 8339 -6942 8409 -6922
rect 8497 -962 8567 -942
rect 8497 -6942 8567 -6922
rect 8655 -962 8725 -942
rect 8655 -6942 8725 -6922
rect 8813 -962 8883 -942
rect 8813 -6942 8883 -6922
rect 8971 -962 9041 -942
rect 8971 -6942 9041 -6922
rect 9129 -962 9199 -942
rect 9129 -6942 9199 -6922
rect 9287 -962 9357 -942
rect 9287 -6942 9357 -6922
rect 9445 -962 9515 -942
rect 9445 -6942 9515 -6922
rect 9603 -962 9673 -942
rect 9603 -6942 9673 -6922
rect 9761 -962 9831 -942
rect 9761 -6942 9831 -6922
rect 9919 -962 9989 -942
rect 9919 -6942 9989 -6922
rect 10077 -962 10147 -942
rect 10077 -6942 10147 -6922
rect 10235 -962 10305 -942
rect 10235 -6942 10305 -6922
rect 10393 -962 10463 -942
rect 10393 -6942 10463 -6922
rect 10551 -962 10621 -942
rect 10551 -6942 10621 -6922
rect 10709 -962 10779 -942
rect 10709 -6942 10779 -6922
rect 10867 -962 10937 -942
rect 10867 -6942 10937 -6922
rect 11025 -962 11095 -942
rect 11025 -6942 11095 -6922
rect 11183 -962 11253 -942
rect 11183 -6942 11253 -6922
rect 11341 -962 11411 -942
rect 11341 -6942 11411 -6922
rect 11499 -962 11569 -942
rect 11499 -6942 11569 -6922
rect 11657 -962 11727 -942
rect 11657 -6942 11727 -6922
rect 11815 -962 11885 -942
rect 11815 -6942 11885 -6922
rect 11973 -962 12043 -942
rect 11973 -6942 12043 -6922
rect 12131 -962 12201 -942
rect 12131 -6942 12201 -6922
rect 12289 -962 12359 -942
rect 12289 -6942 12359 -6922
rect 12447 -962 12517 -942
rect 12447 -6942 12517 -6922
rect 12605 -962 12675 -942
rect 12605 -6942 12675 -6922
rect 7932 -6990 7952 -6974
rect 12586 -6990 12606 -6974
rect 7932 -7060 7940 -6990
rect 12590 -7060 12606 -6990
rect 7932 -7074 7952 -7060
rect 12586 -7074 12606 -7060
rect 7730 -7170 7800 -7100
rect 12810 -900 14030 -780
rect 12810 -1500 14030 -1100
rect 12810 -2100 14030 -1700
rect 12810 -2700 14030 -2300
rect 12810 -3300 14030 -2900
rect 12810 -3900 14030 -3500
rect 12810 -4500 14030 -4100
rect 12810 -5100 14030 -4700
rect 12810 -5700 14030 -5300
rect 12810 -6300 14030 -5900
rect 12810 -6900 14030 -6500
rect 12740 -7170 12810 -7100
rect 19040 -780 20400 -720
rect 14232 -820 14252 -810
rect 18886 -820 18906 -810
rect 14232 -890 14240 -820
rect 18900 -890 18906 -820
rect 14232 -910 14252 -890
rect 18886 -910 18906 -890
rect 14165 -962 14235 -942
rect 14165 -6942 14235 -6922
rect 14323 -962 14393 -942
rect 14323 -6942 14393 -6922
rect 14481 -962 14551 -942
rect 14481 -6942 14551 -6922
rect 14639 -962 14709 -942
rect 14639 -6942 14709 -6922
rect 14797 -962 14867 -942
rect 14797 -6942 14867 -6922
rect 14955 -962 15025 -942
rect 14955 -6942 15025 -6922
rect 15113 -962 15183 -942
rect 15113 -6942 15183 -6922
rect 15271 -962 15341 -942
rect 15271 -6942 15341 -6922
rect 15429 -962 15499 -942
rect 15429 -6942 15499 -6922
rect 15587 -962 15657 -942
rect 15587 -6942 15657 -6922
rect 15745 -962 15815 -942
rect 15745 -6942 15815 -6922
rect 15903 -962 15973 -942
rect 15903 -6942 15973 -6922
rect 16061 -962 16131 -942
rect 16061 -6942 16131 -6922
rect 16219 -962 16289 -942
rect 16219 -6942 16289 -6922
rect 16377 -962 16447 -942
rect 16377 -6942 16447 -6922
rect 16535 -962 16605 -942
rect 16535 -6942 16605 -6922
rect 16693 -962 16763 -942
rect 16693 -6942 16763 -6922
rect 16851 -962 16921 -942
rect 16851 -6942 16921 -6922
rect 17009 -962 17079 -942
rect 17009 -6942 17079 -6922
rect 17167 -962 17237 -942
rect 17167 -6942 17237 -6922
rect 17325 -962 17395 -942
rect 17325 -6942 17395 -6922
rect 17483 -962 17553 -942
rect 17483 -6942 17553 -6922
rect 17641 -962 17711 -942
rect 17641 -6942 17711 -6922
rect 17799 -962 17869 -942
rect 17799 -6942 17869 -6922
rect 17957 -962 18027 -942
rect 17957 -6942 18027 -6922
rect 18115 -962 18185 -942
rect 18115 -6942 18185 -6922
rect 18273 -962 18343 -942
rect 18273 -6942 18343 -6922
rect 18431 -962 18501 -942
rect 18431 -6942 18501 -6922
rect 18589 -962 18659 -942
rect 18589 -6942 18659 -6922
rect 18747 -962 18817 -942
rect 18747 -6942 18817 -6922
rect 18905 -962 18975 -942
rect 18905 -6942 18975 -6922
rect 14232 -6990 14252 -6974
rect 18886 -6990 18906 -6974
rect 14232 -7060 14240 -6990
rect 18890 -7060 18906 -6990
rect 14232 -7074 14252 -7060
rect 18886 -7074 18906 -7060
rect 14030 -7170 14100 -7100
rect 19110 -900 20330 -780
rect 19110 -1500 20330 -1100
rect 19110 -2100 20330 -1700
rect 19110 -2700 20330 -2300
rect 19110 -3300 20330 -2900
rect 19110 -3900 20330 -3500
rect 19110 -4500 20330 -4100
rect 19110 -5100 20330 -4700
rect 19110 -5700 20330 -5300
rect 19110 -6300 20330 -5900
rect 19110 -6900 20330 -6500
rect 19040 -7170 19110 -7100
rect 25340 -780 25410 -720
rect 20532 -820 20552 -810
rect 25186 -820 25206 -810
rect 20532 -890 20540 -820
rect 25200 -890 25206 -820
rect 20532 -910 20552 -890
rect 25186 -910 25206 -890
rect 20465 -962 20535 -942
rect 20465 -6942 20535 -6922
rect 20623 -962 20693 -942
rect 20623 -6942 20693 -6922
rect 20781 -962 20851 -942
rect 20781 -6942 20851 -6922
rect 20939 -962 21009 -942
rect 20939 -6942 21009 -6922
rect 21097 -962 21167 -942
rect 21097 -6942 21167 -6922
rect 21255 -962 21325 -942
rect 21255 -6942 21325 -6922
rect 21413 -962 21483 -942
rect 21413 -6942 21483 -6922
rect 21571 -962 21641 -942
rect 21571 -6942 21641 -6922
rect 21729 -962 21799 -942
rect 21729 -6942 21799 -6922
rect 21887 -962 21957 -942
rect 21887 -6942 21957 -6922
rect 22045 -962 22115 -942
rect 22045 -6942 22115 -6922
rect 22203 -962 22273 -942
rect 22203 -6942 22273 -6922
rect 22361 -962 22431 -942
rect 22361 -6942 22431 -6922
rect 22519 -962 22589 -942
rect 22519 -6942 22589 -6922
rect 22677 -962 22747 -942
rect 22677 -6942 22747 -6922
rect 22835 -962 22905 -942
rect 22835 -6942 22905 -6922
rect 22993 -962 23063 -942
rect 22993 -6942 23063 -6922
rect 23151 -962 23221 -942
rect 23151 -6942 23221 -6922
rect 23309 -962 23379 -942
rect 23309 -6942 23379 -6922
rect 23467 -962 23537 -942
rect 23467 -6942 23537 -6922
rect 23625 -962 23695 -942
rect 23625 -6942 23695 -6922
rect 23783 -962 23853 -942
rect 23783 -6942 23853 -6922
rect 23941 -962 24011 -942
rect 23941 -6942 24011 -6922
rect 24099 -962 24169 -942
rect 24099 -6942 24169 -6922
rect 24257 -962 24327 -942
rect 24257 -6942 24327 -6922
rect 24415 -962 24485 -942
rect 24415 -6942 24485 -6922
rect 24573 -962 24643 -942
rect 24573 -6942 24643 -6922
rect 24731 -962 24801 -942
rect 24731 -6942 24801 -6922
rect 24889 -962 24959 -942
rect 24889 -6942 24959 -6922
rect 25047 -962 25117 -942
rect 25047 -6942 25117 -6922
rect 25205 -962 25275 -942
rect 25205 -6942 25275 -6922
rect 20532 -6990 20552 -6974
rect 25186 -6990 25206 -6974
rect 20532 -7060 20540 -6990
rect 25190 -7060 25206 -6990
rect 20532 -7074 20552 -7060
rect 25186 -7074 25206 -7060
rect 20330 -7170 20400 -7100
rect 25340 -7170 25410 -7100
<< via2 >>
rect 1640 6710 1652 6780
rect 1652 6710 6286 6780
rect 6286 6710 6300 6780
rect 1570 1210 1630 6110
rect 1728 1210 1788 6110
rect 1886 1210 1946 6110
rect 2044 1210 2104 6110
rect 2202 1210 2262 6110
rect 2360 1210 2420 6110
rect 2518 1210 2578 6110
rect 2676 1210 2736 6110
rect 2834 1210 2894 6110
rect 2992 1210 3052 6110
rect 3150 1210 3210 6110
rect 3308 1210 3368 6110
rect 3466 1210 3526 6110
rect 3624 1210 3684 6110
rect 3782 1210 3842 6110
rect 3940 1210 4000 6110
rect 4098 1210 4158 6110
rect 4256 1210 4316 6110
rect 4414 1210 4474 6110
rect 4572 1210 4632 6110
rect 4730 1210 4790 6110
rect 4888 1210 4948 6110
rect 5046 1210 5106 6110
rect 5204 1210 5264 6110
rect 5362 1210 5422 6110
rect 5520 1210 5580 6110
rect 5678 1210 5738 6110
rect 5836 1210 5896 6110
rect 5994 1210 6054 6110
rect 6152 1210 6212 6110
rect 6310 1210 6370 6110
rect 1640 540 1652 610
rect 1652 540 6286 610
rect 6286 540 6290 610
rect 7940 6710 7952 6780
rect 7952 6710 12586 6780
rect 12586 6710 12600 6780
rect 7870 1210 7930 6110
rect 8028 1210 8088 6110
rect 8186 1210 8246 6110
rect 8344 1210 8404 6110
rect 8502 1210 8562 6110
rect 8660 1210 8720 6110
rect 8818 1210 8878 6110
rect 8976 1210 9036 6110
rect 9134 1210 9194 6110
rect 9292 1210 9352 6110
rect 9450 1210 9510 6110
rect 9608 1210 9668 6110
rect 9766 1210 9826 6110
rect 9924 1210 9984 6110
rect 10082 1210 10142 6110
rect 10240 1210 10300 6110
rect 10398 1210 10458 6110
rect 10556 1210 10616 6110
rect 10714 1210 10774 6110
rect 10872 1210 10932 6110
rect 11030 1210 11090 6110
rect 11188 1210 11248 6110
rect 11346 1210 11406 6110
rect 11504 1210 11564 6110
rect 11662 1210 11722 6110
rect 11820 1210 11880 6110
rect 11978 1210 12038 6110
rect 12136 1210 12196 6110
rect 12294 1210 12354 6110
rect 12452 1210 12512 6110
rect 12610 1210 12670 6110
rect 7940 540 7952 610
rect 7952 540 12586 610
rect 12586 540 12590 610
rect 14240 6710 14252 6780
rect 14252 6710 18886 6780
rect 18886 6710 18900 6780
rect 14170 1210 14230 6110
rect 14328 1210 14388 6110
rect 14486 1210 14546 6110
rect 14644 1210 14704 6110
rect 14802 1210 14862 6110
rect 14960 1210 15020 6110
rect 15118 1210 15178 6110
rect 15276 1210 15336 6110
rect 15434 1210 15494 6110
rect 15592 1210 15652 6110
rect 15750 1210 15810 6110
rect 15908 1210 15968 6110
rect 16066 1210 16126 6110
rect 16224 1210 16284 6110
rect 16382 1210 16442 6110
rect 16540 1210 16600 6110
rect 16698 1210 16758 6110
rect 16856 1210 16916 6110
rect 17014 1210 17074 6110
rect 17172 1210 17232 6110
rect 17330 1210 17390 6110
rect 17488 1210 17548 6110
rect 17646 1210 17706 6110
rect 17804 1210 17864 6110
rect 17962 1210 18022 6110
rect 18120 1210 18180 6110
rect 18278 1210 18338 6110
rect 18436 1210 18496 6110
rect 18594 1210 18654 6110
rect 18752 1210 18812 6110
rect 18910 1210 18970 6110
rect 14240 540 14252 610
rect 14252 540 18886 610
rect 18886 540 18890 610
rect 20540 6710 20552 6780
rect 20552 6710 25186 6780
rect 25186 6710 25200 6780
rect 20470 1210 20530 6110
rect 20628 1210 20688 6110
rect 20786 1210 20846 6110
rect 20944 1210 21004 6110
rect 21102 1210 21162 6110
rect 21260 1210 21320 6110
rect 21418 1210 21478 6110
rect 21576 1210 21636 6110
rect 21734 1210 21794 6110
rect 21892 1210 21952 6110
rect 22050 1210 22110 6110
rect 22208 1210 22268 6110
rect 22366 1210 22426 6110
rect 22524 1210 22584 6110
rect 22682 1210 22742 6110
rect 22840 1210 22900 6110
rect 22998 1210 23058 6110
rect 23156 1210 23216 6110
rect 23314 1210 23374 6110
rect 23472 1210 23532 6110
rect 23630 1210 23690 6110
rect 23788 1210 23848 6110
rect 23946 1210 24006 6110
rect 24104 1210 24164 6110
rect 24262 1210 24322 6110
rect 24420 1210 24480 6110
rect 24578 1210 24638 6110
rect 24736 1210 24796 6110
rect 24894 1210 24954 6110
rect 25052 1210 25112 6110
rect 25210 1210 25270 6110
rect 20540 540 20552 610
rect 20552 540 25186 610
rect 25186 540 25190 610
rect 1640 -890 1652 -820
rect 1652 -890 6286 -820
rect 6286 -890 6300 -820
rect 1570 -6390 1630 -1490
rect 1728 -6390 1788 -1490
rect 1886 -6390 1946 -1490
rect 2044 -6390 2104 -1490
rect 2202 -6390 2262 -1490
rect 2360 -6390 2420 -1490
rect 2518 -6390 2578 -1490
rect 2676 -6390 2736 -1490
rect 2834 -6390 2894 -1490
rect 2992 -6390 3052 -1490
rect 3150 -6390 3210 -1490
rect 3308 -6390 3368 -1490
rect 3466 -6390 3526 -1490
rect 3624 -6390 3684 -1490
rect 3782 -6390 3842 -1490
rect 3940 -6390 4000 -1490
rect 4098 -6390 4158 -1490
rect 4256 -6390 4316 -1490
rect 4414 -6390 4474 -1490
rect 4572 -6390 4632 -1490
rect 4730 -6390 4790 -1490
rect 4888 -6390 4948 -1490
rect 5046 -6390 5106 -1490
rect 5204 -6390 5264 -1490
rect 5362 -6390 5422 -1490
rect 5520 -6390 5580 -1490
rect 5678 -6390 5738 -1490
rect 5836 -6390 5896 -1490
rect 5994 -6390 6054 -1490
rect 6152 -6390 6212 -1490
rect 6310 -6390 6370 -1490
rect 1640 -7060 1652 -6990
rect 1652 -7060 6286 -6990
rect 6286 -7060 6290 -6990
rect 7940 -890 7952 -820
rect 7952 -890 12586 -820
rect 12586 -890 12600 -820
rect 7870 -6390 7930 -1490
rect 8028 -6390 8088 -1490
rect 8186 -6390 8246 -1490
rect 8344 -6390 8404 -1490
rect 8502 -6390 8562 -1490
rect 8660 -6390 8720 -1490
rect 8818 -6390 8878 -1490
rect 8976 -6390 9036 -1490
rect 9134 -6390 9194 -1490
rect 9292 -6390 9352 -1490
rect 9450 -6390 9510 -1490
rect 9608 -6390 9668 -1490
rect 9766 -6390 9826 -1490
rect 9924 -6390 9984 -1490
rect 10082 -6390 10142 -1490
rect 10240 -6390 10300 -1490
rect 10398 -6390 10458 -1490
rect 10556 -6390 10616 -1490
rect 10714 -6390 10774 -1490
rect 10872 -6390 10932 -1490
rect 11030 -6390 11090 -1490
rect 11188 -6390 11248 -1490
rect 11346 -6390 11406 -1490
rect 11504 -6390 11564 -1490
rect 11662 -6390 11722 -1490
rect 11820 -6390 11880 -1490
rect 11978 -6390 12038 -1490
rect 12136 -6390 12196 -1490
rect 12294 -6390 12354 -1490
rect 12452 -6390 12512 -1490
rect 12610 -6390 12670 -1490
rect 7940 -7060 7952 -6990
rect 7952 -7060 12586 -6990
rect 12586 -7060 12590 -6990
rect 14240 -890 14252 -820
rect 14252 -890 18886 -820
rect 18886 -890 18900 -820
rect 14170 -6390 14230 -1490
rect 14328 -6390 14388 -1490
rect 14486 -6390 14546 -1490
rect 14644 -6390 14704 -1490
rect 14802 -6390 14862 -1490
rect 14960 -6390 15020 -1490
rect 15118 -6390 15178 -1490
rect 15276 -6390 15336 -1490
rect 15434 -6390 15494 -1490
rect 15592 -6390 15652 -1490
rect 15750 -6390 15810 -1490
rect 15908 -6390 15968 -1490
rect 16066 -6390 16126 -1490
rect 16224 -6390 16284 -1490
rect 16382 -6390 16442 -1490
rect 16540 -6390 16600 -1490
rect 16698 -6390 16758 -1490
rect 16856 -6390 16916 -1490
rect 17014 -6390 17074 -1490
rect 17172 -6390 17232 -1490
rect 17330 -6390 17390 -1490
rect 17488 -6390 17548 -1490
rect 17646 -6390 17706 -1490
rect 17804 -6390 17864 -1490
rect 17962 -6390 18022 -1490
rect 18120 -6390 18180 -1490
rect 18278 -6390 18338 -1490
rect 18436 -6390 18496 -1490
rect 18594 -6390 18654 -1490
rect 18752 -6390 18812 -1490
rect 18910 -6390 18970 -1490
rect 14240 -7060 14252 -6990
rect 14252 -7060 18886 -6990
rect 18886 -7060 18890 -6990
rect 20540 -890 20552 -820
rect 20552 -890 25186 -820
rect 25186 -890 25200 -820
rect 20470 -6390 20530 -1490
rect 20628 -6390 20688 -1490
rect 20786 -6390 20846 -1490
rect 20944 -6390 21004 -1490
rect 21102 -6390 21162 -1490
rect 21260 -6390 21320 -1490
rect 21418 -6390 21478 -1490
rect 21576 -6390 21636 -1490
rect 21734 -6390 21794 -1490
rect 21892 -6390 21952 -1490
rect 22050 -6390 22110 -1490
rect 22208 -6390 22268 -1490
rect 22366 -6390 22426 -1490
rect 22524 -6390 22584 -1490
rect 22682 -6390 22742 -1490
rect 22840 -6390 22900 -1490
rect 22998 -6390 23058 -1490
rect 23156 -6390 23216 -1490
rect 23314 -6390 23374 -1490
rect 23472 -6390 23532 -1490
rect 23630 -6390 23690 -1490
rect 23788 -6390 23848 -1490
rect 23946 -6390 24006 -1490
rect 24104 -6390 24164 -1490
rect 24262 -6390 24322 -1490
rect 24420 -6390 24480 -1490
rect 24578 -6390 24638 -1490
rect 24736 -6390 24796 -1490
rect 24894 -6390 24954 -1490
rect 25052 -6390 25112 -1490
rect 25210 -6390 25270 -1490
rect 20540 -7060 20552 -6990
rect 20552 -7060 25186 -6990
rect 25186 -7060 25190 -6990
<< metal3 >>
rect 1500 6780 6500 6900
rect 1500 6710 1640 6780
rect 6300 6710 6500 6780
rect 1500 6700 6500 6710
rect 7800 6780 12800 6900
rect 7800 6710 7940 6780
rect 12600 6710 12800 6780
rect 7800 6700 12800 6710
rect 14100 6780 19100 6900
rect 14100 6710 14240 6780
rect 18900 6710 19100 6780
rect 14100 6700 19100 6710
rect 20400 6780 25400 6900
rect 20400 6710 20540 6780
rect 25200 6710 25400 6780
rect 20400 6700 25400 6710
rect 1723 6589 1793 6590
rect 2039 6589 2109 6590
rect 2355 6589 2425 6590
rect 2671 6589 2741 6590
rect 2987 6589 3057 6590
rect 3303 6589 3373 6590
rect 3619 6589 3689 6590
rect 3935 6589 4005 6590
rect 4251 6589 4321 6590
rect 4567 6589 4637 6590
rect 4883 6589 4953 6590
rect 5199 6589 5269 6590
rect 5515 6589 5585 6590
rect 5831 6589 5901 6590
rect 6147 6589 6217 6590
rect 8023 6589 8093 6590
rect 8339 6589 8409 6590
rect 8655 6589 8725 6590
rect 8971 6589 9041 6590
rect 9287 6589 9357 6590
rect 9603 6589 9673 6590
rect 9919 6589 9989 6590
rect 10235 6589 10305 6590
rect 10551 6589 10621 6590
rect 10867 6589 10937 6590
rect 11183 6589 11253 6590
rect 11499 6589 11569 6590
rect 11815 6589 11885 6590
rect 12131 6589 12201 6590
rect 12447 6589 12517 6590
rect 14323 6589 14393 6590
rect 14639 6589 14709 6590
rect 14955 6589 15025 6590
rect 15271 6589 15341 6590
rect 15587 6589 15657 6590
rect 15903 6589 15973 6590
rect 16219 6589 16289 6590
rect 16535 6589 16605 6590
rect 16851 6589 16921 6590
rect 17167 6589 17237 6590
rect 17483 6589 17553 6590
rect 17799 6589 17869 6590
rect 18115 6589 18185 6590
rect 18431 6589 18501 6590
rect 18747 6589 18817 6590
rect 20623 6589 20693 6590
rect 20939 6589 21009 6590
rect 21255 6589 21325 6590
rect 21571 6589 21641 6590
rect 21887 6589 21957 6590
rect 22203 6589 22273 6590
rect 22519 6589 22589 6590
rect 22835 6589 22905 6590
rect 23151 6589 23221 6590
rect 23467 6589 23537 6590
rect 23783 6589 23853 6590
rect 24099 6589 24169 6590
rect 24415 6589 24485 6590
rect 24731 6589 24801 6590
rect 25047 6589 25117 6590
rect 1560 6560 6380 6589
rect 1560 6220 1620 6560
rect 5020 6220 6380 6560
rect 1560 6189 6380 6220
rect 7860 6560 12680 6589
rect 7860 6220 7880 6560
rect 9260 6220 12680 6560
rect 7860 6189 12680 6220
rect 14160 6560 18980 6589
rect 14160 6220 14220 6560
rect 17620 6220 18980 6560
rect 14160 6189 18980 6220
rect 20460 6560 25280 6589
rect 20460 6220 20480 6560
rect 21860 6220 25280 6560
rect 20460 6189 25280 6220
rect 1565 6110 1635 6120
rect 1565 1210 1570 6110
rect 1630 1210 1635 6110
rect 1565 1140 1635 1210
rect 1723 6110 1793 6189
rect 1723 1210 1728 6110
rect 1788 1210 1793 6110
rect 1723 1200 1793 1210
rect 1881 6110 1951 6120
rect 1881 1210 1886 6110
rect 1946 1210 1951 6110
rect 1881 1140 1951 1210
rect 2039 6110 2109 6189
rect 2039 1210 2044 6110
rect 2104 1210 2109 6110
rect 2039 1200 2109 1210
rect 2197 6110 2267 6120
rect 2197 1210 2202 6110
rect 2262 1210 2267 6110
rect 2197 1140 2267 1210
rect 2355 6110 2425 6189
rect 2355 1210 2360 6110
rect 2420 1210 2425 6110
rect 2355 1200 2425 1210
rect 2513 6110 2583 6120
rect 2513 1210 2518 6110
rect 2578 1210 2583 6110
rect 2513 1140 2583 1210
rect 2671 6110 2741 6189
rect 2671 1210 2676 6110
rect 2736 1210 2741 6110
rect 2671 1200 2741 1210
rect 2829 6110 2899 6120
rect 2829 1210 2834 6110
rect 2894 1210 2899 6110
rect 2829 1140 2899 1210
rect 2987 6110 3057 6189
rect 2987 1210 2992 6110
rect 3052 1210 3057 6110
rect 2987 1200 3057 1210
rect 3145 6110 3215 6120
rect 3145 1210 3150 6110
rect 3210 1210 3215 6110
rect 3145 1140 3215 1210
rect 3303 6110 3373 6189
rect 3303 1210 3308 6110
rect 3368 1210 3373 6110
rect 3303 1200 3373 1210
rect 3461 6110 3531 6120
rect 3461 1210 3466 6110
rect 3526 1210 3531 6110
rect 3461 1140 3531 1210
rect 3619 6110 3689 6189
rect 3935 6120 4005 6189
rect 3619 1210 3624 6110
rect 3684 1210 3689 6110
rect 3619 1200 3689 1210
rect 3777 6110 3847 6120
rect 3777 1210 3782 6110
rect 3842 1210 3847 6110
rect 3777 1140 3847 1210
rect 3935 6110 4006 6120
rect 3935 1210 3940 6110
rect 4000 1210 4006 6110
rect 3935 1200 4006 1210
rect 4093 6110 4163 6120
rect 4093 1210 4098 6110
rect 4158 1210 4163 6110
rect 4093 1140 4163 1210
rect 4251 6110 4321 6189
rect 4251 1210 4256 6110
rect 4316 1210 4321 6110
rect 4251 1200 4321 1210
rect 4409 6110 4479 6120
rect 4409 1210 4414 6110
rect 4474 1210 4479 6110
rect 4409 1140 4479 1210
rect 4567 6110 4637 6189
rect 4567 1210 4572 6110
rect 4632 1210 4637 6110
rect 4567 1200 4637 1210
rect 4725 6110 4795 6120
rect 4725 1210 4730 6110
rect 4790 1210 4795 6110
rect 4725 1140 4795 1210
rect 4883 6110 4953 6189
rect 4883 1210 4888 6110
rect 4948 1210 4953 6110
rect 4883 1200 4953 1210
rect 5041 6110 5111 6120
rect 5041 1210 5046 6110
rect 5106 1210 5111 6110
rect 5041 1140 5111 1210
rect 5199 6110 5269 6189
rect 5199 1210 5204 6110
rect 5264 1210 5269 6110
rect 5199 1200 5269 1210
rect 5357 6110 5427 6120
rect 5357 1210 5362 6110
rect 5422 1210 5427 6110
rect 5357 1140 5427 1210
rect 5515 6110 5585 6189
rect 5515 1210 5520 6110
rect 5580 1210 5585 6110
rect 5515 1200 5585 1210
rect 5673 6110 5743 6120
rect 5673 1210 5678 6110
rect 5738 1210 5743 6110
rect 5673 1140 5743 1210
rect 5831 6110 5901 6189
rect 5831 1210 5836 6110
rect 5896 1210 5901 6110
rect 5831 1200 5901 1210
rect 5989 6110 6059 6120
rect 5989 1210 5994 6110
rect 6054 1210 6059 6110
rect 5989 1140 6059 1210
rect 6147 6110 6217 6189
rect 6147 1210 6152 6110
rect 6212 1210 6217 6110
rect 6147 1200 6217 1210
rect 6305 6110 6375 6120
rect 6305 1210 6310 6110
rect 6370 1210 6375 6110
rect 6305 1140 6375 1210
rect 7865 6110 7935 6120
rect 7865 1210 7870 6110
rect 7930 1210 7935 6110
rect 7865 1140 7935 1210
rect 8023 6110 8093 6189
rect 8023 1210 8028 6110
rect 8088 1210 8093 6110
rect 8023 1200 8093 1210
rect 8181 6110 8251 6120
rect 8181 1210 8186 6110
rect 8246 1210 8251 6110
rect 8181 1140 8251 1210
rect 8339 6110 8409 6189
rect 8339 1210 8344 6110
rect 8404 1210 8409 6110
rect 8339 1200 8409 1210
rect 8497 6110 8567 6120
rect 8497 1210 8502 6110
rect 8562 1210 8567 6110
rect 8497 1140 8567 1210
rect 8655 6110 8725 6189
rect 8655 1210 8660 6110
rect 8720 1210 8725 6110
rect 8655 1200 8725 1210
rect 8813 6110 8883 6120
rect 8813 1210 8818 6110
rect 8878 1210 8883 6110
rect 8813 1140 8883 1210
rect 8971 6110 9041 6189
rect 8971 1210 8976 6110
rect 9036 1210 9041 6110
rect 8971 1200 9041 1210
rect 9129 6110 9199 6120
rect 9129 1210 9134 6110
rect 9194 1210 9199 6110
rect 9129 1140 9199 1210
rect 9287 6110 9357 6189
rect 9287 1210 9292 6110
rect 9352 1210 9357 6110
rect 9287 1200 9357 1210
rect 9445 6110 9515 6120
rect 9445 1210 9450 6110
rect 9510 1210 9515 6110
rect 9445 1140 9515 1210
rect 9603 6110 9673 6189
rect 9603 1210 9608 6110
rect 9668 1210 9673 6110
rect 9603 1200 9673 1210
rect 9761 6110 9831 6120
rect 9761 1210 9766 6110
rect 9826 1210 9831 6110
rect 9761 1140 9831 1210
rect 9919 6110 9989 6189
rect 10235 6120 10305 6189
rect 9919 1210 9924 6110
rect 9984 1210 9989 6110
rect 9919 1200 9989 1210
rect 10077 6110 10147 6120
rect 10077 1210 10082 6110
rect 10142 1210 10147 6110
rect 10077 1140 10147 1210
rect 10235 6110 10306 6120
rect 10235 1210 10240 6110
rect 10300 1210 10306 6110
rect 10235 1200 10306 1210
rect 10393 6110 10463 6120
rect 10393 1210 10398 6110
rect 10458 1210 10463 6110
rect 10393 1140 10463 1210
rect 10551 6110 10621 6189
rect 10551 1210 10556 6110
rect 10616 1210 10621 6110
rect 10551 1200 10621 1210
rect 10709 6110 10779 6120
rect 10709 1210 10714 6110
rect 10774 1210 10779 6110
rect 10709 1140 10779 1210
rect 10867 6110 10937 6189
rect 10867 1210 10872 6110
rect 10932 1210 10937 6110
rect 10867 1200 10937 1210
rect 11025 6110 11095 6120
rect 11025 1210 11030 6110
rect 11090 1210 11095 6110
rect 11025 1140 11095 1210
rect 11183 6110 11253 6189
rect 11183 1210 11188 6110
rect 11248 1210 11253 6110
rect 11183 1200 11253 1210
rect 11341 6110 11411 6120
rect 11341 1210 11346 6110
rect 11406 1210 11411 6110
rect 11341 1140 11411 1210
rect 11499 6110 11569 6189
rect 11499 1210 11504 6110
rect 11564 1210 11569 6110
rect 11499 1200 11569 1210
rect 11657 6110 11727 6120
rect 11657 1210 11662 6110
rect 11722 1210 11727 6110
rect 11657 1140 11727 1210
rect 11815 6110 11885 6189
rect 11815 1210 11820 6110
rect 11880 1210 11885 6110
rect 11815 1200 11885 1210
rect 11973 6110 12043 6120
rect 11973 1210 11978 6110
rect 12038 1210 12043 6110
rect 11973 1140 12043 1210
rect 12131 6110 12201 6189
rect 12131 1210 12136 6110
rect 12196 1210 12201 6110
rect 12131 1200 12201 1210
rect 12289 6110 12359 6120
rect 12289 1210 12294 6110
rect 12354 1210 12359 6110
rect 12289 1140 12359 1210
rect 12447 6110 12517 6189
rect 12447 1210 12452 6110
rect 12512 1210 12517 6110
rect 12447 1200 12517 1210
rect 12605 6110 12675 6120
rect 12605 1210 12610 6110
rect 12670 1210 12675 6110
rect 12605 1140 12675 1210
rect 14165 6110 14235 6120
rect 14165 1210 14170 6110
rect 14230 1210 14235 6110
rect 14165 1140 14235 1210
rect 14323 6110 14393 6189
rect 14323 1210 14328 6110
rect 14388 1210 14393 6110
rect 14323 1200 14393 1210
rect 14481 6110 14551 6120
rect 14481 1210 14486 6110
rect 14546 1210 14551 6110
rect 14481 1140 14551 1210
rect 14639 6110 14709 6189
rect 14639 1210 14644 6110
rect 14704 1210 14709 6110
rect 14639 1200 14709 1210
rect 14797 6110 14867 6120
rect 14797 1210 14802 6110
rect 14862 1210 14867 6110
rect 14797 1140 14867 1210
rect 14955 6110 15025 6189
rect 14955 1210 14960 6110
rect 15020 1210 15025 6110
rect 14955 1200 15025 1210
rect 15113 6110 15183 6120
rect 15113 1210 15118 6110
rect 15178 1210 15183 6110
rect 15113 1140 15183 1210
rect 15271 6110 15341 6189
rect 15271 1210 15276 6110
rect 15336 1210 15341 6110
rect 15271 1200 15341 1210
rect 15429 6110 15499 6120
rect 15429 1210 15434 6110
rect 15494 1210 15499 6110
rect 15429 1140 15499 1210
rect 15587 6110 15657 6189
rect 15587 1210 15592 6110
rect 15652 1210 15657 6110
rect 15587 1200 15657 1210
rect 15745 6110 15815 6120
rect 15745 1210 15750 6110
rect 15810 1210 15815 6110
rect 15745 1140 15815 1210
rect 15903 6110 15973 6189
rect 15903 1210 15908 6110
rect 15968 1210 15973 6110
rect 15903 1200 15973 1210
rect 16061 6110 16131 6120
rect 16061 1210 16066 6110
rect 16126 1210 16131 6110
rect 16061 1140 16131 1210
rect 16219 6110 16289 6189
rect 16535 6120 16605 6189
rect 16219 1210 16224 6110
rect 16284 1210 16289 6110
rect 16219 1200 16289 1210
rect 16377 6110 16447 6120
rect 16377 1210 16382 6110
rect 16442 1210 16447 6110
rect 16377 1140 16447 1210
rect 16535 6110 16606 6120
rect 16535 1210 16540 6110
rect 16600 1210 16606 6110
rect 16535 1200 16606 1210
rect 16693 6110 16763 6120
rect 16693 1210 16698 6110
rect 16758 1210 16763 6110
rect 16693 1140 16763 1210
rect 16851 6110 16921 6189
rect 16851 1210 16856 6110
rect 16916 1210 16921 6110
rect 16851 1200 16921 1210
rect 17009 6110 17079 6120
rect 17009 1210 17014 6110
rect 17074 1210 17079 6110
rect 17009 1140 17079 1210
rect 17167 6110 17237 6189
rect 17167 1210 17172 6110
rect 17232 1210 17237 6110
rect 17167 1200 17237 1210
rect 17325 6110 17395 6120
rect 17325 1210 17330 6110
rect 17390 1210 17395 6110
rect 17325 1140 17395 1210
rect 17483 6110 17553 6189
rect 17483 1210 17488 6110
rect 17548 1210 17553 6110
rect 17483 1200 17553 1210
rect 17641 6110 17711 6120
rect 17641 1210 17646 6110
rect 17706 1210 17711 6110
rect 17641 1140 17711 1210
rect 17799 6110 17869 6189
rect 17799 1210 17804 6110
rect 17864 1210 17869 6110
rect 17799 1200 17869 1210
rect 17957 6110 18027 6120
rect 17957 1210 17962 6110
rect 18022 1210 18027 6110
rect 17957 1140 18027 1210
rect 18115 6110 18185 6189
rect 18115 1210 18120 6110
rect 18180 1210 18185 6110
rect 18115 1200 18185 1210
rect 18273 6110 18343 6120
rect 18273 1210 18278 6110
rect 18338 1210 18343 6110
rect 18273 1140 18343 1210
rect 18431 6110 18501 6189
rect 18431 1210 18436 6110
rect 18496 1210 18501 6110
rect 18431 1200 18501 1210
rect 18589 6110 18659 6120
rect 18589 1210 18594 6110
rect 18654 1210 18659 6110
rect 18589 1140 18659 1210
rect 18747 6110 18817 6189
rect 18747 1210 18752 6110
rect 18812 1210 18817 6110
rect 18747 1200 18817 1210
rect 18905 6110 18975 6120
rect 18905 1210 18910 6110
rect 18970 1210 18975 6110
rect 18905 1140 18975 1210
rect 20465 6110 20535 6120
rect 20465 1210 20470 6110
rect 20530 1210 20535 6110
rect 20465 1140 20535 1210
rect 20623 6110 20693 6189
rect 20623 1210 20628 6110
rect 20688 1210 20693 6110
rect 20623 1200 20693 1210
rect 20781 6110 20851 6120
rect 20781 1210 20786 6110
rect 20846 1210 20851 6110
rect 20781 1140 20851 1210
rect 20939 6110 21009 6189
rect 20939 1210 20944 6110
rect 21004 1210 21009 6110
rect 20939 1200 21009 1210
rect 21097 6110 21167 6120
rect 21097 1210 21102 6110
rect 21162 1210 21167 6110
rect 21097 1140 21167 1210
rect 21255 6110 21325 6189
rect 21255 1210 21260 6110
rect 21320 1210 21325 6110
rect 21255 1200 21325 1210
rect 21413 6110 21483 6120
rect 21413 1210 21418 6110
rect 21478 1210 21483 6110
rect 21413 1140 21483 1210
rect 21571 6110 21641 6189
rect 21571 1210 21576 6110
rect 21636 1210 21641 6110
rect 21571 1200 21641 1210
rect 21729 6110 21799 6120
rect 21729 1210 21734 6110
rect 21794 1210 21799 6110
rect 21729 1140 21799 1210
rect 21887 6110 21957 6189
rect 21887 1210 21892 6110
rect 21952 1210 21957 6110
rect 21887 1200 21957 1210
rect 22045 6110 22115 6120
rect 22045 1210 22050 6110
rect 22110 1210 22115 6110
rect 22045 1140 22115 1210
rect 22203 6110 22273 6189
rect 22203 1210 22208 6110
rect 22268 1210 22273 6110
rect 22203 1200 22273 1210
rect 22361 6110 22431 6120
rect 22361 1210 22366 6110
rect 22426 1210 22431 6110
rect 22361 1140 22431 1210
rect 22519 6110 22589 6189
rect 22835 6120 22905 6189
rect 22519 1210 22524 6110
rect 22584 1210 22589 6110
rect 22519 1200 22589 1210
rect 22677 6110 22747 6120
rect 22677 1210 22682 6110
rect 22742 1210 22747 6110
rect 22677 1140 22747 1210
rect 22835 6110 22906 6120
rect 22835 1210 22840 6110
rect 22900 1210 22906 6110
rect 22835 1200 22906 1210
rect 22993 6110 23063 6120
rect 22993 1210 22998 6110
rect 23058 1210 23063 6110
rect 22993 1140 23063 1210
rect 23151 6110 23221 6189
rect 23151 1210 23156 6110
rect 23216 1210 23221 6110
rect 23151 1200 23221 1210
rect 23309 6110 23379 6120
rect 23309 1210 23314 6110
rect 23374 1210 23379 6110
rect 23309 1140 23379 1210
rect 23467 6110 23537 6189
rect 23467 1210 23472 6110
rect 23532 1210 23537 6110
rect 23467 1200 23537 1210
rect 23625 6110 23695 6120
rect 23625 1210 23630 6110
rect 23690 1210 23695 6110
rect 23625 1140 23695 1210
rect 23783 6110 23853 6189
rect 23783 1210 23788 6110
rect 23848 1210 23853 6110
rect 23783 1200 23853 1210
rect 23941 6110 24011 6120
rect 23941 1210 23946 6110
rect 24006 1210 24011 6110
rect 23941 1140 24011 1210
rect 24099 6110 24169 6189
rect 24099 1210 24104 6110
rect 24164 1210 24169 6110
rect 24099 1200 24169 1210
rect 24257 6110 24327 6120
rect 24257 1210 24262 6110
rect 24322 1210 24327 6110
rect 24257 1140 24327 1210
rect 24415 6110 24485 6189
rect 24415 1210 24420 6110
rect 24480 1210 24485 6110
rect 24415 1200 24485 1210
rect 24573 6110 24643 6120
rect 24573 1210 24578 6110
rect 24638 1210 24643 6110
rect 24573 1140 24643 1210
rect 24731 6110 24801 6189
rect 24731 1210 24736 6110
rect 24796 1210 24801 6110
rect 24731 1200 24801 1210
rect 24889 6110 24959 6120
rect 24889 1210 24894 6110
rect 24954 1210 24959 6110
rect 24889 1140 24959 1210
rect 25047 6110 25117 6189
rect 25047 1210 25052 6110
rect 25112 1210 25117 6110
rect 25047 1200 25117 1210
rect 25205 6110 25275 6120
rect 25205 1210 25210 6110
rect 25270 1210 25275 6110
rect 25205 1140 25275 1210
rect 1560 1100 6380 1140
rect 1560 780 1700 1100
rect 4900 780 6380 1100
rect 1560 740 6380 780
rect 7860 1100 12680 1140
rect 7860 780 11440 1100
rect 12660 780 12680 1100
rect 7860 740 12680 780
rect 14160 1100 18980 1140
rect 14160 780 14300 1100
rect 17500 780 18980 1100
rect 14160 740 18980 780
rect 20460 1100 25280 1140
rect 20460 780 24040 1100
rect 25260 780 25280 1100
rect 20460 740 25280 780
rect 1500 610 6500 630
rect 1500 540 1640 610
rect 6290 540 6500 610
rect 1500 430 6500 540
rect 7800 610 12800 630
rect 7800 540 7940 610
rect 12590 540 12800 610
rect 3100 400 5000 430
rect 3100 300 3300 400
rect 1400 100 3300 300
rect 4800 300 5000 400
rect 7800 300 12800 540
rect 14100 610 19100 630
rect 14100 540 14240 610
rect 18890 540 19100 610
rect 14100 400 19100 540
rect 14100 300 15900 400
rect 4800 180 7400 300
rect 4800 100 7020 180
rect 1400 20 7020 100
rect 7380 20 7400 180
rect 1400 0 7400 20
rect 7600 180 13700 300
rect 7600 20 13320 180
rect 13680 20 13700 180
rect 7600 0 13700 20
rect 13900 100 15900 300
rect 17400 300 19100 400
rect 20400 610 25400 630
rect 20400 540 20540 610
rect 25190 540 25400 610
rect 20400 300 25400 540
rect 17400 180 20000 300
rect 17400 100 19620 180
rect 13900 20 19620 100
rect 19980 20 20000 180
rect 13900 0 20000 20
rect 20200 0 25400 300
rect 7600 -200 7900 0
rect 9400 -100 12000 0
rect 13900 -100 14100 0
rect 20200 -100 20500 0
rect 22000 -100 24600 0
rect 6500 -400 7900 -200
rect 12800 -300 14100 -100
rect 19100 -300 20500 -100
rect 3100 -500 5000 -400
rect 6500 -500 6800 -400
rect 9400 -500 12000 -400
rect 12800 -500 13100 -300
rect 15700 -500 17600 -400
rect 19100 -500 19400 -300
rect 22000 -500 24600 -400
rect 1400 -800 3300 -500
rect 4800 -800 6800 -500
rect 7000 -520 13100 -500
rect 7000 -680 7020 -520
rect 7380 -680 13100 -520
rect 7000 -800 13100 -680
rect 13300 -520 15900 -500
rect 13300 -680 13320 -520
rect 13680 -680 15900 -520
rect 13300 -800 15900 -680
rect 17400 -800 19400 -500
rect 19600 -520 25400 -500
rect 19600 -680 19620 -520
rect 19980 -680 25400 -520
rect 19600 -800 25400 -680
rect 1500 -820 6500 -800
rect 1500 -890 1640 -820
rect 6300 -890 6500 -820
rect 1500 -900 6500 -890
rect 7800 -820 12800 -800
rect 7800 -890 7940 -820
rect 12600 -890 12800 -820
rect 7800 -900 12800 -890
rect 14100 -820 19100 -800
rect 14100 -890 14240 -820
rect 18900 -890 19100 -820
rect 14100 -900 19100 -890
rect 20400 -820 25400 -800
rect 20400 -890 20540 -820
rect 25200 -890 25400 -820
rect 20400 -900 25400 -890
rect 1723 -1011 1793 -1010
rect 2039 -1011 2109 -1010
rect 2355 -1011 2425 -1010
rect 2671 -1011 2741 -1010
rect 2987 -1011 3057 -1010
rect 3303 -1011 3373 -1010
rect 3619 -1011 3689 -1010
rect 3935 -1011 4005 -1010
rect 4251 -1011 4321 -1010
rect 4567 -1011 4637 -1010
rect 4883 -1011 4953 -1010
rect 5199 -1011 5269 -1010
rect 5515 -1011 5585 -1010
rect 5831 -1011 5901 -1010
rect 6147 -1011 6217 -1010
rect 8023 -1011 8093 -1010
rect 8339 -1011 8409 -1010
rect 8655 -1011 8725 -1010
rect 8971 -1011 9041 -1010
rect 9287 -1011 9357 -1010
rect 9603 -1011 9673 -1010
rect 9919 -1011 9989 -1010
rect 10235 -1011 10305 -1010
rect 10551 -1011 10621 -1010
rect 10867 -1011 10937 -1010
rect 11183 -1011 11253 -1010
rect 11499 -1011 11569 -1010
rect 11815 -1011 11885 -1010
rect 12131 -1011 12201 -1010
rect 12447 -1011 12517 -1010
rect 14323 -1011 14393 -1010
rect 14639 -1011 14709 -1010
rect 14955 -1011 15025 -1010
rect 15271 -1011 15341 -1010
rect 15587 -1011 15657 -1010
rect 15903 -1011 15973 -1010
rect 16219 -1011 16289 -1010
rect 16535 -1011 16605 -1010
rect 16851 -1011 16921 -1010
rect 17167 -1011 17237 -1010
rect 17483 -1011 17553 -1010
rect 17799 -1011 17869 -1010
rect 18115 -1011 18185 -1010
rect 18431 -1011 18501 -1010
rect 18747 -1011 18817 -1010
rect 20623 -1011 20693 -1010
rect 20939 -1011 21009 -1010
rect 21255 -1011 21325 -1010
rect 21571 -1011 21641 -1010
rect 21887 -1011 21957 -1010
rect 22203 -1011 22273 -1010
rect 22519 -1011 22589 -1010
rect 22835 -1011 22905 -1010
rect 23151 -1011 23221 -1010
rect 23467 -1011 23537 -1010
rect 23783 -1011 23853 -1010
rect 24099 -1011 24169 -1010
rect 24415 -1011 24485 -1010
rect 24731 -1011 24801 -1010
rect 25047 -1011 25117 -1010
rect 1560 -1060 6380 -1011
rect 1560 -1360 3260 -1060
rect 4840 -1360 6380 -1060
rect 1560 -1411 6380 -1360
rect 7860 -1040 12680 -1011
rect 7860 -1380 7900 -1040
rect 9260 -1380 12680 -1040
rect 7860 -1411 12680 -1380
rect 14160 -1060 18980 -1011
rect 14160 -1360 15860 -1060
rect 17440 -1360 18980 -1060
rect 14160 -1411 18980 -1360
rect 20460 -1040 25280 -1011
rect 20460 -1380 20500 -1040
rect 21860 -1380 25280 -1040
rect 20460 -1411 25280 -1380
rect 1565 -1490 1635 -1480
rect 1565 -6390 1570 -1490
rect 1630 -6390 1635 -1490
rect 1565 -6460 1635 -6390
rect 1723 -1490 1793 -1411
rect 1723 -6390 1728 -1490
rect 1788 -6390 1793 -1490
rect 1723 -6400 1793 -6390
rect 1881 -1490 1951 -1480
rect 1881 -6390 1886 -1490
rect 1946 -6390 1951 -1490
rect 1881 -6460 1951 -6390
rect 2039 -1490 2109 -1411
rect 2039 -6390 2044 -1490
rect 2104 -6390 2109 -1490
rect 2039 -6400 2109 -6390
rect 2197 -1490 2267 -1480
rect 2197 -6390 2202 -1490
rect 2262 -6390 2267 -1490
rect 2197 -6460 2267 -6390
rect 2355 -1490 2425 -1411
rect 2355 -6390 2360 -1490
rect 2420 -6390 2425 -1490
rect 2355 -6400 2425 -6390
rect 2513 -1490 2583 -1480
rect 2513 -6390 2518 -1490
rect 2578 -6390 2583 -1490
rect 2513 -6460 2583 -6390
rect 2671 -1490 2741 -1411
rect 2671 -6390 2676 -1490
rect 2736 -6390 2741 -1490
rect 2671 -6400 2741 -6390
rect 2829 -1490 2899 -1480
rect 2829 -6390 2834 -1490
rect 2894 -6390 2899 -1490
rect 2829 -6460 2899 -6390
rect 2987 -1490 3057 -1411
rect 2987 -6390 2992 -1490
rect 3052 -6390 3057 -1490
rect 2987 -6400 3057 -6390
rect 3145 -1490 3215 -1480
rect 3145 -6390 3150 -1490
rect 3210 -6390 3215 -1490
rect 3145 -6460 3215 -6390
rect 3303 -1490 3373 -1411
rect 3303 -6390 3308 -1490
rect 3368 -6390 3373 -1490
rect 3303 -6400 3373 -6390
rect 3461 -1490 3531 -1480
rect 3461 -6390 3466 -1490
rect 3526 -6390 3531 -1490
rect 3461 -6460 3531 -6390
rect 3619 -1490 3689 -1411
rect 3935 -1480 4005 -1411
rect 3619 -6390 3624 -1490
rect 3684 -6390 3689 -1490
rect 3619 -6400 3689 -6390
rect 3777 -1490 3847 -1480
rect 3777 -6390 3782 -1490
rect 3842 -6390 3847 -1490
rect 3777 -6460 3847 -6390
rect 3935 -1490 4006 -1480
rect 3935 -6390 3940 -1490
rect 4000 -6390 4006 -1490
rect 3935 -6400 4006 -6390
rect 4093 -1490 4163 -1480
rect 4093 -6390 4098 -1490
rect 4158 -6390 4163 -1490
rect 4093 -6460 4163 -6390
rect 4251 -1490 4321 -1411
rect 4251 -6390 4256 -1490
rect 4316 -6390 4321 -1490
rect 4251 -6400 4321 -6390
rect 4409 -1490 4479 -1480
rect 4409 -6390 4414 -1490
rect 4474 -6390 4479 -1490
rect 4409 -6460 4479 -6390
rect 4567 -1490 4637 -1411
rect 4567 -6390 4572 -1490
rect 4632 -6390 4637 -1490
rect 4567 -6400 4637 -6390
rect 4725 -1490 4795 -1480
rect 4725 -6390 4730 -1490
rect 4790 -6390 4795 -1490
rect 4725 -6460 4795 -6390
rect 4883 -1490 4953 -1411
rect 4883 -6390 4888 -1490
rect 4948 -6390 4953 -1490
rect 4883 -6400 4953 -6390
rect 5041 -1490 5111 -1480
rect 5041 -6390 5046 -1490
rect 5106 -6390 5111 -1490
rect 5041 -6460 5111 -6390
rect 5199 -1490 5269 -1411
rect 5199 -6390 5204 -1490
rect 5264 -6390 5269 -1490
rect 5199 -6400 5269 -6390
rect 5357 -1490 5427 -1480
rect 5357 -6390 5362 -1490
rect 5422 -6390 5427 -1490
rect 5357 -6460 5427 -6390
rect 5515 -1490 5585 -1411
rect 5515 -6390 5520 -1490
rect 5580 -6390 5585 -1490
rect 5515 -6400 5585 -6390
rect 5673 -1490 5743 -1480
rect 5673 -6390 5678 -1490
rect 5738 -6390 5743 -1490
rect 5673 -6460 5743 -6390
rect 5831 -1490 5901 -1411
rect 5831 -6390 5836 -1490
rect 5896 -6390 5901 -1490
rect 5831 -6400 5901 -6390
rect 5989 -1490 6059 -1480
rect 5989 -6390 5994 -1490
rect 6054 -6390 6059 -1490
rect 5989 -6460 6059 -6390
rect 6147 -1490 6217 -1411
rect 6147 -6390 6152 -1490
rect 6212 -6390 6217 -1490
rect 6147 -6400 6217 -6390
rect 6305 -1490 6375 -1480
rect 6305 -6390 6310 -1490
rect 6370 -6390 6375 -1490
rect 6305 -6460 6375 -6390
rect 7865 -1490 7935 -1480
rect 7865 -6390 7870 -1490
rect 7930 -6390 7935 -1490
rect 7865 -6460 7935 -6390
rect 8023 -1490 8093 -1411
rect 8023 -6390 8028 -1490
rect 8088 -6390 8093 -1490
rect 8023 -6400 8093 -6390
rect 8181 -1490 8251 -1480
rect 8181 -6390 8186 -1490
rect 8246 -6390 8251 -1490
rect 8181 -6460 8251 -6390
rect 8339 -1490 8409 -1411
rect 8339 -6390 8344 -1490
rect 8404 -6390 8409 -1490
rect 8339 -6400 8409 -6390
rect 8497 -1490 8567 -1480
rect 8497 -6390 8502 -1490
rect 8562 -6390 8567 -1490
rect 8497 -6460 8567 -6390
rect 8655 -1490 8725 -1411
rect 8655 -6390 8660 -1490
rect 8720 -6390 8725 -1490
rect 8655 -6400 8725 -6390
rect 8813 -1490 8883 -1480
rect 8813 -6390 8818 -1490
rect 8878 -6390 8883 -1490
rect 8813 -6460 8883 -6390
rect 8971 -1490 9041 -1411
rect 8971 -6390 8976 -1490
rect 9036 -6390 9041 -1490
rect 8971 -6400 9041 -6390
rect 9129 -1490 9199 -1480
rect 9129 -6390 9134 -1490
rect 9194 -6390 9199 -1490
rect 9129 -6460 9199 -6390
rect 9287 -1490 9357 -1411
rect 9287 -6390 9292 -1490
rect 9352 -6390 9357 -1490
rect 9287 -6400 9357 -6390
rect 9445 -1490 9515 -1480
rect 9445 -6390 9450 -1490
rect 9510 -6390 9515 -1490
rect 9445 -6460 9515 -6390
rect 9603 -1490 9673 -1411
rect 9603 -6390 9608 -1490
rect 9668 -6390 9673 -1490
rect 9603 -6400 9673 -6390
rect 9761 -1490 9831 -1480
rect 9761 -6390 9766 -1490
rect 9826 -6390 9831 -1490
rect 9761 -6460 9831 -6390
rect 9919 -1490 9989 -1411
rect 10235 -1480 10305 -1411
rect 9919 -6390 9924 -1490
rect 9984 -6390 9989 -1490
rect 9919 -6400 9989 -6390
rect 10077 -1490 10147 -1480
rect 10077 -6390 10082 -1490
rect 10142 -6390 10147 -1490
rect 10077 -6460 10147 -6390
rect 10235 -1490 10306 -1480
rect 10235 -6390 10240 -1490
rect 10300 -6390 10306 -1490
rect 10235 -6400 10306 -6390
rect 10393 -1490 10463 -1480
rect 10393 -6390 10398 -1490
rect 10458 -6390 10463 -1490
rect 10393 -6460 10463 -6390
rect 10551 -1490 10621 -1411
rect 10551 -6390 10556 -1490
rect 10616 -6390 10621 -1490
rect 10551 -6400 10621 -6390
rect 10709 -1490 10779 -1480
rect 10709 -6390 10714 -1490
rect 10774 -6390 10779 -1490
rect 10709 -6460 10779 -6390
rect 10867 -1490 10937 -1411
rect 10867 -6390 10872 -1490
rect 10932 -6390 10937 -1490
rect 10867 -6400 10937 -6390
rect 11025 -1490 11095 -1480
rect 11025 -6390 11030 -1490
rect 11090 -6390 11095 -1490
rect 11025 -6460 11095 -6390
rect 11183 -1490 11253 -1411
rect 11183 -6390 11188 -1490
rect 11248 -6390 11253 -1490
rect 11183 -6400 11253 -6390
rect 11341 -1490 11411 -1480
rect 11341 -6390 11346 -1490
rect 11406 -6390 11411 -1490
rect 11341 -6460 11411 -6390
rect 11499 -1490 11569 -1411
rect 11499 -6390 11504 -1490
rect 11564 -6390 11569 -1490
rect 11499 -6400 11569 -6390
rect 11657 -1490 11727 -1480
rect 11657 -6390 11662 -1490
rect 11722 -6390 11727 -1490
rect 11657 -6460 11727 -6390
rect 11815 -1490 11885 -1411
rect 11815 -6390 11820 -1490
rect 11880 -6390 11885 -1490
rect 11815 -6400 11885 -6390
rect 11973 -1490 12043 -1480
rect 11973 -6390 11978 -1490
rect 12038 -6390 12043 -1490
rect 11973 -6460 12043 -6390
rect 12131 -1490 12201 -1411
rect 12131 -6390 12136 -1490
rect 12196 -6390 12201 -1490
rect 12131 -6400 12201 -6390
rect 12289 -1490 12359 -1480
rect 12289 -6390 12294 -1490
rect 12354 -6390 12359 -1490
rect 12289 -6460 12359 -6390
rect 12447 -1490 12517 -1411
rect 12447 -6390 12452 -1490
rect 12512 -6390 12517 -1490
rect 12447 -6400 12517 -6390
rect 12605 -1490 12675 -1480
rect 12605 -6390 12610 -1490
rect 12670 -6390 12675 -1490
rect 12605 -6460 12675 -6390
rect 14165 -1490 14235 -1480
rect 14165 -6390 14170 -1490
rect 14230 -6390 14235 -1490
rect 14165 -6460 14235 -6390
rect 14323 -1490 14393 -1411
rect 14323 -6390 14328 -1490
rect 14388 -6390 14393 -1490
rect 14323 -6400 14393 -6390
rect 14481 -1490 14551 -1480
rect 14481 -6390 14486 -1490
rect 14546 -6390 14551 -1490
rect 14481 -6460 14551 -6390
rect 14639 -1490 14709 -1411
rect 14639 -6390 14644 -1490
rect 14704 -6390 14709 -1490
rect 14639 -6400 14709 -6390
rect 14797 -1490 14867 -1480
rect 14797 -6390 14802 -1490
rect 14862 -6390 14867 -1490
rect 14797 -6460 14867 -6390
rect 14955 -1490 15025 -1411
rect 14955 -6390 14960 -1490
rect 15020 -6390 15025 -1490
rect 14955 -6400 15025 -6390
rect 15113 -1490 15183 -1480
rect 15113 -6390 15118 -1490
rect 15178 -6390 15183 -1490
rect 15113 -6460 15183 -6390
rect 15271 -1490 15341 -1411
rect 15271 -6390 15276 -1490
rect 15336 -6390 15341 -1490
rect 15271 -6400 15341 -6390
rect 15429 -1490 15499 -1480
rect 15429 -6390 15434 -1490
rect 15494 -6390 15499 -1490
rect 15429 -6460 15499 -6390
rect 15587 -1490 15657 -1411
rect 15587 -6390 15592 -1490
rect 15652 -6390 15657 -1490
rect 15587 -6400 15657 -6390
rect 15745 -1490 15815 -1480
rect 15745 -6390 15750 -1490
rect 15810 -6390 15815 -1490
rect 15745 -6460 15815 -6390
rect 15903 -1490 15973 -1411
rect 15903 -6390 15908 -1490
rect 15968 -6390 15973 -1490
rect 15903 -6400 15973 -6390
rect 16061 -1490 16131 -1480
rect 16061 -6390 16066 -1490
rect 16126 -6390 16131 -1490
rect 16061 -6460 16131 -6390
rect 16219 -1490 16289 -1411
rect 16535 -1480 16605 -1411
rect 16219 -6390 16224 -1490
rect 16284 -6390 16289 -1490
rect 16219 -6400 16289 -6390
rect 16377 -1490 16447 -1480
rect 16377 -6390 16382 -1490
rect 16442 -6390 16447 -1490
rect 16377 -6460 16447 -6390
rect 16535 -1490 16606 -1480
rect 16535 -6390 16540 -1490
rect 16600 -6390 16606 -1490
rect 16535 -6400 16606 -6390
rect 16693 -1490 16763 -1480
rect 16693 -6390 16698 -1490
rect 16758 -6390 16763 -1490
rect 16693 -6460 16763 -6390
rect 16851 -1490 16921 -1411
rect 16851 -6390 16856 -1490
rect 16916 -6390 16921 -1490
rect 16851 -6400 16921 -6390
rect 17009 -1490 17079 -1480
rect 17009 -6390 17014 -1490
rect 17074 -6390 17079 -1490
rect 17009 -6460 17079 -6390
rect 17167 -1490 17237 -1411
rect 17167 -6390 17172 -1490
rect 17232 -6390 17237 -1490
rect 17167 -6400 17237 -6390
rect 17325 -1490 17395 -1480
rect 17325 -6390 17330 -1490
rect 17390 -6390 17395 -1490
rect 17325 -6460 17395 -6390
rect 17483 -1490 17553 -1411
rect 17483 -6390 17488 -1490
rect 17548 -6390 17553 -1490
rect 17483 -6400 17553 -6390
rect 17641 -1490 17711 -1480
rect 17641 -6390 17646 -1490
rect 17706 -6390 17711 -1490
rect 17641 -6460 17711 -6390
rect 17799 -1490 17869 -1411
rect 17799 -6390 17804 -1490
rect 17864 -6390 17869 -1490
rect 17799 -6400 17869 -6390
rect 17957 -1490 18027 -1480
rect 17957 -6390 17962 -1490
rect 18022 -6390 18027 -1490
rect 17957 -6460 18027 -6390
rect 18115 -1490 18185 -1411
rect 18115 -6390 18120 -1490
rect 18180 -6390 18185 -1490
rect 18115 -6400 18185 -6390
rect 18273 -1490 18343 -1480
rect 18273 -6390 18278 -1490
rect 18338 -6390 18343 -1490
rect 18273 -6460 18343 -6390
rect 18431 -1490 18501 -1411
rect 18431 -6390 18436 -1490
rect 18496 -6390 18501 -1490
rect 18431 -6400 18501 -6390
rect 18589 -1490 18659 -1480
rect 18589 -6390 18594 -1490
rect 18654 -6390 18659 -1490
rect 18589 -6460 18659 -6390
rect 18747 -1490 18817 -1411
rect 18747 -6390 18752 -1490
rect 18812 -6390 18817 -1490
rect 18747 -6400 18817 -6390
rect 18905 -1490 18975 -1480
rect 18905 -6390 18910 -1490
rect 18970 -6390 18975 -1490
rect 18905 -6460 18975 -6390
rect 20465 -1490 20535 -1480
rect 20465 -6390 20470 -1490
rect 20530 -6390 20535 -1490
rect 20465 -6460 20535 -6390
rect 20623 -1490 20693 -1411
rect 20623 -6390 20628 -1490
rect 20688 -6390 20693 -1490
rect 20623 -6400 20693 -6390
rect 20781 -1490 20851 -1480
rect 20781 -6390 20786 -1490
rect 20846 -6390 20851 -1490
rect 20781 -6460 20851 -6390
rect 20939 -1490 21009 -1411
rect 20939 -6390 20944 -1490
rect 21004 -6390 21009 -1490
rect 20939 -6400 21009 -6390
rect 21097 -1490 21167 -1480
rect 21097 -6390 21102 -1490
rect 21162 -6390 21167 -1490
rect 21097 -6460 21167 -6390
rect 21255 -1490 21325 -1411
rect 21255 -6390 21260 -1490
rect 21320 -6390 21325 -1490
rect 21255 -6400 21325 -6390
rect 21413 -1490 21483 -1480
rect 21413 -6390 21418 -1490
rect 21478 -6390 21483 -1490
rect 21413 -6460 21483 -6390
rect 21571 -1490 21641 -1411
rect 21571 -6390 21576 -1490
rect 21636 -6390 21641 -1490
rect 21571 -6400 21641 -6390
rect 21729 -1490 21799 -1480
rect 21729 -6390 21734 -1490
rect 21794 -6390 21799 -1490
rect 21729 -6460 21799 -6390
rect 21887 -1490 21957 -1411
rect 21887 -6390 21892 -1490
rect 21952 -6390 21957 -1490
rect 21887 -6400 21957 -6390
rect 22045 -1490 22115 -1480
rect 22045 -6390 22050 -1490
rect 22110 -6390 22115 -1490
rect 22045 -6460 22115 -6390
rect 22203 -1490 22273 -1411
rect 22203 -6390 22208 -1490
rect 22268 -6390 22273 -1490
rect 22203 -6400 22273 -6390
rect 22361 -1490 22431 -1480
rect 22361 -6390 22366 -1490
rect 22426 -6390 22431 -1490
rect 22361 -6460 22431 -6390
rect 22519 -1490 22589 -1411
rect 22835 -1480 22905 -1411
rect 22519 -6390 22524 -1490
rect 22584 -6390 22589 -1490
rect 22519 -6400 22589 -6390
rect 22677 -1490 22747 -1480
rect 22677 -6390 22682 -1490
rect 22742 -6390 22747 -1490
rect 22677 -6460 22747 -6390
rect 22835 -1490 22906 -1480
rect 22835 -6390 22840 -1490
rect 22900 -6390 22906 -1490
rect 22835 -6400 22906 -6390
rect 22993 -1490 23063 -1480
rect 22993 -6390 22998 -1490
rect 23058 -6390 23063 -1490
rect 22993 -6460 23063 -6390
rect 23151 -1490 23221 -1411
rect 23151 -6390 23156 -1490
rect 23216 -6390 23221 -1490
rect 23151 -6400 23221 -6390
rect 23309 -1490 23379 -1480
rect 23309 -6390 23314 -1490
rect 23374 -6390 23379 -1490
rect 23309 -6460 23379 -6390
rect 23467 -1490 23537 -1411
rect 23467 -6390 23472 -1490
rect 23532 -6390 23537 -1490
rect 23467 -6400 23537 -6390
rect 23625 -1490 23695 -1480
rect 23625 -6390 23630 -1490
rect 23690 -6390 23695 -1490
rect 23625 -6460 23695 -6390
rect 23783 -1490 23853 -1411
rect 23783 -6390 23788 -1490
rect 23848 -6390 23853 -1490
rect 23783 -6400 23853 -6390
rect 23941 -1490 24011 -1480
rect 23941 -6390 23946 -1490
rect 24006 -6390 24011 -1490
rect 23941 -6460 24011 -6390
rect 24099 -1490 24169 -1411
rect 24099 -6390 24104 -1490
rect 24164 -6390 24169 -1490
rect 24099 -6400 24169 -6390
rect 24257 -1490 24327 -1480
rect 24257 -6390 24262 -1490
rect 24322 -6390 24327 -1490
rect 24257 -6460 24327 -6390
rect 24415 -1490 24485 -1411
rect 24415 -6390 24420 -1490
rect 24480 -6390 24485 -1490
rect 24415 -6400 24485 -6390
rect 24573 -1490 24643 -1480
rect 24573 -6390 24578 -1490
rect 24638 -6390 24643 -1490
rect 24573 -6460 24643 -6390
rect 24731 -1490 24801 -1411
rect 24731 -6390 24736 -1490
rect 24796 -6390 24801 -1490
rect 24731 -6400 24801 -6390
rect 24889 -1490 24959 -1480
rect 24889 -6390 24894 -1490
rect 24954 -6390 24959 -1490
rect 24889 -6460 24959 -6390
rect 25047 -1490 25117 -1411
rect 25047 -6390 25052 -1490
rect 25112 -6390 25117 -1490
rect 25047 -6400 25117 -6390
rect 25205 -1490 25275 -1480
rect 25205 -6390 25210 -1490
rect 25270 -6390 25275 -1490
rect 25205 -6460 25275 -6390
rect 1560 -6500 6380 -6460
rect 1560 -6820 5140 -6500
rect 6360 -6820 6380 -6500
rect 1560 -6860 6380 -6820
rect 7860 -6480 12680 -6460
rect 7860 -6840 9640 -6480
rect 11060 -6840 12680 -6480
rect 7860 -6860 12680 -6840
rect 14160 -6500 18980 -6460
rect 14160 -6820 17740 -6500
rect 18960 -6820 18980 -6500
rect 14160 -6860 18980 -6820
rect 20460 -6480 25280 -6460
rect 20460 -6840 22240 -6480
rect 23660 -6840 25280 -6480
rect 20460 -6860 25280 -6840
rect 1500 -6990 6500 -6970
rect 1500 -7060 1640 -6990
rect 6290 -7060 6500 -6990
rect 1500 -7170 6500 -7060
rect 7800 -6990 12800 -6970
rect 7800 -7060 7940 -6990
rect 12590 -7060 12800 -6990
rect 7800 -7170 12800 -7060
rect 14100 -6990 19100 -6970
rect 14100 -7060 14240 -6990
rect 18890 -7060 19100 -6990
rect 14100 -7170 19100 -7060
rect 20400 -6990 25400 -6970
rect 20400 -7060 20540 -6990
rect 25190 -7060 25400 -6990
rect 20400 -7170 25400 -7060
<< via3 >>
rect 1620 6220 5020 6560
rect 7880 6220 9260 6560
rect 14220 6220 17620 6560
rect 20480 6220 21860 6560
rect 1700 780 4900 1100
rect 11440 780 12660 1100
rect 14300 780 17500 1100
rect 24040 780 25260 1100
rect 3300 100 4800 400
rect 7020 20 7380 180
rect 13320 20 13680 180
rect 15900 100 17400 400
rect 19620 20 19980 180
rect 3300 -800 4800 -500
rect 7020 -680 7380 -520
rect 13320 -680 13680 -520
rect 15900 -800 17400 -500
rect 19620 -680 19980 -520
rect 3260 -1360 4840 -1060
rect 7900 -1380 9260 -1040
rect 15860 -1360 17440 -1060
rect 20500 -1380 21860 -1040
rect 5140 -6820 6360 -6500
rect 9640 -6840 11060 -6480
rect 17740 -6820 18960 -6500
rect 22240 -6840 23660 -6480
<< metal4 >>
rect 5200 11100 6700 11200
rect 5200 9500 5300 11100
rect 6600 9500 6700 11100
rect 1400 8000 2900 8200
rect 1400 6600 1600 8000
rect 2800 6600 2900 8000
rect 1400 6560 5100 6600
rect 1400 6220 1620 6560
rect 5020 6220 5100 6560
rect 1400 6180 5100 6220
rect 1400 1100 5000 1140
rect 1400 780 1700 1100
rect 4900 780 5000 1100
rect 1400 700 5000 780
rect 1400 -9900 2900 700
rect 3200 400 4900 500
rect 3200 100 3300 400
rect 4800 100 4900 400
rect 3200 0 4900 100
rect 3200 -500 4900 -400
rect 3200 -800 3300 -500
rect 4800 -800 4900 -500
rect 3200 -900 4900 -800
rect 3220 -1060 4880 -1020
rect 3220 -1360 3260 -1060
rect 4840 -1360 4880 -1060
rect 3220 -1400 4880 -1360
rect 3300 -6900 4800 -1400
rect 5200 -6460 6700 9500
rect 7700 11100 9200 11200
rect 7700 9500 7800 11100
rect 9100 9500 9200 11100
rect 7700 6600 9200 9500
rect 17800 11100 19300 11200
rect 17800 9500 17900 11100
rect 19200 9500 19300 11100
rect 9600 8100 11100 8200
rect 7700 6560 9300 6600
rect 7700 6220 7880 6560
rect 9260 6220 9300 6560
rect 7700 6180 9300 6220
rect 9600 6500 9800 8100
rect 11000 6500 11100 8100
rect 7000 180 7400 200
rect 7000 20 7020 180
rect 7380 20 7400 180
rect 7000 -520 7400 20
rect 7000 -680 7020 -520
rect 7380 -680 7400 -520
rect 7000 -700 7400 -680
rect 5100 -6500 6700 -6460
rect 5100 -6820 5140 -6500
rect 6360 -6820 6700 -6500
rect 5100 -6860 6700 -6820
rect 7700 -1040 9300 -1000
rect 7700 -1380 7900 -1040
rect 9260 -1380 9300 -1040
rect 7700 -1420 9300 -1380
rect 3300 -8500 3400 -6900
rect 4700 -8500 4800 -6900
rect 3300 -8600 4800 -8500
rect 1400 -11500 1500 -9900
rect 2800 -11500 2900 -9900
rect 1400 -11600 2900 -11500
rect 7700 -9900 9200 -1420
rect 9600 -6480 11100 6500
rect 14000 8000 15500 8200
rect 14000 6600 14200 8000
rect 15400 6600 15500 8000
rect 14000 6560 17700 6600
rect 14000 6220 14220 6560
rect 17620 6220 17700 6560
rect 14000 6180 17700 6220
rect 14000 6080 15500 6180
rect 11400 1100 13000 1140
rect 11400 780 11440 1100
rect 12660 780 13000 1100
rect 11400 740 13000 780
rect 9600 -6840 9640 -6480
rect 11060 -6840 11100 -6480
rect 9600 -6860 11100 -6840
rect 11500 -6900 13000 740
rect 14000 1100 17600 1140
rect 14000 780 14300 1100
rect 17500 780 17600 1100
rect 14000 700 17600 780
rect 13300 180 13700 200
rect 13300 20 13320 180
rect 13680 20 13700 180
rect 13300 -520 13700 20
rect 13300 -680 13320 -520
rect 13680 -680 13700 -520
rect 13300 -700 13700 -680
rect 11500 -8500 11600 -6900
rect 12900 -8500 13000 -6900
rect 11500 -8600 13000 -8500
rect 7700 -11500 7800 -9900
rect 9100 -11500 9200 -9900
rect 7700 -11600 9200 -11500
rect 14000 -9900 15500 700
rect 15800 400 17500 500
rect 15800 100 15900 400
rect 17400 100 17500 400
rect 15800 0 17500 100
rect 15800 -500 17500 -400
rect 15800 -800 15900 -500
rect 17400 -800 17500 -500
rect 15800 -900 17500 -800
rect 15820 -1060 17480 -1020
rect 15820 -1360 15860 -1060
rect 17440 -1360 17480 -1060
rect 15820 -1400 17480 -1360
rect 15900 -6900 17400 -1400
rect 17800 -6460 19300 9500
rect 20300 11100 21800 11200
rect 20300 9500 20400 11100
rect 21700 9500 21800 11100
rect 20300 8200 21800 9500
rect 20300 6560 21900 8200
rect 20300 6220 20480 6560
rect 21860 6220 21900 6560
rect 20300 6180 21900 6220
rect 22200 8100 23700 8200
rect 22200 6500 22400 8100
rect 23600 6500 23700 8100
rect 20300 6040 21800 6180
rect 19600 180 20000 200
rect 19600 20 19620 180
rect 19980 20 20000 180
rect 19600 -520 20000 20
rect 19600 -680 19620 -520
rect 19980 -680 20000 -520
rect 19600 -700 20000 -680
rect 17700 -6500 19300 -6460
rect 17700 -6820 17740 -6500
rect 18960 -6820 19300 -6500
rect 17700 -6860 19300 -6820
rect 20300 -1040 21900 -1000
rect 20300 -1380 20500 -1040
rect 21860 -1380 21900 -1040
rect 20300 -1420 21900 -1380
rect 15900 -8500 16000 -6900
rect 17300 -8500 17400 -6900
rect 15900 -8600 17400 -8500
rect 14000 -11500 14100 -9900
rect 15400 -11500 15500 -9900
rect 14000 -11600 15500 -11500
rect 20300 -9900 21800 -1420
rect 22200 -6480 23700 6500
rect 24000 1100 25340 1140
rect 24000 780 24040 1100
rect 25260 780 25340 1100
rect 24000 740 25340 780
rect 22200 -6840 22240 -6480
rect 23660 -6840 23700 -6480
rect 22200 -6860 23700 -6840
rect 24100 700 25340 740
rect 24100 -6900 25600 700
rect 24100 -8500 24200 -6900
rect 25500 -8500 25600 -6900
rect 24100 -8600 25600 -8500
rect 20300 -11500 20400 -9900
rect 21700 -11500 21800 -9900
rect 20300 -11600 21800 -11500
<< via4 >>
rect 5300 9500 6600 11100
rect 1600 6600 2800 8000
rect 3300 100 4800 400
rect 3300 -800 4800 -500
rect 7800 9500 9100 11100
rect 17900 9500 19200 11100
rect 9800 6500 11000 8100
rect 3400 -8500 4700 -6900
rect 1500 -11500 2800 -9900
rect 14200 6600 15400 8000
rect 11600 -8500 12900 -6900
rect 7800 -11500 9100 -9900
rect 15900 100 17400 400
rect 15900 -800 17400 -500
rect 20400 9500 21700 11100
rect 22400 6500 23600 8100
rect 16000 -8500 17300 -6900
rect 14100 -11500 15400 -9900
rect 24200 -8500 25500 -6900
rect 20400 -11500 21700 -9900
<< metal5 >>
rect 1400 8200 4200 11400
rect 22800 11200 25600 11400
rect 5200 11100 25600 11200
rect 5200 9500 5300 11100
rect 6600 9500 7800 11100
rect 9100 9500 17900 11100
rect 19200 9500 20400 11100
rect 21700 9500 25600 11100
rect 5200 9400 25600 9500
rect 1400 8100 23700 8200
rect 1400 8000 9800 8100
rect 1400 6600 1600 8000
rect 2800 6600 9800 8000
rect 1400 6500 9800 6600
rect 11000 8000 22400 8100
rect 11000 6600 14200 8000
rect 15400 6600 22400 8000
rect 11000 6500 22400 6600
rect 23600 6500 23700 8100
rect 1400 6400 23700 6500
rect 1300 400 25500 500
rect 1300 100 3300 400
rect 4800 100 15900 400
rect 17400 100 25500 400
rect 1300 0 25500 100
rect 1300 -500 25500 -400
rect 1300 -800 3300 -500
rect 4800 -800 15900 -500
rect 17400 -800 25500 -500
rect 1300 -900 25500 -800
rect 3300 -6900 25600 -6800
rect 3300 -8500 3400 -6900
rect 4700 -8500 11600 -6900
rect 12900 -8500 16000 -6900
rect 17300 -8500 24200 -6900
rect 25500 -8500 25600 -6900
rect 3300 -8600 25600 -8500
rect 1400 -9900 21800 -9800
rect 1400 -11500 1500 -9900
rect 2800 -11500 7800 -9900
rect 9100 -11500 14100 -9900
rect 15400 -11500 20400 -9900
rect 21700 -11500 21800 -9900
rect 1400 -11600 21800 -11500
rect 1400 -11800 4200 -11600
rect 22800 -11800 25600 -8600
<< labels >>
rlabel metal5 1300 0 1400 500 1 GL
rlabel metal5 1300 -900 1400 -400 1 GR
rlabel metal5 1400 -11800 4200 -11600 1 SD2L
rlabel metal5 22800 -11800 25600 -11600 1 SD2R
rlabel metal5 22800 11200 25600 11400 1 SD1R
rlabel metal5 1400 11200 4200 11400 1 SD1L
rlabel metal2 13300 1400 13600 1500 1 SUB
<< end >>
