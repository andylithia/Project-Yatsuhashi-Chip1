* SPICE3 file created from sky130_ef_io__analog_pad.ext - technology: sky130A

.subckt sky130_ef_io__analog_pad P_CORE VSSA VSSD AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO
+ VSWITCH VSSIO VDDA VCCD VCCHIB VSSIO_Q P_PAD
R0 P_CORE P_PAD sky130_fd_pr__res_generic_m5 w=2.5296e+08u l=100000u
C0 VCCHIB P_CORE 13.94fF
C1 AMUXBUS_A VSSA 44.98fF
C2 VSWITCH VSSA 12.85fF
C3 VDDIO_Q VSSIO_Q 11.21fF
C4 VSSA VSSD 21.28fF
C5 VSSIO_Q P_CORE 12.92fF
C6 VSSA P_CORE 15.87fF
C7 VSSIO VSWITCH 10.98fF
C8 AMUXBUS_B VSSA 44.98fF
C9 VDDA VSSA 8.01fF
C10 w_810_9943# VDDIO 3.60fF
C11 VDDIO_Q VDDIO 11.29fF
C12 VDDIO P_CORE 123.70fF
C13 w_810_9943# VSSIO 3.39fF
C14 VDDA VDDIO 18.91fF
C15 VSSIO P_CORE 23.23fF
C16 VSSIO VDDA 10.25fF
C17 VSSIO_Q VSSA 10.26fF
C18 P_CORE sky130_fd_io__simple_pad_and_busses_0/sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1334_20520# 2.02fF
C19 VCCD P_CORE 11.51fF
C20 VCCD VDDA 11.78fF
C21 w_810_9943# P_PAD 20.77fF
C22 AMUXBUS_A P_CORE 6.87fF
C23 VSWITCH P_CORE 8.91fF
C24 P_PAD P_CORE 45.64fF
C25 VCCD VCCHIB 11.43fF
C26 VDDA VSWITCH 4.95fF
C27 VSSD P_CORE 11.54fF
C28 w_810_9943# P_CORE 67.73fF
C29 VDDIO_Q P_CORE 15.90fF
C30 VDDA VSSD 8.46fF
C31 w_810_9943# VDDA 1052.18fF
C32 VSSIO VDDIO 11.30fF
C33 AMUXBUS_B P_CORE 6.73fF
C34 VDDA P_CORE 25.12fF
C35 AMUXBUS_B VDDA 2.17fF
Xsky130_fd_io__simple_pad_and_busses_0/sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0
+ VSSIO VSSA VDDA VSSD VSSIO_Q VSWITCH VCCD VDDIO_Q VDDIO VCCHIB AMUXBUS_B AMUXBUS_A
+ sky130_fd_io__com_bus_hookup
C36 P_PAD VSUBS 26.10fF
C37 P_CORE VSUBS 10.32fF
C38 VCCHIB VSUBS 9.29fF
C39 VCCD VSUBS 4.36fF
C40 VDDA VSUBS 29.93fF
C41 VDDIO VSUBS 13.09fF
C42 VSSIO VSUBS 17.27fF
C43 VSWITCH VSUBS 3.82fF
C44 VSSA VSUBS 7.61fF
C45 VSSD VSUBS 2.81fF
C46 VSSIO_Q VSUBS 2.67fF
C47 VDDIO_Q VSUBS 4.27fF
.ends
