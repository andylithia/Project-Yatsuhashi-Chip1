** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/2stack_1.sch
**.subckt 2stack_1
x1 net8 net1 net10 GND rf_nfet_6xaM02_extracted
L1 net2 net1 2n m=1
V1 VDD GND 1.8
Ldeg5 net3 VDDI 2n m=1
R3 net3 VDD 3 m=1
Ldeg6 net4 GND 2n m=1
R4 net4 GNDI 3 m=1
XC3 net11 GNDI sky130_fd_pr__cap_mim_m3_1 W=40 L=60 MF=8 m=8
C8 GNDI GND 200f m=1
C19 VDD VDDI 200f m=1
R2 net11 VDDI 5 m=1
XC4 net12 GNDI sky130_fd_pr__cap_mim_m3_1 W=40 L=60 MF=8 m=8
R8 net12 VDDI 5 m=1
V2 net6 GND dc 0.9 ac 1 portnum 1 z0 50
V4 net5 GND DC 0.9 AC 0 portnum 2 z0 50
C17 net5 net1 1p m=1
L2 net9 net8 1n m=1
L3 net8 net7 1n m=1
C1 net7 net6 0.4p m=1
x2 vbias vbias GND GND rf_nfet_6xaM02_extracted
I0 VDDI vbias 5m
R1 net9 vbias 1k m=1
C2 vbias GND 2p m=1
V3 net2 GND 0.9
L4 net10 GND 0.3n m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice



.options savecurrents

* .tran 10ps 50ns
.sp dec 1000 1G 10G 1
.control
run
display


.endc


**** end user architecture code
**.ends

* expanding   symbol:  rf_nfet_6xaM02_extracted.sym # of pins=4
** sym_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/rf_nfet_6xaM02_extracted.sym
** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/rf_nfet_6xaM02_extracted.sch
.subckt rf_nfet_6xaM02_extracted  G DS1 DS2 SUB
*.iopin G
*.iopin DS1
*.iopin DS2
*.iopin SUB
**** begin user architecture code


* Extraction of 6xaM02 (12 finger) Transistors
* wt=60um, L=0.15um
.subckt NFET_extract_1 D G S B

 .subckt sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
  X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=1.414e+12p pd=1.066e+07u as=2.828e+12p
+ ps=2.132e+07u w=5.05e+06u l=150000u
  X1 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
  C0 SOURCE DRAIN 3.73fF
  C1 SOURCE SUBSTRATE 2.58fF
 .ends

C0 B G 2.85fF
C1 S D 22.23fF
C2 G D 5.77fF
C3 S G 7.53fF
Xnfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0 D G S B
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xnfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1 D G S B
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xnfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2 D G S B
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xnfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0 D G S B
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xnfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1 D G S B
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xnfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2 D G S B
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
C4 S B 13.70fF
C5 G B 3.35fF

.ends

XM0 DS1 G DS2 SUB NFET_extract_1


**** end user architecture code
.ends

.GLOBAL GND
.GLOBAL GNDI
.end
