magic
tech sky130B
magscale 1 2
timestamp 1659752630
<< metal4 >>
rect -10500 -18786 3200 -18674
rect -10500 -22562 -10388 -18786
rect -6612 -22562 3200 -18786
rect -10500 -22674 3200 -22562
<< via4 >>
rect -10388 -22562 -6612 -18786
<< metal5 >>
tri -36655 1000 -32655 5000 se
rect -32655 1000 -11945 5000
tri -11945 1000 -7945 5000 sw
tri -38502 -847 -36655 1000 se
rect -36655 400 -31598 1000
tri -31598 400 -30998 1000 nw
tri -13602 400 -13002 1000 ne
rect -13002 400 -7945 1000
rect -36655 -448 -32446 400
tri -32446 -448 -31598 400 nw
tri -31598 -448 -30750 400 se
rect -30750 -448 -13850 400
tri -13850 -448 -13002 400 sw
tri -13002 -448 -12154 400 ne
rect -12154 -448 -7945 400
rect -36655 -847 -32845 -448
tri -32845 -847 -32446 -448 nw
tri -31997 -847 -31598 -448 se
rect -31598 -847 -13002 -448
tri -43300 -5645 -38502 -847 se
rect -38502 -1695 -33693 -847
tri -33693 -1695 -32845 -847 nw
tri -32845 -1695 -31997 -847 se
rect -31997 -1296 -13002 -847
tri -13002 -1296 -12154 -448 sw
tri -12154 -1296 -11306 -448 ne
rect -11306 -1296 -7945 -448
rect -31997 -1695 -12154 -1296
rect -38502 -2543 -34541 -1695
tri -34541 -2543 -33693 -1695 nw
tri -33693 -2543 -32845 -1695 se
rect -32845 -2102 -12154 -1695
tri -12154 -2102 -11348 -1296 sw
tri -11306 -2102 -10500 -1296 ne
rect -10500 -2102 -7945 -1296
rect -32845 -2543 -11348 -2102
rect -38502 -2752 -34750 -2543
tri -34750 -2752 -34541 -2543 nw
tri -33902 -2752 -33693 -2543 se
rect -33693 -2752 -11348 -2543
rect -38502 -3600 -35598 -2752
tri -35598 -3600 -34750 -2752 nw
tri -34750 -3600 -33902 -2752 se
rect -33902 -2950 -11348 -2752
tri -11348 -2950 -10500 -2102 sw
tri -10500 -2950 -9652 -2102 ne
rect -9652 -2950 -7945 -2102
rect -33902 -3600 -10500 -2950
rect -38502 -4448 -36446 -3600
tri -36446 -4448 -35598 -3600 nw
tri -35598 -4448 -34750 -3600 se
rect -34750 -4200 -29693 -3600
tri -29693 -4200 -29093 -3600 nw
tri -15507 -4200 -14907 -3600 ne
rect -14907 -3798 -10500 -3600
tri -10500 -3798 -9652 -2950 sw
tri -9652 -3798 -8804 -2950 ne
rect -8804 -3798 -7945 -2950
tri -7945 -3798 -3147 1000 sw
rect -14907 -4200 -9652 -3798
rect -34750 -4448 -30541 -4200
rect -38502 -5296 -37294 -4448
tri -37294 -5296 -36446 -4448 nw
tri -36446 -5296 -35598 -4448 se
rect -35598 -5048 -30541 -4448
tri -30541 -5048 -29693 -4200 nw
tri -29693 -5048 -28845 -4200 se
rect -28845 -5048 -15755 -4200
tri -15755 -5048 -14907 -4200 sw
tri -14907 -5048 -14059 -4200 ne
rect -14059 -4646 -9652 -4200
tri -9652 -4646 -8804 -3798 sw
tri -8804 -4646 -7956 -3798 ne
rect -7956 -4646 -3147 -3798
rect -14059 -5048 -8804 -4646
rect -35598 -5296 -31389 -5048
rect -38502 -5645 -37654 -5296
tri -44159 -6504 -43300 -5645 se
rect -43300 -5656 -37654 -5645
tri -37654 -5656 -37294 -5296 nw
tri -36806 -5656 -36446 -5296 se
rect -36446 -5656 -31389 -5296
rect -43300 -6504 -38502 -5656
tri -38502 -6504 -37654 -5656 nw
tri -37654 -6504 -36806 -5656 se
rect -36806 -5896 -31389 -5656
tri -31389 -5896 -30541 -5048 nw
tri -30541 -5896 -29693 -5048 se
rect -29693 -5896 -14907 -5048
tri -14907 -5896 -14059 -5048 sw
tri -14059 -5896 -13211 -5048 ne
rect -13211 -5494 -8804 -5048
tri -8804 -5494 -7956 -4646 sw
tri -7956 -5494 -7108 -4646 ne
rect -7108 -5494 -3147 -4646
rect -13211 -5896 -7956 -5494
rect -36806 -6504 -31997 -5896
tri -31997 -6504 -31389 -5896 nw
tri -31149 -6504 -30541 -5896 se
rect -30541 -6504 -14059 -5896
tri -14059 -6504 -13451 -5896 sw
tri -13211 -6504 -12603 -5896 ne
rect -12603 -6342 -7956 -5896
tri -7956 -6342 -7108 -5494 sw
tri -7108 -6342 -6260 -5494 ne
rect -6260 -6342 -3147 -5494
rect -12603 -6504 -7108 -6342
tri -47300 -9645 -44159 -6504 se
rect -44159 -7352 -39350 -6504
tri -39350 -7352 -38502 -6504 nw
tri -38502 -7352 -37654 -6504 se
rect -37654 -7352 -32845 -6504
tri -32845 -7352 -31997 -6504 nw
tri -31997 -7352 -31149 -6504 se
rect -31149 -7352 -13451 -6504
tri -13451 -7352 -12603 -6504 sw
tri -12603 -7352 -11755 -6504 ne
rect -11755 -6911 -7108 -6504
tri -7108 -6911 -6539 -6342 sw
tri -6260 -6911 -5691 -6342 ne
rect -5691 -6911 -3147 -6342
rect -11755 -7352 -6539 -6911
rect -44159 -8200 -40198 -7352
tri -40198 -8200 -39350 -7352 nw
tri -39350 -8200 -38502 -7352 se
rect -38502 -8200 -33693 -7352
tri -33693 -8200 -32845 -7352 nw
tri -32845 -8200 -31997 -7352 se
rect -31997 -8200 -12603 -7352
tri -12603 -8200 -11755 -7352 sw
tri -11755 -8200 -10907 -7352 ne
rect -10907 -7759 -6539 -7352
tri -6539 -7759 -5691 -6911 sw
tri -5691 -7759 -4843 -6911 ne
rect -4843 -7759 -3147 -6911
rect -10907 -8200 -5691 -7759
rect -44159 -9048 -41046 -8200
tri -41046 -9048 -40198 -8200 nw
tri -40198 -9048 -39350 -8200 se
rect -39350 -9048 -34541 -8200
tri -34541 -9048 -33693 -8200 nw
tri -33693 -9048 -32845 -8200 se
rect -44159 -9645 -41852 -9048
rect -47300 -9854 -41852 -9645
tri -41852 -9854 -41046 -9048 nw
tri -41004 -9854 -40198 -9048 se
rect -40198 -9854 -35389 -9048
rect -47300 -10702 -42700 -9854
tri -42700 -10702 -41852 -9854 nw
tri -41852 -10702 -41004 -9854 se
rect -41004 -9896 -35389 -9854
tri -35389 -9896 -34541 -9048 nw
tri -34541 -9896 -33693 -9048 se
rect -33693 -9896 -32845 -9048
rect -41004 -10702 -36237 -9896
rect -47300 -18000 -43300 -10702
tri -43300 -11302 -42700 -10702 nw
rect -51300 -22000 -43300 -18000
tri -42700 -11550 -41852 -10702 se
rect -41852 -10744 -36237 -10702
tri -36237 -10744 -35389 -9896 nw
tri -35389 -10744 -34541 -9896 se
rect -34541 -10744 -32845 -9896
rect -41852 -10911 -36404 -10744
tri -36404 -10911 -36237 -10744 nw
tri -35556 -10911 -35389 -10744 se
rect -35389 -10911 -32845 -10744
rect -41852 -11550 -37252 -10911
rect -42700 -11759 -37252 -11550
tri -37252 -11759 -36404 -10911 nw
tri -36404 -11759 -35556 -10911 se
rect -35556 -11759 -32845 -10911
rect -42700 -12607 -38100 -11759
tri -38100 -12607 -37252 -11759 nw
tri -37252 -12607 -36404 -11759 se
rect -36404 -12607 -32845 -11759
rect -42700 -30646 -38700 -12607
tri -38700 -13207 -38100 -12607 nw
tri -38100 -13455 -37252 -12607 se
rect -37252 -13455 -32845 -12607
rect -38100 -13857 -32845 -13455
tri -32845 -13857 -27188 -8200 nw
tri -17412 -13857 -11755 -8200 ne
tri -11755 -8607 -11348 -8200 sw
tri -10907 -8607 -10500 -8200 ne
rect -10500 -8607 -5691 -8200
tri -5691 -8607 -4843 -7759 sw
tri -4843 -8607 -3995 -7759 ne
rect -3995 -8607 -3147 -7759
rect -11755 -9455 -11348 -8607
tri -11348 -9455 -10500 -8607 sw
tri -10500 -9455 -9652 -8607 ne
rect -9652 -9455 -4843 -8607
tri -4843 -9455 -3995 -8607 sw
tri -3995 -9455 -3147 -8607 ne
tri -3147 -9455 2510 -3798 sw
rect -11755 -10303 -10500 -9455
tri -10500 -10303 -9652 -9455 sw
tri -9652 -10303 -8804 -9455 ne
rect -8804 -10303 -3995 -9455
tri -3995 -10303 -3147 -9455 sw
tri -3147 -10303 -2299 -9455 ne
rect -2299 -9645 2510 -9455
tri 2510 -9645 2700 -9455 sw
rect -2299 -10303 2700 -9645
rect -11755 -11151 -9652 -10303
tri -9652 -11151 -8804 -10303 sw
tri -8804 -11151 -7956 -10303 ne
rect -7956 -10702 -3147 -10303
tri -3147 -10702 -2748 -10303 sw
tri -2299 -10702 -1900 -10303 ne
rect -1900 -10702 2700 -10303
rect -7956 -11151 -2748 -10702
rect -11755 -11759 -8804 -11151
tri -8804 -11759 -8196 -11151 sw
tri -7956 -11759 -7348 -11151 ne
rect -7348 -11550 -2748 -11151
tri -2748 -11550 -1900 -10702 sw
tri -1900 -11302 -1300 -10702 ne
rect -7348 -11759 -1900 -11550
rect -11755 -12607 -8196 -11759
tri -8196 -12607 -7348 -11759 sw
tri -7348 -12607 -6500 -11759 ne
rect -6500 -12607 -1900 -11759
rect -11755 -13455 -7348 -12607
tri -7348 -13455 -6500 -12607 sw
tri -6500 -13207 -5900 -12607 ne
rect -11755 -13857 -6500 -13455
rect -38100 -29797 -34100 -13857
tri -34100 -15112 -32845 -13857 nw
tri -11755 -15112 -10500 -13857 ne
rect -10500 -18786 -6500 -13857
rect -10500 -22562 -10388 -18786
rect -6612 -22562 -6500 -18786
rect -10500 -22674 -6500 -22562
tri -38700 -30646 -38100 -30046 sw
tri -38100 -30646 -37251 -29797 ne
rect -37251 -30646 -34100 -29797
rect -42700 -31495 -38100 -30646
tri -38100 -31495 -37251 -30646 sw
tri -37251 -31495 -36402 -30646 ne
rect -36402 -31495 -34100 -30646
rect -42700 -31703 -37251 -31495
tri -42700 -36400 -38003 -31703 ne
rect -38003 -32099 -37251 -31703
tri -37251 -32099 -36647 -31495 sw
tri -36402 -32099 -35798 -31495 ne
rect -35798 -32099 -34100 -31495
rect -38003 -32948 -36647 -32099
tri -36647 -32948 -35798 -32099 sw
tri -35798 -32948 -34949 -32099 ne
rect -34949 -32948 -34100 -32099
rect -38003 -33797 -35798 -32948
tri -35798 -33797 -34949 -32948 sw
tri -34949 -33797 -34100 -32948 ne
tri -34100 -33797 -28443 -28140 sw
tri -8503 -30743 -5900 -28140 se
rect -5900 -29797 -1900 -12607
rect -5900 -30646 -2749 -29797
tri -2749 -30646 -1900 -29797 nw
tri -1900 -30646 -1300 -30046 se
rect -1300 -30646 2700 -10702
rect -5900 -30743 -2846 -30646
tri -2846 -30743 -2749 -30646 nw
tri -1997 -30743 -1900 -30646 se
rect -1900 -30743 2700 -30646
tri -11557 -33797 -8503 -30743 se
rect -8503 -31592 -3695 -30743
tri -3695 -31592 -2846 -30743 nw
tri -2846 -31592 -1997 -30743 se
rect -1997 -31592 2700 -30743
rect -8503 -32099 -4202 -31592
tri -4202 -32099 -3695 -31592 nw
tri -3353 -32099 -2846 -31592 se
rect -2846 -31703 2700 -31592
rect -8503 -32948 -5051 -32099
tri -5051 -32948 -4202 -32099 nw
tri -4202 -32948 -3353 -32099 se
rect -3353 -32948 -2846 -32099
rect -8503 -33797 -5900 -32948
tri -5900 -33797 -5051 -32948 nw
tri -5051 -33797 -4202 -32948 se
rect -4202 -33797 -2846 -32948
rect -38003 -34646 -34949 -33797
tri -34949 -34646 -34100 -33797 sw
tri -34100 -34646 -33251 -33797 ne
rect -33251 -34646 -28443 -33797
rect -38003 -35495 -34100 -34646
tri -34100 -35495 -33251 -34646 sw
tri -33251 -35495 -32402 -34646 ne
rect -32402 -35495 -28443 -34646
rect -38003 -35551 -33251 -35495
tri -33251 -35551 -33195 -35495 sw
tri -32402 -35551 -32346 -35495 ne
rect -32346 -35551 -28443 -35495
rect -38003 -36400 -33195 -35551
tri -33195 -36400 -32346 -35551 sw
tri -32346 -36400 -31497 -35551 ne
rect -31497 -36400 -28443 -35551
tri -28443 -36400 -25840 -33797 sw
tri -14160 -36400 -11557 -33797 se
rect -11557 -34646 -6749 -33797
tri -6749 -34646 -5900 -33797 nw
tri -5900 -34646 -5051 -33797 se
rect -5051 -34646 -2846 -33797
rect -11557 -35495 -7598 -34646
tri -7598 -35495 -6749 -34646 nw
tri -6749 -35495 -5900 -34646 se
rect -5900 -35495 -2846 -34646
rect -11557 -35551 -7654 -35495
tri -7654 -35551 -7598 -35495 nw
tri -6805 -35551 -6749 -35495 se
rect -6749 -35551 -2846 -35495
rect -11557 -36400 -8503 -35551
tri -8503 -36400 -7654 -35551 nw
tri -7654 -36400 -6805 -35551 se
rect -6805 -36400 -2846 -35551
tri -38003 -41000 -33403 -36400 ne
rect -33403 -37249 -32346 -36400
tri -32346 -37249 -31497 -36400 sw
tri -31497 -37249 -30648 -36400 ne
rect -30648 -37249 -9352 -36400
tri -9352 -37249 -8503 -36400 nw
tri -8503 -37249 -7654 -36400 se
rect -7654 -37249 -2846 -36400
tri -2846 -37249 2700 -31703 nw
rect -33403 -38098 -31497 -37249
tri -31497 -38098 -30648 -37249 sw
tri -30648 -38098 -29799 -37249 ne
rect -29799 -38098 -10201 -37249
tri -10201 -38098 -9352 -37249 nw
tri -9352 -38098 -8503 -37249 se
rect -33403 -38702 -30648 -38098
tri -30648 -38702 -30044 -38098 sw
tri -29799 -38702 -29195 -38098 ne
rect -29195 -38702 -10805 -38098
tri -10805 -38702 -10201 -38098 nw
tri -9956 -38702 -9352 -38098 se
rect -9352 -38702 -8503 -38098
rect -33403 -39551 -30044 -38702
tri -30044 -39551 -29195 -38702 sw
tri -29195 -39551 -28346 -38702 ne
rect -28346 -39551 -11654 -38702
tri -11654 -39551 -10805 -38702 nw
tri -10805 -39551 -9956 -38702 se
rect -9956 -39551 -8503 -38702
rect -33403 -40400 -29195 -39551
tri -29195 -40400 -28346 -39551 sw
tri -28346 -40400 -27497 -39551 ne
rect -27497 -40400 -12503 -39551
tri -12503 -40400 -11654 -39551 nw
tri -11654 -40400 -10805 -39551 se
rect -10805 -40400 -8503 -39551
rect -33403 -41000 -28346 -40400
tri -28346 -41000 -27746 -40400 sw
tri -12254 -41000 -11654 -40400 se
rect -11654 -41000 -8503 -40400
tri -33403 -45000 -29403 -41000 ne
rect -29403 -42906 -8503 -41000
tri -8503 -42906 -2846 -37249 nw
rect -29403 -45000 -10597 -42906
tri -10597 -45000 -8503 -42906 nw
<< end >>
