magic
tech sky130B
magscale 1 2
timestamp 1662014484
<< metal1 >>
rect -16000 97980 20000 98000
rect -16000 97910 -15850 97980
rect -15650 97910 -15350 97980
rect -15150 97910 -14850 97980
rect -14650 97910 -14350 97980
rect -14150 97910 -13850 97980
rect -13650 97910 -13350 97980
rect -13150 97910 -12850 97980
rect -12650 97910 -12350 97980
rect -12150 97910 -11850 97980
rect -11650 97910 -11350 97980
rect -11150 97910 -10850 97980
rect -10650 97910 -10350 97980
rect -10150 97910 -9850 97980
rect -9650 97910 -9350 97980
rect -9150 97910 -8850 97980
rect -8650 97910 -8350 97980
rect -8150 97910 -7850 97980
rect -7650 97910 -7350 97980
rect -7150 97910 -6850 97980
rect -6650 97910 -6350 97980
rect -6150 97910 -5850 97980
rect -5650 97910 -5350 97980
rect -5150 97910 -4850 97980
rect -4650 97910 -4350 97980
rect -4150 97910 -3850 97980
rect -3650 97910 -3350 97980
rect -3150 97910 -2850 97980
rect -2650 97910 -2350 97980
rect -2150 97910 -1850 97980
rect -1650 97910 -1350 97980
rect -1150 97910 -850 97980
rect -650 97910 -350 97980
rect -150 97910 150 97980
rect 350 97910 650 97980
rect 850 97910 1150 97980
rect 1350 97910 1650 97980
rect 1850 97910 2150 97980
rect 2350 97910 2650 97980
rect 2850 97910 3150 97980
rect 3350 97910 3650 97980
rect 3850 97910 4150 97980
rect 4350 97910 4650 97980
rect 4850 97910 5150 97980
rect 5350 97910 5650 97980
rect 5850 97910 6150 97980
rect 6350 97910 6650 97980
rect 6850 97910 7150 97980
rect 7350 97910 7650 97980
rect 7850 97910 8150 97980
rect 8350 97910 8650 97980
rect 8850 97910 9150 97980
rect 9350 97910 9650 97980
rect 9850 97910 10150 97980
rect 10350 97910 10650 97980
rect 10850 97910 11150 97980
rect 11350 97910 11650 97980
rect 11850 97910 12150 97980
rect 12350 97910 12650 97980
rect 12850 97910 13150 97980
rect 13350 97910 13650 97980
rect 13850 97910 14150 97980
rect 14350 97910 14650 97980
rect 14850 97910 15150 97980
rect 15350 97910 15650 97980
rect 15850 97910 16150 97980
rect 16350 97910 16650 97980
rect 16850 97910 17150 97980
rect 17350 97910 17650 97980
rect 17850 97910 18150 97980
rect 18350 97910 18650 97980
rect 18850 97910 19150 97980
rect 19350 97910 19650 97980
rect 19850 97910 20000 97980
rect -16000 97900 20000 97910
rect -16000 97880 -15880 97900
rect -15620 97880 -15380 97900
rect -15120 97880 -14880 97900
rect -14620 97880 -14380 97900
rect -14120 97880 -13880 97900
rect -13620 97880 -13380 97900
rect -13120 97880 -12880 97900
rect -12620 97880 -12380 97900
rect -12120 97880 -11880 97900
rect -11620 97880 -11380 97900
rect -11120 97880 -10880 97900
rect -10620 97880 -10380 97900
rect -10120 97880 -9880 97900
rect -9620 97880 -9380 97900
rect -9120 97880 -8880 97900
rect -8620 97880 -8380 97900
rect -8120 97880 -7880 97900
rect -7620 97880 -7380 97900
rect -7120 97880 -6880 97900
rect -6620 97880 -6380 97900
rect -6120 97880 -5880 97900
rect -5620 97880 -5380 97900
rect -5120 97880 -4880 97900
rect -4620 97880 -4380 97900
rect -4120 97880 -3880 97900
rect -3620 97880 -3380 97900
rect -3120 97880 -2880 97900
rect -2620 97880 -2380 97900
rect -2120 97880 -1880 97900
rect -1620 97880 -1380 97900
rect -1120 97880 -880 97900
rect -620 97880 -380 97900
rect -120 97880 120 97900
rect 380 97880 620 97900
rect 880 97880 1120 97900
rect 1380 97880 1620 97900
rect 1880 97880 2120 97900
rect 2380 97880 2620 97900
rect 2880 97880 3120 97900
rect 3380 97880 3620 97900
rect 3880 97880 4120 97900
rect 4380 97880 4620 97900
rect 4880 97880 5120 97900
rect 5380 97880 5620 97900
rect 5880 97880 6120 97900
rect 6380 97880 6620 97900
rect 6880 97880 7120 97900
rect 7380 97880 7620 97900
rect 7880 97880 8120 97900
rect 8380 97880 8620 97900
rect 8880 97880 9120 97900
rect 9380 97880 9620 97900
rect 9880 97880 10120 97900
rect 10380 97880 10620 97900
rect 10880 97880 11120 97900
rect 11380 97880 11620 97900
rect 11880 97880 12120 97900
rect 12380 97880 12620 97900
rect 12880 97880 13120 97900
rect 13380 97880 13620 97900
rect 13880 97880 14120 97900
rect 14380 97880 14620 97900
rect 14880 97880 15120 97900
rect 15380 97880 15620 97900
rect 15880 97880 16120 97900
rect 16380 97880 16620 97900
rect 16880 97880 17120 97900
rect 17380 97880 17620 97900
rect 17880 97880 18120 97900
rect 18380 97880 18620 97900
rect 18880 97880 19120 97900
rect 19380 97880 19620 97900
rect 19880 97880 20000 97900
rect -16000 97850 -15900 97880
rect -16000 97650 -15980 97850
rect -15910 97650 -15900 97850
rect -16000 97620 -15900 97650
rect -15600 97850 -15400 97880
rect -15600 97650 -15590 97850
rect -15520 97650 -15480 97850
rect -15410 97650 -15400 97850
rect -15600 97620 -15400 97650
rect -15100 97850 -14900 97880
rect -15100 97650 -15090 97850
rect -15020 97650 -14980 97850
rect -14910 97650 -14900 97850
rect -15100 97620 -14900 97650
rect -14600 97850 -14400 97880
rect -14600 97650 -14590 97850
rect -14520 97650 -14480 97850
rect -14410 97650 -14400 97850
rect -14600 97620 -14400 97650
rect -14100 97850 -13900 97880
rect -14100 97650 -14090 97850
rect -14020 97650 -13980 97850
rect -13910 97650 -13900 97850
rect -14100 97620 -13900 97650
rect -13600 97850 -13400 97880
rect -13600 97650 -13590 97850
rect -13520 97650 -13480 97850
rect -13410 97650 -13400 97850
rect -13600 97620 -13400 97650
rect -13100 97850 -12900 97880
rect -13100 97650 -13090 97850
rect -13020 97650 -12980 97850
rect -12910 97650 -12900 97850
rect -13100 97620 -12900 97650
rect -12600 97850 -12400 97880
rect -12600 97650 -12590 97850
rect -12520 97650 -12480 97850
rect -12410 97650 -12400 97850
rect -12600 97620 -12400 97650
rect -12100 97850 -11900 97880
rect -12100 97650 -12090 97850
rect -12020 97650 -11980 97850
rect -11910 97650 -11900 97850
rect -12100 97620 -11900 97650
rect -11600 97850 -11400 97880
rect -11600 97650 -11590 97850
rect -11520 97650 -11480 97850
rect -11410 97650 -11400 97850
rect -11600 97620 -11400 97650
rect -11100 97850 -10900 97880
rect -11100 97650 -11090 97850
rect -11020 97650 -10980 97850
rect -10910 97650 -10900 97850
rect -11100 97620 -10900 97650
rect -10600 97850 -10400 97880
rect -10600 97650 -10590 97850
rect -10520 97650 -10480 97850
rect -10410 97650 -10400 97850
rect -10600 97620 -10400 97650
rect -10100 97850 -9900 97880
rect -10100 97650 -10090 97850
rect -10020 97650 -9980 97850
rect -9910 97650 -9900 97850
rect -10100 97620 -9900 97650
rect -9600 97850 -9400 97880
rect -9600 97650 -9590 97850
rect -9520 97650 -9480 97850
rect -9410 97650 -9400 97850
rect -9600 97620 -9400 97650
rect -9100 97850 -8900 97880
rect -9100 97650 -9090 97850
rect -9020 97650 -8980 97850
rect -8910 97650 -8900 97850
rect -9100 97620 -8900 97650
rect -8600 97850 -8400 97880
rect -8600 97650 -8590 97850
rect -8520 97650 -8480 97850
rect -8410 97650 -8400 97850
rect -8600 97620 -8400 97650
rect -8100 97850 -7900 97880
rect -8100 97650 -8090 97850
rect -8020 97650 -7980 97850
rect -7910 97650 -7900 97850
rect -8100 97620 -7900 97650
rect -7600 97850 -7400 97880
rect -7600 97650 -7590 97850
rect -7520 97650 -7480 97850
rect -7410 97650 -7400 97850
rect -7600 97620 -7400 97650
rect -7100 97850 -6900 97880
rect -7100 97650 -7090 97850
rect -7020 97650 -6980 97850
rect -6910 97650 -6900 97850
rect -7100 97620 -6900 97650
rect -6600 97850 -6400 97880
rect -6600 97650 -6590 97850
rect -6520 97650 -6480 97850
rect -6410 97650 -6400 97850
rect -6600 97620 -6400 97650
rect -6100 97850 -5900 97880
rect -6100 97650 -6090 97850
rect -6020 97650 -5980 97850
rect -5910 97650 -5900 97850
rect -6100 97620 -5900 97650
rect -5600 97850 -5400 97880
rect -5600 97650 -5590 97850
rect -5520 97650 -5480 97850
rect -5410 97650 -5400 97850
rect -5600 97620 -5400 97650
rect -5100 97850 -4900 97880
rect -5100 97650 -5090 97850
rect -5020 97650 -4980 97850
rect -4910 97650 -4900 97850
rect -5100 97620 -4900 97650
rect -4600 97850 -4400 97880
rect -4600 97650 -4590 97850
rect -4520 97650 -4480 97850
rect -4410 97650 -4400 97850
rect -4600 97620 -4400 97650
rect -4100 97850 -3900 97880
rect -4100 97650 -4090 97850
rect -4020 97650 -3980 97850
rect -3910 97650 -3900 97850
rect -4100 97620 -3900 97650
rect -3600 97850 -3400 97880
rect -3600 97650 -3590 97850
rect -3520 97650 -3480 97850
rect -3410 97650 -3400 97850
rect -3600 97620 -3400 97650
rect -3100 97850 -2900 97880
rect -3100 97650 -3090 97850
rect -3020 97650 -2980 97850
rect -2910 97650 -2900 97850
rect -3100 97620 -2900 97650
rect -2600 97850 -2400 97880
rect -2600 97650 -2590 97850
rect -2520 97650 -2480 97850
rect -2410 97650 -2400 97850
rect -2600 97620 -2400 97650
rect -2100 97850 -1900 97880
rect -2100 97650 -2090 97850
rect -2020 97650 -1980 97850
rect -1910 97650 -1900 97850
rect -2100 97620 -1900 97650
rect -1600 97850 -1400 97880
rect -1600 97650 -1590 97850
rect -1520 97650 -1480 97850
rect -1410 97650 -1400 97850
rect -1600 97620 -1400 97650
rect -1100 97850 -900 97880
rect -1100 97650 -1090 97850
rect -1020 97650 -980 97850
rect -910 97650 -900 97850
rect -1100 97620 -900 97650
rect -600 97850 -400 97880
rect -600 97650 -590 97850
rect -520 97650 -480 97850
rect -410 97650 -400 97850
rect -600 97620 -400 97650
rect -100 97850 100 97880
rect -100 97650 -90 97850
rect -20 97650 20 97850
rect 90 97650 100 97850
rect -100 97620 100 97650
rect 400 97850 600 97880
rect 400 97650 410 97850
rect 480 97650 520 97850
rect 590 97650 600 97850
rect 400 97620 600 97650
rect 900 97850 1100 97880
rect 900 97650 910 97850
rect 980 97650 1020 97850
rect 1090 97650 1100 97850
rect 900 97620 1100 97650
rect 1400 97850 1600 97880
rect 1400 97650 1410 97850
rect 1480 97650 1520 97850
rect 1590 97650 1600 97850
rect 1400 97620 1600 97650
rect 1900 97850 2100 97880
rect 1900 97650 1910 97850
rect 1980 97650 2020 97850
rect 2090 97650 2100 97850
rect 1900 97620 2100 97650
rect 2400 97850 2600 97880
rect 2400 97650 2410 97850
rect 2480 97650 2520 97850
rect 2590 97650 2600 97850
rect 2400 97620 2600 97650
rect 2900 97850 3100 97880
rect 2900 97650 2910 97850
rect 2980 97650 3020 97850
rect 3090 97650 3100 97850
rect 2900 97620 3100 97650
rect 3400 97850 3600 97880
rect 3400 97650 3410 97850
rect 3480 97650 3520 97850
rect 3590 97650 3600 97850
rect 3400 97620 3600 97650
rect 3900 97850 4100 97880
rect 3900 97650 3910 97850
rect 3980 97650 4020 97850
rect 4090 97650 4100 97850
rect 3900 97620 4100 97650
rect 4400 97850 4600 97880
rect 4400 97650 4410 97850
rect 4480 97650 4520 97850
rect 4590 97650 4600 97850
rect 4400 97620 4600 97650
rect 4900 97850 5100 97880
rect 4900 97650 4910 97850
rect 4980 97650 5020 97850
rect 5090 97650 5100 97850
rect 4900 97620 5100 97650
rect 5400 97850 5600 97880
rect 5400 97650 5410 97850
rect 5480 97650 5520 97850
rect 5590 97650 5600 97850
rect 5400 97620 5600 97650
rect 5900 97850 6100 97880
rect 5900 97650 5910 97850
rect 5980 97650 6020 97850
rect 6090 97650 6100 97850
rect 5900 97620 6100 97650
rect 6400 97850 6600 97880
rect 6400 97650 6410 97850
rect 6480 97650 6520 97850
rect 6590 97650 6600 97850
rect 6400 97620 6600 97650
rect 6900 97850 7100 97880
rect 6900 97650 6910 97850
rect 6980 97650 7020 97850
rect 7090 97650 7100 97850
rect 6900 97620 7100 97650
rect 7400 97850 7600 97880
rect 7400 97650 7410 97850
rect 7480 97650 7520 97850
rect 7590 97650 7600 97850
rect 7400 97620 7600 97650
rect 7900 97850 8100 97880
rect 7900 97650 7910 97850
rect 7980 97650 8020 97850
rect 8090 97650 8100 97850
rect 7900 97620 8100 97650
rect 8400 97850 8600 97880
rect 8400 97650 8410 97850
rect 8480 97650 8520 97850
rect 8590 97650 8600 97850
rect 8400 97620 8600 97650
rect 8900 97850 9100 97880
rect 8900 97650 8910 97850
rect 8980 97650 9020 97850
rect 9090 97650 9100 97850
rect 8900 97620 9100 97650
rect 9400 97850 9600 97880
rect 9400 97650 9410 97850
rect 9480 97650 9520 97850
rect 9590 97650 9600 97850
rect 9400 97620 9600 97650
rect 9900 97850 10100 97880
rect 9900 97650 9910 97850
rect 9980 97650 10020 97850
rect 10090 97650 10100 97850
rect 9900 97620 10100 97650
rect 10400 97850 10600 97880
rect 10400 97650 10410 97850
rect 10480 97650 10520 97850
rect 10590 97650 10600 97850
rect 10400 97620 10600 97650
rect 10900 97850 11100 97880
rect 10900 97650 10910 97850
rect 10980 97650 11020 97850
rect 11090 97650 11100 97850
rect 10900 97620 11100 97650
rect 11400 97850 11600 97880
rect 11400 97650 11410 97850
rect 11480 97650 11520 97850
rect 11590 97650 11600 97850
rect 11400 97620 11600 97650
rect 11900 97850 12100 97880
rect 11900 97650 11910 97850
rect 11980 97650 12020 97850
rect 12090 97650 12100 97850
rect 11900 97620 12100 97650
rect 12400 97850 12600 97880
rect 12400 97650 12410 97850
rect 12480 97650 12520 97850
rect 12590 97650 12600 97850
rect 12400 97620 12600 97650
rect 12900 97850 13100 97880
rect 12900 97650 12910 97850
rect 12980 97650 13020 97850
rect 13090 97650 13100 97850
rect 12900 97620 13100 97650
rect 13400 97850 13600 97880
rect 13400 97650 13410 97850
rect 13480 97650 13520 97850
rect 13590 97650 13600 97850
rect 13400 97620 13600 97650
rect 13900 97850 14100 97880
rect 13900 97650 13910 97850
rect 13980 97650 14020 97850
rect 14090 97650 14100 97850
rect 13900 97620 14100 97650
rect 14400 97850 14600 97880
rect 14400 97650 14410 97850
rect 14480 97650 14520 97850
rect 14590 97650 14600 97850
rect 14400 97620 14600 97650
rect 14900 97850 15100 97880
rect 14900 97650 14910 97850
rect 14980 97650 15020 97850
rect 15090 97650 15100 97850
rect 14900 97620 15100 97650
rect 15400 97850 15600 97880
rect 15400 97650 15410 97850
rect 15480 97650 15520 97850
rect 15590 97650 15600 97850
rect 15400 97620 15600 97650
rect 15900 97850 16100 97880
rect 15900 97650 15910 97850
rect 15980 97650 16020 97850
rect 16090 97650 16100 97850
rect 15900 97620 16100 97650
rect 16400 97850 16600 97880
rect 16400 97650 16410 97850
rect 16480 97650 16520 97850
rect 16590 97650 16600 97850
rect 16400 97620 16600 97650
rect 16900 97850 17100 97880
rect 16900 97650 16910 97850
rect 16980 97650 17020 97850
rect 17090 97650 17100 97850
rect 16900 97620 17100 97650
rect 17400 97850 17600 97880
rect 17400 97650 17410 97850
rect 17480 97650 17520 97850
rect 17590 97650 17600 97850
rect 17400 97620 17600 97650
rect 17900 97850 18100 97880
rect 17900 97650 17910 97850
rect 17980 97650 18020 97850
rect 18090 97650 18100 97850
rect 17900 97620 18100 97650
rect 18400 97850 18600 97880
rect 18400 97650 18410 97850
rect 18480 97650 18520 97850
rect 18590 97650 18600 97850
rect 18400 97620 18600 97650
rect 18900 97850 19100 97880
rect 18900 97650 18910 97850
rect 18980 97650 19020 97850
rect 19090 97650 19100 97850
rect 18900 97620 19100 97650
rect 19400 97850 19600 97880
rect 19400 97650 19410 97850
rect 19480 97650 19520 97850
rect 19590 97650 19600 97850
rect 19400 97620 19600 97650
rect 19900 97850 20000 97880
rect 19900 97650 19910 97850
rect 19980 97650 20000 97850
rect 19900 97620 20000 97650
rect -16000 97600 -15880 97620
rect -15620 97600 -15380 97620
rect -15120 97600 -14880 97620
rect -14620 97600 -14380 97620
rect -14120 97600 -13880 97620
rect -13620 97600 -13380 97620
rect -13120 97600 -12880 97620
rect -12620 97600 -12380 97620
rect -12120 97600 -11880 97620
rect -11620 97600 -11380 97620
rect -11120 97600 -10880 97620
rect -10620 97600 -10380 97620
rect -10120 97600 -9880 97620
rect -9620 97600 -9380 97620
rect -9120 97600 -8880 97620
rect -8620 97600 -8380 97620
rect -8120 97600 -7880 97620
rect -7620 97600 -7380 97620
rect -7120 97600 -6880 97620
rect -6620 97600 -6380 97620
rect -6120 97600 -5880 97620
rect -5620 97600 -5380 97620
rect -5120 97600 -4880 97620
rect -4620 97600 -4380 97620
rect -4120 97600 -3880 97620
rect -3620 97600 -3380 97620
rect -3120 97600 -2880 97620
rect -2620 97600 -2380 97620
rect -2120 97600 -1880 97620
rect -1620 97600 -1380 97620
rect -1120 97600 -880 97620
rect -620 97600 -380 97620
rect -120 97600 120 97620
rect 380 97600 620 97620
rect 880 97600 1120 97620
rect 1380 97600 1620 97620
rect 1880 97600 2120 97620
rect 2380 97600 2620 97620
rect 2880 97600 3120 97620
rect 3380 97600 3620 97620
rect 3880 97600 4120 97620
rect 4380 97600 4620 97620
rect 4880 97600 5120 97620
rect 5380 97600 5620 97620
rect 5880 97600 6120 97620
rect 6380 97600 6620 97620
rect 6880 97600 7120 97620
rect 7380 97600 7620 97620
rect 7880 97600 8120 97620
rect 8380 97600 8620 97620
rect 8880 97600 9120 97620
rect 9380 97600 9620 97620
rect 9880 97600 10120 97620
rect 10380 97600 10620 97620
rect 10880 97600 11120 97620
rect 11380 97600 11620 97620
rect 11880 97600 12120 97620
rect 12380 97600 12620 97620
rect 12880 97600 13120 97620
rect 13380 97600 13620 97620
rect 13880 97600 14120 97620
rect 14380 97600 14620 97620
rect 14880 97600 15120 97620
rect 15380 97600 15620 97620
rect 15880 97600 16120 97620
rect 16380 97600 16620 97620
rect 16880 97600 17120 97620
rect 17380 97600 17620 97620
rect 17880 97600 18120 97620
rect 18380 97600 18620 97620
rect 18880 97600 19120 97620
rect 19380 97600 19620 97620
rect 19880 97600 20000 97620
rect -16000 97590 20000 97600
rect -16000 97520 -15850 97590
rect -15650 97520 -15350 97590
rect -15150 97520 -14850 97590
rect -14650 97520 -14350 97590
rect -14150 97520 -13850 97590
rect -13650 97520 -13350 97590
rect -13150 97520 -12850 97590
rect -12650 97520 -12350 97590
rect -12150 97520 -11850 97590
rect -11650 97520 -11350 97590
rect -11150 97520 -10850 97590
rect -10650 97520 -10350 97590
rect -10150 97520 -9850 97590
rect -9650 97520 -9350 97590
rect -9150 97520 -8850 97590
rect -8650 97520 -8350 97590
rect -8150 97520 -7850 97590
rect -7650 97520 -7350 97590
rect -7150 97520 -6850 97590
rect -6650 97520 -6350 97590
rect -6150 97520 -5850 97590
rect -5650 97520 -5350 97590
rect -5150 97520 -4850 97590
rect -4650 97520 -4350 97590
rect -4150 97520 -3850 97590
rect -3650 97520 -3350 97590
rect -3150 97520 -2850 97590
rect -2650 97520 -2350 97590
rect -2150 97520 -1850 97590
rect -1650 97520 -1350 97590
rect -1150 97520 -850 97590
rect -650 97520 -350 97590
rect -150 97520 150 97590
rect 350 97520 650 97590
rect 850 97520 1150 97590
rect 1350 97520 1650 97590
rect 1850 97520 2150 97590
rect 2350 97520 2650 97590
rect 2850 97520 3150 97590
rect 3350 97520 3650 97590
rect 3850 97520 4150 97590
rect 4350 97520 4650 97590
rect 4850 97520 5150 97590
rect 5350 97520 5650 97590
rect 5850 97520 6150 97590
rect 6350 97520 6650 97590
rect 6850 97520 7150 97590
rect 7350 97520 7650 97590
rect 7850 97520 8150 97590
rect 8350 97520 8650 97590
rect 8850 97520 9150 97590
rect 9350 97520 9650 97590
rect 9850 97520 10150 97590
rect 10350 97520 10650 97590
rect 10850 97520 11150 97590
rect 11350 97520 11650 97590
rect 11850 97520 12150 97590
rect 12350 97520 12650 97590
rect 12850 97520 13150 97590
rect 13350 97520 13650 97590
rect 13850 97520 14150 97590
rect 14350 97520 14650 97590
rect 14850 97520 15150 97590
rect 15350 97520 15650 97590
rect 15850 97520 16150 97590
rect 16350 97520 16650 97590
rect 16850 97520 17150 97590
rect 17350 97520 17650 97590
rect 17850 97520 18150 97590
rect 18350 97520 18650 97590
rect 18850 97520 19150 97590
rect 19350 97520 19650 97590
rect 19850 97520 20000 97590
rect -16000 97480 20000 97520
rect -16000 97410 -15850 97480
rect -15650 97410 -15350 97480
rect -15150 97410 -14850 97480
rect -14650 97410 -14350 97480
rect -14150 97410 -13850 97480
rect -13650 97410 -13350 97480
rect -13150 97410 -12850 97480
rect -12650 97410 -12350 97480
rect -12150 97410 -11850 97480
rect -11650 97410 -11350 97480
rect -11150 97410 -10850 97480
rect -10650 97410 -10350 97480
rect -10150 97410 -9850 97480
rect -9650 97410 -9350 97480
rect -9150 97410 -8850 97480
rect -8650 97410 -8350 97480
rect -8150 97410 -7850 97480
rect -7650 97410 -7350 97480
rect -7150 97410 -6850 97480
rect -6650 97410 -6350 97480
rect -6150 97410 -5850 97480
rect -5650 97410 -5350 97480
rect -5150 97410 -4850 97480
rect -4650 97410 -4350 97480
rect -4150 97410 -3850 97480
rect -3650 97410 -3350 97480
rect -3150 97410 -2850 97480
rect -2650 97410 -2350 97480
rect -2150 97410 -1850 97480
rect -1650 97410 -1350 97480
rect -1150 97410 -850 97480
rect -650 97410 -350 97480
rect -150 97410 150 97480
rect 350 97410 650 97480
rect 850 97410 1150 97480
rect 1350 97410 1650 97480
rect 1850 97410 2150 97480
rect 2350 97410 2650 97480
rect 2850 97410 3150 97480
rect 3350 97410 3650 97480
rect 3850 97410 4150 97480
rect 4350 97410 4650 97480
rect 4850 97410 5150 97480
rect 5350 97410 5650 97480
rect 5850 97410 6150 97480
rect 6350 97410 6650 97480
rect 6850 97410 7150 97480
rect 7350 97410 7650 97480
rect 7850 97410 8150 97480
rect 8350 97410 8650 97480
rect 8850 97410 9150 97480
rect 9350 97410 9650 97480
rect 9850 97410 10150 97480
rect 10350 97410 10650 97480
rect 10850 97410 11150 97480
rect 11350 97410 11650 97480
rect 11850 97410 12150 97480
rect 12350 97410 12650 97480
rect 12850 97410 13150 97480
rect 13350 97410 13650 97480
rect 13850 97410 14150 97480
rect 14350 97410 14650 97480
rect 14850 97410 15150 97480
rect 15350 97410 15650 97480
rect 15850 97410 16150 97480
rect 16350 97410 16650 97480
rect 16850 97410 17150 97480
rect 17350 97410 17650 97480
rect 17850 97410 18150 97480
rect 18350 97410 18650 97480
rect 18850 97410 19150 97480
rect 19350 97410 19650 97480
rect 19850 97410 20000 97480
rect -16000 97400 20000 97410
rect -16000 97380 -15880 97400
rect -15620 97380 -15380 97400
rect -15120 97380 -14880 97400
rect -14620 97380 -14380 97400
rect -14120 97380 -13880 97400
rect -13620 97380 -13380 97400
rect -13120 97380 -12880 97400
rect -12620 97380 -12380 97400
rect -12120 97380 -11880 97400
rect -11620 97380 -11380 97400
rect -11120 97380 -10880 97400
rect -10620 97380 -10380 97400
rect -10120 97380 -9880 97400
rect -9620 97380 -9380 97400
rect -9120 97380 -8880 97400
rect -8620 97380 -8380 97400
rect -8120 97380 -7880 97400
rect -7620 97380 -7380 97400
rect -7120 97380 -6880 97400
rect -6620 97380 -6380 97400
rect -6120 97380 -5880 97400
rect -5620 97380 -5380 97400
rect -5120 97380 -4880 97400
rect -4620 97380 -4380 97400
rect -4120 97380 -3880 97400
rect -3620 97380 -3380 97400
rect -3120 97380 -2880 97400
rect -2620 97380 -2380 97400
rect -2120 97380 -1880 97400
rect -1620 97380 -1380 97400
rect -1120 97380 -880 97400
rect -620 97380 -380 97400
rect -120 97380 120 97400
rect 380 97380 620 97400
rect 880 97380 1120 97400
rect 1380 97380 1620 97400
rect 1880 97380 2120 97400
rect 2380 97380 2620 97400
rect 2880 97380 3120 97400
rect 3380 97380 3620 97400
rect 3880 97380 4120 97400
rect 4380 97380 4620 97400
rect 4880 97380 5120 97400
rect 5380 97380 5620 97400
rect 5880 97380 6120 97400
rect 6380 97380 6620 97400
rect 6880 97380 7120 97400
rect 7380 97380 7620 97400
rect 7880 97380 8120 97400
rect 8380 97380 8620 97400
rect 8880 97380 9120 97400
rect 9380 97380 9620 97400
rect 9880 97380 10120 97400
rect 10380 97380 10620 97400
rect 10880 97380 11120 97400
rect 11380 97380 11620 97400
rect 11880 97380 12120 97400
rect 12380 97380 12620 97400
rect 12880 97380 13120 97400
rect 13380 97380 13620 97400
rect 13880 97380 14120 97400
rect 14380 97380 14620 97400
rect 14880 97380 15120 97400
rect 15380 97380 15620 97400
rect 15880 97380 16120 97400
rect 16380 97380 16620 97400
rect 16880 97380 17120 97400
rect 17380 97380 17620 97400
rect 17880 97380 18120 97400
rect 18380 97380 18620 97400
rect 18880 97380 19120 97400
rect 19380 97380 19620 97400
rect 19880 97380 20000 97400
rect -16000 97350 -15900 97380
rect -16000 97150 -15980 97350
rect -15910 97150 -15900 97350
rect -16000 97120 -15900 97150
rect -15600 97350 -15400 97380
rect -15600 97150 -15590 97350
rect -15520 97150 -15480 97350
rect -15410 97150 -15400 97350
rect -15600 97120 -15400 97150
rect -15100 97350 -14900 97380
rect -15100 97150 -15090 97350
rect -15020 97150 -14980 97350
rect -14910 97150 -14900 97350
rect -15100 97120 -14900 97150
rect -14600 97350 -14400 97380
rect -14600 97150 -14590 97350
rect -14520 97150 -14480 97350
rect -14410 97150 -14400 97350
rect -14600 97120 -14400 97150
rect -14100 97350 -13900 97380
rect -14100 97150 -14090 97350
rect -14020 97150 -13980 97350
rect -13910 97150 -13900 97350
rect -14100 97120 -13900 97150
rect -13600 97350 -13400 97380
rect -13600 97150 -13590 97350
rect -13520 97150 -13480 97350
rect -13410 97150 -13400 97350
rect -13600 97120 -13400 97150
rect -13100 97350 -12900 97380
rect -13100 97150 -13090 97350
rect -13020 97150 -12980 97350
rect -12910 97150 -12900 97350
rect -13100 97120 -12900 97150
rect -12600 97350 -12400 97380
rect -12600 97150 -12590 97350
rect -12520 97150 -12480 97350
rect -12410 97150 -12400 97350
rect -12600 97120 -12400 97150
rect -12100 97350 -11900 97380
rect -12100 97150 -12090 97350
rect -12020 97150 -11980 97350
rect -11910 97150 -11900 97350
rect -12100 97120 -11900 97150
rect -11600 97350 -11400 97380
rect -11600 97150 -11590 97350
rect -11520 97150 -11480 97350
rect -11410 97150 -11400 97350
rect -11600 97120 -11400 97150
rect -11100 97350 -10900 97380
rect -11100 97150 -11090 97350
rect -11020 97150 -10980 97350
rect -10910 97150 -10900 97350
rect -11100 97120 -10900 97150
rect -10600 97350 -10400 97380
rect -10600 97150 -10590 97350
rect -10520 97150 -10480 97350
rect -10410 97150 -10400 97350
rect -10600 97120 -10400 97150
rect -10100 97350 -9900 97380
rect -10100 97150 -10090 97350
rect -10020 97150 -9980 97350
rect -9910 97150 -9900 97350
rect -10100 97120 -9900 97150
rect -9600 97350 -9400 97380
rect -9600 97150 -9590 97350
rect -9520 97150 -9480 97350
rect -9410 97150 -9400 97350
rect -9600 97120 -9400 97150
rect -9100 97350 -8900 97380
rect -9100 97150 -9090 97350
rect -9020 97150 -8980 97350
rect -8910 97150 -8900 97350
rect -9100 97120 -8900 97150
rect -8600 97350 -8400 97380
rect -8600 97150 -8590 97350
rect -8520 97150 -8480 97350
rect -8410 97150 -8400 97350
rect -8600 97120 -8400 97150
rect -8100 97350 -7900 97380
rect -8100 97150 -8090 97350
rect -8020 97150 -7980 97350
rect -7910 97150 -7900 97350
rect -8100 97120 -7900 97150
rect -7600 97350 -7400 97380
rect -7600 97150 -7590 97350
rect -7520 97150 -7480 97350
rect -7410 97150 -7400 97350
rect -7600 97120 -7400 97150
rect -7100 97350 -6900 97380
rect -7100 97150 -7090 97350
rect -7020 97150 -6980 97350
rect -6910 97150 -6900 97350
rect -7100 97120 -6900 97150
rect -6600 97350 -6400 97380
rect -6600 97150 -6590 97350
rect -6520 97150 -6480 97350
rect -6410 97150 -6400 97350
rect -6600 97120 -6400 97150
rect -6100 97350 -5900 97380
rect -6100 97150 -6090 97350
rect -6020 97150 -5980 97350
rect -5910 97150 -5900 97350
rect -6100 97120 -5900 97150
rect -5600 97350 -5400 97380
rect -5600 97150 -5590 97350
rect -5520 97150 -5480 97350
rect -5410 97150 -5400 97350
rect -5600 97120 -5400 97150
rect -5100 97350 -4900 97380
rect -5100 97150 -5090 97350
rect -5020 97150 -4980 97350
rect -4910 97150 -4900 97350
rect -5100 97120 -4900 97150
rect -4600 97350 -4400 97380
rect -4600 97150 -4590 97350
rect -4520 97150 -4480 97350
rect -4410 97150 -4400 97350
rect -4600 97120 -4400 97150
rect -4100 97350 -3900 97380
rect -4100 97150 -4090 97350
rect -4020 97150 -3980 97350
rect -3910 97150 -3900 97350
rect -4100 97120 -3900 97150
rect -3600 97350 -3400 97380
rect -3600 97150 -3590 97350
rect -3520 97150 -3480 97350
rect -3410 97150 -3400 97350
rect -3600 97120 -3400 97150
rect -3100 97350 -2900 97380
rect -3100 97150 -3090 97350
rect -3020 97150 -2980 97350
rect -2910 97150 -2900 97350
rect -3100 97120 -2900 97150
rect -2600 97350 -2400 97380
rect -2600 97150 -2590 97350
rect -2520 97150 -2480 97350
rect -2410 97150 -2400 97350
rect -2600 97120 -2400 97150
rect -2100 97350 -1900 97380
rect -2100 97150 -2090 97350
rect -2020 97150 -1980 97350
rect -1910 97150 -1900 97350
rect -2100 97120 -1900 97150
rect -1600 97350 -1400 97380
rect -1600 97150 -1590 97350
rect -1520 97150 -1480 97350
rect -1410 97150 -1400 97350
rect -1600 97120 -1400 97150
rect -1100 97350 -900 97380
rect -1100 97150 -1090 97350
rect -1020 97150 -980 97350
rect -910 97150 -900 97350
rect -1100 97120 -900 97150
rect -600 97350 -400 97380
rect -600 97150 -590 97350
rect -520 97150 -480 97350
rect -410 97150 -400 97350
rect -600 97120 -400 97150
rect -100 97350 100 97380
rect -100 97150 -90 97350
rect -20 97150 20 97350
rect 90 97150 100 97350
rect -100 97120 100 97150
rect 400 97350 600 97380
rect 400 97150 410 97350
rect 480 97150 520 97350
rect 590 97150 600 97350
rect 400 97120 600 97150
rect 900 97350 1100 97380
rect 900 97150 910 97350
rect 980 97150 1020 97350
rect 1090 97150 1100 97350
rect 900 97120 1100 97150
rect 1400 97350 1600 97380
rect 1400 97150 1410 97350
rect 1480 97150 1520 97350
rect 1590 97150 1600 97350
rect 1400 97120 1600 97150
rect 1900 97350 2100 97380
rect 1900 97150 1910 97350
rect 1980 97150 2020 97350
rect 2090 97150 2100 97350
rect 1900 97120 2100 97150
rect 2400 97350 2600 97380
rect 2400 97150 2410 97350
rect 2480 97150 2520 97350
rect 2590 97150 2600 97350
rect 2400 97120 2600 97150
rect 2900 97350 3100 97380
rect 2900 97150 2910 97350
rect 2980 97150 3020 97350
rect 3090 97150 3100 97350
rect 2900 97120 3100 97150
rect 3400 97350 3600 97380
rect 3400 97150 3410 97350
rect 3480 97150 3520 97350
rect 3590 97150 3600 97350
rect 3400 97120 3600 97150
rect 3900 97350 4100 97380
rect 3900 97150 3910 97350
rect 3980 97150 4020 97350
rect 4090 97150 4100 97350
rect 3900 97120 4100 97150
rect 4400 97350 4600 97380
rect 4400 97150 4410 97350
rect 4480 97150 4520 97350
rect 4590 97150 4600 97350
rect 4400 97120 4600 97150
rect 4900 97350 5100 97380
rect 4900 97150 4910 97350
rect 4980 97150 5020 97350
rect 5090 97150 5100 97350
rect 4900 97120 5100 97150
rect 5400 97350 5600 97380
rect 5400 97150 5410 97350
rect 5480 97150 5520 97350
rect 5590 97150 5600 97350
rect 5400 97120 5600 97150
rect 5900 97350 6100 97380
rect 5900 97150 5910 97350
rect 5980 97150 6020 97350
rect 6090 97150 6100 97350
rect 5900 97120 6100 97150
rect 6400 97350 6600 97380
rect 6400 97150 6410 97350
rect 6480 97150 6520 97350
rect 6590 97150 6600 97350
rect 6400 97120 6600 97150
rect 6900 97350 7100 97380
rect 6900 97150 6910 97350
rect 6980 97150 7020 97350
rect 7090 97150 7100 97350
rect 6900 97120 7100 97150
rect 7400 97350 7600 97380
rect 7400 97150 7410 97350
rect 7480 97150 7520 97350
rect 7590 97150 7600 97350
rect 7400 97120 7600 97150
rect 7900 97350 8100 97380
rect 7900 97150 7910 97350
rect 7980 97150 8020 97350
rect 8090 97150 8100 97350
rect 7900 97120 8100 97150
rect 8400 97350 8600 97380
rect 8400 97150 8410 97350
rect 8480 97150 8520 97350
rect 8590 97150 8600 97350
rect 8400 97120 8600 97150
rect 8900 97350 9100 97380
rect 8900 97150 8910 97350
rect 8980 97150 9020 97350
rect 9090 97150 9100 97350
rect 8900 97120 9100 97150
rect 9400 97350 9600 97380
rect 9400 97150 9410 97350
rect 9480 97150 9520 97350
rect 9590 97150 9600 97350
rect 9400 97120 9600 97150
rect 9900 97350 10100 97380
rect 9900 97150 9910 97350
rect 9980 97150 10020 97350
rect 10090 97150 10100 97350
rect 9900 97120 10100 97150
rect 10400 97350 10600 97380
rect 10400 97150 10410 97350
rect 10480 97150 10520 97350
rect 10590 97150 10600 97350
rect 10400 97120 10600 97150
rect 10900 97350 11100 97380
rect 10900 97150 10910 97350
rect 10980 97150 11020 97350
rect 11090 97150 11100 97350
rect 10900 97120 11100 97150
rect 11400 97350 11600 97380
rect 11400 97150 11410 97350
rect 11480 97150 11520 97350
rect 11590 97150 11600 97350
rect 11400 97120 11600 97150
rect 11900 97350 12100 97380
rect 11900 97150 11910 97350
rect 11980 97150 12020 97350
rect 12090 97150 12100 97350
rect 11900 97120 12100 97150
rect 12400 97350 12600 97380
rect 12400 97150 12410 97350
rect 12480 97150 12520 97350
rect 12590 97150 12600 97350
rect 12400 97120 12600 97150
rect 12900 97350 13100 97380
rect 12900 97150 12910 97350
rect 12980 97150 13020 97350
rect 13090 97150 13100 97350
rect 12900 97120 13100 97150
rect 13400 97350 13600 97380
rect 13400 97150 13410 97350
rect 13480 97150 13520 97350
rect 13590 97150 13600 97350
rect 13400 97120 13600 97150
rect 13900 97350 14100 97380
rect 13900 97150 13910 97350
rect 13980 97150 14020 97350
rect 14090 97150 14100 97350
rect 13900 97120 14100 97150
rect 14400 97350 14600 97380
rect 14400 97150 14410 97350
rect 14480 97150 14520 97350
rect 14590 97150 14600 97350
rect 14400 97120 14600 97150
rect 14900 97350 15100 97380
rect 14900 97150 14910 97350
rect 14980 97150 15020 97350
rect 15090 97150 15100 97350
rect 14900 97120 15100 97150
rect 15400 97350 15600 97380
rect 15400 97150 15410 97350
rect 15480 97150 15520 97350
rect 15590 97150 15600 97350
rect 15400 97120 15600 97150
rect 15900 97350 16100 97380
rect 15900 97150 15910 97350
rect 15980 97150 16020 97350
rect 16090 97150 16100 97350
rect 15900 97120 16100 97150
rect 16400 97350 16600 97380
rect 16400 97150 16410 97350
rect 16480 97150 16520 97350
rect 16590 97150 16600 97350
rect 16400 97120 16600 97150
rect 16900 97350 17100 97380
rect 16900 97150 16910 97350
rect 16980 97150 17020 97350
rect 17090 97150 17100 97350
rect 16900 97120 17100 97150
rect 17400 97350 17600 97380
rect 17400 97150 17410 97350
rect 17480 97150 17520 97350
rect 17590 97150 17600 97350
rect 17400 97120 17600 97150
rect 17900 97350 18100 97380
rect 17900 97150 17910 97350
rect 17980 97150 18020 97350
rect 18090 97150 18100 97350
rect 17900 97120 18100 97150
rect 18400 97350 18600 97380
rect 18400 97150 18410 97350
rect 18480 97150 18520 97350
rect 18590 97150 18600 97350
rect 18400 97120 18600 97150
rect 18900 97350 19100 97380
rect 18900 97150 18910 97350
rect 18980 97150 19020 97350
rect 19090 97150 19100 97350
rect 18900 97120 19100 97150
rect 19400 97350 19600 97380
rect 19400 97150 19410 97350
rect 19480 97150 19520 97350
rect 19590 97150 19600 97350
rect 19400 97120 19600 97150
rect 19900 97350 20000 97380
rect 19900 97150 19910 97350
rect 19980 97150 20000 97350
rect 19900 97120 20000 97150
rect -16000 97100 -15880 97120
rect -15620 97100 -15380 97120
rect -15120 97100 -14880 97120
rect -14620 97100 -14380 97120
rect -14120 97100 -13880 97120
rect -13620 97100 -13380 97120
rect -13120 97100 -12880 97120
rect -12620 97100 -12380 97120
rect -12120 97100 -11880 97120
rect -11620 97100 -11380 97120
rect -11120 97100 -10880 97120
rect -10620 97100 -10380 97120
rect -10120 97100 -9880 97120
rect -9620 97100 -9380 97120
rect -9120 97100 -8880 97120
rect -8620 97100 -8380 97120
rect -8120 97100 -7880 97120
rect -7620 97100 -7380 97120
rect -7120 97100 -6880 97120
rect -6620 97100 -6380 97120
rect -6120 97100 -5880 97120
rect -5620 97100 -5380 97120
rect -5120 97100 -4880 97120
rect -4620 97100 -4380 97120
rect -4120 97100 -3880 97120
rect -3620 97100 -3380 97120
rect -3120 97100 -2880 97120
rect -2620 97100 -2380 97120
rect -2120 97100 -1880 97120
rect -1620 97100 -1380 97120
rect -1120 97100 -880 97120
rect -620 97100 -380 97120
rect -120 97100 120 97120
rect 380 97100 620 97120
rect 880 97100 1120 97120
rect 1380 97100 1620 97120
rect 1880 97100 2120 97120
rect 2380 97100 2620 97120
rect 2880 97100 3120 97120
rect 3380 97100 3620 97120
rect 3880 97100 4120 97120
rect 4380 97100 4620 97120
rect 4880 97100 5120 97120
rect 5380 97100 5620 97120
rect 5880 97100 6120 97120
rect 6380 97100 6620 97120
rect 6880 97100 7120 97120
rect 7380 97100 7620 97120
rect 7880 97100 8120 97120
rect 8380 97100 8620 97120
rect 8880 97100 9120 97120
rect 9380 97100 9620 97120
rect 9880 97100 10120 97120
rect 10380 97100 10620 97120
rect 10880 97100 11120 97120
rect 11380 97100 11620 97120
rect 11880 97100 12120 97120
rect 12380 97100 12620 97120
rect 12880 97100 13120 97120
rect 13380 97100 13620 97120
rect 13880 97100 14120 97120
rect 14380 97100 14620 97120
rect 14880 97100 15120 97120
rect 15380 97100 15620 97120
rect 15880 97100 16120 97120
rect 16380 97100 16620 97120
rect 16880 97100 17120 97120
rect 17380 97100 17620 97120
rect 17880 97100 18120 97120
rect 18380 97100 18620 97120
rect 18880 97100 19120 97120
rect 19380 97100 19620 97120
rect 19880 97100 20000 97120
rect -16000 97090 20000 97100
rect -16000 97020 -15850 97090
rect -15650 97020 -15350 97090
rect -15150 97020 -14850 97090
rect -14650 97020 -14350 97090
rect -14150 97020 -13850 97090
rect -13650 97020 -13350 97090
rect -13150 97020 -12850 97090
rect -12650 97020 -12350 97090
rect -12150 97020 -11850 97090
rect -11650 97020 -11350 97090
rect -11150 97020 -10850 97090
rect -10650 97020 -10350 97090
rect -10150 97020 -9850 97090
rect -9650 97020 -9350 97090
rect -9150 97020 -8850 97090
rect -8650 97020 -8350 97090
rect -8150 97020 -7850 97090
rect -7650 97020 -7350 97090
rect -7150 97020 -6850 97090
rect -6650 97020 -6350 97090
rect -6150 97020 -5850 97090
rect -5650 97020 -5350 97090
rect -5150 97020 -4850 97090
rect -4650 97020 -4350 97090
rect -4150 97020 -3850 97090
rect -3650 97020 -3350 97090
rect -3150 97020 -2850 97090
rect -2650 97020 -2350 97090
rect -2150 97020 -1850 97090
rect -1650 97020 -1350 97090
rect -1150 97020 -850 97090
rect -650 97020 -350 97090
rect -150 97020 150 97090
rect 350 97020 650 97090
rect 850 97020 1150 97090
rect 1350 97020 1650 97090
rect 1850 97020 2150 97090
rect 2350 97020 2650 97090
rect 2850 97020 3150 97090
rect 3350 97020 3650 97090
rect 3850 97020 4150 97090
rect 4350 97020 4650 97090
rect 4850 97020 5150 97090
rect 5350 97020 5650 97090
rect 5850 97020 6150 97090
rect 6350 97020 6650 97090
rect 6850 97020 7150 97090
rect 7350 97020 7650 97090
rect 7850 97020 8150 97090
rect 8350 97020 8650 97090
rect 8850 97020 9150 97090
rect 9350 97020 9650 97090
rect 9850 97020 10150 97090
rect 10350 97020 10650 97090
rect 10850 97020 11150 97090
rect 11350 97020 11650 97090
rect 11850 97020 12150 97090
rect 12350 97020 12650 97090
rect 12850 97020 13150 97090
rect 13350 97020 13650 97090
rect 13850 97020 14150 97090
rect 14350 97020 14650 97090
rect 14850 97020 15150 97090
rect 15350 97020 15650 97090
rect 15850 97020 16150 97090
rect 16350 97020 16650 97090
rect 16850 97020 17150 97090
rect 17350 97020 17650 97090
rect 17850 97020 18150 97090
rect 18350 97020 18650 97090
rect 18850 97020 19150 97090
rect 19350 97020 19650 97090
rect 19850 97020 20000 97090
rect -16000 96980 20000 97020
rect -16000 96910 -15850 96980
rect -15650 96910 -15350 96980
rect -15150 96910 -14850 96980
rect -14650 96910 -14350 96980
rect -14150 96910 -13850 96980
rect -13650 96910 -13350 96980
rect -13150 96910 -12850 96980
rect -12650 96910 -12350 96980
rect -12150 96910 -11850 96980
rect -11650 96910 -11350 96980
rect -11150 96910 -10850 96980
rect -10650 96910 -10350 96980
rect -10150 96910 -9850 96980
rect -9650 96910 -9350 96980
rect -9150 96910 -8850 96980
rect -8650 96910 -8350 96980
rect -8150 96910 -7850 96980
rect -7650 96910 -7350 96980
rect -7150 96910 -6850 96980
rect -6650 96910 -6350 96980
rect -6150 96910 -5850 96980
rect -5650 96910 -5350 96980
rect -5150 96910 -4850 96980
rect -4650 96910 -4350 96980
rect -4150 96910 -3850 96980
rect -3650 96910 -3350 96980
rect -3150 96910 -2850 96980
rect -2650 96910 -2350 96980
rect -2150 96910 -1850 96980
rect -1650 96910 -1350 96980
rect -1150 96910 -850 96980
rect -650 96910 -350 96980
rect -150 96910 150 96980
rect 350 96910 650 96980
rect 850 96910 1150 96980
rect 1350 96910 1650 96980
rect 1850 96910 2150 96980
rect 2350 96910 2650 96980
rect 2850 96910 3150 96980
rect 3350 96910 3650 96980
rect 3850 96910 4150 96980
rect 4350 96910 4650 96980
rect 4850 96910 5150 96980
rect 5350 96910 5650 96980
rect 5850 96910 6150 96980
rect 6350 96910 6650 96980
rect 6850 96910 7150 96980
rect 7350 96910 7650 96980
rect 7850 96910 8150 96980
rect 8350 96910 8650 96980
rect 8850 96910 9150 96980
rect 9350 96910 9650 96980
rect 9850 96910 10150 96980
rect 10350 96910 10650 96980
rect 10850 96910 11150 96980
rect 11350 96910 11650 96980
rect 11850 96910 12150 96980
rect 12350 96910 12650 96980
rect 12850 96910 13150 96980
rect 13350 96910 13650 96980
rect 13850 96910 14150 96980
rect 14350 96910 14650 96980
rect 14850 96910 15150 96980
rect 15350 96910 15650 96980
rect 15850 96910 16150 96980
rect 16350 96910 16650 96980
rect 16850 96910 17150 96980
rect 17350 96910 17650 96980
rect 17850 96910 18150 96980
rect 18350 96910 18650 96980
rect 18850 96910 19150 96980
rect 19350 96910 19650 96980
rect 19850 96910 20000 96980
rect -16000 96900 20000 96910
rect -16000 96880 -15880 96900
rect -15620 96880 -15380 96900
rect -15120 96880 -14880 96900
rect -14620 96880 -14380 96900
rect -14120 96880 -13880 96900
rect -13620 96880 -13380 96900
rect -13120 96880 -12880 96900
rect -12620 96880 -12380 96900
rect -12120 96880 -11880 96900
rect -11620 96880 -11380 96900
rect -11120 96880 -10880 96900
rect -10620 96880 -10380 96900
rect -10120 96880 -9880 96900
rect -9620 96880 -9380 96900
rect -9120 96880 -8880 96900
rect -8620 96880 -8380 96900
rect -8120 96880 -7880 96900
rect -7620 96880 -7380 96900
rect -7120 96880 -6880 96900
rect -6620 96880 -6380 96900
rect -6120 96880 -5880 96900
rect -5620 96880 -5380 96900
rect -5120 96880 -4880 96900
rect -4620 96880 -4380 96900
rect -4120 96880 -3880 96900
rect -3620 96880 -3380 96900
rect -3120 96880 -2880 96900
rect -2620 96880 -2380 96900
rect -2120 96880 -1880 96900
rect -1620 96880 -1380 96900
rect -1120 96880 -880 96900
rect -620 96880 -380 96900
rect -120 96880 120 96900
rect 380 96880 620 96900
rect 880 96880 1120 96900
rect 1380 96880 1620 96900
rect 1880 96880 2120 96900
rect 2380 96880 2620 96900
rect 2880 96880 3120 96900
rect 3380 96880 3620 96900
rect 3880 96880 4120 96900
rect 4380 96880 4620 96900
rect 4880 96880 5120 96900
rect 5380 96880 5620 96900
rect 5880 96880 6120 96900
rect 6380 96880 6620 96900
rect 6880 96880 7120 96900
rect 7380 96880 7620 96900
rect 7880 96880 8120 96900
rect 8380 96880 8620 96900
rect 8880 96880 9120 96900
rect 9380 96880 9620 96900
rect 9880 96880 10120 96900
rect 10380 96880 10620 96900
rect 10880 96880 11120 96900
rect 11380 96880 11620 96900
rect 11880 96880 12120 96900
rect 12380 96880 12620 96900
rect 12880 96880 13120 96900
rect 13380 96880 13620 96900
rect 13880 96880 14120 96900
rect 14380 96880 14620 96900
rect 14880 96880 15120 96900
rect 15380 96880 15620 96900
rect 15880 96880 16120 96900
rect 16380 96880 16620 96900
rect 16880 96880 17120 96900
rect 17380 96880 17620 96900
rect 17880 96880 18120 96900
rect 18380 96880 18620 96900
rect 18880 96880 19120 96900
rect 19380 96880 19620 96900
rect 19880 96880 20000 96900
rect -16000 96850 -15900 96880
rect -16000 96650 -15980 96850
rect -15910 96650 -15900 96850
rect -16000 96620 -15900 96650
rect -15600 96850 -15400 96880
rect -15600 96650 -15590 96850
rect -15520 96650 -15480 96850
rect -15410 96650 -15400 96850
rect -15600 96620 -15400 96650
rect -15100 96850 -14900 96880
rect -15100 96650 -15090 96850
rect -15020 96650 -14980 96850
rect -14910 96650 -14900 96850
rect -15100 96620 -14900 96650
rect -14600 96850 -14400 96880
rect -14600 96650 -14590 96850
rect -14520 96650 -14480 96850
rect -14410 96650 -14400 96850
rect -14600 96620 -14400 96650
rect -14100 96850 -13900 96880
rect -14100 96650 -14090 96850
rect -14020 96650 -13980 96850
rect -13910 96650 -13900 96850
rect -14100 96620 -13900 96650
rect -13600 96850 -13400 96880
rect -13600 96650 -13590 96850
rect -13520 96650 -13480 96850
rect -13410 96650 -13400 96850
rect -13600 96620 -13400 96650
rect -13100 96850 -12900 96880
rect -13100 96650 -13090 96850
rect -13020 96650 -12980 96850
rect -12910 96650 -12900 96850
rect -13100 96620 -12900 96650
rect -12600 96850 -12400 96880
rect -12600 96650 -12590 96850
rect -12520 96650 -12480 96850
rect -12410 96650 -12400 96850
rect -12600 96620 -12400 96650
rect -12100 96850 -11900 96880
rect -12100 96650 -12090 96850
rect -12020 96650 -11980 96850
rect -11910 96650 -11900 96850
rect -12100 96620 -11900 96650
rect -11600 96850 -11400 96880
rect -11600 96650 -11590 96850
rect -11520 96650 -11480 96850
rect -11410 96650 -11400 96850
rect -11600 96620 -11400 96650
rect -11100 96850 -10900 96880
rect -11100 96650 -11090 96850
rect -11020 96650 -10980 96850
rect -10910 96650 -10900 96850
rect -11100 96620 -10900 96650
rect -10600 96850 -10400 96880
rect -10600 96650 -10590 96850
rect -10520 96650 -10480 96850
rect -10410 96650 -10400 96850
rect -10600 96620 -10400 96650
rect -10100 96850 -9900 96880
rect -10100 96650 -10090 96850
rect -10020 96650 -9980 96850
rect -9910 96650 -9900 96850
rect -10100 96620 -9900 96650
rect -9600 96850 -9400 96880
rect -9600 96650 -9590 96850
rect -9520 96650 -9480 96850
rect -9410 96650 -9400 96850
rect -9600 96620 -9400 96650
rect -9100 96850 -8900 96880
rect -9100 96650 -9090 96850
rect -9020 96650 -8980 96850
rect -8910 96650 -8900 96850
rect -9100 96620 -8900 96650
rect -8600 96850 -8400 96880
rect -8600 96650 -8590 96850
rect -8520 96650 -8480 96850
rect -8410 96650 -8400 96850
rect -8600 96620 -8400 96650
rect -8100 96850 -7900 96880
rect -8100 96650 -8090 96850
rect -8020 96650 -7980 96850
rect -7910 96650 -7900 96850
rect -8100 96620 -7900 96650
rect -7600 96850 -7400 96880
rect -7600 96650 -7590 96850
rect -7520 96650 -7480 96850
rect -7410 96650 -7400 96850
rect -7600 96620 -7400 96650
rect -7100 96850 -6900 96880
rect -7100 96650 -7090 96850
rect -7020 96650 -6980 96850
rect -6910 96650 -6900 96850
rect -7100 96620 -6900 96650
rect -6600 96850 -6400 96880
rect -6600 96650 -6590 96850
rect -6520 96650 -6480 96850
rect -6410 96650 -6400 96850
rect -6600 96620 -6400 96650
rect -6100 96850 -5900 96880
rect -6100 96650 -6090 96850
rect -6020 96650 -5980 96850
rect -5910 96650 -5900 96850
rect -6100 96620 -5900 96650
rect -5600 96850 -5400 96880
rect -5600 96650 -5590 96850
rect -5520 96650 -5480 96850
rect -5410 96650 -5400 96850
rect -5600 96620 -5400 96650
rect -5100 96850 -4900 96880
rect -5100 96650 -5090 96850
rect -5020 96650 -4980 96850
rect -4910 96650 -4900 96850
rect -5100 96620 -4900 96650
rect -4600 96850 -4400 96880
rect -4600 96650 -4590 96850
rect -4520 96650 -4480 96850
rect -4410 96650 -4400 96850
rect -4600 96620 -4400 96650
rect -4100 96850 -3900 96880
rect -4100 96650 -4090 96850
rect -4020 96650 -3980 96850
rect -3910 96650 -3900 96850
rect -4100 96620 -3900 96650
rect -3600 96850 -3400 96880
rect -3600 96650 -3590 96850
rect -3520 96650 -3480 96850
rect -3410 96650 -3400 96850
rect -3600 96620 -3400 96650
rect -3100 96850 -2900 96880
rect -3100 96650 -3090 96850
rect -3020 96650 -2980 96850
rect -2910 96650 -2900 96850
rect -3100 96620 -2900 96650
rect -2600 96850 -2400 96880
rect -2600 96650 -2590 96850
rect -2520 96650 -2480 96850
rect -2410 96650 -2400 96850
rect -2600 96620 -2400 96650
rect -2100 96850 -1900 96880
rect -2100 96650 -2090 96850
rect -2020 96650 -1980 96850
rect -1910 96650 -1900 96850
rect -2100 96620 -1900 96650
rect -1600 96850 -1400 96880
rect -1600 96650 -1590 96850
rect -1520 96650 -1480 96850
rect -1410 96650 -1400 96850
rect -1600 96620 -1400 96650
rect -1100 96850 -900 96880
rect -1100 96650 -1090 96850
rect -1020 96650 -980 96850
rect -910 96650 -900 96850
rect -1100 96620 -900 96650
rect -600 96850 -400 96880
rect -600 96650 -590 96850
rect -520 96650 -480 96850
rect -410 96650 -400 96850
rect -600 96620 -400 96650
rect -100 96850 100 96880
rect -100 96650 -90 96850
rect -20 96650 20 96850
rect 90 96650 100 96850
rect -100 96620 100 96650
rect 400 96850 600 96880
rect 400 96650 410 96850
rect 480 96650 520 96850
rect 590 96650 600 96850
rect 400 96620 600 96650
rect 900 96850 1100 96880
rect 900 96650 910 96850
rect 980 96650 1020 96850
rect 1090 96650 1100 96850
rect 900 96620 1100 96650
rect 1400 96850 1600 96880
rect 1400 96650 1410 96850
rect 1480 96650 1520 96850
rect 1590 96650 1600 96850
rect 1400 96620 1600 96650
rect 1900 96850 2100 96880
rect 1900 96650 1910 96850
rect 1980 96650 2020 96850
rect 2090 96650 2100 96850
rect 1900 96620 2100 96650
rect 2400 96850 2600 96880
rect 2400 96650 2410 96850
rect 2480 96650 2520 96850
rect 2590 96650 2600 96850
rect 2400 96620 2600 96650
rect 2900 96850 3100 96880
rect 2900 96650 2910 96850
rect 2980 96650 3020 96850
rect 3090 96650 3100 96850
rect 2900 96620 3100 96650
rect 3400 96850 3600 96880
rect 3400 96650 3410 96850
rect 3480 96650 3520 96850
rect 3590 96650 3600 96850
rect 3400 96620 3600 96650
rect 3900 96850 4100 96880
rect 3900 96650 3910 96850
rect 3980 96650 4020 96850
rect 4090 96650 4100 96850
rect 3900 96620 4100 96650
rect 4400 96850 4600 96880
rect 4400 96650 4410 96850
rect 4480 96650 4520 96850
rect 4590 96650 4600 96850
rect 4400 96620 4600 96650
rect 4900 96850 5100 96880
rect 4900 96650 4910 96850
rect 4980 96650 5020 96850
rect 5090 96650 5100 96850
rect 4900 96620 5100 96650
rect 5400 96850 5600 96880
rect 5400 96650 5410 96850
rect 5480 96650 5520 96850
rect 5590 96650 5600 96850
rect 5400 96620 5600 96650
rect 5900 96850 6100 96880
rect 5900 96650 5910 96850
rect 5980 96650 6020 96850
rect 6090 96650 6100 96850
rect 5900 96620 6100 96650
rect 6400 96850 6600 96880
rect 6400 96650 6410 96850
rect 6480 96650 6520 96850
rect 6590 96650 6600 96850
rect 6400 96620 6600 96650
rect 6900 96850 7100 96880
rect 6900 96650 6910 96850
rect 6980 96650 7020 96850
rect 7090 96650 7100 96850
rect 6900 96620 7100 96650
rect 7400 96850 7600 96880
rect 7400 96650 7410 96850
rect 7480 96650 7520 96850
rect 7590 96650 7600 96850
rect 7400 96620 7600 96650
rect 7900 96850 8100 96880
rect 7900 96650 7910 96850
rect 7980 96650 8020 96850
rect 8090 96650 8100 96850
rect 7900 96620 8100 96650
rect 8400 96850 8600 96880
rect 8400 96650 8410 96850
rect 8480 96650 8520 96850
rect 8590 96650 8600 96850
rect 8400 96620 8600 96650
rect 8900 96850 9100 96880
rect 8900 96650 8910 96850
rect 8980 96650 9020 96850
rect 9090 96650 9100 96850
rect 8900 96620 9100 96650
rect 9400 96850 9600 96880
rect 9400 96650 9410 96850
rect 9480 96650 9520 96850
rect 9590 96650 9600 96850
rect 9400 96620 9600 96650
rect 9900 96850 10100 96880
rect 9900 96650 9910 96850
rect 9980 96650 10020 96850
rect 10090 96650 10100 96850
rect 9900 96620 10100 96650
rect 10400 96850 10600 96880
rect 10400 96650 10410 96850
rect 10480 96650 10520 96850
rect 10590 96650 10600 96850
rect 10400 96620 10600 96650
rect 10900 96850 11100 96880
rect 10900 96650 10910 96850
rect 10980 96650 11020 96850
rect 11090 96650 11100 96850
rect 10900 96620 11100 96650
rect 11400 96850 11600 96880
rect 11400 96650 11410 96850
rect 11480 96650 11520 96850
rect 11590 96650 11600 96850
rect 11400 96620 11600 96650
rect 11900 96850 12100 96880
rect 11900 96650 11910 96850
rect 11980 96650 12020 96850
rect 12090 96650 12100 96850
rect 11900 96620 12100 96650
rect 12400 96850 12600 96880
rect 12400 96650 12410 96850
rect 12480 96650 12520 96850
rect 12590 96650 12600 96850
rect 12400 96620 12600 96650
rect 12900 96850 13100 96880
rect 12900 96650 12910 96850
rect 12980 96650 13020 96850
rect 13090 96650 13100 96850
rect 12900 96620 13100 96650
rect 13400 96850 13600 96880
rect 13400 96650 13410 96850
rect 13480 96650 13520 96850
rect 13590 96650 13600 96850
rect 13400 96620 13600 96650
rect 13900 96850 14100 96880
rect 13900 96650 13910 96850
rect 13980 96650 14020 96850
rect 14090 96650 14100 96850
rect 13900 96620 14100 96650
rect 14400 96850 14600 96880
rect 14400 96650 14410 96850
rect 14480 96650 14520 96850
rect 14590 96650 14600 96850
rect 14400 96620 14600 96650
rect 14900 96850 15100 96880
rect 14900 96650 14910 96850
rect 14980 96650 15020 96850
rect 15090 96650 15100 96850
rect 14900 96620 15100 96650
rect 15400 96850 15600 96880
rect 15400 96650 15410 96850
rect 15480 96650 15520 96850
rect 15590 96650 15600 96850
rect 15400 96620 15600 96650
rect 15900 96850 16100 96880
rect 15900 96650 15910 96850
rect 15980 96650 16020 96850
rect 16090 96650 16100 96850
rect 15900 96620 16100 96650
rect 16400 96850 16600 96880
rect 16400 96650 16410 96850
rect 16480 96650 16520 96850
rect 16590 96650 16600 96850
rect 16400 96620 16600 96650
rect 16900 96850 17100 96880
rect 16900 96650 16910 96850
rect 16980 96650 17020 96850
rect 17090 96650 17100 96850
rect 16900 96620 17100 96650
rect 17400 96850 17600 96880
rect 17400 96650 17410 96850
rect 17480 96650 17520 96850
rect 17590 96650 17600 96850
rect 17400 96620 17600 96650
rect 17900 96850 18100 96880
rect 17900 96650 17910 96850
rect 17980 96650 18020 96850
rect 18090 96650 18100 96850
rect 17900 96620 18100 96650
rect 18400 96850 18600 96880
rect 18400 96650 18410 96850
rect 18480 96650 18520 96850
rect 18590 96650 18600 96850
rect 18400 96620 18600 96650
rect 18900 96850 19100 96880
rect 18900 96650 18910 96850
rect 18980 96650 19020 96850
rect 19090 96650 19100 96850
rect 18900 96620 19100 96650
rect 19400 96850 19600 96880
rect 19400 96650 19410 96850
rect 19480 96650 19520 96850
rect 19590 96650 19600 96850
rect 19400 96620 19600 96650
rect 19900 96850 20000 96880
rect 19900 96650 19910 96850
rect 19980 96650 20000 96850
rect 19900 96620 20000 96650
rect -16000 96600 -15880 96620
rect -15620 96600 -15380 96620
rect -15120 96600 -14880 96620
rect -14620 96600 -14380 96620
rect -14120 96600 -13880 96620
rect -13620 96600 -13380 96620
rect -13120 96600 -12880 96620
rect -12620 96600 -12380 96620
rect -12120 96600 -11880 96620
rect -11620 96600 -11380 96620
rect -11120 96600 -10880 96620
rect -10620 96600 -10380 96620
rect -10120 96600 -9880 96620
rect -9620 96600 -9380 96620
rect -9120 96600 -8880 96620
rect -8620 96600 -8380 96620
rect -8120 96600 -7880 96620
rect -7620 96600 -7380 96620
rect -7120 96600 -6880 96620
rect -6620 96600 -6380 96620
rect -6120 96600 -5880 96620
rect -5620 96600 -5380 96620
rect -5120 96600 -4880 96620
rect -4620 96600 -4380 96620
rect -4120 96600 -3880 96620
rect -3620 96600 -3380 96620
rect -3120 96600 -2880 96620
rect -2620 96600 -2380 96620
rect -2120 96600 -1880 96620
rect -1620 96600 -1380 96620
rect -1120 96600 -880 96620
rect -620 96600 -380 96620
rect -120 96600 120 96620
rect 380 96600 620 96620
rect 880 96600 1120 96620
rect 1380 96600 1620 96620
rect 1880 96600 2120 96620
rect 2380 96600 2620 96620
rect 2880 96600 3120 96620
rect 3380 96600 3620 96620
rect 3880 96600 4120 96620
rect 4380 96600 4620 96620
rect 4880 96600 5120 96620
rect 5380 96600 5620 96620
rect 5880 96600 6120 96620
rect 6380 96600 6620 96620
rect 6880 96600 7120 96620
rect 7380 96600 7620 96620
rect 7880 96600 8120 96620
rect 8380 96600 8620 96620
rect 8880 96600 9120 96620
rect 9380 96600 9620 96620
rect 9880 96600 10120 96620
rect 10380 96600 10620 96620
rect 10880 96600 11120 96620
rect 11380 96600 11620 96620
rect 11880 96600 12120 96620
rect 12380 96600 12620 96620
rect 12880 96600 13120 96620
rect 13380 96600 13620 96620
rect 13880 96600 14120 96620
rect 14380 96600 14620 96620
rect 14880 96600 15120 96620
rect 15380 96600 15620 96620
rect 15880 96600 16120 96620
rect 16380 96600 16620 96620
rect 16880 96600 17120 96620
rect 17380 96600 17620 96620
rect 17880 96600 18120 96620
rect 18380 96600 18620 96620
rect 18880 96600 19120 96620
rect 19380 96600 19620 96620
rect 19880 96600 20000 96620
rect -16000 96590 20000 96600
rect -16000 96520 -15850 96590
rect -15650 96520 -15350 96590
rect -15150 96520 -14850 96590
rect -14650 96520 -14350 96590
rect -14150 96520 -13850 96590
rect -13650 96520 -13350 96590
rect -13150 96520 -12850 96590
rect -12650 96520 -12350 96590
rect -12150 96520 -11850 96590
rect -11650 96520 -11350 96590
rect -11150 96520 -10850 96590
rect -10650 96520 -10350 96590
rect -10150 96520 -9850 96590
rect -9650 96520 -9350 96590
rect -9150 96520 -8850 96590
rect -8650 96520 -8350 96590
rect -8150 96520 -7850 96590
rect -7650 96520 -7350 96590
rect -7150 96520 -6850 96590
rect -6650 96520 -6350 96590
rect -6150 96520 -5850 96590
rect -5650 96520 -5350 96590
rect -5150 96520 -4850 96590
rect -4650 96520 -4350 96590
rect -4150 96520 -3850 96590
rect -3650 96520 -3350 96590
rect -3150 96520 -2850 96590
rect -2650 96520 -2350 96590
rect -2150 96520 -1850 96590
rect -1650 96520 -1350 96590
rect -1150 96520 -850 96590
rect -650 96520 -350 96590
rect -150 96520 150 96590
rect 350 96520 650 96590
rect 850 96520 1150 96590
rect 1350 96520 1650 96590
rect 1850 96520 2150 96590
rect 2350 96520 2650 96590
rect 2850 96520 3150 96590
rect 3350 96520 3650 96590
rect 3850 96520 4150 96590
rect 4350 96520 4650 96590
rect 4850 96520 5150 96590
rect 5350 96520 5650 96590
rect 5850 96520 6150 96590
rect 6350 96520 6650 96590
rect 6850 96520 7150 96590
rect 7350 96520 7650 96590
rect 7850 96520 8150 96590
rect 8350 96520 8650 96590
rect 8850 96520 9150 96590
rect 9350 96520 9650 96590
rect 9850 96520 10150 96590
rect 10350 96520 10650 96590
rect 10850 96520 11150 96590
rect 11350 96520 11650 96590
rect 11850 96520 12150 96590
rect 12350 96520 12650 96590
rect 12850 96520 13150 96590
rect 13350 96520 13650 96590
rect 13850 96520 14150 96590
rect 14350 96520 14650 96590
rect 14850 96520 15150 96590
rect 15350 96520 15650 96590
rect 15850 96520 16150 96590
rect 16350 96520 16650 96590
rect 16850 96520 17150 96590
rect 17350 96520 17650 96590
rect 17850 96520 18150 96590
rect 18350 96520 18650 96590
rect 18850 96520 19150 96590
rect 19350 96520 19650 96590
rect 19850 96520 20000 96590
rect -16000 96480 20000 96520
rect -16000 96410 -15850 96480
rect -15650 96410 -15350 96480
rect -15150 96410 -14850 96480
rect -14650 96410 -14350 96480
rect -14150 96410 -13850 96480
rect -13650 96410 -13350 96480
rect -13150 96410 -12850 96480
rect -12650 96410 -12350 96480
rect -12150 96410 -11850 96480
rect -11650 96410 -11350 96480
rect -11150 96410 -10850 96480
rect -10650 96410 -10350 96480
rect -10150 96410 -9850 96480
rect -9650 96410 -9350 96480
rect -9150 96410 -8850 96480
rect -8650 96410 -8350 96480
rect -8150 96410 -7850 96480
rect -7650 96410 -7350 96480
rect -7150 96410 -6850 96480
rect -6650 96410 -6350 96480
rect -6150 96410 -5850 96480
rect -5650 96410 -5350 96480
rect -5150 96410 -4850 96480
rect -4650 96410 -4350 96480
rect -4150 96410 -3850 96480
rect -3650 96410 -3350 96480
rect -3150 96410 -2850 96480
rect -2650 96410 -2350 96480
rect -2150 96410 -1850 96480
rect -1650 96410 -1350 96480
rect -1150 96410 -850 96480
rect -650 96410 -350 96480
rect -150 96410 150 96480
rect 350 96410 650 96480
rect 850 96410 1150 96480
rect 1350 96410 1650 96480
rect 1850 96410 2150 96480
rect 2350 96410 2650 96480
rect 2850 96410 3150 96480
rect 3350 96410 3650 96480
rect 3850 96410 4150 96480
rect 4350 96410 4650 96480
rect 4850 96410 5150 96480
rect 5350 96410 5650 96480
rect 5850 96410 6150 96480
rect 6350 96410 6650 96480
rect 6850 96410 7150 96480
rect 7350 96410 7650 96480
rect 7850 96410 8150 96480
rect 8350 96410 8650 96480
rect 8850 96410 9150 96480
rect 9350 96410 9650 96480
rect 9850 96410 10150 96480
rect 10350 96410 10650 96480
rect 10850 96410 11150 96480
rect 11350 96410 11650 96480
rect 11850 96410 12150 96480
rect 12350 96410 12650 96480
rect 12850 96410 13150 96480
rect 13350 96410 13650 96480
rect 13850 96410 14150 96480
rect 14350 96410 14650 96480
rect 14850 96410 15150 96480
rect 15350 96410 15650 96480
rect 15850 96410 16150 96480
rect 16350 96410 16650 96480
rect 16850 96410 17150 96480
rect 17350 96410 17650 96480
rect 17850 96410 18150 96480
rect 18350 96410 18650 96480
rect 18850 96410 19150 96480
rect 19350 96410 19650 96480
rect 19850 96410 20000 96480
rect -16000 96400 20000 96410
rect -16000 96380 -15880 96400
rect -15620 96380 -15380 96400
rect -15120 96380 -14880 96400
rect -14620 96380 -14380 96400
rect -14120 96380 -13880 96400
rect -13620 96380 -13380 96400
rect -13120 96380 -12880 96400
rect -12620 96380 -12380 96400
rect -12120 96380 -11880 96400
rect -11620 96380 -11380 96400
rect -11120 96380 -10880 96400
rect -10620 96380 -10380 96400
rect -10120 96380 -9880 96400
rect -9620 96380 -9380 96400
rect -9120 96380 -8880 96400
rect -8620 96380 -8380 96400
rect -8120 96380 -7880 96400
rect -7620 96380 -7380 96400
rect -7120 96380 -6880 96400
rect -6620 96380 -6380 96400
rect -6120 96380 -5880 96400
rect -5620 96380 -5380 96400
rect -5120 96380 -4880 96400
rect -4620 96380 -4380 96400
rect -4120 96380 -3880 96400
rect -3620 96380 -3380 96400
rect -3120 96380 -2880 96400
rect -2620 96380 -2380 96400
rect -2120 96380 -1880 96400
rect -1620 96380 -1380 96400
rect -1120 96380 -880 96400
rect -620 96380 -380 96400
rect -120 96380 120 96400
rect 380 96380 620 96400
rect 880 96380 1120 96400
rect 1380 96380 1620 96400
rect 1880 96380 2120 96400
rect 2380 96380 2620 96400
rect 2880 96380 3120 96400
rect 3380 96380 3620 96400
rect 3880 96380 4120 96400
rect 4380 96380 4620 96400
rect 4880 96380 5120 96400
rect 5380 96380 5620 96400
rect 5880 96380 6120 96400
rect 6380 96380 6620 96400
rect 6880 96380 7120 96400
rect 7380 96380 7620 96400
rect 7880 96380 8120 96400
rect 8380 96380 8620 96400
rect 8880 96380 9120 96400
rect 9380 96380 9620 96400
rect 9880 96380 10120 96400
rect 10380 96380 10620 96400
rect 10880 96380 11120 96400
rect 11380 96380 11620 96400
rect 11880 96380 12120 96400
rect 12380 96380 12620 96400
rect 12880 96380 13120 96400
rect 13380 96380 13620 96400
rect 13880 96380 14120 96400
rect 14380 96380 14620 96400
rect 14880 96380 15120 96400
rect 15380 96380 15620 96400
rect 15880 96380 16120 96400
rect 16380 96380 16620 96400
rect 16880 96380 17120 96400
rect 17380 96380 17620 96400
rect 17880 96380 18120 96400
rect 18380 96380 18620 96400
rect 18880 96380 19120 96400
rect 19380 96380 19620 96400
rect 19880 96380 20000 96400
rect -16000 96350 -15900 96380
rect -16000 96150 -15980 96350
rect -15910 96150 -15900 96350
rect -16000 96120 -15900 96150
rect -15600 96350 -15400 96380
rect -15600 96150 -15590 96350
rect -15520 96150 -15480 96350
rect -15410 96150 -15400 96350
rect -15600 96120 -15400 96150
rect -15100 96350 -14900 96380
rect -15100 96150 -15090 96350
rect -15020 96150 -14980 96350
rect -14910 96150 -14900 96350
rect -15100 96120 -14900 96150
rect -14600 96350 -14400 96380
rect -14600 96150 -14590 96350
rect -14520 96150 -14480 96350
rect -14410 96150 -14400 96350
rect -14600 96120 -14400 96150
rect -14100 96350 -13900 96380
rect -14100 96150 -14090 96350
rect -14020 96150 -13980 96350
rect -13910 96150 -13900 96350
rect -14100 96120 -13900 96150
rect -13600 96350 -13400 96380
rect -13600 96150 -13590 96350
rect -13520 96150 -13480 96350
rect -13410 96150 -13400 96350
rect -13600 96120 -13400 96150
rect -13100 96350 -12900 96380
rect -13100 96150 -13090 96350
rect -13020 96150 -12980 96350
rect -12910 96150 -12900 96350
rect -13100 96120 -12900 96150
rect -12600 96350 -12400 96380
rect -12600 96150 -12590 96350
rect -12520 96150 -12480 96350
rect -12410 96150 -12400 96350
rect -12600 96120 -12400 96150
rect -12100 96350 -11900 96380
rect -12100 96150 -12090 96350
rect -12020 96150 -11980 96350
rect -11910 96150 -11900 96350
rect -12100 96120 -11900 96150
rect -11600 96350 -11400 96380
rect -11600 96150 -11590 96350
rect -11520 96150 -11480 96350
rect -11410 96150 -11400 96350
rect -11600 96120 -11400 96150
rect -11100 96350 -10900 96380
rect -11100 96150 -11090 96350
rect -11020 96150 -10980 96350
rect -10910 96150 -10900 96350
rect -11100 96120 -10900 96150
rect -10600 96350 -10400 96380
rect -10600 96150 -10590 96350
rect -10520 96150 -10480 96350
rect -10410 96150 -10400 96350
rect -10600 96120 -10400 96150
rect -10100 96350 -9900 96380
rect -10100 96150 -10090 96350
rect -10020 96150 -9980 96350
rect -9910 96150 -9900 96350
rect -10100 96120 -9900 96150
rect -9600 96350 -9400 96380
rect -9600 96150 -9590 96350
rect -9520 96150 -9480 96350
rect -9410 96150 -9400 96350
rect -9600 96120 -9400 96150
rect -9100 96350 -8900 96380
rect -9100 96150 -9090 96350
rect -9020 96150 -8980 96350
rect -8910 96150 -8900 96350
rect -9100 96120 -8900 96150
rect -8600 96350 -8400 96380
rect -8600 96150 -8590 96350
rect -8520 96150 -8480 96350
rect -8410 96150 -8400 96350
rect -8600 96120 -8400 96150
rect -8100 96350 -7900 96380
rect -8100 96150 -8090 96350
rect -8020 96150 -7980 96350
rect -7910 96150 -7900 96350
rect -8100 96120 -7900 96150
rect -7600 96350 -7400 96380
rect -7600 96150 -7590 96350
rect -7520 96150 -7480 96350
rect -7410 96150 -7400 96350
rect -7600 96120 -7400 96150
rect -7100 96350 -6900 96380
rect -7100 96150 -7090 96350
rect -7020 96150 -6980 96350
rect -6910 96150 -6900 96350
rect -7100 96120 -6900 96150
rect -6600 96350 -6400 96380
rect -6600 96150 -6590 96350
rect -6520 96150 -6480 96350
rect -6410 96150 -6400 96350
rect -6600 96120 -6400 96150
rect -6100 96350 -5900 96380
rect -6100 96150 -6090 96350
rect -6020 96150 -5980 96350
rect -5910 96150 -5900 96350
rect -6100 96120 -5900 96150
rect -5600 96350 -5400 96380
rect -5600 96150 -5590 96350
rect -5520 96150 -5480 96350
rect -5410 96150 -5400 96350
rect -5600 96120 -5400 96150
rect -5100 96350 -4900 96380
rect -5100 96150 -5090 96350
rect -5020 96150 -4980 96350
rect -4910 96150 -4900 96350
rect -5100 96120 -4900 96150
rect -4600 96350 -4400 96380
rect -4600 96150 -4590 96350
rect -4520 96150 -4480 96350
rect -4410 96150 -4400 96350
rect -4600 96120 -4400 96150
rect -4100 96350 -3900 96380
rect -4100 96150 -4090 96350
rect -4020 96150 -3980 96350
rect -3910 96150 -3900 96350
rect -4100 96120 -3900 96150
rect -3600 96350 -3400 96380
rect -3600 96150 -3590 96350
rect -3520 96150 -3480 96350
rect -3410 96150 -3400 96350
rect -3600 96120 -3400 96150
rect -3100 96350 -2900 96380
rect -3100 96150 -3090 96350
rect -3020 96150 -2980 96350
rect -2910 96150 -2900 96350
rect -3100 96120 -2900 96150
rect -2600 96350 -2400 96380
rect -2600 96150 -2590 96350
rect -2520 96150 -2480 96350
rect -2410 96150 -2400 96350
rect -2600 96120 -2400 96150
rect -2100 96350 -1900 96380
rect -2100 96150 -2090 96350
rect -2020 96150 -1980 96350
rect -1910 96150 -1900 96350
rect -2100 96120 -1900 96150
rect -1600 96350 -1400 96380
rect -1600 96150 -1590 96350
rect -1520 96150 -1480 96350
rect -1410 96150 -1400 96350
rect -1600 96120 -1400 96150
rect -1100 96350 -900 96380
rect -1100 96150 -1090 96350
rect -1020 96150 -980 96350
rect -910 96150 -900 96350
rect -1100 96120 -900 96150
rect -600 96350 -400 96380
rect -600 96150 -590 96350
rect -520 96150 -480 96350
rect -410 96150 -400 96350
rect -600 96120 -400 96150
rect -100 96350 100 96380
rect -100 96150 -90 96350
rect -20 96150 20 96350
rect 90 96150 100 96350
rect -100 96120 100 96150
rect 400 96350 600 96380
rect 400 96150 410 96350
rect 480 96150 520 96350
rect 590 96150 600 96350
rect 400 96120 600 96150
rect 900 96350 1100 96380
rect 900 96150 910 96350
rect 980 96150 1020 96350
rect 1090 96150 1100 96350
rect 900 96120 1100 96150
rect 1400 96350 1600 96380
rect 1400 96150 1410 96350
rect 1480 96150 1520 96350
rect 1590 96150 1600 96350
rect 1400 96120 1600 96150
rect 1900 96350 2100 96380
rect 1900 96150 1910 96350
rect 1980 96150 2020 96350
rect 2090 96150 2100 96350
rect 1900 96120 2100 96150
rect 2400 96350 2600 96380
rect 2400 96150 2410 96350
rect 2480 96150 2520 96350
rect 2590 96150 2600 96350
rect 2400 96120 2600 96150
rect 2900 96350 3100 96380
rect 2900 96150 2910 96350
rect 2980 96150 3020 96350
rect 3090 96150 3100 96350
rect 2900 96120 3100 96150
rect 3400 96350 3600 96380
rect 3400 96150 3410 96350
rect 3480 96150 3520 96350
rect 3590 96150 3600 96350
rect 3400 96120 3600 96150
rect 3900 96350 4100 96380
rect 3900 96150 3910 96350
rect 3980 96150 4020 96350
rect 4090 96150 4100 96350
rect 3900 96120 4100 96150
rect 4400 96350 4600 96380
rect 4400 96150 4410 96350
rect 4480 96150 4520 96350
rect 4590 96150 4600 96350
rect 4400 96120 4600 96150
rect 4900 96350 5100 96380
rect 4900 96150 4910 96350
rect 4980 96150 5020 96350
rect 5090 96150 5100 96350
rect 4900 96120 5100 96150
rect 5400 96350 5600 96380
rect 5400 96150 5410 96350
rect 5480 96150 5520 96350
rect 5590 96150 5600 96350
rect 5400 96120 5600 96150
rect 5900 96350 6100 96380
rect 5900 96150 5910 96350
rect 5980 96150 6020 96350
rect 6090 96150 6100 96350
rect 5900 96120 6100 96150
rect 6400 96350 6600 96380
rect 6400 96150 6410 96350
rect 6480 96150 6520 96350
rect 6590 96150 6600 96350
rect 6400 96120 6600 96150
rect 6900 96350 7100 96380
rect 6900 96150 6910 96350
rect 6980 96150 7020 96350
rect 7090 96150 7100 96350
rect 6900 96120 7100 96150
rect 7400 96350 7600 96380
rect 7400 96150 7410 96350
rect 7480 96150 7520 96350
rect 7590 96150 7600 96350
rect 7400 96120 7600 96150
rect 7900 96350 8100 96380
rect 7900 96150 7910 96350
rect 7980 96150 8020 96350
rect 8090 96150 8100 96350
rect 7900 96120 8100 96150
rect 8400 96350 8600 96380
rect 8400 96150 8410 96350
rect 8480 96150 8520 96350
rect 8590 96150 8600 96350
rect 8400 96120 8600 96150
rect 8900 96350 9100 96380
rect 8900 96150 8910 96350
rect 8980 96150 9020 96350
rect 9090 96150 9100 96350
rect 8900 96120 9100 96150
rect 9400 96350 9600 96380
rect 9400 96150 9410 96350
rect 9480 96150 9520 96350
rect 9590 96150 9600 96350
rect 9400 96120 9600 96150
rect 9900 96350 10100 96380
rect 9900 96150 9910 96350
rect 9980 96150 10020 96350
rect 10090 96150 10100 96350
rect 9900 96120 10100 96150
rect 10400 96350 10600 96380
rect 10400 96150 10410 96350
rect 10480 96150 10520 96350
rect 10590 96150 10600 96350
rect 10400 96120 10600 96150
rect 10900 96350 11100 96380
rect 10900 96150 10910 96350
rect 10980 96150 11020 96350
rect 11090 96150 11100 96350
rect 10900 96120 11100 96150
rect 11400 96350 11600 96380
rect 11400 96150 11410 96350
rect 11480 96150 11520 96350
rect 11590 96150 11600 96350
rect 11400 96120 11600 96150
rect 11900 96350 12100 96380
rect 11900 96150 11910 96350
rect 11980 96150 12020 96350
rect 12090 96150 12100 96350
rect 11900 96120 12100 96150
rect 12400 96350 12600 96380
rect 12400 96150 12410 96350
rect 12480 96150 12520 96350
rect 12590 96150 12600 96350
rect 12400 96120 12600 96150
rect 12900 96350 13100 96380
rect 12900 96150 12910 96350
rect 12980 96150 13020 96350
rect 13090 96150 13100 96350
rect 12900 96120 13100 96150
rect 13400 96350 13600 96380
rect 13400 96150 13410 96350
rect 13480 96150 13520 96350
rect 13590 96150 13600 96350
rect 13400 96120 13600 96150
rect 13900 96350 14100 96380
rect 13900 96150 13910 96350
rect 13980 96150 14020 96350
rect 14090 96150 14100 96350
rect 13900 96120 14100 96150
rect 14400 96350 14600 96380
rect 14400 96150 14410 96350
rect 14480 96150 14520 96350
rect 14590 96150 14600 96350
rect 14400 96120 14600 96150
rect 14900 96350 15100 96380
rect 14900 96150 14910 96350
rect 14980 96150 15020 96350
rect 15090 96150 15100 96350
rect 14900 96120 15100 96150
rect 15400 96350 15600 96380
rect 15400 96150 15410 96350
rect 15480 96150 15520 96350
rect 15590 96150 15600 96350
rect 15400 96120 15600 96150
rect 15900 96350 16100 96380
rect 15900 96150 15910 96350
rect 15980 96150 16020 96350
rect 16090 96150 16100 96350
rect 15900 96120 16100 96150
rect 16400 96350 16600 96380
rect 16400 96150 16410 96350
rect 16480 96150 16520 96350
rect 16590 96150 16600 96350
rect 16400 96120 16600 96150
rect 16900 96350 17100 96380
rect 16900 96150 16910 96350
rect 16980 96150 17020 96350
rect 17090 96150 17100 96350
rect 16900 96120 17100 96150
rect 17400 96350 17600 96380
rect 17400 96150 17410 96350
rect 17480 96150 17520 96350
rect 17590 96150 17600 96350
rect 17400 96120 17600 96150
rect 17900 96350 18100 96380
rect 17900 96150 17910 96350
rect 17980 96150 18020 96350
rect 18090 96150 18100 96350
rect 17900 96120 18100 96150
rect 18400 96350 18600 96380
rect 18400 96150 18410 96350
rect 18480 96150 18520 96350
rect 18590 96150 18600 96350
rect 18400 96120 18600 96150
rect 18900 96350 19100 96380
rect 18900 96150 18910 96350
rect 18980 96150 19020 96350
rect 19090 96150 19100 96350
rect 18900 96120 19100 96150
rect 19400 96350 19600 96380
rect 19400 96150 19410 96350
rect 19480 96150 19520 96350
rect 19590 96150 19600 96350
rect 19400 96120 19600 96150
rect 19900 96350 20000 96380
rect 19900 96150 19910 96350
rect 19980 96150 20000 96350
rect 19900 96120 20000 96150
rect -16000 96100 -15880 96120
rect -15620 96100 -15380 96120
rect -15120 96100 -14880 96120
rect -14620 96100 -14380 96120
rect -14120 96100 -13880 96120
rect -13620 96100 -13380 96120
rect -13120 96100 -12880 96120
rect -12620 96100 -12380 96120
rect -12120 96100 -11880 96120
rect -11620 96100 -11380 96120
rect -11120 96100 -10880 96120
rect -10620 96100 -10380 96120
rect -10120 96100 -9880 96120
rect -9620 96100 -9380 96120
rect -9120 96100 -8880 96120
rect -8620 96100 -8380 96120
rect -8120 96100 -7880 96120
rect -7620 96100 -7380 96120
rect -7120 96100 -6880 96120
rect -6620 96100 -6380 96120
rect -6120 96100 -5880 96120
rect -5620 96100 -5380 96120
rect -5120 96100 -4880 96120
rect -4620 96100 -4380 96120
rect -4120 96100 -3880 96120
rect -3620 96100 -3380 96120
rect -3120 96100 -2880 96120
rect -2620 96100 -2380 96120
rect -2120 96100 -1880 96120
rect -1620 96100 -1380 96120
rect -1120 96100 -880 96120
rect -620 96100 -380 96120
rect -120 96100 120 96120
rect 380 96100 620 96120
rect 880 96100 1120 96120
rect 1380 96100 1620 96120
rect 1880 96100 2120 96120
rect 2380 96100 2620 96120
rect 2880 96100 3120 96120
rect 3380 96100 3620 96120
rect 3880 96100 4120 96120
rect 4380 96100 4620 96120
rect 4880 96100 5120 96120
rect 5380 96100 5620 96120
rect 5880 96100 6120 96120
rect 6380 96100 6620 96120
rect 6880 96100 7120 96120
rect 7380 96100 7620 96120
rect 7880 96100 8120 96120
rect 8380 96100 8620 96120
rect 8880 96100 9120 96120
rect 9380 96100 9620 96120
rect 9880 96100 10120 96120
rect 10380 96100 10620 96120
rect 10880 96100 11120 96120
rect 11380 96100 11620 96120
rect 11880 96100 12120 96120
rect 12380 96100 12620 96120
rect 12880 96100 13120 96120
rect 13380 96100 13620 96120
rect 13880 96100 14120 96120
rect 14380 96100 14620 96120
rect 14880 96100 15120 96120
rect 15380 96100 15620 96120
rect 15880 96100 16120 96120
rect 16380 96100 16620 96120
rect 16880 96100 17120 96120
rect 17380 96100 17620 96120
rect 17880 96100 18120 96120
rect 18380 96100 18620 96120
rect 18880 96100 19120 96120
rect 19380 96100 19620 96120
rect 19880 96100 20000 96120
rect -16000 96090 20000 96100
rect -16000 96020 -15850 96090
rect -15650 96020 -15350 96090
rect -15150 96020 -14850 96090
rect -14650 96020 -14350 96090
rect -14150 96020 -13850 96090
rect -13650 96020 -13350 96090
rect -13150 96020 -12850 96090
rect -12650 96020 -12350 96090
rect -12150 96020 -11850 96090
rect -11650 96020 -11350 96090
rect -11150 96020 -10850 96090
rect -10650 96020 -10350 96090
rect -10150 96020 -9850 96090
rect -9650 96020 -9350 96090
rect -9150 96020 -8850 96090
rect -8650 96020 -8350 96090
rect -8150 96020 -7850 96090
rect -7650 96020 -7350 96090
rect -7150 96020 -6850 96090
rect -6650 96020 -6350 96090
rect -6150 96020 -5850 96090
rect -5650 96020 -5350 96090
rect -5150 96020 -4850 96090
rect -4650 96020 -4350 96090
rect -4150 96020 -3850 96090
rect -3650 96020 -3350 96090
rect -3150 96020 -2850 96090
rect -2650 96020 -2350 96090
rect -2150 96020 -1850 96090
rect -1650 96020 -1350 96090
rect -1150 96020 -850 96090
rect -650 96020 -350 96090
rect -150 96020 150 96090
rect 350 96020 650 96090
rect 850 96020 1150 96090
rect 1350 96020 1650 96090
rect 1850 96020 2150 96090
rect 2350 96020 2650 96090
rect 2850 96020 3150 96090
rect 3350 96020 3650 96090
rect 3850 96020 4150 96090
rect 4350 96020 4650 96090
rect 4850 96020 5150 96090
rect 5350 96020 5650 96090
rect 5850 96020 6150 96090
rect 6350 96020 6650 96090
rect 6850 96020 7150 96090
rect 7350 96020 7650 96090
rect 7850 96020 8150 96090
rect 8350 96020 8650 96090
rect 8850 96020 9150 96090
rect 9350 96020 9650 96090
rect 9850 96020 10150 96090
rect 10350 96020 10650 96090
rect 10850 96020 11150 96090
rect 11350 96020 11650 96090
rect 11850 96020 12150 96090
rect 12350 96020 12650 96090
rect 12850 96020 13150 96090
rect 13350 96020 13650 96090
rect 13850 96020 14150 96090
rect 14350 96020 14650 96090
rect 14850 96020 15150 96090
rect 15350 96020 15650 96090
rect 15850 96020 16150 96090
rect 16350 96020 16650 96090
rect 16850 96020 17150 96090
rect 17350 96020 17650 96090
rect 17850 96020 18150 96090
rect 18350 96020 18650 96090
rect 18850 96020 19150 96090
rect 19350 96020 19650 96090
rect 19850 96020 20000 96090
rect -16000 95980 20000 96020
rect -16000 95910 -15850 95980
rect -15650 95910 -15350 95980
rect -15150 95910 -14850 95980
rect -14650 95910 -14350 95980
rect -14150 95910 -13850 95980
rect -13650 95910 -13350 95980
rect -13150 95910 -12850 95980
rect -12650 95910 -12350 95980
rect -12150 95910 -11850 95980
rect -11650 95910 -11350 95980
rect -11150 95910 -10850 95980
rect -10650 95910 -10350 95980
rect -10150 95910 -9850 95980
rect -9650 95910 -9350 95980
rect -9150 95910 -8850 95980
rect -8650 95910 -8350 95980
rect -8150 95910 -7850 95980
rect -7650 95910 -7350 95980
rect -7150 95910 -6850 95980
rect -6650 95910 -6350 95980
rect -6150 95910 -5850 95980
rect -5650 95910 -5350 95980
rect -5150 95910 -4850 95980
rect -4650 95910 -4350 95980
rect -4150 95910 -3850 95980
rect -3650 95910 -3350 95980
rect -3150 95910 -2850 95980
rect -2650 95910 -2350 95980
rect -2150 95910 -1850 95980
rect -1650 95910 -1350 95980
rect -1150 95910 -850 95980
rect -650 95910 -350 95980
rect -150 95910 150 95980
rect 350 95910 650 95980
rect 850 95910 1150 95980
rect 1350 95910 1650 95980
rect 1850 95910 2150 95980
rect 2350 95910 2650 95980
rect 2850 95910 3150 95980
rect 3350 95910 3650 95980
rect 3850 95910 4150 95980
rect 4350 95910 4650 95980
rect 4850 95910 5150 95980
rect 5350 95910 5650 95980
rect 5850 95910 6150 95980
rect 6350 95910 6650 95980
rect 6850 95910 7150 95980
rect 7350 95910 7650 95980
rect 7850 95910 8150 95980
rect 8350 95910 8650 95980
rect 8850 95910 9150 95980
rect 9350 95910 9650 95980
rect 9850 95910 10150 95980
rect 10350 95910 10650 95980
rect 10850 95910 11150 95980
rect 11350 95910 11650 95980
rect 11850 95910 12150 95980
rect 12350 95910 12650 95980
rect 12850 95910 13150 95980
rect 13350 95910 13650 95980
rect 13850 95910 14150 95980
rect 14350 95910 14650 95980
rect 14850 95910 15150 95980
rect 15350 95910 15650 95980
rect 15850 95910 16150 95980
rect 16350 95910 16650 95980
rect 16850 95910 17150 95980
rect 17350 95910 17650 95980
rect 17850 95910 18150 95980
rect 18350 95910 18650 95980
rect 18850 95910 19150 95980
rect 19350 95910 19650 95980
rect 19850 95910 20000 95980
rect -16000 95900 20000 95910
rect -16000 95880 -15880 95900
rect -15620 95880 -15380 95900
rect -15120 95880 -14880 95900
rect -14620 95880 -14380 95900
rect -14120 95880 -13880 95900
rect -13620 95880 -13380 95900
rect -13120 95880 -12880 95900
rect -12620 95880 -12380 95900
rect -12120 95880 -11880 95900
rect -11620 95880 -11380 95900
rect -11120 95880 -10880 95900
rect -10620 95880 -10380 95900
rect -10120 95880 -9880 95900
rect -9620 95880 -9380 95900
rect -9120 95880 -8880 95900
rect -8620 95880 -8380 95900
rect -8120 95880 -7880 95900
rect -7620 95880 -7380 95900
rect -7120 95880 -6880 95900
rect -6620 95880 -6380 95900
rect -6120 95880 -5880 95900
rect -5620 95880 -5380 95900
rect -5120 95880 -4880 95900
rect -4620 95880 -4380 95900
rect -4120 95880 -3880 95900
rect -3620 95880 -3380 95900
rect -3120 95880 -2880 95900
rect -2620 95880 -2380 95900
rect -2120 95880 -1880 95900
rect -1620 95880 -1380 95900
rect -1120 95880 -880 95900
rect -620 95880 -380 95900
rect -120 95880 120 95900
rect 380 95880 620 95900
rect 880 95880 1120 95900
rect 1380 95880 1620 95900
rect 1880 95880 2120 95900
rect 2380 95880 2620 95900
rect 2880 95880 3120 95900
rect 3380 95880 3620 95900
rect 3880 95880 4120 95900
rect 4380 95880 4620 95900
rect 4880 95880 5120 95900
rect 5380 95880 5620 95900
rect 5880 95880 6120 95900
rect 6380 95880 6620 95900
rect 6880 95880 7120 95900
rect 7380 95880 7620 95900
rect 7880 95880 8120 95900
rect 8380 95880 8620 95900
rect 8880 95880 9120 95900
rect 9380 95880 9620 95900
rect 9880 95880 10120 95900
rect 10380 95880 10620 95900
rect 10880 95880 11120 95900
rect 11380 95880 11620 95900
rect 11880 95880 12120 95900
rect 12380 95880 12620 95900
rect 12880 95880 13120 95900
rect 13380 95880 13620 95900
rect 13880 95880 14120 95900
rect 14380 95880 14620 95900
rect 14880 95880 15120 95900
rect 15380 95880 15620 95900
rect 15880 95880 16120 95900
rect 16380 95880 16620 95900
rect 16880 95880 17120 95900
rect 17380 95880 17620 95900
rect 17880 95880 18120 95900
rect 18380 95880 18620 95900
rect 18880 95880 19120 95900
rect 19380 95880 19620 95900
rect 19880 95880 20000 95900
rect -16000 95850 -15900 95880
rect -16000 95650 -15980 95850
rect -15910 95650 -15900 95850
rect -16000 95620 -15900 95650
rect -15600 95850 -15400 95880
rect -15600 95650 -15590 95850
rect -15520 95650 -15480 95850
rect -15410 95650 -15400 95850
rect -15600 95620 -15400 95650
rect -15100 95850 -14900 95880
rect -15100 95650 -15090 95850
rect -15020 95650 -14980 95850
rect -14910 95650 -14900 95850
rect -15100 95620 -14900 95650
rect -14600 95850 -14400 95880
rect -14600 95650 -14590 95850
rect -14520 95650 -14480 95850
rect -14410 95650 -14400 95850
rect -14600 95620 -14400 95650
rect -14100 95850 -13900 95880
rect -14100 95650 -14090 95850
rect -14020 95650 -13980 95850
rect -13910 95650 -13900 95850
rect -14100 95620 -13900 95650
rect -13600 95850 -13400 95880
rect -13600 95650 -13590 95850
rect -13520 95650 -13480 95850
rect -13410 95650 -13400 95850
rect -13600 95620 -13400 95650
rect -13100 95850 -12900 95880
rect -13100 95650 -13090 95850
rect -13020 95650 -12980 95850
rect -12910 95650 -12900 95850
rect -13100 95620 -12900 95650
rect -12600 95850 -12400 95880
rect -12600 95650 -12590 95850
rect -12520 95650 -12480 95850
rect -12410 95650 -12400 95850
rect -12600 95620 -12400 95650
rect -12100 95850 -11900 95880
rect -12100 95650 -12090 95850
rect -12020 95650 -11980 95850
rect -11910 95650 -11900 95850
rect -12100 95620 -11900 95650
rect -11600 95850 -11400 95880
rect -11600 95650 -11590 95850
rect -11520 95650 -11480 95850
rect -11410 95650 -11400 95850
rect -11600 95620 -11400 95650
rect -11100 95850 -10900 95880
rect -11100 95650 -11090 95850
rect -11020 95650 -10980 95850
rect -10910 95650 -10900 95850
rect -11100 95620 -10900 95650
rect -10600 95850 -10400 95880
rect -10600 95650 -10590 95850
rect -10520 95650 -10480 95850
rect -10410 95650 -10400 95850
rect -10600 95620 -10400 95650
rect -10100 95850 -9900 95880
rect -10100 95650 -10090 95850
rect -10020 95650 -9980 95850
rect -9910 95650 -9900 95850
rect -10100 95620 -9900 95650
rect -9600 95850 -9400 95880
rect -9600 95650 -9590 95850
rect -9520 95650 -9480 95850
rect -9410 95650 -9400 95850
rect -9600 95620 -9400 95650
rect -9100 95850 -8900 95880
rect -9100 95650 -9090 95850
rect -9020 95650 -8980 95850
rect -8910 95650 -8900 95850
rect -9100 95620 -8900 95650
rect -8600 95850 -8400 95880
rect -8600 95650 -8590 95850
rect -8520 95650 -8480 95850
rect -8410 95650 -8400 95850
rect -8600 95620 -8400 95650
rect -8100 95850 -7900 95880
rect -8100 95650 -8090 95850
rect -8020 95650 -7980 95850
rect -7910 95650 -7900 95850
rect -8100 95620 -7900 95650
rect -7600 95850 -7400 95880
rect -7600 95650 -7590 95850
rect -7520 95650 -7480 95850
rect -7410 95650 -7400 95850
rect -7600 95620 -7400 95650
rect -7100 95850 -6900 95880
rect -7100 95650 -7090 95850
rect -7020 95650 -6980 95850
rect -6910 95650 -6900 95850
rect -7100 95620 -6900 95650
rect -6600 95850 -6400 95880
rect -6600 95650 -6590 95850
rect -6520 95650 -6480 95850
rect -6410 95650 -6400 95850
rect -6600 95620 -6400 95650
rect -6100 95850 -5900 95880
rect -6100 95650 -6090 95850
rect -6020 95650 -5980 95850
rect -5910 95650 -5900 95850
rect -6100 95620 -5900 95650
rect -5600 95850 -5400 95880
rect -5600 95650 -5590 95850
rect -5520 95650 -5480 95850
rect -5410 95650 -5400 95850
rect -5600 95620 -5400 95650
rect -5100 95850 -4900 95880
rect -5100 95650 -5090 95850
rect -5020 95650 -4980 95850
rect -4910 95650 -4900 95850
rect -5100 95620 -4900 95650
rect -4600 95850 -4400 95880
rect -4600 95650 -4590 95850
rect -4520 95650 -4480 95850
rect -4410 95650 -4400 95850
rect -4600 95620 -4400 95650
rect -4100 95850 -3900 95880
rect -4100 95650 -4090 95850
rect -4020 95650 -3980 95850
rect -3910 95650 -3900 95850
rect -4100 95620 -3900 95650
rect -3600 95850 -3400 95880
rect -3600 95650 -3590 95850
rect -3520 95650 -3480 95850
rect -3410 95650 -3400 95850
rect -3600 95620 -3400 95650
rect -3100 95850 -2900 95880
rect -3100 95650 -3090 95850
rect -3020 95650 -2980 95850
rect -2910 95650 -2900 95850
rect -3100 95620 -2900 95650
rect -2600 95850 -2400 95880
rect -2600 95650 -2590 95850
rect -2520 95650 -2480 95850
rect -2410 95650 -2400 95850
rect -2600 95620 -2400 95650
rect -2100 95850 -1900 95880
rect -2100 95650 -2090 95850
rect -2020 95650 -1980 95850
rect -1910 95650 -1900 95850
rect -2100 95620 -1900 95650
rect -1600 95850 -1400 95880
rect -1600 95650 -1590 95850
rect -1520 95650 -1480 95850
rect -1410 95650 -1400 95850
rect -1600 95620 -1400 95650
rect -1100 95850 -900 95880
rect -1100 95650 -1090 95850
rect -1020 95650 -980 95850
rect -910 95650 -900 95850
rect -1100 95620 -900 95650
rect -600 95850 -400 95880
rect -600 95650 -590 95850
rect -520 95650 -480 95850
rect -410 95650 -400 95850
rect -600 95620 -400 95650
rect -100 95850 100 95880
rect -100 95650 -90 95850
rect -20 95650 20 95850
rect 90 95650 100 95850
rect -100 95620 100 95650
rect 400 95850 600 95880
rect 400 95650 410 95850
rect 480 95650 520 95850
rect 590 95650 600 95850
rect 400 95620 600 95650
rect 900 95850 1100 95880
rect 900 95650 910 95850
rect 980 95650 1020 95850
rect 1090 95650 1100 95850
rect 900 95620 1100 95650
rect 1400 95850 1600 95880
rect 1400 95650 1410 95850
rect 1480 95650 1520 95850
rect 1590 95650 1600 95850
rect 1400 95620 1600 95650
rect 1900 95850 2100 95880
rect 1900 95650 1910 95850
rect 1980 95650 2020 95850
rect 2090 95650 2100 95850
rect 1900 95620 2100 95650
rect 2400 95850 2600 95880
rect 2400 95650 2410 95850
rect 2480 95650 2520 95850
rect 2590 95650 2600 95850
rect 2400 95620 2600 95650
rect 2900 95850 3100 95880
rect 2900 95650 2910 95850
rect 2980 95650 3020 95850
rect 3090 95650 3100 95850
rect 2900 95620 3100 95650
rect 3400 95850 3600 95880
rect 3400 95650 3410 95850
rect 3480 95650 3520 95850
rect 3590 95650 3600 95850
rect 3400 95620 3600 95650
rect 3900 95850 4100 95880
rect 3900 95650 3910 95850
rect 3980 95650 4020 95850
rect 4090 95650 4100 95850
rect 3900 95620 4100 95650
rect 4400 95850 4600 95880
rect 4400 95650 4410 95850
rect 4480 95650 4520 95850
rect 4590 95650 4600 95850
rect 4400 95620 4600 95650
rect 4900 95850 5100 95880
rect 4900 95650 4910 95850
rect 4980 95650 5020 95850
rect 5090 95650 5100 95850
rect 4900 95620 5100 95650
rect 5400 95850 5600 95880
rect 5400 95650 5410 95850
rect 5480 95650 5520 95850
rect 5590 95650 5600 95850
rect 5400 95620 5600 95650
rect 5900 95850 6100 95880
rect 5900 95650 5910 95850
rect 5980 95650 6020 95850
rect 6090 95650 6100 95850
rect 5900 95620 6100 95650
rect 6400 95850 6600 95880
rect 6400 95650 6410 95850
rect 6480 95650 6520 95850
rect 6590 95650 6600 95850
rect 6400 95620 6600 95650
rect 6900 95850 7100 95880
rect 6900 95650 6910 95850
rect 6980 95650 7020 95850
rect 7090 95650 7100 95850
rect 6900 95620 7100 95650
rect 7400 95850 7600 95880
rect 7400 95650 7410 95850
rect 7480 95650 7520 95850
rect 7590 95650 7600 95850
rect 7400 95620 7600 95650
rect 7900 95850 8100 95880
rect 7900 95650 7910 95850
rect 7980 95650 8020 95850
rect 8090 95650 8100 95850
rect 7900 95620 8100 95650
rect 8400 95850 8600 95880
rect 8400 95650 8410 95850
rect 8480 95650 8520 95850
rect 8590 95650 8600 95850
rect 8400 95620 8600 95650
rect 8900 95850 9100 95880
rect 8900 95650 8910 95850
rect 8980 95650 9020 95850
rect 9090 95650 9100 95850
rect 8900 95620 9100 95650
rect 9400 95850 9600 95880
rect 9400 95650 9410 95850
rect 9480 95650 9520 95850
rect 9590 95650 9600 95850
rect 9400 95620 9600 95650
rect 9900 95850 10100 95880
rect 9900 95650 9910 95850
rect 9980 95650 10020 95850
rect 10090 95650 10100 95850
rect 9900 95620 10100 95650
rect 10400 95850 10600 95880
rect 10400 95650 10410 95850
rect 10480 95650 10520 95850
rect 10590 95650 10600 95850
rect 10400 95620 10600 95650
rect 10900 95850 11100 95880
rect 10900 95650 10910 95850
rect 10980 95650 11020 95850
rect 11090 95650 11100 95850
rect 10900 95620 11100 95650
rect 11400 95850 11600 95880
rect 11400 95650 11410 95850
rect 11480 95650 11520 95850
rect 11590 95650 11600 95850
rect 11400 95620 11600 95650
rect 11900 95850 12100 95880
rect 11900 95650 11910 95850
rect 11980 95650 12020 95850
rect 12090 95650 12100 95850
rect 11900 95620 12100 95650
rect 12400 95850 12600 95880
rect 12400 95650 12410 95850
rect 12480 95650 12520 95850
rect 12590 95650 12600 95850
rect 12400 95620 12600 95650
rect 12900 95850 13100 95880
rect 12900 95650 12910 95850
rect 12980 95650 13020 95850
rect 13090 95650 13100 95850
rect 12900 95620 13100 95650
rect 13400 95850 13600 95880
rect 13400 95650 13410 95850
rect 13480 95650 13520 95850
rect 13590 95650 13600 95850
rect 13400 95620 13600 95650
rect 13900 95850 14100 95880
rect 13900 95650 13910 95850
rect 13980 95650 14020 95850
rect 14090 95650 14100 95850
rect 13900 95620 14100 95650
rect 14400 95850 14600 95880
rect 14400 95650 14410 95850
rect 14480 95650 14520 95850
rect 14590 95650 14600 95850
rect 14400 95620 14600 95650
rect 14900 95850 15100 95880
rect 14900 95650 14910 95850
rect 14980 95650 15020 95850
rect 15090 95650 15100 95850
rect 14900 95620 15100 95650
rect 15400 95850 15600 95880
rect 15400 95650 15410 95850
rect 15480 95650 15520 95850
rect 15590 95650 15600 95850
rect 15400 95620 15600 95650
rect 15900 95850 16100 95880
rect 15900 95650 15910 95850
rect 15980 95650 16020 95850
rect 16090 95650 16100 95850
rect 15900 95620 16100 95650
rect 16400 95850 16600 95880
rect 16400 95650 16410 95850
rect 16480 95650 16520 95850
rect 16590 95650 16600 95850
rect 16400 95620 16600 95650
rect 16900 95850 17100 95880
rect 16900 95650 16910 95850
rect 16980 95650 17020 95850
rect 17090 95650 17100 95850
rect 16900 95620 17100 95650
rect 17400 95850 17600 95880
rect 17400 95650 17410 95850
rect 17480 95650 17520 95850
rect 17590 95650 17600 95850
rect 17400 95620 17600 95650
rect 17900 95850 18100 95880
rect 17900 95650 17910 95850
rect 17980 95650 18020 95850
rect 18090 95650 18100 95850
rect 17900 95620 18100 95650
rect 18400 95850 18600 95880
rect 18400 95650 18410 95850
rect 18480 95650 18520 95850
rect 18590 95650 18600 95850
rect 18400 95620 18600 95650
rect 18900 95850 19100 95880
rect 18900 95650 18910 95850
rect 18980 95650 19020 95850
rect 19090 95650 19100 95850
rect 18900 95620 19100 95650
rect 19400 95850 19600 95880
rect 19400 95650 19410 95850
rect 19480 95650 19520 95850
rect 19590 95650 19600 95850
rect 19400 95620 19600 95650
rect 19900 95850 20000 95880
rect 19900 95650 19910 95850
rect 19980 95650 20000 95850
rect 19900 95620 20000 95650
rect -16000 95600 -15880 95620
rect -15620 95600 -15380 95620
rect -15120 95600 -14880 95620
rect -14620 95600 -14380 95620
rect -14120 95600 -13880 95620
rect -13620 95600 -13380 95620
rect -13120 95600 -12880 95620
rect -12620 95600 -12380 95620
rect -12120 95600 -11880 95620
rect -11620 95600 -11380 95620
rect -11120 95600 -10880 95620
rect -10620 95600 -10380 95620
rect -10120 95600 -9880 95620
rect -9620 95600 -9380 95620
rect -9120 95600 -8880 95620
rect -8620 95600 -8380 95620
rect -8120 95600 -7880 95620
rect -7620 95600 -7380 95620
rect -7120 95600 -6880 95620
rect -6620 95600 -6380 95620
rect -6120 95600 -5880 95620
rect -5620 95600 -5380 95620
rect -5120 95600 -4880 95620
rect -4620 95600 -4380 95620
rect -4120 95600 -3880 95620
rect -3620 95600 -3380 95620
rect -3120 95600 -2880 95620
rect -2620 95600 -2380 95620
rect -2120 95600 -1880 95620
rect -1620 95600 -1380 95620
rect -1120 95600 -880 95620
rect -620 95600 -380 95620
rect -120 95600 120 95620
rect 380 95600 620 95620
rect 880 95600 1120 95620
rect 1380 95600 1620 95620
rect 1880 95600 2120 95620
rect 2380 95600 2620 95620
rect 2880 95600 3120 95620
rect 3380 95600 3620 95620
rect 3880 95600 4120 95620
rect 4380 95600 4620 95620
rect 4880 95600 5120 95620
rect 5380 95600 5620 95620
rect 5880 95600 6120 95620
rect 6380 95600 6620 95620
rect 6880 95600 7120 95620
rect 7380 95600 7620 95620
rect 7880 95600 8120 95620
rect 8380 95600 8620 95620
rect 8880 95600 9120 95620
rect 9380 95600 9620 95620
rect 9880 95600 10120 95620
rect 10380 95600 10620 95620
rect 10880 95600 11120 95620
rect 11380 95600 11620 95620
rect 11880 95600 12120 95620
rect 12380 95600 12620 95620
rect 12880 95600 13120 95620
rect 13380 95600 13620 95620
rect 13880 95600 14120 95620
rect 14380 95600 14620 95620
rect 14880 95600 15120 95620
rect 15380 95600 15620 95620
rect 15880 95600 16120 95620
rect 16380 95600 16620 95620
rect 16880 95600 17120 95620
rect 17380 95600 17620 95620
rect 17880 95600 18120 95620
rect 18380 95600 18620 95620
rect 18880 95600 19120 95620
rect 19380 95600 19620 95620
rect 19880 95600 20000 95620
rect -16000 95590 20000 95600
rect -16000 95520 -15850 95590
rect -15650 95520 -15350 95590
rect -15150 95520 -14850 95590
rect -14650 95520 -14350 95590
rect -14150 95520 -13850 95590
rect -13650 95520 -13350 95590
rect -13150 95520 -12850 95590
rect -12650 95520 -12350 95590
rect -12150 95520 -11850 95590
rect -11650 95520 -11350 95590
rect -11150 95520 -10850 95590
rect -10650 95520 -10350 95590
rect -10150 95520 -9850 95590
rect -9650 95520 -9350 95590
rect -9150 95520 -8850 95590
rect -8650 95520 -8350 95590
rect -8150 95520 -7850 95590
rect -7650 95520 -7350 95590
rect -7150 95520 -6850 95590
rect -6650 95520 -6350 95590
rect -6150 95520 -5850 95590
rect -5650 95520 -5350 95590
rect -5150 95520 -4850 95590
rect -4650 95520 -4350 95590
rect -4150 95520 -3850 95590
rect -3650 95520 -3350 95590
rect -3150 95520 -2850 95590
rect -2650 95520 -2350 95590
rect -2150 95520 -1850 95590
rect -1650 95520 -1350 95590
rect -1150 95520 -850 95590
rect -650 95520 -350 95590
rect -150 95520 150 95590
rect 350 95520 650 95590
rect 850 95520 1150 95590
rect 1350 95520 1650 95590
rect 1850 95520 2150 95590
rect 2350 95520 2650 95590
rect 2850 95520 3150 95590
rect 3350 95520 3650 95590
rect 3850 95520 4150 95590
rect 4350 95520 4650 95590
rect 4850 95520 5150 95590
rect 5350 95520 5650 95590
rect 5850 95520 6150 95590
rect 6350 95520 6650 95590
rect 6850 95520 7150 95590
rect 7350 95520 7650 95590
rect 7850 95520 8150 95590
rect 8350 95520 8650 95590
rect 8850 95520 9150 95590
rect 9350 95520 9650 95590
rect 9850 95520 10150 95590
rect 10350 95520 10650 95590
rect 10850 95520 11150 95590
rect 11350 95520 11650 95590
rect 11850 95520 12150 95590
rect 12350 95520 12650 95590
rect 12850 95520 13150 95590
rect 13350 95520 13650 95590
rect 13850 95520 14150 95590
rect 14350 95520 14650 95590
rect 14850 95520 15150 95590
rect 15350 95520 15650 95590
rect 15850 95520 16150 95590
rect 16350 95520 16650 95590
rect 16850 95520 17150 95590
rect 17350 95520 17650 95590
rect 17850 95520 18150 95590
rect 18350 95520 18650 95590
rect 18850 95520 19150 95590
rect 19350 95520 19650 95590
rect 19850 95520 20000 95590
rect -16000 95480 20000 95520
rect -16000 95410 -15850 95480
rect -15650 95410 -15350 95480
rect -15150 95410 -14850 95480
rect -14650 95410 -14350 95480
rect -14150 95410 -13850 95480
rect -13650 95410 -13350 95480
rect -13150 95410 -12850 95480
rect -12650 95410 -12350 95480
rect -12150 95410 -11850 95480
rect -11650 95410 -11350 95480
rect -11150 95410 -10850 95480
rect -10650 95410 -10350 95480
rect -10150 95410 -9850 95480
rect -9650 95410 -9350 95480
rect -9150 95410 -8850 95480
rect -8650 95410 -8350 95480
rect -8150 95410 -7850 95480
rect -7650 95410 -7350 95480
rect -7150 95410 -6850 95480
rect -6650 95410 -6350 95480
rect -6150 95410 -5850 95480
rect -5650 95410 -5350 95480
rect -5150 95410 -4850 95480
rect -4650 95410 -4350 95480
rect -4150 95410 -3850 95480
rect -3650 95410 -3350 95480
rect -3150 95410 -2850 95480
rect -2650 95410 -2350 95480
rect -2150 95410 -1850 95480
rect -1650 95410 -1350 95480
rect -1150 95410 -850 95480
rect -650 95410 -350 95480
rect -150 95410 150 95480
rect 350 95410 650 95480
rect 850 95410 1150 95480
rect 1350 95410 1650 95480
rect 1850 95410 2150 95480
rect 2350 95410 2650 95480
rect 2850 95410 3150 95480
rect 3350 95410 3650 95480
rect 3850 95410 4150 95480
rect 4350 95410 4650 95480
rect 4850 95410 5150 95480
rect 5350 95410 5650 95480
rect 5850 95410 6150 95480
rect 6350 95410 6650 95480
rect 6850 95410 7150 95480
rect 7350 95410 7650 95480
rect 7850 95410 8150 95480
rect 8350 95410 8650 95480
rect 8850 95410 9150 95480
rect 9350 95410 9650 95480
rect 9850 95410 10150 95480
rect 10350 95410 10650 95480
rect 10850 95410 11150 95480
rect 11350 95410 11650 95480
rect 11850 95410 12150 95480
rect 12350 95410 12650 95480
rect 12850 95410 13150 95480
rect 13350 95410 13650 95480
rect 13850 95410 14150 95480
rect 14350 95410 14650 95480
rect 14850 95410 15150 95480
rect 15350 95410 15650 95480
rect 15850 95410 16150 95480
rect 16350 95410 16650 95480
rect 16850 95410 17150 95480
rect 17350 95410 17650 95480
rect 17850 95410 18150 95480
rect 18350 95410 18650 95480
rect 18850 95410 19150 95480
rect 19350 95410 19650 95480
rect 19850 95410 20000 95480
rect -16000 95400 20000 95410
rect -16000 95380 -15880 95400
rect -15620 95380 -15380 95400
rect -15120 95380 -14880 95400
rect -14620 95380 -14380 95400
rect -14120 95380 -13880 95400
rect -13620 95380 -13380 95400
rect -13120 95380 -12880 95400
rect -12620 95380 -12380 95400
rect -12120 95380 -11880 95400
rect -11620 95380 -11380 95400
rect -11120 95380 -10880 95400
rect -10620 95380 -10380 95400
rect -10120 95380 -9880 95400
rect -9620 95380 -9380 95400
rect -9120 95380 -8880 95400
rect -8620 95380 -8380 95400
rect -8120 95380 -7880 95400
rect -7620 95380 -7380 95400
rect -7120 95380 -6880 95400
rect -6620 95380 -6380 95400
rect -6120 95380 -5880 95400
rect -5620 95380 -5380 95400
rect -5120 95380 -4880 95400
rect -4620 95380 -4380 95400
rect -4120 95380 -3880 95400
rect -3620 95380 -3380 95400
rect -3120 95380 -2880 95400
rect -2620 95380 -2380 95400
rect -2120 95380 -1880 95400
rect -1620 95380 -1380 95400
rect -1120 95380 -880 95400
rect -620 95380 -380 95400
rect -120 95380 120 95400
rect 380 95380 620 95400
rect 880 95380 1120 95400
rect 1380 95380 1620 95400
rect 1880 95380 2120 95400
rect 2380 95380 2620 95400
rect 2880 95380 3120 95400
rect 3380 95380 3620 95400
rect 3880 95380 4120 95400
rect 4380 95380 4620 95400
rect 4880 95380 5120 95400
rect 5380 95380 5620 95400
rect 5880 95380 6120 95400
rect 6380 95380 6620 95400
rect 6880 95380 7120 95400
rect 7380 95380 7620 95400
rect 7880 95380 8120 95400
rect 8380 95380 8620 95400
rect 8880 95380 9120 95400
rect 9380 95380 9620 95400
rect 9880 95380 10120 95400
rect 10380 95380 10620 95400
rect 10880 95380 11120 95400
rect 11380 95380 11620 95400
rect 11880 95380 12120 95400
rect 12380 95380 12620 95400
rect 12880 95380 13120 95400
rect 13380 95380 13620 95400
rect 13880 95380 14120 95400
rect 14380 95380 14620 95400
rect 14880 95380 15120 95400
rect 15380 95380 15620 95400
rect 15880 95380 16120 95400
rect 16380 95380 16620 95400
rect 16880 95380 17120 95400
rect 17380 95380 17620 95400
rect 17880 95380 18120 95400
rect 18380 95380 18620 95400
rect 18880 95380 19120 95400
rect 19380 95380 19620 95400
rect 19880 95380 20000 95400
rect -16000 95350 -15900 95380
rect -16000 95150 -15980 95350
rect -15910 95150 -15900 95350
rect -16000 95120 -15900 95150
rect -15600 95350 -15400 95380
rect -15600 95150 -15590 95350
rect -15520 95150 -15480 95350
rect -15410 95150 -15400 95350
rect -15600 95120 -15400 95150
rect -15100 95350 -14900 95380
rect -15100 95150 -15090 95350
rect -15020 95150 -14980 95350
rect -14910 95150 -14900 95350
rect -15100 95120 -14900 95150
rect -14600 95350 -14400 95380
rect -14600 95150 -14590 95350
rect -14520 95150 -14480 95350
rect -14410 95150 -14400 95350
rect -14600 95120 -14400 95150
rect -14100 95350 -13900 95380
rect -14100 95150 -14090 95350
rect -14020 95150 -13980 95350
rect -13910 95150 -13900 95350
rect -14100 95120 -13900 95150
rect -13600 95350 -13400 95380
rect -13600 95150 -13590 95350
rect -13520 95150 -13480 95350
rect -13410 95150 -13400 95350
rect -13600 95120 -13400 95150
rect -13100 95350 -12900 95380
rect -13100 95150 -13090 95350
rect -13020 95150 -12980 95350
rect -12910 95150 -12900 95350
rect -13100 95120 -12900 95150
rect -12600 95350 -12400 95380
rect -12600 95150 -12590 95350
rect -12520 95150 -12480 95350
rect -12410 95150 -12400 95350
rect -12600 95120 -12400 95150
rect -12100 95350 -11900 95380
rect -12100 95150 -12090 95350
rect -12020 95150 -11980 95350
rect -11910 95150 -11900 95350
rect -12100 95120 -11900 95150
rect -11600 95350 -11400 95380
rect -11600 95150 -11590 95350
rect -11520 95150 -11480 95350
rect -11410 95150 -11400 95350
rect -11600 95120 -11400 95150
rect -11100 95350 -10900 95380
rect -11100 95150 -11090 95350
rect -11020 95150 -10980 95350
rect -10910 95150 -10900 95350
rect -11100 95120 -10900 95150
rect -10600 95350 -10400 95380
rect -10600 95150 -10590 95350
rect -10520 95150 -10480 95350
rect -10410 95150 -10400 95350
rect -10600 95120 -10400 95150
rect -10100 95350 -9900 95380
rect -10100 95150 -10090 95350
rect -10020 95150 -9980 95350
rect -9910 95150 -9900 95350
rect -10100 95120 -9900 95150
rect -9600 95350 -9400 95380
rect -9600 95150 -9590 95350
rect -9520 95150 -9480 95350
rect -9410 95150 -9400 95350
rect -9600 95120 -9400 95150
rect -9100 95350 -8900 95380
rect -9100 95150 -9090 95350
rect -9020 95150 -8980 95350
rect -8910 95150 -8900 95350
rect -9100 95120 -8900 95150
rect -8600 95350 -8400 95380
rect -8600 95150 -8590 95350
rect -8520 95150 -8480 95350
rect -8410 95150 -8400 95350
rect -8600 95120 -8400 95150
rect -8100 95350 -7900 95380
rect -8100 95150 -8090 95350
rect -8020 95150 -7980 95350
rect -7910 95150 -7900 95350
rect -8100 95120 -7900 95150
rect -7600 95350 -7400 95380
rect -7600 95150 -7590 95350
rect -7520 95150 -7480 95350
rect -7410 95150 -7400 95350
rect -7600 95120 -7400 95150
rect -7100 95350 -6900 95380
rect -7100 95150 -7090 95350
rect -7020 95150 -6980 95350
rect -6910 95150 -6900 95350
rect -7100 95120 -6900 95150
rect -6600 95350 -6400 95380
rect -6600 95150 -6590 95350
rect -6520 95150 -6480 95350
rect -6410 95150 -6400 95350
rect -6600 95120 -6400 95150
rect -6100 95350 -5900 95380
rect -6100 95150 -6090 95350
rect -6020 95150 -5980 95350
rect -5910 95150 -5900 95350
rect -6100 95120 -5900 95150
rect -5600 95350 -5400 95380
rect -5600 95150 -5590 95350
rect -5520 95150 -5480 95350
rect -5410 95150 -5400 95350
rect -5600 95120 -5400 95150
rect -5100 95350 -4900 95380
rect -5100 95150 -5090 95350
rect -5020 95150 -4980 95350
rect -4910 95150 -4900 95350
rect -5100 95120 -4900 95150
rect -4600 95350 -4400 95380
rect -4600 95150 -4590 95350
rect -4520 95150 -4480 95350
rect -4410 95150 -4400 95350
rect -4600 95120 -4400 95150
rect -4100 95350 -3900 95380
rect -4100 95150 -4090 95350
rect -4020 95150 -3980 95350
rect -3910 95150 -3900 95350
rect -4100 95120 -3900 95150
rect -3600 95350 -3400 95380
rect -3600 95150 -3590 95350
rect -3520 95150 -3480 95350
rect -3410 95150 -3400 95350
rect -3600 95120 -3400 95150
rect -3100 95350 -2900 95380
rect -3100 95150 -3090 95350
rect -3020 95150 -2980 95350
rect -2910 95150 -2900 95350
rect -3100 95120 -2900 95150
rect -2600 95350 -2400 95380
rect -2600 95150 -2590 95350
rect -2520 95150 -2480 95350
rect -2410 95150 -2400 95350
rect -2600 95120 -2400 95150
rect -2100 95350 -1900 95380
rect -2100 95150 -2090 95350
rect -2020 95150 -1980 95350
rect -1910 95150 -1900 95350
rect -2100 95120 -1900 95150
rect -1600 95350 -1400 95380
rect -1600 95150 -1590 95350
rect -1520 95150 -1480 95350
rect -1410 95150 -1400 95350
rect -1600 95120 -1400 95150
rect -1100 95350 -900 95380
rect -1100 95150 -1090 95350
rect -1020 95150 -980 95350
rect -910 95150 -900 95350
rect -1100 95120 -900 95150
rect -600 95350 -400 95380
rect -600 95150 -590 95350
rect -520 95150 -480 95350
rect -410 95150 -400 95350
rect -600 95120 -400 95150
rect -100 95350 100 95380
rect -100 95150 -90 95350
rect -20 95150 20 95350
rect 90 95150 100 95350
rect -100 95120 100 95150
rect 400 95350 600 95380
rect 400 95150 410 95350
rect 480 95150 520 95350
rect 590 95150 600 95350
rect 400 95120 600 95150
rect 900 95350 1100 95380
rect 900 95150 910 95350
rect 980 95150 1020 95350
rect 1090 95150 1100 95350
rect 900 95120 1100 95150
rect 1400 95350 1600 95380
rect 1400 95150 1410 95350
rect 1480 95150 1520 95350
rect 1590 95150 1600 95350
rect 1400 95120 1600 95150
rect 1900 95350 2100 95380
rect 1900 95150 1910 95350
rect 1980 95150 2020 95350
rect 2090 95150 2100 95350
rect 1900 95120 2100 95150
rect 2400 95350 2600 95380
rect 2400 95150 2410 95350
rect 2480 95150 2520 95350
rect 2590 95150 2600 95350
rect 2400 95120 2600 95150
rect 2900 95350 3100 95380
rect 2900 95150 2910 95350
rect 2980 95150 3020 95350
rect 3090 95150 3100 95350
rect 2900 95120 3100 95150
rect 3400 95350 3600 95380
rect 3400 95150 3410 95350
rect 3480 95150 3520 95350
rect 3590 95150 3600 95350
rect 3400 95120 3600 95150
rect 3900 95350 4100 95380
rect 3900 95150 3910 95350
rect 3980 95150 4020 95350
rect 4090 95150 4100 95350
rect 3900 95120 4100 95150
rect 4400 95350 4600 95380
rect 4400 95150 4410 95350
rect 4480 95150 4520 95350
rect 4590 95150 4600 95350
rect 4400 95120 4600 95150
rect 4900 95350 5100 95380
rect 4900 95150 4910 95350
rect 4980 95150 5020 95350
rect 5090 95150 5100 95350
rect 4900 95120 5100 95150
rect 5400 95350 5600 95380
rect 5400 95150 5410 95350
rect 5480 95150 5520 95350
rect 5590 95150 5600 95350
rect 5400 95120 5600 95150
rect 5900 95350 6100 95380
rect 5900 95150 5910 95350
rect 5980 95150 6020 95350
rect 6090 95150 6100 95350
rect 5900 95120 6100 95150
rect 6400 95350 6600 95380
rect 6400 95150 6410 95350
rect 6480 95150 6520 95350
rect 6590 95150 6600 95350
rect 6400 95120 6600 95150
rect 6900 95350 7100 95380
rect 6900 95150 6910 95350
rect 6980 95150 7020 95350
rect 7090 95150 7100 95350
rect 6900 95120 7100 95150
rect 7400 95350 7600 95380
rect 7400 95150 7410 95350
rect 7480 95150 7520 95350
rect 7590 95150 7600 95350
rect 7400 95120 7600 95150
rect 7900 95350 8100 95380
rect 7900 95150 7910 95350
rect 7980 95150 8020 95350
rect 8090 95150 8100 95350
rect 7900 95120 8100 95150
rect 8400 95350 8600 95380
rect 8400 95150 8410 95350
rect 8480 95150 8520 95350
rect 8590 95150 8600 95350
rect 8400 95120 8600 95150
rect 8900 95350 9100 95380
rect 8900 95150 8910 95350
rect 8980 95150 9020 95350
rect 9090 95150 9100 95350
rect 8900 95120 9100 95150
rect 9400 95350 9600 95380
rect 9400 95150 9410 95350
rect 9480 95150 9520 95350
rect 9590 95150 9600 95350
rect 9400 95120 9600 95150
rect 9900 95350 10100 95380
rect 9900 95150 9910 95350
rect 9980 95150 10020 95350
rect 10090 95150 10100 95350
rect 9900 95120 10100 95150
rect 10400 95350 10600 95380
rect 10400 95150 10410 95350
rect 10480 95150 10520 95350
rect 10590 95150 10600 95350
rect 10400 95120 10600 95150
rect 10900 95350 11100 95380
rect 10900 95150 10910 95350
rect 10980 95150 11020 95350
rect 11090 95150 11100 95350
rect 10900 95120 11100 95150
rect 11400 95350 11600 95380
rect 11400 95150 11410 95350
rect 11480 95150 11520 95350
rect 11590 95150 11600 95350
rect 11400 95120 11600 95150
rect 11900 95350 12100 95380
rect 11900 95150 11910 95350
rect 11980 95150 12020 95350
rect 12090 95150 12100 95350
rect 11900 95120 12100 95150
rect 12400 95350 12600 95380
rect 12400 95150 12410 95350
rect 12480 95150 12520 95350
rect 12590 95150 12600 95350
rect 12400 95120 12600 95150
rect 12900 95350 13100 95380
rect 12900 95150 12910 95350
rect 12980 95150 13020 95350
rect 13090 95150 13100 95350
rect 12900 95120 13100 95150
rect 13400 95350 13600 95380
rect 13400 95150 13410 95350
rect 13480 95150 13520 95350
rect 13590 95150 13600 95350
rect 13400 95120 13600 95150
rect 13900 95350 14100 95380
rect 13900 95150 13910 95350
rect 13980 95150 14020 95350
rect 14090 95150 14100 95350
rect 13900 95120 14100 95150
rect 14400 95350 14600 95380
rect 14400 95150 14410 95350
rect 14480 95150 14520 95350
rect 14590 95150 14600 95350
rect 14400 95120 14600 95150
rect 14900 95350 15100 95380
rect 14900 95150 14910 95350
rect 14980 95150 15020 95350
rect 15090 95150 15100 95350
rect 14900 95120 15100 95150
rect 15400 95350 15600 95380
rect 15400 95150 15410 95350
rect 15480 95150 15520 95350
rect 15590 95150 15600 95350
rect 15400 95120 15600 95150
rect 15900 95350 16100 95380
rect 15900 95150 15910 95350
rect 15980 95150 16020 95350
rect 16090 95150 16100 95350
rect 15900 95120 16100 95150
rect 16400 95350 16600 95380
rect 16400 95150 16410 95350
rect 16480 95150 16520 95350
rect 16590 95150 16600 95350
rect 16400 95120 16600 95150
rect 16900 95350 17100 95380
rect 16900 95150 16910 95350
rect 16980 95150 17020 95350
rect 17090 95150 17100 95350
rect 16900 95120 17100 95150
rect 17400 95350 17600 95380
rect 17400 95150 17410 95350
rect 17480 95150 17520 95350
rect 17590 95150 17600 95350
rect 17400 95120 17600 95150
rect 17900 95350 18100 95380
rect 17900 95150 17910 95350
rect 17980 95150 18020 95350
rect 18090 95150 18100 95350
rect 17900 95120 18100 95150
rect 18400 95350 18600 95380
rect 18400 95150 18410 95350
rect 18480 95150 18520 95350
rect 18590 95150 18600 95350
rect 18400 95120 18600 95150
rect 18900 95350 19100 95380
rect 18900 95150 18910 95350
rect 18980 95150 19020 95350
rect 19090 95150 19100 95350
rect 18900 95120 19100 95150
rect 19400 95350 19600 95380
rect 19400 95150 19410 95350
rect 19480 95150 19520 95350
rect 19590 95150 19600 95350
rect 19400 95120 19600 95150
rect 19900 95350 20000 95380
rect 19900 95150 19910 95350
rect 19980 95150 20000 95350
rect 19900 95120 20000 95150
rect -16000 95100 -15880 95120
rect -15620 95100 -15380 95120
rect -15120 95100 -14880 95120
rect -14620 95100 -14380 95120
rect -14120 95100 -13880 95120
rect -13620 95100 -13380 95120
rect -13120 95100 -12880 95120
rect -12620 95100 -12380 95120
rect -12120 95100 -11880 95120
rect -11620 95100 -11380 95120
rect -11120 95100 -10880 95120
rect -10620 95100 -10380 95120
rect -10120 95100 -9880 95120
rect -9620 95100 -9380 95120
rect -9120 95100 -8880 95120
rect -8620 95100 -8380 95120
rect -8120 95100 -7880 95120
rect -7620 95100 -7380 95120
rect -7120 95100 -6880 95120
rect -6620 95100 -6380 95120
rect -6120 95100 -5880 95120
rect -5620 95100 -5380 95120
rect -5120 95100 -4880 95120
rect -4620 95100 -4380 95120
rect -4120 95100 -3880 95120
rect -3620 95100 -3380 95120
rect -3120 95100 -2880 95120
rect -2620 95100 -2380 95120
rect -2120 95100 -1880 95120
rect -1620 95100 -1380 95120
rect -1120 95100 -880 95120
rect -620 95100 -380 95120
rect -120 95100 120 95120
rect 380 95100 620 95120
rect 880 95100 1120 95120
rect 1380 95100 1620 95120
rect 1880 95100 2120 95120
rect 2380 95100 2620 95120
rect 2880 95100 3120 95120
rect 3380 95100 3620 95120
rect 3880 95100 4120 95120
rect 4380 95100 4620 95120
rect 4880 95100 5120 95120
rect 5380 95100 5620 95120
rect 5880 95100 6120 95120
rect 6380 95100 6620 95120
rect 6880 95100 7120 95120
rect 7380 95100 7620 95120
rect 7880 95100 8120 95120
rect 8380 95100 8620 95120
rect 8880 95100 9120 95120
rect 9380 95100 9620 95120
rect 9880 95100 10120 95120
rect 10380 95100 10620 95120
rect 10880 95100 11120 95120
rect 11380 95100 11620 95120
rect 11880 95100 12120 95120
rect 12380 95100 12620 95120
rect 12880 95100 13120 95120
rect 13380 95100 13620 95120
rect 13880 95100 14120 95120
rect 14380 95100 14620 95120
rect 14880 95100 15120 95120
rect 15380 95100 15620 95120
rect 15880 95100 16120 95120
rect 16380 95100 16620 95120
rect 16880 95100 17120 95120
rect 17380 95100 17620 95120
rect 17880 95100 18120 95120
rect 18380 95100 18620 95120
rect 18880 95100 19120 95120
rect 19380 95100 19620 95120
rect 19880 95100 20000 95120
rect -16000 95090 20000 95100
rect -16000 95020 -15850 95090
rect -15650 95020 -15350 95090
rect -15150 95020 -14850 95090
rect -14650 95020 -14350 95090
rect -14150 95020 -13850 95090
rect -13650 95020 -13350 95090
rect -13150 95020 -12850 95090
rect -12650 95020 -12350 95090
rect -12150 95020 -11850 95090
rect -11650 95020 -11350 95090
rect -11150 95020 -10850 95090
rect -10650 95020 -10350 95090
rect -10150 95020 -9850 95090
rect -9650 95020 -9350 95090
rect -9150 95020 -8850 95090
rect -8650 95020 -8350 95090
rect -8150 95020 -7850 95090
rect -7650 95020 -7350 95090
rect -7150 95020 -6850 95090
rect -6650 95020 -6350 95090
rect -6150 95020 -5850 95090
rect -5650 95020 -5350 95090
rect -5150 95020 -4850 95090
rect -4650 95020 -4350 95090
rect -4150 95020 -3850 95090
rect -3650 95020 -3350 95090
rect -3150 95020 -2850 95090
rect -2650 95020 -2350 95090
rect -2150 95020 -1850 95090
rect -1650 95020 -1350 95090
rect -1150 95020 -850 95090
rect -650 95020 -350 95090
rect -150 95020 150 95090
rect 350 95020 650 95090
rect 850 95020 1150 95090
rect 1350 95020 1650 95090
rect 1850 95020 2150 95090
rect 2350 95020 2650 95090
rect 2850 95020 3150 95090
rect 3350 95020 3650 95090
rect 3850 95020 4150 95090
rect 4350 95020 4650 95090
rect 4850 95020 5150 95090
rect 5350 95020 5650 95090
rect 5850 95020 6150 95090
rect 6350 95020 6650 95090
rect 6850 95020 7150 95090
rect 7350 95020 7650 95090
rect 7850 95020 8150 95090
rect 8350 95020 8650 95090
rect 8850 95020 9150 95090
rect 9350 95020 9650 95090
rect 9850 95020 10150 95090
rect 10350 95020 10650 95090
rect 10850 95020 11150 95090
rect 11350 95020 11650 95090
rect 11850 95020 12150 95090
rect 12350 95020 12650 95090
rect 12850 95020 13150 95090
rect 13350 95020 13650 95090
rect 13850 95020 14150 95090
rect 14350 95020 14650 95090
rect 14850 95020 15150 95090
rect 15350 95020 15650 95090
rect 15850 95020 16150 95090
rect 16350 95020 16650 95090
rect 16850 95020 17150 95090
rect 17350 95020 17650 95090
rect 17850 95020 18150 95090
rect 18350 95020 18650 95090
rect 18850 95020 19150 95090
rect 19350 95020 19650 95090
rect 19850 95020 20000 95090
rect -16000 94980 20000 95020
rect -16000 94910 -15850 94980
rect -15650 94910 -15350 94980
rect -15150 94910 -14850 94980
rect -14650 94910 -14350 94980
rect -14150 94910 -13850 94980
rect -13650 94910 -13350 94980
rect -13150 94910 -12850 94980
rect -12650 94910 -12350 94980
rect -12150 94910 -11850 94980
rect -11650 94910 -11350 94980
rect -11150 94910 -10850 94980
rect -10650 94910 -10350 94980
rect -10150 94910 -9850 94980
rect -9650 94910 -9350 94980
rect -9150 94910 -8850 94980
rect -8650 94910 -8350 94980
rect -8150 94910 -7850 94980
rect -7650 94910 -7350 94980
rect -7150 94910 -6850 94980
rect -6650 94910 -6350 94980
rect -6150 94910 -5850 94980
rect -5650 94910 -5350 94980
rect -5150 94910 -4850 94980
rect -4650 94910 -4350 94980
rect -4150 94910 -3850 94980
rect -3650 94910 -3350 94980
rect -3150 94910 -2850 94980
rect -2650 94910 -2350 94980
rect -2150 94910 -1850 94980
rect -1650 94910 -1350 94980
rect -1150 94910 -850 94980
rect -650 94910 -350 94980
rect -150 94910 150 94980
rect 350 94910 650 94980
rect 850 94910 1150 94980
rect 1350 94910 1650 94980
rect 1850 94910 2150 94980
rect 2350 94910 2650 94980
rect 2850 94910 3150 94980
rect 3350 94910 3650 94980
rect 3850 94910 4150 94980
rect 4350 94910 4650 94980
rect 4850 94910 5150 94980
rect 5350 94910 5650 94980
rect 5850 94910 6150 94980
rect 6350 94910 6650 94980
rect 6850 94910 7150 94980
rect 7350 94910 7650 94980
rect 7850 94910 8150 94980
rect 8350 94910 8650 94980
rect 8850 94910 9150 94980
rect 9350 94910 9650 94980
rect 9850 94910 10150 94980
rect 10350 94910 10650 94980
rect 10850 94910 11150 94980
rect 11350 94910 11650 94980
rect 11850 94910 12150 94980
rect 12350 94910 12650 94980
rect 12850 94910 13150 94980
rect 13350 94910 13650 94980
rect 13850 94910 14150 94980
rect 14350 94910 14650 94980
rect 14850 94910 15150 94980
rect 15350 94910 15650 94980
rect 15850 94910 16150 94980
rect 16350 94910 16650 94980
rect 16850 94910 17150 94980
rect 17350 94910 17650 94980
rect 17850 94910 18150 94980
rect 18350 94910 18650 94980
rect 18850 94910 19150 94980
rect 19350 94910 19650 94980
rect 19850 94910 20000 94980
rect -16000 94900 20000 94910
rect -16000 94880 -15880 94900
rect -15620 94880 -15380 94900
rect -15120 94880 -14880 94900
rect -14620 94880 -14380 94900
rect -14120 94880 -13880 94900
rect -13620 94880 -13380 94900
rect -13120 94880 -12880 94900
rect -12620 94880 -12380 94900
rect -12120 94880 -11880 94900
rect -11620 94880 -11380 94900
rect -11120 94880 -10880 94900
rect -10620 94880 -10380 94900
rect -10120 94880 -9880 94900
rect -9620 94880 -9380 94900
rect -9120 94880 -8880 94900
rect -8620 94880 -8380 94900
rect -8120 94880 -7880 94900
rect -7620 94880 -7380 94900
rect -7120 94880 -6880 94900
rect -6620 94880 -6380 94900
rect -6120 94880 -5880 94900
rect -5620 94880 -5380 94900
rect -5120 94880 -4880 94900
rect -4620 94880 -4380 94900
rect -4120 94880 -3880 94900
rect -3620 94880 -3380 94900
rect -3120 94880 -2880 94900
rect -2620 94880 -2380 94900
rect -2120 94880 -1880 94900
rect -1620 94880 -1380 94900
rect -1120 94880 -880 94900
rect -620 94880 -380 94900
rect -120 94880 120 94900
rect 380 94880 620 94900
rect 880 94880 1120 94900
rect 1380 94880 1620 94900
rect 1880 94880 2120 94900
rect 2380 94880 2620 94900
rect 2880 94880 3120 94900
rect 3380 94880 3620 94900
rect 3880 94880 4120 94900
rect 4380 94880 4620 94900
rect 4880 94880 5120 94900
rect 5380 94880 5620 94900
rect 5880 94880 6120 94900
rect 6380 94880 6620 94900
rect 6880 94880 7120 94900
rect 7380 94880 7620 94900
rect 7880 94880 8120 94900
rect 8380 94880 8620 94900
rect 8880 94880 9120 94900
rect 9380 94880 9620 94900
rect 9880 94880 10120 94900
rect 10380 94880 10620 94900
rect 10880 94880 11120 94900
rect 11380 94880 11620 94900
rect 11880 94880 12120 94900
rect 12380 94880 12620 94900
rect 12880 94880 13120 94900
rect 13380 94880 13620 94900
rect 13880 94880 14120 94900
rect 14380 94880 14620 94900
rect 14880 94880 15120 94900
rect 15380 94880 15620 94900
rect 15880 94880 16120 94900
rect 16380 94880 16620 94900
rect 16880 94880 17120 94900
rect 17380 94880 17620 94900
rect 17880 94880 18120 94900
rect 18380 94880 18620 94900
rect 18880 94880 19120 94900
rect 19380 94880 19620 94900
rect 19880 94880 20000 94900
rect -16000 94850 -15900 94880
rect -16000 94650 -15980 94850
rect -15910 94650 -15900 94850
rect -16000 94620 -15900 94650
rect -15600 94850 -15400 94880
rect -15600 94650 -15590 94850
rect -15520 94650 -15480 94850
rect -15410 94650 -15400 94850
rect -15600 94620 -15400 94650
rect -15100 94850 -14900 94880
rect -15100 94650 -15090 94850
rect -15020 94650 -14980 94850
rect -14910 94650 -14900 94850
rect -15100 94620 -14900 94650
rect -14600 94850 -14400 94880
rect -14600 94650 -14590 94850
rect -14520 94650 -14480 94850
rect -14410 94650 -14400 94850
rect -14600 94620 -14400 94650
rect -14100 94850 -13900 94880
rect -14100 94650 -14090 94850
rect -14020 94650 -13980 94850
rect -13910 94650 -13900 94850
rect -14100 94620 -13900 94650
rect -13600 94850 -13400 94880
rect -13600 94650 -13590 94850
rect -13520 94650 -13480 94850
rect -13410 94650 -13400 94850
rect -13600 94620 -13400 94650
rect -13100 94850 -12900 94880
rect -13100 94650 -13090 94850
rect -13020 94650 -12980 94850
rect -12910 94650 -12900 94850
rect -13100 94620 -12900 94650
rect -12600 94850 -12400 94880
rect -12600 94650 -12590 94850
rect -12520 94650 -12480 94850
rect -12410 94650 -12400 94850
rect -12600 94620 -12400 94650
rect -12100 94850 -11900 94880
rect -12100 94650 -12090 94850
rect -12020 94650 -11980 94850
rect -11910 94650 -11900 94850
rect -12100 94620 -11900 94650
rect -11600 94850 -11400 94880
rect -11600 94650 -11590 94850
rect -11520 94650 -11480 94850
rect -11410 94650 -11400 94850
rect -11600 94620 -11400 94650
rect -11100 94850 -10900 94880
rect -11100 94650 -11090 94850
rect -11020 94650 -10980 94850
rect -10910 94650 -10900 94850
rect -11100 94620 -10900 94650
rect -10600 94850 -10400 94880
rect -10600 94650 -10590 94850
rect -10520 94650 -10480 94850
rect -10410 94650 -10400 94850
rect -10600 94620 -10400 94650
rect -10100 94850 -9900 94880
rect -10100 94650 -10090 94850
rect -10020 94650 -9980 94850
rect -9910 94650 -9900 94850
rect -10100 94620 -9900 94650
rect -9600 94850 -9400 94880
rect -9600 94650 -9590 94850
rect -9520 94650 -9480 94850
rect -9410 94650 -9400 94850
rect -9600 94620 -9400 94650
rect -9100 94850 -8900 94880
rect -9100 94650 -9090 94850
rect -9020 94650 -8980 94850
rect -8910 94650 -8900 94850
rect -9100 94620 -8900 94650
rect -8600 94850 -8400 94880
rect -8600 94650 -8590 94850
rect -8520 94650 -8480 94850
rect -8410 94650 -8400 94850
rect -8600 94620 -8400 94650
rect -8100 94850 -7900 94880
rect -8100 94650 -8090 94850
rect -8020 94650 -7980 94850
rect -7910 94650 -7900 94850
rect -8100 94620 -7900 94650
rect -7600 94850 -7400 94880
rect -7600 94650 -7590 94850
rect -7520 94650 -7480 94850
rect -7410 94650 -7400 94850
rect -7600 94620 -7400 94650
rect -7100 94850 -6900 94880
rect -7100 94650 -7090 94850
rect -7020 94650 -6980 94850
rect -6910 94650 -6900 94850
rect -7100 94620 -6900 94650
rect -6600 94850 -6400 94880
rect -6600 94650 -6590 94850
rect -6520 94650 -6480 94850
rect -6410 94650 -6400 94850
rect -6600 94620 -6400 94650
rect -6100 94850 -5900 94880
rect -6100 94650 -6090 94850
rect -6020 94650 -5980 94850
rect -5910 94650 -5900 94850
rect -6100 94620 -5900 94650
rect -5600 94850 -5400 94880
rect -5600 94650 -5590 94850
rect -5520 94650 -5480 94850
rect -5410 94650 -5400 94850
rect -5600 94620 -5400 94650
rect -5100 94850 -4900 94880
rect -5100 94650 -5090 94850
rect -5020 94650 -4980 94850
rect -4910 94650 -4900 94850
rect -5100 94620 -4900 94650
rect -4600 94850 -4400 94880
rect -4600 94650 -4590 94850
rect -4520 94650 -4480 94850
rect -4410 94650 -4400 94850
rect -4600 94620 -4400 94650
rect -4100 94850 -3900 94880
rect -4100 94650 -4090 94850
rect -4020 94650 -3980 94850
rect -3910 94650 -3900 94850
rect -4100 94620 -3900 94650
rect -3600 94850 -3400 94880
rect -3600 94650 -3590 94850
rect -3520 94650 -3480 94850
rect -3410 94650 -3400 94850
rect -3600 94620 -3400 94650
rect -3100 94850 -2900 94880
rect -3100 94650 -3090 94850
rect -3020 94650 -2980 94850
rect -2910 94650 -2900 94850
rect -3100 94620 -2900 94650
rect -2600 94850 -2400 94880
rect -2600 94650 -2590 94850
rect -2520 94650 -2480 94850
rect -2410 94650 -2400 94850
rect -2600 94620 -2400 94650
rect -2100 94850 -1900 94880
rect -2100 94650 -2090 94850
rect -2020 94650 -1980 94850
rect -1910 94650 -1900 94850
rect -2100 94620 -1900 94650
rect -1600 94850 -1400 94880
rect -1600 94650 -1590 94850
rect -1520 94650 -1480 94850
rect -1410 94650 -1400 94850
rect -1600 94620 -1400 94650
rect -1100 94850 -900 94880
rect -1100 94650 -1090 94850
rect -1020 94650 -980 94850
rect -910 94650 -900 94850
rect -1100 94620 -900 94650
rect -600 94850 -400 94880
rect -600 94650 -590 94850
rect -520 94650 -480 94850
rect -410 94650 -400 94850
rect -600 94620 -400 94650
rect -100 94850 100 94880
rect -100 94650 -90 94850
rect -20 94650 20 94850
rect 90 94650 100 94850
rect -100 94620 100 94650
rect 400 94850 600 94880
rect 400 94650 410 94850
rect 480 94650 520 94850
rect 590 94650 600 94850
rect 400 94620 600 94650
rect 900 94850 1100 94880
rect 900 94650 910 94850
rect 980 94650 1020 94850
rect 1090 94650 1100 94850
rect 900 94620 1100 94650
rect 1400 94850 1600 94880
rect 1400 94650 1410 94850
rect 1480 94650 1520 94850
rect 1590 94650 1600 94850
rect 1400 94620 1600 94650
rect 1900 94850 2100 94880
rect 1900 94650 1910 94850
rect 1980 94650 2020 94850
rect 2090 94650 2100 94850
rect 1900 94620 2100 94650
rect 2400 94850 2600 94880
rect 2400 94650 2410 94850
rect 2480 94650 2520 94850
rect 2590 94650 2600 94850
rect 2400 94620 2600 94650
rect 2900 94850 3100 94880
rect 2900 94650 2910 94850
rect 2980 94650 3020 94850
rect 3090 94650 3100 94850
rect 2900 94620 3100 94650
rect 3400 94850 3600 94880
rect 3400 94650 3410 94850
rect 3480 94650 3520 94850
rect 3590 94650 3600 94850
rect 3400 94620 3600 94650
rect 3900 94850 4100 94880
rect 3900 94650 3910 94850
rect 3980 94650 4020 94850
rect 4090 94650 4100 94850
rect 3900 94620 4100 94650
rect 4400 94850 4600 94880
rect 4400 94650 4410 94850
rect 4480 94650 4520 94850
rect 4590 94650 4600 94850
rect 4400 94620 4600 94650
rect 4900 94850 5100 94880
rect 4900 94650 4910 94850
rect 4980 94650 5020 94850
rect 5090 94650 5100 94850
rect 4900 94620 5100 94650
rect 5400 94850 5600 94880
rect 5400 94650 5410 94850
rect 5480 94650 5520 94850
rect 5590 94650 5600 94850
rect 5400 94620 5600 94650
rect 5900 94850 6100 94880
rect 5900 94650 5910 94850
rect 5980 94650 6020 94850
rect 6090 94650 6100 94850
rect 5900 94620 6100 94650
rect 6400 94850 6600 94880
rect 6400 94650 6410 94850
rect 6480 94650 6520 94850
rect 6590 94650 6600 94850
rect 6400 94620 6600 94650
rect 6900 94850 7100 94880
rect 6900 94650 6910 94850
rect 6980 94650 7020 94850
rect 7090 94650 7100 94850
rect 6900 94620 7100 94650
rect 7400 94850 7600 94880
rect 7400 94650 7410 94850
rect 7480 94650 7520 94850
rect 7590 94650 7600 94850
rect 7400 94620 7600 94650
rect 7900 94850 8100 94880
rect 7900 94650 7910 94850
rect 7980 94650 8020 94850
rect 8090 94650 8100 94850
rect 7900 94620 8100 94650
rect 8400 94850 8600 94880
rect 8400 94650 8410 94850
rect 8480 94650 8520 94850
rect 8590 94650 8600 94850
rect 8400 94620 8600 94650
rect 8900 94850 9100 94880
rect 8900 94650 8910 94850
rect 8980 94650 9020 94850
rect 9090 94650 9100 94850
rect 8900 94620 9100 94650
rect 9400 94850 9600 94880
rect 9400 94650 9410 94850
rect 9480 94650 9520 94850
rect 9590 94650 9600 94850
rect 9400 94620 9600 94650
rect 9900 94850 10100 94880
rect 9900 94650 9910 94850
rect 9980 94650 10020 94850
rect 10090 94650 10100 94850
rect 9900 94620 10100 94650
rect 10400 94850 10600 94880
rect 10400 94650 10410 94850
rect 10480 94650 10520 94850
rect 10590 94650 10600 94850
rect 10400 94620 10600 94650
rect 10900 94850 11100 94880
rect 10900 94650 10910 94850
rect 10980 94650 11020 94850
rect 11090 94650 11100 94850
rect 10900 94620 11100 94650
rect 11400 94850 11600 94880
rect 11400 94650 11410 94850
rect 11480 94650 11520 94850
rect 11590 94650 11600 94850
rect 11400 94620 11600 94650
rect 11900 94850 12100 94880
rect 11900 94650 11910 94850
rect 11980 94650 12020 94850
rect 12090 94650 12100 94850
rect 11900 94620 12100 94650
rect 12400 94850 12600 94880
rect 12400 94650 12410 94850
rect 12480 94650 12520 94850
rect 12590 94650 12600 94850
rect 12400 94620 12600 94650
rect 12900 94850 13100 94880
rect 12900 94650 12910 94850
rect 12980 94650 13020 94850
rect 13090 94650 13100 94850
rect 12900 94620 13100 94650
rect 13400 94850 13600 94880
rect 13400 94650 13410 94850
rect 13480 94650 13520 94850
rect 13590 94650 13600 94850
rect 13400 94620 13600 94650
rect 13900 94850 14100 94880
rect 13900 94650 13910 94850
rect 13980 94650 14020 94850
rect 14090 94650 14100 94850
rect 13900 94620 14100 94650
rect 14400 94850 14600 94880
rect 14400 94650 14410 94850
rect 14480 94650 14520 94850
rect 14590 94650 14600 94850
rect 14400 94620 14600 94650
rect 14900 94850 15100 94880
rect 14900 94650 14910 94850
rect 14980 94650 15020 94850
rect 15090 94650 15100 94850
rect 14900 94620 15100 94650
rect 15400 94850 15600 94880
rect 15400 94650 15410 94850
rect 15480 94650 15520 94850
rect 15590 94650 15600 94850
rect 15400 94620 15600 94650
rect 15900 94850 16100 94880
rect 15900 94650 15910 94850
rect 15980 94650 16020 94850
rect 16090 94650 16100 94850
rect 15900 94620 16100 94650
rect 16400 94850 16600 94880
rect 16400 94650 16410 94850
rect 16480 94650 16520 94850
rect 16590 94650 16600 94850
rect 16400 94620 16600 94650
rect 16900 94850 17100 94880
rect 16900 94650 16910 94850
rect 16980 94650 17020 94850
rect 17090 94650 17100 94850
rect 16900 94620 17100 94650
rect 17400 94850 17600 94880
rect 17400 94650 17410 94850
rect 17480 94650 17520 94850
rect 17590 94650 17600 94850
rect 17400 94620 17600 94650
rect 17900 94850 18100 94880
rect 17900 94650 17910 94850
rect 17980 94650 18020 94850
rect 18090 94650 18100 94850
rect 17900 94620 18100 94650
rect 18400 94850 18600 94880
rect 18400 94650 18410 94850
rect 18480 94650 18520 94850
rect 18590 94650 18600 94850
rect 18400 94620 18600 94650
rect 18900 94850 19100 94880
rect 18900 94650 18910 94850
rect 18980 94650 19020 94850
rect 19090 94650 19100 94850
rect 18900 94620 19100 94650
rect 19400 94850 19600 94880
rect 19400 94650 19410 94850
rect 19480 94650 19520 94850
rect 19590 94650 19600 94850
rect 19400 94620 19600 94650
rect 19900 94850 20000 94880
rect 19900 94650 19910 94850
rect 19980 94650 20000 94850
rect 19900 94620 20000 94650
rect -16000 94600 -15880 94620
rect -15620 94600 -15380 94620
rect -15120 94600 -14880 94620
rect -14620 94600 -14380 94620
rect -14120 94600 -13880 94620
rect -13620 94600 -13380 94620
rect -13120 94600 -12880 94620
rect -12620 94600 -12380 94620
rect -12120 94600 -11880 94620
rect -11620 94600 -11380 94620
rect -11120 94600 -10880 94620
rect -10620 94600 -10380 94620
rect -10120 94600 -9880 94620
rect -9620 94600 -9380 94620
rect -9120 94600 -8880 94620
rect -8620 94600 -8380 94620
rect -8120 94600 -7880 94620
rect -7620 94600 -7380 94620
rect -7120 94600 -6880 94620
rect -6620 94600 -6380 94620
rect -6120 94600 -5880 94620
rect -5620 94600 -5380 94620
rect -5120 94600 -4880 94620
rect -4620 94600 -4380 94620
rect -4120 94600 -3880 94620
rect -3620 94600 -3380 94620
rect -3120 94600 -2880 94620
rect -2620 94600 -2380 94620
rect -2120 94600 -1880 94620
rect -1620 94600 -1380 94620
rect -1120 94600 -880 94620
rect -620 94600 -380 94620
rect -120 94600 120 94620
rect 380 94600 620 94620
rect 880 94600 1120 94620
rect 1380 94600 1620 94620
rect 1880 94600 2120 94620
rect 2380 94600 2620 94620
rect 2880 94600 3120 94620
rect 3380 94600 3620 94620
rect 3880 94600 4120 94620
rect 4380 94600 4620 94620
rect 4880 94600 5120 94620
rect 5380 94600 5620 94620
rect 5880 94600 6120 94620
rect 6380 94600 6620 94620
rect 6880 94600 7120 94620
rect 7380 94600 7620 94620
rect 7880 94600 8120 94620
rect 8380 94600 8620 94620
rect 8880 94600 9120 94620
rect 9380 94600 9620 94620
rect 9880 94600 10120 94620
rect 10380 94600 10620 94620
rect 10880 94600 11120 94620
rect 11380 94600 11620 94620
rect 11880 94600 12120 94620
rect 12380 94600 12620 94620
rect 12880 94600 13120 94620
rect 13380 94600 13620 94620
rect 13880 94600 14120 94620
rect 14380 94600 14620 94620
rect 14880 94600 15120 94620
rect 15380 94600 15620 94620
rect 15880 94600 16120 94620
rect 16380 94600 16620 94620
rect 16880 94600 17120 94620
rect 17380 94600 17620 94620
rect 17880 94600 18120 94620
rect 18380 94600 18620 94620
rect 18880 94600 19120 94620
rect 19380 94600 19620 94620
rect 19880 94600 20000 94620
rect -16000 94590 20000 94600
rect -16000 94520 -15850 94590
rect -15650 94520 -15350 94590
rect -15150 94520 -14850 94590
rect -14650 94520 -14350 94590
rect -14150 94520 -13850 94590
rect -13650 94520 -13350 94590
rect -13150 94520 -12850 94590
rect -12650 94520 -12350 94590
rect -12150 94520 -11850 94590
rect -11650 94520 -11350 94590
rect -11150 94520 -10850 94590
rect -10650 94520 -10350 94590
rect -10150 94520 -9850 94590
rect -9650 94520 -9350 94590
rect -9150 94520 -8850 94590
rect -8650 94520 -8350 94590
rect -8150 94520 -7850 94590
rect -7650 94520 -7350 94590
rect -7150 94520 -6850 94590
rect -6650 94520 -6350 94590
rect -6150 94520 -5850 94590
rect -5650 94520 -5350 94590
rect -5150 94520 -4850 94590
rect -4650 94520 -4350 94590
rect -4150 94520 -3850 94590
rect -3650 94520 -3350 94590
rect -3150 94520 -2850 94590
rect -2650 94520 -2350 94590
rect -2150 94520 -1850 94590
rect -1650 94520 -1350 94590
rect -1150 94520 -850 94590
rect -650 94520 -350 94590
rect -150 94520 150 94590
rect 350 94520 650 94590
rect 850 94520 1150 94590
rect 1350 94520 1650 94590
rect 1850 94520 2150 94590
rect 2350 94520 2650 94590
rect 2850 94520 3150 94590
rect 3350 94520 3650 94590
rect 3850 94520 4150 94590
rect 4350 94520 4650 94590
rect 4850 94520 5150 94590
rect 5350 94520 5650 94590
rect 5850 94520 6150 94590
rect 6350 94520 6650 94590
rect 6850 94520 7150 94590
rect 7350 94520 7650 94590
rect 7850 94520 8150 94590
rect 8350 94520 8650 94590
rect 8850 94520 9150 94590
rect 9350 94520 9650 94590
rect 9850 94520 10150 94590
rect 10350 94520 10650 94590
rect 10850 94520 11150 94590
rect 11350 94520 11650 94590
rect 11850 94520 12150 94590
rect 12350 94520 12650 94590
rect 12850 94520 13150 94590
rect 13350 94520 13650 94590
rect 13850 94520 14150 94590
rect 14350 94520 14650 94590
rect 14850 94520 15150 94590
rect 15350 94520 15650 94590
rect 15850 94520 16150 94590
rect 16350 94520 16650 94590
rect 16850 94520 17150 94590
rect 17350 94520 17650 94590
rect 17850 94520 18150 94590
rect 18350 94520 18650 94590
rect 18850 94520 19150 94590
rect 19350 94520 19650 94590
rect 19850 94520 20000 94590
rect -16000 94480 20000 94520
rect -16000 94410 -15850 94480
rect -15650 94410 -15350 94480
rect -15150 94410 -14850 94480
rect -14650 94410 -14350 94480
rect -14150 94410 -13850 94480
rect -13650 94410 -13350 94480
rect -13150 94410 -12850 94480
rect -12650 94410 -12350 94480
rect -12150 94410 -11850 94480
rect -11650 94410 -11350 94480
rect -11150 94410 -10850 94480
rect -10650 94410 -10350 94480
rect -10150 94410 -9850 94480
rect -9650 94410 -9350 94480
rect -9150 94410 -8850 94480
rect -8650 94410 -8350 94480
rect -8150 94410 -7850 94480
rect -7650 94410 -7350 94480
rect -7150 94410 -6850 94480
rect -6650 94410 -6350 94480
rect -6150 94410 -5850 94480
rect -5650 94410 -5350 94480
rect -5150 94410 -4850 94480
rect -4650 94410 -4350 94480
rect -4150 94410 -3850 94480
rect -3650 94410 -3350 94480
rect -3150 94410 -2850 94480
rect -2650 94410 -2350 94480
rect -2150 94410 -1850 94480
rect -1650 94410 -1350 94480
rect -1150 94410 -850 94480
rect -650 94410 -350 94480
rect -150 94410 150 94480
rect 350 94410 650 94480
rect 850 94410 1150 94480
rect 1350 94410 1650 94480
rect 1850 94410 2150 94480
rect 2350 94410 2650 94480
rect 2850 94410 3150 94480
rect 3350 94410 3650 94480
rect 3850 94410 4150 94480
rect 4350 94410 4650 94480
rect 4850 94410 5150 94480
rect 5350 94410 5650 94480
rect 5850 94410 6150 94480
rect 6350 94410 6650 94480
rect 6850 94410 7150 94480
rect 7350 94410 7650 94480
rect 7850 94410 8150 94480
rect 8350 94410 8650 94480
rect 8850 94410 9150 94480
rect 9350 94410 9650 94480
rect 9850 94410 10150 94480
rect 10350 94410 10650 94480
rect 10850 94410 11150 94480
rect 11350 94410 11650 94480
rect 11850 94410 12150 94480
rect 12350 94410 12650 94480
rect 12850 94410 13150 94480
rect 13350 94410 13650 94480
rect 13850 94410 14150 94480
rect 14350 94410 14650 94480
rect 14850 94410 15150 94480
rect 15350 94410 15650 94480
rect 15850 94410 16150 94480
rect 16350 94410 16650 94480
rect 16850 94410 17150 94480
rect 17350 94410 17650 94480
rect 17850 94410 18150 94480
rect 18350 94410 18650 94480
rect 18850 94410 19150 94480
rect 19350 94410 19650 94480
rect 19850 94410 20000 94480
rect -16000 94400 20000 94410
rect -16000 94380 -15880 94400
rect -15620 94380 -15380 94400
rect -15120 94380 -14880 94400
rect -14620 94380 -14380 94400
rect -14120 94380 -13880 94400
rect -13620 94380 -13380 94400
rect -13120 94380 -12880 94400
rect -12620 94380 -12380 94400
rect -12120 94380 -11880 94400
rect -11620 94380 -11380 94400
rect -11120 94380 -10880 94400
rect -10620 94380 -10380 94400
rect -10120 94380 -9880 94400
rect -9620 94380 -9380 94400
rect -9120 94380 -8880 94400
rect -8620 94380 -8380 94400
rect -8120 94380 -7880 94400
rect -7620 94380 -7380 94400
rect -7120 94380 -6880 94400
rect -6620 94380 -6380 94400
rect -6120 94380 -5880 94400
rect -5620 94380 -5380 94400
rect -5120 94380 -4880 94400
rect -4620 94380 -4380 94400
rect -4120 94380 -3880 94400
rect -3620 94380 -3380 94400
rect -3120 94380 -2880 94400
rect -2620 94380 -2380 94400
rect -2120 94380 -1880 94400
rect -1620 94380 -1380 94400
rect -1120 94380 -880 94400
rect -620 94380 -380 94400
rect -120 94380 120 94400
rect 380 94380 620 94400
rect 880 94380 1120 94400
rect 1380 94380 1620 94400
rect 1880 94380 2120 94400
rect 2380 94380 2620 94400
rect 2880 94380 3120 94400
rect 3380 94380 3620 94400
rect 3880 94380 4120 94400
rect 4380 94380 4620 94400
rect 4880 94380 5120 94400
rect 5380 94380 5620 94400
rect 5880 94380 6120 94400
rect 6380 94380 6620 94400
rect 6880 94380 7120 94400
rect 7380 94380 7620 94400
rect 7880 94380 8120 94400
rect 8380 94380 8620 94400
rect 8880 94380 9120 94400
rect 9380 94380 9620 94400
rect 9880 94380 10120 94400
rect 10380 94380 10620 94400
rect 10880 94380 11120 94400
rect 11380 94380 11620 94400
rect 11880 94380 12120 94400
rect 12380 94380 12620 94400
rect 12880 94380 13120 94400
rect 13380 94380 13620 94400
rect 13880 94380 14120 94400
rect 14380 94380 14620 94400
rect 14880 94380 15120 94400
rect 15380 94380 15620 94400
rect 15880 94380 16120 94400
rect 16380 94380 16620 94400
rect 16880 94380 17120 94400
rect 17380 94380 17620 94400
rect 17880 94380 18120 94400
rect 18380 94380 18620 94400
rect 18880 94380 19120 94400
rect 19380 94380 19620 94400
rect 19880 94380 20000 94400
rect -16000 94350 -15900 94380
rect -16000 94150 -15980 94350
rect -15910 94150 -15900 94350
rect -16000 94120 -15900 94150
rect -15600 94350 -15400 94380
rect -15600 94150 -15590 94350
rect -15520 94150 -15480 94350
rect -15410 94150 -15400 94350
rect -15600 94120 -15400 94150
rect -15100 94350 -14900 94380
rect -15100 94150 -15090 94350
rect -15020 94150 -14980 94350
rect -14910 94150 -14900 94350
rect -15100 94120 -14900 94150
rect -14600 94350 -14400 94380
rect -14600 94150 -14590 94350
rect -14520 94150 -14480 94350
rect -14410 94150 -14400 94350
rect -14600 94120 -14400 94150
rect -14100 94350 -13900 94380
rect -14100 94150 -14090 94350
rect -14020 94150 -13980 94350
rect -13910 94150 -13900 94350
rect -14100 94120 -13900 94150
rect -13600 94350 -13400 94380
rect -13600 94150 -13590 94350
rect -13520 94150 -13480 94350
rect -13410 94150 -13400 94350
rect -13600 94120 -13400 94150
rect -13100 94350 -12900 94380
rect -13100 94150 -13090 94350
rect -13020 94150 -12980 94350
rect -12910 94150 -12900 94350
rect -13100 94120 -12900 94150
rect -12600 94350 -12400 94380
rect -12600 94150 -12590 94350
rect -12520 94150 -12480 94350
rect -12410 94150 -12400 94350
rect -12600 94120 -12400 94150
rect -12100 94350 -11900 94380
rect -12100 94150 -12090 94350
rect -12020 94150 -11980 94350
rect -11910 94150 -11900 94350
rect -12100 94120 -11900 94150
rect -11600 94350 -11400 94380
rect -11600 94150 -11590 94350
rect -11520 94150 -11480 94350
rect -11410 94150 -11400 94350
rect -11600 94120 -11400 94150
rect -11100 94350 -10900 94380
rect -11100 94150 -11090 94350
rect -11020 94150 -10980 94350
rect -10910 94150 -10900 94350
rect -11100 94120 -10900 94150
rect -10600 94350 -10400 94380
rect -10600 94150 -10590 94350
rect -10520 94150 -10480 94350
rect -10410 94150 -10400 94350
rect -10600 94120 -10400 94150
rect -10100 94350 -9900 94380
rect -10100 94150 -10090 94350
rect -10020 94150 -9980 94350
rect -9910 94150 -9900 94350
rect -10100 94120 -9900 94150
rect -9600 94350 -9400 94380
rect -9600 94150 -9590 94350
rect -9520 94150 -9480 94350
rect -9410 94150 -9400 94350
rect -9600 94120 -9400 94150
rect -9100 94350 -8900 94380
rect -9100 94150 -9090 94350
rect -9020 94150 -8980 94350
rect -8910 94150 -8900 94350
rect -9100 94120 -8900 94150
rect -8600 94350 -8400 94380
rect -8600 94150 -8590 94350
rect -8520 94150 -8480 94350
rect -8410 94150 -8400 94350
rect -8600 94120 -8400 94150
rect -8100 94350 -7900 94380
rect -8100 94150 -8090 94350
rect -8020 94150 -7980 94350
rect -7910 94150 -7900 94350
rect -8100 94120 -7900 94150
rect -7600 94350 -7400 94380
rect -7600 94150 -7590 94350
rect -7520 94150 -7480 94350
rect -7410 94150 -7400 94350
rect -7600 94120 -7400 94150
rect -7100 94350 -6900 94380
rect -7100 94150 -7090 94350
rect -7020 94150 -6980 94350
rect -6910 94150 -6900 94350
rect -7100 94120 -6900 94150
rect -6600 94350 -6400 94380
rect -6600 94150 -6590 94350
rect -6520 94150 -6480 94350
rect -6410 94150 -6400 94350
rect -6600 94120 -6400 94150
rect -6100 94350 -5900 94380
rect -6100 94150 -6090 94350
rect -6020 94150 -5980 94350
rect -5910 94150 -5900 94350
rect -6100 94120 -5900 94150
rect -5600 94350 -5400 94380
rect -5600 94150 -5590 94350
rect -5520 94150 -5480 94350
rect -5410 94150 -5400 94350
rect -5600 94120 -5400 94150
rect -5100 94350 -4900 94380
rect -5100 94150 -5090 94350
rect -5020 94150 -4980 94350
rect -4910 94150 -4900 94350
rect -5100 94120 -4900 94150
rect -4600 94350 -4400 94380
rect -4600 94150 -4590 94350
rect -4520 94150 -4480 94350
rect -4410 94150 -4400 94350
rect -4600 94120 -4400 94150
rect -4100 94350 -3900 94380
rect -4100 94150 -4090 94350
rect -4020 94150 -3980 94350
rect -3910 94150 -3900 94350
rect -4100 94120 -3900 94150
rect -3600 94350 -3400 94380
rect -3600 94150 -3590 94350
rect -3520 94150 -3480 94350
rect -3410 94150 -3400 94350
rect -3600 94120 -3400 94150
rect -3100 94350 -2900 94380
rect -3100 94150 -3090 94350
rect -3020 94150 -2980 94350
rect -2910 94150 -2900 94350
rect -3100 94120 -2900 94150
rect -2600 94350 -2400 94380
rect -2600 94150 -2590 94350
rect -2520 94150 -2480 94350
rect -2410 94150 -2400 94350
rect -2600 94120 -2400 94150
rect -2100 94350 -1900 94380
rect -2100 94150 -2090 94350
rect -2020 94150 -1980 94350
rect -1910 94150 -1900 94350
rect -2100 94120 -1900 94150
rect -1600 94350 -1400 94380
rect -1600 94150 -1590 94350
rect -1520 94150 -1480 94350
rect -1410 94150 -1400 94350
rect -1600 94120 -1400 94150
rect -1100 94350 -900 94380
rect -1100 94150 -1090 94350
rect -1020 94150 -980 94350
rect -910 94150 -900 94350
rect -1100 94120 -900 94150
rect -600 94350 -400 94380
rect -600 94150 -590 94350
rect -520 94150 -480 94350
rect -410 94150 -400 94350
rect -600 94120 -400 94150
rect -100 94350 100 94380
rect -100 94150 -90 94350
rect -20 94150 20 94350
rect 90 94150 100 94350
rect -100 94120 100 94150
rect 400 94350 600 94380
rect 400 94150 410 94350
rect 480 94150 520 94350
rect 590 94150 600 94350
rect 400 94120 600 94150
rect 900 94350 1100 94380
rect 900 94150 910 94350
rect 980 94150 1020 94350
rect 1090 94150 1100 94350
rect 900 94120 1100 94150
rect 1400 94350 1600 94380
rect 1400 94150 1410 94350
rect 1480 94150 1520 94350
rect 1590 94150 1600 94350
rect 1400 94120 1600 94150
rect 1900 94350 2100 94380
rect 1900 94150 1910 94350
rect 1980 94150 2020 94350
rect 2090 94150 2100 94350
rect 1900 94120 2100 94150
rect 2400 94350 2600 94380
rect 2400 94150 2410 94350
rect 2480 94150 2520 94350
rect 2590 94150 2600 94350
rect 2400 94120 2600 94150
rect 2900 94350 3100 94380
rect 2900 94150 2910 94350
rect 2980 94150 3020 94350
rect 3090 94150 3100 94350
rect 2900 94120 3100 94150
rect 3400 94350 3600 94380
rect 3400 94150 3410 94350
rect 3480 94150 3520 94350
rect 3590 94150 3600 94350
rect 3400 94120 3600 94150
rect 3900 94350 4100 94380
rect 3900 94150 3910 94350
rect 3980 94150 4020 94350
rect 4090 94150 4100 94350
rect 3900 94120 4100 94150
rect 4400 94350 4600 94380
rect 4400 94150 4410 94350
rect 4480 94150 4520 94350
rect 4590 94150 4600 94350
rect 4400 94120 4600 94150
rect 4900 94350 5100 94380
rect 4900 94150 4910 94350
rect 4980 94150 5020 94350
rect 5090 94150 5100 94350
rect 4900 94120 5100 94150
rect 5400 94350 5600 94380
rect 5400 94150 5410 94350
rect 5480 94150 5520 94350
rect 5590 94150 5600 94350
rect 5400 94120 5600 94150
rect 5900 94350 6100 94380
rect 5900 94150 5910 94350
rect 5980 94150 6020 94350
rect 6090 94150 6100 94350
rect 5900 94120 6100 94150
rect 6400 94350 6600 94380
rect 6400 94150 6410 94350
rect 6480 94150 6520 94350
rect 6590 94150 6600 94350
rect 6400 94120 6600 94150
rect 6900 94350 7100 94380
rect 6900 94150 6910 94350
rect 6980 94150 7020 94350
rect 7090 94150 7100 94350
rect 6900 94120 7100 94150
rect 7400 94350 7600 94380
rect 7400 94150 7410 94350
rect 7480 94150 7520 94350
rect 7590 94150 7600 94350
rect 7400 94120 7600 94150
rect 7900 94350 8100 94380
rect 7900 94150 7910 94350
rect 7980 94150 8020 94350
rect 8090 94150 8100 94350
rect 7900 94120 8100 94150
rect 8400 94350 8600 94380
rect 8400 94150 8410 94350
rect 8480 94150 8520 94350
rect 8590 94150 8600 94350
rect 8400 94120 8600 94150
rect 8900 94350 9100 94380
rect 8900 94150 8910 94350
rect 8980 94150 9020 94350
rect 9090 94150 9100 94350
rect 8900 94120 9100 94150
rect 9400 94350 9600 94380
rect 9400 94150 9410 94350
rect 9480 94150 9520 94350
rect 9590 94150 9600 94350
rect 9400 94120 9600 94150
rect 9900 94350 10100 94380
rect 9900 94150 9910 94350
rect 9980 94150 10020 94350
rect 10090 94150 10100 94350
rect 9900 94120 10100 94150
rect 10400 94350 10600 94380
rect 10400 94150 10410 94350
rect 10480 94150 10520 94350
rect 10590 94150 10600 94350
rect 10400 94120 10600 94150
rect 10900 94350 11100 94380
rect 10900 94150 10910 94350
rect 10980 94150 11020 94350
rect 11090 94150 11100 94350
rect 10900 94120 11100 94150
rect 11400 94350 11600 94380
rect 11400 94150 11410 94350
rect 11480 94150 11520 94350
rect 11590 94150 11600 94350
rect 11400 94120 11600 94150
rect 11900 94350 12100 94380
rect 11900 94150 11910 94350
rect 11980 94150 12020 94350
rect 12090 94150 12100 94350
rect 11900 94120 12100 94150
rect 12400 94350 12600 94380
rect 12400 94150 12410 94350
rect 12480 94150 12520 94350
rect 12590 94150 12600 94350
rect 12400 94120 12600 94150
rect 12900 94350 13100 94380
rect 12900 94150 12910 94350
rect 12980 94150 13020 94350
rect 13090 94150 13100 94350
rect 12900 94120 13100 94150
rect 13400 94350 13600 94380
rect 13400 94150 13410 94350
rect 13480 94150 13520 94350
rect 13590 94150 13600 94350
rect 13400 94120 13600 94150
rect 13900 94350 14100 94380
rect 13900 94150 13910 94350
rect 13980 94150 14020 94350
rect 14090 94150 14100 94350
rect 13900 94120 14100 94150
rect 14400 94350 14600 94380
rect 14400 94150 14410 94350
rect 14480 94150 14520 94350
rect 14590 94150 14600 94350
rect 14400 94120 14600 94150
rect 14900 94350 15100 94380
rect 14900 94150 14910 94350
rect 14980 94150 15020 94350
rect 15090 94150 15100 94350
rect 14900 94120 15100 94150
rect 15400 94350 15600 94380
rect 15400 94150 15410 94350
rect 15480 94150 15520 94350
rect 15590 94150 15600 94350
rect 15400 94120 15600 94150
rect 15900 94350 16100 94380
rect 15900 94150 15910 94350
rect 15980 94150 16020 94350
rect 16090 94150 16100 94350
rect 15900 94120 16100 94150
rect 16400 94350 16600 94380
rect 16400 94150 16410 94350
rect 16480 94150 16520 94350
rect 16590 94150 16600 94350
rect 16400 94120 16600 94150
rect 16900 94350 17100 94380
rect 16900 94150 16910 94350
rect 16980 94150 17020 94350
rect 17090 94150 17100 94350
rect 16900 94120 17100 94150
rect 17400 94350 17600 94380
rect 17400 94150 17410 94350
rect 17480 94150 17520 94350
rect 17590 94150 17600 94350
rect 17400 94120 17600 94150
rect 17900 94350 18100 94380
rect 17900 94150 17910 94350
rect 17980 94150 18020 94350
rect 18090 94150 18100 94350
rect 17900 94120 18100 94150
rect 18400 94350 18600 94380
rect 18400 94150 18410 94350
rect 18480 94150 18520 94350
rect 18590 94150 18600 94350
rect 18400 94120 18600 94150
rect 18900 94350 19100 94380
rect 18900 94150 18910 94350
rect 18980 94150 19020 94350
rect 19090 94150 19100 94350
rect 18900 94120 19100 94150
rect 19400 94350 19600 94380
rect 19400 94150 19410 94350
rect 19480 94150 19520 94350
rect 19590 94150 19600 94350
rect 19400 94120 19600 94150
rect 19900 94350 20000 94380
rect 19900 94150 19910 94350
rect 19980 94150 20000 94350
rect 19900 94120 20000 94150
rect -16000 94100 -15880 94120
rect -15620 94100 -15380 94120
rect -15120 94100 -14880 94120
rect -14620 94100 -14380 94120
rect -14120 94100 -13880 94120
rect -13620 94100 -13380 94120
rect -13120 94100 -12880 94120
rect -12620 94100 -12380 94120
rect -12120 94100 -11880 94120
rect -11620 94100 -11380 94120
rect -11120 94100 -10880 94120
rect -10620 94100 -10380 94120
rect -10120 94100 -9880 94120
rect -9620 94100 -9380 94120
rect -9120 94100 -8880 94120
rect -8620 94100 -8380 94120
rect -8120 94100 -7880 94120
rect -7620 94100 -7380 94120
rect -7120 94100 -6880 94120
rect -6620 94100 -6380 94120
rect -6120 94100 -5880 94120
rect -5620 94100 -5380 94120
rect -5120 94100 -4880 94120
rect -4620 94100 -4380 94120
rect -4120 94100 -3880 94120
rect -3620 94100 -3380 94120
rect -3120 94100 -2880 94120
rect -2620 94100 -2380 94120
rect -2120 94100 -1880 94120
rect -1620 94100 -1380 94120
rect -1120 94100 -880 94120
rect -620 94100 -380 94120
rect -120 94100 120 94120
rect 380 94100 620 94120
rect 880 94100 1120 94120
rect 1380 94100 1620 94120
rect 1880 94100 2120 94120
rect 2380 94100 2620 94120
rect 2880 94100 3120 94120
rect 3380 94100 3620 94120
rect 3880 94100 4120 94120
rect 4380 94100 4620 94120
rect 4880 94100 5120 94120
rect 5380 94100 5620 94120
rect 5880 94100 6120 94120
rect 6380 94100 6620 94120
rect 6880 94100 7120 94120
rect 7380 94100 7620 94120
rect 7880 94100 8120 94120
rect 8380 94100 8620 94120
rect 8880 94100 9120 94120
rect 9380 94100 9620 94120
rect 9880 94100 10120 94120
rect 10380 94100 10620 94120
rect 10880 94100 11120 94120
rect 11380 94100 11620 94120
rect 11880 94100 12120 94120
rect 12380 94100 12620 94120
rect 12880 94100 13120 94120
rect 13380 94100 13620 94120
rect 13880 94100 14120 94120
rect 14380 94100 14620 94120
rect 14880 94100 15120 94120
rect 15380 94100 15620 94120
rect 15880 94100 16120 94120
rect 16380 94100 16620 94120
rect 16880 94100 17120 94120
rect 17380 94100 17620 94120
rect 17880 94100 18120 94120
rect 18380 94100 18620 94120
rect 18880 94100 19120 94120
rect 19380 94100 19620 94120
rect 19880 94100 20000 94120
rect -16000 94090 20000 94100
rect -16000 94020 -15850 94090
rect -15650 94020 -15350 94090
rect -15150 94020 -14850 94090
rect -14650 94020 -14350 94090
rect -14150 94020 -13850 94090
rect -13650 94020 -13350 94090
rect -13150 94020 -12850 94090
rect -12650 94020 -12350 94090
rect -12150 94020 -11850 94090
rect -11650 94020 -11350 94090
rect -11150 94020 -10850 94090
rect -10650 94020 -10350 94090
rect -10150 94020 -9850 94090
rect -9650 94020 -9350 94090
rect -9150 94020 -8850 94090
rect -8650 94020 -8350 94090
rect -8150 94020 -7850 94090
rect -7650 94020 -7350 94090
rect -7150 94020 -6850 94090
rect -6650 94020 -6350 94090
rect -6150 94020 -5850 94090
rect -5650 94020 -5350 94090
rect -5150 94020 -4850 94090
rect -4650 94020 -4350 94090
rect -4150 94020 -3850 94090
rect -3650 94020 -3350 94090
rect -3150 94020 -2850 94090
rect -2650 94020 -2350 94090
rect -2150 94020 -1850 94090
rect -1650 94020 -1350 94090
rect -1150 94020 -850 94090
rect -650 94020 -350 94090
rect -150 94020 150 94090
rect 350 94020 650 94090
rect 850 94020 1150 94090
rect 1350 94020 1650 94090
rect 1850 94020 2150 94090
rect 2350 94020 2650 94090
rect 2850 94020 3150 94090
rect 3350 94020 3650 94090
rect 3850 94020 4150 94090
rect 4350 94020 4650 94090
rect 4850 94020 5150 94090
rect 5350 94020 5650 94090
rect 5850 94020 6150 94090
rect 6350 94020 6650 94090
rect 6850 94020 7150 94090
rect 7350 94020 7650 94090
rect 7850 94020 8150 94090
rect 8350 94020 8650 94090
rect 8850 94020 9150 94090
rect 9350 94020 9650 94090
rect 9850 94020 10150 94090
rect 10350 94020 10650 94090
rect 10850 94020 11150 94090
rect 11350 94020 11650 94090
rect 11850 94020 12150 94090
rect 12350 94020 12650 94090
rect 12850 94020 13150 94090
rect 13350 94020 13650 94090
rect 13850 94020 14150 94090
rect 14350 94020 14650 94090
rect 14850 94020 15150 94090
rect 15350 94020 15650 94090
rect 15850 94020 16150 94090
rect 16350 94020 16650 94090
rect 16850 94020 17150 94090
rect 17350 94020 17650 94090
rect 17850 94020 18150 94090
rect 18350 94020 18650 94090
rect 18850 94020 19150 94090
rect 19350 94020 19650 94090
rect 19850 94020 20000 94090
rect -16000 94000 20000 94020
rect -16000 93980 -12000 94000
rect -16000 93910 -15850 93980
rect -15650 93910 -15350 93980
rect -15150 93910 -14850 93980
rect -14650 93910 -14350 93980
rect -14150 93910 -13850 93980
rect -13650 93910 -13350 93980
rect -13150 93910 -12850 93980
rect -12650 93910 -12350 93980
rect -12150 93910 -12000 93980
rect -16000 93900 -12000 93910
rect -16000 93880 -15880 93900
rect -15620 93880 -15380 93900
rect -15120 93880 -14880 93900
rect -14620 93880 -14380 93900
rect -14120 93880 -13880 93900
rect -13620 93880 -13380 93900
rect -13120 93880 -12880 93900
rect -12620 93880 -12380 93900
rect -12120 93880 -12000 93900
rect -16000 93850 -15900 93880
rect -16000 93650 -15980 93850
rect -15910 93650 -15900 93850
rect -16000 93620 -15900 93650
rect -15600 93850 -15400 93880
rect -15600 93650 -15590 93850
rect -15520 93650 -15480 93850
rect -15410 93650 -15400 93850
rect -15600 93620 -15400 93650
rect -15100 93850 -14900 93880
rect -15100 93650 -15090 93850
rect -15020 93650 -14980 93850
rect -14910 93650 -14900 93850
rect -15100 93620 -14900 93650
rect -14600 93850 -14400 93880
rect -14600 93650 -14590 93850
rect -14520 93650 -14480 93850
rect -14410 93650 -14400 93850
rect -14600 93620 -14400 93650
rect -14100 93850 -13900 93880
rect -14100 93650 -14090 93850
rect -14020 93650 -13980 93850
rect -13910 93650 -13900 93850
rect -14100 93620 -13900 93650
rect -13600 93850 -13400 93880
rect -13600 93650 -13590 93850
rect -13520 93650 -13480 93850
rect -13410 93650 -13400 93850
rect -13600 93620 -13400 93650
rect -13100 93850 -12900 93880
rect -13100 93650 -13090 93850
rect -13020 93650 -12980 93850
rect -12910 93650 -12900 93850
rect -13100 93620 -12900 93650
rect -12600 93850 -12400 93880
rect -12600 93650 -12590 93850
rect -12520 93650 -12480 93850
rect -12410 93650 -12400 93850
rect -12600 93620 -12400 93650
rect -12100 93850 -12000 93880
rect -12100 93650 -12090 93850
rect -12020 93650 -12000 93850
rect -12100 93620 -12000 93650
rect -16000 93600 -15880 93620
rect -15620 93600 -15380 93620
rect -15120 93600 -14880 93620
rect -14620 93600 -14380 93620
rect -14120 93600 -13880 93620
rect -13620 93600 -13380 93620
rect -13120 93600 -12880 93620
rect -12620 93600 -12380 93620
rect -12120 93600 -12000 93620
rect -16000 93590 -12000 93600
rect -16000 93520 -15850 93590
rect -15650 93520 -15350 93590
rect -15150 93520 -14850 93590
rect -14650 93520 -14350 93590
rect -14150 93520 -13850 93590
rect -13650 93520 -13350 93590
rect -13150 93520 -12850 93590
rect -12650 93520 -12350 93590
rect -12150 93520 -12000 93590
rect -16000 93480 -12000 93520
rect -16000 93410 -15850 93480
rect -15650 93410 -15350 93480
rect -15150 93410 -14850 93480
rect -14650 93410 -14350 93480
rect -14150 93410 -13850 93480
rect -13650 93410 -13350 93480
rect -13150 93410 -12850 93480
rect -12650 93410 -12350 93480
rect -12150 93410 -12000 93480
rect -16000 93400 -12000 93410
rect -16000 93380 -15880 93400
rect -15620 93380 -15380 93400
rect -15120 93380 -14880 93400
rect -14620 93380 -14380 93400
rect -14120 93380 -13880 93400
rect -13620 93380 -13380 93400
rect -13120 93380 -12880 93400
rect -12620 93380 -12380 93400
rect -12120 93380 -12000 93400
rect -16000 93350 -15900 93380
rect -16000 93150 -15980 93350
rect -15910 93150 -15900 93350
rect -16000 93120 -15900 93150
rect -15600 93350 -15400 93380
rect -15600 93150 -15590 93350
rect -15520 93150 -15480 93350
rect -15410 93150 -15400 93350
rect -15600 93120 -15400 93150
rect -15100 93350 -14900 93380
rect -15100 93150 -15090 93350
rect -15020 93150 -14980 93350
rect -14910 93150 -14900 93350
rect -15100 93120 -14900 93150
rect -14600 93350 -14400 93380
rect -14600 93150 -14590 93350
rect -14520 93150 -14480 93350
rect -14410 93150 -14400 93350
rect -14600 93120 -14400 93150
rect -14100 93350 -13900 93380
rect -14100 93150 -14090 93350
rect -14020 93150 -13980 93350
rect -13910 93150 -13900 93350
rect -14100 93120 -13900 93150
rect -13600 93350 -13400 93380
rect -13600 93150 -13590 93350
rect -13520 93150 -13480 93350
rect -13410 93150 -13400 93350
rect -13600 93120 -13400 93150
rect -13100 93350 -12900 93380
rect -13100 93150 -13090 93350
rect -13020 93150 -12980 93350
rect -12910 93150 -12900 93350
rect -13100 93120 -12900 93150
rect -12600 93350 -12400 93380
rect -12600 93150 -12590 93350
rect -12520 93150 -12480 93350
rect -12410 93150 -12400 93350
rect -12600 93120 -12400 93150
rect -12100 93350 -12000 93380
rect -12100 93150 -12090 93350
rect -12020 93150 -12000 93350
rect -12100 93120 -12000 93150
rect -16000 93100 -15880 93120
rect -15620 93100 -15380 93120
rect -15120 93100 -14880 93120
rect -14620 93100 -14380 93120
rect -14120 93100 -13880 93120
rect -13620 93100 -13380 93120
rect -13120 93100 -12880 93120
rect -12620 93100 -12380 93120
rect -12120 93100 -12000 93120
rect -16000 93090 -12000 93100
rect -16000 93020 -15850 93090
rect -15650 93020 -15350 93090
rect -15150 93020 -14850 93090
rect -14650 93020 -14350 93090
rect -14150 93020 -13850 93090
rect -13650 93020 -13350 93090
rect -13150 93020 -12850 93090
rect -12650 93020 -12350 93090
rect -12150 93020 -12000 93090
rect -16000 92980 -12000 93020
rect -16000 92910 -15850 92980
rect -15650 92910 -15350 92980
rect -15150 92910 -14850 92980
rect -14650 92910 -14350 92980
rect -14150 92910 -13850 92980
rect -13650 92910 -13350 92980
rect -13150 92910 -12850 92980
rect -12650 92910 -12350 92980
rect -12150 92910 -12000 92980
rect -16000 92900 -12000 92910
rect -16000 92880 -15880 92900
rect -15620 92880 -15380 92900
rect -15120 92880 -14880 92900
rect -14620 92880 -14380 92900
rect -14120 92880 -13880 92900
rect -13620 92880 -13380 92900
rect -13120 92880 -12880 92900
rect -12620 92880 -12380 92900
rect -12120 92880 -12000 92900
rect -16000 92850 -15900 92880
rect -16000 92650 -15980 92850
rect -15910 92650 -15900 92850
rect -16000 92620 -15900 92650
rect -15600 92850 -15400 92880
rect -15600 92650 -15590 92850
rect -15520 92650 -15480 92850
rect -15410 92650 -15400 92850
rect -15600 92620 -15400 92650
rect -15100 92850 -14900 92880
rect -15100 92650 -15090 92850
rect -15020 92650 -14980 92850
rect -14910 92650 -14900 92850
rect -15100 92620 -14900 92650
rect -14600 92850 -14400 92880
rect -14600 92650 -14590 92850
rect -14520 92650 -14480 92850
rect -14410 92650 -14400 92850
rect -14600 92620 -14400 92650
rect -14100 92850 -13900 92880
rect -14100 92650 -14090 92850
rect -14020 92650 -13980 92850
rect -13910 92650 -13900 92850
rect -14100 92620 -13900 92650
rect -13600 92850 -13400 92880
rect -13600 92650 -13590 92850
rect -13520 92650 -13480 92850
rect -13410 92650 -13400 92850
rect -13600 92620 -13400 92650
rect -13100 92850 -12900 92880
rect -13100 92650 -13090 92850
rect -13020 92650 -12980 92850
rect -12910 92650 -12900 92850
rect -13100 92620 -12900 92650
rect -12600 92850 -12400 92880
rect -12600 92650 -12590 92850
rect -12520 92650 -12480 92850
rect -12410 92650 -12400 92850
rect -12600 92620 -12400 92650
rect -12100 92850 -12000 92880
rect -12100 92650 -12090 92850
rect -12020 92650 -12000 92850
rect -12100 92620 -12000 92650
rect -16000 92600 -15880 92620
rect -15620 92600 -15380 92620
rect -15120 92600 -14880 92620
rect -14620 92600 -14380 92620
rect -14120 92600 -13880 92620
rect -13620 92600 -13380 92620
rect -13120 92600 -12880 92620
rect -12620 92600 -12380 92620
rect -12120 92600 -12000 92620
rect -16000 92590 -12000 92600
rect -16000 92520 -15850 92590
rect -15650 92520 -15350 92590
rect -15150 92520 -14850 92590
rect -14650 92520 -14350 92590
rect -14150 92520 -13850 92590
rect -13650 92520 -13350 92590
rect -13150 92520 -12850 92590
rect -12650 92520 -12350 92590
rect -12150 92520 -12000 92590
rect -16000 92480 -12000 92520
rect -16000 92410 -15850 92480
rect -15650 92410 -15350 92480
rect -15150 92410 -14850 92480
rect -14650 92410 -14350 92480
rect -14150 92410 -13850 92480
rect -13650 92410 -13350 92480
rect -13150 92410 -12850 92480
rect -12650 92410 -12350 92480
rect -12150 92410 -12000 92480
rect -16000 92400 -12000 92410
rect -16000 92380 -15880 92400
rect -15620 92380 -15380 92400
rect -15120 92380 -14880 92400
rect -14620 92380 -14380 92400
rect -14120 92380 -13880 92400
rect -13620 92380 -13380 92400
rect -13120 92380 -12880 92400
rect -12620 92380 -12380 92400
rect -12120 92380 -12000 92400
rect -16000 92350 -15900 92380
rect -16000 92150 -15980 92350
rect -15910 92150 -15900 92350
rect -16000 92120 -15900 92150
rect -15600 92350 -15400 92380
rect -15600 92150 -15590 92350
rect -15520 92150 -15480 92350
rect -15410 92150 -15400 92350
rect -15600 92120 -15400 92150
rect -15100 92350 -14900 92380
rect -15100 92150 -15090 92350
rect -15020 92150 -14980 92350
rect -14910 92150 -14900 92350
rect -15100 92120 -14900 92150
rect -14600 92350 -14400 92380
rect -14600 92150 -14590 92350
rect -14520 92150 -14480 92350
rect -14410 92150 -14400 92350
rect -14600 92120 -14400 92150
rect -14100 92350 -13900 92380
rect -14100 92150 -14090 92350
rect -14020 92150 -13980 92350
rect -13910 92150 -13900 92350
rect -14100 92120 -13900 92150
rect -13600 92350 -13400 92380
rect -13600 92150 -13590 92350
rect -13520 92150 -13480 92350
rect -13410 92150 -13400 92350
rect -13600 92120 -13400 92150
rect -13100 92350 -12900 92380
rect -13100 92150 -13090 92350
rect -13020 92150 -12980 92350
rect -12910 92150 -12900 92350
rect -13100 92120 -12900 92150
rect -12600 92350 -12400 92380
rect -12600 92150 -12590 92350
rect -12520 92150 -12480 92350
rect -12410 92150 -12400 92350
rect -12600 92120 -12400 92150
rect -12100 92350 -12000 92380
rect -12100 92150 -12090 92350
rect -12020 92150 -12000 92350
rect -12100 92120 -12000 92150
rect -16000 92100 -15880 92120
rect -15620 92100 -15380 92120
rect -15120 92100 -14880 92120
rect -14620 92100 -14380 92120
rect -14120 92100 -13880 92120
rect -13620 92100 -13380 92120
rect -13120 92100 -12880 92120
rect -12620 92100 -12380 92120
rect -12120 92100 -12000 92120
rect -16000 92090 -12000 92100
rect -16000 92020 -15850 92090
rect -15650 92020 -15350 92090
rect -15150 92020 -14850 92090
rect -14650 92020 -14350 92090
rect -14150 92020 -13850 92090
rect -13650 92020 -13350 92090
rect -13150 92020 -12850 92090
rect -12650 92020 -12350 92090
rect -12150 92020 -12000 92090
rect -16000 91980 -12000 92020
rect -16000 91910 -15850 91980
rect -15650 91910 -15350 91980
rect -15150 91910 -14850 91980
rect -14650 91910 -14350 91980
rect -14150 91910 -13850 91980
rect -13650 91910 -13350 91980
rect -13150 91910 -12850 91980
rect -12650 91910 -12350 91980
rect -12150 91910 -12000 91980
rect -16000 91900 -12000 91910
rect -16000 91880 -15880 91900
rect -15620 91880 -15380 91900
rect -15120 91880 -14880 91900
rect -14620 91880 -14380 91900
rect -14120 91880 -13880 91900
rect -13620 91880 -13380 91900
rect -13120 91880 -12880 91900
rect -12620 91880 -12380 91900
rect -12120 91880 -12000 91900
rect -16000 91850 -15900 91880
rect -16000 91650 -15980 91850
rect -15910 91650 -15900 91850
rect -16000 91620 -15900 91650
rect -15600 91850 -15400 91880
rect -15600 91650 -15590 91850
rect -15520 91650 -15480 91850
rect -15410 91650 -15400 91850
rect -15600 91620 -15400 91650
rect -15100 91850 -14900 91880
rect -15100 91650 -15090 91850
rect -15020 91650 -14980 91850
rect -14910 91650 -14900 91850
rect -15100 91620 -14900 91650
rect -14600 91850 -14400 91880
rect -14600 91650 -14590 91850
rect -14520 91650 -14480 91850
rect -14410 91650 -14400 91850
rect -14600 91620 -14400 91650
rect -14100 91850 -13900 91880
rect -14100 91650 -14090 91850
rect -14020 91650 -13980 91850
rect -13910 91650 -13900 91850
rect -14100 91620 -13900 91650
rect -13600 91850 -13400 91880
rect -13600 91650 -13590 91850
rect -13520 91650 -13480 91850
rect -13410 91650 -13400 91850
rect -13600 91620 -13400 91650
rect -13100 91850 -12900 91880
rect -13100 91650 -13090 91850
rect -13020 91650 -12980 91850
rect -12910 91650 -12900 91850
rect -13100 91620 -12900 91650
rect -12600 91850 -12400 91880
rect -12600 91650 -12590 91850
rect -12520 91650 -12480 91850
rect -12410 91650 -12400 91850
rect -12600 91620 -12400 91650
rect -12100 91850 -12000 91880
rect -12100 91650 -12090 91850
rect -12020 91650 -12000 91850
rect -12100 91620 -12000 91650
rect -16000 91600 -15880 91620
rect -15620 91600 -15380 91620
rect -15120 91600 -14880 91620
rect -14620 91600 -14380 91620
rect -14120 91600 -13880 91620
rect -13620 91600 -13380 91620
rect -13120 91600 -12880 91620
rect -12620 91600 -12380 91620
rect -12120 91600 -12000 91620
rect -16000 91590 -12000 91600
rect -16000 91520 -15850 91590
rect -15650 91520 -15350 91590
rect -15150 91520 -14850 91590
rect -14650 91520 -14350 91590
rect -14150 91520 -13850 91590
rect -13650 91520 -13350 91590
rect -13150 91520 -12850 91590
rect -12650 91520 -12350 91590
rect -12150 91520 -12000 91590
rect -16000 91480 -12000 91520
rect -16000 91410 -15850 91480
rect -15650 91410 -15350 91480
rect -15150 91410 -14850 91480
rect -14650 91410 -14350 91480
rect -14150 91410 -13850 91480
rect -13650 91410 -13350 91480
rect -13150 91410 -12850 91480
rect -12650 91410 -12350 91480
rect -12150 91410 -12000 91480
rect -16000 91400 -12000 91410
rect -16000 91380 -15880 91400
rect -15620 91380 -15380 91400
rect -15120 91380 -14880 91400
rect -14620 91380 -14380 91400
rect -14120 91380 -13880 91400
rect -13620 91380 -13380 91400
rect -13120 91380 -12880 91400
rect -12620 91380 -12380 91400
rect -12120 91380 -12000 91400
rect -16000 91350 -15900 91380
rect -16000 91150 -15980 91350
rect -15910 91150 -15900 91350
rect -16000 91120 -15900 91150
rect -15600 91350 -15400 91380
rect -15600 91150 -15590 91350
rect -15520 91150 -15480 91350
rect -15410 91150 -15400 91350
rect -15600 91120 -15400 91150
rect -15100 91350 -14900 91380
rect -15100 91150 -15090 91350
rect -15020 91150 -14980 91350
rect -14910 91150 -14900 91350
rect -15100 91120 -14900 91150
rect -14600 91350 -14400 91380
rect -14600 91150 -14590 91350
rect -14520 91150 -14480 91350
rect -14410 91150 -14400 91350
rect -14600 91120 -14400 91150
rect -14100 91350 -13900 91380
rect -14100 91150 -14090 91350
rect -14020 91150 -13980 91350
rect -13910 91150 -13900 91350
rect -14100 91120 -13900 91150
rect -13600 91350 -13400 91380
rect -13600 91150 -13590 91350
rect -13520 91150 -13480 91350
rect -13410 91150 -13400 91350
rect -13600 91120 -13400 91150
rect -13100 91350 -12900 91380
rect -13100 91150 -13090 91350
rect -13020 91150 -12980 91350
rect -12910 91150 -12900 91350
rect -13100 91120 -12900 91150
rect -12600 91350 -12400 91380
rect -12600 91150 -12590 91350
rect -12520 91150 -12480 91350
rect -12410 91150 -12400 91350
rect -12600 91120 -12400 91150
rect -12100 91350 -12000 91380
rect -12100 91150 -12090 91350
rect -12020 91150 -12000 91350
rect -12100 91120 -12000 91150
rect -16000 91100 -15880 91120
rect -15620 91100 -15380 91120
rect -15120 91100 -14880 91120
rect -14620 91100 -14380 91120
rect -14120 91100 -13880 91120
rect -13620 91100 -13380 91120
rect -13120 91100 -12880 91120
rect -12620 91100 -12380 91120
rect -12120 91100 -12000 91120
rect -16000 91090 -12000 91100
rect -16000 91020 -15850 91090
rect -15650 91020 -15350 91090
rect -15150 91020 -14850 91090
rect -14650 91020 -14350 91090
rect -14150 91020 -13850 91090
rect -13650 91020 -13350 91090
rect -13150 91020 -12850 91090
rect -12650 91020 -12350 91090
rect -12150 91020 -12000 91090
rect -16000 90980 -12000 91020
rect -16000 90910 -15850 90980
rect -15650 90910 -15350 90980
rect -15150 90910 -14850 90980
rect -14650 90910 -14350 90980
rect -14150 90910 -13850 90980
rect -13650 90910 -13350 90980
rect -13150 90910 -12850 90980
rect -12650 90910 -12350 90980
rect -12150 90910 -12000 90980
rect -16000 90900 -12000 90910
rect -16000 90880 -15880 90900
rect -15620 90880 -15380 90900
rect -15120 90880 -14880 90900
rect -14620 90880 -14380 90900
rect -14120 90880 -13880 90900
rect -13620 90880 -13380 90900
rect -13120 90880 -12880 90900
rect -12620 90880 -12380 90900
rect -12120 90880 -12000 90900
rect -16000 90850 -15900 90880
rect -16000 90650 -15980 90850
rect -15910 90650 -15900 90850
rect -16000 90620 -15900 90650
rect -15600 90850 -15400 90880
rect -15600 90650 -15590 90850
rect -15520 90650 -15480 90850
rect -15410 90650 -15400 90850
rect -15600 90620 -15400 90650
rect -15100 90850 -14900 90880
rect -15100 90650 -15090 90850
rect -15020 90650 -14980 90850
rect -14910 90650 -14900 90850
rect -15100 90620 -14900 90650
rect -14600 90850 -14400 90880
rect -14600 90650 -14590 90850
rect -14520 90650 -14480 90850
rect -14410 90650 -14400 90850
rect -14600 90620 -14400 90650
rect -14100 90850 -13900 90880
rect -14100 90650 -14090 90850
rect -14020 90650 -13980 90850
rect -13910 90650 -13900 90850
rect -14100 90620 -13900 90650
rect -13600 90850 -13400 90880
rect -13600 90650 -13590 90850
rect -13520 90650 -13480 90850
rect -13410 90650 -13400 90850
rect -13600 90620 -13400 90650
rect -13100 90850 -12900 90880
rect -13100 90650 -13090 90850
rect -13020 90650 -12980 90850
rect -12910 90650 -12900 90850
rect -13100 90620 -12900 90650
rect -12600 90850 -12400 90880
rect -12600 90650 -12590 90850
rect -12520 90650 -12480 90850
rect -12410 90650 -12400 90850
rect -12600 90620 -12400 90650
rect -12100 90850 -12000 90880
rect -12100 90650 -12090 90850
rect -12020 90650 -12000 90850
rect -12100 90620 -12000 90650
rect -16000 90600 -15880 90620
rect -15620 90600 -15380 90620
rect -15120 90600 -14880 90620
rect -14620 90600 -14380 90620
rect -14120 90600 -13880 90620
rect -13620 90600 -13380 90620
rect -13120 90600 -12880 90620
rect -12620 90600 -12380 90620
rect -12120 90600 -12000 90620
rect -16000 90590 -12000 90600
rect -16000 90520 -15850 90590
rect -15650 90520 -15350 90590
rect -15150 90520 -14850 90590
rect -14650 90520 -14350 90590
rect -14150 90520 -13850 90590
rect -13650 90520 -13350 90590
rect -13150 90520 -12850 90590
rect -12650 90520 -12350 90590
rect -12150 90520 -12000 90590
rect -16000 90480 -12000 90520
rect -16000 90410 -15850 90480
rect -15650 90410 -15350 90480
rect -15150 90410 -14850 90480
rect -14650 90410 -14350 90480
rect -14150 90410 -13850 90480
rect -13650 90410 -13350 90480
rect -13150 90410 -12850 90480
rect -12650 90410 -12350 90480
rect -12150 90410 -12000 90480
rect -16000 90400 -12000 90410
rect -16000 90380 -15880 90400
rect -15620 90380 -15380 90400
rect -15120 90380 -14880 90400
rect -14620 90380 -14380 90400
rect -14120 90380 -13880 90400
rect -13620 90380 -13380 90400
rect -13120 90380 -12880 90400
rect -12620 90380 -12380 90400
rect -12120 90380 -12000 90400
rect -16000 90350 -15900 90380
rect -16000 90150 -15980 90350
rect -15910 90150 -15900 90350
rect -16000 90120 -15900 90150
rect -15600 90350 -15400 90380
rect -15600 90150 -15590 90350
rect -15520 90150 -15480 90350
rect -15410 90150 -15400 90350
rect -15600 90120 -15400 90150
rect -15100 90350 -14900 90380
rect -15100 90150 -15090 90350
rect -15020 90150 -14980 90350
rect -14910 90150 -14900 90350
rect -15100 90120 -14900 90150
rect -14600 90350 -14400 90380
rect -14600 90150 -14590 90350
rect -14520 90150 -14480 90350
rect -14410 90150 -14400 90350
rect -14600 90120 -14400 90150
rect -14100 90350 -13900 90380
rect -14100 90150 -14090 90350
rect -14020 90150 -13980 90350
rect -13910 90150 -13900 90350
rect -14100 90120 -13900 90150
rect -13600 90350 -13400 90380
rect -13600 90150 -13590 90350
rect -13520 90150 -13480 90350
rect -13410 90150 -13400 90350
rect -13600 90120 -13400 90150
rect -13100 90350 -12900 90380
rect -13100 90150 -13090 90350
rect -13020 90150 -12980 90350
rect -12910 90150 -12900 90350
rect -13100 90120 -12900 90150
rect -12600 90350 -12400 90380
rect -12600 90150 -12590 90350
rect -12520 90150 -12480 90350
rect -12410 90150 -12400 90350
rect -12600 90120 -12400 90150
rect -12100 90350 -12000 90380
rect -12100 90150 -12090 90350
rect -12020 90150 -12000 90350
rect -12100 90120 -12000 90150
rect -16000 90100 -15880 90120
rect -15620 90100 -15380 90120
rect -15120 90100 -14880 90120
rect -14620 90100 -14380 90120
rect -14120 90100 -13880 90120
rect -13620 90100 -13380 90120
rect -13120 90100 -12880 90120
rect -12620 90100 -12380 90120
rect -12120 90100 -12000 90120
rect -16000 90090 -12000 90100
rect -16000 90020 -15850 90090
rect -15650 90020 -15350 90090
rect -15150 90020 -14850 90090
rect -14650 90020 -14350 90090
rect -14150 90020 -13850 90090
rect -13650 90020 -13350 90090
rect -13150 90020 -12850 90090
rect -12650 90020 -12350 90090
rect -12150 90020 -12000 90090
rect -16000 89980 -12000 90020
rect -16000 89910 -15850 89980
rect -15650 89910 -15350 89980
rect -15150 89910 -14850 89980
rect -14650 89910 -14350 89980
rect -14150 89910 -13850 89980
rect -13650 89910 -13350 89980
rect -13150 89910 -12850 89980
rect -12650 89910 -12350 89980
rect -12150 89910 -12000 89980
rect -16000 89900 -12000 89910
rect -16000 89880 -15880 89900
rect -15620 89880 -15380 89900
rect -15120 89880 -14880 89900
rect -14620 89880 -14380 89900
rect -14120 89880 -13880 89900
rect -13620 89880 -13380 89900
rect -13120 89880 -12880 89900
rect -12620 89880 -12380 89900
rect -12120 89880 -12000 89900
rect -16000 89850 -15900 89880
rect -16000 89650 -15980 89850
rect -15910 89650 -15900 89850
rect -16000 89620 -15900 89650
rect -15600 89850 -15400 89880
rect -15600 89650 -15590 89850
rect -15520 89650 -15480 89850
rect -15410 89650 -15400 89850
rect -15600 89620 -15400 89650
rect -15100 89850 -14900 89880
rect -15100 89650 -15090 89850
rect -15020 89650 -14980 89850
rect -14910 89650 -14900 89850
rect -15100 89620 -14900 89650
rect -14600 89850 -14400 89880
rect -14600 89650 -14590 89850
rect -14520 89650 -14480 89850
rect -14410 89650 -14400 89850
rect -14600 89620 -14400 89650
rect -14100 89850 -13900 89880
rect -14100 89650 -14090 89850
rect -14020 89650 -13980 89850
rect -13910 89650 -13900 89850
rect -14100 89620 -13900 89650
rect -13600 89850 -13400 89880
rect -13600 89650 -13590 89850
rect -13520 89650 -13480 89850
rect -13410 89650 -13400 89850
rect -13600 89620 -13400 89650
rect -13100 89850 -12900 89880
rect -13100 89650 -13090 89850
rect -13020 89650 -12980 89850
rect -12910 89650 -12900 89850
rect -13100 89620 -12900 89650
rect -12600 89850 -12400 89880
rect -12600 89650 -12590 89850
rect -12520 89650 -12480 89850
rect -12410 89650 -12400 89850
rect -12600 89620 -12400 89650
rect -12100 89850 -12000 89880
rect -12100 89650 -12090 89850
rect -12020 89650 -12000 89850
rect -12100 89620 -12000 89650
rect -16000 89600 -15880 89620
rect -15620 89600 -15380 89620
rect -15120 89600 -14880 89620
rect -14620 89600 -14380 89620
rect -14120 89600 -13880 89620
rect -13620 89600 -13380 89620
rect -13120 89600 -12880 89620
rect -12620 89600 -12380 89620
rect -12120 89600 -12000 89620
rect -16000 89590 -12000 89600
rect -16000 89520 -15850 89590
rect -15650 89520 -15350 89590
rect -15150 89520 -14850 89590
rect -14650 89520 -14350 89590
rect -14150 89520 -13850 89590
rect -13650 89520 -13350 89590
rect -13150 89520 -12850 89590
rect -12650 89520 -12350 89590
rect -12150 89520 -12000 89590
rect -16000 89480 -12000 89520
rect -16000 89410 -15850 89480
rect -15650 89410 -15350 89480
rect -15150 89410 -14850 89480
rect -14650 89410 -14350 89480
rect -14150 89410 -13850 89480
rect -13650 89410 -13350 89480
rect -13150 89410 -12850 89480
rect -12650 89410 -12350 89480
rect -12150 89410 -12000 89480
rect -16000 89400 -12000 89410
rect -16000 89380 -15880 89400
rect -15620 89380 -15380 89400
rect -15120 89380 -14880 89400
rect -14620 89380 -14380 89400
rect -14120 89380 -13880 89400
rect -13620 89380 -13380 89400
rect -13120 89380 -12880 89400
rect -12620 89380 -12380 89400
rect -12120 89380 -12000 89400
rect -16000 89350 -15900 89380
rect -16000 89150 -15980 89350
rect -15910 89150 -15900 89350
rect -16000 89120 -15900 89150
rect -15600 89350 -15400 89380
rect -15600 89150 -15590 89350
rect -15520 89150 -15480 89350
rect -15410 89150 -15400 89350
rect -15600 89120 -15400 89150
rect -15100 89350 -14900 89380
rect -15100 89150 -15090 89350
rect -15020 89150 -14980 89350
rect -14910 89150 -14900 89350
rect -15100 89120 -14900 89150
rect -14600 89350 -14400 89380
rect -14600 89150 -14590 89350
rect -14520 89150 -14480 89350
rect -14410 89150 -14400 89350
rect -14600 89120 -14400 89150
rect -14100 89350 -13900 89380
rect -14100 89150 -14090 89350
rect -14020 89150 -13980 89350
rect -13910 89150 -13900 89350
rect -14100 89120 -13900 89150
rect -13600 89350 -13400 89380
rect -13600 89150 -13590 89350
rect -13520 89150 -13480 89350
rect -13410 89150 -13400 89350
rect -13600 89120 -13400 89150
rect -13100 89350 -12900 89380
rect -13100 89150 -13090 89350
rect -13020 89150 -12980 89350
rect -12910 89150 -12900 89350
rect -13100 89120 -12900 89150
rect -12600 89350 -12400 89380
rect -12600 89150 -12590 89350
rect -12520 89150 -12480 89350
rect -12410 89150 -12400 89350
rect -12600 89120 -12400 89150
rect -12100 89350 -12000 89380
rect -12100 89150 -12090 89350
rect -12020 89150 -12000 89350
rect -12100 89120 -12000 89150
rect -16000 89100 -15880 89120
rect -15620 89100 -15380 89120
rect -15120 89100 -14880 89120
rect -14620 89100 -14380 89120
rect -14120 89100 -13880 89120
rect -13620 89100 -13380 89120
rect -13120 89100 -12880 89120
rect -12620 89100 -12380 89120
rect -12120 89100 -12000 89120
rect -16000 89090 -12000 89100
rect -16000 89020 -15850 89090
rect -15650 89020 -15350 89090
rect -15150 89020 -14850 89090
rect -14650 89020 -14350 89090
rect -14150 89020 -13850 89090
rect -13650 89020 -13350 89090
rect -13150 89020 -12850 89090
rect -12650 89020 -12350 89090
rect -12150 89020 -12000 89090
rect -16000 88980 -12000 89020
rect -16000 88910 -15850 88980
rect -15650 88910 -15350 88980
rect -15150 88910 -14850 88980
rect -14650 88910 -14350 88980
rect -14150 88910 -13850 88980
rect -13650 88910 -13350 88980
rect -13150 88910 -12850 88980
rect -12650 88910 -12350 88980
rect -12150 88910 -12000 88980
rect -16000 88900 -12000 88910
rect -16000 88880 -15880 88900
rect -15620 88880 -15380 88900
rect -15120 88880 -14880 88900
rect -14620 88880 -14380 88900
rect -14120 88880 -13880 88900
rect -13620 88880 -13380 88900
rect -13120 88880 -12880 88900
rect -12620 88880 -12380 88900
rect -12120 88880 -12000 88900
rect -16000 88850 -15900 88880
rect -16000 88650 -15980 88850
rect -15910 88650 -15900 88850
rect -16000 88620 -15900 88650
rect -15600 88850 -15400 88880
rect -15600 88650 -15590 88850
rect -15520 88650 -15480 88850
rect -15410 88650 -15400 88850
rect -15600 88620 -15400 88650
rect -15100 88850 -14900 88880
rect -15100 88650 -15090 88850
rect -15020 88650 -14980 88850
rect -14910 88650 -14900 88850
rect -15100 88620 -14900 88650
rect -14600 88850 -14400 88880
rect -14600 88650 -14590 88850
rect -14520 88650 -14480 88850
rect -14410 88650 -14400 88850
rect -14600 88620 -14400 88650
rect -14100 88850 -13900 88880
rect -14100 88650 -14090 88850
rect -14020 88650 -13980 88850
rect -13910 88650 -13900 88850
rect -14100 88620 -13900 88650
rect -13600 88850 -13400 88880
rect -13600 88650 -13590 88850
rect -13520 88650 -13480 88850
rect -13410 88650 -13400 88850
rect -13600 88620 -13400 88650
rect -13100 88850 -12900 88880
rect -13100 88650 -13090 88850
rect -13020 88650 -12980 88850
rect -12910 88650 -12900 88850
rect -13100 88620 -12900 88650
rect -12600 88850 -12400 88880
rect -12600 88650 -12590 88850
rect -12520 88650 -12480 88850
rect -12410 88650 -12400 88850
rect -12600 88620 -12400 88650
rect -12100 88850 -12000 88880
rect -12100 88650 -12090 88850
rect -12020 88650 -12000 88850
rect -12100 88620 -12000 88650
rect -16000 88600 -15880 88620
rect -15620 88600 -15380 88620
rect -15120 88600 -14880 88620
rect -14620 88600 -14380 88620
rect -14120 88600 -13880 88620
rect -13620 88600 -13380 88620
rect -13120 88600 -12880 88620
rect -12620 88600 -12380 88620
rect -12120 88600 -12000 88620
rect -16000 88590 -12000 88600
rect -16000 88520 -15850 88590
rect -15650 88520 -15350 88590
rect -15150 88520 -14850 88590
rect -14650 88520 -14350 88590
rect -14150 88520 -13850 88590
rect -13650 88520 -13350 88590
rect -13150 88520 -12850 88590
rect -12650 88520 -12350 88590
rect -12150 88520 -12000 88590
rect -16000 88480 -12000 88520
rect -16000 88410 -15850 88480
rect -15650 88410 -15350 88480
rect -15150 88410 -14850 88480
rect -14650 88410 -14350 88480
rect -14150 88410 -13850 88480
rect -13650 88410 -13350 88480
rect -13150 88410 -12850 88480
rect -12650 88410 -12350 88480
rect -12150 88410 -12000 88480
rect -16000 88400 -12000 88410
rect -16000 88380 -15880 88400
rect -15620 88380 -15380 88400
rect -15120 88380 -14880 88400
rect -14620 88380 -14380 88400
rect -14120 88380 -13880 88400
rect -13620 88380 -13380 88400
rect -13120 88380 -12880 88400
rect -12620 88380 -12380 88400
rect -12120 88380 -12000 88400
rect -16000 88350 -15900 88380
rect -16000 88150 -15980 88350
rect -15910 88150 -15900 88350
rect -16000 88120 -15900 88150
rect -15600 88350 -15400 88380
rect -15600 88150 -15590 88350
rect -15520 88150 -15480 88350
rect -15410 88150 -15400 88350
rect -15600 88120 -15400 88150
rect -15100 88350 -14900 88380
rect -15100 88150 -15090 88350
rect -15020 88150 -14980 88350
rect -14910 88150 -14900 88350
rect -15100 88120 -14900 88150
rect -14600 88350 -14400 88380
rect -14600 88150 -14590 88350
rect -14520 88150 -14480 88350
rect -14410 88150 -14400 88350
rect -14600 88120 -14400 88150
rect -14100 88350 -13900 88380
rect -14100 88150 -14090 88350
rect -14020 88150 -13980 88350
rect -13910 88150 -13900 88350
rect -14100 88120 -13900 88150
rect -13600 88350 -13400 88380
rect -13600 88150 -13590 88350
rect -13520 88150 -13480 88350
rect -13410 88150 -13400 88350
rect -13600 88120 -13400 88150
rect -13100 88350 -12900 88380
rect -13100 88150 -13090 88350
rect -13020 88150 -12980 88350
rect -12910 88150 -12900 88350
rect -13100 88120 -12900 88150
rect -12600 88350 -12400 88380
rect -12600 88150 -12590 88350
rect -12520 88150 -12480 88350
rect -12410 88150 -12400 88350
rect -12600 88120 -12400 88150
rect -12100 88350 -12000 88380
rect -12100 88150 -12090 88350
rect -12020 88150 -12000 88350
rect -12100 88120 -12000 88150
rect -16000 88100 -15880 88120
rect -15620 88100 -15380 88120
rect -15120 88100 -14880 88120
rect -14620 88100 -14380 88120
rect -14120 88100 -13880 88120
rect -13620 88100 -13380 88120
rect -13120 88100 -12880 88120
rect -12620 88100 -12380 88120
rect -12120 88100 -12000 88120
rect -16000 88090 -12000 88100
rect -16000 88020 -15850 88090
rect -15650 88020 -15350 88090
rect -15150 88020 -14850 88090
rect -14650 88020 -14350 88090
rect -14150 88020 -13850 88090
rect -13650 88020 -13350 88090
rect -13150 88020 -12850 88090
rect -12650 88020 -12350 88090
rect -12150 88020 -12000 88090
rect -16000 87980 -12000 88020
rect -16000 87910 -15850 87980
rect -15650 87910 -15350 87980
rect -15150 87910 -14850 87980
rect -14650 87910 -14350 87980
rect -14150 87910 -13850 87980
rect -13650 87910 -13350 87980
rect -13150 87910 -12850 87980
rect -12650 87910 -12350 87980
rect -12150 87910 -12000 87980
rect -16000 87900 -12000 87910
rect -16000 87880 -15880 87900
rect -15620 87880 -15380 87900
rect -15120 87880 -14880 87900
rect -14620 87880 -14380 87900
rect -14120 87880 -13880 87900
rect -13620 87880 -13380 87900
rect -13120 87880 -12880 87900
rect -12620 87880 -12380 87900
rect -12120 87880 -12000 87900
rect -16000 87850 -15900 87880
rect -16000 87650 -15980 87850
rect -15910 87650 -15900 87850
rect -16000 87620 -15900 87650
rect -15600 87850 -15400 87880
rect -15600 87650 -15590 87850
rect -15520 87650 -15480 87850
rect -15410 87650 -15400 87850
rect -15600 87620 -15400 87650
rect -15100 87850 -14900 87880
rect -15100 87650 -15090 87850
rect -15020 87650 -14980 87850
rect -14910 87650 -14900 87850
rect -15100 87620 -14900 87650
rect -14600 87850 -14400 87880
rect -14600 87650 -14590 87850
rect -14520 87650 -14480 87850
rect -14410 87650 -14400 87850
rect -14600 87620 -14400 87650
rect -14100 87850 -13900 87880
rect -14100 87650 -14090 87850
rect -14020 87650 -13980 87850
rect -13910 87650 -13900 87850
rect -14100 87620 -13900 87650
rect -13600 87850 -13400 87880
rect -13600 87650 -13590 87850
rect -13520 87650 -13480 87850
rect -13410 87650 -13400 87850
rect -13600 87620 -13400 87650
rect -13100 87850 -12900 87880
rect -13100 87650 -13090 87850
rect -13020 87650 -12980 87850
rect -12910 87650 -12900 87850
rect -13100 87620 -12900 87650
rect -12600 87850 -12400 87880
rect -12600 87650 -12590 87850
rect -12520 87650 -12480 87850
rect -12410 87650 -12400 87850
rect -12600 87620 -12400 87650
rect -12100 87850 -12000 87880
rect -12100 87650 -12090 87850
rect -12020 87650 -12000 87850
rect -12100 87620 -12000 87650
rect -16000 87600 -15880 87620
rect -15620 87600 -15380 87620
rect -15120 87600 -14880 87620
rect -14620 87600 -14380 87620
rect -14120 87600 -13880 87620
rect -13620 87600 -13380 87620
rect -13120 87600 -12880 87620
rect -12620 87600 -12380 87620
rect -12120 87600 -12000 87620
rect -16000 87590 -12000 87600
rect -16000 87520 -15850 87590
rect -15650 87520 -15350 87590
rect -15150 87520 -14850 87590
rect -14650 87520 -14350 87590
rect -14150 87520 -13850 87590
rect -13650 87520 -13350 87590
rect -13150 87520 -12850 87590
rect -12650 87520 -12350 87590
rect -12150 87520 -12000 87590
rect -16000 87480 -12000 87520
rect -16000 87410 -15850 87480
rect -15650 87410 -15350 87480
rect -15150 87410 -14850 87480
rect -14650 87410 -14350 87480
rect -14150 87410 -13850 87480
rect -13650 87410 -13350 87480
rect -13150 87410 -12850 87480
rect -12650 87410 -12350 87480
rect -12150 87410 -12000 87480
rect -16000 87400 -12000 87410
rect -16000 87380 -15880 87400
rect -15620 87380 -15380 87400
rect -15120 87380 -14880 87400
rect -14620 87380 -14380 87400
rect -14120 87380 -13880 87400
rect -13620 87380 -13380 87400
rect -13120 87380 -12880 87400
rect -12620 87380 -12380 87400
rect -12120 87380 -12000 87400
rect -16000 87350 -15900 87380
rect -16000 87150 -15980 87350
rect -15910 87150 -15900 87350
rect -16000 87120 -15900 87150
rect -15600 87350 -15400 87380
rect -15600 87150 -15590 87350
rect -15520 87150 -15480 87350
rect -15410 87150 -15400 87350
rect -15600 87120 -15400 87150
rect -15100 87350 -14900 87380
rect -15100 87150 -15090 87350
rect -15020 87150 -14980 87350
rect -14910 87150 -14900 87350
rect -15100 87120 -14900 87150
rect -14600 87350 -14400 87380
rect -14600 87150 -14590 87350
rect -14520 87150 -14480 87350
rect -14410 87150 -14400 87350
rect -14600 87120 -14400 87150
rect -14100 87350 -13900 87380
rect -14100 87150 -14090 87350
rect -14020 87150 -13980 87350
rect -13910 87150 -13900 87350
rect -14100 87120 -13900 87150
rect -13600 87350 -13400 87380
rect -13600 87150 -13590 87350
rect -13520 87150 -13480 87350
rect -13410 87150 -13400 87350
rect -13600 87120 -13400 87150
rect -13100 87350 -12900 87380
rect -13100 87150 -13090 87350
rect -13020 87150 -12980 87350
rect -12910 87150 -12900 87350
rect -13100 87120 -12900 87150
rect -12600 87350 -12400 87380
rect -12600 87150 -12590 87350
rect -12520 87150 -12480 87350
rect -12410 87150 -12400 87350
rect -12600 87120 -12400 87150
rect -12100 87350 -12000 87380
rect -12100 87150 -12090 87350
rect -12020 87150 -12000 87350
rect -12100 87120 -12000 87150
rect -16000 87100 -15880 87120
rect -15620 87100 -15380 87120
rect -15120 87100 -14880 87120
rect -14620 87100 -14380 87120
rect -14120 87100 -13880 87120
rect -13620 87100 -13380 87120
rect -13120 87100 -12880 87120
rect -12620 87100 -12380 87120
rect -12120 87100 -12000 87120
rect -16000 87090 -12000 87100
rect -16000 87020 -15850 87090
rect -15650 87020 -15350 87090
rect -15150 87020 -14850 87090
rect -14650 87020 -14350 87090
rect -14150 87020 -13850 87090
rect -13650 87020 -13350 87090
rect -13150 87020 -12850 87090
rect -12650 87020 -12350 87090
rect -12150 87020 -12000 87090
rect -16000 86980 -12000 87020
rect -16000 86910 -15850 86980
rect -15650 86910 -15350 86980
rect -15150 86910 -14850 86980
rect -14650 86910 -14350 86980
rect -14150 86910 -13850 86980
rect -13650 86910 -13350 86980
rect -13150 86910 -12850 86980
rect -12650 86910 -12350 86980
rect -12150 86910 -12000 86980
rect -16000 86900 -12000 86910
rect -16000 86880 -15880 86900
rect -15620 86880 -15380 86900
rect -15120 86880 -14880 86900
rect -14620 86880 -14380 86900
rect -14120 86880 -13880 86900
rect -13620 86880 -13380 86900
rect -13120 86880 -12880 86900
rect -12620 86880 -12380 86900
rect -12120 86880 -12000 86900
rect -16000 86850 -15900 86880
rect -16000 86650 -15980 86850
rect -15910 86650 -15900 86850
rect -16000 86620 -15900 86650
rect -15600 86850 -15400 86880
rect -15600 86650 -15590 86850
rect -15520 86650 -15480 86850
rect -15410 86650 -15400 86850
rect -15600 86620 -15400 86650
rect -15100 86850 -14900 86880
rect -15100 86650 -15090 86850
rect -15020 86650 -14980 86850
rect -14910 86650 -14900 86850
rect -15100 86620 -14900 86650
rect -14600 86850 -14400 86880
rect -14600 86650 -14590 86850
rect -14520 86650 -14480 86850
rect -14410 86650 -14400 86850
rect -14600 86620 -14400 86650
rect -14100 86850 -13900 86880
rect -14100 86650 -14090 86850
rect -14020 86650 -13980 86850
rect -13910 86650 -13900 86850
rect -14100 86620 -13900 86650
rect -13600 86850 -13400 86880
rect -13600 86650 -13590 86850
rect -13520 86650 -13480 86850
rect -13410 86650 -13400 86850
rect -13600 86620 -13400 86650
rect -13100 86850 -12900 86880
rect -13100 86650 -13090 86850
rect -13020 86650 -12980 86850
rect -12910 86650 -12900 86850
rect -13100 86620 -12900 86650
rect -12600 86850 -12400 86880
rect -12600 86650 -12590 86850
rect -12520 86650 -12480 86850
rect -12410 86650 -12400 86850
rect -12600 86620 -12400 86650
rect -12100 86850 -12000 86880
rect -12100 86650 -12090 86850
rect -12020 86650 -12000 86850
rect -12100 86620 -12000 86650
rect -16000 86600 -15880 86620
rect -15620 86600 -15380 86620
rect -15120 86600 -14880 86620
rect -14620 86600 -14380 86620
rect -14120 86600 -13880 86620
rect -13620 86600 -13380 86620
rect -13120 86600 -12880 86620
rect -12620 86600 -12380 86620
rect -12120 86600 -12000 86620
rect -16000 86590 -12000 86600
rect -16000 86520 -15850 86590
rect -15650 86520 -15350 86590
rect -15150 86520 -14850 86590
rect -14650 86520 -14350 86590
rect -14150 86520 -13850 86590
rect -13650 86520 -13350 86590
rect -13150 86520 -12850 86590
rect -12650 86520 -12350 86590
rect -12150 86520 -12000 86590
rect -16000 86480 -12000 86520
rect -16000 86410 -15850 86480
rect -15650 86410 -15350 86480
rect -15150 86410 -14850 86480
rect -14650 86410 -14350 86480
rect -14150 86410 -13850 86480
rect -13650 86410 -13350 86480
rect -13150 86410 -12850 86480
rect -12650 86410 -12350 86480
rect -12150 86410 -12000 86480
rect -16000 86400 -12000 86410
rect -16000 86380 -15880 86400
rect -15620 86380 -15380 86400
rect -15120 86380 -14880 86400
rect -14620 86380 -14380 86400
rect -14120 86380 -13880 86400
rect -13620 86380 -13380 86400
rect -13120 86380 -12880 86400
rect -12620 86380 -12380 86400
rect -12120 86380 -12000 86400
rect -16000 86350 -15900 86380
rect -16000 86150 -15980 86350
rect -15910 86150 -15900 86350
rect -16000 86120 -15900 86150
rect -15600 86350 -15400 86380
rect -15600 86150 -15590 86350
rect -15520 86150 -15480 86350
rect -15410 86150 -15400 86350
rect -15600 86120 -15400 86150
rect -15100 86350 -14900 86380
rect -15100 86150 -15090 86350
rect -15020 86150 -14980 86350
rect -14910 86150 -14900 86350
rect -15100 86120 -14900 86150
rect -14600 86350 -14400 86380
rect -14600 86150 -14590 86350
rect -14520 86150 -14480 86350
rect -14410 86150 -14400 86350
rect -14600 86120 -14400 86150
rect -14100 86350 -13900 86380
rect -14100 86150 -14090 86350
rect -14020 86150 -13980 86350
rect -13910 86150 -13900 86350
rect -14100 86120 -13900 86150
rect -13600 86350 -13400 86380
rect -13600 86150 -13590 86350
rect -13520 86150 -13480 86350
rect -13410 86150 -13400 86350
rect -13600 86120 -13400 86150
rect -13100 86350 -12900 86380
rect -13100 86150 -13090 86350
rect -13020 86150 -12980 86350
rect -12910 86150 -12900 86350
rect -13100 86120 -12900 86150
rect -12600 86350 -12400 86380
rect -12600 86150 -12590 86350
rect -12520 86150 -12480 86350
rect -12410 86150 -12400 86350
rect -12600 86120 -12400 86150
rect -12100 86350 -12000 86380
rect -12100 86150 -12090 86350
rect -12020 86150 -12000 86350
rect -12100 86120 -12000 86150
rect -16000 86100 -15880 86120
rect -15620 86100 -15380 86120
rect -15120 86100 -14880 86120
rect -14620 86100 -14380 86120
rect -14120 86100 -13880 86120
rect -13620 86100 -13380 86120
rect -13120 86100 -12880 86120
rect -12620 86100 -12380 86120
rect -12120 86100 -12000 86120
rect -16000 86090 -12000 86100
rect -16000 86020 -15850 86090
rect -15650 86020 -15350 86090
rect -15150 86020 -14850 86090
rect -14650 86020 -14350 86090
rect -14150 86020 -13850 86090
rect -13650 86020 -13350 86090
rect -13150 86020 -12850 86090
rect -12650 86020 -12350 86090
rect -12150 86020 -12000 86090
rect -16000 85980 -12000 86020
rect -16000 85910 -15850 85980
rect -15650 85910 -15350 85980
rect -15150 85910 -14850 85980
rect -14650 85910 -14350 85980
rect -14150 85910 -13850 85980
rect -13650 85910 -13350 85980
rect -13150 85910 -12850 85980
rect -12650 85910 -12350 85980
rect -12150 85910 -12000 85980
rect -16000 85900 -12000 85910
rect -16000 85880 -15880 85900
rect -15620 85880 -15380 85900
rect -15120 85880 -14880 85900
rect -14620 85880 -14380 85900
rect -14120 85880 -13880 85900
rect -13620 85880 -13380 85900
rect -13120 85880 -12880 85900
rect -12620 85880 -12380 85900
rect -12120 85880 -12000 85900
rect -16000 85850 -15900 85880
rect -16000 85650 -15980 85850
rect -15910 85650 -15900 85850
rect -16000 85620 -15900 85650
rect -15600 85850 -15400 85880
rect -15600 85650 -15590 85850
rect -15520 85650 -15480 85850
rect -15410 85650 -15400 85850
rect -15600 85620 -15400 85650
rect -15100 85850 -14900 85880
rect -15100 85650 -15090 85850
rect -15020 85650 -14980 85850
rect -14910 85650 -14900 85850
rect -15100 85620 -14900 85650
rect -14600 85850 -14400 85880
rect -14600 85650 -14590 85850
rect -14520 85650 -14480 85850
rect -14410 85650 -14400 85850
rect -14600 85620 -14400 85650
rect -14100 85850 -13900 85880
rect -14100 85650 -14090 85850
rect -14020 85650 -13980 85850
rect -13910 85650 -13900 85850
rect -14100 85620 -13900 85650
rect -13600 85850 -13400 85880
rect -13600 85650 -13590 85850
rect -13520 85650 -13480 85850
rect -13410 85650 -13400 85850
rect -13600 85620 -13400 85650
rect -13100 85850 -12900 85880
rect -13100 85650 -13090 85850
rect -13020 85650 -12980 85850
rect -12910 85650 -12900 85850
rect -13100 85620 -12900 85650
rect -12600 85850 -12400 85880
rect -12600 85650 -12590 85850
rect -12520 85650 -12480 85850
rect -12410 85650 -12400 85850
rect -12600 85620 -12400 85650
rect -12100 85850 -12000 85880
rect -12100 85650 -12090 85850
rect -12020 85650 -12000 85850
rect -12100 85620 -12000 85650
rect -16000 85600 -15880 85620
rect -15620 85600 -15380 85620
rect -15120 85600 -14880 85620
rect -14620 85600 -14380 85620
rect -14120 85600 -13880 85620
rect -13620 85600 -13380 85620
rect -13120 85600 -12880 85620
rect -12620 85600 -12380 85620
rect -12120 85600 -12000 85620
rect -16000 85590 -12000 85600
rect -16000 85520 -15850 85590
rect -15650 85520 -15350 85590
rect -15150 85520 -14850 85590
rect -14650 85520 -14350 85590
rect -14150 85520 -13850 85590
rect -13650 85520 -13350 85590
rect -13150 85520 -12850 85590
rect -12650 85520 -12350 85590
rect -12150 85520 -12000 85590
rect -16000 85480 -12000 85520
rect -16000 85410 -15850 85480
rect -15650 85410 -15350 85480
rect -15150 85410 -14850 85480
rect -14650 85410 -14350 85480
rect -14150 85410 -13850 85480
rect -13650 85410 -13350 85480
rect -13150 85410 -12850 85480
rect -12650 85410 -12350 85480
rect -12150 85410 -12000 85480
rect -16000 85400 -12000 85410
rect -16000 85380 -15880 85400
rect -15620 85380 -15380 85400
rect -15120 85380 -14880 85400
rect -14620 85380 -14380 85400
rect -14120 85380 -13880 85400
rect -13620 85380 -13380 85400
rect -13120 85380 -12880 85400
rect -12620 85380 -12380 85400
rect -12120 85380 -12000 85400
rect -16000 85350 -15900 85380
rect -16000 85150 -15980 85350
rect -15910 85150 -15900 85350
rect -16000 85120 -15900 85150
rect -15600 85350 -15400 85380
rect -15600 85150 -15590 85350
rect -15520 85150 -15480 85350
rect -15410 85150 -15400 85350
rect -15600 85120 -15400 85150
rect -15100 85350 -14900 85380
rect -15100 85150 -15090 85350
rect -15020 85150 -14980 85350
rect -14910 85150 -14900 85350
rect -15100 85120 -14900 85150
rect -14600 85350 -14400 85380
rect -14600 85150 -14590 85350
rect -14520 85150 -14480 85350
rect -14410 85150 -14400 85350
rect -14600 85120 -14400 85150
rect -14100 85350 -13900 85380
rect -14100 85150 -14090 85350
rect -14020 85150 -13980 85350
rect -13910 85150 -13900 85350
rect -14100 85120 -13900 85150
rect -13600 85350 -13400 85380
rect -13600 85150 -13590 85350
rect -13520 85150 -13480 85350
rect -13410 85150 -13400 85350
rect -13600 85120 -13400 85150
rect -13100 85350 -12900 85380
rect -13100 85150 -13090 85350
rect -13020 85150 -12980 85350
rect -12910 85150 -12900 85350
rect -13100 85120 -12900 85150
rect -12600 85350 -12400 85380
rect -12600 85150 -12590 85350
rect -12520 85150 -12480 85350
rect -12410 85150 -12400 85350
rect -12600 85120 -12400 85150
rect -12100 85350 -12000 85380
rect -12100 85150 -12090 85350
rect -12020 85150 -12000 85350
rect -12100 85120 -12000 85150
rect -16000 85100 -15880 85120
rect -15620 85100 -15380 85120
rect -15120 85100 -14880 85120
rect -14620 85100 -14380 85120
rect -14120 85100 -13880 85120
rect -13620 85100 -13380 85120
rect -13120 85100 -12880 85120
rect -12620 85100 -12380 85120
rect -12120 85100 -12000 85120
rect -16000 85090 -12000 85100
rect -16000 85020 -15850 85090
rect -15650 85020 -15350 85090
rect -15150 85020 -14850 85090
rect -14650 85020 -14350 85090
rect -14150 85020 -13850 85090
rect -13650 85020 -13350 85090
rect -13150 85020 -12850 85090
rect -12650 85020 -12350 85090
rect -12150 85020 -12000 85090
rect -16000 84980 -12000 85020
rect -16000 84910 -15850 84980
rect -15650 84910 -15350 84980
rect -15150 84910 -14850 84980
rect -14650 84910 -14350 84980
rect -14150 84910 -13850 84980
rect -13650 84910 -13350 84980
rect -13150 84910 -12850 84980
rect -12650 84910 -12350 84980
rect -12150 84910 -12000 84980
rect -16000 84900 -12000 84910
rect -16000 84880 -15880 84900
rect -15620 84880 -15380 84900
rect -15120 84880 -14880 84900
rect -14620 84880 -14380 84900
rect -14120 84880 -13880 84900
rect -13620 84880 -13380 84900
rect -13120 84880 -12880 84900
rect -12620 84880 -12380 84900
rect -12120 84880 -12000 84900
rect -16000 84850 -15900 84880
rect -16000 84650 -15980 84850
rect -15910 84650 -15900 84850
rect -16000 84620 -15900 84650
rect -15600 84850 -15400 84880
rect -15600 84650 -15590 84850
rect -15520 84650 -15480 84850
rect -15410 84650 -15400 84850
rect -15600 84620 -15400 84650
rect -15100 84850 -14900 84880
rect -15100 84650 -15090 84850
rect -15020 84650 -14980 84850
rect -14910 84650 -14900 84850
rect -15100 84620 -14900 84650
rect -14600 84850 -14400 84880
rect -14600 84650 -14590 84850
rect -14520 84650 -14480 84850
rect -14410 84650 -14400 84850
rect -14600 84620 -14400 84650
rect -14100 84850 -13900 84880
rect -14100 84650 -14090 84850
rect -14020 84650 -13980 84850
rect -13910 84650 -13900 84850
rect -14100 84620 -13900 84650
rect -13600 84850 -13400 84880
rect -13600 84650 -13590 84850
rect -13520 84650 -13480 84850
rect -13410 84650 -13400 84850
rect -13600 84620 -13400 84650
rect -13100 84850 -12900 84880
rect -13100 84650 -13090 84850
rect -13020 84650 -12980 84850
rect -12910 84650 -12900 84850
rect -13100 84620 -12900 84650
rect -12600 84850 -12400 84880
rect -12600 84650 -12590 84850
rect -12520 84650 -12480 84850
rect -12410 84650 -12400 84850
rect -12600 84620 -12400 84650
rect -12100 84850 -12000 84880
rect -12100 84650 -12090 84850
rect -12020 84650 -12000 84850
rect -12100 84620 -12000 84650
rect -16000 84600 -15880 84620
rect -15620 84600 -15380 84620
rect -15120 84600 -14880 84620
rect -14620 84600 -14380 84620
rect -14120 84600 -13880 84620
rect -13620 84600 -13380 84620
rect -13120 84600 -12880 84620
rect -12620 84600 -12380 84620
rect -12120 84600 -12000 84620
rect -16000 84590 -12000 84600
rect -16000 84520 -15850 84590
rect -15650 84520 -15350 84590
rect -15150 84520 -14850 84590
rect -14650 84520 -14350 84590
rect -14150 84520 -13850 84590
rect -13650 84520 -13350 84590
rect -13150 84520 -12850 84590
rect -12650 84520 -12350 84590
rect -12150 84520 -12000 84590
rect -16000 84480 -12000 84520
rect -16000 84410 -15850 84480
rect -15650 84410 -15350 84480
rect -15150 84410 -14850 84480
rect -14650 84410 -14350 84480
rect -14150 84410 -13850 84480
rect -13650 84410 -13350 84480
rect -13150 84410 -12850 84480
rect -12650 84410 -12350 84480
rect -12150 84410 -12000 84480
rect -16000 84400 -12000 84410
rect -16000 84380 -15880 84400
rect -15620 84380 -15380 84400
rect -15120 84380 -14880 84400
rect -14620 84380 -14380 84400
rect -14120 84380 -13880 84400
rect -13620 84380 -13380 84400
rect -13120 84380 -12880 84400
rect -12620 84380 -12380 84400
rect -12120 84380 -12000 84400
rect -16000 84350 -15900 84380
rect -16000 84150 -15980 84350
rect -15910 84150 -15900 84350
rect -16000 84120 -15900 84150
rect -15600 84350 -15400 84380
rect -15600 84150 -15590 84350
rect -15520 84150 -15480 84350
rect -15410 84150 -15400 84350
rect -15600 84120 -15400 84150
rect -15100 84350 -14900 84380
rect -15100 84150 -15090 84350
rect -15020 84150 -14980 84350
rect -14910 84150 -14900 84350
rect -15100 84120 -14900 84150
rect -14600 84350 -14400 84380
rect -14600 84150 -14590 84350
rect -14520 84150 -14480 84350
rect -14410 84150 -14400 84350
rect -14600 84120 -14400 84150
rect -14100 84350 -13900 84380
rect -14100 84150 -14090 84350
rect -14020 84150 -13980 84350
rect -13910 84150 -13900 84350
rect -14100 84120 -13900 84150
rect -13600 84350 -13400 84380
rect -13600 84150 -13590 84350
rect -13520 84150 -13480 84350
rect -13410 84150 -13400 84350
rect -13600 84120 -13400 84150
rect -13100 84350 -12900 84380
rect -13100 84150 -13090 84350
rect -13020 84150 -12980 84350
rect -12910 84150 -12900 84350
rect -13100 84120 -12900 84150
rect -12600 84350 -12400 84380
rect -12600 84150 -12590 84350
rect -12520 84150 -12480 84350
rect -12410 84150 -12400 84350
rect -12600 84120 -12400 84150
rect -12100 84350 -12000 84380
rect -12100 84150 -12090 84350
rect -12020 84150 -12000 84350
rect -12100 84120 -12000 84150
rect -16000 84100 -15880 84120
rect -15620 84100 -15380 84120
rect -15120 84100 -14880 84120
rect -14620 84100 -14380 84120
rect -14120 84100 -13880 84120
rect -13620 84100 -13380 84120
rect -13120 84100 -12880 84120
rect -12620 84100 -12380 84120
rect -12120 84100 -12000 84120
rect -16000 84090 -12000 84100
rect -16000 84020 -15850 84090
rect -15650 84020 -15350 84090
rect -15150 84020 -14850 84090
rect -14650 84020 -14350 84090
rect -14150 84020 -13850 84090
rect -13650 84020 -13350 84090
rect -13150 84020 -12850 84090
rect -12650 84020 -12350 84090
rect -12150 84020 -12000 84090
rect -16000 83980 -12000 84020
rect -16000 83910 -15850 83980
rect -15650 83910 -15350 83980
rect -15150 83910 -14850 83980
rect -14650 83910 -14350 83980
rect -14150 83910 -13850 83980
rect -13650 83910 -13350 83980
rect -13150 83910 -12850 83980
rect -12650 83910 -12350 83980
rect -12150 83910 -12000 83980
rect -16000 83900 -12000 83910
rect -16000 83880 -15880 83900
rect -15620 83880 -15380 83900
rect -15120 83880 -14880 83900
rect -14620 83880 -14380 83900
rect -14120 83880 -13880 83900
rect -13620 83880 -13380 83900
rect -13120 83880 -12880 83900
rect -12620 83880 -12380 83900
rect -12120 83880 -12000 83900
rect -16000 83850 -15900 83880
rect -16000 83650 -15980 83850
rect -15910 83650 -15900 83850
rect -16000 83620 -15900 83650
rect -15600 83850 -15400 83880
rect -15600 83650 -15590 83850
rect -15520 83650 -15480 83850
rect -15410 83650 -15400 83850
rect -15600 83620 -15400 83650
rect -15100 83850 -14900 83880
rect -15100 83650 -15090 83850
rect -15020 83650 -14980 83850
rect -14910 83650 -14900 83850
rect -15100 83620 -14900 83650
rect -14600 83850 -14400 83880
rect -14600 83650 -14590 83850
rect -14520 83650 -14480 83850
rect -14410 83650 -14400 83850
rect -14600 83620 -14400 83650
rect -14100 83850 -13900 83880
rect -14100 83650 -14090 83850
rect -14020 83650 -13980 83850
rect -13910 83650 -13900 83850
rect -14100 83620 -13900 83650
rect -13600 83850 -13400 83880
rect -13600 83650 -13590 83850
rect -13520 83650 -13480 83850
rect -13410 83650 -13400 83850
rect -13600 83620 -13400 83650
rect -13100 83850 -12900 83880
rect -13100 83650 -13090 83850
rect -13020 83650 -12980 83850
rect -12910 83650 -12900 83850
rect -13100 83620 -12900 83650
rect -12600 83850 -12400 83880
rect -12600 83650 -12590 83850
rect -12520 83650 -12480 83850
rect -12410 83650 -12400 83850
rect -12600 83620 -12400 83650
rect -12100 83850 -12000 83880
rect -12100 83650 -12090 83850
rect -12020 83650 -12000 83850
rect -12100 83620 -12000 83650
rect -16000 83600 -15880 83620
rect -15620 83600 -15380 83620
rect -15120 83600 -14880 83620
rect -14620 83600 -14380 83620
rect -14120 83600 -13880 83620
rect -13620 83600 -13380 83620
rect -13120 83600 -12880 83620
rect -12620 83600 -12380 83620
rect -12120 83600 -12000 83620
rect -16000 83590 -12000 83600
rect -16000 83520 -15850 83590
rect -15650 83520 -15350 83590
rect -15150 83520 -14850 83590
rect -14650 83520 -14350 83590
rect -14150 83520 -13850 83590
rect -13650 83520 -13350 83590
rect -13150 83520 -12850 83590
rect -12650 83520 -12350 83590
rect -12150 83520 -12000 83590
rect -16000 83480 -12000 83520
rect -16000 83410 -15850 83480
rect -15650 83410 -15350 83480
rect -15150 83410 -14850 83480
rect -14650 83410 -14350 83480
rect -14150 83410 -13850 83480
rect -13650 83410 -13350 83480
rect -13150 83410 -12850 83480
rect -12650 83410 -12350 83480
rect -12150 83410 -12000 83480
rect -16000 83400 -12000 83410
rect -16000 83380 -15880 83400
rect -15620 83380 -15380 83400
rect -15120 83380 -14880 83400
rect -14620 83380 -14380 83400
rect -14120 83380 -13880 83400
rect -13620 83380 -13380 83400
rect -13120 83380 -12880 83400
rect -12620 83380 -12380 83400
rect -12120 83380 -12000 83400
rect -16000 83350 -15900 83380
rect -16000 83150 -15980 83350
rect -15910 83150 -15900 83350
rect -16000 83120 -15900 83150
rect -15600 83350 -15400 83380
rect -15600 83150 -15590 83350
rect -15520 83150 -15480 83350
rect -15410 83150 -15400 83350
rect -15600 83120 -15400 83150
rect -15100 83350 -14900 83380
rect -15100 83150 -15090 83350
rect -15020 83150 -14980 83350
rect -14910 83150 -14900 83350
rect -15100 83120 -14900 83150
rect -14600 83350 -14400 83380
rect -14600 83150 -14590 83350
rect -14520 83150 -14480 83350
rect -14410 83150 -14400 83350
rect -14600 83120 -14400 83150
rect -14100 83350 -13900 83380
rect -14100 83150 -14090 83350
rect -14020 83150 -13980 83350
rect -13910 83150 -13900 83350
rect -14100 83120 -13900 83150
rect -13600 83350 -13400 83380
rect -13600 83150 -13590 83350
rect -13520 83150 -13480 83350
rect -13410 83150 -13400 83350
rect -13600 83120 -13400 83150
rect -13100 83350 -12900 83380
rect -13100 83150 -13090 83350
rect -13020 83150 -12980 83350
rect -12910 83150 -12900 83350
rect -13100 83120 -12900 83150
rect -12600 83350 -12400 83380
rect -12600 83150 -12590 83350
rect -12520 83150 -12480 83350
rect -12410 83150 -12400 83350
rect -12600 83120 -12400 83150
rect -12100 83350 -12000 83380
rect -12100 83150 -12090 83350
rect -12020 83150 -12000 83350
rect -12100 83120 -12000 83150
rect -16000 83100 -15880 83120
rect -15620 83100 -15380 83120
rect -15120 83100 -14880 83120
rect -14620 83100 -14380 83120
rect -14120 83100 -13880 83120
rect -13620 83100 -13380 83120
rect -13120 83100 -12880 83120
rect -12620 83100 -12380 83120
rect -12120 83100 -12000 83120
rect -16000 83090 -12000 83100
rect -16000 83020 -15850 83090
rect -15650 83020 -15350 83090
rect -15150 83020 -14850 83090
rect -14650 83020 -14350 83090
rect -14150 83020 -13850 83090
rect -13650 83020 -13350 83090
rect -13150 83020 -12850 83090
rect -12650 83020 -12350 83090
rect -12150 83020 -12000 83090
rect -16000 82980 -12000 83020
rect -16000 82910 -15850 82980
rect -15650 82910 -15350 82980
rect -15150 82910 -14850 82980
rect -14650 82910 -14350 82980
rect -14150 82910 -13850 82980
rect -13650 82910 -13350 82980
rect -13150 82910 -12850 82980
rect -12650 82910 -12350 82980
rect -12150 82910 -12000 82980
rect -16000 82900 -12000 82910
rect -16000 82880 -15880 82900
rect -15620 82880 -15380 82900
rect -15120 82880 -14880 82900
rect -14620 82880 -14380 82900
rect -14120 82880 -13880 82900
rect -13620 82880 -13380 82900
rect -13120 82880 -12880 82900
rect -12620 82880 -12380 82900
rect -12120 82880 -12000 82900
rect -16000 82850 -15900 82880
rect -16000 82650 -15980 82850
rect -15910 82650 -15900 82850
rect -16000 82620 -15900 82650
rect -15600 82850 -15400 82880
rect -15600 82650 -15590 82850
rect -15520 82650 -15480 82850
rect -15410 82650 -15400 82850
rect -15600 82620 -15400 82650
rect -15100 82850 -14900 82880
rect -15100 82650 -15090 82850
rect -15020 82650 -14980 82850
rect -14910 82650 -14900 82850
rect -15100 82620 -14900 82650
rect -14600 82850 -14400 82880
rect -14600 82650 -14590 82850
rect -14520 82650 -14480 82850
rect -14410 82650 -14400 82850
rect -14600 82620 -14400 82650
rect -14100 82850 -13900 82880
rect -14100 82650 -14090 82850
rect -14020 82650 -13980 82850
rect -13910 82650 -13900 82850
rect -14100 82620 -13900 82650
rect -13600 82850 -13400 82880
rect -13600 82650 -13590 82850
rect -13520 82650 -13480 82850
rect -13410 82650 -13400 82850
rect -13600 82620 -13400 82650
rect -13100 82850 -12900 82880
rect -13100 82650 -13090 82850
rect -13020 82650 -12980 82850
rect -12910 82650 -12900 82850
rect -13100 82620 -12900 82650
rect -12600 82850 -12400 82880
rect -12600 82650 -12590 82850
rect -12520 82650 -12480 82850
rect -12410 82650 -12400 82850
rect -12600 82620 -12400 82650
rect -12100 82850 -12000 82880
rect -12100 82650 -12090 82850
rect -12020 82650 -12000 82850
rect -12100 82620 -12000 82650
rect -16000 82600 -15880 82620
rect -15620 82600 -15380 82620
rect -15120 82600 -14880 82620
rect -14620 82600 -14380 82620
rect -14120 82600 -13880 82620
rect -13620 82600 -13380 82620
rect -13120 82600 -12880 82620
rect -12620 82600 -12380 82620
rect -12120 82600 -12000 82620
rect -16000 82590 -12000 82600
rect -16000 82520 -15850 82590
rect -15650 82520 -15350 82590
rect -15150 82520 -14850 82590
rect -14650 82520 -14350 82590
rect -14150 82520 -13850 82590
rect -13650 82520 -13350 82590
rect -13150 82520 -12850 82590
rect -12650 82520 -12350 82590
rect -12150 82520 -12000 82590
rect -16000 82480 -12000 82520
rect -16000 82410 -15850 82480
rect -15650 82410 -15350 82480
rect -15150 82410 -14850 82480
rect -14650 82410 -14350 82480
rect -14150 82410 -13850 82480
rect -13650 82410 -13350 82480
rect -13150 82410 -12850 82480
rect -12650 82410 -12350 82480
rect -12150 82410 -12000 82480
rect -16000 82400 -12000 82410
rect -16000 82380 -15880 82400
rect -15620 82380 -15380 82400
rect -15120 82380 -14880 82400
rect -14620 82380 -14380 82400
rect -14120 82380 -13880 82400
rect -13620 82380 -13380 82400
rect -13120 82380 -12880 82400
rect -12620 82380 -12380 82400
rect -12120 82380 -12000 82400
rect -16000 82350 -15900 82380
rect -16000 82150 -15980 82350
rect -15910 82150 -15900 82350
rect -16000 82120 -15900 82150
rect -15600 82350 -15400 82380
rect -15600 82150 -15590 82350
rect -15520 82150 -15480 82350
rect -15410 82150 -15400 82350
rect -15600 82120 -15400 82150
rect -15100 82350 -14900 82380
rect -15100 82150 -15090 82350
rect -15020 82150 -14980 82350
rect -14910 82150 -14900 82350
rect -15100 82120 -14900 82150
rect -14600 82350 -14400 82380
rect -14600 82150 -14590 82350
rect -14520 82150 -14480 82350
rect -14410 82150 -14400 82350
rect -14600 82120 -14400 82150
rect -14100 82350 -13900 82380
rect -14100 82150 -14090 82350
rect -14020 82150 -13980 82350
rect -13910 82150 -13900 82350
rect -14100 82120 -13900 82150
rect -13600 82350 -13400 82380
rect -13600 82150 -13590 82350
rect -13520 82150 -13480 82350
rect -13410 82150 -13400 82350
rect -13600 82120 -13400 82150
rect -13100 82350 -12900 82380
rect -13100 82150 -13090 82350
rect -13020 82150 -12980 82350
rect -12910 82150 -12900 82350
rect -13100 82120 -12900 82150
rect -12600 82350 -12400 82380
rect -12600 82150 -12590 82350
rect -12520 82150 -12480 82350
rect -12410 82150 -12400 82350
rect -12600 82120 -12400 82150
rect -12100 82350 -12000 82380
rect -12100 82150 -12090 82350
rect -12020 82150 -12000 82350
rect -12100 82120 -12000 82150
rect -16000 82100 -15880 82120
rect -15620 82100 -15380 82120
rect -15120 82100 -14880 82120
rect -14620 82100 -14380 82120
rect -14120 82100 -13880 82120
rect -13620 82100 -13380 82120
rect -13120 82100 -12880 82120
rect -12620 82100 -12380 82120
rect -12120 82100 -12000 82120
rect -16000 82090 -12000 82100
rect -16000 82020 -15850 82090
rect -15650 82020 -15350 82090
rect -15150 82020 -14850 82090
rect -14650 82020 -14350 82090
rect -14150 82020 -13850 82090
rect -13650 82020 -13350 82090
rect -13150 82020 -12850 82090
rect -12650 82020 -12350 82090
rect -12150 82020 -12000 82090
rect -16000 81980 -12000 82020
rect -16000 81910 -15850 81980
rect -15650 81910 -15350 81980
rect -15150 81910 -14850 81980
rect -14650 81910 -14350 81980
rect -14150 81910 -13850 81980
rect -13650 81910 -13350 81980
rect -13150 81910 -12850 81980
rect -12650 81910 -12350 81980
rect -12150 81910 -12000 81980
rect -16000 81900 -12000 81910
rect -16000 81880 -15880 81900
rect -15620 81880 -15380 81900
rect -15120 81880 -14880 81900
rect -14620 81880 -14380 81900
rect -14120 81880 -13880 81900
rect -13620 81880 -13380 81900
rect -13120 81880 -12880 81900
rect -12620 81880 -12380 81900
rect -12120 81880 -12000 81900
rect -16000 81850 -15900 81880
rect -16000 81650 -15980 81850
rect -15910 81650 -15900 81850
rect -16000 81620 -15900 81650
rect -15600 81850 -15400 81880
rect -15600 81650 -15590 81850
rect -15520 81650 -15480 81850
rect -15410 81650 -15400 81850
rect -15600 81620 -15400 81650
rect -15100 81850 -14900 81880
rect -15100 81650 -15090 81850
rect -15020 81650 -14980 81850
rect -14910 81650 -14900 81850
rect -15100 81620 -14900 81650
rect -14600 81850 -14400 81880
rect -14600 81650 -14590 81850
rect -14520 81650 -14480 81850
rect -14410 81650 -14400 81850
rect -14600 81620 -14400 81650
rect -14100 81850 -13900 81880
rect -14100 81650 -14090 81850
rect -14020 81650 -13980 81850
rect -13910 81650 -13900 81850
rect -14100 81620 -13900 81650
rect -13600 81850 -13400 81880
rect -13600 81650 -13590 81850
rect -13520 81650 -13480 81850
rect -13410 81650 -13400 81850
rect -13600 81620 -13400 81650
rect -13100 81850 -12900 81880
rect -13100 81650 -13090 81850
rect -13020 81650 -12980 81850
rect -12910 81650 -12900 81850
rect -13100 81620 -12900 81650
rect -12600 81850 -12400 81880
rect -12600 81650 -12590 81850
rect -12520 81650 -12480 81850
rect -12410 81650 -12400 81850
rect -12600 81620 -12400 81650
rect -12100 81850 -12000 81880
rect -12100 81650 -12090 81850
rect -12020 81650 -12000 81850
rect -12100 81620 -12000 81650
rect -16000 81600 -15880 81620
rect -15620 81600 -15380 81620
rect -15120 81600 -14880 81620
rect -14620 81600 -14380 81620
rect -14120 81600 -13880 81620
rect -13620 81600 -13380 81620
rect -13120 81600 -12880 81620
rect -12620 81600 -12380 81620
rect -12120 81600 -12000 81620
rect -16000 81590 -12000 81600
rect -16000 81520 -15850 81590
rect -15650 81520 -15350 81590
rect -15150 81520 -14850 81590
rect -14650 81520 -14350 81590
rect -14150 81520 -13850 81590
rect -13650 81520 -13350 81590
rect -13150 81520 -12850 81590
rect -12650 81520 -12350 81590
rect -12150 81520 -12000 81590
rect -16000 81480 -12000 81520
rect -16000 81410 -15850 81480
rect -15650 81410 -15350 81480
rect -15150 81410 -14850 81480
rect -14650 81410 -14350 81480
rect -14150 81410 -13850 81480
rect -13650 81410 -13350 81480
rect -13150 81410 -12850 81480
rect -12650 81410 -12350 81480
rect -12150 81410 -12000 81480
rect -16000 81400 -12000 81410
rect -16000 81380 -15880 81400
rect -15620 81380 -15380 81400
rect -15120 81380 -14880 81400
rect -14620 81380 -14380 81400
rect -14120 81380 -13880 81400
rect -13620 81380 -13380 81400
rect -13120 81380 -12880 81400
rect -12620 81380 -12380 81400
rect -12120 81380 -12000 81400
rect -16000 81350 -15900 81380
rect -16000 81150 -15980 81350
rect -15910 81150 -15900 81350
rect -16000 81120 -15900 81150
rect -15600 81350 -15400 81380
rect -15600 81150 -15590 81350
rect -15520 81150 -15480 81350
rect -15410 81150 -15400 81350
rect -15600 81120 -15400 81150
rect -15100 81350 -14900 81380
rect -15100 81150 -15090 81350
rect -15020 81150 -14980 81350
rect -14910 81150 -14900 81350
rect -15100 81120 -14900 81150
rect -14600 81350 -14400 81380
rect -14600 81150 -14590 81350
rect -14520 81150 -14480 81350
rect -14410 81150 -14400 81350
rect -14600 81120 -14400 81150
rect -14100 81350 -13900 81380
rect -14100 81150 -14090 81350
rect -14020 81150 -13980 81350
rect -13910 81150 -13900 81350
rect -14100 81120 -13900 81150
rect -13600 81350 -13400 81380
rect -13600 81150 -13590 81350
rect -13520 81150 -13480 81350
rect -13410 81150 -13400 81350
rect -13600 81120 -13400 81150
rect -13100 81350 -12900 81380
rect -13100 81150 -13090 81350
rect -13020 81150 -12980 81350
rect -12910 81150 -12900 81350
rect -13100 81120 -12900 81150
rect -12600 81350 -12400 81380
rect -12600 81150 -12590 81350
rect -12520 81150 -12480 81350
rect -12410 81150 -12400 81350
rect -12600 81120 -12400 81150
rect -12100 81350 -12000 81380
rect -12100 81150 -12090 81350
rect -12020 81150 -12000 81350
rect -12100 81120 -12000 81150
rect -16000 81100 -15880 81120
rect -15620 81100 -15380 81120
rect -15120 81100 -14880 81120
rect -14620 81100 -14380 81120
rect -14120 81100 -13880 81120
rect -13620 81100 -13380 81120
rect -13120 81100 -12880 81120
rect -12620 81100 -12380 81120
rect -12120 81100 -12000 81120
rect -16000 81090 -12000 81100
rect -16000 81020 -15850 81090
rect -15650 81020 -15350 81090
rect -15150 81020 -14850 81090
rect -14650 81020 -14350 81090
rect -14150 81020 -13850 81090
rect -13650 81020 -13350 81090
rect -13150 81020 -12850 81090
rect -12650 81020 -12350 81090
rect -12150 81020 -12000 81090
rect -16000 80980 -12000 81020
rect -16000 80910 -15850 80980
rect -15650 80910 -15350 80980
rect -15150 80910 -14850 80980
rect -14650 80910 -14350 80980
rect -14150 80910 -13850 80980
rect -13650 80910 -13350 80980
rect -13150 80910 -12850 80980
rect -12650 80910 -12350 80980
rect -12150 80910 -12000 80980
rect -16000 80900 -12000 80910
rect -16000 80880 -15880 80900
rect -15620 80880 -15380 80900
rect -15120 80880 -14880 80900
rect -14620 80880 -14380 80900
rect -14120 80880 -13880 80900
rect -13620 80880 -13380 80900
rect -13120 80880 -12880 80900
rect -12620 80880 -12380 80900
rect -12120 80880 -12000 80900
rect -16000 80850 -15900 80880
rect -16000 80650 -15980 80850
rect -15910 80650 -15900 80850
rect -16000 80620 -15900 80650
rect -15600 80850 -15400 80880
rect -15600 80650 -15590 80850
rect -15520 80650 -15480 80850
rect -15410 80650 -15400 80850
rect -15600 80620 -15400 80650
rect -15100 80850 -14900 80880
rect -15100 80650 -15090 80850
rect -15020 80650 -14980 80850
rect -14910 80650 -14900 80850
rect -15100 80620 -14900 80650
rect -14600 80850 -14400 80880
rect -14600 80650 -14590 80850
rect -14520 80650 -14480 80850
rect -14410 80650 -14400 80850
rect -14600 80620 -14400 80650
rect -14100 80850 -13900 80880
rect -14100 80650 -14090 80850
rect -14020 80650 -13980 80850
rect -13910 80650 -13900 80850
rect -14100 80620 -13900 80650
rect -13600 80850 -13400 80880
rect -13600 80650 -13590 80850
rect -13520 80650 -13480 80850
rect -13410 80650 -13400 80850
rect -13600 80620 -13400 80650
rect -13100 80850 -12900 80880
rect -13100 80650 -13090 80850
rect -13020 80650 -12980 80850
rect -12910 80650 -12900 80850
rect -13100 80620 -12900 80650
rect -12600 80850 -12400 80880
rect -12600 80650 -12590 80850
rect -12520 80650 -12480 80850
rect -12410 80650 -12400 80850
rect -12600 80620 -12400 80650
rect -12100 80850 -12000 80880
rect -12100 80650 -12090 80850
rect -12020 80650 -12000 80850
rect -12100 80620 -12000 80650
rect -16000 80600 -15880 80620
rect -15620 80600 -15380 80620
rect -15120 80600 -14880 80620
rect -14620 80600 -14380 80620
rect -14120 80600 -13880 80620
rect -13620 80600 -13380 80620
rect -13120 80600 -12880 80620
rect -12620 80600 -12380 80620
rect -12120 80600 -12000 80620
rect -16000 80590 -12000 80600
rect -16000 80520 -15850 80590
rect -15650 80520 -15350 80590
rect -15150 80520 -14850 80590
rect -14650 80520 -14350 80590
rect -14150 80520 -13850 80590
rect -13650 80520 -13350 80590
rect -13150 80520 -12850 80590
rect -12650 80520 -12350 80590
rect -12150 80520 -12000 80590
rect -16000 80480 -12000 80520
rect -16000 80410 -15850 80480
rect -15650 80410 -15350 80480
rect -15150 80410 -14850 80480
rect -14650 80410 -14350 80480
rect -14150 80410 -13850 80480
rect -13650 80410 -13350 80480
rect -13150 80410 -12850 80480
rect -12650 80410 -12350 80480
rect -12150 80410 -12000 80480
rect -16000 80400 -12000 80410
rect -16000 80380 -15880 80400
rect -15620 80380 -15380 80400
rect -15120 80380 -14880 80400
rect -14620 80380 -14380 80400
rect -14120 80380 -13880 80400
rect -13620 80380 -13380 80400
rect -13120 80380 -12880 80400
rect -12620 80380 -12380 80400
rect -12120 80380 -12000 80400
rect -16000 80350 -15900 80380
rect -16000 80150 -15980 80350
rect -15910 80150 -15900 80350
rect -16000 80120 -15900 80150
rect -15600 80350 -15400 80380
rect -15600 80150 -15590 80350
rect -15520 80150 -15480 80350
rect -15410 80150 -15400 80350
rect -15600 80120 -15400 80150
rect -15100 80350 -14900 80380
rect -15100 80150 -15090 80350
rect -15020 80150 -14980 80350
rect -14910 80150 -14900 80350
rect -15100 80120 -14900 80150
rect -14600 80350 -14400 80380
rect -14600 80150 -14590 80350
rect -14520 80150 -14480 80350
rect -14410 80150 -14400 80350
rect -14600 80120 -14400 80150
rect -14100 80350 -13900 80380
rect -14100 80150 -14090 80350
rect -14020 80150 -13980 80350
rect -13910 80150 -13900 80350
rect -14100 80120 -13900 80150
rect -13600 80350 -13400 80380
rect -13600 80150 -13590 80350
rect -13520 80150 -13480 80350
rect -13410 80150 -13400 80350
rect -13600 80120 -13400 80150
rect -13100 80350 -12900 80380
rect -13100 80150 -13090 80350
rect -13020 80150 -12980 80350
rect -12910 80150 -12900 80350
rect -13100 80120 -12900 80150
rect -12600 80350 -12400 80380
rect -12600 80150 -12590 80350
rect -12520 80150 -12480 80350
rect -12410 80150 -12400 80350
rect -12600 80120 -12400 80150
rect -12100 80350 -12000 80380
rect -12100 80150 -12090 80350
rect -12020 80150 -12000 80350
rect -12100 80120 -12000 80150
rect -16000 80100 -15880 80120
rect -15620 80100 -15380 80120
rect -15120 80100 -14880 80120
rect -14620 80100 -14380 80120
rect -14120 80100 -13880 80120
rect -13620 80100 -13380 80120
rect -13120 80100 -12880 80120
rect -12620 80100 -12380 80120
rect -12120 80100 -12000 80120
rect -16000 80090 -12000 80100
rect -16000 80020 -15850 80090
rect -15650 80020 -15350 80090
rect -15150 80020 -14850 80090
rect -14650 80020 -14350 80090
rect -14150 80020 -13850 80090
rect -13650 80020 -13350 80090
rect -13150 80020 -12850 80090
rect -12650 80020 -12350 80090
rect -12150 80020 -12000 80090
rect -16000 79980 -12000 80020
rect -16000 79910 -15850 79980
rect -15650 79910 -15350 79980
rect -15150 79910 -14850 79980
rect -14650 79910 -14350 79980
rect -14150 79910 -13850 79980
rect -13650 79910 -13350 79980
rect -13150 79910 -12850 79980
rect -12650 79910 -12350 79980
rect -12150 79910 -12000 79980
rect -16000 79900 -12000 79910
rect -16000 79880 -15880 79900
rect -15620 79880 -15380 79900
rect -15120 79880 -14880 79900
rect -14620 79880 -14380 79900
rect -14120 79880 -13880 79900
rect -13620 79880 -13380 79900
rect -13120 79880 -12880 79900
rect -12620 79880 -12380 79900
rect -12120 79880 -12000 79900
rect -16000 79850 -15900 79880
rect -16000 79650 -15980 79850
rect -15910 79650 -15900 79850
rect -16000 79620 -15900 79650
rect -15600 79850 -15400 79880
rect -15600 79650 -15590 79850
rect -15520 79650 -15480 79850
rect -15410 79650 -15400 79850
rect -15600 79620 -15400 79650
rect -15100 79850 -14900 79880
rect -15100 79650 -15090 79850
rect -15020 79650 -14980 79850
rect -14910 79650 -14900 79850
rect -15100 79620 -14900 79650
rect -14600 79850 -14400 79880
rect -14600 79650 -14590 79850
rect -14520 79650 -14480 79850
rect -14410 79650 -14400 79850
rect -14600 79620 -14400 79650
rect -14100 79850 -13900 79880
rect -14100 79650 -14090 79850
rect -14020 79650 -13980 79850
rect -13910 79650 -13900 79850
rect -14100 79620 -13900 79650
rect -13600 79850 -13400 79880
rect -13600 79650 -13590 79850
rect -13520 79650 -13480 79850
rect -13410 79650 -13400 79850
rect -13600 79620 -13400 79650
rect -13100 79850 -12900 79880
rect -13100 79650 -13090 79850
rect -13020 79650 -12980 79850
rect -12910 79650 -12900 79850
rect -13100 79620 -12900 79650
rect -12600 79850 -12400 79880
rect -12600 79650 -12590 79850
rect -12520 79650 -12480 79850
rect -12410 79650 -12400 79850
rect -12600 79620 -12400 79650
rect -12100 79850 -12000 79880
rect -12100 79650 -12090 79850
rect -12020 79650 -12000 79850
rect -12100 79620 -12000 79650
rect -16000 79600 -15880 79620
rect -15620 79600 -15380 79620
rect -15120 79600 -14880 79620
rect -14620 79600 -14380 79620
rect -14120 79600 -13880 79620
rect -13620 79600 -13380 79620
rect -13120 79600 -12880 79620
rect -12620 79600 -12380 79620
rect -12120 79600 -12000 79620
rect -16000 79590 -12000 79600
rect -16000 79520 -15850 79590
rect -15650 79520 -15350 79590
rect -15150 79520 -14850 79590
rect -14650 79520 -14350 79590
rect -14150 79520 -13850 79590
rect -13650 79520 -13350 79590
rect -13150 79520 -12850 79590
rect -12650 79520 -12350 79590
rect -12150 79520 -12000 79590
rect -16000 79480 -12000 79520
rect -16000 79410 -15850 79480
rect -15650 79410 -15350 79480
rect -15150 79410 -14850 79480
rect -14650 79410 -14350 79480
rect -14150 79410 -13850 79480
rect -13650 79410 -13350 79480
rect -13150 79410 -12850 79480
rect -12650 79410 -12350 79480
rect -12150 79410 -12000 79480
rect -16000 79400 -12000 79410
rect -16000 79380 -15880 79400
rect -15620 79380 -15380 79400
rect -15120 79380 -14880 79400
rect -14620 79380 -14380 79400
rect -14120 79380 -13880 79400
rect -13620 79380 -13380 79400
rect -13120 79380 -12880 79400
rect -12620 79380 -12380 79400
rect -12120 79380 -12000 79400
rect -16000 79350 -15900 79380
rect -16000 79150 -15980 79350
rect -15910 79150 -15900 79350
rect -16000 79120 -15900 79150
rect -15600 79350 -15400 79380
rect -15600 79150 -15590 79350
rect -15520 79150 -15480 79350
rect -15410 79150 -15400 79350
rect -15600 79120 -15400 79150
rect -15100 79350 -14900 79380
rect -15100 79150 -15090 79350
rect -15020 79150 -14980 79350
rect -14910 79150 -14900 79350
rect -15100 79120 -14900 79150
rect -14600 79350 -14400 79380
rect -14600 79150 -14590 79350
rect -14520 79150 -14480 79350
rect -14410 79150 -14400 79350
rect -14600 79120 -14400 79150
rect -14100 79350 -13900 79380
rect -14100 79150 -14090 79350
rect -14020 79150 -13980 79350
rect -13910 79150 -13900 79350
rect -14100 79120 -13900 79150
rect -13600 79350 -13400 79380
rect -13600 79150 -13590 79350
rect -13520 79150 -13480 79350
rect -13410 79150 -13400 79350
rect -13600 79120 -13400 79150
rect -13100 79350 -12900 79380
rect -13100 79150 -13090 79350
rect -13020 79150 -12980 79350
rect -12910 79150 -12900 79350
rect -13100 79120 -12900 79150
rect -12600 79350 -12400 79380
rect -12600 79150 -12590 79350
rect -12520 79150 -12480 79350
rect -12410 79150 -12400 79350
rect -12600 79120 -12400 79150
rect -12100 79350 -12000 79380
rect -12100 79150 -12090 79350
rect -12020 79150 -12000 79350
rect -12100 79120 -12000 79150
rect -16000 79100 -15880 79120
rect -15620 79100 -15380 79120
rect -15120 79100 -14880 79120
rect -14620 79100 -14380 79120
rect -14120 79100 -13880 79120
rect -13620 79100 -13380 79120
rect -13120 79100 -12880 79120
rect -12620 79100 -12380 79120
rect -12120 79100 -12000 79120
rect -16000 79090 -12000 79100
rect -16000 79020 -15850 79090
rect -15650 79020 -15350 79090
rect -15150 79020 -14850 79090
rect -14650 79020 -14350 79090
rect -14150 79020 -13850 79090
rect -13650 79020 -13350 79090
rect -13150 79020 -12850 79090
rect -12650 79020 -12350 79090
rect -12150 79020 -12000 79090
rect -16000 78980 -12000 79020
rect -16000 78910 -15850 78980
rect -15650 78910 -15350 78980
rect -15150 78910 -14850 78980
rect -14650 78910 -14350 78980
rect -14150 78910 -13850 78980
rect -13650 78910 -13350 78980
rect -13150 78910 -12850 78980
rect -12650 78910 -12350 78980
rect -12150 78910 -12000 78980
rect -16000 78900 -12000 78910
rect -16000 78880 -15880 78900
rect -15620 78880 -15380 78900
rect -15120 78880 -14880 78900
rect -14620 78880 -14380 78900
rect -14120 78880 -13880 78900
rect -13620 78880 -13380 78900
rect -13120 78880 -12880 78900
rect -12620 78880 -12380 78900
rect -12120 78880 -12000 78900
rect -16000 78850 -15900 78880
rect -16000 78650 -15980 78850
rect -15910 78650 -15900 78850
rect -16000 78620 -15900 78650
rect -15600 78850 -15400 78880
rect -15600 78650 -15590 78850
rect -15520 78650 -15480 78850
rect -15410 78650 -15400 78850
rect -15600 78620 -15400 78650
rect -15100 78850 -14900 78880
rect -15100 78650 -15090 78850
rect -15020 78650 -14980 78850
rect -14910 78650 -14900 78850
rect -15100 78620 -14900 78650
rect -14600 78850 -14400 78880
rect -14600 78650 -14590 78850
rect -14520 78650 -14480 78850
rect -14410 78650 -14400 78850
rect -14600 78620 -14400 78650
rect -14100 78850 -13900 78880
rect -14100 78650 -14090 78850
rect -14020 78650 -13980 78850
rect -13910 78650 -13900 78850
rect -14100 78620 -13900 78650
rect -13600 78850 -13400 78880
rect -13600 78650 -13590 78850
rect -13520 78650 -13480 78850
rect -13410 78650 -13400 78850
rect -13600 78620 -13400 78650
rect -13100 78850 -12900 78880
rect -13100 78650 -13090 78850
rect -13020 78650 -12980 78850
rect -12910 78650 -12900 78850
rect -13100 78620 -12900 78650
rect -12600 78850 -12400 78880
rect -12600 78650 -12590 78850
rect -12520 78650 -12480 78850
rect -12410 78650 -12400 78850
rect -12600 78620 -12400 78650
rect -12100 78850 -12000 78880
rect -12100 78650 -12090 78850
rect -12020 78650 -12000 78850
rect -12100 78620 -12000 78650
rect -16000 78600 -15880 78620
rect -15620 78600 -15380 78620
rect -15120 78600 -14880 78620
rect -14620 78600 -14380 78620
rect -14120 78600 -13880 78620
rect -13620 78600 -13380 78620
rect -13120 78600 -12880 78620
rect -12620 78600 -12380 78620
rect -12120 78600 -12000 78620
rect -16000 78590 -12000 78600
rect -16000 78520 -15850 78590
rect -15650 78520 -15350 78590
rect -15150 78520 -14850 78590
rect -14650 78520 -14350 78590
rect -14150 78520 -13850 78590
rect -13650 78520 -13350 78590
rect -13150 78520 -12850 78590
rect -12650 78520 -12350 78590
rect -12150 78520 -12000 78590
rect -16000 78480 -12000 78520
rect -16000 78410 -15850 78480
rect -15650 78410 -15350 78480
rect -15150 78410 -14850 78480
rect -14650 78410 -14350 78480
rect -14150 78410 -13850 78480
rect -13650 78410 -13350 78480
rect -13150 78410 -12850 78480
rect -12650 78410 -12350 78480
rect -12150 78410 -12000 78480
rect -16000 78400 -12000 78410
rect -16000 78380 -15880 78400
rect -15620 78380 -15380 78400
rect -15120 78380 -14880 78400
rect -14620 78380 -14380 78400
rect -14120 78380 -13880 78400
rect -13620 78380 -13380 78400
rect -13120 78380 -12880 78400
rect -12620 78380 -12380 78400
rect -12120 78380 -12000 78400
rect -16000 78350 -15900 78380
rect -16000 78150 -15980 78350
rect -15910 78150 -15900 78350
rect -16000 78120 -15900 78150
rect -15600 78350 -15400 78380
rect -15600 78150 -15590 78350
rect -15520 78150 -15480 78350
rect -15410 78150 -15400 78350
rect -15600 78120 -15400 78150
rect -15100 78350 -14900 78380
rect -15100 78150 -15090 78350
rect -15020 78150 -14980 78350
rect -14910 78150 -14900 78350
rect -15100 78120 -14900 78150
rect -14600 78350 -14400 78380
rect -14600 78150 -14590 78350
rect -14520 78150 -14480 78350
rect -14410 78150 -14400 78350
rect -14600 78120 -14400 78150
rect -14100 78350 -13900 78380
rect -14100 78150 -14090 78350
rect -14020 78150 -13980 78350
rect -13910 78150 -13900 78350
rect -14100 78120 -13900 78150
rect -13600 78350 -13400 78380
rect -13600 78150 -13590 78350
rect -13520 78150 -13480 78350
rect -13410 78150 -13400 78350
rect -13600 78120 -13400 78150
rect -13100 78350 -12900 78380
rect -13100 78150 -13090 78350
rect -13020 78150 -12980 78350
rect -12910 78150 -12900 78350
rect -13100 78120 -12900 78150
rect -12600 78350 -12400 78380
rect -12600 78150 -12590 78350
rect -12520 78150 -12480 78350
rect -12410 78150 -12400 78350
rect -12600 78120 -12400 78150
rect -12100 78350 -12000 78380
rect -12100 78150 -12090 78350
rect -12020 78150 -12000 78350
rect -12100 78120 -12000 78150
rect -16000 78100 -15880 78120
rect -15620 78100 -15380 78120
rect -15120 78100 -14880 78120
rect -14620 78100 -14380 78120
rect -14120 78100 -13880 78120
rect -13620 78100 -13380 78120
rect -13120 78100 -12880 78120
rect -12620 78100 -12380 78120
rect -12120 78100 -12000 78120
rect -16000 78090 -12000 78100
rect -16000 78020 -15850 78090
rect -15650 78020 -15350 78090
rect -15150 78020 -14850 78090
rect -14650 78020 -14350 78090
rect -14150 78020 -13850 78090
rect -13650 78020 -13350 78090
rect -13150 78020 -12850 78090
rect -12650 78020 -12350 78090
rect -12150 78020 -12000 78090
rect -16000 77980 -12000 78020
rect -16000 77910 -15850 77980
rect -15650 77910 -15350 77980
rect -15150 77910 -14850 77980
rect -14650 77910 -14350 77980
rect -14150 77910 -13850 77980
rect -13650 77910 -13350 77980
rect -13150 77910 -12850 77980
rect -12650 77910 -12350 77980
rect -12150 77910 -12000 77980
rect -16000 77900 -12000 77910
rect -16000 77880 -15880 77900
rect -15620 77880 -15380 77900
rect -15120 77880 -14880 77900
rect -14620 77880 -14380 77900
rect -14120 77880 -13880 77900
rect -13620 77880 -13380 77900
rect -13120 77880 -12880 77900
rect -12620 77880 -12380 77900
rect -12120 77880 -12000 77900
rect -16000 77850 -15900 77880
rect -16000 77650 -15980 77850
rect -15910 77650 -15900 77850
rect -16000 77620 -15900 77650
rect -15600 77850 -15400 77880
rect -15600 77650 -15590 77850
rect -15520 77650 -15480 77850
rect -15410 77650 -15400 77850
rect -15600 77620 -15400 77650
rect -15100 77850 -14900 77880
rect -15100 77650 -15090 77850
rect -15020 77650 -14980 77850
rect -14910 77650 -14900 77850
rect -15100 77620 -14900 77650
rect -14600 77850 -14400 77880
rect -14600 77650 -14590 77850
rect -14520 77650 -14480 77850
rect -14410 77650 -14400 77850
rect -14600 77620 -14400 77650
rect -14100 77850 -13900 77880
rect -14100 77650 -14090 77850
rect -14020 77650 -13980 77850
rect -13910 77650 -13900 77850
rect -14100 77620 -13900 77650
rect -13600 77850 -13400 77880
rect -13600 77650 -13590 77850
rect -13520 77650 -13480 77850
rect -13410 77650 -13400 77850
rect -13600 77620 -13400 77650
rect -13100 77850 -12900 77880
rect -13100 77650 -13090 77850
rect -13020 77650 -12980 77850
rect -12910 77650 -12900 77850
rect -13100 77620 -12900 77650
rect -12600 77850 -12400 77880
rect -12600 77650 -12590 77850
rect -12520 77650 -12480 77850
rect -12410 77650 -12400 77850
rect -12600 77620 -12400 77650
rect -12100 77850 -12000 77880
rect -12100 77650 -12090 77850
rect -12020 77650 -12000 77850
rect -12100 77620 -12000 77650
rect -16000 77600 -15880 77620
rect -15620 77600 -15380 77620
rect -15120 77600 -14880 77620
rect -14620 77600 -14380 77620
rect -14120 77600 -13880 77620
rect -13620 77600 -13380 77620
rect -13120 77600 -12880 77620
rect -12620 77600 -12380 77620
rect -12120 77600 -12000 77620
rect -16000 77590 -12000 77600
rect -16000 77520 -15850 77590
rect -15650 77520 -15350 77590
rect -15150 77520 -14850 77590
rect -14650 77520 -14350 77590
rect -14150 77520 -13850 77590
rect -13650 77520 -13350 77590
rect -13150 77520 -12850 77590
rect -12650 77520 -12350 77590
rect -12150 77520 -12000 77590
rect -16000 77480 -12000 77520
rect -16000 77410 -15850 77480
rect -15650 77410 -15350 77480
rect -15150 77410 -14850 77480
rect -14650 77410 -14350 77480
rect -14150 77410 -13850 77480
rect -13650 77410 -13350 77480
rect -13150 77410 -12850 77480
rect -12650 77410 -12350 77480
rect -12150 77410 -12000 77480
rect -16000 77400 -12000 77410
rect -16000 77380 -15880 77400
rect -15620 77380 -15380 77400
rect -15120 77380 -14880 77400
rect -14620 77380 -14380 77400
rect -14120 77380 -13880 77400
rect -13620 77380 -13380 77400
rect -13120 77380 -12880 77400
rect -12620 77380 -12380 77400
rect -12120 77380 -12000 77400
rect -16000 77350 -15900 77380
rect -16000 77150 -15980 77350
rect -15910 77150 -15900 77350
rect -16000 77120 -15900 77150
rect -15600 77350 -15400 77380
rect -15600 77150 -15590 77350
rect -15520 77150 -15480 77350
rect -15410 77150 -15400 77350
rect -15600 77120 -15400 77150
rect -15100 77350 -14900 77380
rect -15100 77150 -15090 77350
rect -15020 77150 -14980 77350
rect -14910 77150 -14900 77350
rect -15100 77120 -14900 77150
rect -14600 77350 -14400 77380
rect -14600 77150 -14590 77350
rect -14520 77150 -14480 77350
rect -14410 77150 -14400 77350
rect -14600 77120 -14400 77150
rect -14100 77350 -13900 77380
rect -14100 77150 -14090 77350
rect -14020 77150 -13980 77350
rect -13910 77150 -13900 77350
rect -14100 77120 -13900 77150
rect -13600 77350 -13400 77380
rect -13600 77150 -13590 77350
rect -13520 77150 -13480 77350
rect -13410 77150 -13400 77350
rect -13600 77120 -13400 77150
rect -13100 77350 -12900 77380
rect -13100 77150 -13090 77350
rect -13020 77150 -12980 77350
rect -12910 77150 -12900 77350
rect -13100 77120 -12900 77150
rect -12600 77350 -12400 77380
rect -12600 77150 -12590 77350
rect -12520 77150 -12480 77350
rect -12410 77150 -12400 77350
rect -12600 77120 -12400 77150
rect -12100 77350 -12000 77380
rect -12100 77150 -12090 77350
rect -12020 77150 -12000 77350
rect -12100 77120 -12000 77150
rect -16000 77100 -15880 77120
rect -15620 77100 -15380 77120
rect -15120 77100 -14880 77120
rect -14620 77100 -14380 77120
rect -14120 77100 -13880 77120
rect -13620 77100 -13380 77120
rect -13120 77100 -12880 77120
rect -12620 77100 -12380 77120
rect -12120 77100 -12000 77120
rect -16000 77090 -12000 77100
rect -16000 77020 -15850 77090
rect -15650 77020 -15350 77090
rect -15150 77020 -14850 77090
rect -14650 77020 -14350 77090
rect -14150 77020 -13850 77090
rect -13650 77020 -13350 77090
rect -13150 77020 -12850 77090
rect -12650 77020 -12350 77090
rect -12150 77020 -12000 77090
rect -16000 76980 -12000 77020
rect -16000 76910 -15850 76980
rect -15650 76910 -15350 76980
rect -15150 76910 -14850 76980
rect -14650 76910 -14350 76980
rect -14150 76910 -13850 76980
rect -13650 76910 -13350 76980
rect -13150 76910 -12850 76980
rect -12650 76910 -12350 76980
rect -12150 76910 -12000 76980
rect -16000 76900 -12000 76910
rect -16000 76880 -15880 76900
rect -15620 76880 -15380 76900
rect -15120 76880 -14880 76900
rect -14620 76880 -14380 76900
rect -14120 76880 -13880 76900
rect -13620 76880 -13380 76900
rect -13120 76880 -12880 76900
rect -12620 76880 -12380 76900
rect -12120 76880 -12000 76900
rect -16000 76850 -15900 76880
rect -16000 76650 -15980 76850
rect -15910 76650 -15900 76850
rect -16000 76620 -15900 76650
rect -15600 76850 -15400 76880
rect -15600 76650 -15590 76850
rect -15520 76650 -15480 76850
rect -15410 76650 -15400 76850
rect -15600 76620 -15400 76650
rect -15100 76850 -14900 76880
rect -15100 76650 -15090 76850
rect -15020 76650 -14980 76850
rect -14910 76650 -14900 76850
rect -15100 76620 -14900 76650
rect -14600 76850 -14400 76880
rect -14600 76650 -14590 76850
rect -14520 76650 -14480 76850
rect -14410 76650 -14400 76850
rect -14600 76620 -14400 76650
rect -14100 76850 -13900 76880
rect -14100 76650 -14090 76850
rect -14020 76650 -13980 76850
rect -13910 76650 -13900 76850
rect -14100 76620 -13900 76650
rect -13600 76850 -13400 76880
rect -13600 76650 -13590 76850
rect -13520 76650 -13480 76850
rect -13410 76650 -13400 76850
rect -13600 76620 -13400 76650
rect -13100 76850 -12900 76880
rect -13100 76650 -13090 76850
rect -13020 76650 -12980 76850
rect -12910 76650 -12900 76850
rect -13100 76620 -12900 76650
rect -12600 76850 -12400 76880
rect -12600 76650 -12590 76850
rect -12520 76650 -12480 76850
rect -12410 76650 -12400 76850
rect -12600 76620 -12400 76650
rect -12100 76850 -12000 76880
rect -12100 76650 -12090 76850
rect -12020 76650 -12000 76850
rect -12100 76620 -12000 76650
rect -16000 76600 -15880 76620
rect -15620 76600 -15380 76620
rect -15120 76600 -14880 76620
rect -14620 76600 -14380 76620
rect -14120 76600 -13880 76620
rect -13620 76600 -13380 76620
rect -13120 76600 -12880 76620
rect -12620 76600 -12380 76620
rect -12120 76600 -12000 76620
rect -16000 76590 -12000 76600
rect -16000 76520 -15850 76590
rect -15650 76520 -15350 76590
rect -15150 76520 -14850 76590
rect -14650 76520 -14350 76590
rect -14150 76520 -13850 76590
rect -13650 76520 -13350 76590
rect -13150 76520 -12850 76590
rect -12650 76520 -12350 76590
rect -12150 76520 -12000 76590
rect -16000 76480 -12000 76520
rect -16000 76410 -15850 76480
rect -15650 76410 -15350 76480
rect -15150 76410 -14850 76480
rect -14650 76410 -14350 76480
rect -14150 76410 -13850 76480
rect -13650 76410 -13350 76480
rect -13150 76410 -12850 76480
rect -12650 76410 -12350 76480
rect -12150 76410 -12000 76480
rect -16000 76400 -12000 76410
rect -16000 76380 -15880 76400
rect -15620 76380 -15380 76400
rect -15120 76380 -14880 76400
rect -14620 76380 -14380 76400
rect -14120 76380 -13880 76400
rect -13620 76380 -13380 76400
rect -13120 76380 -12880 76400
rect -12620 76380 -12380 76400
rect -12120 76380 -12000 76400
rect -16000 76350 -15900 76380
rect -16000 76150 -15980 76350
rect -15910 76150 -15900 76350
rect -16000 76120 -15900 76150
rect -15600 76350 -15400 76380
rect -15600 76150 -15590 76350
rect -15520 76150 -15480 76350
rect -15410 76150 -15400 76350
rect -15600 76120 -15400 76150
rect -15100 76350 -14900 76380
rect -15100 76150 -15090 76350
rect -15020 76150 -14980 76350
rect -14910 76150 -14900 76350
rect -15100 76120 -14900 76150
rect -14600 76350 -14400 76380
rect -14600 76150 -14590 76350
rect -14520 76150 -14480 76350
rect -14410 76150 -14400 76350
rect -14600 76120 -14400 76150
rect -14100 76350 -13900 76380
rect -14100 76150 -14090 76350
rect -14020 76150 -13980 76350
rect -13910 76150 -13900 76350
rect -14100 76120 -13900 76150
rect -13600 76350 -13400 76380
rect -13600 76150 -13590 76350
rect -13520 76150 -13480 76350
rect -13410 76150 -13400 76350
rect -13600 76120 -13400 76150
rect -13100 76350 -12900 76380
rect -13100 76150 -13090 76350
rect -13020 76150 -12980 76350
rect -12910 76150 -12900 76350
rect -13100 76120 -12900 76150
rect -12600 76350 -12400 76380
rect -12600 76150 -12590 76350
rect -12520 76150 -12480 76350
rect -12410 76150 -12400 76350
rect -12600 76120 -12400 76150
rect -12100 76350 -12000 76380
rect -12100 76150 -12090 76350
rect -12020 76150 -12000 76350
rect -12100 76120 -12000 76150
rect -16000 76100 -15880 76120
rect -15620 76100 -15380 76120
rect -15120 76100 -14880 76120
rect -14620 76100 -14380 76120
rect -14120 76100 -13880 76120
rect -13620 76100 -13380 76120
rect -13120 76100 -12880 76120
rect -12620 76100 -12380 76120
rect -12120 76100 -12000 76120
rect -16000 76090 -12000 76100
rect -16000 76020 -15850 76090
rect -15650 76020 -15350 76090
rect -15150 76020 -14850 76090
rect -14650 76020 -14350 76090
rect -14150 76020 -13850 76090
rect -13650 76020 -13350 76090
rect -13150 76020 -12850 76090
rect -12650 76020 -12350 76090
rect -12150 76020 -12000 76090
rect -16000 75980 -12000 76020
rect -16000 75910 -15850 75980
rect -15650 75910 -15350 75980
rect -15150 75910 -14850 75980
rect -14650 75910 -14350 75980
rect -14150 75910 -13850 75980
rect -13650 75910 -13350 75980
rect -13150 75910 -12850 75980
rect -12650 75910 -12350 75980
rect -12150 75910 -12000 75980
rect -16000 75900 -12000 75910
rect -16000 75880 -15880 75900
rect -15620 75880 -15380 75900
rect -15120 75880 -14880 75900
rect -14620 75880 -14380 75900
rect -14120 75880 -13880 75900
rect -13620 75880 -13380 75900
rect -13120 75880 -12880 75900
rect -12620 75880 -12380 75900
rect -12120 75880 -12000 75900
rect -16000 75850 -15900 75880
rect -16000 75650 -15980 75850
rect -15910 75650 -15900 75850
rect -16000 75620 -15900 75650
rect -15600 75850 -15400 75880
rect -15600 75650 -15590 75850
rect -15520 75650 -15480 75850
rect -15410 75650 -15400 75850
rect -15600 75620 -15400 75650
rect -15100 75850 -14900 75880
rect -15100 75650 -15090 75850
rect -15020 75650 -14980 75850
rect -14910 75650 -14900 75850
rect -15100 75620 -14900 75650
rect -14600 75850 -14400 75880
rect -14600 75650 -14590 75850
rect -14520 75650 -14480 75850
rect -14410 75650 -14400 75850
rect -14600 75620 -14400 75650
rect -14100 75850 -13900 75880
rect -14100 75650 -14090 75850
rect -14020 75650 -13980 75850
rect -13910 75650 -13900 75850
rect -14100 75620 -13900 75650
rect -13600 75850 -13400 75880
rect -13600 75650 -13590 75850
rect -13520 75650 -13480 75850
rect -13410 75650 -13400 75850
rect -13600 75620 -13400 75650
rect -13100 75850 -12900 75880
rect -13100 75650 -13090 75850
rect -13020 75650 -12980 75850
rect -12910 75650 -12900 75850
rect -13100 75620 -12900 75650
rect -12600 75850 -12400 75880
rect -12600 75650 -12590 75850
rect -12520 75650 -12480 75850
rect -12410 75650 -12400 75850
rect -12600 75620 -12400 75650
rect -12100 75850 -12000 75880
rect -12100 75650 -12090 75850
rect -12020 75650 -12000 75850
rect -12100 75620 -12000 75650
rect -16000 75600 -15880 75620
rect -15620 75600 -15380 75620
rect -15120 75600 -14880 75620
rect -14620 75600 -14380 75620
rect -14120 75600 -13880 75620
rect -13620 75600 -13380 75620
rect -13120 75600 -12880 75620
rect -12620 75600 -12380 75620
rect -12120 75600 -12000 75620
rect -16000 75590 -12000 75600
rect -16000 75520 -15850 75590
rect -15650 75520 -15350 75590
rect -15150 75520 -14850 75590
rect -14650 75520 -14350 75590
rect -14150 75520 -13850 75590
rect -13650 75520 -13350 75590
rect -13150 75520 -12850 75590
rect -12650 75520 -12350 75590
rect -12150 75520 -12000 75590
rect -16000 75480 -12000 75520
rect -16000 75410 -15850 75480
rect -15650 75410 -15350 75480
rect -15150 75410 -14850 75480
rect -14650 75410 -14350 75480
rect -14150 75410 -13850 75480
rect -13650 75410 -13350 75480
rect -13150 75410 -12850 75480
rect -12650 75410 -12350 75480
rect -12150 75410 -12000 75480
rect -16000 75400 -12000 75410
rect -16000 75380 -15880 75400
rect -15620 75380 -15380 75400
rect -15120 75380 -14880 75400
rect -14620 75380 -14380 75400
rect -14120 75380 -13880 75400
rect -13620 75380 -13380 75400
rect -13120 75380 -12880 75400
rect -12620 75380 -12380 75400
rect -12120 75380 -12000 75400
rect -16000 75350 -15900 75380
rect -16000 75150 -15980 75350
rect -15910 75150 -15900 75350
rect -16000 75120 -15900 75150
rect -15600 75350 -15400 75380
rect -15600 75150 -15590 75350
rect -15520 75150 -15480 75350
rect -15410 75150 -15400 75350
rect -15600 75120 -15400 75150
rect -15100 75350 -14900 75380
rect -15100 75150 -15090 75350
rect -15020 75150 -14980 75350
rect -14910 75150 -14900 75350
rect -15100 75120 -14900 75150
rect -14600 75350 -14400 75380
rect -14600 75150 -14590 75350
rect -14520 75150 -14480 75350
rect -14410 75150 -14400 75350
rect -14600 75120 -14400 75150
rect -14100 75350 -13900 75380
rect -14100 75150 -14090 75350
rect -14020 75150 -13980 75350
rect -13910 75150 -13900 75350
rect -14100 75120 -13900 75150
rect -13600 75350 -13400 75380
rect -13600 75150 -13590 75350
rect -13520 75150 -13480 75350
rect -13410 75150 -13400 75350
rect -13600 75120 -13400 75150
rect -13100 75350 -12900 75380
rect -13100 75150 -13090 75350
rect -13020 75150 -12980 75350
rect -12910 75150 -12900 75350
rect -13100 75120 -12900 75150
rect -12600 75350 -12400 75380
rect -12600 75150 -12590 75350
rect -12520 75150 -12480 75350
rect -12410 75150 -12400 75350
rect -12600 75120 -12400 75150
rect -12100 75350 -12000 75380
rect -12100 75150 -12090 75350
rect -12020 75150 -12000 75350
rect -12100 75120 -12000 75150
rect -16000 75100 -15880 75120
rect -15620 75100 -15380 75120
rect -15120 75100 -14880 75120
rect -14620 75100 -14380 75120
rect -14120 75100 -13880 75120
rect -13620 75100 -13380 75120
rect -13120 75100 -12880 75120
rect -12620 75100 -12380 75120
rect -12120 75100 -12000 75120
rect -16000 75090 -12000 75100
rect -16000 75020 -15850 75090
rect -15650 75020 -15350 75090
rect -15150 75020 -14850 75090
rect -14650 75020 -14350 75090
rect -14150 75020 -13850 75090
rect -13650 75020 -13350 75090
rect -13150 75020 -12850 75090
rect -12650 75020 -12350 75090
rect -12150 75020 -12000 75090
rect -16000 74980 -12000 75020
rect -16000 74910 -15850 74980
rect -15650 74910 -15350 74980
rect -15150 74910 -14850 74980
rect -14650 74910 -14350 74980
rect -14150 74910 -13850 74980
rect -13650 74910 -13350 74980
rect -13150 74910 -12850 74980
rect -12650 74910 -12350 74980
rect -12150 74910 -12000 74980
rect -16000 74900 -12000 74910
rect -16000 74880 -15880 74900
rect -15620 74880 -15380 74900
rect -15120 74880 -14880 74900
rect -14620 74880 -14380 74900
rect -14120 74880 -13880 74900
rect -13620 74880 -13380 74900
rect -13120 74880 -12880 74900
rect -12620 74880 -12380 74900
rect -12120 74880 -12000 74900
rect -16000 74850 -15900 74880
rect -16000 74650 -15980 74850
rect -15910 74650 -15900 74850
rect -16000 74620 -15900 74650
rect -15600 74850 -15400 74880
rect -15600 74650 -15590 74850
rect -15520 74650 -15480 74850
rect -15410 74650 -15400 74850
rect -15600 74620 -15400 74650
rect -15100 74850 -14900 74880
rect -15100 74650 -15090 74850
rect -15020 74650 -14980 74850
rect -14910 74650 -14900 74850
rect -15100 74620 -14900 74650
rect -14600 74850 -14400 74880
rect -14600 74650 -14590 74850
rect -14520 74650 -14480 74850
rect -14410 74650 -14400 74850
rect -14600 74620 -14400 74650
rect -14100 74850 -13900 74880
rect -14100 74650 -14090 74850
rect -14020 74650 -13980 74850
rect -13910 74650 -13900 74850
rect -14100 74620 -13900 74650
rect -13600 74850 -13400 74880
rect -13600 74650 -13590 74850
rect -13520 74650 -13480 74850
rect -13410 74650 -13400 74850
rect -13600 74620 -13400 74650
rect -13100 74850 -12900 74880
rect -13100 74650 -13090 74850
rect -13020 74650 -12980 74850
rect -12910 74650 -12900 74850
rect -13100 74620 -12900 74650
rect -12600 74850 -12400 74880
rect -12600 74650 -12590 74850
rect -12520 74650 -12480 74850
rect -12410 74650 -12400 74850
rect -12600 74620 -12400 74650
rect -12100 74850 -12000 74880
rect -12100 74650 -12090 74850
rect -12020 74650 -12000 74850
rect -12100 74620 -12000 74650
rect -16000 74600 -15880 74620
rect -15620 74600 -15380 74620
rect -15120 74600 -14880 74620
rect -14620 74600 -14380 74620
rect -14120 74600 -13880 74620
rect -13620 74600 -13380 74620
rect -13120 74600 -12880 74620
rect -12620 74600 -12380 74620
rect -12120 74600 -12000 74620
rect -16000 74590 -12000 74600
rect -16000 74520 -15850 74590
rect -15650 74520 -15350 74590
rect -15150 74520 -14850 74590
rect -14650 74520 -14350 74590
rect -14150 74520 -13850 74590
rect -13650 74520 -13350 74590
rect -13150 74520 -12850 74590
rect -12650 74520 -12350 74590
rect -12150 74520 -12000 74590
rect -16000 74480 -12000 74520
rect -16000 74410 -15850 74480
rect -15650 74410 -15350 74480
rect -15150 74410 -14850 74480
rect -14650 74410 -14350 74480
rect -14150 74410 -13850 74480
rect -13650 74410 -13350 74480
rect -13150 74410 -12850 74480
rect -12650 74410 -12350 74480
rect -12150 74410 -12000 74480
rect -16000 74400 -12000 74410
rect -16000 74380 -15880 74400
rect -15620 74380 -15380 74400
rect -15120 74380 -14880 74400
rect -14620 74380 -14380 74400
rect -14120 74380 -13880 74400
rect -13620 74380 -13380 74400
rect -13120 74380 -12880 74400
rect -12620 74380 -12380 74400
rect -12120 74380 -12000 74400
rect -16000 74350 -15900 74380
rect -16000 74150 -15980 74350
rect -15910 74150 -15900 74350
rect -16000 74120 -15900 74150
rect -15600 74350 -15400 74380
rect -15600 74150 -15590 74350
rect -15520 74150 -15480 74350
rect -15410 74150 -15400 74350
rect -15600 74120 -15400 74150
rect -15100 74350 -14900 74380
rect -15100 74150 -15090 74350
rect -15020 74150 -14980 74350
rect -14910 74150 -14900 74350
rect -15100 74120 -14900 74150
rect -14600 74350 -14400 74380
rect -14600 74150 -14590 74350
rect -14520 74150 -14480 74350
rect -14410 74150 -14400 74350
rect -14600 74120 -14400 74150
rect -14100 74350 -13900 74380
rect -14100 74150 -14090 74350
rect -14020 74150 -13980 74350
rect -13910 74150 -13900 74350
rect -14100 74120 -13900 74150
rect -13600 74350 -13400 74380
rect -13600 74150 -13590 74350
rect -13520 74150 -13480 74350
rect -13410 74150 -13400 74350
rect -13600 74120 -13400 74150
rect -13100 74350 -12900 74380
rect -13100 74150 -13090 74350
rect -13020 74150 -12980 74350
rect -12910 74150 -12900 74350
rect -13100 74120 -12900 74150
rect -12600 74350 -12400 74380
rect -12600 74150 -12590 74350
rect -12520 74150 -12480 74350
rect -12410 74150 -12400 74350
rect -12600 74120 -12400 74150
rect -12100 74350 -12000 74380
rect -12100 74150 -12090 74350
rect -12020 74150 -12000 74350
rect -12100 74120 -12000 74150
rect -16000 74100 -15880 74120
rect -15620 74100 -15380 74120
rect -15120 74100 -14880 74120
rect -14620 74100 -14380 74120
rect -14120 74100 -13880 74120
rect -13620 74100 -13380 74120
rect -13120 74100 -12880 74120
rect -12620 74100 -12380 74120
rect -12120 74100 -12000 74120
rect -16000 74090 -12000 74100
rect -16000 74020 -15850 74090
rect -15650 74020 -15350 74090
rect -15150 74020 -14850 74090
rect -14650 74020 -14350 74090
rect -14150 74020 -13850 74090
rect -13650 74020 -13350 74090
rect -13150 74020 -12850 74090
rect -12650 74020 -12350 74090
rect -12150 74020 -12000 74090
rect -16000 73980 -12000 74020
rect -16000 73910 -15850 73980
rect -15650 73910 -15350 73980
rect -15150 73910 -14850 73980
rect -14650 73910 -14350 73980
rect -14150 73910 -13850 73980
rect -13650 73910 -13350 73980
rect -13150 73910 -12850 73980
rect -12650 73910 -12350 73980
rect -12150 73910 -12000 73980
rect -16000 73900 -12000 73910
rect -16000 73880 -15880 73900
rect -15620 73880 -15380 73900
rect -15120 73880 -14880 73900
rect -14620 73880 -14380 73900
rect -14120 73880 -13880 73900
rect -13620 73880 -13380 73900
rect -13120 73880 -12880 73900
rect -12620 73880 -12380 73900
rect -12120 73880 -12000 73900
rect -16000 73850 -15900 73880
rect -16000 73650 -15980 73850
rect -15910 73650 -15900 73850
rect -16000 73620 -15900 73650
rect -15600 73850 -15400 73880
rect -15600 73650 -15590 73850
rect -15520 73650 -15480 73850
rect -15410 73650 -15400 73850
rect -15600 73620 -15400 73650
rect -15100 73850 -14900 73880
rect -15100 73650 -15090 73850
rect -15020 73650 -14980 73850
rect -14910 73650 -14900 73850
rect -15100 73620 -14900 73650
rect -14600 73850 -14400 73880
rect -14600 73650 -14590 73850
rect -14520 73650 -14480 73850
rect -14410 73650 -14400 73850
rect -14600 73620 -14400 73650
rect -14100 73850 -13900 73880
rect -14100 73650 -14090 73850
rect -14020 73650 -13980 73850
rect -13910 73650 -13900 73850
rect -14100 73620 -13900 73650
rect -13600 73850 -13400 73880
rect -13600 73650 -13590 73850
rect -13520 73650 -13480 73850
rect -13410 73650 -13400 73850
rect -13600 73620 -13400 73650
rect -13100 73850 -12900 73880
rect -13100 73650 -13090 73850
rect -13020 73650 -12980 73850
rect -12910 73650 -12900 73850
rect -13100 73620 -12900 73650
rect -12600 73850 -12400 73880
rect -12600 73650 -12590 73850
rect -12520 73650 -12480 73850
rect -12410 73650 -12400 73850
rect -12600 73620 -12400 73650
rect -12100 73850 -12000 73880
rect -12100 73650 -12090 73850
rect -12020 73650 -12000 73850
rect -12100 73620 -12000 73650
rect -16000 73600 -15880 73620
rect -15620 73600 -15380 73620
rect -15120 73600 -14880 73620
rect -14620 73600 -14380 73620
rect -14120 73600 -13880 73620
rect -13620 73600 -13380 73620
rect -13120 73600 -12880 73620
rect -12620 73600 -12380 73620
rect -12120 73600 -12000 73620
rect -16000 73590 -12000 73600
rect -16000 73520 -15850 73590
rect -15650 73520 -15350 73590
rect -15150 73520 -14850 73590
rect -14650 73520 -14350 73590
rect -14150 73520 -13850 73590
rect -13650 73520 -13350 73590
rect -13150 73520 -12850 73590
rect -12650 73520 -12350 73590
rect -12150 73520 -12000 73590
rect -16000 73480 -12000 73520
rect -16000 73410 -15850 73480
rect -15650 73410 -15350 73480
rect -15150 73410 -14850 73480
rect -14650 73410 -14350 73480
rect -14150 73410 -13850 73480
rect -13650 73410 -13350 73480
rect -13150 73410 -12850 73480
rect -12650 73410 -12350 73480
rect -12150 73410 -12000 73480
rect -16000 73400 -12000 73410
rect -16000 73380 -15880 73400
rect -15620 73380 -15380 73400
rect -15120 73380 -14880 73400
rect -14620 73380 -14380 73400
rect -14120 73380 -13880 73400
rect -13620 73380 -13380 73400
rect -13120 73380 -12880 73400
rect -12620 73380 -12380 73400
rect -12120 73380 -12000 73400
rect -16000 73350 -15900 73380
rect -16000 73150 -15980 73350
rect -15910 73150 -15900 73350
rect -16000 73120 -15900 73150
rect -15600 73350 -15400 73380
rect -15600 73150 -15590 73350
rect -15520 73150 -15480 73350
rect -15410 73150 -15400 73350
rect -15600 73120 -15400 73150
rect -15100 73350 -14900 73380
rect -15100 73150 -15090 73350
rect -15020 73150 -14980 73350
rect -14910 73150 -14900 73350
rect -15100 73120 -14900 73150
rect -14600 73350 -14400 73380
rect -14600 73150 -14590 73350
rect -14520 73150 -14480 73350
rect -14410 73150 -14400 73350
rect -14600 73120 -14400 73150
rect -14100 73350 -13900 73380
rect -14100 73150 -14090 73350
rect -14020 73150 -13980 73350
rect -13910 73150 -13900 73350
rect -14100 73120 -13900 73150
rect -13600 73350 -13400 73380
rect -13600 73150 -13590 73350
rect -13520 73150 -13480 73350
rect -13410 73150 -13400 73350
rect -13600 73120 -13400 73150
rect -13100 73350 -12900 73380
rect -13100 73150 -13090 73350
rect -13020 73150 -12980 73350
rect -12910 73150 -12900 73350
rect -13100 73120 -12900 73150
rect -12600 73350 -12400 73380
rect -12600 73150 -12590 73350
rect -12520 73150 -12480 73350
rect -12410 73150 -12400 73350
rect -12600 73120 -12400 73150
rect -12100 73350 -12000 73380
rect -12100 73150 -12090 73350
rect -12020 73150 -12000 73350
rect -12100 73120 -12000 73150
rect -16000 73100 -15880 73120
rect -15620 73100 -15380 73120
rect -15120 73100 -14880 73120
rect -14620 73100 -14380 73120
rect -14120 73100 -13880 73120
rect -13620 73100 -13380 73120
rect -13120 73100 -12880 73120
rect -12620 73100 -12380 73120
rect -12120 73100 -12000 73120
rect -16000 73090 -12000 73100
rect -16000 73020 -15850 73090
rect -15650 73020 -15350 73090
rect -15150 73020 -14850 73090
rect -14650 73020 -14350 73090
rect -14150 73020 -13850 73090
rect -13650 73020 -13350 73090
rect -13150 73020 -12850 73090
rect -12650 73020 -12350 73090
rect -12150 73020 -12000 73090
rect -16000 72980 -12000 73020
rect -16000 72910 -15850 72980
rect -15650 72910 -15350 72980
rect -15150 72910 -14850 72980
rect -14650 72910 -14350 72980
rect -14150 72910 -13850 72980
rect -13650 72910 -13350 72980
rect -13150 72910 -12850 72980
rect -12650 72910 -12350 72980
rect -12150 72910 -12000 72980
rect -16000 72900 -12000 72910
rect -16000 72880 -15880 72900
rect -15620 72880 -15380 72900
rect -15120 72880 -14880 72900
rect -14620 72880 -14380 72900
rect -14120 72880 -13880 72900
rect -13620 72880 -13380 72900
rect -13120 72880 -12880 72900
rect -12620 72880 -12380 72900
rect -12120 72880 -12000 72900
rect -16000 72850 -15900 72880
rect -16000 72650 -15980 72850
rect -15910 72650 -15900 72850
rect -16000 72620 -15900 72650
rect -15600 72850 -15400 72880
rect -15600 72650 -15590 72850
rect -15520 72650 -15480 72850
rect -15410 72650 -15400 72850
rect -15600 72620 -15400 72650
rect -15100 72850 -14900 72880
rect -15100 72650 -15090 72850
rect -15020 72650 -14980 72850
rect -14910 72650 -14900 72850
rect -15100 72620 -14900 72650
rect -14600 72850 -14400 72880
rect -14600 72650 -14590 72850
rect -14520 72650 -14480 72850
rect -14410 72650 -14400 72850
rect -14600 72620 -14400 72650
rect -14100 72850 -13900 72880
rect -14100 72650 -14090 72850
rect -14020 72650 -13980 72850
rect -13910 72650 -13900 72850
rect -14100 72620 -13900 72650
rect -13600 72850 -13400 72880
rect -13600 72650 -13590 72850
rect -13520 72650 -13480 72850
rect -13410 72650 -13400 72850
rect -13600 72620 -13400 72650
rect -13100 72850 -12900 72880
rect -13100 72650 -13090 72850
rect -13020 72650 -12980 72850
rect -12910 72650 -12900 72850
rect -13100 72620 -12900 72650
rect -12600 72850 -12400 72880
rect -12600 72650 -12590 72850
rect -12520 72650 -12480 72850
rect -12410 72650 -12400 72850
rect -12600 72620 -12400 72650
rect -12100 72850 -12000 72880
rect -12100 72650 -12090 72850
rect -12020 72650 -12000 72850
rect -12100 72620 -12000 72650
rect -16000 72600 -15880 72620
rect -15620 72600 -15380 72620
rect -15120 72600 -14880 72620
rect -14620 72600 -14380 72620
rect -14120 72600 -13880 72620
rect -13620 72600 -13380 72620
rect -13120 72600 -12880 72620
rect -12620 72600 -12380 72620
rect -12120 72600 -12000 72620
rect -16000 72590 -12000 72600
rect -16000 72520 -15850 72590
rect -15650 72520 -15350 72590
rect -15150 72520 -14850 72590
rect -14650 72520 -14350 72590
rect -14150 72520 -13850 72590
rect -13650 72520 -13350 72590
rect -13150 72520 -12850 72590
rect -12650 72520 -12350 72590
rect -12150 72520 -12000 72590
rect -16000 72480 -12000 72520
rect -16000 72410 -15850 72480
rect -15650 72410 -15350 72480
rect -15150 72410 -14850 72480
rect -14650 72410 -14350 72480
rect -14150 72410 -13850 72480
rect -13650 72410 -13350 72480
rect -13150 72410 -12850 72480
rect -12650 72410 -12350 72480
rect -12150 72410 -12000 72480
rect -16000 72400 -12000 72410
rect -16000 72380 -15880 72400
rect -15620 72380 -15380 72400
rect -15120 72380 -14880 72400
rect -14620 72380 -14380 72400
rect -14120 72380 -13880 72400
rect -13620 72380 -13380 72400
rect -13120 72380 -12880 72400
rect -12620 72380 -12380 72400
rect -12120 72380 -12000 72400
rect -16000 72350 -15900 72380
rect -16000 72150 -15980 72350
rect -15910 72150 -15900 72350
rect -16000 72120 -15900 72150
rect -15600 72350 -15400 72380
rect -15600 72150 -15590 72350
rect -15520 72150 -15480 72350
rect -15410 72150 -15400 72350
rect -15600 72120 -15400 72150
rect -15100 72350 -14900 72380
rect -15100 72150 -15090 72350
rect -15020 72150 -14980 72350
rect -14910 72150 -14900 72350
rect -15100 72120 -14900 72150
rect -14600 72350 -14400 72380
rect -14600 72150 -14590 72350
rect -14520 72150 -14480 72350
rect -14410 72150 -14400 72350
rect -14600 72120 -14400 72150
rect -14100 72350 -13900 72380
rect -14100 72150 -14090 72350
rect -14020 72150 -13980 72350
rect -13910 72150 -13900 72350
rect -14100 72120 -13900 72150
rect -13600 72350 -13400 72380
rect -13600 72150 -13590 72350
rect -13520 72150 -13480 72350
rect -13410 72150 -13400 72350
rect -13600 72120 -13400 72150
rect -13100 72350 -12900 72380
rect -13100 72150 -13090 72350
rect -13020 72150 -12980 72350
rect -12910 72150 -12900 72350
rect -13100 72120 -12900 72150
rect -12600 72350 -12400 72380
rect -12600 72150 -12590 72350
rect -12520 72150 -12480 72350
rect -12410 72150 -12400 72350
rect -12600 72120 -12400 72150
rect -12100 72350 -12000 72380
rect -12100 72150 -12090 72350
rect -12020 72150 -12000 72350
rect -12100 72120 -12000 72150
rect -16000 72100 -15880 72120
rect -15620 72100 -15380 72120
rect -15120 72100 -14880 72120
rect -14620 72100 -14380 72120
rect -14120 72100 -13880 72120
rect -13620 72100 -13380 72120
rect -13120 72100 -12880 72120
rect -12620 72100 -12380 72120
rect -12120 72100 -12000 72120
rect -16000 72090 -12000 72100
rect -16000 72020 -15850 72090
rect -15650 72020 -15350 72090
rect -15150 72020 -14850 72090
rect -14650 72020 -14350 72090
rect -14150 72020 -13850 72090
rect -13650 72020 -13350 72090
rect -13150 72020 -12850 72090
rect -12650 72020 -12350 72090
rect -12150 72020 -12000 72090
rect -16000 71980 -12000 72020
rect -16000 71910 -15850 71980
rect -15650 71910 -15350 71980
rect -15150 71910 -14850 71980
rect -14650 71910 -14350 71980
rect -14150 71910 -13850 71980
rect -13650 71910 -13350 71980
rect -13150 71910 -12850 71980
rect -12650 71910 -12350 71980
rect -12150 71910 -12000 71980
rect -16000 71900 -12000 71910
rect -16000 71880 -15880 71900
rect -15620 71880 -15380 71900
rect -15120 71880 -14880 71900
rect -14620 71880 -14380 71900
rect -14120 71880 -13880 71900
rect -13620 71880 -13380 71900
rect -13120 71880 -12880 71900
rect -12620 71880 -12380 71900
rect -12120 71880 -12000 71900
rect -16000 71850 -15900 71880
rect -16000 71650 -15980 71850
rect -15910 71650 -15900 71850
rect -16000 71620 -15900 71650
rect -15600 71850 -15400 71880
rect -15600 71650 -15590 71850
rect -15520 71650 -15480 71850
rect -15410 71650 -15400 71850
rect -15600 71620 -15400 71650
rect -15100 71850 -14900 71880
rect -15100 71650 -15090 71850
rect -15020 71650 -14980 71850
rect -14910 71650 -14900 71850
rect -15100 71620 -14900 71650
rect -14600 71850 -14400 71880
rect -14600 71650 -14590 71850
rect -14520 71650 -14480 71850
rect -14410 71650 -14400 71850
rect -14600 71620 -14400 71650
rect -14100 71850 -13900 71880
rect -14100 71650 -14090 71850
rect -14020 71650 -13980 71850
rect -13910 71650 -13900 71850
rect -14100 71620 -13900 71650
rect -13600 71850 -13400 71880
rect -13600 71650 -13590 71850
rect -13520 71650 -13480 71850
rect -13410 71650 -13400 71850
rect -13600 71620 -13400 71650
rect -13100 71850 -12900 71880
rect -13100 71650 -13090 71850
rect -13020 71650 -12980 71850
rect -12910 71650 -12900 71850
rect -13100 71620 -12900 71650
rect -12600 71850 -12400 71880
rect -12600 71650 -12590 71850
rect -12520 71650 -12480 71850
rect -12410 71650 -12400 71850
rect -12600 71620 -12400 71650
rect -12100 71850 -12000 71880
rect -12100 71650 -12090 71850
rect -12020 71650 -12000 71850
rect -12100 71620 -12000 71650
rect -16000 71600 -15880 71620
rect -15620 71600 -15380 71620
rect -15120 71600 -14880 71620
rect -14620 71600 -14380 71620
rect -14120 71600 -13880 71620
rect -13620 71600 -13380 71620
rect -13120 71600 -12880 71620
rect -12620 71600 -12380 71620
rect -12120 71600 -12000 71620
rect -16000 71590 -12000 71600
rect -16000 71520 -15850 71590
rect -15650 71520 -15350 71590
rect -15150 71520 -14850 71590
rect -14650 71520 -14350 71590
rect -14150 71520 -13850 71590
rect -13650 71520 -13350 71590
rect -13150 71520 -12850 71590
rect -12650 71520 -12350 71590
rect -12150 71520 -12000 71590
rect -16000 71480 -12000 71520
rect -16000 71410 -15850 71480
rect -15650 71410 -15350 71480
rect -15150 71410 -14850 71480
rect -14650 71410 -14350 71480
rect -14150 71410 -13850 71480
rect -13650 71410 -13350 71480
rect -13150 71410 -12850 71480
rect -12650 71410 -12350 71480
rect -12150 71410 -12000 71480
rect -16000 71400 -12000 71410
rect -16000 71380 -15880 71400
rect -15620 71380 -15380 71400
rect -15120 71380 -14880 71400
rect -14620 71380 -14380 71400
rect -14120 71380 -13880 71400
rect -13620 71380 -13380 71400
rect -13120 71380 -12880 71400
rect -12620 71380 -12380 71400
rect -12120 71380 -12000 71400
rect -16000 71350 -15900 71380
rect -16000 71150 -15980 71350
rect -15910 71150 -15900 71350
rect -16000 71120 -15900 71150
rect -15600 71350 -15400 71380
rect -15600 71150 -15590 71350
rect -15520 71150 -15480 71350
rect -15410 71150 -15400 71350
rect -15600 71120 -15400 71150
rect -15100 71350 -14900 71380
rect -15100 71150 -15090 71350
rect -15020 71150 -14980 71350
rect -14910 71150 -14900 71350
rect -15100 71120 -14900 71150
rect -14600 71350 -14400 71380
rect -14600 71150 -14590 71350
rect -14520 71150 -14480 71350
rect -14410 71150 -14400 71350
rect -14600 71120 -14400 71150
rect -14100 71350 -13900 71380
rect -14100 71150 -14090 71350
rect -14020 71150 -13980 71350
rect -13910 71150 -13900 71350
rect -14100 71120 -13900 71150
rect -13600 71350 -13400 71380
rect -13600 71150 -13590 71350
rect -13520 71150 -13480 71350
rect -13410 71150 -13400 71350
rect -13600 71120 -13400 71150
rect -13100 71350 -12900 71380
rect -13100 71150 -13090 71350
rect -13020 71150 -12980 71350
rect -12910 71150 -12900 71350
rect -13100 71120 -12900 71150
rect -12600 71350 -12400 71380
rect -12600 71150 -12590 71350
rect -12520 71150 -12480 71350
rect -12410 71150 -12400 71350
rect -12600 71120 -12400 71150
rect -12100 71350 -12000 71380
rect -12100 71150 -12090 71350
rect -12020 71150 -12000 71350
rect -12100 71120 -12000 71150
rect -16000 71100 -15880 71120
rect -15620 71100 -15380 71120
rect -15120 71100 -14880 71120
rect -14620 71100 -14380 71120
rect -14120 71100 -13880 71120
rect -13620 71100 -13380 71120
rect -13120 71100 -12880 71120
rect -12620 71100 -12380 71120
rect -12120 71100 -12000 71120
rect -16000 71090 -12000 71100
rect -16000 71020 -15850 71090
rect -15650 71020 -15350 71090
rect -15150 71020 -14850 71090
rect -14650 71020 -14350 71090
rect -14150 71020 -13850 71090
rect -13650 71020 -13350 71090
rect -13150 71020 -12850 71090
rect -12650 71020 -12350 71090
rect -12150 71020 -12000 71090
rect -16000 70980 -12000 71020
rect -16000 70910 -15850 70980
rect -15650 70910 -15350 70980
rect -15150 70910 -14850 70980
rect -14650 70910 -14350 70980
rect -14150 70910 -13850 70980
rect -13650 70910 -13350 70980
rect -13150 70910 -12850 70980
rect -12650 70910 -12350 70980
rect -12150 70910 -12000 70980
rect -16000 70900 -12000 70910
rect -16000 70880 -15880 70900
rect -15620 70880 -15380 70900
rect -15120 70880 -14880 70900
rect -14620 70880 -14380 70900
rect -14120 70880 -13880 70900
rect -13620 70880 -13380 70900
rect -13120 70880 -12880 70900
rect -12620 70880 -12380 70900
rect -12120 70880 -12000 70900
rect -16000 70850 -15900 70880
rect -16000 70650 -15980 70850
rect -15910 70650 -15900 70850
rect -16000 70620 -15900 70650
rect -15600 70850 -15400 70880
rect -15600 70650 -15590 70850
rect -15520 70650 -15480 70850
rect -15410 70650 -15400 70850
rect -15600 70620 -15400 70650
rect -15100 70850 -14900 70880
rect -15100 70650 -15090 70850
rect -15020 70650 -14980 70850
rect -14910 70650 -14900 70850
rect -15100 70620 -14900 70650
rect -14600 70850 -14400 70880
rect -14600 70650 -14590 70850
rect -14520 70650 -14480 70850
rect -14410 70650 -14400 70850
rect -14600 70620 -14400 70650
rect -14100 70850 -13900 70880
rect -14100 70650 -14090 70850
rect -14020 70650 -13980 70850
rect -13910 70650 -13900 70850
rect -14100 70620 -13900 70650
rect -13600 70850 -13400 70880
rect -13600 70650 -13590 70850
rect -13520 70650 -13480 70850
rect -13410 70650 -13400 70850
rect -13600 70620 -13400 70650
rect -13100 70850 -12900 70880
rect -13100 70650 -13090 70850
rect -13020 70650 -12980 70850
rect -12910 70650 -12900 70850
rect -13100 70620 -12900 70650
rect -12600 70850 -12400 70880
rect -12600 70650 -12590 70850
rect -12520 70650 -12480 70850
rect -12410 70650 -12400 70850
rect -12600 70620 -12400 70650
rect -12100 70850 -12000 70880
rect -12100 70650 -12090 70850
rect -12020 70650 -12000 70850
rect -12100 70620 -12000 70650
rect -16000 70600 -15880 70620
rect -15620 70600 -15380 70620
rect -15120 70600 -14880 70620
rect -14620 70600 -14380 70620
rect -14120 70600 -13880 70620
rect -13620 70600 -13380 70620
rect -13120 70600 -12880 70620
rect -12620 70600 -12380 70620
rect -12120 70600 -12000 70620
rect -16000 70590 -12000 70600
rect -16000 70520 -15850 70590
rect -15650 70520 -15350 70590
rect -15150 70520 -14850 70590
rect -14650 70520 -14350 70590
rect -14150 70520 -13850 70590
rect -13650 70520 -13350 70590
rect -13150 70520 -12850 70590
rect -12650 70520 -12350 70590
rect -12150 70520 -12000 70590
rect -16000 70480 -12000 70520
rect -16000 70410 -15850 70480
rect -15650 70410 -15350 70480
rect -15150 70410 -14850 70480
rect -14650 70410 -14350 70480
rect -14150 70410 -13850 70480
rect -13650 70410 -13350 70480
rect -13150 70410 -12850 70480
rect -12650 70410 -12350 70480
rect -12150 70410 -12000 70480
rect -16000 70400 -12000 70410
rect -16000 70380 -15880 70400
rect -15620 70380 -15380 70400
rect -15120 70380 -14880 70400
rect -14620 70380 -14380 70400
rect -14120 70380 -13880 70400
rect -13620 70380 -13380 70400
rect -13120 70380 -12880 70400
rect -12620 70380 -12380 70400
rect -12120 70380 -12000 70400
rect -16000 70350 -15900 70380
rect -16000 70150 -15980 70350
rect -15910 70150 -15900 70350
rect -16000 70120 -15900 70150
rect -15600 70350 -15400 70380
rect -15600 70150 -15590 70350
rect -15520 70150 -15480 70350
rect -15410 70150 -15400 70350
rect -15600 70120 -15400 70150
rect -15100 70350 -14900 70380
rect -15100 70150 -15090 70350
rect -15020 70150 -14980 70350
rect -14910 70150 -14900 70350
rect -15100 70120 -14900 70150
rect -14600 70350 -14400 70380
rect -14600 70150 -14590 70350
rect -14520 70150 -14480 70350
rect -14410 70150 -14400 70350
rect -14600 70120 -14400 70150
rect -14100 70350 -13900 70380
rect -14100 70150 -14090 70350
rect -14020 70150 -13980 70350
rect -13910 70150 -13900 70350
rect -14100 70120 -13900 70150
rect -13600 70350 -13400 70380
rect -13600 70150 -13590 70350
rect -13520 70150 -13480 70350
rect -13410 70150 -13400 70350
rect -13600 70120 -13400 70150
rect -13100 70350 -12900 70380
rect -13100 70150 -13090 70350
rect -13020 70150 -12980 70350
rect -12910 70150 -12900 70350
rect -13100 70120 -12900 70150
rect -12600 70350 -12400 70380
rect -12600 70150 -12590 70350
rect -12520 70150 -12480 70350
rect -12410 70150 -12400 70350
rect -12600 70120 -12400 70150
rect -12100 70350 -12000 70380
rect -12100 70150 -12090 70350
rect -12020 70150 -12000 70350
rect -12100 70120 -12000 70150
rect -16000 70100 -15880 70120
rect -15620 70100 -15380 70120
rect -15120 70100 -14880 70120
rect -14620 70100 -14380 70120
rect -14120 70100 -13880 70120
rect -13620 70100 -13380 70120
rect -13120 70100 -12880 70120
rect -12620 70100 -12380 70120
rect -12120 70100 -12000 70120
rect -16000 70090 -12000 70100
rect -16000 70020 -15850 70090
rect -15650 70020 -15350 70090
rect -15150 70020 -14850 70090
rect -14650 70020 -14350 70090
rect -14150 70020 -13850 70090
rect -13650 70020 -13350 70090
rect -13150 70020 -12850 70090
rect -12650 70020 -12350 70090
rect -12150 70020 -12000 70090
rect -16000 69980 -12000 70020
rect -16000 69910 -15850 69980
rect -15650 69910 -15350 69980
rect -15150 69910 -14850 69980
rect -14650 69910 -14350 69980
rect -14150 69910 -13850 69980
rect -13650 69910 -13350 69980
rect -13150 69910 -12850 69980
rect -12650 69910 -12350 69980
rect -12150 69910 -12000 69980
rect -16000 69900 -12000 69910
rect -16000 69880 -15880 69900
rect -15620 69880 -15380 69900
rect -15120 69880 -14880 69900
rect -14620 69880 -14380 69900
rect -14120 69880 -13880 69900
rect -13620 69880 -13380 69900
rect -13120 69880 -12880 69900
rect -12620 69880 -12380 69900
rect -12120 69880 -12000 69900
rect -16000 69850 -15900 69880
rect -16000 69650 -15980 69850
rect -15910 69650 -15900 69850
rect -16000 69620 -15900 69650
rect -15600 69850 -15400 69880
rect -15600 69650 -15590 69850
rect -15520 69650 -15480 69850
rect -15410 69650 -15400 69850
rect -15600 69620 -15400 69650
rect -15100 69850 -14900 69880
rect -15100 69650 -15090 69850
rect -15020 69650 -14980 69850
rect -14910 69650 -14900 69850
rect -15100 69620 -14900 69650
rect -14600 69850 -14400 69880
rect -14600 69650 -14590 69850
rect -14520 69650 -14480 69850
rect -14410 69650 -14400 69850
rect -14600 69620 -14400 69650
rect -14100 69850 -13900 69880
rect -14100 69650 -14090 69850
rect -14020 69650 -13980 69850
rect -13910 69650 -13900 69850
rect -14100 69620 -13900 69650
rect -13600 69850 -13400 69880
rect -13600 69650 -13590 69850
rect -13520 69650 -13480 69850
rect -13410 69650 -13400 69850
rect -13600 69620 -13400 69650
rect -13100 69850 -12900 69880
rect -13100 69650 -13090 69850
rect -13020 69650 -12980 69850
rect -12910 69650 -12900 69850
rect -13100 69620 -12900 69650
rect -12600 69850 -12400 69880
rect -12600 69650 -12590 69850
rect -12520 69650 -12480 69850
rect -12410 69650 -12400 69850
rect -12600 69620 -12400 69650
rect -12100 69850 -12000 69880
rect -12100 69650 -12090 69850
rect -12020 69650 -12000 69850
rect -12100 69620 -12000 69650
rect -16000 69600 -15880 69620
rect -15620 69600 -15380 69620
rect -15120 69600 -14880 69620
rect -14620 69600 -14380 69620
rect -14120 69600 -13880 69620
rect -13620 69600 -13380 69620
rect -13120 69600 -12880 69620
rect -12620 69600 -12380 69620
rect -12120 69600 -12000 69620
rect -16000 69590 -12000 69600
rect -16000 69520 -15850 69590
rect -15650 69520 -15350 69590
rect -15150 69520 -14850 69590
rect -14650 69520 -14350 69590
rect -14150 69520 -13850 69590
rect -13650 69520 -13350 69590
rect -13150 69520 -12850 69590
rect -12650 69520 -12350 69590
rect -12150 69520 -12000 69590
rect -16000 69480 -12000 69520
rect -16000 69410 -15850 69480
rect -15650 69410 -15350 69480
rect -15150 69410 -14850 69480
rect -14650 69410 -14350 69480
rect -14150 69410 -13850 69480
rect -13650 69410 -13350 69480
rect -13150 69410 -12850 69480
rect -12650 69410 -12350 69480
rect -12150 69410 -12000 69480
rect -16000 69400 -12000 69410
rect -16000 69380 -15880 69400
rect -15620 69380 -15380 69400
rect -15120 69380 -14880 69400
rect -14620 69380 -14380 69400
rect -14120 69380 -13880 69400
rect -13620 69380 -13380 69400
rect -13120 69380 -12880 69400
rect -12620 69380 -12380 69400
rect -12120 69380 -12000 69400
rect -16000 69350 -15900 69380
rect -16000 69150 -15980 69350
rect -15910 69150 -15900 69350
rect -16000 69120 -15900 69150
rect -15600 69350 -15400 69380
rect -15600 69150 -15590 69350
rect -15520 69150 -15480 69350
rect -15410 69150 -15400 69350
rect -15600 69120 -15400 69150
rect -15100 69350 -14900 69380
rect -15100 69150 -15090 69350
rect -15020 69150 -14980 69350
rect -14910 69150 -14900 69350
rect -15100 69120 -14900 69150
rect -14600 69350 -14400 69380
rect -14600 69150 -14590 69350
rect -14520 69150 -14480 69350
rect -14410 69150 -14400 69350
rect -14600 69120 -14400 69150
rect -14100 69350 -13900 69380
rect -14100 69150 -14090 69350
rect -14020 69150 -13980 69350
rect -13910 69150 -13900 69350
rect -14100 69120 -13900 69150
rect -13600 69350 -13400 69380
rect -13600 69150 -13590 69350
rect -13520 69150 -13480 69350
rect -13410 69150 -13400 69350
rect -13600 69120 -13400 69150
rect -13100 69350 -12900 69380
rect -13100 69150 -13090 69350
rect -13020 69150 -12980 69350
rect -12910 69150 -12900 69350
rect -13100 69120 -12900 69150
rect -12600 69350 -12400 69380
rect -12600 69150 -12590 69350
rect -12520 69150 -12480 69350
rect -12410 69150 -12400 69350
rect -12600 69120 -12400 69150
rect -12100 69350 -12000 69380
rect -12100 69150 -12090 69350
rect -12020 69150 -12000 69350
rect -12100 69120 -12000 69150
rect -16000 69100 -15880 69120
rect -15620 69100 -15380 69120
rect -15120 69100 -14880 69120
rect -14620 69100 -14380 69120
rect -14120 69100 -13880 69120
rect -13620 69100 -13380 69120
rect -13120 69100 -12880 69120
rect -12620 69100 -12380 69120
rect -12120 69100 -12000 69120
rect -16000 69090 -12000 69100
rect -16000 69020 -15850 69090
rect -15650 69020 -15350 69090
rect -15150 69020 -14850 69090
rect -14650 69020 -14350 69090
rect -14150 69020 -13850 69090
rect -13650 69020 -13350 69090
rect -13150 69020 -12850 69090
rect -12650 69020 -12350 69090
rect -12150 69020 -12000 69090
rect -16000 68980 -12000 69020
rect -16000 68910 -15850 68980
rect -15650 68910 -15350 68980
rect -15150 68910 -14850 68980
rect -14650 68910 -14350 68980
rect -14150 68910 -13850 68980
rect -13650 68910 -13350 68980
rect -13150 68910 -12850 68980
rect -12650 68910 -12350 68980
rect -12150 68910 -12000 68980
rect -16000 68900 -12000 68910
rect -16000 68880 -15880 68900
rect -15620 68880 -15380 68900
rect -15120 68880 -14880 68900
rect -14620 68880 -14380 68900
rect -14120 68880 -13880 68900
rect -13620 68880 -13380 68900
rect -13120 68880 -12880 68900
rect -12620 68880 -12380 68900
rect -12120 68880 -12000 68900
rect -16000 68850 -15900 68880
rect -16000 68650 -15980 68850
rect -15910 68650 -15900 68850
rect -16000 68620 -15900 68650
rect -15600 68850 -15400 68880
rect -15600 68650 -15590 68850
rect -15520 68650 -15480 68850
rect -15410 68650 -15400 68850
rect -15600 68620 -15400 68650
rect -15100 68850 -14900 68880
rect -15100 68650 -15090 68850
rect -15020 68650 -14980 68850
rect -14910 68650 -14900 68850
rect -15100 68620 -14900 68650
rect -14600 68850 -14400 68880
rect -14600 68650 -14590 68850
rect -14520 68650 -14480 68850
rect -14410 68650 -14400 68850
rect -14600 68620 -14400 68650
rect -14100 68850 -13900 68880
rect -14100 68650 -14090 68850
rect -14020 68650 -13980 68850
rect -13910 68650 -13900 68850
rect -14100 68620 -13900 68650
rect -13600 68850 -13400 68880
rect -13600 68650 -13590 68850
rect -13520 68650 -13480 68850
rect -13410 68650 -13400 68850
rect -13600 68620 -13400 68650
rect -13100 68850 -12900 68880
rect -13100 68650 -13090 68850
rect -13020 68650 -12980 68850
rect -12910 68650 -12900 68850
rect -13100 68620 -12900 68650
rect -12600 68850 -12400 68880
rect -12600 68650 -12590 68850
rect -12520 68650 -12480 68850
rect -12410 68650 -12400 68850
rect -12600 68620 -12400 68650
rect -12100 68850 -12000 68880
rect -12100 68650 -12090 68850
rect -12020 68650 -12000 68850
rect -12100 68620 -12000 68650
rect -16000 68600 -15880 68620
rect -15620 68600 -15380 68620
rect -15120 68600 -14880 68620
rect -14620 68600 -14380 68620
rect -14120 68600 -13880 68620
rect -13620 68600 -13380 68620
rect -13120 68600 -12880 68620
rect -12620 68600 -12380 68620
rect -12120 68600 -12000 68620
rect -16000 68590 -12000 68600
rect -16000 68520 -15850 68590
rect -15650 68520 -15350 68590
rect -15150 68520 -14850 68590
rect -14650 68520 -14350 68590
rect -14150 68520 -13850 68590
rect -13650 68520 -13350 68590
rect -13150 68520 -12850 68590
rect -12650 68520 -12350 68590
rect -12150 68520 -12000 68590
rect -16000 68480 -12000 68520
rect -16000 68410 -15850 68480
rect -15650 68410 -15350 68480
rect -15150 68410 -14850 68480
rect -14650 68410 -14350 68480
rect -14150 68410 -13850 68480
rect -13650 68410 -13350 68480
rect -13150 68410 -12850 68480
rect -12650 68410 -12350 68480
rect -12150 68410 -12000 68480
rect -16000 68400 -12000 68410
rect -16000 68380 -15880 68400
rect -15620 68380 -15380 68400
rect -15120 68380 -14880 68400
rect -14620 68380 -14380 68400
rect -14120 68380 -13880 68400
rect -13620 68380 -13380 68400
rect -13120 68380 -12880 68400
rect -12620 68380 -12380 68400
rect -12120 68380 -12000 68400
rect -16000 68350 -15900 68380
rect -16000 68150 -15980 68350
rect -15910 68150 -15900 68350
rect -16000 68120 -15900 68150
rect -15600 68350 -15400 68380
rect -15600 68150 -15590 68350
rect -15520 68150 -15480 68350
rect -15410 68150 -15400 68350
rect -15600 68120 -15400 68150
rect -15100 68350 -14900 68380
rect -15100 68150 -15090 68350
rect -15020 68150 -14980 68350
rect -14910 68150 -14900 68350
rect -15100 68120 -14900 68150
rect -14600 68350 -14400 68380
rect -14600 68150 -14590 68350
rect -14520 68150 -14480 68350
rect -14410 68150 -14400 68350
rect -14600 68120 -14400 68150
rect -14100 68350 -13900 68380
rect -14100 68150 -14090 68350
rect -14020 68150 -13980 68350
rect -13910 68150 -13900 68350
rect -14100 68120 -13900 68150
rect -13600 68350 -13400 68380
rect -13600 68150 -13590 68350
rect -13520 68150 -13480 68350
rect -13410 68150 -13400 68350
rect -13600 68120 -13400 68150
rect -13100 68350 -12900 68380
rect -13100 68150 -13090 68350
rect -13020 68150 -12980 68350
rect -12910 68150 -12900 68350
rect -13100 68120 -12900 68150
rect -12600 68350 -12400 68380
rect -12600 68150 -12590 68350
rect -12520 68150 -12480 68350
rect -12410 68150 -12400 68350
rect -12600 68120 -12400 68150
rect -12100 68350 -12000 68380
rect -12100 68150 -12090 68350
rect -12020 68150 -12000 68350
rect -12100 68120 -12000 68150
rect -16000 68100 -15880 68120
rect -15620 68100 -15380 68120
rect -15120 68100 -14880 68120
rect -14620 68100 -14380 68120
rect -14120 68100 -13880 68120
rect -13620 68100 -13380 68120
rect -13120 68100 -12880 68120
rect -12620 68100 -12380 68120
rect -12120 68100 -12000 68120
rect -16000 68090 -12000 68100
rect -16000 68020 -15850 68090
rect -15650 68020 -15350 68090
rect -15150 68020 -14850 68090
rect -14650 68020 -14350 68090
rect -14150 68020 -13850 68090
rect -13650 68020 -13350 68090
rect -13150 68020 -12850 68090
rect -12650 68020 -12350 68090
rect -12150 68020 -12000 68090
rect -16000 67980 -12000 68020
rect -16000 67910 -15850 67980
rect -15650 67910 -15350 67980
rect -15150 67910 -14850 67980
rect -14650 67910 -14350 67980
rect -14150 67910 -13850 67980
rect -13650 67910 -13350 67980
rect -13150 67910 -12850 67980
rect -12650 67910 -12350 67980
rect -12150 67910 -12000 67980
rect -16000 67900 -12000 67910
rect -16000 67880 -15880 67900
rect -15620 67880 -15380 67900
rect -15120 67880 -14880 67900
rect -14620 67880 -14380 67900
rect -14120 67880 -13880 67900
rect -13620 67880 -13380 67900
rect -13120 67880 -12880 67900
rect -12620 67880 -12380 67900
rect -12120 67880 -12000 67900
rect -16000 67850 -15900 67880
rect -16000 67650 -15980 67850
rect -15910 67650 -15900 67850
rect -16000 67620 -15900 67650
rect -15600 67850 -15400 67880
rect -15600 67650 -15590 67850
rect -15520 67650 -15480 67850
rect -15410 67650 -15400 67850
rect -15600 67620 -15400 67650
rect -15100 67850 -14900 67880
rect -15100 67650 -15090 67850
rect -15020 67650 -14980 67850
rect -14910 67650 -14900 67850
rect -15100 67620 -14900 67650
rect -14600 67850 -14400 67880
rect -14600 67650 -14590 67850
rect -14520 67650 -14480 67850
rect -14410 67650 -14400 67850
rect -14600 67620 -14400 67650
rect -14100 67850 -13900 67880
rect -14100 67650 -14090 67850
rect -14020 67650 -13980 67850
rect -13910 67650 -13900 67850
rect -14100 67620 -13900 67650
rect -13600 67850 -13400 67880
rect -13600 67650 -13590 67850
rect -13520 67650 -13480 67850
rect -13410 67650 -13400 67850
rect -13600 67620 -13400 67650
rect -13100 67850 -12900 67880
rect -13100 67650 -13090 67850
rect -13020 67650 -12980 67850
rect -12910 67650 -12900 67850
rect -13100 67620 -12900 67650
rect -12600 67850 -12400 67880
rect -12600 67650 -12590 67850
rect -12520 67650 -12480 67850
rect -12410 67650 -12400 67850
rect -12600 67620 -12400 67650
rect -12100 67850 -12000 67880
rect -12100 67650 -12090 67850
rect -12020 67650 -12000 67850
rect -12100 67620 -12000 67650
rect -16000 67600 -15880 67620
rect -15620 67600 -15380 67620
rect -15120 67600 -14880 67620
rect -14620 67600 -14380 67620
rect -14120 67600 -13880 67620
rect -13620 67600 -13380 67620
rect -13120 67600 -12880 67620
rect -12620 67600 -12380 67620
rect -12120 67600 -12000 67620
rect -16000 67590 -12000 67600
rect -16000 67520 -15850 67590
rect -15650 67520 -15350 67590
rect -15150 67520 -14850 67590
rect -14650 67520 -14350 67590
rect -14150 67520 -13850 67590
rect -13650 67520 -13350 67590
rect -13150 67520 -12850 67590
rect -12650 67520 -12350 67590
rect -12150 67520 -12000 67590
rect -16000 67480 -12000 67520
rect -16000 67410 -15850 67480
rect -15650 67410 -15350 67480
rect -15150 67410 -14850 67480
rect -14650 67410 -14350 67480
rect -14150 67410 -13850 67480
rect -13650 67410 -13350 67480
rect -13150 67410 -12850 67480
rect -12650 67410 -12350 67480
rect -12150 67410 -12000 67480
rect -16000 67400 -12000 67410
rect -16000 67380 -15880 67400
rect -15620 67380 -15380 67400
rect -15120 67380 -14880 67400
rect -14620 67380 -14380 67400
rect -14120 67380 -13880 67400
rect -13620 67380 -13380 67400
rect -13120 67380 -12880 67400
rect -12620 67380 -12380 67400
rect -12120 67380 -12000 67400
rect -16000 67350 -15900 67380
rect -16000 67150 -15980 67350
rect -15910 67150 -15900 67350
rect -16000 67120 -15900 67150
rect -15600 67350 -15400 67380
rect -15600 67150 -15590 67350
rect -15520 67150 -15480 67350
rect -15410 67150 -15400 67350
rect -15600 67120 -15400 67150
rect -15100 67350 -14900 67380
rect -15100 67150 -15090 67350
rect -15020 67150 -14980 67350
rect -14910 67150 -14900 67350
rect -15100 67120 -14900 67150
rect -14600 67350 -14400 67380
rect -14600 67150 -14590 67350
rect -14520 67150 -14480 67350
rect -14410 67150 -14400 67350
rect -14600 67120 -14400 67150
rect -14100 67350 -13900 67380
rect -14100 67150 -14090 67350
rect -14020 67150 -13980 67350
rect -13910 67150 -13900 67350
rect -14100 67120 -13900 67150
rect -13600 67350 -13400 67380
rect -13600 67150 -13590 67350
rect -13520 67150 -13480 67350
rect -13410 67150 -13400 67350
rect -13600 67120 -13400 67150
rect -13100 67350 -12900 67380
rect -13100 67150 -13090 67350
rect -13020 67150 -12980 67350
rect -12910 67150 -12900 67350
rect -13100 67120 -12900 67150
rect -12600 67350 -12400 67380
rect -12600 67150 -12590 67350
rect -12520 67150 -12480 67350
rect -12410 67150 -12400 67350
rect -12600 67120 -12400 67150
rect -12100 67350 -12000 67380
rect -12100 67150 -12090 67350
rect -12020 67150 -12000 67350
rect -12100 67120 -12000 67150
rect -16000 67100 -15880 67120
rect -15620 67100 -15380 67120
rect -15120 67100 -14880 67120
rect -14620 67100 -14380 67120
rect -14120 67100 -13880 67120
rect -13620 67100 -13380 67120
rect -13120 67100 -12880 67120
rect -12620 67100 -12380 67120
rect -12120 67100 -12000 67120
rect -16000 67090 -12000 67100
rect -16000 67020 -15850 67090
rect -15650 67020 -15350 67090
rect -15150 67020 -14850 67090
rect -14650 67020 -14350 67090
rect -14150 67020 -13850 67090
rect -13650 67020 -13350 67090
rect -13150 67020 -12850 67090
rect -12650 67020 -12350 67090
rect -12150 67020 -12000 67090
rect -16000 66980 -12000 67020
rect -16000 66910 -15850 66980
rect -15650 66910 -15350 66980
rect -15150 66910 -14850 66980
rect -14650 66910 -14350 66980
rect -14150 66910 -13850 66980
rect -13650 66910 -13350 66980
rect -13150 66910 -12850 66980
rect -12650 66910 -12350 66980
rect -12150 66910 -12000 66980
rect -16000 66900 -12000 66910
rect -16000 66880 -15880 66900
rect -15620 66880 -15380 66900
rect -15120 66880 -14880 66900
rect -14620 66880 -14380 66900
rect -14120 66880 -13880 66900
rect -13620 66880 -13380 66900
rect -13120 66880 -12880 66900
rect -12620 66880 -12380 66900
rect -12120 66880 -12000 66900
rect -16000 66850 -15900 66880
rect -16000 66650 -15980 66850
rect -15910 66650 -15900 66850
rect -16000 66620 -15900 66650
rect -15600 66850 -15400 66880
rect -15600 66650 -15590 66850
rect -15520 66650 -15480 66850
rect -15410 66650 -15400 66850
rect -15600 66620 -15400 66650
rect -15100 66850 -14900 66880
rect -15100 66650 -15090 66850
rect -15020 66650 -14980 66850
rect -14910 66650 -14900 66850
rect -15100 66620 -14900 66650
rect -14600 66850 -14400 66880
rect -14600 66650 -14590 66850
rect -14520 66650 -14480 66850
rect -14410 66650 -14400 66850
rect -14600 66620 -14400 66650
rect -14100 66850 -13900 66880
rect -14100 66650 -14090 66850
rect -14020 66650 -13980 66850
rect -13910 66650 -13900 66850
rect -14100 66620 -13900 66650
rect -13600 66850 -13400 66880
rect -13600 66650 -13590 66850
rect -13520 66650 -13480 66850
rect -13410 66650 -13400 66850
rect -13600 66620 -13400 66650
rect -13100 66850 -12900 66880
rect -13100 66650 -13090 66850
rect -13020 66650 -12980 66850
rect -12910 66650 -12900 66850
rect -13100 66620 -12900 66650
rect -12600 66850 -12400 66880
rect -12600 66650 -12590 66850
rect -12520 66650 -12480 66850
rect -12410 66650 -12400 66850
rect -12600 66620 -12400 66650
rect -12100 66850 -12000 66880
rect -12100 66650 -12090 66850
rect -12020 66650 -12000 66850
rect -12100 66620 -12000 66650
rect -16000 66600 -15880 66620
rect -15620 66600 -15380 66620
rect -15120 66600 -14880 66620
rect -14620 66600 -14380 66620
rect -14120 66600 -13880 66620
rect -13620 66600 -13380 66620
rect -13120 66600 -12880 66620
rect -12620 66600 -12380 66620
rect -12120 66600 -12000 66620
rect -16000 66590 -12000 66600
rect -16000 66520 -15850 66590
rect -15650 66520 -15350 66590
rect -15150 66520 -14850 66590
rect -14650 66520 -14350 66590
rect -14150 66520 -13850 66590
rect -13650 66520 -13350 66590
rect -13150 66520 -12850 66590
rect -12650 66520 -12350 66590
rect -12150 66520 -12000 66590
rect -16000 66480 -12000 66520
rect -16000 66410 -15850 66480
rect -15650 66410 -15350 66480
rect -15150 66410 -14850 66480
rect -14650 66410 -14350 66480
rect -14150 66410 -13850 66480
rect -13650 66410 -13350 66480
rect -13150 66410 -12850 66480
rect -12650 66410 -12350 66480
rect -12150 66410 -12000 66480
rect -16000 66400 -12000 66410
rect -16000 66380 -15880 66400
rect -15620 66380 -15380 66400
rect -15120 66380 -14880 66400
rect -14620 66380 -14380 66400
rect -14120 66380 -13880 66400
rect -13620 66380 -13380 66400
rect -13120 66380 -12880 66400
rect -12620 66380 -12380 66400
rect -12120 66380 -12000 66400
rect -16000 66350 -15900 66380
rect -16000 66150 -15980 66350
rect -15910 66150 -15900 66350
rect -16000 66120 -15900 66150
rect -15600 66350 -15400 66380
rect -15600 66150 -15590 66350
rect -15520 66150 -15480 66350
rect -15410 66150 -15400 66350
rect -15600 66120 -15400 66150
rect -15100 66350 -14900 66380
rect -15100 66150 -15090 66350
rect -15020 66150 -14980 66350
rect -14910 66150 -14900 66350
rect -15100 66120 -14900 66150
rect -14600 66350 -14400 66380
rect -14600 66150 -14590 66350
rect -14520 66150 -14480 66350
rect -14410 66150 -14400 66350
rect -14600 66120 -14400 66150
rect -14100 66350 -13900 66380
rect -14100 66150 -14090 66350
rect -14020 66150 -13980 66350
rect -13910 66150 -13900 66350
rect -14100 66120 -13900 66150
rect -13600 66350 -13400 66380
rect -13600 66150 -13590 66350
rect -13520 66150 -13480 66350
rect -13410 66150 -13400 66350
rect -13600 66120 -13400 66150
rect -13100 66350 -12900 66380
rect -13100 66150 -13090 66350
rect -13020 66150 -12980 66350
rect -12910 66150 -12900 66350
rect -13100 66120 -12900 66150
rect -12600 66350 -12400 66380
rect -12600 66150 -12590 66350
rect -12520 66150 -12480 66350
rect -12410 66150 -12400 66350
rect -12600 66120 -12400 66150
rect -12100 66350 -12000 66380
rect -12100 66150 -12090 66350
rect -12020 66150 -12000 66350
rect -12100 66120 -12000 66150
rect -16000 66100 -15880 66120
rect -15620 66100 -15380 66120
rect -15120 66100 -14880 66120
rect -14620 66100 -14380 66120
rect -14120 66100 -13880 66120
rect -13620 66100 -13380 66120
rect -13120 66100 -12880 66120
rect -12620 66100 -12380 66120
rect -12120 66100 -12000 66120
rect -16000 66090 -12000 66100
rect -16000 66020 -15850 66090
rect -15650 66020 -15350 66090
rect -15150 66020 -14850 66090
rect -14650 66020 -14350 66090
rect -14150 66020 -13850 66090
rect -13650 66020 -13350 66090
rect -13150 66020 -12850 66090
rect -12650 66020 -12350 66090
rect -12150 66020 -12000 66090
rect -16000 65980 -12000 66020
rect -16000 65910 -15850 65980
rect -15650 65910 -15350 65980
rect -15150 65910 -14850 65980
rect -14650 65910 -14350 65980
rect -14150 65910 -13850 65980
rect -13650 65910 -13350 65980
rect -13150 65910 -12850 65980
rect -12650 65910 -12350 65980
rect -12150 65910 -12000 65980
rect -16000 65900 -12000 65910
rect -16000 65880 -15880 65900
rect -15620 65880 -15380 65900
rect -15120 65880 -14880 65900
rect -14620 65880 -14380 65900
rect -14120 65880 -13880 65900
rect -13620 65880 -13380 65900
rect -13120 65880 -12880 65900
rect -12620 65880 -12380 65900
rect -12120 65880 -12000 65900
rect -16000 65850 -15900 65880
rect -16000 65650 -15980 65850
rect -15910 65650 -15900 65850
rect -16000 65620 -15900 65650
rect -15600 65850 -15400 65880
rect -15600 65650 -15590 65850
rect -15520 65650 -15480 65850
rect -15410 65650 -15400 65850
rect -15600 65620 -15400 65650
rect -15100 65850 -14900 65880
rect -15100 65650 -15090 65850
rect -15020 65650 -14980 65850
rect -14910 65650 -14900 65850
rect -15100 65620 -14900 65650
rect -14600 65850 -14400 65880
rect -14600 65650 -14590 65850
rect -14520 65650 -14480 65850
rect -14410 65650 -14400 65850
rect -14600 65620 -14400 65650
rect -14100 65850 -13900 65880
rect -14100 65650 -14090 65850
rect -14020 65650 -13980 65850
rect -13910 65650 -13900 65850
rect -14100 65620 -13900 65650
rect -13600 65850 -13400 65880
rect -13600 65650 -13590 65850
rect -13520 65650 -13480 65850
rect -13410 65650 -13400 65850
rect -13600 65620 -13400 65650
rect -13100 65850 -12900 65880
rect -13100 65650 -13090 65850
rect -13020 65650 -12980 65850
rect -12910 65650 -12900 65850
rect -13100 65620 -12900 65650
rect -12600 65850 -12400 65880
rect -12600 65650 -12590 65850
rect -12520 65650 -12480 65850
rect -12410 65650 -12400 65850
rect -12600 65620 -12400 65650
rect -12100 65850 -12000 65880
rect -12100 65650 -12090 65850
rect -12020 65650 -12000 65850
rect -12100 65620 -12000 65650
rect -16000 65600 -15880 65620
rect -15620 65600 -15380 65620
rect -15120 65600 -14880 65620
rect -14620 65600 -14380 65620
rect -14120 65600 -13880 65620
rect -13620 65600 -13380 65620
rect -13120 65600 -12880 65620
rect -12620 65600 -12380 65620
rect -12120 65600 -12000 65620
rect -16000 65590 -12000 65600
rect -16000 65520 -15850 65590
rect -15650 65520 -15350 65590
rect -15150 65520 -14850 65590
rect -14650 65520 -14350 65590
rect -14150 65520 -13850 65590
rect -13650 65520 -13350 65590
rect -13150 65520 -12850 65590
rect -12650 65520 -12350 65590
rect -12150 65520 -12000 65590
rect -16000 65480 -12000 65520
rect -16000 65410 -15850 65480
rect -15650 65410 -15350 65480
rect -15150 65410 -14850 65480
rect -14650 65410 -14350 65480
rect -14150 65410 -13850 65480
rect -13650 65410 -13350 65480
rect -13150 65410 -12850 65480
rect -12650 65410 -12350 65480
rect -12150 65410 -12000 65480
rect -16000 65400 -12000 65410
rect -16000 65380 -15880 65400
rect -15620 65380 -15380 65400
rect -15120 65380 -14880 65400
rect -14620 65380 -14380 65400
rect -14120 65380 -13880 65400
rect -13620 65380 -13380 65400
rect -13120 65380 -12880 65400
rect -12620 65380 -12380 65400
rect -12120 65380 -12000 65400
rect -16000 65350 -15900 65380
rect -16000 65150 -15980 65350
rect -15910 65150 -15900 65350
rect -16000 65120 -15900 65150
rect -15600 65350 -15400 65380
rect -15600 65150 -15590 65350
rect -15520 65150 -15480 65350
rect -15410 65150 -15400 65350
rect -15600 65120 -15400 65150
rect -15100 65350 -14900 65380
rect -15100 65150 -15090 65350
rect -15020 65150 -14980 65350
rect -14910 65150 -14900 65350
rect -15100 65120 -14900 65150
rect -14600 65350 -14400 65380
rect -14600 65150 -14590 65350
rect -14520 65150 -14480 65350
rect -14410 65150 -14400 65350
rect -14600 65120 -14400 65150
rect -14100 65350 -13900 65380
rect -14100 65150 -14090 65350
rect -14020 65150 -13980 65350
rect -13910 65150 -13900 65350
rect -14100 65120 -13900 65150
rect -13600 65350 -13400 65380
rect -13600 65150 -13590 65350
rect -13520 65150 -13480 65350
rect -13410 65150 -13400 65350
rect -13600 65120 -13400 65150
rect -13100 65350 -12900 65380
rect -13100 65150 -13090 65350
rect -13020 65150 -12980 65350
rect -12910 65150 -12900 65350
rect -13100 65120 -12900 65150
rect -12600 65350 -12400 65380
rect -12600 65150 -12590 65350
rect -12520 65150 -12480 65350
rect -12410 65150 -12400 65350
rect -12600 65120 -12400 65150
rect -12100 65350 -12000 65380
rect -12100 65150 -12090 65350
rect -12020 65150 -12000 65350
rect -12100 65120 -12000 65150
rect -16000 65100 -15880 65120
rect -15620 65100 -15380 65120
rect -15120 65100 -14880 65120
rect -14620 65100 -14380 65120
rect -14120 65100 -13880 65120
rect -13620 65100 -13380 65120
rect -13120 65100 -12880 65120
rect -12620 65100 -12380 65120
rect -12120 65100 -12000 65120
rect -16000 65090 -12000 65100
rect -16000 65020 -15850 65090
rect -15650 65020 -15350 65090
rect -15150 65020 -14850 65090
rect -14650 65020 -14350 65090
rect -14150 65020 -13850 65090
rect -13650 65020 -13350 65090
rect -13150 65020 -12850 65090
rect -12650 65020 -12350 65090
rect -12150 65020 -12000 65090
rect -16000 64980 -12000 65020
rect -16000 64910 -15850 64980
rect -15650 64910 -15350 64980
rect -15150 64910 -14850 64980
rect -14650 64910 -14350 64980
rect -14150 64910 -13850 64980
rect -13650 64910 -13350 64980
rect -13150 64910 -12850 64980
rect -12650 64910 -12350 64980
rect -12150 64910 -12000 64980
rect -16000 64900 -12000 64910
rect -16000 64880 -15880 64900
rect -15620 64880 -15380 64900
rect -15120 64880 -14880 64900
rect -14620 64880 -14380 64900
rect -14120 64880 -13880 64900
rect -13620 64880 -13380 64900
rect -13120 64880 -12880 64900
rect -12620 64880 -12380 64900
rect -12120 64880 -12000 64900
rect -16000 64850 -15900 64880
rect -16000 64650 -15980 64850
rect -15910 64650 -15900 64850
rect -16000 64620 -15900 64650
rect -15600 64850 -15400 64880
rect -15600 64650 -15590 64850
rect -15520 64650 -15480 64850
rect -15410 64650 -15400 64850
rect -15600 64620 -15400 64650
rect -15100 64850 -14900 64880
rect -15100 64650 -15090 64850
rect -15020 64650 -14980 64850
rect -14910 64650 -14900 64850
rect -15100 64620 -14900 64650
rect -14600 64850 -14400 64880
rect -14600 64650 -14590 64850
rect -14520 64650 -14480 64850
rect -14410 64650 -14400 64850
rect -14600 64620 -14400 64650
rect -14100 64850 -13900 64880
rect -14100 64650 -14090 64850
rect -14020 64650 -13980 64850
rect -13910 64650 -13900 64850
rect -14100 64620 -13900 64650
rect -13600 64850 -13400 64880
rect -13600 64650 -13590 64850
rect -13520 64650 -13480 64850
rect -13410 64650 -13400 64850
rect -13600 64620 -13400 64650
rect -13100 64850 -12900 64880
rect -13100 64650 -13090 64850
rect -13020 64650 -12980 64850
rect -12910 64650 -12900 64850
rect -13100 64620 -12900 64650
rect -12600 64850 -12400 64880
rect -12600 64650 -12590 64850
rect -12520 64650 -12480 64850
rect -12410 64650 -12400 64850
rect -12600 64620 -12400 64650
rect -12100 64850 -12000 64880
rect -12100 64650 -12090 64850
rect -12020 64650 -12000 64850
rect -12100 64620 -12000 64650
rect -16000 64600 -15880 64620
rect -15620 64600 -15380 64620
rect -15120 64600 -14880 64620
rect -14620 64600 -14380 64620
rect -14120 64600 -13880 64620
rect -13620 64600 -13380 64620
rect -13120 64600 -12880 64620
rect -12620 64600 -12380 64620
rect -12120 64600 -12000 64620
rect -16000 64590 -12000 64600
rect -16000 64520 -15850 64590
rect -15650 64520 -15350 64590
rect -15150 64520 -14850 64590
rect -14650 64520 -14350 64590
rect -14150 64520 -13850 64590
rect -13650 64520 -13350 64590
rect -13150 64520 -12850 64590
rect -12650 64520 -12350 64590
rect -12150 64520 -12000 64590
rect -16000 64480 -12000 64520
rect -16000 64410 -15850 64480
rect -15650 64410 -15350 64480
rect -15150 64410 -14850 64480
rect -14650 64410 -14350 64480
rect -14150 64410 -13850 64480
rect -13650 64410 -13350 64480
rect -13150 64410 -12850 64480
rect -12650 64410 -12350 64480
rect -12150 64410 -12000 64480
rect -16000 64400 -12000 64410
rect -16000 64380 -15880 64400
rect -15620 64380 -15380 64400
rect -15120 64380 -14880 64400
rect -14620 64380 -14380 64400
rect -14120 64380 -13880 64400
rect -13620 64380 -13380 64400
rect -13120 64380 -12880 64400
rect -12620 64380 -12380 64400
rect -12120 64380 -12000 64400
rect -16000 64350 -15900 64380
rect -16000 64150 -15980 64350
rect -15910 64150 -15900 64350
rect -16000 64120 -15900 64150
rect -15600 64350 -15400 64380
rect -15600 64150 -15590 64350
rect -15520 64150 -15480 64350
rect -15410 64150 -15400 64350
rect -15600 64120 -15400 64150
rect -15100 64350 -14900 64380
rect -15100 64150 -15090 64350
rect -15020 64150 -14980 64350
rect -14910 64150 -14900 64350
rect -15100 64120 -14900 64150
rect -14600 64350 -14400 64380
rect -14600 64150 -14590 64350
rect -14520 64150 -14480 64350
rect -14410 64150 -14400 64350
rect -14600 64120 -14400 64150
rect -14100 64350 -13900 64380
rect -14100 64150 -14090 64350
rect -14020 64150 -13980 64350
rect -13910 64150 -13900 64350
rect -14100 64120 -13900 64150
rect -13600 64350 -13400 64380
rect -13600 64150 -13590 64350
rect -13520 64150 -13480 64350
rect -13410 64150 -13400 64350
rect -13600 64120 -13400 64150
rect -13100 64350 -12900 64380
rect -13100 64150 -13090 64350
rect -13020 64150 -12980 64350
rect -12910 64150 -12900 64350
rect -13100 64120 -12900 64150
rect -12600 64350 -12400 64380
rect -12600 64150 -12590 64350
rect -12520 64150 -12480 64350
rect -12410 64150 -12400 64350
rect -12600 64120 -12400 64150
rect -12100 64350 -12000 64380
rect -12100 64150 -12090 64350
rect -12020 64150 -12000 64350
rect -12100 64120 -12000 64150
rect -16000 64100 -15880 64120
rect -15620 64100 -15380 64120
rect -15120 64100 -14880 64120
rect -14620 64100 -14380 64120
rect -14120 64100 -13880 64120
rect -13620 64100 -13380 64120
rect -13120 64100 -12880 64120
rect -12620 64100 -12380 64120
rect -12120 64100 -12000 64120
rect -16000 64090 -12000 64100
rect -16000 64020 -15850 64090
rect -15650 64020 -15350 64090
rect -15150 64020 -14850 64090
rect -14650 64020 -14350 64090
rect -14150 64020 -13850 64090
rect -13650 64020 -13350 64090
rect -13150 64020 -12850 64090
rect -12650 64020 -12350 64090
rect -12150 64020 -12000 64090
rect -16000 63980 -12000 64020
rect -16000 63910 -15850 63980
rect -15650 63910 -15350 63980
rect -15150 63910 -14850 63980
rect -14650 63910 -14350 63980
rect -14150 63910 -13850 63980
rect -13650 63910 -13350 63980
rect -13150 63910 -12850 63980
rect -12650 63910 -12350 63980
rect -12150 63910 -12000 63980
rect -16000 63900 -12000 63910
rect -16000 63880 -15880 63900
rect -15620 63880 -15380 63900
rect -15120 63880 -14880 63900
rect -14620 63880 -14380 63900
rect -14120 63880 -13880 63900
rect -13620 63880 -13380 63900
rect -13120 63880 -12880 63900
rect -12620 63880 -12380 63900
rect -12120 63880 -12000 63900
rect -16000 63850 -15900 63880
rect -16000 63650 -15980 63850
rect -15910 63650 -15900 63850
rect -16000 63620 -15900 63650
rect -15600 63850 -15400 63880
rect -15600 63650 -15590 63850
rect -15520 63650 -15480 63850
rect -15410 63650 -15400 63850
rect -15600 63620 -15400 63650
rect -15100 63850 -14900 63880
rect -15100 63650 -15090 63850
rect -15020 63650 -14980 63850
rect -14910 63650 -14900 63850
rect -15100 63620 -14900 63650
rect -14600 63850 -14400 63880
rect -14600 63650 -14590 63850
rect -14520 63650 -14480 63850
rect -14410 63650 -14400 63850
rect -14600 63620 -14400 63650
rect -14100 63850 -13900 63880
rect -14100 63650 -14090 63850
rect -14020 63650 -13980 63850
rect -13910 63650 -13900 63850
rect -14100 63620 -13900 63650
rect -13600 63850 -13400 63880
rect -13600 63650 -13590 63850
rect -13520 63650 -13480 63850
rect -13410 63650 -13400 63850
rect -13600 63620 -13400 63650
rect -13100 63850 -12900 63880
rect -13100 63650 -13090 63850
rect -13020 63650 -12980 63850
rect -12910 63650 -12900 63850
rect -13100 63620 -12900 63650
rect -12600 63850 -12400 63880
rect -12600 63650 -12590 63850
rect -12520 63650 -12480 63850
rect -12410 63650 -12400 63850
rect -12600 63620 -12400 63650
rect -12100 63850 -12000 63880
rect -12100 63650 -12090 63850
rect -12020 63650 -12000 63850
rect -12100 63620 -12000 63650
rect -16000 63600 -15880 63620
rect -15620 63600 -15380 63620
rect -15120 63600 -14880 63620
rect -14620 63600 -14380 63620
rect -14120 63600 -13880 63620
rect -13620 63600 -13380 63620
rect -13120 63600 -12880 63620
rect -12620 63600 -12380 63620
rect -12120 63600 -12000 63620
rect -16000 63590 -12000 63600
rect -16000 63520 -15850 63590
rect -15650 63520 -15350 63590
rect -15150 63520 -14850 63590
rect -14650 63520 -14350 63590
rect -14150 63520 -13850 63590
rect -13650 63520 -13350 63590
rect -13150 63520 -12850 63590
rect -12650 63520 -12350 63590
rect -12150 63520 -12000 63590
rect -16000 63480 -12000 63520
rect -16000 63410 -15850 63480
rect -15650 63410 -15350 63480
rect -15150 63410 -14850 63480
rect -14650 63410 -14350 63480
rect -14150 63410 -13850 63480
rect -13650 63410 -13350 63480
rect -13150 63410 -12850 63480
rect -12650 63410 -12350 63480
rect -12150 63410 -12000 63480
rect -16000 63400 -12000 63410
rect -16000 63380 -15880 63400
rect -15620 63380 -15380 63400
rect -15120 63380 -14880 63400
rect -14620 63380 -14380 63400
rect -14120 63380 -13880 63400
rect -13620 63380 -13380 63400
rect -13120 63380 -12880 63400
rect -12620 63380 -12380 63400
rect -12120 63380 -12000 63400
rect -16000 63350 -15900 63380
rect -16000 63150 -15980 63350
rect -15910 63150 -15900 63350
rect -16000 63120 -15900 63150
rect -15600 63350 -15400 63380
rect -15600 63150 -15590 63350
rect -15520 63150 -15480 63350
rect -15410 63150 -15400 63350
rect -15600 63120 -15400 63150
rect -15100 63350 -14900 63380
rect -15100 63150 -15090 63350
rect -15020 63150 -14980 63350
rect -14910 63150 -14900 63350
rect -15100 63120 -14900 63150
rect -14600 63350 -14400 63380
rect -14600 63150 -14590 63350
rect -14520 63150 -14480 63350
rect -14410 63150 -14400 63350
rect -14600 63120 -14400 63150
rect -14100 63350 -13900 63380
rect -14100 63150 -14090 63350
rect -14020 63150 -13980 63350
rect -13910 63150 -13900 63350
rect -14100 63120 -13900 63150
rect -13600 63350 -13400 63380
rect -13600 63150 -13590 63350
rect -13520 63150 -13480 63350
rect -13410 63150 -13400 63350
rect -13600 63120 -13400 63150
rect -13100 63350 -12900 63380
rect -13100 63150 -13090 63350
rect -13020 63150 -12980 63350
rect -12910 63150 -12900 63350
rect -13100 63120 -12900 63150
rect -12600 63350 -12400 63380
rect -12600 63150 -12590 63350
rect -12520 63150 -12480 63350
rect -12410 63150 -12400 63350
rect -12600 63120 -12400 63150
rect -12100 63350 -12000 63380
rect -12100 63150 -12090 63350
rect -12020 63150 -12000 63350
rect -12100 63120 -12000 63150
rect -16000 63100 -15880 63120
rect -15620 63100 -15380 63120
rect -15120 63100 -14880 63120
rect -14620 63100 -14380 63120
rect -14120 63100 -13880 63120
rect -13620 63100 -13380 63120
rect -13120 63100 -12880 63120
rect -12620 63100 -12380 63120
rect -12120 63100 -12000 63120
rect -16000 63090 -12000 63100
rect -16000 63020 -15850 63090
rect -15650 63020 -15350 63090
rect -15150 63020 -14850 63090
rect -14650 63020 -14350 63090
rect -14150 63020 -13850 63090
rect -13650 63020 -13350 63090
rect -13150 63020 -12850 63090
rect -12650 63020 -12350 63090
rect -12150 63020 -12000 63090
rect -16000 62980 -12000 63020
rect -16000 62910 -15850 62980
rect -15650 62910 -15350 62980
rect -15150 62910 -14850 62980
rect -14650 62910 -14350 62980
rect -14150 62910 -13850 62980
rect -13650 62910 -13350 62980
rect -13150 62910 -12850 62980
rect -12650 62910 -12350 62980
rect -12150 62910 -12000 62980
rect -16000 62900 -12000 62910
rect -16000 62880 -15880 62900
rect -15620 62880 -15380 62900
rect -15120 62880 -14880 62900
rect -14620 62880 -14380 62900
rect -14120 62880 -13880 62900
rect -13620 62880 -13380 62900
rect -13120 62880 -12880 62900
rect -12620 62880 -12380 62900
rect -12120 62880 -12000 62900
rect -16000 62850 -15900 62880
rect -16000 62650 -15980 62850
rect -15910 62650 -15900 62850
rect -16000 62620 -15900 62650
rect -15600 62850 -15400 62880
rect -15600 62650 -15590 62850
rect -15520 62650 -15480 62850
rect -15410 62650 -15400 62850
rect -15600 62620 -15400 62650
rect -15100 62850 -14900 62880
rect -15100 62650 -15090 62850
rect -15020 62650 -14980 62850
rect -14910 62650 -14900 62850
rect -15100 62620 -14900 62650
rect -14600 62850 -14400 62880
rect -14600 62650 -14590 62850
rect -14520 62650 -14480 62850
rect -14410 62650 -14400 62850
rect -14600 62620 -14400 62650
rect -14100 62850 -13900 62880
rect -14100 62650 -14090 62850
rect -14020 62650 -13980 62850
rect -13910 62650 -13900 62850
rect -14100 62620 -13900 62650
rect -13600 62850 -13400 62880
rect -13600 62650 -13590 62850
rect -13520 62650 -13480 62850
rect -13410 62650 -13400 62850
rect -13600 62620 -13400 62650
rect -13100 62850 -12900 62880
rect -13100 62650 -13090 62850
rect -13020 62650 -12980 62850
rect -12910 62650 -12900 62850
rect -13100 62620 -12900 62650
rect -12600 62850 -12400 62880
rect -12600 62650 -12590 62850
rect -12520 62650 -12480 62850
rect -12410 62650 -12400 62850
rect -12600 62620 -12400 62650
rect -12100 62850 -12000 62880
rect -12100 62650 -12090 62850
rect -12020 62650 -12000 62850
rect -12100 62620 -12000 62650
rect -16000 62600 -15880 62620
rect -15620 62600 -15380 62620
rect -15120 62600 -14880 62620
rect -14620 62600 -14380 62620
rect -14120 62600 -13880 62620
rect -13620 62600 -13380 62620
rect -13120 62600 -12880 62620
rect -12620 62600 -12380 62620
rect -12120 62600 -12000 62620
rect -16000 62590 -12000 62600
rect -16000 62520 -15850 62590
rect -15650 62520 -15350 62590
rect -15150 62520 -14850 62590
rect -14650 62520 -14350 62590
rect -14150 62520 -13850 62590
rect -13650 62520 -13350 62590
rect -13150 62520 -12850 62590
rect -12650 62520 -12350 62590
rect -12150 62520 -12000 62590
rect -16000 62480 -12000 62520
rect -16000 62410 -15850 62480
rect -15650 62410 -15350 62480
rect -15150 62410 -14850 62480
rect -14650 62410 -14350 62480
rect -14150 62410 -13850 62480
rect -13650 62410 -13350 62480
rect -13150 62410 -12850 62480
rect -12650 62410 -12350 62480
rect -12150 62410 -12000 62480
rect -16000 62400 -12000 62410
rect -16000 62380 -15880 62400
rect -15620 62380 -15380 62400
rect -15120 62380 -14880 62400
rect -14620 62380 -14380 62400
rect -14120 62380 -13880 62400
rect -13620 62380 -13380 62400
rect -13120 62380 -12880 62400
rect -12620 62380 -12380 62400
rect -12120 62380 -12000 62400
rect -16000 62350 -15900 62380
rect -16000 62150 -15980 62350
rect -15910 62150 -15900 62350
rect -16000 62120 -15900 62150
rect -15600 62350 -15400 62380
rect -15600 62150 -15590 62350
rect -15520 62150 -15480 62350
rect -15410 62150 -15400 62350
rect -15600 62120 -15400 62150
rect -15100 62350 -14900 62380
rect -15100 62150 -15090 62350
rect -15020 62150 -14980 62350
rect -14910 62150 -14900 62350
rect -15100 62120 -14900 62150
rect -14600 62350 -14400 62380
rect -14600 62150 -14590 62350
rect -14520 62150 -14480 62350
rect -14410 62150 -14400 62350
rect -14600 62120 -14400 62150
rect -14100 62350 -13900 62380
rect -14100 62150 -14090 62350
rect -14020 62150 -13980 62350
rect -13910 62150 -13900 62350
rect -14100 62120 -13900 62150
rect -13600 62350 -13400 62380
rect -13600 62150 -13590 62350
rect -13520 62150 -13480 62350
rect -13410 62150 -13400 62350
rect -13600 62120 -13400 62150
rect -13100 62350 -12900 62380
rect -13100 62150 -13090 62350
rect -13020 62150 -12980 62350
rect -12910 62150 -12900 62350
rect -13100 62120 -12900 62150
rect -12600 62350 -12400 62380
rect -12600 62150 -12590 62350
rect -12520 62150 -12480 62350
rect -12410 62150 -12400 62350
rect -12600 62120 -12400 62150
rect -12100 62350 -12000 62380
rect -12100 62150 -12090 62350
rect -12020 62150 -12000 62350
rect -12100 62120 -12000 62150
rect -16000 62100 -15880 62120
rect -15620 62100 -15380 62120
rect -15120 62100 -14880 62120
rect -14620 62100 -14380 62120
rect -14120 62100 -13880 62120
rect -13620 62100 -13380 62120
rect -13120 62100 -12880 62120
rect -12620 62100 -12380 62120
rect -12120 62100 -12000 62120
rect -16000 62090 -12000 62100
rect -16000 62020 -15850 62090
rect -15650 62020 -15350 62090
rect -15150 62020 -14850 62090
rect -14650 62020 -14350 62090
rect -14150 62020 -13850 62090
rect -13650 62020 -13350 62090
rect -13150 62020 -12850 62090
rect -12650 62020 -12350 62090
rect -12150 62020 -12000 62090
rect -16000 61980 -12000 62020
rect -16000 61910 -15850 61980
rect -15650 61910 -15350 61980
rect -15150 61910 -14850 61980
rect -14650 61910 -14350 61980
rect -14150 61910 -13850 61980
rect -13650 61910 -13350 61980
rect -13150 61910 -12850 61980
rect -12650 61910 -12350 61980
rect -12150 61910 -12000 61980
rect -16000 61900 -12000 61910
rect -16000 61880 -15880 61900
rect -15620 61880 -15380 61900
rect -15120 61880 -14880 61900
rect -14620 61880 -14380 61900
rect -14120 61880 -13880 61900
rect -13620 61880 -13380 61900
rect -13120 61880 -12880 61900
rect -12620 61880 -12380 61900
rect -12120 61880 -12000 61900
rect -16000 61850 -15900 61880
rect -16000 61650 -15980 61850
rect -15910 61650 -15900 61850
rect -16000 61620 -15900 61650
rect -15600 61850 -15400 61880
rect -15600 61650 -15590 61850
rect -15520 61650 -15480 61850
rect -15410 61650 -15400 61850
rect -15600 61620 -15400 61650
rect -15100 61850 -14900 61880
rect -15100 61650 -15090 61850
rect -15020 61650 -14980 61850
rect -14910 61650 -14900 61850
rect -15100 61620 -14900 61650
rect -14600 61850 -14400 61880
rect -14600 61650 -14590 61850
rect -14520 61650 -14480 61850
rect -14410 61650 -14400 61850
rect -14600 61620 -14400 61650
rect -14100 61850 -13900 61880
rect -14100 61650 -14090 61850
rect -14020 61650 -13980 61850
rect -13910 61650 -13900 61850
rect -14100 61620 -13900 61650
rect -13600 61850 -13400 61880
rect -13600 61650 -13590 61850
rect -13520 61650 -13480 61850
rect -13410 61650 -13400 61850
rect -13600 61620 -13400 61650
rect -13100 61850 -12900 61880
rect -13100 61650 -13090 61850
rect -13020 61650 -12980 61850
rect -12910 61650 -12900 61850
rect -13100 61620 -12900 61650
rect -12600 61850 -12400 61880
rect -12600 61650 -12590 61850
rect -12520 61650 -12480 61850
rect -12410 61650 -12400 61850
rect -12600 61620 -12400 61650
rect -12100 61850 -12000 61880
rect -12100 61650 -12090 61850
rect -12020 61650 -12000 61850
rect -12100 61620 -12000 61650
rect -16000 61600 -15880 61620
rect -15620 61600 -15380 61620
rect -15120 61600 -14880 61620
rect -14620 61600 -14380 61620
rect -14120 61600 -13880 61620
rect -13620 61600 -13380 61620
rect -13120 61600 -12880 61620
rect -12620 61600 -12380 61620
rect -12120 61600 -12000 61620
rect -16000 61590 -12000 61600
rect -16000 61520 -15850 61590
rect -15650 61520 -15350 61590
rect -15150 61520 -14850 61590
rect -14650 61520 -14350 61590
rect -14150 61520 -13850 61590
rect -13650 61520 -13350 61590
rect -13150 61520 -12850 61590
rect -12650 61520 -12350 61590
rect -12150 61520 -12000 61590
rect -16000 61480 -12000 61520
rect -16000 61410 -15850 61480
rect -15650 61410 -15350 61480
rect -15150 61410 -14850 61480
rect -14650 61410 -14350 61480
rect -14150 61410 -13850 61480
rect -13650 61410 -13350 61480
rect -13150 61410 -12850 61480
rect -12650 61410 -12350 61480
rect -12150 61410 -12000 61480
rect -16000 61400 -12000 61410
rect -16000 61380 -15880 61400
rect -15620 61380 -15380 61400
rect -15120 61380 -14880 61400
rect -14620 61380 -14380 61400
rect -14120 61380 -13880 61400
rect -13620 61380 -13380 61400
rect -13120 61380 -12880 61400
rect -12620 61380 -12380 61400
rect -12120 61380 -12000 61400
rect -16000 61350 -15900 61380
rect -16000 61150 -15980 61350
rect -15910 61150 -15900 61350
rect -16000 61120 -15900 61150
rect -15600 61350 -15400 61380
rect -15600 61150 -15590 61350
rect -15520 61150 -15480 61350
rect -15410 61150 -15400 61350
rect -15600 61120 -15400 61150
rect -15100 61350 -14900 61380
rect -15100 61150 -15090 61350
rect -15020 61150 -14980 61350
rect -14910 61150 -14900 61350
rect -15100 61120 -14900 61150
rect -14600 61350 -14400 61380
rect -14600 61150 -14590 61350
rect -14520 61150 -14480 61350
rect -14410 61150 -14400 61350
rect -14600 61120 -14400 61150
rect -14100 61350 -13900 61380
rect -14100 61150 -14090 61350
rect -14020 61150 -13980 61350
rect -13910 61150 -13900 61350
rect -14100 61120 -13900 61150
rect -13600 61350 -13400 61380
rect -13600 61150 -13590 61350
rect -13520 61150 -13480 61350
rect -13410 61150 -13400 61350
rect -13600 61120 -13400 61150
rect -13100 61350 -12900 61380
rect -13100 61150 -13090 61350
rect -13020 61150 -12980 61350
rect -12910 61150 -12900 61350
rect -13100 61120 -12900 61150
rect -12600 61350 -12400 61380
rect -12600 61150 -12590 61350
rect -12520 61150 -12480 61350
rect -12410 61150 -12400 61350
rect -12600 61120 -12400 61150
rect -12100 61350 -12000 61380
rect -12100 61150 -12090 61350
rect -12020 61150 -12000 61350
rect -12100 61120 -12000 61150
rect -16000 61100 -15880 61120
rect -15620 61100 -15380 61120
rect -15120 61100 -14880 61120
rect -14620 61100 -14380 61120
rect -14120 61100 -13880 61120
rect -13620 61100 -13380 61120
rect -13120 61100 -12880 61120
rect -12620 61100 -12380 61120
rect -12120 61100 -12000 61120
rect -16000 61090 -12000 61100
rect -16000 61020 -15850 61090
rect -15650 61020 -15350 61090
rect -15150 61020 -14850 61090
rect -14650 61020 -14350 61090
rect -14150 61020 -13850 61090
rect -13650 61020 -13350 61090
rect -13150 61020 -12850 61090
rect -12650 61020 -12350 61090
rect -12150 61020 -12000 61090
rect -16000 60980 -12000 61020
rect -16000 60910 -15850 60980
rect -15650 60910 -15350 60980
rect -15150 60910 -14850 60980
rect -14650 60910 -14350 60980
rect -14150 60910 -13850 60980
rect -13650 60910 -13350 60980
rect -13150 60910 -12850 60980
rect -12650 60910 -12350 60980
rect -12150 60910 -12000 60980
rect -16000 60900 -12000 60910
rect -16000 60880 -15880 60900
rect -15620 60880 -15380 60900
rect -15120 60880 -14880 60900
rect -14620 60880 -14380 60900
rect -14120 60880 -13880 60900
rect -13620 60880 -13380 60900
rect -13120 60880 -12880 60900
rect -12620 60880 -12380 60900
rect -12120 60880 -12000 60900
rect -16000 60850 -15900 60880
rect -16000 60650 -15980 60850
rect -15910 60650 -15900 60850
rect -16000 60620 -15900 60650
rect -15600 60850 -15400 60880
rect -15600 60650 -15590 60850
rect -15520 60650 -15480 60850
rect -15410 60650 -15400 60850
rect -15600 60620 -15400 60650
rect -15100 60850 -14900 60880
rect -15100 60650 -15090 60850
rect -15020 60650 -14980 60850
rect -14910 60650 -14900 60850
rect -15100 60620 -14900 60650
rect -14600 60850 -14400 60880
rect -14600 60650 -14590 60850
rect -14520 60650 -14480 60850
rect -14410 60650 -14400 60850
rect -14600 60620 -14400 60650
rect -14100 60850 -13900 60880
rect -14100 60650 -14090 60850
rect -14020 60650 -13980 60850
rect -13910 60650 -13900 60850
rect -14100 60620 -13900 60650
rect -13600 60850 -13400 60880
rect -13600 60650 -13590 60850
rect -13520 60650 -13480 60850
rect -13410 60650 -13400 60850
rect -13600 60620 -13400 60650
rect -13100 60850 -12900 60880
rect -13100 60650 -13090 60850
rect -13020 60650 -12980 60850
rect -12910 60650 -12900 60850
rect -13100 60620 -12900 60650
rect -12600 60850 -12400 60880
rect -12600 60650 -12590 60850
rect -12520 60650 -12480 60850
rect -12410 60650 -12400 60850
rect -12600 60620 -12400 60650
rect -12100 60850 -12000 60880
rect -12100 60650 -12090 60850
rect -12020 60650 -12000 60850
rect -12100 60620 -12000 60650
rect -16000 60600 -15880 60620
rect -15620 60600 -15380 60620
rect -15120 60600 -14880 60620
rect -14620 60600 -14380 60620
rect -14120 60600 -13880 60620
rect -13620 60600 -13380 60620
rect -13120 60600 -12880 60620
rect -12620 60600 -12380 60620
rect -12120 60600 -12000 60620
rect -16000 60590 -12000 60600
rect -16000 60520 -15850 60590
rect -15650 60520 -15350 60590
rect -15150 60520 -14850 60590
rect -14650 60520 -14350 60590
rect -14150 60520 -13850 60590
rect -13650 60520 -13350 60590
rect -13150 60520 -12850 60590
rect -12650 60520 -12350 60590
rect -12150 60520 -12000 60590
rect -16000 60480 -12000 60520
rect -16000 60410 -15850 60480
rect -15650 60410 -15350 60480
rect -15150 60410 -14850 60480
rect -14650 60410 -14350 60480
rect -14150 60410 -13850 60480
rect -13650 60410 -13350 60480
rect -13150 60410 -12850 60480
rect -12650 60410 -12350 60480
rect -12150 60410 -12000 60480
rect -16000 60400 -12000 60410
rect -16000 60380 -15880 60400
rect -15620 60380 -15380 60400
rect -15120 60380 -14880 60400
rect -14620 60380 -14380 60400
rect -14120 60380 -13880 60400
rect -13620 60380 -13380 60400
rect -13120 60380 -12880 60400
rect -12620 60380 -12380 60400
rect -12120 60380 -12000 60400
rect -16000 60350 -15900 60380
rect -16000 60150 -15980 60350
rect -15910 60150 -15900 60350
rect -16000 60120 -15900 60150
rect -15600 60350 -15400 60380
rect -15600 60150 -15590 60350
rect -15520 60150 -15480 60350
rect -15410 60150 -15400 60350
rect -15600 60120 -15400 60150
rect -15100 60350 -14900 60380
rect -15100 60150 -15090 60350
rect -15020 60150 -14980 60350
rect -14910 60150 -14900 60350
rect -15100 60120 -14900 60150
rect -14600 60350 -14400 60380
rect -14600 60150 -14590 60350
rect -14520 60150 -14480 60350
rect -14410 60150 -14400 60350
rect -14600 60120 -14400 60150
rect -14100 60350 -13900 60380
rect -14100 60150 -14090 60350
rect -14020 60150 -13980 60350
rect -13910 60150 -13900 60350
rect -14100 60120 -13900 60150
rect -13600 60350 -13400 60380
rect -13600 60150 -13590 60350
rect -13520 60150 -13480 60350
rect -13410 60150 -13400 60350
rect -13600 60120 -13400 60150
rect -13100 60350 -12900 60380
rect -13100 60150 -13090 60350
rect -13020 60150 -12980 60350
rect -12910 60150 -12900 60350
rect -13100 60120 -12900 60150
rect -12600 60350 -12400 60380
rect -12600 60150 -12590 60350
rect -12520 60150 -12480 60350
rect -12410 60150 -12400 60350
rect -12600 60120 -12400 60150
rect -12100 60350 -12000 60380
rect -12100 60150 -12090 60350
rect -12020 60150 -12000 60350
rect -12100 60120 -12000 60150
rect -16000 60100 -15880 60120
rect -15620 60100 -15380 60120
rect -15120 60100 -14880 60120
rect -14620 60100 -14380 60120
rect -14120 60100 -13880 60120
rect -13620 60100 -13380 60120
rect -13120 60100 -12880 60120
rect -12620 60100 -12380 60120
rect -12120 60100 -12000 60120
rect -16000 60090 -12000 60100
rect -16000 60020 -15850 60090
rect -15650 60020 -15350 60090
rect -15150 60020 -14850 60090
rect -14650 60020 -14350 60090
rect -14150 60020 -13850 60090
rect -13650 60020 -13350 60090
rect -13150 60020 -12850 60090
rect -12650 60020 -12350 60090
rect -12150 60020 -12000 60090
rect -16000 59980 -12000 60020
rect -16000 59910 -15850 59980
rect -15650 59910 -15350 59980
rect -15150 59910 -14850 59980
rect -14650 59910 -14350 59980
rect -14150 59910 -13850 59980
rect -13650 59910 -13350 59980
rect -13150 59910 -12850 59980
rect -12650 59910 -12350 59980
rect -12150 59910 -12000 59980
rect -16000 59900 -12000 59910
rect -16000 59880 -15880 59900
rect -15620 59880 -15380 59900
rect -15120 59880 -14880 59900
rect -14620 59880 -14380 59900
rect -14120 59880 -13880 59900
rect -13620 59880 -13380 59900
rect -13120 59880 -12880 59900
rect -12620 59880 -12380 59900
rect -12120 59880 -12000 59900
rect -16000 59850 -15900 59880
rect -16000 59650 -15980 59850
rect -15910 59650 -15900 59850
rect -16000 59620 -15900 59650
rect -15600 59850 -15400 59880
rect -15600 59650 -15590 59850
rect -15520 59650 -15480 59850
rect -15410 59650 -15400 59850
rect -15600 59620 -15400 59650
rect -15100 59850 -14900 59880
rect -15100 59650 -15090 59850
rect -15020 59650 -14980 59850
rect -14910 59650 -14900 59850
rect -15100 59620 -14900 59650
rect -14600 59850 -14400 59880
rect -14600 59650 -14590 59850
rect -14520 59650 -14480 59850
rect -14410 59650 -14400 59850
rect -14600 59620 -14400 59650
rect -14100 59850 -13900 59880
rect -14100 59650 -14090 59850
rect -14020 59650 -13980 59850
rect -13910 59650 -13900 59850
rect -14100 59620 -13900 59650
rect -13600 59850 -13400 59880
rect -13600 59650 -13590 59850
rect -13520 59650 -13480 59850
rect -13410 59650 -13400 59850
rect -13600 59620 -13400 59650
rect -13100 59850 -12900 59880
rect -13100 59650 -13090 59850
rect -13020 59650 -12980 59850
rect -12910 59650 -12900 59850
rect -13100 59620 -12900 59650
rect -12600 59850 -12400 59880
rect -12600 59650 -12590 59850
rect -12520 59650 -12480 59850
rect -12410 59650 -12400 59850
rect -12600 59620 -12400 59650
rect -12100 59850 -12000 59880
rect -12100 59650 -12090 59850
rect -12020 59650 -12000 59850
rect -12100 59620 -12000 59650
rect -16000 59600 -15880 59620
rect -15620 59600 -15380 59620
rect -15120 59600 -14880 59620
rect -14620 59600 -14380 59620
rect -14120 59600 -13880 59620
rect -13620 59600 -13380 59620
rect -13120 59600 -12880 59620
rect -12620 59600 -12380 59620
rect -12120 59600 -12000 59620
rect -16000 59590 -12000 59600
rect -16000 59520 -15850 59590
rect -15650 59520 -15350 59590
rect -15150 59520 -14850 59590
rect -14650 59520 -14350 59590
rect -14150 59520 -13850 59590
rect -13650 59520 -13350 59590
rect -13150 59520 -12850 59590
rect -12650 59520 -12350 59590
rect -12150 59520 -12000 59590
rect -16000 59480 -12000 59520
rect -16000 59410 -15850 59480
rect -15650 59410 -15350 59480
rect -15150 59410 -14850 59480
rect -14650 59410 -14350 59480
rect -14150 59410 -13850 59480
rect -13650 59410 -13350 59480
rect -13150 59410 -12850 59480
rect -12650 59410 -12350 59480
rect -12150 59410 -12000 59480
rect -16000 59400 -12000 59410
rect -16000 59380 -15880 59400
rect -15620 59380 -15380 59400
rect -15120 59380 -14880 59400
rect -14620 59380 -14380 59400
rect -14120 59380 -13880 59400
rect -13620 59380 -13380 59400
rect -13120 59380 -12880 59400
rect -12620 59380 -12380 59400
rect -12120 59380 -12000 59400
rect -16000 59350 -15900 59380
rect -16000 59150 -15980 59350
rect -15910 59150 -15900 59350
rect -16000 59120 -15900 59150
rect -15600 59350 -15400 59380
rect -15600 59150 -15590 59350
rect -15520 59150 -15480 59350
rect -15410 59150 -15400 59350
rect -15600 59120 -15400 59150
rect -15100 59350 -14900 59380
rect -15100 59150 -15090 59350
rect -15020 59150 -14980 59350
rect -14910 59150 -14900 59350
rect -15100 59120 -14900 59150
rect -14600 59350 -14400 59380
rect -14600 59150 -14590 59350
rect -14520 59150 -14480 59350
rect -14410 59150 -14400 59350
rect -14600 59120 -14400 59150
rect -14100 59350 -13900 59380
rect -14100 59150 -14090 59350
rect -14020 59150 -13980 59350
rect -13910 59150 -13900 59350
rect -14100 59120 -13900 59150
rect -13600 59350 -13400 59380
rect -13600 59150 -13590 59350
rect -13520 59150 -13480 59350
rect -13410 59150 -13400 59350
rect -13600 59120 -13400 59150
rect -13100 59350 -12900 59380
rect -13100 59150 -13090 59350
rect -13020 59150 -12980 59350
rect -12910 59150 -12900 59350
rect -13100 59120 -12900 59150
rect -12600 59350 -12400 59380
rect -12600 59150 -12590 59350
rect -12520 59150 -12480 59350
rect -12410 59150 -12400 59350
rect -12600 59120 -12400 59150
rect -12100 59350 -12000 59380
rect -12100 59150 -12090 59350
rect -12020 59150 -12000 59350
rect -12100 59120 -12000 59150
rect -16000 59100 -15880 59120
rect -15620 59100 -15380 59120
rect -15120 59100 -14880 59120
rect -14620 59100 -14380 59120
rect -14120 59100 -13880 59120
rect -13620 59100 -13380 59120
rect -13120 59100 -12880 59120
rect -12620 59100 -12380 59120
rect -12120 59100 -12000 59120
rect -16000 59090 -12000 59100
rect -16000 59020 -15850 59090
rect -15650 59020 -15350 59090
rect -15150 59020 -14850 59090
rect -14650 59020 -14350 59090
rect -14150 59020 -13850 59090
rect -13650 59020 -13350 59090
rect -13150 59020 -12850 59090
rect -12650 59020 -12350 59090
rect -12150 59020 -12000 59090
rect -16000 58980 -12000 59020
rect -16000 58910 -15850 58980
rect -15650 58910 -15350 58980
rect -15150 58910 -14850 58980
rect -14650 58910 -14350 58980
rect -14150 58910 -13850 58980
rect -13650 58910 -13350 58980
rect -13150 58910 -12850 58980
rect -12650 58910 -12350 58980
rect -12150 58910 -12000 58980
rect -16000 58900 -12000 58910
rect -16000 58880 -15880 58900
rect -15620 58880 -15380 58900
rect -15120 58880 -14880 58900
rect -14620 58880 -14380 58900
rect -14120 58880 -13880 58900
rect -13620 58880 -13380 58900
rect -13120 58880 -12880 58900
rect -12620 58880 -12380 58900
rect -12120 58880 -12000 58900
rect -16000 58850 -15900 58880
rect -16000 58650 -15980 58850
rect -15910 58650 -15900 58850
rect -16000 58620 -15900 58650
rect -15600 58850 -15400 58880
rect -15600 58650 -15590 58850
rect -15520 58650 -15480 58850
rect -15410 58650 -15400 58850
rect -15600 58620 -15400 58650
rect -15100 58850 -14900 58880
rect -15100 58650 -15090 58850
rect -15020 58650 -14980 58850
rect -14910 58650 -14900 58850
rect -15100 58620 -14900 58650
rect -14600 58850 -14400 58880
rect -14600 58650 -14590 58850
rect -14520 58650 -14480 58850
rect -14410 58650 -14400 58850
rect -14600 58620 -14400 58650
rect -14100 58850 -13900 58880
rect -14100 58650 -14090 58850
rect -14020 58650 -13980 58850
rect -13910 58650 -13900 58850
rect -14100 58620 -13900 58650
rect -13600 58850 -13400 58880
rect -13600 58650 -13590 58850
rect -13520 58650 -13480 58850
rect -13410 58650 -13400 58850
rect -13600 58620 -13400 58650
rect -13100 58850 -12900 58880
rect -13100 58650 -13090 58850
rect -13020 58650 -12980 58850
rect -12910 58650 -12900 58850
rect -13100 58620 -12900 58650
rect -12600 58850 -12400 58880
rect -12600 58650 -12590 58850
rect -12520 58650 -12480 58850
rect -12410 58650 -12400 58850
rect -12600 58620 -12400 58650
rect -12100 58850 -12000 58880
rect -12100 58650 -12090 58850
rect -12020 58650 -12000 58850
rect -12100 58620 -12000 58650
rect -16000 58600 -15880 58620
rect -15620 58600 -15380 58620
rect -15120 58600 -14880 58620
rect -14620 58600 -14380 58620
rect -14120 58600 -13880 58620
rect -13620 58600 -13380 58620
rect -13120 58600 -12880 58620
rect -12620 58600 -12380 58620
rect -12120 58600 -12000 58620
rect -16000 58590 -12000 58600
rect -16000 58520 -15850 58590
rect -15650 58520 -15350 58590
rect -15150 58520 -14850 58590
rect -14650 58520 -14350 58590
rect -14150 58520 -13850 58590
rect -13650 58520 -13350 58590
rect -13150 58520 -12850 58590
rect -12650 58520 -12350 58590
rect -12150 58520 -12000 58590
rect -16000 58480 -12000 58520
rect -16000 58410 -15850 58480
rect -15650 58410 -15350 58480
rect -15150 58410 -14850 58480
rect -14650 58410 -14350 58480
rect -14150 58410 -13850 58480
rect -13650 58410 -13350 58480
rect -13150 58410 -12850 58480
rect -12650 58410 -12350 58480
rect -12150 58410 -12000 58480
rect -16000 58400 -12000 58410
rect -16000 58380 -15880 58400
rect -15620 58380 -15380 58400
rect -15120 58380 -14880 58400
rect -14620 58380 -14380 58400
rect -14120 58380 -13880 58400
rect -13620 58380 -13380 58400
rect -13120 58380 -12880 58400
rect -12620 58380 -12380 58400
rect -12120 58380 -12000 58400
rect -16000 58350 -15900 58380
rect -16000 58150 -15980 58350
rect -15910 58150 -15900 58350
rect -16000 58120 -15900 58150
rect -15600 58350 -15400 58380
rect -15600 58150 -15590 58350
rect -15520 58150 -15480 58350
rect -15410 58150 -15400 58350
rect -15600 58120 -15400 58150
rect -15100 58350 -14900 58380
rect -15100 58150 -15090 58350
rect -15020 58150 -14980 58350
rect -14910 58150 -14900 58350
rect -15100 58120 -14900 58150
rect -14600 58350 -14400 58380
rect -14600 58150 -14590 58350
rect -14520 58150 -14480 58350
rect -14410 58150 -14400 58350
rect -14600 58120 -14400 58150
rect -14100 58350 -13900 58380
rect -14100 58150 -14090 58350
rect -14020 58150 -13980 58350
rect -13910 58150 -13900 58350
rect -14100 58120 -13900 58150
rect -13600 58350 -13400 58380
rect -13600 58150 -13590 58350
rect -13520 58150 -13480 58350
rect -13410 58150 -13400 58350
rect -13600 58120 -13400 58150
rect -13100 58350 -12900 58380
rect -13100 58150 -13090 58350
rect -13020 58150 -12980 58350
rect -12910 58150 -12900 58350
rect -13100 58120 -12900 58150
rect -12600 58350 -12400 58380
rect -12600 58150 -12590 58350
rect -12520 58150 -12480 58350
rect -12410 58150 -12400 58350
rect -12600 58120 -12400 58150
rect -12100 58350 -12000 58380
rect -12100 58150 -12090 58350
rect -12020 58150 -12000 58350
rect -12100 58120 -12000 58150
rect -16000 58100 -15880 58120
rect -15620 58100 -15380 58120
rect -15120 58100 -14880 58120
rect -14620 58100 -14380 58120
rect -14120 58100 -13880 58120
rect -13620 58100 -13380 58120
rect -13120 58100 -12880 58120
rect -12620 58100 -12380 58120
rect -12120 58100 -12000 58120
rect -16000 58090 -12000 58100
rect -16000 58020 -15850 58090
rect -15650 58020 -15350 58090
rect -15150 58020 -14850 58090
rect -14650 58020 -14350 58090
rect -14150 58020 -13850 58090
rect -13650 58020 -13350 58090
rect -13150 58020 -12850 58090
rect -12650 58020 -12350 58090
rect -12150 58020 -12000 58090
rect -16000 57980 -12000 58020
rect -16000 57910 -15850 57980
rect -15650 57910 -15350 57980
rect -15150 57910 -14850 57980
rect -14650 57910 -14350 57980
rect -14150 57910 -13850 57980
rect -13650 57910 -13350 57980
rect -13150 57910 -12850 57980
rect -12650 57910 -12350 57980
rect -12150 57910 -12000 57980
rect -16000 57900 -12000 57910
rect -16000 57880 -15880 57900
rect -15620 57880 -15380 57900
rect -15120 57880 -14880 57900
rect -14620 57880 -14380 57900
rect -14120 57880 -13880 57900
rect -13620 57880 -13380 57900
rect -13120 57880 -12880 57900
rect -12620 57880 -12380 57900
rect -12120 57880 -12000 57900
rect -16000 57850 -15900 57880
rect -16000 57650 -15980 57850
rect -15910 57650 -15900 57850
rect -16000 57620 -15900 57650
rect -15600 57850 -15400 57880
rect -15600 57650 -15590 57850
rect -15520 57650 -15480 57850
rect -15410 57650 -15400 57850
rect -15600 57620 -15400 57650
rect -15100 57850 -14900 57880
rect -15100 57650 -15090 57850
rect -15020 57650 -14980 57850
rect -14910 57650 -14900 57850
rect -15100 57620 -14900 57650
rect -14600 57850 -14400 57880
rect -14600 57650 -14590 57850
rect -14520 57650 -14480 57850
rect -14410 57650 -14400 57850
rect -14600 57620 -14400 57650
rect -14100 57850 -13900 57880
rect -14100 57650 -14090 57850
rect -14020 57650 -13980 57850
rect -13910 57650 -13900 57850
rect -14100 57620 -13900 57650
rect -13600 57850 -13400 57880
rect -13600 57650 -13590 57850
rect -13520 57650 -13480 57850
rect -13410 57650 -13400 57850
rect -13600 57620 -13400 57650
rect -13100 57850 -12900 57880
rect -13100 57650 -13090 57850
rect -13020 57650 -12980 57850
rect -12910 57650 -12900 57850
rect -13100 57620 -12900 57650
rect -12600 57850 -12400 57880
rect -12600 57650 -12590 57850
rect -12520 57650 -12480 57850
rect -12410 57650 -12400 57850
rect -12600 57620 -12400 57650
rect -12100 57850 -12000 57880
rect -12100 57650 -12090 57850
rect -12020 57650 -12000 57850
rect -12100 57620 -12000 57650
rect -16000 57600 -15880 57620
rect -15620 57600 -15380 57620
rect -15120 57600 -14880 57620
rect -14620 57600 -14380 57620
rect -14120 57600 -13880 57620
rect -13620 57600 -13380 57620
rect -13120 57600 -12880 57620
rect -12620 57600 -12380 57620
rect -12120 57600 -12000 57620
rect -16000 57590 -12000 57600
rect -16000 57520 -15850 57590
rect -15650 57520 -15350 57590
rect -15150 57520 -14850 57590
rect -14650 57520 -14350 57590
rect -14150 57520 -13850 57590
rect -13650 57520 -13350 57590
rect -13150 57520 -12850 57590
rect -12650 57520 -12350 57590
rect -12150 57520 -12000 57590
rect -16000 57480 -12000 57520
rect -16000 57410 -15850 57480
rect -15650 57410 -15350 57480
rect -15150 57410 -14850 57480
rect -14650 57410 -14350 57480
rect -14150 57410 -13850 57480
rect -13650 57410 -13350 57480
rect -13150 57410 -12850 57480
rect -12650 57410 -12350 57480
rect -12150 57410 -12000 57480
rect -16000 57400 -12000 57410
rect -16000 57380 -15880 57400
rect -15620 57380 -15380 57400
rect -15120 57380 -14880 57400
rect -14620 57380 -14380 57400
rect -14120 57380 -13880 57400
rect -13620 57380 -13380 57400
rect -13120 57380 -12880 57400
rect -12620 57380 -12380 57400
rect -12120 57380 -12000 57400
rect -16000 57350 -15900 57380
rect -16000 57150 -15980 57350
rect -15910 57150 -15900 57350
rect -16000 57120 -15900 57150
rect -15600 57350 -15400 57380
rect -15600 57150 -15590 57350
rect -15520 57150 -15480 57350
rect -15410 57150 -15400 57350
rect -15600 57120 -15400 57150
rect -15100 57350 -14900 57380
rect -15100 57150 -15090 57350
rect -15020 57150 -14980 57350
rect -14910 57150 -14900 57350
rect -15100 57120 -14900 57150
rect -14600 57350 -14400 57380
rect -14600 57150 -14590 57350
rect -14520 57150 -14480 57350
rect -14410 57150 -14400 57350
rect -14600 57120 -14400 57150
rect -14100 57350 -13900 57380
rect -14100 57150 -14090 57350
rect -14020 57150 -13980 57350
rect -13910 57150 -13900 57350
rect -14100 57120 -13900 57150
rect -13600 57350 -13400 57380
rect -13600 57150 -13590 57350
rect -13520 57150 -13480 57350
rect -13410 57150 -13400 57350
rect -13600 57120 -13400 57150
rect -13100 57350 -12900 57380
rect -13100 57150 -13090 57350
rect -13020 57150 -12980 57350
rect -12910 57150 -12900 57350
rect -13100 57120 -12900 57150
rect -12600 57350 -12400 57380
rect -12600 57150 -12590 57350
rect -12520 57150 -12480 57350
rect -12410 57150 -12400 57350
rect -12600 57120 -12400 57150
rect -12100 57350 -12000 57380
rect -12100 57150 -12090 57350
rect -12020 57150 -12000 57350
rect -12100 57120 -12000 57150
rect -16000 57100 -15880 57120
rect -15620 57100 -15380 57120
rect -15120 57100 -14880 57120
rect -14620 57100 -14380 57120
rect -14120 57100 -13880 57120
rect -13620 57100 -13380 57120
rect -13120 57100 -12880 57120
rect -12620 57100 -12380 57120
rect -12120 57100 -12000 57120
rect -16000 57090 -12000 57100
rect -16000 57020 -15850 57090
rect -15650 57020 -15350 57090
rect -15150 57020 -14850 57090
rect -14650 57020 -14350 57090
rect -14150 57020 -13850 57090
rect -13650 57020 -13350 57090
rect -13150 57020 -12850 57090
rect -12650 57020 -12350 57090
rect -12150 57020 -12000 57090
rect -16000 56980 -12000 57020
rect -16000 56910 -15850 56980
rect -15650 56910 -15350 56980
rect -15150 56910 -14850 56980
rect -14650 56910 -14350 56980
rect -14150 56910 -13850 56980
rect -13650 56910 -13350 56980
rect -13150 56910 -12850 56980
rect -12650 56910 -12350 56980
rect -12150 56910 -12000 56980
rect -16000 56900 -12000 56910
rect -16000 56880 -15880 56900
rect -15620 56880 -15380 56900
rect -15120 56880 -14880 56900
rect -14620 56880 -14380 56900
rect -14120 56880 -13880 56900
rect -13620 56880 -13380 56900
rect -13120 56880 -12880 56900
rect -12620 56880 -12380 56900
rect -12120 56880 -12000 56900
rect -16000 56850 -15900 56880
rect -16000 56650 -15980 56850
rect -15910 56650 -15900 56850
rect -16000 56620 -15900 56650
rect -15600 56850 -15400 56880
rect -15600 56650 -15590 56850
rect -15520 56650 -15480 56850
rect -15410 56650 -15400 56850
rect -15600 56620 -15400 56650
rect -15100 56850 -14900 56880
rect -15100 56650 -15090 56850
rect -15020 56650 -14980 56850
rect -14910 56650 -14900 56850
rect -15100 56620 -14900 56650
rect -14600 56850 -14400 56880
rect -14600 56650 -14590 56850
rect -14520 56650 -14480 56850
rect -14410 56650 -14400 56850
rect -14600 56620 -14400 56650
rect -14100 56850 -13900 56880
rect -14100 56650 -14090 56850
rect -14020 56650 -13980 56850
rect -13910 56650 -13900 56850
rect -14100 56620 -13900 56650
rect -13600 56850 -13400 56880
rect -13600 56650 -13590 56850
rect -13520 56650 -13480 56850
rect -13410 56650 -13400 56850
rect -13600 56620 -13400 56650
rect -13100 56850 -12900 56880
rect -13100 56650 -13090 56850
rect -13020 56650 -12980 56850
rect -12910 56650 -12900 56850
rect -13100 56620 -12900 56650
rect -12600 56850 -12400 56880
rect -12600 56650 -12590 56850
rect -12520 56650 -12480 56850
rect -12410 56650 -12400 56850
rect -12600 56620 -12400 56650
rect -12100 56850 -12000 56880
rect -12100 56650 -12090 56850
rect -12020 56650 -12000 56850
rect -12100 56620 -12000 56650
rect -16000 56600 -15880 56620
rect -15620 56600 -15380 56620
rect -15120 56600 -14880 56620
rect -14620 56600 -14380 56620
rect -14120 56600 -13880 56620
rect -13620 56600 -13380 56620
rect -13120 56600 -12880 56620
rect -12620 56600 -12380 56620
rect -12120 56600 -12000 56620
rect -16000 56590 -12000 56600
rect -16000 56520 -15850 56590
rect -15650 56520 -15350 56590
rect -15150 56520 -14850 56590
rect -14650 56520 -14350 56590
rect -14150 56520 -13850 56590
rect -13650 56520 -13350 56590
rect -13150 56520 -12850 56590
rect -12650 56520 -12350 56590
rect -12150 56520 -12000 56590
rect -16000 56480 -12000 56520
rect -16000 56410 -15850 56480
rect -15650 56410 -15350 56480
rect -15150 56410 -14850 56480
rect -14650 56410 -14350 56480
rect -14150 56410 -13850 56480
rect -13650 56410 -13350 56480
rect -13150 56410 -12850 56480
rect -12650 56410 -12350 56480
rect -12150 56410 -12000 56480
rect -16000 56400 -12000 56410
rect -16000 56380 -15880 56400
rect -15620 56380 -15380 56400
rect -15120 56380 -14880 56400
rect -14620 56380 -14380 56400
rect -14120 56380 -13880 56400
rect -13620 56380 -13380 56400
rect -13120 56380 -12880 56400
rect -12620 56380 -12380 56400
rect -12120 56380 -12000 56400
rect -16000 56350 -15900 56380
rect -16000 56150 -15980 56350
rect -15910 56150 -15900 56350
rect -16000 56120 -15900 56150
rect -15600 56350 -15400 56380
rect -15600 56150 -15590 56350
rect -15520 56150 -15480 56350
rect -15410 56150 -15400 56350
rect -15600 56120 -15400 56150
rect -15100 56350 -14900 56380
rect -15100 56150 -15090 56350
rect -15020 56150 -14980 56350
rect -14910 56150 -14900 56350
rect -15100 56120 -14900 56150
rect -14600 56350 -14400 56380
rect -14600 56150 -14590 56350
rect -14520 56150 -14480 56350
rect -14410 56150 -14400 56350
rect -14600 56120 -14400 56150
rect -14100 56350 -13900 56380
rect -14100 56150 -14090 56350
rect -14020 56150 -13980 56350
rect -13910 56150 -13900 56350
rect -14100 56120 -13900 56150
rect -13600 56350 -13400 56380
rect -13600 56150 -13590 56350
rect -13520 56150 -13480 56350
rect -13410 56150 -13400 56350
rect -13600 56120 -13400 56150
rect -13100 56350 -12900 56380
rect -13100 56150 -13090 56350
rect -13020 56150 -12980 56350
rect -12910 56150 -12900 56350
rect -13100 56120 -12900 56150
rect -12600 56350 -12400 56380
rect -12600 56150 -12590 56350
rect -12520 56150 -12480 56350
rect -12410 56150 -12400 56350
rect -12600 56120 -12400 56150
rect -12100 56350 -12000 56380
rect -12100 56150 -12090 56350
rect -12020 56150 -12000 56350
rect -12100 56120 -12000 56150
rect -16000 56100 -15880 56120
rect -15620 56100 -15380 56120
rect -15120 56100 -14880 56120
rect -14620 56100 -14380 56120
rect -14120 56100 -13880 56120
rect -13620 56100 -13380 56120
rect -13120 56100 -12880 56120
rect -12620 56100 -12380 56120
rect -12120 56100 -12000 56120
rect -16000 56090 -12000 56100
rect -16000 56020 -15850 56090
rect -15650 56020 -15350 56090
rect -15150 56020 -14850 56090
rect -14650 56020 -14350 56090
rect -14150 56020 -13850 56090
rect -13650 56020 -13350 56090
rect -13150 56020 -12850 56090
rect -12650 56020 -12350 56090
rect -12150 56020 -12000 56090
rect -16000 55980 -12000 56020
rect -16000 55910 -15850 55980
rect -15650 55910 -15350 55980
rect -15150 55910 -14850 55980
rect -14650 55910 -14350 55980
rect -14150 55910 -13850 55980
rect -13650 55910 -13350 55980
rect -13150 55910 -12850 55980
rect -12650 55910 -12350 55980
rect -12150 55910 -12000 55980
rect -16000 55900 -12000 55910
rect -16000 55880 -15880 55900
rect -15620 55880 -15380 55900
rect -15120 55880 -14880 55900
rect -14620 55880 -14380 55900
rect -14120 55880 -13880 55900
rect -13620 55880 -13380 55900
rect -13120 55880 -12880 55900
rect -12620 55880 -12380 55900
rect -12120 55880 -12000 55900
rect -16000 55850 -15900 55880
rect -16000 55650 -15980 55850
rect -15910 55650 -15900 55850
rect -16000 55620 -15900 55650
rect -15600 55850 -15400 55880
rect -15600 55650 -15590 55850
rect -15520 55650 -15480 55850
rect -15410 55650 -15400 55850
rect -15600 55620 -15400 55650
rect -15100 55850 -14900 55880
rect -15100 55650 -15090 55850
rect -15020 55650 -14980 55850
rect -14910 55650 -14900 55850
rect -15100 55620 -14900 55650
rect -14600 55850 -14400 55880
rect -14600 55650 -14590 55850
rect -14520 55650 -14480 55850
rect -14410 55650 -14400 55850
rect -14600 55620 -14400 55650
rect -14100 55850 -13900 55880
rect -14100 55650 -14090 55850
rect -14020 55650 -13980 55850
rect -13910 55650 -13900 55850
rect -14100 55620 -13900 55650
rect -13600 55850 -13400 55880
rect -13600 55650 -13590 55850
rect -13520 55650 -13480 55850
rect -13410 55650 -13400 55850
rect -13600 55620 -13400 55650
rect -13100 55850 -12900 55880
rect -13100 55650 -13090 55850
rect -13020 55650 -12980 55850
rect -12910 55650 -12900 55850
rect -13100 55620 -12900 55650
rect -12600 55850 -12400 55880
rect -12600 55650 -12590 55850
rect -12520 55650 -12480 55850
rect -12410 55650 -12400 55850
rect -12600 55620 -12400 55650
rect -12100 55850 -12000 55880
rect -12100 55650 -12090 55850
rect -12020 55650 -12000 55850
rect -12100 55620 -12000 55650
rect -16000 55600 -15880 55620
rect -15620 55600 -15380 55620
rect -15120 55600 -14880 55620
rect -14620 55600 -14380 55620
rect -14120 55600 -13880 55620
rect -13620 55600 -13380 55620
rect -13120 55600 -12880 55620
rect -12620 55600 -12380 55620
rect -12120 55600 -12000 55620
rect -16000 55590 -12000 55600
rect -16000 55520 -15850 55590
rect -15650 55520 -15350 55590
rect -15150 55520 -14850 55590
rect -14650 55520 -14350 55590
rect -14150 55520 -13850 55590
rect -13650 55520 -13350 55590
rect -13150 55520 -12850 55590
rect -12650 55520 -12350 55590
rect -12150 55520 -12000 55590
rect -16000 55480 -12000 55520
rect -16000 55410 -15850 55480
rect -15650 55410 -15350 55480
rect -15150 55410 -14850 55480
rect -14650 55410 -14350 55480
rect -14150 55410 -13850 55480
rect -13650 55410 -13350 55480
rect -13150 55410 -12850 55480
rect -12650 55410 -12350 55480
rect -12150 55410 -12000 55480
rect -16000 55400 -12000 55410
rect -16000 55380 -15880 55400
rect -15620 55380 -15380 55400
rect -15120 55380 -14880 55400
rect -14620 55380 -14380 55400
rect -14120 55380 -13880 55400
rect -13620 55380 -13380 55400
rect -13120 55380 -12880 55400
rect -12620 55380 -12380 55400
rect -12120 55380 -12000 55400
rect -16000 55350 -15900 55380
rect -16000 55150 -15980 55350
rect -15910 55150 -15900 55350
rect -16000 55120 -15900 55150
rect -15600 55350 -15400 55380
rect -15600 55150 -15590 55350
rect -15520 55150 -15480 55350
rect -15410 55150 -15400 55350
rect -15600 55120 -15400 55150
rect -15100 55350 -14900 55380
rect -15100 55150 -15090 55350
rect -15020 55150 -14980 55350
rect -14910 55150 -14900 55350
rect -15100 55120 -14900 55150
rect -14600 55350 -14400 55380
rect -14600 55150 -14590 55350
rect -14520 55150 -14480 55350
rect -14410 55150 -14400 55350
rect -14600 55120 -14400 55150
rect -14100 55350 -13900 55380
rect -14100 55150 -14090 55350
rect -14020 55150 -13980 55350
rect -13910 55150 -13900 55350
rect -14100 55120 -13900 55150
rect -13600 55350 -13400 55380
rect -13600 55150 -13590 55350
rect -13520 55150 -13480 55350
rect -13410 55150 -13400 55350
rect -13600 55120 -13400 55150
rect -13100 55350 -12900 55380
rect -13100 55150 -13090 55350
rect -13020 55150 -12980 55350
rect -12910 55150 -12900 55350
rect -13100 55120 -12900 55150
rect -12600 55350 -12400 55380
rect -12600 55150 -12590 55350
rect -12520 55150 -12480 55350
rect -12410 55150 -12400 55350
rect -12600 55120 -12400 55150
rect -12100 55350 -12000 55380
rect -12100 55150 -12090 55350
rect -12020 55150 -12000 55350
rect -12100 55120 -12000 55150
rect -16000 55100 -15880 55120
rect -15620 55100 -15380 55120
rect -15120 55100 -14880 55120
rect -14620 55100 -14380 55120
rect -14120 55100 -13880 55120
rect -13620 55100 -13380 55120
rect -13120 55100 -12880 55120
rect -12620 55100 -12380 55120
rect -12120 55100 -12000 55120
rect -16000 55090 -12000 55100
rect -16000 55020 -15850 55090
rect -15650 55020 -15350 55090
rect -15150 55020 -14850 55090
rect -14650 55020 -14350 55090
rect -14150 55020 -13850 55090
rect -13650 55020 -13350 55090
rect -13150 55020 -12850 55090
rect -12650 55020 -12350 55090
rect -12150 55020 -12000 55090
rect -16000 54980 -12000 55020
rect -16000 54910 -15850 54980
rect -15650 54910 -15350 54980
rect -15150 54910 -14850 54980
rect -14650 54910 -14350 54980
rect -14150 54910 -13850 54980
rect -13650 54910 -13350 54980
rect -13150 54910 -12850 54980
rect -12650 54910 -12350 54980
rect -12150 54910 -12000 54980
rect -16000 54900 -12000 54910
rect -16000 54880 -15880 54900
rect -15620 54880 -15380 54900
rect -15120 54880 -14880 54900
rect -14620 54880 -14380 54900
rect -14120 54880 -13880 54900
rect -13620 54880 -13380 54900
rect -13120 54880 -12880 54900
rect -12620 54880 -12380 54900
rect -12120 54880 -12000 54900
rect -16000 54850 -15900 54880
rect -16000 54650 -15980 54850
rect -15910 54650 -15900 54850
rect -16000 54620 -15900 54650
rect -15600 54850 -15400 54880
rect -15600 54650 -15590 54850
rect -15520 54650 -15480 54850
rect -15410 54650 -15400 54850
rect -15600 54620 -15400 54650
rect -15100 54850 -14900 54880
rect -15100 54650 -15090 54850
rect -15020 54650 -14980 54850
rect -14910 54650 -14900 54850
rect -15100 54620 -14900 54650
rect -14600 54850 -14400 54880
rect -14600 54650 -14590 54850
rect -14520 54650 -14480 54850
rect -14410 54650 -14400 54850
rect -14600 54620 -14400 54650
rect -14100 54850 -13900 54880
rect -14100 54650 -14090 54850
rect -14020 54650 -13980 54850
rect -13910 54650 -13900 54850
rect -14100 54620 -13900 54650
rect -13600 54850 -13400 54880
rect -13600 54650 -13590 54850
rect -13520 54650 -13480 54850
rect -13410 54650 -13400 54850
rect -13600 54620 -13400 54650
rect -13100 54850 -12900 54880
rect -13100 54650 -13090 54850
rect -13020 54650 -12980 54850
rect -12910 54650 -12900 54850
rect -13100 54620 -12900 54650
rect -12600 54850 -12400 54880
rect -12600 54650 -12590 54850
rect -12520 54650 -12480 54850
rect -12410 54650 -12400 54850
rect -12600 54620 -12400 54650
rect -12100 54850 -12000 54880
rect -12100 54650 -12090 54850
rect -12020 54650 -12000 54850
rect -12100 54620 -12000 54650
rect -16000 54600 -15880 54620
rect -15620 54600 -15380 54620
rect -15120 54600 -14880 54620
rect -14620 54600 -14380 54620
rect -14120 54600 -13880 54620
rect -13620 54600 -13380 54620
rect -13120 54600 -12880 54620
rect -12620 54600 -12380 54620
rect -12120 54600 -12000 54620
rect -16000 54590 -12000 54600
rect -16000 54520 -15850 54590
rect -15650 54520 -15350 54590
rect -15150 54520 -14850 54590
rect -14650 54520 -14350 54590
rect -14150 54520 -13850 54590
rect -13650 54520 -13350 54590
rect -13150 54520 -12850 54590
rect -12650 54520 -12350 54590
rect -12150 54520 -12000 54590
rect -16000 54480 -12000 54520
rect -16000 54410 -15850 54480
rect -15650 54410 -15350 54480
rect -15150 54410 -14850 54480
rect -14650 54410 -14350 54480
rect -14150 54410 -13850 54480
rect -13650 54410 -13350 54480
rect -13150 54410 -12850 54480
rect -12650 54410 -12350 54480
rect -12150 54410 -12000 54480
rect -16000 54400 -12000 54410
rect -16000 54380 -15880 54400
rect -15620 54380 -15380 54400
rect -15120 54380 -14880 54400
rect -14620 54380 -14380 54400
rect -14120 54380 -13880 54400
rect -13620 54380 -13380 54400
rect -13120 54380 -12880 54400
rect -12620 54380 -12380 54400
rect -12120 54380 -12000 54400
rect -16000 54350 -15900 54380
rect -16000 54150 -15980 54350
rect -15910 54150 -15900 54350
rect -16000 54120 -15900 54150
rect -15600 54350 -15400 54380
rect -15600 54150 -15590 54350
rect -15520 54150 -15480 54350
rect -15410 54150 -15400 54350
rect -15600 54120 -15400 54150
rect -15100 54350 -14900 54380
rect -15100 54150 -15090 54350
rect -15020 54150 -14980 54350
rect -14910 54150 -14900 54350
rect -15100 54120 -14900 54150
rect -14600 54350 -14400 54380
rect -14600 54150 -14590 54350
rect -14520 54150 -14480 54350
rect -14410 54150 -14400 54350
rect -14600 54120 -14400 54150
rect -14100 54350 -13900 54380
rect -14100 54150 -14090 54350
rect -14020 54150 -13980 54350
rect -13910 54150 -13900 54350
rect -14100 54120 -13900 54150
rect -13600 54350 -13400 54380
rect -13600 54150 -13590 54350
rect -13520 54150 -13480 54350
rect -13410 54150 -13400 54350
rect -13600 54120 -13400 54150
rect -13100 54350 -12900 54380
rect -13100 54150 -13090 54350
rect -13020 54150 -12980 54350
rect -12910 54150 -12900 54350
rect -13100 54120 -12900 54150
rect -12600 54350 -12400 54380
rect -12600 54150 -12590 54350
rect -12520 54150 -12480 54350
rect -12410 54150 -12400 54350
rect -12600 54120 -12400 54150
rect -12100 54350 -12000 54380
rect -12100 54150 -12090 54350
rect -12020 54150 -12000 54350
rect -12100 54120 -12000 54150
rect -16000 54100 -15880 54120
rect -15620 54100 -15380 54120
rect -15120 54100 -14880 54120
rect -14620 54100 -14380 54120
rect -14120 54100 -13880 54120
rect -13620 54100 -13380 54120
rect -13120 54100 -12880 54120
rect -12620 54100 -12380 54120
rect -12120 54100 -12000 54120
rect -16000 54090 -12000 54100
rect -16000 54020 -15850 54090
rect -15650 54020 -15350 54090
rect -15150 54020 -14850 54090
rect -14650 54020 -14350 54090
rect -14150 54020 -13850 54090
rect -13650 54020 -13350 54090
rect -13150 54020 -12850 54090
rect -12650 54020 -12350 54090
rect -12150 54020 -12000 54090
rect -16000 53980 -12000 54020
rect -16000 53910 -15850 53980
rect -15650 53910 -15350 53980
rect -15150 53910 -14850 53980
rect -14650 53910 -14350 53980
rect -14150 53910 -13850 53980
rect -13650 53910 -13350 53980
rect -13150 53910 -12850 53980
rect -12650 53910 -12350 53980
rect -12150 53910 -12000 53980
rect -16000 53900 -12000 53910
rect -16000 53880 -15880 53900
rect -15620 53880 -15380 53900
rect -15120 53880 -14880 53900
rect -14620 53880 -14380 53900
rect -14120 53880 -13880 53900
rect -13620 53880 -13380 53900
rect -13120 53880 -12880 53900
rect -12620 53880 -12380 53900
rect -12120 53880 -12000 53900
rect -16000 53850 -15900 53880
rect -16000 53650 -15980 53850
rect -15910 53650 -15900 53850
rect -16000 53620 -15900 53650
rect -15600 53850 -15400 53880
rect -15600 53650 -15590 53850
rect -15520 53650 -15480 53850
rect -15410 53650 -15400 53850
rect -15600 53620 -15400 53650
rect -15100 53850 -14900 53880
rect -15100 53650 -15090 53850
rect -15020 53650 -14980 53850
rect -14910 53650 -14900 53850
rect -15100 53620 -14900 53650
rect -14600 53850 -14400 53880
rect -14600 53650 -14590 53850
rect -14520 53650 -14480 53850
rect -14410 53650 -14400 53850
rect -14600 53620 -14400 53650
rect -14100 53850 -13900 53880
rect -14100 53650 -14090 53850
rect -14020 53650 -13980 53850
rect -13910 53650 -13900 53850
rect -14100 53620 -13900 53650
rect -13600 53850 -13400 53880
rect -13600 53650 -13590 53850
rect -13520 53650 -13480 53850
rect -13410 53650 -13400 53850
rect -13600 53620 -13400 53650
rect -13100 53850 -12900 53880
rect -13100 53650 -13090 53850
rect -13020 53650 -12980 53850
rect -12910 53650 -12900 53850
rect -13100 53620 -12900 53650
rect -12600 53850 -12400 53880
rect -12600 53650 -12590 53850
rect -12520 53650 -12480 53850
rect -12410 53650 -12400 53850
rect -12600 53620 -12400 53650
rect -12100 53850 -12000 53880
rect -12100 53650 -12090 53850
rect -12020 53650 -12000 53850
rect -12100 53620 -12000 53650
rect -16000 53600 -15880 53620
rect -15620 53600 -15380 53620
rect -15120 53600 -14880 53620
rect -14620 53600 -14380 53620
rect -14120 53600 -13880 53620
rect -13620 53600 -13380 53620
rect -13120 53600 -12880 53620
rect -12620 53600 -12380 53620
rect -12120 53600 -12000 53620
rect -16000 53590 -12000 53600
rect -16000 53520 -15850 53590
rect -15650 53520 -15350 53590
rect -15150 53520 -14850 53590
rect -14650 53520 -14350 53590
rect -14150 53520 -13850 53590
rect -13650 53520 -13350 53590
rect -13150 53520 -12850 53590
rect -12650 53520 -12350 53590
rect -12150 53520 -12000 53590
rect -16000 53480 -12000 53520
rect -16000 53410 -15850 53480
rect -15650 53410 -15350 53480
rect -15150 53410 -14850 53480
rect -14650 53410 -14350 53480
rect -14150 53410 -13850 53480
rect -13650 53410 -13350 53480
rect -13150 53410 -12850 53480
rect -12650 53410 -12350 53480
rect -12150 53410 -12000 53480
rect -16000 53400 -12000 53410
rect -16000 53380 -15880 53400
rect -15620 53380 -15380 53400
rect -15120 53380 -14880 53400
rect -14620 53380 -14380 53400
rect -14120 53380 -13880 53400
rect -13620 53380 -13380 53400
rect -13120 53380 -12880 53400
rect -12620 53380 -12380 53400
rect -12120 53380 -12000 53400
rect -16000 53350 -15900 53380
rect -16000 53150 -15980 53350
rect -15910 53150 -15900 53350
rect -16000 53120 -15900 53150
rect -15600 53350 -15400 53380
rect -15600 53150 -15590 53350
rect -15520 53150 -15480 53350
rect -15410 53150 -15400 53350
rect -15600 53120 -15400 53150
rect -15100 53350 -14900 53380
rect -15100 53150 -15090 53350
rect -15020 53150 -14980 53350
rect -14910 53150 -14900 53350
rect -15100 53120 -14900 53150
rect -14600 53350 -14400 53380
rect -14600 53150 -14590 53350
rect -14520 53150 -14480 53350
rect -14410 53150 -14400 53350
rect -14600 53120 -14400 53150
rect -14100 53350 -13900 53380
rect -14100 53150 -14090 53350
rect -14020 53150 -13980 53350
rect -13910 53150 -13900 53350
rect -14100 53120 -13900 53150
rect -13600 53350 -13400 53380
rect -13600 53150 -13590 53350
rect -13520 53150 -13480 53350
rect -13410 53150 -13400 53350
rect -13600 53120 -13400 53150
rect -13100 53350 -12900 53380
rect -13100 53150 -13090 53350
rect -13020 53150 -12980 53350
rect -12910 53150 -12900 53350
rect -13100 53120 -12900 53150
rect -12600 53350 -12400 53380
rect -12600 53150 -12590 53350
rect -12520 53150 -12480 53350
rect -12410 53150 -12400 53350
rect -12600 53120 -12400 53150
rect -12100 53350 -12000 53380
rect -12100 53150 -12090 53350
rect -12020 53150 -12000 53350
rect -12100 53120 -12000 53150
rect -16000 53100 -15880 53120
rect -15620 53100 -15380 53120
rect -15120 53100 -14880 53120
rect -14620 53100 -14380 53120
rect -14120 53100 -13880 53120
rect -13620 53100 -13380 53120
rect -13120 53100 -12880 53120
rect -12620 53100 -12380 53120
rect -12120 53100 -12000 53120
rect -16000 53090 -12000 53100
rect -16000 53020 -15850 53090
rect -15650 53020 -15350 53090
rect -15150 53020 -14850 53090
rect -14650 53020 -14350 53090
rect -14150 53020 -13850 53090
rect -13650 53020 -13350 53090
rect -13150 53020 -12850 53090
rect -12650 53020 -12350 53090
rect -12150 53020 -12000 53090
rect -16000 52980 -12000 53020
rect -16000 52910 -15850 52980
rect -15650 52910 -15350 52980
rect -15150 52910 -14850 52980
rect -14650 52910 -14350 52980
rect -14150 52910 -13850 52980
rect -13650 52910 -13350 52980
rect -13150 52910 -12850 52980
rect -12650 52910 -12350 52980
rect -12150 52910 -12000 52980
rect -16000 52900 -12000 52910
rect -16000 52880 -15880 52900
rect -15620 52880 -15380 52900
rect -15120 52880 -14880 52900
rect -14620 52880 -14380 52900
rect -14120 52880 -13880 52900
rect -13620 52880 -13380 52900
rect -13120 52880 -12880 52900
rect -12620 52880 -12380 52900
rect -12120 52880 -12000 52900
rect -16000 52850 -15900 52880
rect -16000 52650 -15980 52850
rect -15910 52650 -15900 52850
rect -16000 52620 -15900 52650
rect -15600 52850 -15400 52880
rect -15600 52650 -15590 52850
rect -15520 52650 -15480 52850
rect -15410 52650 -15400 52850
rect -15600 52620 -15400 52650
rect -15100 52850 -14900 52880
rect -15100 52650 -15090 52850
rect -15020 52650 -14980 52850
rect -14910 52650 -14900 52850
rect -15100 52620 -14900 52650
rect -14600 52850 -14400 52880
rect -14600 52650 -14590 52850
rect -14520 52650 -14480 52850
rect -14410 52650 -14400 52850
rect -14600 52620 -14400 52650
rect -14100 52850 -13900 52880
rect -14100 52650 -14090 52850
rect -14020 52650 -13980 52850
rect -13910 52650 -13900 52850
rect -14100 52620 -13900 52650
rect -13600 52850 -13400 52880
rect -13600 52650 -13590 52850
rect -13520 52650 -13480 52850
rect -13410 52650 -13400 52850
rect -13600 52620 -13400 52650
rect -13100 52850 -12900 52880
rect -13100 52650 -13090 52850
rect -13020 52650 -12980 52850
rect -12910 52650 -12900 52850
rect -13100 52620 -12900 52650
rect -12600 52850 -12400 52880
rect -12600 52650 -12590 52850
rect -12520 52650 -12480 52850
rect -12410 52650 -12400 52850
rect -12600 52620 -12400 52650
rect -12100 52850 -12000 52880
rect -12100 52650 -12090 52850
rect -12020 52650 -12000 52850
rect -12100 52620 -12000 52650
rect -16000 52600 -15880 52620
rect -15620 52600 -15380 52620
rect -15120 52600 -14880 52620
rect -14620 52600 -14380 52620
rect -14120 52600 -13880 52620
rect -13620 52600 -13380 52620
rect -13120 52600 -12880 52620
rect -12620 52600 -12380 52620
rect -12120 52600 -12000 52620
rect -16000 52590 -12000 52600
rect -16000 52520 -15850 52590
rect -15650 52520 -15350 52590
rect -15150 52520 -14850 52590
rect -14650 52520 -14350 52590
rect -14150 52520 -13850 52590
rect -13650 52520 -13350 52590
rect -13150 52520 -12850 52590
rect -12650 52520 -12350 52590
rect -12150 52520 -12000 52590
rect -16000 52480 -12000 52520
rect -16000 52410 -15850 52480
rect -15650 52410 -15350 52480
rect -15150 52410 -14850 52480
rect -14650 52410 -14350 52480
rect -14150 52410 -13850 52480
rect -13650 52410 -13350 52480
rect -13150 52410 -12850 52480
rect -12650 52410 -12350 52480
rect -12150 52410 -12000 52480
rect -16000 52400 -12000 52410
rect -16000 52380 -15880 52400
rect -15620 52380 -15380 52400
rect -15120 52380 -14880 52400
rect -14620 52380 -14380 52400
rect -14120 52380 -13880 52400
rect -13620 52380 -13380 52400
rect -13120 52380 -12880 52400
rect -12620 52380 -12380 52400
rect -12120 52380 -12000 52400
rect -16000 52350 -15900 52380
rect -16000 52150 -15980 52350
rect -15910 52150 -15900 52350
rect -16000 52120 -15900 52150
rect -15600 52350 -15400 52380
rect -15600 52150 -15590 52350
rect -15520 52150 -15480 52350
rect -15410 52150 -15400 52350
rect -15600 52120 -15400 52150
rect -15100 52350 -14900 52380
rect -15100 52150 -15090 52350
rect -15020 52150 -14980 52350
rect -14910 52150 -14900 52350
rect -15100 52120 -14900 52150
rect -14600 52350 -14400 52380
rect -14600 52150 -14590 52350
rect -14520 52150 -14480 52350
rect -14410 52150 -14400 52350
rect -14600 52120 -14400 52150
rect -14100 52350 -13900 52380
rect -14100 52150 -14090 52350
rect -14020 52150 -13980 52350
rect -13910 52150 -13900 52350
rect -14100 52120 -13900 52150
rect -13600 52350 -13400 52380
rect -13600 52150 -13590 52350
rect -13520 52150 -13480 52350
rect -13410 52150 -13400 52350
rect -13600 52120 -13400 52150
rect -13100 52350 -12900 52380
rect -13100 52150 -13090 52350
rect -13020 52150 -12980 52350
rect -12910 52150 -12900 52350
rect -13100 52120 -12900 52150
rect -12600 52350 -12400 52380
rect -12600 52150 -12590 52350
rect -12520 52150 -12480 52350
rect -12410 52150 -12400 52350
rect -12600 52120 -12400 52150
rect -12100 52350 -12000 52380
rect -12100 52150 -12090 52350
rect -12020 52150 -12000 52350
rect -12100 52120 -12000 52150
rect -16000 52100 -15880 52120
rect -15620 52100 -15380 52120
rect -15120 52100 -14880 52120
rect -14620 52100 -14380 52120
rect -14120 52100 -13880 52120
rect -13620 52100 -13380 52120
rect -13120 52100 -12880 52120
rect -12620 52100 -12380 52120
rect -12120 52100 -12000 52120
rect -16000 52090 -12000 52100
rect -16000 52020 -15850 52090
rect -15650 52020 -15350 52090
rect -15150 52020 -14850 52090
rect -14650 52020 -14350 52090
rect -14150 52020 -13850 52090
rect -13650 52020 -13350 52090
rect -13150 52020 -12850 52090
rect -12650 52020 -12350 52090
rect -12150 52020 -12000 52090
rect -16000 51980 -12000 52020
rect -16000 51910 -15850 51980
rect -15650 51910 -15350 51980
rect -15150 51910 -14850 51980
rect -14650 51910 -14350 51980
rect -14150 51910 -13850 51980
rect -13650 51910 -13350 51980
rect -13150 51910 -12850 51980
rect -12650 51910 -12350 51980
rect -12150 51910 -12000 51980
rect -16000 51900 -12000 51910
rect -16000 51880 -15880 51900
rect -15620 51880 -15380 51900
rect -15120 51880 -14880 51900
rect -14620 51880 -14380 51900
rect -14120 51880 -13880 51900
rect -13620 51880 -13380 51900
rect -13120 51880 -12880 51900
rect -12620 51880 -12380 51900
rect -12120 51880 -12000 51900
rect -16000 51850 -15900 51880
rect -16000 51650 -15980 51850
rect -15910 51650 -15900 51850
rect -16000 51620 -15900 51650
rect -15600 51850 -15400 51880
rect -15600 51650 -15590 51850
rect -15520 51650 -15480 51850
rect -15410 51650 -15400 51850
rect -15600 51620 -15400 51650
rect -15100 51850 -14900 51880
rect -15100 51650 -15090 51850
rect -15020 51650 -14980 51850
rect -14910 51650 -14900 51850
rect -15100 51620 -14900 51650
rect -14600 51850 -14400 51880
rect -14600 51650 -14590 51850
rect -14520 51650 -14480 51850
rect -14410 51650 -14400 51850
rect -14600 51620 -14400 51650
rect -14100 51850 -13900 51880
rect -14100 51650 -14090 51850
rect -14020 51650 -13980 51850
rect -13910 51650 -13900 51850
rect -14100 51620 -13900 51650
rect -13600 51850 -13400 51880
rect -13600 51650 -13590 51850
rect -13520 51650 -13480 51850
rect -13410 51650 -13400 51850
rect -13600 51620 -13400 51650
rect -13100 51850 -12900 51880
rect -13100 51650 -13090 51850
rect -13020 51650 -12980 51850
rect -12910 51650 -12900 51850
rect -13100 51620 -12900 51650
rect -12600 51850 -12400 51880
rect -12600 51650 -12590 51850
rect -12520 51650 -12480 51850
rect -12410 51650 -12400 51850
rect -12600 51620 -12400 51650
rect -12100 51850 -12000 51880
rect -12100 51650 -12090 51850
rect -12020 51650 -12000 51850
rect -12100 51620 -12000 51650
rect -16000 51600 -15880 51620
rect -15620 51600 -15380 51620
rect -15120 51600 -14880 51620
rect -14620 51600 -14380 51620
rect -14120 51600 -13880 51620
rect -13620 51600 -13380 51620
rect -13120 51600 -12880 51620
rect -12620 51600 -12380 51620
rect -12120 51600 -12000 51620
rect -16000 51590 -12000 51600
rect -16000 51520 -15850 51590
rect -15650 51520 -15350 51590
rect -15150 51520 -14850 51590
rect -14650 51520 -14350 51590
rect -14150 51520 -13850 51590
rect -13650 51520 -13350 51590
rect -13150 51520 -12850 51590
rect -12650 51520 -12350 51590
rect -12150 51520 -12000 51590
rect -16000 51480 -12000 51520
rect -16000 51410 -15850 51480
rect -15650 51410 -15350 51480
rect -15150 51410 -14850 51480
rect -14650 51410 -14350 51480
rect -14150 51410 -13850 51480
rect -13650 51410 -13350 51480
rect -13150 51410 -12850 51480
rect -12650 51410 -12350 51480
rect -12150 51410 -12000 51480
rect -16000 51400 -12000 51410
rect -16000 51380 -15880 51400
rect -15620 51380 -15380 51400
rect -15120 51380 -14880 51400
rect -14620 51380 -14380 51400
rect -14120 51380 -13880 51400
rect -13620 51380 -13380 51400
rect -13120 51380 -12880 51400
rect -12620 51380 -12380 51400
rect -12120 51380 -12000 51400
rect -16000 51350 -15900 51380
rect -16000 51150 -15980 51350
rect -15910 51150 -15900 51350
rect -16000 51120 -15900 51150
rect -15600 51350 -15400 51380
rect -15600 51150 -15590 51350
rect -15520 51150 -15480 51350
rect -15410 51150 -15400 51350
rect -15600 51120 -15400 51150
rect -15100 51350 -14900 51380
rect -15100 51150 -15090 51350
rect -15020 51150 -14980 51350
rect -14910 51150 -14900 51350
rect -15100 51120 -14900 51150
rect -14600 51350 -14400 51380
rect -14600 51150 -14590 51350
rect -14520 51150 -14480 51350
rect -14410 51150 -14400 51350
rect -14600 51120 -14400 51150
rect -14100 51350 -13900 51380
rect -14100 51150 -14090 51350
rect -14020 51150 -13980 51350
rect -13910 51150 -13900 51350
rect -14100 51120 -13900 51150
rect -13600 51350 -13400 51380
rect -13600 51150 -13590 51350
rect -13520 51150 -13480 51350
rect -13410 51150 -13400 51350
rect -13600 51120 -13400 51150
rect -13100 51350 -12900 51380
rect -13100 51150 -13090 51350
rect -13020 51150 -12980 51350
rect -12910 51150 -12900 51350
rect -13100 51120 -12900 51150
rect -12600 51350 -12400 51380
rect -12600 51150 -12590 51350
rect -12520 51150 -12480 51350
rect -12410 51150 -12400 51350
rect -12600 51120 -12400 51150
rect -12100 51350 -12000 51380
rect -12100 51150 -12090 51350
rect -12020 51150 -12000 51350
rect -12100 51120 -12000 51150
rect -16000 51100 -15880 51120
rect -15620 51100 -15380 51120
rect -15120 51100 -14880 51120
rect -14620 51100 -14380 51120
rect -14120 51100 -13880 51120
rect -13620 51100 -13380 51120
rect -13120 51100 -12880 51120
rect -12620 51100 -12380 51120
rect -12120 51100 -12000 51120
rect -16000 51090 -12000 51100
rect -16000 51020 -15850 51090
rect -15650 51020 -15350 51090
rect -15150 51020 -14850 51090
rect -14650 51020 -14350 51090
rect -14150 51020 -13850 51090
rect -13650 51020 -13350 51090
rect -13150 51020 -12850 51090
rect -12650 51020 -12350 51090
rect -12150 51020 -12000 51090
rect -16000 50980 -12000 51020
rect -16000 50910 -15850 50980
rect -15650 50910 -15350 50980
rect -15150 50910 -14850 50980
rect -14650 50910 -14350 50980
rect -14150 50910 -13850 50980
rect -13650 50910 -13350 50980
rect -13150 50910 -12850 50980
rect -12650 50910 -12350 50980
rect -12150 50910 -12000 50980
rect -16000 50900 -12000 50910
rect -16000 50880 -15880 50900
rect -15620 50880 -15380 50900
rect -15120 50880 -14880 50900
rect -14620 50880 -14380 50900
rect -14120 50880 -13880 50900
rect -13620 50880 -13380 50900
rect -13120 50880 -12880 50900
rect -12620 50880 -12380 50900
rect -12120 50880 -12000 50900
rect -16000 50850 -15900 50880
rect -16000 50650 -15980 50850
rect -15910 50650 -15900 50850
rect -16000 50620 -15900 50650
rect -15600 50850 -15400 50880
rect -15600 50650 -15590 50850
rect -15520 50650 -15480 50850
rect -15410 50650 -15400 50850
rect -15600 50620 -15400 50650
rect -15100 50850 -14900 50880
rect -15100 50650 -15090 50850
rect -15020 50650 -14980 50850
rect -14910 50650 -14900 50850
rect -15100 50620 -14900 50650
rect -14600 50850 -14400 50880
rect -14600 50650 -14590 50850
rect -14520 50650 -14480 50850
rect -14410 50650 -14400 50850
rect -14600 50620 -14400 50650
rect -14100 50850 -13900 50880
rect -14100 50650 -14090 50850
rect -14020 50650 -13980 50850
rect -13910 50650 -13900 50850
rect -14100 50620 -13900 50650
rect -13600 50850 -13400 50880
rect -13600 50650 -13590 50850
rect -13520 50650 -13480 50850
rect -13410 50650 -13400 50850
rect -13600 50620 -13400 50650
rect -13100 50850 -12900 50880
rect -13100 50650 -13090 50850
rect -13020 50650 -12980 50850
rect -12910 50650 -12900 50850
rect -13100 50620 -12900 50650
rect -12600 50850 -12400 50880
rect -12600 50650 -12590 50850
rect -12520 50650 -12480 50850
rect -12410 50650 -12400 50850
rect -12600 50620 -12400 50650
rect -12100 50850 -12000 50880
rect -12100 50650 -12090 50850
rect -12020 50650 -12000 50850
rect -12100 50620 -12000 50650
rect -16000 50600 -15880 50620
rect -15620 50600 -15380 50620
rect -15120 50600 -14880 50620
rect -14620 50600 -14380 50620
rect -14120 50600 -13880 50620
rect -13620 50600 -13380 50620
rect -13120 50600 -12880 50620
rect -12620 50600 -12380 50620
rect -12120 50600 -12000 50620
rect -16000 50590 -12000 50600
rect -16000 50520 -15850 50590
rect -15650 50520 -15350 50590
rect -15150 50520 -14850 50590
rect -14650 50520 -14350 50590
rect -14150 50520 -13850 50590
rect -13650 50520 -13350 50590
rect -13150 50520 -12850 50590
rect -12650 50520 -12350 50590
rect -12150 50520 -12000 50590
rect -16000 50480 -12000 50520
rect -16000 50410 -15850 50480
rect -15650 50410 -15350 50480
rect -15150 50410 -14850 50480
rect -14650 50410 -14350 50480
rect -14150 50410 -13850 50480
rect -13650 50410 -13350 50480
rect -13150 50410 -12850 50480
rect -12650 50410 -12350 50480
rect -12150 50410 -12000 50480
rect -16000 50400 -12000 50410
rect -16000 50380 -15880 50400
rect -15620 50380 -15380 50400
rect -15120 50380 -14880 50400
rect -14620 50380 -14380 50400
rect -14120 50380 -13880 50400
rect -13620 50380 -13380 50400
rect -13120 50380 -12880 50400
rect -12620 50380 -12380 50400
rect -12120 50380 -12000 50400
rect -16000 50350 -15900 50380
rect -16000 50150 -15980 50350
rect -15910 50150 -15900 50350
rect -16000 50120 -15900 50150
rect -15600 50350 -15400 50380
rect -15600 50150 -15590 50350
rect -15520 50150 -15480 50350
rect -15410 50150 -15400 50350
rect -15600 50120 -15400 50150
rect -15100 50350 -14900 50380
rect -15100 50150 -15090 50350
rect -15020 50150 -14980 50350
rect -14910 50150 -14900 50350
rect -15100 50120 -14900 50150
rect -14600 50350 -14400 50380
rect -14600 50150 -14590 50350
rect -14520 50150 -14480 50350
rect -14410 50150 -14400 50350
rect -14600 50120 -14400 50150
rect -14100 50350 -13900 50380
rect -14100 50150 -14090 50350
rect -14020 50150 -13980 50350
rect -13910 50150 -13900 50350
rect -14100 50120 -13900 50150
rect -13600 50350 -13400 50380
rect -13600 50150 -13590 50350
rect -13520 50150 -13480 50350
rect -13410 50150 -13400 50350
rect -13600 50120 -13400 50150
rect -13100 50350 -12900 50380
rect -13100 50150 -13090 50350
rect -13020 50150 -12980 50350
rect -12910 50150 -12900 50350
rect -13100 50120 -12900 50150
rect -12600 50350 -12400 50380
rect -12600 50150 -12590 50350
rect -12520 50150 -12480 50350
rect -12410 50150 -12400 50350
rect -12600 50120 -12400 50150
rect -12100 50350 -12000 50380
rect -12100 50150 -12090 50350
rect -12020 50150 -12000 50350
rect -12100 50120 -12000 50150
rect -16000 50100 -15880 50120
rect -15620 50100 -15380 50120
rect -15120 50100 -14880 50120
rect -14620 50100 -14380 50120
rect -14120 50100 -13880 50120
rect -13620 50100 -13380 50120
rect -13120 50100 -12880 50120
rect -12620 50100 -12380 50120
rect -12120 50100 -12000 50120
rect -16000 50090 -12000 50100
rect -16000 50020 -15850 50090
rect -15650 50020 -15350 50090
rect -15150 50020 -14850 50090
rect -14650 50020 -14350 50090
rect -14150 50020 -13850 50090
rect -13650 50020 -13350 50090
rect -13150 50020 -12850 50090
rect -12650 50020 -12350 50090
rect -12150 50020 -12000 50090
rect -16000 49980 -12000 50020
rect 96000 85980 100000 86000
rect 96000 85910 96150 85980
rect 96350 85910 96650 85980
rect 96850 85910 97150 85980
rect 97350 85910 97650 85980
rect 97850 85910 98150 85980
rect 98350 85910 98650 85980
rect 98850 85910 99150 85980
rect 99350 85910 99650 85980
rect 99850 85910 100000 85980
rect 96000 85900 100000 85910
rect 96000 85880 96120 85900
rect 96380 85880 96620 85900
rect 96880 85880 97120 85900
rect 97380 85880 97620 85900
rect 97880 85880 98120 85900
rect 98380 85880 98620 85900
rect 98880 85880 99120 85900
rect 99380 85880 99620 85900
rect 99880 85880 100000 85900
rect 96000 85850 96100 85880
rect 96000 85650 96020 85850
rect 96090 85650 96100 85850
rect 96000 85620 96100 85650
rect 96400 85850 96600 85880
rect 96400 85650 96410 85850
rect 96480 85650 96520 85850
rect 96590 85650 96600 85850
rect 96400 85620 96600 85650
rect 96900 85850 97100 85880
rect 96900 85650 96910 85850
rect 96980 85650 97020 85850
rect 97090 85650 97100 85850
rect 96900 85620 97100 85650
rect 97400 85850 97600 85880
rect 97400 85650 97410 85850
rect 97480 85650 97520 85850
rect 97590 85650 97600 85850
rect 97400 85620 97600 85650
rect 97900 85850 98100 85880
rect 97900 85650 97910 85850
rect 97980 85650 98020 85850
rect 98090 85650 98100 85850
rect 97900 85620 98100 85650
rect 98400 85850 98600 85880
rect 98400 85650 98410 85850
rect 98480 85650 98520 85850
rect 98590 85650 98600 85850
rect 98400 85620 98600 85650
rect 98900 85850 99100 85880
rect 98900 85650 98910 85850
rect 98980 85650 99020 85850
rect 99090 85650 99100 85850
rect 98900 85620 99100 85650
rect 99400 85850 99600 85880
rect 99400 85650 99410 85850
rect 99480 85650 99520 85850
rect 99590 85650 99600 85850
rect 99400 85620 99600 85650
rect 99900 85850 100000 85880
rect 99900 85650 99910 85850
rect 99980 85650 100000 85850
rect 99900 85620 100000 85650
rect 96000 85600 96120 85620
rect 96380 85600 96620 85620
rect 96880 85600 97120 85620
rect 97380 85600 97620 85620
rect 97880 85600 98120 85620
rect 98380 85600 98620 85620
rect 98880 85600 99120 85620
rect 99380 85600 99620 85620
rect 99880 85600 100000 85620
rect 96000 85590 100000 85600
rect 96000 85520 96150 85590
rect 96350 85520 96650 85590
rect 96850 85520 97150 85590
rect 97350 85520 97650 85590
rect 97850 85520 98150 85590
rect 98350 85520 98650 85590
rect 98850 85520 99150 85590
rect 99350 85520 99650 85590
rect 99850 85520 100000 85590
rect 96000 85480 100000 85520
rect 96000 85410 96150 85480
rect 96350 85410 96650 85480
rect 96850 85410 97150 85480
rect 97350 85410 97650 85480
rect 97850 85410 98150 85480
rect 98350 85410 98650 85480
rect 98850 85410 99150 85480
rect 99350 85410 99650 85480
rect 99850 85410 100000 85480
rect 96000 85400 100000 85410
rect 96000 85380 96120 85400
rect 96380 85380 96620 85400
rect 96880 85380 97120 85400
rect 97380 85380 97620 85400
rect 97880 85380 98120 85400
rect 98380 85380 98620 85400
rect 98880 85380 99120 85400
rect 99380 85380 99620 85400
rect 99880 85380 100000 85400
rect 96000 85350 96100 85380
rect 96000 85150 96020 85350
rect 96090 85150 96100 85350
rect 96000 85120 96100 85150
rect 96400 85350 96600 85380
rect 96400 85150 96410 85350
rect 96480 85150 96520 85350
rect 96590 85150 96600 85350
rect 96400 85120 96600 85150
rect 96900 85350 97100 85380
rect 96900 85150 96910 85350
rect 96980 85150 97020 85350
rect 97090 85150 97100 85350
rect 96900 85120 97100 85150
rect 97400 85350 97600 85380
rect 97400 85150 97410 85350
rect 97480 85150 97520 85350
rect 97590 85150 97600 85350
rect 97400 85120 97600 85150
rect 97900 85350 98100 85380
rect 97900 85150 97910 85350
rect 97980 85150 98020 85350
rect 98090 85150 98100 85350
rect 97900 85120 98100 85150
rect 98400 85350 98600 85380
rect 98400 85150 98410 85350
rect 98480 85150 98520 85350
rect 98590 85150 98600 85350
rect 98400 85120 98600 85150
rect 98900 85350 99100 85380
rect 98900 85150 98910 85350
rect 98980 85150 99020 85350
rect 99090 85150 99100 85350
rect 98900 85120 99100 85150
rect 99400 85350 99600 85380
rect 99400 85150 99410 85350
rect 99480 85150 99520 85350
rect 99590 85150 99600 85350
rect 99400 85120 99600 85150
rect 99900 85350 100000 85380
rect 99900 85150 99910 85350
rect 99980 85150 100000 85350
rect 99900 85120 100000 85150
rect 96000 85100 96120 85120
rect 96380 85100 96620 85120
rect 96880 85100 97120 85120
rect 97380 85100 97620 85120
rect 97880 85100 98120 85120
rect 98380 85100 98620 85120
rect 98880 85100 99120 85120
rect 99380 85100 99620 85120
rect 99880 85100 100000 85120
rect 96000 85090 100000 85100
rect 96000 85020 96150 85090
rect 96350 85020 96650 85090
rect 96850 85020 97150 85090
rect 97350 85020 97650 85090
rect 97850 85020 98150 85090
rect 98350 85020 98650 85090
rect 98850 85020 99150 85090
rect 99350 85020 99650 85090
rect 99850 85020 100000 85090
rect 96000 84980 100000 85020
rect 96000 84910 96150 84980
rect 96350 84910 96650 84980
rect 96850 84910 97150 84980
rect 97350 84910 97650 84980
rect 97850 84910 98150 84980
rect 98350 84910 98650 84980
rect 98850 84910 99150 84980
rect 99350 84910 99650 84980
rect 99850 84910 100000 84980
rect 96000 84900 100000 84910
rect 96000 84880 96120 84900
rect 96380 84880 96620 84900
rect 96880 84880 97120 84900
rect 97380 84880 97620 84900
rect 97880 84880 98120 84900
rect 98380 84880 98620 84900
rect 98880 84880 99120 84900
rect 99380 84880 99620 84900
rect 99880 84880 100000 84900
rect 96000 84850 96100 84880
rect 96000 84650 96020 84850
rect 96090 84650 96100 84850
rect 96000 84620 96100 84650
rect 96400 84850 96600 84880
rect 96400 84650 96410 84850
rect 96480 84650 96520 84850
rect 96590 84650 96600 84850
rect 96400 84620 96600 84650
rect 96900 84850 97100 84880
rect 96900 84650 96910 84850
rect 96980 84650 97020 84850
rect 97090 84650 97100 84850
rect 96900 84620 97100 84650
rect 97400 84850 97600 84880
rect 97400 84650 97410 84850
rect 97480 84650 97520 84850
rect 97590 84650 97600 84850
rect 97400 84620 97600 84650
rect 97900 84850 98100 84880
rect 97900 84650 97910 84850
rect 97980 84650 98020 84850
rect 98090 84650 98100 84850
rect 97900 84620 98100 84650
rect 98400 84850 98600 84880
rect 98400 84650 98410 84850
rect 98480 84650 98520 84850
rect 98590 84650 98600 84850
rect 98400 84620 98600 84650
rect 98900 84850 99100 84880
rect 98900 84650 98910 84850
rect 98980 84650 99020 84850
rect 99090 84650 99100 84850
rect 98900 84620 99100 84650
rect 99400 84850 99600 84880
rect 99400 84650 99410 84850
rect 99480 84650 99520 84850
rect 99590 84650 99600 84850
rect 99400 84620 99600 84650
rect 99900 84850 100000 84880
rect 99900 84650 99910 84850
rect 99980 84650 100000 84850
rect 99900 84620 100000 84650
rect 96000 84600 96120 84620
rect 96380 84600 96620 84620
rect 96880 84600 97120 84620
rect 97380 84600 97620 84620
rect 97880 84600 98120 84620
rect 98380 84600 98620 84620
rect 98880 84600 99120 84620
rect 99380 84600 99620 84620
rect 99880 84600 100000 84620
rect 96000 84590 100000 84600
rect 96000 84520 96150 84590
rect 96350 84520 96650 84590
rect 96850 84520 97150 84590
rect 97350 84520 97650 84590
rect 97850 84520 98150 84590
rect 98350 84520 98650 84590
rect 98850 84520 99150 84590
rect 99350 84520 99650 84590
rect 99850 84520 100000 84590
rect 96000 84480 100000 84520
rect 96000 84410 96150 84480
rect 96350 84410 96650 84480
rect 96850 84410 97150 84480
rect 97350 84410 97650 84480
rect 97850 84410 98150 84480
rect 98350 84410 98650 84480
rect 98850 84410 99150 84480
rect 99350 84410 99650 84480
rect 99850 84410 100000 84480
rect 96000 84400 100000 84410
rect 96000 84380 96120 84400
rect 96380 84380 96620 84400
rect 96880 84380 97120 84400
rect 97380 84380 97620 84400
rect 97880 84380 98120 84400
rect 98380 84380 98620 84400
rect 98880 84380 99120 84400
rect 99380 84380 99620 84400
rect 99880 84380 100000 84400
rect 96000 84350 96100 84380
rect 96000 84150 96020 84350
rect 96090 84150 96100 84350
rect 96000 84120 96100 84150
rect 96400 84350 96600 84380
rect 96400 84150 96410 84350
rect 96480 84150 96520 84350
rect 96590 84150 96600 84350
rect 96400 84120 96600 84150
rect 96900 84350 97100 84380
rect 96900 84150 96910 84350
rect 96980 84150 97020 84350
rect 97090 84150 97100 84350
rect 96900 84120 97100 84150
rect 97400 84350 97600 84380
rect 97400 84150 97410 84350
rect 97480 84150 97520 84350
rect 97590 84150 97600 84350
rect 97400 84120 97600 84150
rect 97900 84350 98100 84380
rect 97900 84150 97910 84350
rect 97980 84150 98020 84350
rect 98090 84150 98100 84350
rect 97900 84120 98100 84150
rect 98400 84350 98600 84380
rect 98400 84150 98410 84350
rect 98480 84150 98520 84350
rect 98590 84150 98600 84350
rect 98400 84120 98600 84150
rect 98900 84350 99100 84380
rect 98900 84150 98910 84350
rect 98980 84150 99020 84350
rect 99090 84150 99100 84350
rect 98900 84120 99100 84150
rect 99400 84350 99600 84380
rect 99400 84150 99410 84350
rect 99480 84150 99520 84350
rect 99590 84150 99600 84350
rect 99400 84120 99600 84150
rect 99900 84350 100000 84380
rect 99900 84150 99910 84350
rect 99980 84150 100000 84350
rect 99900 84120 100000 84150
rect 96000 84100 96120 84120
rect 96380 84100 96620 84120
rect 96880 84100 97120 84120
rect 97380 84100 97620 84120
rect 97880 84100 98120 84120
rect 98380 84100 98620 84120
rect 98880 84100 99120 84120
rect 99380 84100 99620 84120
rect 99880 84100 100000 84120
rect 96000 84090 100000 84100
rect 96000 84020 96150 84090
rect 96350 84020 96650 84090
rect 96850 84020 97150 84090
rect 97350 84020 97650 84090
rect 97850 84020 98150 84090
rect 98350 84020 98650 84090
rect 98850 84020 99150 84090
rect 99350 84020 99650 84090
rect 99850 84020 100000 84090
rect 96000 83980 100000 84020
rect 96000 83910 96150 83980
rect 96350 83910 96650 83980
rect 96850 83910 97150 83980
rect 97350 83910 97650 83980
rect 97850 83910 98150 83980
rect 98350 83910 98650 83980
rect 98850 83910 99150 83980
rect 99350 83910 99650 83980
rect 99850 83910 100000 83980
rect 96000 83900 100000 83910
rect 96000 83880 96120 83900
rect 96380 83880 96620 83900
rect 96880 83880 97120 83900
rect 97380 83880 97620 83900
rect 97880 83880 98120 83900
rect 98380 83880 98620 83900
rect 98880 83880 99120 83900
rect 99380 83880 99620 83900
rect 99880 83880 100000 83900
rect 96000 83850 96100 83880
rect 96000 83650 96020 83850
rect 96090 83650 96100 83850
rect 96000 83620 96100 83650
rect 96400 83850 96600 83880
rect 96400 83650 96410 83850
rect 96480 83650 96520 83850
rect 96590 83650 96600 83850
rect 96400 83620 96600 83650
rect 96900 83850 97100 83880
rect 96900 83650 96910 83850
rect 96980 83650 97020 83850
rect 97090 83650 97100 83850
rect 96900 83620 97100 83650
rect 97400 83850 97600 83880
rect 97400 83650 97410 83850
rect 97480 83650 97520 83850
rect 97590 83650 97600 83850
rect 97400 83620 97600 83650
rect 97900 83850 98100 83880
rect 97900 83650 97910 83850
rect 97980 83650 98020 83850
rect 98090 83650 98100 83850
rect 97900 83620 98100 83650
rect 98400 83850 98600 83880
rect 98400 83650 98410 83850
rect 98480 83650 98520 83850
rect 98590 83650 98600 83850
rect 98400 83620 98600 83650
rect 98900 83850 99100 83880
rect 98900 83650 98910 83850
rect 98980 83650 99020 83850
rect 99090 83650 99100 83850
rect 98900 83620 99100 83650
rect 99400 83850 99600 83880
rect 99400 83650 99410 83850
rect 99480 83650 99520 83850
rect 99590 83650 99600 83850
rect 99400 83620 99600 83650
rect 99900 83850 100000 83880
rect 99900 83650 99910 83850
rect 99980 83650 100000 83850
rect 99900 83620 100000 83650
rect 96000 83600 96120 83620
rect 96380 83600 96620 83620
rect 96880 83600 97120 83620
rect 97380 83600 97620 83620
rect 97880 83600 98120 83620
rect 98380 83600 98620 83620
rect 98880 83600 99120 83620
rect 99380 83600 99620 83620
rect 99880 83600 100000 83620
rect 96000 83590 100000 83600
rect 96000 83520 96150 83590
rect 96350 83520 96650 83590
rect 96850 83520 97150 83590
rect 97350 83520 97650 83590
rect 97850 83520 98150 83590
rect 98350 83520 98650 83590
rect 98850 83520 99150 83590
rect 99350 83520 99650 83590
rect 99850 83520 100000 83590
rect 96000 83480 100000 83520
rect 96000 83410 96150 83480
rect 96350 83410 96650 83480
rect 96850 83410 97150 83480
rect 97350 83410 97650 83480
rect 97850 83410 98150 83480
rect 98350 83410 98650 83480
rect 98850 83410 99150 83480
rect 99350 83410 99650 83480
rect 99850 83410 100000 83480
rect 96000 83400 100000 83410
rect 96000 83380 96120 83400
rect 96380 83380 96620 83400
rect 96880 83380 97120 83400
rect 97380 83380 97620 83400
rect 97880 83380 98120 83400
rect 98380 83380 98620 83400
rect 98880 83380 99120 83400
rect 99380 83380 99620 83400
rect 99880 83380 100000 83400
rect 96000 83350 96100 83380
rect 96000 83150 96020 83350
rect 96090 83150 96100 83350
rect 96000 83120 96100 83150
rect 96400 83350 96600 83380
rect 96400 83150 96410 83350
rect 96480 83150 96520 83350
rect 96590 83150 96600 83350
rect 96400 83120 96600 83150
rect 96900 83350 97100 83380
rect 96900 83150 96910 83350
rect 96980 83150 97020 83350
rect 97090 83150 97100 83350
rect 96900 83120 97100 83150
rect 97400 83350 97600 83380
rect 97400 83150 97410 83350
rect 97480 83150 97520 83350
rect 97590 83150 97600 83350
rect 97400 83120 97600 83150
rect 97900 83350 98100 83380
rect 97900 83150 97910 83350
rect 97980 83150 98020 83350
rect 98090 83150 98100 83350
rect 97900 83120 98100 83150
rect 98400 83350 98600 83380
rect 98400 83150 98410 83350
rect 98480 83150 98520 83350
rect 98590 83150 98600 83350
rect 98400 83120 98600 83150
rect 98900 83350 99100 83380
rect 98900 83150 98910 83350
rect 98980 83150 99020 83350
rect 99090 83150 99100 83350
rect 98900 83120 99100 83150
rect 99400 83350 99600 83380
rect 99400 83150 99410 83350
rect 99480 83150 99520 83350
rect 99590 83150 99600 83350
rect 99400 83120 99600 83150
rect 99900 83350 100000 83380
rect 99900 83150 99910 83350
rect 99980 83150 100000 83350
rect 99900 83120 100000 83150
rect 96000 83100 96120 83120
rect 96380 83100 96620 83120
rect 96880 83100 97120 83120
rect 97380 83100 97620 83120
rect 97880 83100 98120 83120
rect 98380 83100 98620 83120
rect 98880 83100 99120 83120
rect 99380 83100 99620 83120
rect 99880 83100 100000 83120
rect 96000 83090 100000 83100
rect 96000 83020 96150 83090
rect 96350 83020 96650 83090
rect 96850 83020 97150 83090
rect 97350 83020 97650 83090
rect 97850 83020 98150 83090
rect 98350 83020 98650 83090
rect 98850 83020 99150 83090
rect 99350 83020 99650 83090
rect 99850 83020 100000 83090
rect 96000 82980 100000 83020
rect 96000 82910 96150 82980
rect 96350 82910 96650 82980
rect 96850 82910 97150 82980
rect 97350 82910 97650 82980
rect 97850 82910 98150 82980
rect 98350 82910 98650 82980
rect 98850 82910 99150 82980
rect 99350 82910 99650 82980
rect 99850 82910 100000 82980
rect 96000 82900 100000 82910
rect 96000 82880 96120 82900
rect 96380 82880 96620 82900
rect 96880 82880 97120 82900
rect 97380 82880 97620 82900
rect 97880 82880 98120 82900
rect 98380 82880 98620 82900
rect 98880 82880 99120 82900
rect 99380 82880 99620 82900
rect 99880 82880 100000 82900
rect 96000 82850 96100 82880
rect 96000 82650 96020 82850
rect 96090 82650 96100 82850
rect 96000 82620 96100 82650
rect 96400 82850 96600 82880
rect 96400 82650 96410 82850
rect 96480 82650 96520 82850
rect 96590 82650 96600 82850
rect 96400 82620 96600 82650
rect 96900 82850 97100 82880
rect 96900 82650 96910 82850
rect 96980 82650 97020 82850
rect 97090 82650 97100 82850
rect 96900 82620 97100 82650
rect 97400 82850 97600 82880
rect 97400 82650 97410 82850
rect 97480 82650 97520 82850
rect 97590 82650 97600 82850
rect 97400 82620 97600 82650
rect 97900 82850 98100 82880
rect 97900 82650 97910 82850
rect 97980 82650 98020 82850
rect 98090 82650 98100 82850
rect 97900 82620 98100 82650
rect 98400 82850 98600 82880
rect 98400 82650 98410 82850
rect 98480 82650 98520 82850
rect 98590 82650 98600 82850
rect 98400 82620 98600 82650
rect 98900 82850 99100 82880
rect 98900 82650 98910 82850
rect 98980 82650 99020 82850
rect 99090 82650 99100 82850
rect 98900 82620 99100 82650
rect 99400 82850 99600 82880
rect 99400 82650 99410 82850
rect 99480 82650 99520 82850
rect 99590 82650 99600 82850
rect 99400 82620 99600 82650
rect 99900 82850 100000 82880
rect 99900 82650 99910 82850
rect 99980 82650 100000 82850
rect 99900 82620 100000 82650
rect 96000 82600 96120 82620
rect 96380 82600 96620 82620
rect 96880 82600 97120 82620
rect 97380 82600 97620 82620
rect 97880 82600 98120 82620
rect 98380 82600 98620 82620
rect 98880 82600 99120 82620
rect 99380 82600 99620 82620
rect 99880 82600 100000 82620
rect 96000 82590 100000 82600
rect 96000 82520 96150 82590
rect 96350 82520 96650 82590
rect 96850 82520 97150 82590
rect 97350 82520 97650 82590
rect 97850 82520 98150 82590
rect 98350 82520 98650 82590
rect 98850 82520 99150 82590
rect 99350 82520 99650 82590
rect 99850 82520 100000 82590
rect 96000 82480 100000 82520
rect 96000 82410 96150 82480
rect 96350 82410 96650 82480
rect 96850 82410 97150 82480
rect 97350 82410 97650 82480
rect 97850 82410 98150 82480
rect 98350 82410 98650 82480
rect 98850 82410 99150 82480
rect 99350 82410 99650 82480
rect 99850 82410 100000 82480
rect 96000 82400 100000 82410
rect 96000 82380 96120 82400
rect 96380 82380 96620 82400
rect 96880 82380 97120 82400
rect 97380 82380 97620 82400
rect 97880 82380 98120 82400
rect 98380 82380 98620 82400
rect 98880 82380 99120 82400
rect 99380 82380 99620 82400
rect 99880 82380 100000 82400
rect 96000 82350 96100 82380
rect 96000 82150 96020 82350
rect 96090 82150 96100 82350
rect 96000 82120 96100 82150
rect 96400 82350 96600 82380
rect 96400 82150 96410 82350
rect 96480 82150 96520 82350
rect 96590 82150 96600 82350
rect 96400 82120 96600 82150
rect 96900 82350 97100 82380
rect 96900 82150 96910 82350
rect 96980 82150 97020 82350
rect 97090 82150 97100 82350
rect 96900 82120 97100 82150
rect 97400 82350 97600 82380
rect 97400 82150 97410 82350
rect 97480 82150 97520 82350
rect 97590 82150 97600 82350
rect 97400 82120 97600 82150
rect 97900 82350 98100 82380
rect 97900 82150 97910 82350
rect 97980 82150 98020 82350
rect 98090 82150 98100 82350
rect 97900 82120 98100 82150
rect 98400 82350 98600 82380
rect 98400 82150 98410 82350
rect 98480 82150 98520 82350
rect 98590 82150 98600 82350
rect 98400 82120 98600 82150
rect 98900 82350 99100 82380
rect 98900 82150 98910 82350
rect 98980 82150 99020 82350
rect 99090 82150 99100 82350
rect 98900 82120 99100 82150
rect 99400 82350 99600 82380
rect 99400 82150 99410 82350
rect 99480 82150 99520 82350
rect 99590 82150 99600 82350
rect 99400 82120 99600 82150
rect 99900 82350 100000 82380
rect 99900 82150 99910 82350
rect 99980 82150 100000 82350
rect 99900 82120 100000 82150
rect 96000 82100 96120 82120
rect 96380 82100 96620 82120
rect 96880 82100 97120 82120
rect 97380 82100 97620 82120
rect 97880 82100 98120 82120
rect 98380 82100 98620 82120
rect 98880 82100 99120 82120
rect 99380 82100 99620 82120
rect 99880 82100 100000 82120
rect 96000 82090 100000 82100
rect 96000 82020 96150 82090
rect 96350 82020 96650 82090
rect 96850 82020 97150 82090
rect 97350 82020 97650 82090
rect 97850 82020 98150 82090
rect 98350 82020 98650 82090
rect 98850 82020 99150 82090
rect 99350 82020 99650 82090
rect 99850 82020 100000 82090
rect 96000 81980 100000 82020
rect 96000 81910 96150 81980
rect 96350 81910 96650 81980
rect 96850 81910 97150 81980
rect 97350 81910 97650 81980
rect 97850 81910 98150 81980
rect 98350 81910 98650 81980
rect 98850 81910 99150 81980
rect 99350 81910 99650 81980
rect 99850 81910 100000 81980
rect 96000 81900 100000 81910
rect 96000 81880 96120 81900
rect 96380 81880 96620 81900
rect 96880 81880 97120 81900
rect 97380 81880 97620 81900
rect 97880 81880 98120 81900
rect 98380 81880 98620 81900
rect 98880 81880 99120 81900
rect 99380 81880 99620 81900
rect 99880 81880 100000 81900
rect 96000 81850 96100 81880
rect 96000 81650 96020 81850
rect 96090 81650 96100 81850
rect 96000 81620 96100 81650
rect 96400 81850 96600 81880
rect 96400 81650 96410 81850
rect 96480 81650 96520 81850
rect 96590 81650 96600 81850
rect 96400 81620 96600 81650
rect 96900 81850 97100 81880
rect 96900 81650 96910 81850
rect 96980 81650 97020 81850
rect 97090 81650 97100 81850
rect 96900 81620 97100 81650
rect 97400 81850 97600 81880
rect 97400 81650 97410 81850
rect 97480 81650 97520 81850
rect 97590 81650 97600 81850
rect 97400 81620 97600 81650
rect 97900 81850 98100 81880
rect 97900 81650 97910 81850
rect 97980 81650 98020 81850
rect 98090 81650 98100 81850
rect 97900 81620 98100 81650
rect 98400 81850 98600 81880
rect 98400 81650 98410 81850
rect 98480 81650 98520 81850
rect 98590 81650 98600 81850
rect 98400 81620 98600 81650
rect 98900 81850 99100 81880
rect 98900 81650 98910 81850
rect 98980 81650 99020 81850
rect 99090 81650 99100 81850
rect 98900 81620 99100 81650
rect 99400 81850 99600 81880
rect 99400 81650 99410 81850
rect 99480 81650 99520 81850
rect 99590 81650 99600 81850
rect 99400 81620 99600 81650
rect 99900 81850 100000 81880
rect 99900 81650 99910 81850
rect 99980 81650 100000 81850
rect 99900 81620 100000 81650
rect 96000 81600 96120 81620
rect 96380 81600 96620 81620
rect 96880 81600 97120 81620
rect 97380 81600 97620 81620
rect 97880 81600 98120 81620
rect 98380 81600 98620 81620
rect 98880 81600 99120 81620
rect 99380 81600 99620 81620
rect 99880 81600 100000 81620
rect 96000 81590 100000 81600
rect 96000 81520 96150 81590
rect 96350 81520 96650 81590
rect 96850 81520 97150 81590
rect 97350 81520 97650 81590
rect 97850 81520 98150 81590
rect 98350 81520 98650 81590
rect 98850 81520 99150 81590
rect 99350 81520 99650 81590
rect 99850 81520 100000 81590
rect 96000 81480 100000 81520
rect 96000 81410 96150 81480
rect 96350 81410 96650 81480
rect 96850 81410 97150 81480
rect 97350 81410 97650 81480
rect 97850 81410 98150 81480
rect 98350 81410 98650 81480
rect 98850 81410 99150 81480
rect 99350 81410 99650 81480
rect 99850 81410 100000 81480
rect 96000 81400 100000 81410
rect 96000 81380 96120 81400
rect 96380 81380 96620 81400
rect 96880 81380 97120 81400
rect 97380 81380 97620 81400
rect 97880 81380 98120 81400
rect 98380 81380 98620 81400
rect 98880 81380 99120 81400
rect 99380 81380 99620 81400
rect 99880 81380 100000 81400
rect 96000 81350 96100 81380
rect 96000 81150 96020 81350
rect 96090 81150 96100 81350
rect 96000 81120 96100 81150
rect 96400 81350 96600 81380
rect 96400 81150 96410 81350
rect 96480 81150 96520 81350
rect 96590 81150 96600 81350
rect 96400 81120 96600 81150
rect 96900 81350 97100 81380
rect 96900 81150 96910 81350
rect 96980 81150 97020 81350
rect 97090 81150 97100 81350
rect 96900 81120 97100 81150
rect 97400 81350 97600 81380
rect 97400 81150 97410 81350
rect 97480 81150 97520 81350
rect 97590 81150 97600 81350
rect 97400 81120 97600 81150
rect 97900 81350 98100 81380
rect 97900 81150 97910 81350
rect 97980 81150 98020 81350
rect 98090 81150 98100 81350
rect 97900 81120 98100 81150
rect 98400 81350 98600 81380
rect 98400 81150 98410 81350
rect 98480 81150 98520 81350
rect 98590 81150 98600 81350
rect 98400 81120 98600 81150
rect 98900 81350 99100 81380
rect 98900 81150 98910 81350
rect 98980 81150 99020 81350
rect 99090 81150 99100 81350
rect 98900 81120 99100 81150
rect 99400 81350 99600 81380
rect 99400 81150 99410 81350
rect 99480 81150 99520 81350
rect 99590 81150 99600 81350
rect 99400 81120 99600 81150
rect 99900 81350 100000 81380
rect 99900 81150 99910 81350
rect 99980 81150 100000 81350
rect 99900 81120 100000 81150
rect 96000 81100 96120 81120
rect 96380 81100 96620 81120
rect 96880 81100 97120 81120
rect 97380 81100 97620 81120
rect 97880 81100 98120 81120
rect 98380 81100 98620 81120
rect 98880 81100 99120 81120
rect 99380 81100 99620 81120
rect 99880 81100 100000 81120
rect 96000 81090 100000 81100
rect 96000 81020 96150 81090
rect 96350 81020 96650 81090
rect 96850 81020 97150 81090
rect 97350 81020 97650 81090
rect 97850 81020 98150 81090
rect 98350 81020 98650 81090
rect 98850 81020 99150 81090
rect 99350 81020 99650 81090
rect 99850 81020 100000 81090
rect 96000 80980 100000 81020
rect 96000 80910 96150 80980
rect 96350 80910 96650 80980
rect 96850 80910 97150 80980
rect 97350 80910 97650 80980
rect 97850 80910 98150 80980
rect 98350 80910 98650 80980
rect 98850 80910 99150 80980
rect 99350 80910 99650 80980
rect 99850 80910 100000 80980
rect 96000 80900 100000 80910
rect 96000 80880 96120 80900
rect 96380 80880 96620 80900
rect 96880 80880 97120 80900
rect 97380 80880 97620 80900
rect 97880 80880 98120 80900
rect 98380 80880 98620 80900
rect 98880 80880 99120 80900
rect 99380 80880 99620 80900
rect 99880 80880 100000 80900
rect 96000 80850 96100 80880
rect 96000 80650 96020 80850
rect 96090 80650 96100 80850
rect 96000 80620 96100 80650
rect 96400 80850 96600 80880
rect 96400 80650 96410 80850
rect 96480 80650 96520 80850
rect 96590 80650 96600 80850
rect 96400 80620 96600 80650
rect 96900 80850 97100 80880
rect 96900 80650 96910 80850
rect 96980 80650 97020 80850
rect 97090 80650 97100 80850
rect 96900 80620 97100 80650
rect 97400 80850 97600 80880
rect 97400 80650 97410 80850
rect 97480 80650 97520 80850
rect 97590 80650 97600 80850
rect 97400 80620 97600 80650
rect 97900 80850 98100 80880
rect 97900 80650 97910 80850
rect 97980 80650 98020 80850
rect 98090 80650 98100 80850
rect 97900 80620 98100 80650
rect 98400 80850 98600 80880
rect 98400 80650 98410 80850
rect 98480 80650 98520 80850
rect 98590 80650 98600 80850
rect 98400 80620 98600 80650
rect 98900 80850 99100 80880
rect 98900 80650 98910 80850
rect 98980 80650 99020 80850
rect 99090 80650 99100 80850
rect 98900 80620 99100 80650
rect 99400 80850 99600 80880
rect 99400 80650 99410 80850
rect 99480 80650 99520 80850
rect 99590 80650 99600 80850
rect 99400 80620 99600 80650
rect 99900 80850 100000 80880
rect 99900 80650 99910 80850
rect 99980 80650 100000 80850
rect 99900 80620 100000 80650
rect 96000 80600 96120 80620
rect 96380 80600 96620 80620
rect 96880 80600 97120 80620
rect 97380 80600 97620 80620
rect 97880 80600 98120 80620
rect 98380 80600 98620 80620
rect 98880 80600 99120 80620
rect 99380 80600 99620 80620
rect 99880 80600 100000 80620
rect 96000 80590 100000 80600
rect 96000 80520 96150 80590
rect 96350 80520 96650 80590
rect 96850 80520 97150 80590
rect 97350 80520 97650 80590
rect 97850 80520 98150 80590
rect 98350 80520 98650 80590
rect 98850 80520 99150 80590
rect 99350 80520 99650 80590
rect 99850 80520 100000 80590
rect 96000 80480 100000 80520
rect 96000 80410 96150 80480
rect 96350 80410 96650 80480
rect 96850 80410 97150 80480
rect 97350 80410 97650 80480
rect 97850 80410 98150 80480
rect 98350 80410 98650 80480
rect 98850 80410 99150 80480
rect 99350 80410 99650 80480
rect 99850 80410 100000 80480
rect 96000 80400 100000 80410
rect 96000 80380 96120 80400
rect 96380 80380 96620 80400
rect 96880 80380 97120 80400
rect 97380 80380 97620 80400
rect 97880 80380 98120 80400
rect 98380 80380 98620 80400
rect 98880 80380 99120 80400
rect 99380 80380 99620 80400
rect 99880 80380 100000 80400
rect 96000 80350 96100 80380
rect 96000 80150 96020 80350
rect 96090 80150 96100 80350
rect 96000 80120 96100 80150
rect 96400 80350 96600 80380
rect 96400 80150 96410 80350
rect 96480 80150 96520 80350
rect 96590 80150 96600 80350
rect 96400 80120 96600 80150
rect 96900 80350 97100 80380
rect 96900 80150 96910 80350
rect 96980 80150 97020 80350
rect 97090 80150 97100 80350
rect 96900 80120 97100 80150
rect 97400 80350 97600 80380
rect 97400 80150 97410 80350
rect 97480 80150 97520 80350
rect 97590 80150 97600 80350
rect 97400 80120 97600 80150
rect 97900 80350 98100 80380
rect 97900 80150 97910 80350
rect 97980 80150 98020 80350
rect 98090 80150 98100 80350
rect 97900 80120 98100 80150
rect 98400 80350 98600 80380
rect 98400 80150 98410 80350
rect 98480 80150 98520 80350
rect 98590 80150 98600 80350
rect 98400 80120 98600 80150
rect 98900 80350 99100 80380
rect 98900 80150 98910 80350
rect 98980 80150 99020 80350
rect 99090 80150 99100 80350
rect 98900 80120 99100 80150
rect 99400 80350 99600 80380
rect 99400 80150 99410 80350
rect 99480 80150 99520 80350
rect 99590 80150 99600 80350
rect 99400 80120 99600 80150
rect 99900 80350 100000 80380
rect 99900 80150 99910 80350
rect 99980 80150 100000 80350
rect 99900 80120 100000 80150
rect 96000 80100 96120 80120
rect 96380 80100 96620 80120
rect 96880 80100 97120 80120
rect 97380 80100 97620 80120
rect 97880 80100 98120 80120
rect 98380 80100 98620 80120
rect 98880 80100 99120 80120
rect 99380 80100 99620 80120
rect 99880 80100 100000 80120
rect 96000 80090 100000 80100
rect 96000 80020 96150 80090
rect 96350 80020 96650 80090
rect 96850 80020 97150 80090
rect 97350 80020 97650 80090
rect 97850 80020 98150 80090
rect 98350 80020 98650 80090
rect 98850 80020 99150 80090
rect 99350 80020 99650 80090
rect 99850 80020 100000 80090
rect 96000 79980 100000 80020
rect 96000 79910 96150 79980
rect 96350 79910 96650 79980
rect 96850 79910 97150 79980
rect 97350 79910 97650 79980
rect 97850 79910 98150 79980
rect 98350 79910 98650 79980
rect 98850 79910 99150 79980
rect 99350 79910 99650 79980
rect 99850 79910 100000 79980
rect 96000 79900 100000 79910
rect 96000 79880 96120 79900
rect 96380 79880 96620 79900
rect 96880 79880 97120 79900
rect 97380 79880 97620 79900
rect 97880 79880 98120 79900
rect 98380 79880 98620 79900
rect 98880 79880 99120 79900
rect 99380 79880 99620 79900
rect 99880 79880 100000 79900
rect 96000 79850 96100 79880
rect 96000 79650 96020 79850
rect 96090 79650 96100 79850
rect 96000 79620 96100 79650
rect 96400 79850 96600 79880
rect 96400 79650 96410 79850
rect 96480 79650 96520 79850
rect 96590 79650 96600 79850
rect 96400 79620 96600 79650
rect 96900 79850 97100 79880
rect 96900 79650 96910 79850
rect 96980 79650 97020 79850
rect 97090 79650 97100 79850
rect 96900 79620 97100 79650
rect 97400 79850 97600 79880
rect 97400 79650 97410 79850
rect 97480 79650 97520 79850
rect 97590 79650 97600 79850
rect 97400 79620 97600 79650
rect 97900 79850 98100 79880
rect 97900 79650 97910 79850
rect 97980 79650 98020 79850
rect 98090 79650 98100 79850
rect 97900 79620 98100 79650
rect 98400 79850 98600 79880
rect 98400 79650 98410 79850
rect 98480 79650 98520 79850
rect 98590 79650 98600 79850
rect 98400 79620 98600 79650
rect 98900 79850 99100 79880
rect 98900 79650 98910 79850
rect 98980 79650 99020 79850
rect 99090 79650 99100 79850
rect 98900 79620 99100 79650
rect 99400 79850 99600 79880
rect 99400 79650 99410 79850
rect 99480 79650 99520 79850
rect 99590 79650 99600 79850
rect 99400 79620 99600 79650
rect 99900 79850 100000 79880
rect 99900 79650 99910 79850
rect 99980 79650 100000 79850
rect 99900 79620 100000 79650
rect 96000 79600 96120 79620
rect 96380 79600 96620 79620
rect 96880 79600 97120 79620
rect 97380 79600 97620 79620
rect 97880 79600 98120 79620
rect 98380 79600 98620 79620
rect 98880 79600 99120 79620
rect 99380 79600 99620 79620
rect 99880 79600 100000 79620
rect 96000 79590 100000 79600
rect 96000 79520 96150 79590
rect 96350 79520 96650 79590
rect 96850 79520 97150 79590
rect 97350 79520 97650 79590
rect 97850 79520 98150 79590
rect 98350 79520 98650 79590
rect 98850 79520 99150 79590
rect 99350 79520 99650 79590
rect 99850 79520 100000 79590
rect 96000 79480 100000 79520
rect 96000 79410 96150 79480
rect 96350 79410 96650 79480
rect 96850 79410 97150 79480
rect 97350 79410 97650 79480
rect 97850 79410 98150 79480
rect 98350 79410 98650 79480
rect 98850 79410 99150 79480
rect 99350 79410 99650 79480
rect 99850 79410 100000 79480
rect 96000 79400 100000 79410
rect 96000 79380 96120 79400
rect 96380 79380 96620 79400
rect 96880 79380 97120 79400
rect 97380 79380 97620 79400
rect 97880 79380 98120 79400
rect 98380 79380 98620 79400
rect 98880 79380 99120 79400
rect 99380 79380 99620 79400
rect 99880 79380 100000 79400
rect 96000 79350 96100 79380
rect 96000 79150 96020 79350
rect 96090 79150 96100 79350
rect 96000 79120 96100 79150
rect 96400 79350 96600 79380
rect 96400 79150 96410 79350
rect 96480 79150 96520 79350
rect 96590 79150 96600 79350
rect 96400 79120 96600 79150
rect 96900 79350 97100 79380
rect 96900 79150 96910 79350
rect 96980 79150 97020 79350
rect 97090 79150 97100 79350
rect 96900 79120 97100 79150
rect 97400 79350 97600 79380
rect 97400 79150 97410 79350
rect 97480 79150 97520 79350
rect 97590 79150 97600 79350
rect 97400 79120 97600 79150
rect 97900 79350 98100 79380
rect 97900 79150 97910 79350
rect 97980 79150 98020 79350
rect 98090 79150 98100 79350
rect 97900 79120 98100 79150
rect 98400 79350 98600 79380
rect 98400 79150 98410 79350
rect 98480 79150 98520 79350
rect 98590 79150 98600 79350
rect 98400 79120 98600 79150
rect 98900 79350 99100 79380
rect 98900 79150 98910 79350
rect 98980 79150 99020 79350
rect 99090 79150 99100 79350
rect 98900 79120 99100 79150
rect 99400 79350 99600 79380
rect 99400 79150 99410 79350
rect 99480 79150 99520 79350
rect 99590 79150 99600 79350
rect 99400 79120 99600 79150
rect 99900 79350 100000 79380
rect 99900 79150 99910 79350
rect 99980 79150 100000 79350
rect 99900 79120 100000 79150
rect 96000 79100 96120 79120
rect 96380 79100 96620 79120
rect 96880 79100 97120 79120
rect 97380 79100 97620 79120
rect 97880 79100 98120 79120
rect 98380 79100 98620 79120
rect 98880 79100 99120 79120
rect 99380 79100 99620 79120
rect 99880 79100 100000 79120
rect 96000 79090 100000 79100
rect 96000 79020 96150 79090
rect 96350 79020 96650 79090
rect 96850 79020 97150 79090
rect 97350 79020 97650 79090
rect 97850 79020 98150 79090
rect 98350 79020 98650 79090
rect 98850 79020 99150 79090
rect 99350 79020 99650 79090
rect 99850 79020 100000 79090
rect 96000 78980 100000 79020
rect 96000 78910 96150 78980
rect 96350 78910 96650 78980
rect 96850 78910 97150 78980
rect 97350 78910 97650 78980
rect 97850 78910 98150 78980
rect 98350 78910 98650 78980
rect 98850 78910 99150 78980
rect 99350 78910 99650 78980
rect 99850 78910 100000 78980
rect 96000 78900 100000 78910
rect 96000 78880 96120 78900
rect 96380 78880 96620 78900
rect 96880 78880 97120 78900
rect 97380 78880 97620 78900
rect 97880 78880 98120 78900
rect 98380 78880 98620 78900
rect 98880 78880 99120 78900
rect 99380 78880 99620 78900
rect 99880 78880 100000 78900
rect 96000 78850 96100 78880
rect 96000 78650 96020 78850
rect 96090 78650 96100 78850
rect 96000 78620 96100 78650
rect 96400 78850 96600 78880
rect 96400 78650 96410 78850
rect 96480 78650 96520 78850
rect 96590 78650 96600 78850
rect 96400 78620 96600 78650
rect 96900 78850 97100 78880
rect 96900 78650 96910 78850
rect 96980 78650 97020 78850
rect 97090 78650 97100 78850
rect 96900 78620 97100 78650
rect 97400 78850 97600 78880
rect 97400 78650 97410 78850
rect 97480 78650 97520 78850
rect 97590 78650 97600 78850
rect 97400 78620 97600 78650
rect 97900 78850 98100 78880
rect 97900 78650 97910 78850
rect 97980 78650 98020 78850
rect 98090 78650 98100 78850
rect 97900 78620 98100 78650
rect 98400 78850 98600 78880
rect 98400 78650 98410 78850
rect 98480 78650 98520 78850
rect 98590 78650 98600 78850
rect 98400 78620 98600 78650
rect 98900 78850 99100 78880
rect 98900 78650 98910 78850
rect 98980 78650 99020 78850
rect 99090 78650 99100 78850
rect 98900 78620 99100 78650
rect 99400 78850 99600 78880
rect 99400 78650 99410 78850
rect 99480 78650 99520 78850
rect 99590 78650 99600 78850
rect 99400 78620 99600 78650
rect 99900 78850 100000 78880
rect 99900 78650 99910 78850
rect 99980 78650 100000 78850
rect 99900 78620 100000 78650
rect 96000 78600 96120 78620
rect 96380 78600 96620 78620
rect 96880 78600 97120 78620
rect 97380 78600 97620 78620
rect 97880 78600 98120 78620
rect 98380 78600 98620 78620
rect 98880 78600 99120 78620
rect 99380 78600 99620 78620
rect 99880 78600 100000 78620
rect 96000 78590 100000 78600
rect 96000 78520 96150 78590
rect 96350 78520 96650 78590
rect 96850 78520 97150 78590
rect 97350 78520 97650 78590
rect 97850 78520 98150 78590
rect 98350 78520 98650 78590
rect 98850 78520 99150 78590
rect 99350 78520 99650 78590
rect 99850 78520 100000 78590
rect 96000 78480 100000 78520
rect 96000 78410 96150 78480
rect 96350 78410 96650 78480
rect 96850 78410 97150 78480
rect 97350 78410 97650 78480
rect 97850 78410 98150 78480
rect 98350 78410 98650 78480
rect 98850 78410 99150 78480
rect 99350 78410 99650 78480
rect 99850 78410 100000 78480
rect 96000 78400 100000 78410
rect 96000 78380 96120 78400
rect 96380 78380 96620 78400
rect 96880 78380 97120 78400
rect 97380 78380 97620 78400
rect 97880 78380 98120 78400
rect 98380 78380 98620 78400
rect 98880 78380 99120 78400
rect 99380 78380 99620 78400
rect 99880 78380 100000 78400
rect 96000 78350 96100 78380
rect 96000 78150 96020 78350
rect 96090 78150 96100 78350
rect 96000 78120 96100 78150
rect 96400 78350 96600 78380
rect 96400 78150 96410 78350
rect 96480 78150 96520 78350
rect 96590 78150 96600 78350
rect 96400 78120 96600 78150
rect 96900 78350 97100 78380
rect 96900 78150 96910 78350
rect 96980 78150 97020 78350
rect 97090 78150 97100 78350
rect 96900 78120 97100 78150
rect 97400 78350 97600 78380
rect 97400 78150 97410 78350
rect 97480 78150 97520 78350
rect 97590 78150 97600 78350
rect 97400 78120 97600 78150
rect 97900 78350 98100 78380
rect 97900 78150 97910 78350
rect 97980 78150 98020 78350
rect 98090 78150 98100 78350
rect 97900 78120 98100 78150
rect 98400 78350 98600 78380
rect 98400 78150 98410 78350
rect 98480 78150 98520 78350
rect 98590 78150 98600 78350
rect 98400 78120 98600 78150
rect 98900 78350 99100 78380
rect 98900 78150 98910 78350
rect 98980 78150 99020 78350
rect 99090 78150 99100 78350
rect 98900 78120 99100 78150
rect 99400 78350 99600 78380
rect 99400 78150 99410 78350
rect 99480 78150 99520 78350
rect 99590 78150 99600 78350
rect 99400 78120 99600 78150
rect 99900 78350 100000 78380
rect 99900 78150 99910 78350
rect 99980 78150 100000 78350
rect 99900 78120 100000 78150
rect 96000 78100 96120 78120
rect 96380 78100 96620 78120
rect 96880 78100 97120 78120
rect 97380 78100 97620 78120
rect 97880 78100 98120 78120
rect 98380 78100 98620 78120
rect 98880 78100 99120 78120
rect 99380 78100 99620 78120
rect 99880 78100 100000 78120
rect 96000 78090 100000 78100
rect 96000 78020 96150 78090
rect 96350 78020 96650 78090
rect 96850 78020 97150 78090
rect 97350 78020 97650 78090
rect 97850 78020 98150 78090
rect 98350 78020 98650 78090
rect 98850 78020 99150 78090
rect 99350 78020 99650 78090
rect 99850 78020 100000 78090
rect 96000 77980 100000 78020
rect 96000 77910 96150 77980
rect 96350 77910 96650 77980
rect 96850 77910 97150 77980
rect 97350 77910 97650 77980
rect 97850 77910 98150 77980
rect 98350 77910 98650 77980
rect 98850 77910 99150 77980
rect 99350 77910 99650 77980
rect 99850 77910 100000 77980
rect 96000 77900 100000 77910
rect 96000 77880 96120 77900
rect 96380 77880 96620 77900
rect 96880 77880 97120 77900
rect 97380 77880 97620 77900
rect 97880 77880 98120 77900
rect 98380 77880 98620 77900
rect 98880 77880 99120 77900
rect 99380 77880 99620 77900
rect 99880 77880 100000 77900
rect 96000 77850 96100 77880
rect 96000 77650 96020 77850
rect 96090 77650 96100 77850
rect 96000 77620 96100 77650
rect 96400 77850 96600 77880
rect 96400 77650 96410 77850
rect 96480 77650 96520 77850
rect 96590 77650 96600 77850
rect 96400 77620 96600 77650
rect 96900 77850 97100 77880
rect 96900 77650 96910 77850
rect 96980 77650 97020 77850
rect 97090 77650 97100 77850
rect 96900 77620 97100 77650
rect 97400 77850 97600 77880
rect 97400 77650 97410 77850
rect 97480 77650 97520 77850
rect 97590 77650 97600 77850
rect 97400 77620 97600 77650
rect 97900 77850 98100 77880
rect 97900 77650 97910 77850
rect 97980 77650 98020 77850
rect 98090 77650 98100 77850
rect 97900 77620 98100 77650
rect 98400 77850 98600 77880
rect 98400 77650 98410 77850
rect 98480 77650 98520 77850
rect 98590 77650 98600 77850
rect 98400 77620 98600 77650
rect 98900 77850 99100 77880
rect 98900 77650 98910 77850
rect 98980 77650 99020 77850
rect 99090 77650 99100 77850
rect 98900 77620 99100 77650
rect 99400 77850 99600 77880
rect 99400 77650 99410 77850
rect 99480 77650 99520 77850
rect 99590 77650 99600 77850
rect 99400 77620 99600 77650
rect 99900 77850 100000 77880
rect 99900 77650 99910 77850
rect 99980 77650 100000 77850
rect 99900 77620 100000 77650
rect 96000 77600 96120 77620
rect 96380 77600 96620 77620
rect 96880 77600 97120 77620
rect 97380 77600 97620 77620
rect 97880 77600 98120 77620
rect 98380 77600 98620 77620
rect 98880 77600 99120 77620
rect 99380 77600 99620 77620
rect 99880 77600 100000 77620
rect 96000 77590 100000 77600
rect 96000 77520 96150 77590
rect 96350 77520 96650 77590
rect 96850 77520 97150 77590
rect 97350 77520 97650 77590
rect 97850 77520 98150 77590
rect 98350 77520 98650 77590
rect 98850 77520 99150 77590
rect 99350 77520 99650 77590
rect 99850 77520 100000 77590
rect 96000 77480 100000 77520
rect 96000 77410 96150 77480
rect 96350 77410 96650 77480
rect 96850 77410 97150 77480
rect 97350 77410 97650 77480
rect 97850 77410 98150 77480
rect 98350 77410 98650 77480
rect 98850 77410 99150 77480
rect 99350 77410 99650 77480
rect 99850 77410 100000 77480
rect 96000 77400 100000 77410
rect 96000 77380 96120 77400
rect 96380 77380 96620 77400
rect 96880 77380 97120 77400
rect 97380 77380 97620 77400
rect 97880 77380 98120 77400
rect 98380 77380 98620 77400
rect 98880 77380 99120 77400
rect 99380 77380 99620 77400
rect 99880 77380 100000 77400
rect 96000 77350 96100 77380
rect 96000 77150 96020 77350
rect 96090 77150 96100 77350
rect 96000 77120 96100 77150
rect 96400 77350 96600 77380
rect 96400 77150 96410 77350
rect 96480 77150 96520 77350
rect 96590 77150 96600 77350
rect 96400 77120 96600 77150
rect 96900 77350 97100 77380
rect 96900 77150 96910 77350
rect 96980 77150 97020 77350
rect 97090 77150 97100 77350
rect 96900 77120 97100 77150
rect 97400 77350 97600 77380
rect 97400 77150 97410 77350
rect 97480 77150 97520 77350
rect 97590 77150 97600 77350
rect 97400 77120 97600 77150
rect 97900 77350 98100 77380
rect 97900 77150 97910 77350
rect 97980 77150 98020 77350
rect 98090 77150 98100 77350
rect 97900 77120 98100 77150
rect 98400 77350 98600 77380
rect 98400 77150 98410 77350
rect 98480 77150 98520 77350
rect 98590 77150 98600 77350
rect 98400 77120 98600 77150
rect 98900 77350 99100 77380
rect 98900 77150 98910 77350
rect 98980 77150 99020 77350
rect 99090 77150 99100 77350
rect 98900 77120 99100 77150
rect 99400 77350 99600 77380
rect 99400 77150 99410 77350
rect 99480 77150 99520 77350
rect 99590 77150 99600 77350
rect 99400 77120 99600 77150
rect 99900 77350 100000 77380
rect 99900 77150 99910 77350
rect 99980 77150 100000 77350
rect 99900 77120 100000 77150
rect 96000 77100 96120 77120
rect 96380 77100 96620 77120
rect 96880 77100 97120 77120
rect 97380 77100 97620 77120
rect 97880 77100 98120 77120
rect 98380 77100 98620 77120
rect 98880 77100 99120 77120
rect 99380 77100 99620 77120
rect 99880 77100 100000 77120
rect 96000 77090 100000 77100
rect 96000 77020 96150 77090
rect 96350 77020 96650 77090
rect 96850 77020 97150 77090
rect 97350 77020 97650 77090
rect 97850 77020 98150 77090
rect 98350 77020 98650 77090
rect 98850 77020 99150 77090
rect 99350 77020 99650 77090
rect 99850 77020 100000 77090
rect 96000 76980 100000 77020
rect 96000 76910 96150 76980
rect 96350 76910 96650 76980
rect 96850 76910 97150 76980
rect 97350 76910 97650 76980
rect 97850 76910 98150 76980
rect 98350 76910 98650 76980
rect 98850 76910 99150 76980
rect 99350 76910 99650 76980
rect 99850 76910 100000 76980
rect 96000 76900 100000 76910
rect 96000 76880 96120 76900
rect 96380 76880 96620 76900
rect 96880 76880 97120 76900
rect 97380 76880 97620 76900
rect 97880 76880 98120 76900
rect 98380 76880 98620 76900
rect 98880 76880 99120 76900
rect 99380 76880 99620 76900
rect 99880 76880 100000 76900
rect 96000 76850 96100 76880
rect 96000 76650 96020 76850
rect 96090 76650 96100 76850
rect 96000 76620 96100 76650
rect 96400 76850 96600 76880
rect 96400 76650 96410 76850
rect 96480 76650 96520 76850
rect 96590 76650 96600 76850
rect 96400 76620 96600 76650
rect 96900 76850 97100 76880
rect 96900 76650 96910 76850
rect 96980 76650 97020 76850
rect 97090 76650 97100 76850
rect 96900 76620 97100 76650
rect 97400 76850 97600 76880
rect 97400 76650 97410 76850
rect 97480 76650 97520 76850
rect 97590 76650 97600 76850
rect 97400 76620 97600 76650
rect 97900 76850 98100 76880
rect 97900 76650 97910 76850
rect 97980 76650 98020 76850
rect 98090 76650 98100 76850
rect 97900 76620 98100 76650
rect 98400 76850 98600 76880
rect 98400 76650 98410 76850
rect 98480 76650 98520 76850
rect 98590 76650 98600 76850
rect 98400 76620 98600 76650
rect 98900 76850 99100 76880
rect 98900 76650 98910 76850
rect 98980 76650 99020 76850
rect 99090 76650 99100 76850
rect 98900 76620 99100 76650
rect 99400 76850 99600 76880
rect 99400 76650 99410 76850
rect 99480 76650 99520 76850
rect 99590 76650 99600 76850
rect 99400 76620 99600 76650
rect 99900 76850 100000 76880
rect 99900 76650 99910 76850
rect 99980 76650 100000 76850
rect 99900 76620 100000 76650
rect 96000 76600 96120 76620
rect 96380 76600 96620 76620
rect 96880 76600 97120 76620
rect 97380 76600 97620 76620
rect 97880 76600 98120 76620
rect 98380 76600 98620 76620
rect 98880 76600 99120 76620
rect 99380 76600 99620 76620
rect 99880 76600 100000 76620
rect 96000 76590 100000 76600
rect 96000 76520 96150 76590
rect 96350 76520 96650 76590
rect 96850 76520 97150 76590
rect 97350 76520 97650 76590
rect 97850 76520 98150 76590
rect 98350 76520 98650 76590
rect 98850 76520 99150 76590
rect 99350 76520 99650 76590
rect 99850 76520 100000 76590
rect 96000 76480 100000 76520
rect 96000 76410 96150 76480
rect 96350 76410 96650 76480
rect 96850 76410 97150 76480
rect 97350 76410 97650 76480
rect 97850 76410 98150 76480
rect 98350 76410 98650 76480
rect 98850 76410 99150 76480
rect 99350 76410 99650 76480
rect 99850 76410 100000 76480
rect 96000 76400 100000 76410
rect 96000 76380 96120 76400
rect 96380 76380 96620 76400
rect 96880 76380 97120 76400
rect 97380 76380 97620 76400
rect 97880 76380 98120 76400
rect 98380 76380 98620 76400
rect 98880 76380 99120 76400
rect 99380 76380 99620 76400
rect 99880 76380 100000 76400
rect 96000 76350 96100 76380
rect 96000 76150 96020 76350
rect 96090 76150 96100 76350
rect 96000 76120 96100 76150
rect 96400 76350 96600 76380
rect 96400 76150 96410 76350
rect 96480 76150 96520 76350
rect 96590 76150 96600 76350
rect 96400 76120 96600 76150
rect 96900 76350 97100 76380
rect 96900 76150 96910 76350
rect 96980 76150 97020 76350
rect 97090 76150 97100 76350
rect 96900 76120 97100 76150
rect 97400 76350 97600 76380
rect 97400 76150 97410 76350
rect 97480 76150 97520 76350
rect 97590 76150 97600 76350
rect 97400 76120 97600 76150
rect 97900 76350 98100 76380
rect 97900 76150 97910 76350
rect 97980 76150 98020 76350
rect 98090 76150 98100 76350
rect 97900 76120 98100 76150
rect 98400 76350 98600 76380
rect 98400 76150 98410 76350
rect 98480 76150 98520 76350
rect 98590 76150 98600 76350
rect 98400 76120 98600 76150
rect 98900 76350 99100 76380
rect 98900 76150 98910 76350
rect 98980 76150 99020 76350
rect 99090 76150 99100 76350
rect 98900 76120 99100 76150
rect 99400 76350 99600 76380
rect 99400 76150 99410 76350
rect 99480 76150 99520 76350
rect 99590 76150 99600 76350
rect 99400 76120 99600 76150
rect 99900 76350 100000 76380
rect 99900 76150 99910 76350
rect 99980 76150 100000 76350
rect 99900 76120 100000 76150
rect 96000 76100 96120 76120
rect 96380 76100 96620 76120
rect 96880 76100 97120 76120
rect 97380 76100 97620 76120
rect 97880 76100 98120 76120
rect 98380 76100 98620 76120
rect 98880 76100 99120 76120
rect 99380 76100 99620 76120
rect 99880 76100 100000 76120
rect 96000 76090 100000 76100
rect 96000 76020 96150 76090
rect 96350 76020 96650 76090
rect 96850 76020 97150 76090
rect 97350 76020 97650 76090
rect 97850 76020 98150 76090
rect 98350 76020 98650 76090
rect 98850 76020 99150 76090
rect 99350 76020 99650 76090
rect 99850 76020 100000 76090
rect 96000 75980 100000 76020
rect 96000 75910 96150 75980
rect 96350 75910 96650 75980
rect 96850 75910 97150 75980
rect 97350 75910 97650 75980
rect 97850 75910 98150 75980
rect 98350 75910 98650 75980
rect 98850 75910 99150 75980
rect 99350 75910 99650 75980
rect 99850 75910 100000 75980
rect 96000 75900 100000 75910
rect 96000 75880 96120 75900
rect 96380 75880 96620 75900
rect 96880 75880 97120 75900
rect 97380 75880 97620 75900
rect 97880 75880 98120 75900
rect 98380 75880 98620 75900
rect 98880 75880 99120 75900
rect 99380 75880 99620 75900
rect 99880 75880 100000 75900
rect 96000 75850 96100 75880
rect 96000 75650 96020 75850
rect 96090 75650 96100 75850
rect 96000 75620 96100 75650
rect 96400 75850 96600 75880
rect 96400 75650 96410 75850
rect 96480 75650 96520 75850
rect 96590 75650 96600 75850
rect 96400 75620 96600 75650
rect 96900 75850 97100 75880
rect 96900 75650 96910 75850
rect 96980 75650 97020 75850
rect 97090 75650 97100 75850
rect 96900 75620 97100 75650
rect 97400 75850 97600 75880
rect 97400 75650 97410 75850
rect 97480 75650 97520 75850
rect 97590 75650 97600 75850
rect 97400 75620 97600 75650
rect 97900 75850 98100 75880
rect 97900 75650 97910 75850
rect 97980 75650 98020 75850
rect 98090 75650 98100 75850
rect 97900 75620 98100 75650
rect 98400 75850 98600 75880
rect 98400 75650 98410 75850
rect 98480 75650 98520 75850
rect 98590 75650 98600 75850
rect 98400 75620 98600 75650
rect 98900 75850 99100 75880
rect 98900 75650 98910 75850
rect 98980 75650 99020 75850
rect 99090 75650 99100 75850
rect 98900 75620 99100 75650
rect 99400 75850 99600 75880
rect 99400 75650 99410 75850
rect 99480 75650 99520 75850
rect 99590 75650 99600 75850
rect 99400 75620 99600 75650
rect 99900 75850 100000 75880
rect 99900 75650 99910 75850
rect 99980 75650 100000 75850
rect 99900 75620 100000 75650
rect 96000 75600 96120 75620
rect 96380 75600 96620 75620
rect 96880 75600 97120 75620
rect 97380 75600 97620 75620
rect 97880 75600 98120 75620
rect 98380 75600 98620 75620
rect 98880 75600 99120 75620
rect 99380 75600 99620 75620
rect 99880 75600 100000 75620
rect 96000 75590 100000 75600
rect 96000 75520 96150 75590
rect 96350 75520 96650 75590
rect 96850 75520 97150 75590
rect 97350 75520 97650 75590
rect 97850 75520 98150 75590
rect 98350 75520 98650 75590
rect 98850 75520 99150 75590
rect 99350 75520 99650 75590
rect 99850 75520 100000 75590
rect 96000 75480 100000 75520
rect 96000 75410 96150 75480
rect 96350 75410 96650 75480
rect 96850 75410 97150 75480
rect 97350 75410 97650 75480
rect 97850 75410 98150 75480
rect 98350 75410 98650 75480
rect 98850 75410 99150 75480
rect 99350 75410 99650 75480
rect 99850 75410 100000 75480
rect 96000 75400 100000 75410
rect 96000 75380 96120 75400
rect 96380 75380 96620 75400
rect 96880 75380 97120 75400
rect 97380 75380 97620 75400
rect 97880 75380 98120 75400
rect 98380 75380 98620 75400
rect 98880 75380 99120 75400
rect 99380 75380 99620 75400
rect 99880 75380 100000 75400
rect 96000 75350 96100 75380
rect 96000 75150 96020 75350
rect 96090 75150 96100 75350
rect 96000 75120 96100 75150
rect 96400 75350 96600 75380
rect 96400 75150 96410 75350
rect 96480 75150 96520 75350
rect 96590 75150 96600 75350
rect 96400 75120 96600 75150
rect 96900 75350 97100 75380
rect 96900 75150 96910 75350
rect 96980 75150 97020 75350
rect 97090 75150 97100 75350
rect 96900 75120 97100 75150
rect 97400 75350 97600 75380
rect 97400 75150 97410 75350
rect 97480 75150 97520 75350
rect 97590 75150 97600 75350
rect 97400 75120 97600 75150
rect 97900 75350 98100 75380
rect 97900 75150 97910 75350
rect 97980 75150 98020 75350
rect 98090 75150 98100 75350
rect 97900 75120 98100 75150
rect 98400 75350 98600 75380
rect 98400 75150 98410 75350
rect 98480 75150 98520 75350
rect 98590 75150 98600 75350
rect 98400 75120 98600 75150
rect 98900 75350 99100 75380
rect 98900 75150 98910 75350
rect 98980 75150 99020 75350
rect 99090 75150 99100 75350
rect 98900 75120 99100 75150
rect 99400 75350 99600 75380
rect 99400 75150 99410 75350
rect 99480 75150 99520 75350
rect 99590 75150 99600 75350
rect 99400 75120 99600 75150
rect 99900 75350 100000 75380
rect 99900 75150 99910 75350
rect 99980 75150 100000 75350
rect 99900 75120 100000 75150
rect 96000 75100 96120 75120
rect 96380 75100 96620 75120
rect 96880 75100 97120 75120
rect 97380 75100 97620 75120
rect 97880 75100 98120 75120
rect 98380 75100 98620 75120
rect 98880 75100 99120 75120
rect 99380 75100 99620 75120
rect 99880 75100 100000 75120
rect 96000 75090 100000 75100
rect 96000 75020 96150 75090
rect 96350 75020 96650 75090
rect 96850 75020 97150 75090
rect 97350 75020 97650 75090
rect 97850 75020 98150 75090
rect 98350 75020 98650 75090
rect 98850 75020 99150 75090
rect 99350 75020 99650 75090
rect 99850 75020 100000 75090
rect 96000 74980 100000 75020
rect 96000 74910 96150 74980
rect 96350 74910 96650 74980
rect 96850 74910 97150 74980
rect 97350 74910 97650 74980
rect 97850 74910 98150 74980
rect 98350 74910 98650 74980
rect 98850 74910 99150 74980
rect 99350 74910 99650 74980
rect 99850 74910 100000 74980
rect 96000 74900 100000 74910
rect 96000 74880 96120 74900
rect 96380 74880 96620 74900
rect 96880 74880 97120 74900
rect 97380 74880 97620 74900
rect 97880 74880 98120 74900
rect 98380 74880 98620 74900
rect 98880 74880 99120 74900
rect 99380 74880 99620 74900
rect 99880 74880 100000 74900
rect 96000 74850 96100 74880
rect 96000 74650 96020 74850
rect 96090 74650 96100 74850
rect 96000 74620 96100 74650
rect 96400 74850 96600 74880
rect 96400 74650 96410 74850
rect 96480 74650 96520 74850
rect 96590 74650 96600 74850
rect 96400 74620 96600 74650
rect 96900 74850 97100 74880
rect 96900 74650 96910 74850
rect 96980 74650 97020 74850
rect 97090 74650 97100 74850
rect 96900 74620 97100 74650
rect 97400 74850 97600 74880
rect 97400 74650 97410 74850
rect 97480 74650 97520 74850
rect 97590 74650 97600 74850
rect 97400 74620 97600 74650
rect 97900 74850 98100 74880
rect 97900 74650 97910 74850
rect 97980 74650 98020 74850
rect 98090 74650 98100 74850
rect 97900 74620 98100 74650
rect 98400 74850 98600 74880
rect 98400 74650 98410 74850
rect 98480 74650 98520 74850
rect 98590 74650 98600 74850
rect 98400 74620 98600 74650
rect 98900 74850 99100 74880
rect 98900 74650 98910 74850
rect 98980 74650 99020 74850
rect 99090 74650 99100 74850
rect 98900 74620 99100 74650
rect 99400 74850 99600 74880
rect 99400 74650 99410 74850
rect 99480 74650 99520 74850
rect 99590 74650 99600 74850
rect 99400 74620 99600 74650
rect 99900 74850 100000 74880
rect 99900 74650 99910 74850
rect 99980 74650 100000 74850
rect 99900 74620 100000 74650
rect 96000 74600 96120 74620
rect 96380 74600 96620 74620
rect 96880 74600 97120 74620
rect 97380 74600 97620 74620
rect 97880 74600 98120 74620
rect 98380 74600 98620 74620
rect 98880 74600 99120 74620
rect 99380 74600 99620 74620
rect 99880 74600 100000 74620
rect 96000 74590 100000 74600
rect 96000 74520 96150 74590
rect 96350 74520 96650 74590
rect 96850 74520 97150 74590
rect 97350 74520 97650 74590
rect 97850 74520 98150 74590
rect 98350 74520 98650 74590
rect 98850 74520 99150 74590
rect 99350 74520 99650 74590
rect 99850 74520 100000 74590
rect 96000 74480 100000 74520
rect 96000 74410 96150 74480
rect 96350 74410 96650 74480
rect 96850 74410 97150 74480
rect 97350 74410 97650 74480
rect 97850 74410 98150 74480
rect 98350 74410 98650 74480
rect 98850 74410 99150 74480
rect 99350 74410 99650 74480
rect 99850 74410 100000 74480
rect 96000 74400 100000 74410
rect 96000 74380 96120 74400
rect 96380 74380 96620 74400
rect 96880 74380 97120 74400
rect 97380 74380 97620 74400
rect 97880 74380 98120 74400
rect 98380 74380 98620 74400
rect 98880 74380 99120 74400
rect 99380 74380 99620 74400
rect 99880 74380 100000 74400
rect 96000 74350 96100 74380
rect 96000 74150 96020 74350
rect 96090 74150 96100 74350
rect 96000 74120 96100 74150
rect 96400 74350 96600 74380
rect 96400 74150 96410 74350
rect 96480 74150 96520 74350
rect 96590 74150 96600 74350
rect 96400 74120 96600 74150
rect 96900 74350 97100 74380
rect 96900 74150 96910 74350
rect 96980 74150 97020 74350
rect 97090 74150 97100 74350
rect 96900 74120 97100 74150
rect 97400 74350 97600 74380
rect 97400 74150 97410 74350
rect 97480 74150 97520 74350
rect 97590 74150 97600 74350
rect 97400 74120 97600 74150
rect 97900 74350 98100 74380
rect 97900 74150 97910 74350
rect 97980 74150 98020 74350
rect 98090 74150 98100 74350
rect 97900 74120 98100 74150
rect 98400 74350 98600 74380
rect 98400 74150 98410 74350
rect 98480 74150 98520 74350
rect 98590 74150 98600 74350
rect 98400 74120 98600 74150
rect 98900 74350 99100 74380
rect 98900 74150 98910 74350
rect 98980 74150 99020 74350
rect 99090 74150 99100 74350
rect 98900 74120 99100 74150
rect 99400 74350 99600 74380
rect 99400 74150 99410 74350
rect 99480 74150 99520 74350
rect 99590 74150 99600 74350
rect 99400 74120 99600 74150
rect 99900 74350 100000 74380
rect 99900 74150 99910 74350
rect 99980 74150 100000 74350
rect 99900 74120 100000 74150
rect 96000 74100 96120 74120
rect 96380 74100 96620 74120
rect 96880 74100 97120 74120
rect 97380 74100 97620 74120
rect 97880 74100 98120 74120
rect 98380 74100 98620 74120
rect 98880 74100 99120 74120
rect 99380 74100 99620 74120
rect 99880 74100 100000 74120
rect 96000 74090 100000 74100
rect 96000 74020 96150 74090
rect 96350 74020 96650 74090
rect 96850 74020 97150 74090
rect 97350 74020 97650 74090
rect 97850 74020 98150 74090
rect 98350 74020 98650 74090
rect 98850 74020 99150 74090
rect 99350 74020 99650 74090
rect 99850 74020 100000 74090
rect 96000 73980 100000 74020
rect 96000 73910 96150 73980
rect 96350 73910 96650 73980
rect 96850 73910 97150 73980
rect 97350 73910 97650 73980
rect 97850 73910 98150 73980
rect 98350 73910 98650 73980
rect 98850 73910 99150 73980
rect 99350 73910 99650 73980
rect 99850 73910 100000 73980
rect 96000 73900 100000 73910
rect 96000 73880 96120 73900
rect 96380 73880 96620 73900
rect 96880 73880 97120 73900
rect 97380 73880 97620 73900
rect 97880 73880 98120 73900
rect 98380 73880 98620 73900
rect 98880 73880 99120 73900
rect 99380 73880 99620 73900
rect 99880 73880 100000 73900
rect 96000 73850 96100 73880
rect 96000 73650 96020 73850
rect 96090 73650 96100 73850
rect 96000 73620 96100 73650
rect 96400 73850 96600 73880
rect 96400 73650 96410 73850
rect 96480 73650 96520 73850
rect 96590 73650 96600 73850
rect 96400 73620 96600 73650
rect 96900 73850 97100 73880
rect 96900 73650 96910 73850
rect 96980 73650 97020 73850
rect 97090 73650 97100 73850
rect 96900 73620 97100 73650
rect 97400 73850 97600 73880
rect 97400 73650 97410 73850
rect 97480 73650 97520 73850
rect 97590 73650 97600 73850
rect 97400 73620 97600 73650
rect 97900 73850 98100 73880
rect 97900 73650 97910 73850
rect 97980 73650 98020 73850
rect 98090 73650 98100 73850
rect 97900 73620 98100 73650
rect 98400 73850 98600 73880
rect 98400 73650 98410 73850
rect 98480 73650 98520 73850
rect 98590 73650 98600 73850
rect 98400 73620 98600 73650
rect 98900 73850 99100 73880
rect 98900 73650 98910 73850
rect 98980 73650 99020 73850
rect 99090 73650 99100 73850
rect 98900 73620 99100 73650
rect 99400 73850 99600 73880
rect 99400 73650 99410 73850
rect 99480 73650 99520 73850
rect 99590 73650 99600 73850
rect 99400 73620 99600 73650
rect 99900 73850 100000 73880
rect 99900 73650 99910 73850
rect 99980 73650 100000 73850
rect 99900 73620 100000 73650
rect 96000 73600 96120 73620
rect 96380 73600 96620 73620
rect 96880 73600 97120 73620
rect 97380 73600 97620 73620
rect 97880 73600 98120 73620
rect 98380 73600 98620 73620
rect 98880 73600 99120 73620
rect 99380 73600 99620 73620
rect 99880 73600 100000 73620
rect 96000 73590 100000 73600
rect 96000 73520 96150 73590
rect 96350 73520 96650 73590
rect 96850 73520 97150 73590
rect 97350 73520 97650 73590
rect 97850 73520 98150 73590
rect 98350 73520 98650 73590
rect 98850 73520 99150 73590
rect 99350 73520 99650 73590
rect 99850 73520 100000 73590
rect 96000 73480 100000 73520
rect 96000 73410 96150 73480
rect 96350 73410 96650 73480
rect 96850 73410 97150 73480
rect 97350 73410 97650 73480
rect 97850 73410 98150 73480
rect 98350 73410 98650 73480
rect 98850 73410 99150 73480
rect 99350 73410 99650 73480
rect 99850 73410 100000 73480
rect 96000 73400 100000 73410
rect 96000 73380 96120 73400
rect 96380 73380 96620 73400
rect 96880 73380 97120 73400
rect 97380 73380 97620 73400
rect 97880 73380 98120 73400
rect 98380 73380 98620 73400
rect 98880 73380 99120 73400
rect 99380 73380 99620 73400
rect 99880 73380 100000 73400
rect 96000 73350 96100 73380
rect 96000 73150 96020 73350
rect 96090 73150 96100 73350
rect 96000 73120 96100 73150
rect 96400 73350 96600 73380
rect 96400 73150 96410 73350
rect 96480 73150 96520 73350
rect 96590 73150 96600 73350
rect 96400 73120 96600 73150
rect 96900 73350 97100 73380
rect 96900 73150 96910 73350
rect 96980 73150 97020 73350
rect 97090 73150 97100 73350
rect 96900 73120 97100 73150
rect 97400 73350 97600 73380
rect 97400 73150 97410 73350
rect 97480 73150 97520 73350
rect 97590 73150 97600 73350
rect 97400 73120 97600 73150
rect 97900 73350 98100 73380
rect 97900 73150 97910 73350
rect 97980 73150 98020 73350
rect 98090 73150 98100 73350
rect 97900 73120 98100 73150
rect 98400 73350 98600 73380
rect 98400 73150 98410 73350
rect 98480 73150 98520 73350
rect 98590 73150 98600 73350
rect 98400 73120 98600 73150
rect 98900 73350 99100 73380
rect 98900 73150 98910 73350
rect 98980 73150 99020 73350
rect 99090 73150 99100 73350
rect 98900 73120 99100 73150
rect 99400 73350 99600 73380
rect 99400 73150 99410 73350
rect 99480 73150 99520 73350
rect 99590 73150 99600 73350
rect 99400 73120 99600 73150
rect 99900 73350 100000 73380
rect 99900 73150 99910 73350
rect 99980 73150 100000 73350
rect 99900 73120 100000 73150
rect 96000 73100 96120 73120
rect 96380 73100 96620 73120
rect 96880 73100 97120 73120
rect 97380 73100 97620 73120
rect 97880 73100 98120 73120
rect 98380 73100 98620 73120
rect 98880 73100 99120 73120
rect 99380 73100 99620 73120
rect 99880 73100 100000 73120
rect 96000 73090 100000 73100
rect 96000 73020 96150 73090
rect 96350 73020 96650 73090
rect 96850 73020 97150 73090
rect 97350 73020 97650 73090
rect 97850 73020 98150 73090
rect 98350 73020 98650 73090
rect 98850 73020 99150 73090
rect 99350 73020 99650 73090
rect 99850 73020 100000 73090
rect 96000 72980 100000 73020
rect 96000 72910 96150 72980
rect 96350 72910 96650 72980
rect 96850 72910 97150 72980
rect 97350 72910 97650 72980
rect 97850 72910 98150 72980
rect 98350 72910 98650 72980
rect 98850 72910 99150 72980
rect 99350 72910 99650 72980
rect 99850 72910 100000 72980
rect 96000 72900 100000 72910
rect 96000 72880 96120 72900
rect 96380 72880 96620 72900
rect 96880 72880 97120 72900
rect 97380 72880 97620 72900
rect 97880 72880 98120 72900
rect 98380 72880 98620 72900
rect 98880 72880 99120 72900
rect 99380 72880 99620 72900
rect 99880 72880 100000 72900
rect 96000 72850 96100 72880
rect 96000 72650 96020 72850
rect 96090 72650 96100 72850
rect 96000 72620 96100 72650
rect 96400 72850 96600 72880
rect 96400 72650 96410 72850
rect 96480 72650 96520 72850
rect 96590 72650 96600 72850
rect 96400 72620 96600 72650
rect 96900 72850 97100 72880
rect 96900 72650 96910 72850
rect 96980 72650 97020 72850
rect 97090 72650 97100 72850
rect 96900 72620 97100 72650
rect 97400 72850 97600 72880
rect 97400 72650 97410 72850
rect 97480 72650 97520 72850
rect 97590 72650 97600 72850
rect 97400 72620 97600 72650
rect 97900 72850 98100 72880
rect 97900 72650 97910 72850
rect 97980 72650 98020 72850
rect 98090 72650 98100 72850
rect 97900 72620 98100 72650
rect 98400 72850 98600 72880
rect 98400 72650 98410 72850
rect 98480 72650 98520 72850
rect 98590 72650 98600 72850
rect 98400 72620 98600 72650
rect 98900 72850 99100 72880
rect 98900 72650 98910 72850
rect 98980 72650 99020 72850
rect 99090 72650 99100 72850
rect 98900 72620 99100 72650
rect 99400 72850 99600 72880
rect 99400 72650 99410 72850
rect 99480 72650 99520 72850
rect 99590 72650 99600 72850
rect 99400 72620 99600 72650
rect 99900 72850 100000 72880
rect 99900 72650 99910 72850
rect 99980 72650 100000 72850
rect 99900 72620 100000 72650
rect 96000 72600 96120 72620
rect 96380 72600 96620 72620
rect 96880 72600 97120 72620
rect 97380 72600 97620 72620
rect 97880 72600 98120 72620
rect 98380 72600 98620 72620
rect 98880 72600 99120 72620
rect 99380 72600 99620 72620
rect 99880 72600 100000 72620
rect 96000 72590 100000 72600
rect 96000 72520 96150 72590
rect 96350 72520 96650 72590
rect 96850 72520 97150 72590
rect 97350 72520 97650 72590
rect 97850 72520 98150 72590
rect 98350 72520 98650 72590
rect 98850 72520 99150 72590
rect 99350 72520 99650 72590
rect 99850 72520 100000 72590
rect 96000 72480 100000 72520
rect 96000 72410 96150 72480
rect 96350 72410 96650 72480
rect 96850 72410 97150 72480
rect 97350 72410 97650 72480
rect 97850 72410 98150 72480
rect 98350 72410 98650 72480
rect 98850 72410 99150 72480
rect 99350 72410 99650 72480
rect 99850 72410 100000 72480
rect 96000 72400 100000 72410
rect 96000 72380 96120 72400
rect 96380 72380 96620 72400
rect 96880 72380 97120 72400
rect 97380 72380 97620 72400
rect 97880 72380 98120 72400
rect 98380 72380 98620 72400
rect 98880 72380 99120 72400
rect 99380 72380 99620 72400
rect 99880 72380 100000 72400
rect 96000 72350 96100 72380
rect 96000 72150 96020 72350
rect 96090 72150 96100 72350
rect 96000 72120 96100 72150
rect 96400 72350 96600 72380
rect 96400 72150 96410 72350
rect 96480 72150 96520 72350
rect 96590 72150 96600 72350
rect 96400 72120 96600 72150
rect 96900 72350 97100 72380
rect 96900 72150 96910 72350
rect 96980 72150 97020 72350
rect 97090 72150 97100 72350
rect 96900 72120 97100 72150
rect 97400 72350 97600 72380
rect 97400 72150 97410 72350
rect 97480 72150 97520 72350
rect 97590 72150 97600 72350
rect 97400 72120 97600 72150
rect 97900 72350 98100 72380
rect 97900 72150 97910 72350
rect 97980 72150 98020 72350
rect 98090 72150 98100 72350
rect 97900 72120 98100 72150
rect 98400 72350 98600 72380
rect 98400 72150 98410 72350
rect 98480 72150 98520 72350
rect 98590 72150 98600 72350
rect 98400 72120 98600 72150
rect 98900 72350 99100 72380
rect 98900 72150 98910 72350
rect 98980 72150 99020 72350
rect 99090 72150 99100 72350
rect 98900 72120 99100 72150
rect 99400 72350 99600 72380
rect 99400 72150 99410 72350
rect 99480 72150 99520 72350
rect 99590 72150 99600 72350
rect 99400 72120 99600 72150
rect 99900 72350 100000 72380
rect 99900 72150 99910 72350
rect 99980 72150 100000 72350
rect 99900 72120 100000 72150
rect 96000 72100 96120 72120
rect 96380 72100 96620 72120
rect 96880 72100 97120 72120
rect 97380 72100 97620 72120
rect 97880 72100 98120 72120
rect 98380 72100 98620 72120
rect 98880 72100 99120 72120
rect 99380 72100 99620 72120
rect 99880 72100 100000 72120
rect 96000 72090 100000 72100
rect 96000 72020 96150 72090
rect 96350 72020 96650 72090
rect 96850 72020 97150 72090
rect 97350 72020 97650 72090
rect 97850 72020 98150 72090
rect 98350 72020 98650 72090
rect 98850 72020 99150 72090
rect 99350 72020 99650 72090
rect 99850 72020 100000 72090
rect 96000 71980 100000 72020
rect 96000 71910 96150 71980
rect 96350 71910 96650 71980
rect 96850 71910 97150 71980
rect 97350 71910 97650 71980
rect 97850 71910 98150 71980
rect 98350 71910 98650 71980
rect 98850 71910 99150 71980
rect 99350 71910 99650 71980
rect 99850 71910 100000 71980
rect 96000 71900 100000 71910
rect 96000 71880 96120 71900
rect 96380 71880 96620 71900
rect 96880 71880 97120 71900
rect 97380 71880 97620 71900
rect 97880 71880 98120 71900
rect 98380 71880 98620 71900
rect 98880 71880 99120 71900
rect 99380 71880 99620 71900
rect 99880 71880 100000 71900
rect 96000 71850 96100 71880
rect 96000 71650 96020 71850
rect 96090 71650 96100 71850
rect 96000 71620 96100 71650
rect 96400 71850 96600 71880
rect 96400 71650 96410 71850
rect 96480 71650 96520 71850
rect 96590 71650 96600 71850
rect 96400 71620 96600 71650
rect 96900 71850 97100 71880
rect 96900 71650 96910 71850
rect 96980 71650 97020 71850
rect 97090 71650 97100 71850
rect 96900 71620 97100 71650
rect 97400 71850 97600 71880
rect 97400 71650 97410 71850
rect 97480 71650 97520 71850
rect 97590 71650 97600 71850
rect 97400 71620 97600 71650
rect 97900 71850 98100 71880
rect 97900 71650 97910 71850
rect 97980 71650 98020 71850
rect 98090 71650 98100 71850
rect 97900 71620 98100 71650
rect 98400 71850 98600 71880
rect 98400 71650 98410 71850
rect 98480 71650 98520 71850
rect 98590 71650 98600 71850
rect 98400 71620 98600 71650
rect 98900 71850 99100 71880
rect 98900 71650 98910 71850
rect 98980 71650 99020 71850
rect 99090 71650 99100 71850
rect 98900 71620 99100 71650
rect 99400 71850 99600 71880
rect 99400 71650 99410 71850
rect 99480 71650 99520 71850
rect 99590 71650 99600 71850
rect 99400 71620 99600 71650
rect 99900 71850 100000 71880
rect 99900 71650 99910 71850
rect 99980 71650 100000 71850
rect 99900 71620 100000 71650
rect 96000 71600 96120 71620
rect 96380 71600 96620 71620
rect 96880 71600 97120 71620
rect 97380 71600 97620 71620
rect 97880 71600 98120 71620
rect 98380 71600 98620 71620
rect 98880 71600 99120 71620
rect 99380 71600 99620 71620
rect 99880 71600 100000 71620
rect 96000 71590 100000 71600
rect 96000 71520 96150 71590
rect 96350 71520 96650 71590
rect 96850 71520 97150 71590
rect 97350 71520 97650 71590
rect 97850 71520 98150 71590
rect 98350 71520 98650 71590
rect 98850 71520 99150 71590
rect 99350 71520 99650 71590
rect 99850 71520 100000 71590
rect 96000 71480 100000 71520
rect 96000 71410 96150 71480
rect 96350 71410 96650 71480
rect 96850 71410 97150 71480
rect 97350 71410 97650 71480
rect 97850 71410 98150 71480
rect 98350 71410 98650 71480
rect 98850 71410 99150 71480
rect 99350 71410 99650 71480
rect 99850 71410 100000 71480
rect 96000 71400 100000 71410
rect 96000 71380 96120 71400
rect 96380 71380 96620 71400
rect 96880 71380 97120 71400
rect 97380 71380 97620 71400
rect 97880 71380 98120 71400
rect 98380 71380 98620 71400
rect 98880 71380 99120 71400
rect 99380 71380 99620 71400
rect 99880 71380 100000 71400
rect 96000 71350 96100 71380
rect 96000 71150 96020 71350
rect 96090 71150 96100 71350
rect 96000 71120 96100 71150
rect 96400 71350 96600 71380
rect 96400 71150 96410 71350
rect 96480 71150 96520 71350
rect 96590 71150 96600 71350
rect 96400 71120 96600 71150
rect 96900 71350 97100 71380
rect 96900 71150 96910 71350
rect 96980 71150 97020 71350
rect 97090 71150 97100 71350
rect 96900 71120 97100 71150
rect 97400 71350 97600 71380
rect 97400 71150 97410 71350
rect 97480 71150 97520 71350
rect 97590 71150 97600 71350
rect 97400 71120 97600 71150
rect 97900 71350 98100 71380
rect 97900 71150 97910 71350
rect 97980 71150 98020 71350
rect 98090 71150 98100 71350
rect 97900 71120 98100 71150
rect 98400 71350 98600 71380
rect 98400 71150 98410 71350
rect 98480 71150 98520 71350
rect 98590 71150 98600 71350
rect 98400 71120 98600 71150
rect 98900 71350 99100 71380
rect 98900 71150 98910 71350
rect 98980 71150 99020 71350
rect 99090 71150 99100 71350
rect 98900 71120 99100 71150
rect 99400 71350 99600 71380
rect 99400 71150 99410 71350
rect 99480 71150 99520 71350
rect 99590 71150 99600 71350
rect 99400 71120 99600 71150
rect 99900 71350 100000 71380
rect 99900 71150 99910 71350
rect 99980 71150 100000 71350
rect 99900 71120 100000 71150
rect 96000 71100 96120 71120
rect 96380 71100 96620 71120
rect 96880 71100 97120 71120
rect 97380 71100 97620 71120
rect 97880 71100 98120 71120
rect 98380 71100 98620 71120
rect 98880 71100 99120 71120
rect 99380 71100 99620 71120
rect 99880 71100 100000 71120
rect 96000 71090 100000 71100
rect 96000 71020 96150 71090
rect 96350 71020 96650 71090
rect 96850 71020 97150 71090
rect 97350 71020 97650 71090
rect 97850 71020 98150 71090
rect 98350 71020 98650 71090
rect 98850 71020 99150 71090
rect 99350 71020 99650 71090
rect 99850 71020 100000 71090
rect 96000 70980 100000 71020
rect 96000 70910 96150 70980
rect 96350 70910 96650 70980
rect 96850 70910 97150 70980
rect 97350 70910 97650 70980
rect 97850 70910 98150 70980
rect 98350 70910 98650 70980
rect 98850 70910 99150 70980
rect 99350 70910 99650 70980
rect 99850 70910 100000 70980
rect 96000 70900 100000 70910
rect 96000 70880 96120 70900
rect 96380 70880 96620 70900
rect 96880 70880 97120 70900
rect 97380 70880 97620 70900
rect 97880 70880 98120 70900
rect 98380 70880 98620 70900
rect 98880 70880 99120 70900
rect 99380 70880 99620 70900
rect 99880 70880 100000 70900
rect 96000 70850 96100 70880
rect 96000 70650 96020 70850
rect 96090 70650 96100 70850
rect 96000 70620 96100 70650
rect 96400 70850 96600 70880
rect 96400 70650 96410 70850
rect 96480 70650 96520 70850
rect 96590 70650 96600 70850
rect 96400 70620 96600 70650
rect 96900 70850 97100 70880
rect 96900 70650 96910 70850
rect 96980 70650 97020 70850
rect 97090 70650 97100 70850
rect 96900 70620 97100 70650
rect 97400 70850 97600 70880
rect 97400 70650 97410 70850
rect 97480 70650 97520 70850
rect 97590 70650 97600 70850
rect 97400 70620 97600 70650
rect 97900 70850 98100 70880
rect 97900 70650 97910 70850
rect 97980 70650 98020 70850
rect 98090 70650 98100 70850
rect 97900 70620 98100 70650
rect 98400 70850 98600 70880
rect 98400 70650 98410 70850
rect 98480 70650 98520 70850
rect 98590 70650 98600 70850
rect 98400 70620 98600 70650
rect 98900 70850 99100 70880
rect 98900 70650 98910 70850
rect 98980 70650 99020 70850
rect 99090 70650 99100 70850
rect 98900 70620 99100 70650
rect 99400 70850 99600 70880
rect 99400 70650 99410 70850
rect 99480 70650 99520 70850
rect 99590 70650 99600 70850
rect 99400 70620 99600 70650
rect 99900 70850 100000 70880
rect 99900 70650 99910 70850
rect 99980 70650 100000 70850
rect 99900 70620 100000 70650
rect 96000 70600 96120 70620
rect 96380 70600 96620 70620
rect 96880 70600 97120 70620
rect 97380 70600 97620 70620
rect 97880 70600 98120 70620
rect 98380 70600 98620 70620
rect 98880 70600 99120 70620
rect 99380 70600 99620 70620
rect 99880 70600 100000 70620
rect 96000 70590 100000 70600
rect 96000 70520 96150 70590
rect 96350 70520 96650 70590
rect 96850 70520 97150 70590
rect 97350 70520 97650 70590
rect 97850 70520 98150 70590
rect 98350 70520 98650 70590
rect 98850 70520 99150 70590
rect 99350 70520 99650 70590
rect 99850 70520 100000 70590
rect 96000 70480 100000 70520
rect 96000 70410 96150 70480
rect 96350 70410 96650 70480
rect 96850 70410 97150 70480
rect 97350 70410 97650 70480
rect 97850 70410 98150 70480
rect 98350 70410 98650 70480
rect 98850 70410 99150 70480
rect 99350 70410 99650 70480
rect 99850 70410 100000 70480
rect 96000 70400 100000 70410
rect 96000 70380 96120 70400
rect 96380 70380 96620 70400
rect 96880 70380 97120 70400
rect 97380 70380 97620 70400
rect 97880 70380 98120 70400
rect 98380 70380 98620 70400
rect 98880 70380 99120 70400
rect 99380 70380 99620 70400
rect 99880 70380 100000 70400
rect 96000 70350 96100 70380
rect 96000 70150 96020 70350
rect 96090 70150 96100 70350
rect 96000 70120 96100 70150
rect 96400 70350 96600 70380
rect 96400 70150 96410 70350
rect 96480 70150 96520 70350
rect 96590 70150 96600 70350
rect 96400 70120 96600 70150
rect 96900 70350 97100 70380
rect 96900 70150 96910 70350
rect 96980 70150 97020 70350
rect 97090 70150 97100 70350
rect 96900 70120 97100 70150
rect 97400 70350 97600 70380
rect 97400 70150 97410 70350
rect 97480 70150 97520 70350
rect 97590 70150 97600 70350
rect 97400 70120 97600 70150
rect 97900 70350 98100 70380
rect 97900 70150 97910 70350
rect 97980 70150 98020 70350
rect 98090 70150 98100 70350
rect 97900 70120 98100 70150
rect 98400 70350 98600 70380
rect 98400 70150 98410 70350
rect 98480 70150 98520 70350
rect 98590 70150 98600 70350
rect 98400 70120 98600 70150
rect 98900 70350 99100 70380
rect 98900 70150 98910 70350
rect 98980 70150 99020 70350
rect 99090 70150 99100 70350
rect 98900 70120 99100 70150
rect 99400 70350 99600 70380
rect 99400 70150 99410 70350
rect 99480 70150 99520 70350
rect 99590 70150 99600 70350
rect 99400 70120 99600 70150
rect 99900 70350 100000 70380
rect 99900 70150 99910 70350
rect 99980 70150 100000 70350
rect 99900 70120 100000 70150
rect 96000 70100 96120 70120
rect 96380 70100 96620 70120
rect 96880 70100 97120 70120
rect 97380 70100 97620 70120
rect 97880 70100 98120 70120
rect 98380 70100 98620 70120
rect 98880 70100 99120 70120
rect 99380 70100 99620 70120
rect 99880 70100 100000 70120
rect 96000 70090 100000 70100
rect 96000 70020 96150 70090
rect 96350 70020 96650 70090
rect 96850 70020 97150 70090
rect 97350 70020 97650 70090
rect 97850 70020 98150 70090
rect 98350 70020 98650 70090
rect 98850 70020 99150 70090
rect 99350 70020 99650 70090
rect 99850 70020 100000 70090
rect 96000 69980 100000 70020
rect 96000 69910 96150 69980
rect 96350 69910 96650 69980
rect 96850 69910 97150 69980
rect 97350 69910 97650 69980
rect 97850 69910 98150 69980
rect 98350 69910 98650 69980
rect 98850 69910 99150 69980
rect 99350 69910 99650 69980
rect 99850 69910 100000 69980
rect 96000 69900 100000 69910
rect 96000 69880 96120 69900
rect 96380 69880 96620 69900
rect 96880 69880 97120 69900
rect 97380 69880 97620 69900
rect 97880 69880 98120 69900
rect 98380 69880 98620 69900
rect 98880 69880 99120 69900
rect 99380 69880 99620 69900
rect 99880 69880 100000 69900
rect 96000 69850 96100 69880
rect 96000 69650 96020 69850
rect 96090 69650 96100 69850
rect 96000 69620 96100 69650
rect 96400 69850 96600 69880
rect 96400 69650 96410 69850
rect 96480 69650 96520 69850
rect 96590 69650 96600 69850
rect 96400 69620 96600 69650
rect 96900 69850 97100 69880
rect 96900 69650 96910 69850
rect 96980 69650 97020 69850
rect 97090 69650 97100 69850
rect 96900 69620 97100 69650
rect 97400 69850 97600 69880
rect 97400 69650 97410 69850
rect 97480 69650 97520 69850
rect 97590 69650 97600 69850
rect 97400 69620 97600 69650
rect 97900 69850 98100 69880
rect 97900 69650 97910 69850
rect 97980 69650 98020 69850
rect 98090 69650 98100 69850
rect 97900 69620 98100 69650
rect 98400 69850 98600 69880
rect 98400 69650 98410 69850
rect 98480 69650 98520 69850
rect 98590 69650 98600 69850
rect 98400 69620 98600 69650
rect 98900 69850 99100 69880
rect 98900 69650 98910 69850
rect 98980 69650 99020 69850
rect 99090 69650 99100 69850
rect 98900 69620 99100 69650
rect 99400 69850 99600 69880
rect 99400 69650 99410 69850
rect 99480 69650 99520 69850
rect 99590 69650 99600 69850
rect 99400 69620 99600 69650
rect 99900 69850 100000 69880
rect 99900 69650 99910 69850
rect 99980 69650 100000 69850
rect 99900 69620 100000 69650
rect 96000 69600 96120 69620
rect 96380 69600 96620 69620
rect 96880 69600 97120 69620
rect 97380 69600 97620 69620
rect 97880 69600 98120 69620
rect 98380 69600 98620 69620
rect 98880 69600 99120 69620
rect 99380 69600 99620 69620
rect 99880 69600 100000 69620
rect 96000 69590 100000 69600
rect 96000 69520 96150 69590
rect 96350 69520 96650 69590
rect 96850 69520 97150 69590
rect 97350 69520 97650 69590
rect 97850 69520 98150 69590
rect 98350 69520 98650 69590
rect 98850 69520 99150 69590
rect 99350 69520 99650 69590
rect 99850 69520 100000 69590
rect 96000 69480 100000 69520
rect 96000 69410 96150 69480
rect 96350 69410 96650 69480
rect 96850 69410 97150 69480
rect 97350 69410 97650 69480
rect 97850 69410 98150 69480
rect 98350 69410 98650 69480
rect 98850 69410 99150 69480
rect 99350 69410 99650 69480
rect 99850 69410 100000 69480
rect 96000 69400 100000 69410
rect 96000 69380 96120 69400
rect 96380 69380 96620 69400
rect 96880 69380 97120 69400
rect 97380 69380 97620 69400
rect 97880 69380 98120 69400
rect 98380 69380 98620 69400
rect 98880 69380 99120 69400
rect 99380 69380 99620 69400
rect 99880 69380 100000 69400
rect 96000 69350 96100 69380
rect 96000 69150 96020 69350
rect 96090 69150 96100 69350
rect 96000 69120 96100 69150
rect 96400 69350 96600 69380
rect 96400 69150 96410 69350
rect 96480 69150 96520 69350
rect 96590 69150 96600 69350
rect 96400 69120 96600 69150
rect 96900 69350 97100 69380
rect 96900 69150 96910 69350
rect 96980 69150 97020 69350
rect 97090 69150 97100 69350
rect 96900 69120 97100 69150
rect 97400 69350 97600 69380
rect 97400 69150 97410 69350
rect 97480 69150 97520 69350
rect 97590 69150 97600 69350
rect 97400 69120 97600 69150
rect 97900 69350 98100 69380
rect 97900 69150 97910 69350
rect 97980 69150 98020 69350
rect 98090 69150 98100 69350
rect 97900 69120 98100 69150
rect 98400 69350 98600 69380
rect 98400 69150 98410 69350
rect 98480 69150 98520 69350
rect 98590 69150 98600 69350
rect 98400 69120 98600 69150
rect 98900 69350 99100 69380
rect 98900 69150 98910 69350
rect 98980 69150 99020 69350
rect 99090 69150 99100 69350
rect 98900 69120 99100 69150
rect 99400 69350 99600 69380
rect 99400 69150 99410 69350
rect 99480 69150 99520 69350
rect 99590 69150 99600 69350
rect 99400 69120 99600 69150
rect 99900 69350 100000 69380
rect 99900 69150 99910 69350
rect 99980 69150 100000 69350
rect 99900 69120 100000 69150
rect 96000 69100 96120 69120
rect 96380 69100 96620 69120
rect 96880 69100 97120 69120
rect 97380 69100 97620 69120
rect 97880 69100 98120 69120
rect 98380 69100 98620 69120
rect 98880 69100 99120 69120
rect 99380 69100 99620 69120
rect 99880 69100 100000 69120
rect 96000 69090 100000 69100
rect 96000 69020 96150 69090
rect 96350 69020 96650 69090
rect 96850 69020 97150 69090
rect 97350 69020 97650 69090
rect 97850 69020 98150 69090
rect 98350 69020 98650 69090
rect 98850 69020 99150 69090
rect 99350 69020 99650 69090
rect 99850 69020 100000 69090
rect 96000 68980 100000 69020
rect 96000 68910 96150 68980
rect 96350 68910 96650 68980
rect 96850 68910 97150 68980
rect 97350 68910 97650 68980
rect 97850 68910 98150 68980
rect 98350 68910 98650 68980
rect 98850 68910 99150 68980
rect 99350 68910 99650 68980
rect 99850 68910 100000 68980
rect 96000 68900 100000 68910
rect 96000 68880 96120 68900
rect 96380 68880 96620 68900
rect 96880 68880 97120 68900
rect 97380 68880 97620 68900
rect 97880 68880 98120 68900
rect 98380 68880 98620 68900
rect 98880 68880 99120 68900
rect 99380 68880 99620 68900
rect 99880 68880 100000 68900
rect 96000 68850 96100 68880
rect 96000 68650 96020 68850
rect 96090 68650 96100 68850
rect 96000 68620 96100 68650
rect 96400 68850 96600 68880
rect 96400 68650 96410 68850
rect 96480 68650 96520 68850
rect 96590 68650 96600 68850
rect 96400 68620 96600 68650
rect 96900 68850 97100 68880
rect 96900 68650 96910 68850
rect 96980 68650 97020 68850
rect 97090 68650 97100 68850
rect 96900 68620 97100 68650
rect 97400 68850 97600 68880
rect 97400 68650 97410 68850
rect 97480 68650 97520 68850
rect 97590 68650 97600 68850
rect 97400 68620 97600 68650
rect 97900 68850 98100 68880
rect 97900 68650 97910 68850
rect 97980 68650 98020 68850
rect 98090 68650 98100 68850
rect 97900 68620 98100 68650
rect 98400 68850 98600 68880
rect 98400 68650 98410 68850
rect 98480 68650 98520 68850
rect 98590 68650 98600 68850
rect 98400 68620 98600 68650
rect 98900 68850 99100 68880
rect 98900 68650 98910 68850
rect 98980 68650 99020 68850
rect 99090 68650 99100 68850
rect 98900 68620 99100 68650
rect 99400 68850 99600 68880
rect 99400 68650 99410 68850
rect 99480 68650 99520 68850
rect 99590 68650 99600 68850
rect 99400 68620 99600 68650
rect 99900 68850 100000 68880
rect 99900 68650 99910 68850
rect 99980 68650 100000 68850
rect 99900 68620 100000 68650
rect 96000 68600 96120 68620
rect 96380 68600 96620 68620
rect 96880 68600 97120 68620
rect 97380 68600 97620 68620
rect 97880 68600 98120 68620
rect 98380 68600 98620 68620
rect 98880 68600 99120 68620
rect 99380 68600 99620 68620
rect 99880 68600 100000 68620
rect 96000 68590 100000 68600
rect 96000 68520 96150 68590
rect 96350 68520 96650 68590
rect 96850 68520 97150 68590
rect 97350 68520 97650 68590
rect 97850 68520 98150 68590
rect 98350 68520 98650 68590
rect 98850 68520 99150 68590
rect 99350 68520 99650 68590
rect 99850 68520 100000 68590
rect 96000 68480 100000 68520
rect 96000 68410 96150 68480
rect 96350 68410 96650 68480
rect 96850 68410 97150 68480
rect 97350 68410 97650 68480
rect 97850 68410 98150 68480
rect 98350 68410 98650 68480
rect 98850 68410 99150 68480
rect 99350 68410 99650 68480
rect 99850 68410 100000 68480
rect 96000 68400 100000 68410
rect 96000 68380 96120 68400
rect 96380 68380 96620 68400
rect 96880 68380 97120 68400
rect 97380 68380 97620 68400
rect 97880 68380 98120 68400
rect 98380 68380 98620 68400
rect 98880 68380 99120 68400
rect 99380 68380 99620 68400
rect 99880 68380 100000 68400
rect 96000 68350 96100 68380
rect 96000 68150 96020 68350
rect 96090 68150 96100 68350
rect 96000 68120 96100 68150
rect 96400 68350 96600 68380
rect 96400 68150 96410 68350
rect 96480 68150 96520 68350
rect 96590 68150 96600 68350
rect 96400 68120 96600 68150
rect 96900 68350 97100 68380
rect 96900 68150 96910 68350
rect 96980 68150 97020 68350
rect 97090 68150 97100 68350
rect 96900 68120 97100 68150
rect 97400 68350 97600 68380
rect 97400 68150 97410 68350
rect 97480 68150 97520 68350
rect 97590 68150 97600 68350
rect 97400 68120 97600 68150
rect 97900 68350 98100 68380
rect 97900 68150 97910 68350
rect 97980 68150 98020 68350
rect 98090 68150 98100 68350
rect 97900 68120 98100 68150
rect 98400 68350 98600 68380
rect 98400 68150 98410 68350
rect 98480 68150 98520 68350
rect 98590 68150 98600 68350
rect 98400 68120 98600 68150
rect 98900 68350 99100 68380
rect 98900 68150 98910 68350
rect 98980 68150 99020 68350
rect 99090 68150 99100 68350
rect 98900 68120 99100 68150
rect 99400 68350 99600 68380
rect 99400 68150 99410 68350
rect 99480 68150 99520 68350
rect 99590 68150 99600 68350
rect 99400 68120 99600 68150
rect 99900 68350 100000 68380
rect 99900 68150 99910 68350
rect 99980 68150 100000 68350
rect 99900 68120 100000 68150
rect 96000 68100 96120 68120
rect 96380 68100 96620 68120
rect 96880 68100 97120 68120
rect 97380 68100 97620 68120
rect 97880 68100 98120 68120
rect 98380 68100 98620 68120
rect 98880 68100 99120 68120
rect 99380 68100 99620 68120
rect 99880 68100 100000 68120
rect 96000 68090 100000 68100
rect 96000 68020 96150 68090
rect 96350 68020 96650 68090
rect 96850 68020 97150 68090
rect 97350 68020 97650 68090
rect 97850 68020 98150 68090
rect 98350 68020 98650 68090
rect 98850 68020 99150 68090
rect 99350 68020 99650 68090
rect 99850 68020 100000 68090
rect 96000 67980 100000 68020
rect 96000 67910 96150 67980
rect 96350 67910 96650 67980
rect 96850 67910 97150 67980
rect 97350 67910 97650 67980
rect 97850 67910 98150 67980
rect 98350 67910 98650 67980
rect 98850 67910 99150 67980
rect 99350 67910 99650 67980
rect 99850 67910 100000 67980
rect 96000 67900 100000 67910
rect 96000 67880 96120 67900
rect 96380 67880 96620 67900
rect 96880 67880 97120 67900
rect 97380 67880 97620 67900
rect 97880 67880 98120 67900
rect 98380 67880 98620 67900
rect 98880 67880 99120 67900
rect 99380 67880 99620 67900
rect 99880 67880 100000 67900
rect 96000 67850 96100 67880
rect 96000 67650 96020 67850
rect 96090 67650 96100 67850
rect 96000 67620 96100 67650
rect 96400 67850 96600 67880
rect 96400 67650 96410 67850
rect 96480 67650 96520 67850
rect 96590 67650 96600 67850
rect 96400 67620 96600 67650
rect 96900 67850 97100 67880
rect 96900 67650 96910 67850
rect 96980 67650 97020 67850
rect 97090 67650 97100 67850
rect 96900 67620 97100 67650
rect 97400 67850 97600 67880
rect 97400 67650 97410 67850
rect 97480 67650 97520 67850
rect 97590 67650 97600 67850
rect 97400 67620 97600 67650
rect 97900 67850 98100 67880
rect 97900 67650 97910 67850
rect 97980 67650 98020 67850
rect 98090 67650 98100 67850
rect 97900 67620 98100 67650
rect 98400 67850 98600 67880
rect 98400 67650 98410 67850
rect 98480 67650 98520 67850
rect 98590 67650 98600 67850
rect 98400 67620 98600 67650
rect 98900 67850 99100 67880
rect 98900 67650 98910 67850
rect 98980 67650 99020 67850
rect 99090 67650 99100 67850
rect 98900 67620 99100 67650
rect 99400 67850 99600 67880
rect 99400 67650 99410 67850
rect 99480 67650 99520 67850
rect 99590 67650 99600 67850
rect 99400 67620 99600 67650
rect 99900 67850 100000 67880
rect 99900 67650 99910 67850
rect 99980 67650 100000 67850
rect 99900 67620 100000 67650
rect 96000 67600 96120 67620
rect 96380 67600 96620 67620
rect 96880 67600 97120 67620
rect 97380 67600 97620 67620
rect 97880 67600 98120 67620
rect 98380 67600 98620 67620
rect 98880 67600 99120 67620
rect 99380 67600 99620 67620
rect 99880 67600 100000 67620
rect 96000 67590 100000 67600
rect 96000 67520 96150 67590
rect 96350 67520 96650 67590
rect 96850 67520 97150 67590
rect 97350 67520 97650 67590
rect 97850 67520 98150 67590
rect 98350 67520 98650 67590
rect 98850 67520 99150 67590
rect 99350 67520 99650 67590
rect 99850 67520 100000 67590
rect 96000 67480 100000 67520
rect 96000 67410 96150 67480
rect 96350 67410 96650 67480
rect 96850 67410 97150 67480
rect 97350 67410 97650 67480
rect 97850 67410 98150 67480
rect 98350 67410 98650 67480
rect 98850 67410 99150 67480
rect 99350 67410 99650 67480
rect 99850 67410 100000 67480
rect 96000 67400 100000 67410
rect 96000 67380 96120 67400
rect 96380 67380 96620 67400
rect 96880 67380 97120 67400
rect 97380 67380 97620 67400
rect 97880 67380 98120 67400
rect 98380 67380 98620 67400
rect 98880 67380 99120 67400
rect 99380 67380 99620 67400
rect 99880 67380 100000 67400
rect 96000 67350 96100 67380
rect 96000 67150 96020 67350
rect 96090 67150 96100 67350
rect 96000 67120 96100 67150
rect 96400 67350 96600 67380
rect 96400 67150 96410 67350
rect 96480 67150 96520 67350
rect 96590 67150 96600 67350
rect 96400 67120 96600 67150
rect 96900 67350 97100 67380
rect 96900 67150 96910 67350
rect 96980 67150 97020 67350
rect 97090 67150 97100 67350
rect 96900 67120 97100 67150
rect 97400 67350 97600 67380
rect 97400 67150 97410 67350
rect 97480 67150 97520 67350
rect 97590 67150 97600 67350
rect 97400 67120 97600 67150
rect 97900 67350 98100 67380
rect 97900 67150 97910 67350
rect 97980 67150 98020 67350
rect 98090 67150 98100 67350
rect 97900 67120 98100 67150
rect 98400 67350 98600 67380
rect 98400 67150 98410 67350
rect 98480 67150 98520 67350
rect 98590 67150 98600 67350
rect 98400 67120 98600 67150
rect 98900 67350 99100 67380
rect 98900 67150 98910 67350
rect 98980 67150 99020 67350
rect 99090 67150 99100 67350
rect 98900 67120 99100 67150
rect 99400 67350 99600 67380
rect 99400 67150 99410 67350
rect 99480 67150 99520 67350
rect 99590 67150 99600 67350
rect 99400 67120 99600 67150
rect 99900 67350 100000 67380
rect 99900 67150 99910 67350
rect 99980 67150 100000 67350
rect 99900 67120 100000 67150
rect 96000 67100 96120 67120
rect 96380 67100 96620 67120
rect 96880 67100 97120 67120
rect 97380 67100 97620 67120
rect 97880 67100 98120 67120
rect 98380 67100 98620 67120
rect 98880 67100 99120 67120
rect 99380 67100 99620 67120
rect 99880 67100 100000 67120
rect 96000 67090 100000 67100
rect 96000 67020 96150 67090
rect 96350 67020 96650 67090
rect 96850 67020 97150 67090
rect 97350 67020 97650 67090
rect 97850 67020 98150 67090
rect 98350 67020 98650 67090
rect 98850 67020 99150 67090
rect 99350 67020 99650 67090
rect 99850 67020 100000 67090
rect 96000 66980 100000 67020
rect 96000 66910 96150 66980
rect 96350 66910 96650 66980
rect 96850 66910 97150 66980
rect 97350 66910 97650 66980
rect 97850 66910 98150 66980
rect 98350 66910 98650 66980
rect 98850 66910 99150 66980
rect 99350 66910 99650 66980
rect 99850 66910 100000 66980
rect 96000 66900 100000 66910
rect 96000 66880 96120 66900
rect 96380 66880 96620 66900
rect 96880 66880 97120 66900
rect 97380 66880 97620 66900
rect 97880 66880 98120 66900
rect 98380 66880 98620 66900
rect 98880 66880 99120 66900
rect 99380 66880 99620 66900
rect 99880 66880 100000 66900
rect 96000 66850 96100 66880
rect 96000 66650 96020 66850
rect 96090 66650 96100 66850
rect 96000 66620 96100 66650
rect 96400 66850 96600 66880
rect 96400 66650 96410 66850
rect 96480 66650 96520 66850
rect 96590 66650 96600 66850
rect 96400 66620 96600 66650
rect 96900 66850 97100 66880
rect 96900 66650 96910 66850
rect 96980 66650 97020 66850
rect 97090 66650 97100 66850
rect 96900 66620 97100 66650
rect 97400 66850 97600 66880
rect 97400 66650 97410 66850
rect 97480 66650 97520 66850
rect 97590 66650 97600 66850
rect 97400 66620 97600 66650
rect 97900 66850 98100 66880
rect 97900 66650 97910 66850
rect 97980 66650 98020 66850
rect 98090 66650 98100 66850
rect 97900 66620 98100 66650
rect 98400 66850 98600 66880
rect 98400 66650 98410 66850
rect 98480 66650 98520 66850
rect 98590 66650 98600 66850
rect 98400 66620 98600 66650
rect 98900 66850 99100 66880
rect 98900 66650 98910 66850
rect 98980 66650 99020 66850
rect 99090 66650 99100 66850
rect 98900 66620 99100 66650
rect 99400 66850 99600 66880
rect 99400 66650 99410 66850
rect 99480 66650 99520 66850
rect 99590 66650 99600 66850
rect 99400 66620 99600 66650
rect 99900 66850 100000 66880
rect 99900 66650 99910 66850
rect 99980 66650 100000 66850
rect 99900 66620 100000 66650
rect 96000 66600 96120 66620
rect 96380 66600 96620 66620
rect 96880 66600 97120 66620
rect 97380 66600 97620 66620
rect 97880 66600 98120 66620
rect 98380 66600 98620 66620
rect 98880 66600 99120 66620
rect 99380 66600 99620 66620
rect 99880 66600 100000 66620
rect 96000 66590 100000 66600
rect 96000 66520 96150 66590
rect 96350 66520 96650 66590
rect 96850 66520 97150 66590
rect 97350 66520 97650 66590
rect 97850 66520 98150 66590
rect 98350 66520 98650 66590
rect 98850 66520 99150 66590
rect 99350 66520 99650 66590
rect 99850 66520 100000 66590
rect 96000 66480 100000 66520
rect 96000 66410 96150 66480
rect 96350 66410 96650 66480
rect 96850 66410 97150 66480
rect 97350 66410 97650 66480
rect 97850 66410 98150 66480
rect 98350 66410 98650 66480
rect 98850 66410 99150 66480
rect 99350 66410 99650 66480
rect 99850 66410 100000 66480
rect 96000 66400 100000 66410
rect 96000 66380 96120 66400
rect 96380 66380 96620 66400
rect 96880 66380 97120 66400
rect 97380 66380 97620 66400
rect 97880 66380 98120 66400
rect 98380 66380 98620 66400
rect 98880 66380 99120 66400
rect 99380 66380 99620 66400
rect 99880 66380 100000 66400
rect 96000 66350 96100 66380
rect 96000 66150 96020 66350
rect 96090 66150 96100 66350
rect 96000 66120 96100 66150
rect 96400 66350 96600 66380
rect 96400 66150 96410 66350
rect 96480 66150 96520 66350
rect 96590 66150 96600 66350
rect 96400 66120 96600 66150
rect 96900 66350 97100 66380
rect 96900 66150 96910 66350
rect 96980 66150 97020 66350
rect 97090 66150 97100 66350
rect 96900 66120 97100 66150
rect 97400 66350 97600 66380
rect 97400 66150 97410 66350
rect 97480 66150 97520 66350
rect 97590 66150 97600 66350
rect 97400 66120 97600 66150
rect 97900 66350 98100 66380
rect 97900 66150 97910 66350
rect 97980 66150 98020 66350
rect 98090 66150 98100 66350
rect 97900 66120 98100 66150
rect 98400 66350 98600 66380
rect 98400 66150 98410 66350
rect 98480 66150 98520 66350
rect 98590 66150 98600 66350
rect 98400 66120 98600 66150
rect 98900 66350 99100 66380
rect 98900 66150 98910 66350
rect 98980 66150 99020 66350
rect 99090 66150 99100 66350
rect 98900 66120 99100 66150
rect 99400 66350 99600 66380
rect 99400 66150 99410 66350
rect 99480 66150 99520 66350
rect 99590 66150 99600 66350
rect 99400 66120 99600 66150
rect 99900 66350 100000 66380
rect 99900 66150 99910 66350
rect 99980 66150 100000 66350
rect 99900 66120 100000 66150
rect 96000 66100 96120 66120
rect 96380 66100 96620 66120
rect 96880 66100 97120 66120
rect 97380 66100 97620 66120
rect 97880 66100 98120 66120
rect 98380 66100 98620 66120
rect 98880 66100 99120 66120
rect 99380 66100 99620 66120
rect 99880 66100 100000 66120
rect 96000 66090 100000 66100
rect 96000 66020 96150 66090
rect 96350 66020 96650 66090
rect 96850 66020 97150 66090
rect 97350 66020 97650 66090
rect 97850 66020 98150 66090
rect 98350 66020 98650 66090
rect 98850 66020 99150 66090
rect 99350 66020 99650 66090
rect 99850 66020 100000 66090
rect 96000 65980 100000 66020
rect 96000 65910 96150 65980
rect 96350 65910 96650 65980
rect 96850 65910 97150 65980
rect 97350 65910 97650 65980
rect 97850 65910 98150 65980
rect 98350 65910 98650 65980
rect 98850 65910 99150 65980
rect 99350 65910 99650 65980
rect 99850 65910 100000 65980
rect 96000 65900 100000 65910
rect 96000 65880 96120 65900
rect 96380 65880 96620 65900
rect 96880 65880 97120 65900
rect 97380 65880 97620 65900
rect 97880 65880 98120 65900
rect 98380 65880 98620 65900
rect 98880 65880 99120 65900
rect 99380 65880 99620 65900
rect 99880 65880 100000 65900
rect 96000 65850 96100 65880
rect 96000 65650 96020 65850
rect 96090 65650 96100 65850
rect 96000 65620 96100 65650
rect 96400 65850 96600 65880
rect 96400 65650 96410 65850
rect 96480 65650 96520 65850
rect 96590 65650 96600 65850
rect 96400 65620 96600 65650
rect 96900 65850 97100 65880
rect 96900 65650 96910 65850
rect 96980 65650 97020 65850
rect 97090 65650 97100 65850
rect 96900 65620 97100 65650
rect 97400 65850 97600 65880
rect 97400 65650 97410 65850
rect 97480 65650 97520 65850
rect 97590 65650 97600 65850
rect 97400 65620 97600 65650
rect 97900 65850 98100 65880
rect 97900 65650 97910 65850
rect 97980 65650 98020 65850
rect 98090 65650 98100 65850
rect 97900 65620 98100 65650
rect 98400 65850 98600 65880
rect 98400 65650 98410 65850
rect 98480 65650 98520 65850
rect 98590 65650 98600 65850
rect 98400 65620 98600 65650
rect 98900 65850 99100 65880
rect 98900 65650 98910 65850
rect 98980 65650 99020 65850
rect 99090 65650 99100 65850
rect 98900 65620 99100 65650
rect 99400 65850 99600 65880
rect 99400 65650 99410 65850
rect 99480 65650 99520 65850
rect 99590 65650 99600 65850
rect 99400 65620 99600 65650
rect 99900 65850 100000 65880
rect 99900 65650 99910 65850
rect 99980 65650 100000 65850
rect 99900 65620 100000 65650
rect 96000 65600 96120 65620
rect 96380 65600 96620 65620
rect 96880 65600 97120 65620
rect 97380 65600 97620 65620
rect 97880 65600 98120 65620
rect 98380 65600 98620 65620
rect 98880 65600 99120 65620
rect 99380 65600 99620 65620
rect 99880 65600 100000 65620
rect 96000 65590 100000 65600
rect 96000 65520 96150 65590
rect 96350 65520 96650 65590
rect 96850 65520 97150 65590
rect 97350 65520 97650 65590
rect 97850 65520 98150 65590
rect 98350 65520 98650 65590
rect 98850 65520 99150 65590
rect 99350 65520 99650 65590
rect 99850 65520 100000 65590
rect 96000 65480 100000 65520
rect 96000 65410 96150 65480
rect 96350 65410 96650 65480
rect 96850 65410 97150 65480
rect 97350 65410 97650 65480
rect 97850 65410 98150 65480
rect 98350 65410 98650 65480
rect 98850 65410 99150 65480
rect 99350 65410 99650 65480
rect 99850 65410 100000 65480
rect 96000 65400 100000 65410
rect 96000 65380 96120 65400
rect 96380 65380 96620 65400
rect 96880 65380 97120 65400
rect 97380 65380 97620 65400
rect 97880 65380 98120 65400
rect 98380 65380 98620 65400
rect 98880 65380 99120 65400
rect 99380 65380 99620 65400
rect 99880 65380 100000 65400
rect 96000 65350 96100 65380
rect 96000 65150 96020 65350
rect 96090 65150 96100 65350
rect 96000 65120 96100 65150
rect 96400 65350 96600 65380
rect 96400 65150 96410 65350
rect 96480 65150 96520 65350
rect 96590 65150 96600 65350
rect 96400 65120 96600 65150
rect 96900 65350 97100 65380
rect 96900 65150 96910 65350
rect 96980 65150 97020 65350
rect 97090 65150 97100 65350
rect 96900 65120 97100 65150
rect 97400 65350 97600 65380
rect 97400 65150 97410 65350
rect 97480 65150 97520 65350
rect 97590 65150 97600 65350
rect 97400 65120 97600 65150
rect 97900 65350 98100 65380
rect 97900 65150 97910 65350
rect 97980 65150 98020 65350
rect 98090 65150 98100 65350
rect 97900 65120 98100 65150
rect 98400 65350 98600 65380
rect 98400 65150 98410 65350
rect 98480 65150 98520 65350
rect 98590 65150 98600 65350
rect 98400 65120 98600 65150
rect 98900 65350 99100 65380
rect 98900 65150 98910 65350
rect 98980 65150 99020 65350
rect 99090 65150 99100 65350
rect 98900 65120 99100 65150
rect 99400 65350 99600 65380
rect 99400 65150 99410 65350
rect 99480 65150 99520 65350
rect 99590 65150 99600 65350
rect 99400 65120 99600 65150
rect 99900 65350 100000 65380
rect 99900 65150 99910 65350
rect 99980 65150 100000 65350
rect 99900 65120 100000 65150
rect 96000 65100 96120 65120
rect 96380 65100 96620 65120
rect 96880 65100 97120 65120
rect 97380 65100 97620 65120
rect 97880 65100 98120 65120
rect 98380 65100 98620 65120
rect 98880 65100 99120 65120
rect 99380 65100 99620 65120
rect 99880 65100 100000 65120
rect 96000 65090 100000 65100
rect 96000 65020 96150 65090
rect 96350 65020 96650 65090
rect 96850 65020 97150 65090
rect 97350 65020 97650 65090
rect 97850 65020 98150 65090
rect 98350 65020 98650 65090
rect 98850 65020 99150 65090
rect 99350 65020 99650 65090
rect 99850 65020 100000 65090
rect 96000 64980 100000 65020
rect 96000 64910 96150 64980
rect 96350 64910 96650 64980
rect 96850 64910 97150 64980
rect 97350 64910 97650 64980
rect 97850 64910 98150 64980
rect 98350 64910 98650 64980
rect 98850 64910 99150 64980
rect 99350 64910 99650 64980
rect 99850 64910 100000 64980
rect 96000 64900 100000 64910
rect 96000 64880 96120 64900
rect 96380 64880 96620 64900
rect 96880 64880 97120 64900
rect 97380 64880 97620 64900
rect 97880 64880 98120 64900
rect 98380 64880 98620 64900
rect 98880 64880 99120 64900
rect 99380 64880 99620 64900
rect 99880 64880 100000 64900
rect 96000 64850 96100 64880
rect 96000 64650 96020 64850
rect 96090 64650 96100 64850
rect 96000 64620 96100 64650
rect 96400 64850 96600 64880
rect 96400 64650 96410 64850
rect 96480 64650 96520 64850
rect 96590 64650 96600 64850
rect 96400 64620 96600 64650
rect 96900 64850 97100 64880
rect 96900 64650 96910 64850
rect 96980 64650 97020 64850
rect 97090 64650 97100 64850
rect 96900 64620 97100 64650
rect 97400 64850 97600 64880
rect 97400 64650 97410 64850
rect 97480 64650 97520 64850
rect 97590 64650 97600 64850
rect 97400 64620 97600 64650
rect 97900 64850 98100 64880
rect 97900 64650 97910 64850
rect 97980 64650 98020 64850
rect 98090 64650 98100 64850
rect 97900 64620 98100 64650
rect 98400 64850 98600 64880
rect 98400 64650 98410 64850
rect 98480 64650 98520 64850
rect 98590 64650 98600 64850
rect 98400 64620 98600 64650
rect 98900 64850 99100 64880
rect 98900 64650 98910 64850
rect 98980 64650 99020 64850
rect 99090 64650 99100 64850
rect 98900 64620 99100 64650
rect 99400 64850 99600 64880
rect 99400 64650 99410 64850
rect 99480 64650 99520 64850
rect 99590 64650 99600 64850
rect 99400 64620 99600 64650
rect 99900 64850 100000 64880
rect 99900 64650 99910 64850
rect 99980 64650 100000 64850
rect 99900 64620 100000 64650
rect 96000 64600 96120 64620
rect 96380 64600 96620 64620
rect 96880 64600 97120 64620
rect 97380 64600 97620 64620
rect 97880 64600 98120 64620
rect 98380 64600 98620 64620
rect 98880 64600 99120 64620
rect 99380 64600 99620 64620
rect 99880 64600 100000 64620
rect 96000 64590 100000 64600
rect 96000 64520 96150 64590
rect 96350 64520 96650 64590
rect 96850 64520 97150 64590
rect 97350 64520 97650 64590
rect 97850 64520 98150 64590
rect 98350 64520 98650 64590
rect 98850 64520 99150 64590
rect 99350 64520 99650 64590
rect 99850 64520 100000 64590
rect 96000 64480 100000 64520
rect 96000 64410 96150 64480
rect 96350 64410 96650 64480
rect 96850 64410 97150 64480
rect 97350 64410 97650 64480
rect 97850 64410 98150 64480
rect 98350 64410 98650 64480
rect 98850 64410 99150 64480
rect 99350 64410 99650 64480
rect 99850 64410 100000 64480
rect 96000 64400 100000 64410
rect 96000 64380 96120 64400
rect 96380 64380 96620 64400
rect 96880 64380 97120 64400
rect 97380 64380 97620 64400
rect 97880 64380 98120 64400
rect 98380 64380 98620 64400
rect 98880 64380 99120 64400
rect 99380 64380 99620 64400
rect 99880 64380 100000 64400
rect 96000 64350 96100 64380
rect 96000 64150 96020 64350
rect 96090 64150 96100 64350
rect 96000 64120 96100 64150
rect 96400 64350 96600 64380
rect 96400 64150 96410 64350
rect 96480 64150 96520 64350
rect 96590 64150 96600 64350
rect 96400 64120 96600 64150
rect 96900 64350 97100 64380
rect 96900 64150 96910 64350
rect 96980 64150 97020 64350
rect 97090 64150 97100 64350
rect 96900 64120 97100 64150
rect 97400 64350 97600 64380
rect 97400 64150 97410 64350
rect 97480 64150 97520 64350
rect 97590 64150 97600 64350
rect 97400 64120 97600 64150
rect 97900 64350 98100 64380
rect 97900 64150 97910 64350
rect 97980 64150 98020 64350
rect 98090 64150 98100 64350
rect 97900 64120 98100 64150
rect 98400 64350 98600 64380
rect 98400 64150 98410 64350
rect 98480 64150 98520 64350
rect 98590 64150 98600 64350
rect 98400 64120 98600 64150
rect 98900 64350 99100 64380
rect 98900 64150 98910 64350
rect 98980 64150 99020 64350
rect 99090 64150 99100 64350
rect 98900 64120 99100 64150
rect 99400 64350 99600 64380
rect 99400 64150 99410 64350
rect 99480 64150 99520 64350
rect 99590 64150 99600 64350
rect 99400 64120 99600 64150
rect 99900 64350 100000 64380
rect 99900 64150 99910 64350
rect 99980 64150 100000 64350
rect 99900 64120 100000 64150
rect 96000 64100 96120 64120
rect 96380 64100 96620 64120
rect 96880 64100 97120 64120
rect 97380 64100 97620 64120
rect 97880 64100 98120 64120
rect 98380 64100 98620 64120
rect 98880 64100 99120 64120
rect 99380 64100 99620 64120
rect 99880 64100 100000 64120
rect 96000 64090 100000 64100
rect 96000 64020 96150 64090
rect 96350 64020 96650 64090
rect 96850 64020 97150 64090
rect 97350 64020 97650 64090
rect 97850 64020 98150 64090
rect 98350 64020 98650 64090
rect 98850 64020 99150 64090
rect 99350 64020 99650 64090
rect 99850 64020 100000 64090
rect 96000 63980 100000 64020
rect 96000 63910 96150 63980
rect 96350 63910 96650 63980
rect 96850 63910 97150 63980
rect 97350 63910 97650 63980
rect 97850 63910 98150 63980
rect 98350 63910 98650 63980
rect 98850 63910 99150 63980
rect 99350 63910 99650 63980
rect 99850 63910 100000 63980
rect 96000 63900 100000 63910
rect 96000 63880 96120 63900
rect 96380 63880 96620 63900
rect 96880 63880 97120 63900
rect 97380 63880 97620 63900
rect 97880 63880 98120 63900
rect 98380 63880 98620 63900
rect 98880 63880 99120 63900
rect 99380 63880 99620 63900
rect 99880 63880 100000 63900
rect 96000 63850 96100 63880
rect 96000 63650 96020 63850
rect 96090 63650 96100 63850
rect 96000 63620 96100 63650
rect 96400 63850 96600 63880
rect 96400 63650 96410 63850
rect 96480 63650 96520 63850
rect 96590 63650 96600 63850
rect 96400 63620 96600 63650
rect 96900 63850 97100 63880
rect 96900 63650 96910 63850
rect 96980 63650 97020 63850
rect 97090 63650 97100 63850
rect 96900 63620 97100 63650
rect 97400 63850 97600 63880
rect 97400 63650 97410 63850
rect 97480 63650 97520 63850
rect 97590 63650 97600 63850
rect 97400 63620 97600 63650
rect 97900 63850 98100 63880
rect 97900 63650 97910 63850
rect 97980 63650 98020 63850
rect 98090 63650 98100 63850
rect 97900 63620 98100 63650
rect 98400 63850 98600 63880
rect 98400 63650 98410 63850
rect 98480 63650 98520 63850
rect 98590 63650 98600 63850
rect 98400 63620 98600 63650
rect 98900 63850 99100 63880
rect 98900 63650 98910 63850
rect 98980 63650 99020 63850
rect 99090 63650 99100 63850
rect 98900 63620 99100 63650
rect 99400 63850 99600 63880
rect 99400 63650 99410 63850
rect 99480 63650 99520 63850
rect 99590 63650 99600 63850
rect 99400 63620 99600 63650
rect 99900 63850 100000 63880
rect 99900 63650 99910 63850
rect 99980 63650 100000 63850
rect 99900 63620 100000 63650
rect 96000 63600 96120 63620
rect 96380 63600 96620 63620
rect 96880 63600 97120 63620
rect 97380 63600 97620 63620
rect 97880 63600 98120 63620
rect 98380 63600 98620 63620
rect 98880 63600 99120 63620
rect 99380 63600 99620 63620
rect 99880 63600 100000 63620
rect 96000 63590 100000 63600
rect 96000 63520 96150 63590
rect 96350 63520 96650 63590
rect 96850 63520 97150 63590
rect 97350 63520 97650 63590
rect 97850 63520 98150 63590
rect 98350 63520 98650 63590
rect 98850 63520 99150 63590
rect 99350 63520 99650 63590
rect 99850 63520 100000 63590
rect 96000 63480 100000 63520
rect 96000 63410 96150 63480
rect 96350 63410 96650 63480
rect 96850 63410 97150 63480
rect 97350 63410 97650 63480
rect 97850 63410 98150 63480
rect 98350 63410 98650 63480
rect 98850 63410 99150 63480
rect 99350 63410 99650 63480
rect 99850 63410 100000 63480
rect 96000 63400 100000 63410
rect 96000 63380 96120 63400
rect 96380 63380 96620 63400
rect 96880 63380 97120 63400
rect 97380 63380 97620 63400
rect 97880 63380 98120 63400
rect 98380 63380 98620 63400
rect 98880 63380 99120 63400
rect 99380 63380 99620 63400
rect 99880 63380 100000 63400
rect 96000 63350 96100 63380
rect 96000 63150 96020 63350
rect 96090 63150 96100 63350
rect 96000 63120 96100 63150
rect 96400 63350 96600 63380
rect 96400 63150 96410 63350
rect 96480 63150 96520 63350
rect 96590 63150 96600 63350
rect 96400 63120 96600 63150
rect 96900 63350 97100 63380
rect 96900 63150 96910 63350
rect 96980 63150 97020 63350
rect 97090 63150 97100 63350
rect 96900 63120 97100 63150
rect 97400 63350 97600 63380
rect 97400 63150 97410 63350
rect 97480 63150 97520 63350
rect 97590 63150 97600 63350
rect 97400 63120 97600 63150
rect 97900 63350 98100 63380
rect 97900 63150 97910 63350
rect 97980 63150 98020 63350
rect 98090 63150 98100 63350
rect 97900 63120 98100 63150
rect 98400 63350 98600 63380
rect 98400 63150 98410 63350
rect 98480 63150 98520 63350
rect 98590 63150 98600 63350
rect 98400 63120 98600 63150
rect 98900 63350 99100 63380
rect 98900 63150 98910 63350
rect 98980 63150 99020 63350
rect 99090 63150 99100 63350
rect 98900 63120 99100 63150
rect 99400 63350 99600 63380
rect 99400 63150 99410 63350
rect 99480 63150 99520 63350
rect 99590 63150 99600 63350
rect 99400 63120 99600 63150
rect 99900 63350 100000 63380
rect 99900 63150 99910 63350
rect 99980 63150 100000 63350
rect 99900 63120 100000 63150
rect 96000 63100 96120 63120
rect 96380 63100 96620 63120
rect 96880 63100 97120 63120
rect 97380 63100 97620 63120
rect 97880 63100 98120 63120
rect 98380 63100 98620 63120
rect 98880 63100 99120 63120
rect 99380 63100 99620 63120
rect 99880 63100 100000 63120
rect 96000 63090 100000 63100
rect 96000 63020 96150 63090
rect 96350 63020 96650 63090
rect 96850 63020 97150 63090
rect 97350 63020 97650 63090
rect 97850 63020 98150 63090
rect 98350 63020 98650 63090
rect 98850 63020 99150 63090
rect 99350 63020 99650 63090
rect 99850 63020 100000 63090
rect 96000 62980 100000 63020
rect 96000 62910 96150 62980
rect 96350 62910 96650 62980
rect 96850 62910 97150 62980
rect 97350 62910 97650 62980
rect 97850 62910 98150 62980
rect 98350 62910 98650 62980
rect 98850 62910 99150 62980
rect 99350 62910 99650 62980
rect 99850 62910 100000 62980
rect 96000 62900 100000 62910
rect 96000 62880 96120 62900
rect 96380 62880 96620 62900
rect 96880 62880 97120 62900
rect 97380 62880 97620 62900
rect 97880 62880 98120 62900
rect 98380 62880 98620 62900
rect 98880 62880 99120 62900
rect 99380 62880 99620 62900
rect 99880 62880 100000 62900
rect 96000 62850 96100 62880
rect 96000 62650 96020 62850
rect 96090 62650 96100 62850
rect 96000 62620 96100 62650
rect 96400 62850 96600 62880
rect 96400 62650 96410 62850
rect 96480 62650 96520 62850
rect 96590 62650 96600 62850
rect 96400 62620 96600 62650
rect 96900 62850 97100 62880
rect 96900 62650 96910 62850
rect 96980 62650 97020 62850
rect 97090 62650 97100 62850
rect 96900 62620 97100 62650
rect 97400 62850 97600 62880
rect 97400 62650 97410 62850
rect 97480 62650 97520 62850
rect 97590 62650 97600 62850
rect 97400 62620 97600 62650
rect 97900 62850 98100 62880
rect 97900 62650 97910 62850
rect 97980 62650 98020 62850
rect 98090 62650 98100 62850
rect 97900 62620 98100 62650
rect 98400 62850 98600 62880
rect 98400 62650 98410 62850
rect 98480 62650 98520 62850
rect 98590 62650 98600 62850
rect 98400 62620 98600 62650
rect 98900 62850 99100 62880
rect 98900 62650 98910 62850
rect 98980 62650 99020 62850
rect 99090 62650 99100 62850
rect 98900 62620 99100 62650
rect 99400 62850 99600 62880
rect 99400 62650 99410 62850
rect 99480 62650 99520 62850
rect 99590 62650 99600 62850
rect 99400 62620 99600 62650
rect 99900 62850 100000 62880
rect 99900 62650 99910 62850
rect 99980 62650 100000 62850
rect 99900 62620 100000 62650
rect 96000 62600 96120 62620
rect 96380 62600 96620 62620
rect 96880 62600 97120 62620
rect 97380 62600 97620 62620
rect 97880 62600 98120 62620
rect 98380 62600 98620 62620
rect 98880 62600 99120 62620
rect 99380 62600 99620 62620
rect 99880 62600 100000 62620
rect 96000 62590 100000 62600
rect 96000 62520 96150 62590
rect 96350 62520 96650 62590
rect 96850 62520 97150 62590
rect 97350 62520 97650 62590
rect 97850 62520 98150 62590
rect 98350 62520 98650 62590
rect 98850 62520 99150 62590
rect 99350 62520 99650 62590
rect 99850 62520 100000 62590
rect 96000 62480 100000 62520
rect 96000 62410 96150 62480
rect 96350 62410 96650 62480
rect 96850 62410 97150 62480
rect 97350 62410 97650 62480
rect 97850 62410 98150 62480
rect 98350 62410 98650 62480
rect 98850 62410 99150 62480
rect 99350 62410 99650 62480
rect 99850 62410 100000 62480
rect 96000 62400 100000 62410
rect 96000 62380 96120 62400
rect 96380 62380 96620 62400
rect 96880 62380 97120 62400
rect 97380 62380 97620 62400
rect 97880 62380 98120 62400
rect 98380 62380 98620 62400
rect 98880 62380 99120 62400
rect 99380 62380 99620 62400
rect 99880 62380 100000 62400
rect 96000 62350 96100 62380
rect 96000 62150 96020 62350
rect 96090 62150 96100 62350
rect 96000 62120 96100 62150
rect 96400 62350 96600 62380
rect 96400 62150 96410 62350
rect 96480 62150 96520 62350
rect 96590 62150 96600 62350
rect 96400 62120 96600 62150
rect 96900 62350 97100 62380
rect 96900 62150 96910 62350
rect 96980 62150 97020 62350
rect 97090 62150 97100 62350
rect 96900 62120 97100 62150
rect 97400 62350 97600 62380
rect 97400 62150 97410 62350
rect 97480 62150 97520 62350
rect 97590 62150 97600 62350
rect 97400 62120 97600 62150
rect 97900 62350 98100 62380
rect 97900 62150 97910 62350
rect 97980 62150 98020 62350
rect 98090 62150 98100 62350
rect 97900 62120 98100 62150
rect 98400 62350 98600 62380
rect 98400 62150 98410 62350
rect 98480 62150 98520 62350
rect 98590 62150 98600 62350
rect 98400 62120 98600 62150
rect 98900 62350 99100 62380
rect 98900 62150 98910 62350
rect 98980 62150 99020 62350
rect 99090 62150 99100 62350
rect 98900 62120 99100 62150
rect 99400 62350 99600 62380
rect 99400 62150 99410 62350
rect 99480 62150 99520 62350
rect 99590 62150 99600 62350
rect 99400 62120 99600 62150
rect 99900 62350 100000 62380
rect 99900 62150 99910 62350
rect 99980 62150 100000 62350
rect 99900 62120 100000 62150
rect 96000 62100 96120 62120
rect 96380 62100 96620 62120
rect 96880 62100 97120 62120
rect 97380 62100 97620 62120
rect 97880 62100 98120 62120
rect 98380 62100 98620 62120
rect 98880 62100 99120 62120
rect 99380 62100 99620 62120
rect 99880 62100 100000 62120
rect 96000 62090 100000 62100
rect 96000 62020 96150 62090
rect 96350 62020 96650 62090
rect 96850 62020 97150 62090
rect 97350 62020 97650 62090
rect 97850 62020 98150 62090
rect 98350 62020 98650 62090
rect 98850 62020 99150 62090
rect 99350 62020 99650 62090
rect 99850 62020 100000 62090
rect 96000 61980 100000 62020
rect 96000 61910 96150 61980
rect 96350 61910 96650 61980
rect 96850 61910 97150 61980
rect 97350 61910 97650 61980
rect 97850 61910 98150 61980
rect 98350 61910 98650 61980
rect 98850 61910 99150 61980
rect 99350 61910 99650 61980
rect 99850 61910 100000 61980
rect 96000 61900 100000 61910
rect 96000 61880 96120 61900
rect 96380 61880 96620 61900
rect 96880 61880 97120 61900
rect 97380 61880 97620 61900
rect 97880 61880 98120 61900
rect 98380 61880 98620 61900
rect 98880 61880 99120 61900
rect 99380 61880 99620 61900
rect 99880 61880 100000 61900
rect 96000 61850 96100 61880
rect 96000 61650 96020 61850
rect 96090 61650 96100 61850
rect 96000 61620 96100 61650
rect 96400 61850 96600 61880
rect 96400 61650 96410 61850
rect 96480 61650 96520 61850
rect 96590 61650 96600 61850
rect 96400 61620 96600 61650
rect 96900 61850 97100 61880
rect 96900 61650 96910 61850
rect 96980 61650 97020 61850
rect 97090 61650 97100 61850
rect 96900 61620 97100 61650
rect 97400 61850 97600 61880
rect 97400 61650 97410 61850
rect 97480 61650 97520 61850
rect 97590 61650 97600 61850
rect 97400 61620 97600 61650
rect 97900 61850 98100 61880
rect 97900 61650 97910 61850
rect 97980 61650 98020 61850
rect 98090 61650 98100 61850
rect 97900 61620 98100 61650
rect 98400 61850 98600 61880
rect 98400 61650 98410 61850
rect 98480 61650 98520 61850
rect 98590 61650 98600 61850
rect 98400 61620 98600 61650
rect 98900 61850 99100 61880
rect 98900 61650 98910 61850
rect 98980 61650 99020 61850
rect 99090 61650 99100 61850
rect 98900 61620 99100 61650
rect 99400 61850 99600 61880
rect 99400 61650 99410 61850
rect 99480 61650 99520 61850
rect 99590 61650 99600 61850
rect 99400 61620 99600 61650
rect 99900 61850 100000 61880
rect 99900 61650 99910 61850
rect 99980 61650 100000 61850
rect 99900 61620 100000 61650
rect 96000 61600 96120 61620
rect 96380 61600 96620 61620
rect 96880 61600 97120 61620
rect 97380 61600 97620 61620
rect 97880 61600 98120 61620
rect 98380 61600 98620 61620
rect 98880 61600 99120 61620
rect 99380 61600 99620 61620
rect 99880 61600 100000 61620
rect 96000 61590 100000 61600
rect 96000 61520 96150 61590
rect 96350 61520 96650 61590
rect 96850 61520 97150 61590
rect 97350 61520 97650 61590
rect 97850 61520 98150 61590
rect 98350 61520 98650 61590
rect 98850 61520 99150 61590
rect 99350 61520 99650 61590
rect 99850 61520 100000 61590
rect 96000 61480 100000 61520
rect 96000 61410 96150 61480
rect 96350 61410 96650 61480
rect 96850 61410 97150 61480
rect 97350 61410 97650 61480
rect 97850 61410 98150 61480
rect 98350 61410 98650 61480
rect 98850 61410 99150 61480
rect 99350 61410 99650 61480
rect 99850 61410 100000 61480
rect 96000 61400 100000 61410
rect 96000 61380 96120 61400
rect 96380 61380 96620 61400
rect 96880 61380 97120 61400
rect 97380 61380 97620 61400
rect 97880 61380 98120 61400
rect 98380 61380 98620 61400
rect 98880 61380 99120 61400
rect 99380 61380 99620 61400
rect 99880 61380 100000 61400
rect 96000 61350 96100 61380
rect 96000 61150 96020 61350
rect 96090 61150 96100 61350
rect 96000 61120 96100 61150
rect 96400 61350 96600 61380
rect 96400 61150 96410 61350
rect 96480 61150 96520 61350
rect 96590 61150 96600 61350
rect 96400 61120 96600 61150
rect 96900 61350 97100 61380
rect 96900 61150 96910 61350
rect 96980 61150 97020 61350
rect 97090 61150 97100 61350
rect 96900 61120 97100 61150
rect 97400 61350 97600 61380
rect 97400 61150 97410 61350
rect 97480 61150 97520 61350
rect 97590 61150 97600 61350
rect 97400 61120 97600 61150
rect 97900 61350 98100 61380
rect 97900 61150 97910 61350
rect 97980 61150 98020 61350
rect 98090 61150 98100 61350
rect 97900 61120 98100 61150
rect 98400 61350 98600 61380
rect 98400 61150 98410 61350
rect 98480 61150 98520 61350
rect 98590 61150 98600 61350
rect 98400 61120 98600 61150
rect 98900 61350 99100 61380
rect 98900 61150 98910 61350
rect 98980 61150 99020 61350
rect 99090 61150 99100 61350
rect 98900 61120 99100 61150
rect 99400 61350 99600 61380
rect 99400 61150 99410 61350
rect 99480 61150 99520 61350
rect 99590 61150 99600 61350
rect 99400 61120 99600 61150
rect 99900 61350 100000 61380
rect 99900 61150 99910 61350
rect 99980 61150 100000 61350
rect 99900 61120 100000 61150
rect 96000 61100 96120 61120
rect 96380 61100 96620 61120
rect 96880 61100 97120 61120
rect 97380 61100 97620 61120
rect 97880 61100 98120 61120
rect 98380 61100 98620 61120
rect 98880 61100 99120 61120
rect 99380 61100 99620 61120
rect 99880 61100 100000 61120
rect 96000 61090 100000 61100
rect 96000 61020 96150 61090
rect 96350 61020 96650 61090
rect 96850 61020 97150 61090
rect 97350 61020 97650 61090
rect 97850 61020 98150 61090
rect 98350 61020 98650 61090
rect 98850 61020 99150 61090
rect 99350 61020 99650 61090
rect 99850 61020 100000 61090
rect 96000 60980 100000 61020
rect 96000 60910 96150 60980
rect 96350 60910 96650 60980
rect 96850 60910 97150 60980
rect 97350 60910 97650 60980
rect 97850 60910 98150 60980
rect 98350 60910 98650 60980
rect 98850 60910 99150 60980
rect 99350 60910 99650 60980
rect 99850 60910 100000 60980
rect 96000 60900 100000 60910
rect 96000 60880 96120 60900
rect 96380 60880 96620 60900
rect 96880 60880 97120 60900
rect 97380 60880 97620 60900
rect 97880 60880 98120 60900
rect 98380 60880 98620 60900
rect 98880 60880 99120 60900
rect 99380 60880 99620 60900
rect 99880 60880 100000 60900
rect 96000 60850 96100 60880
rect 96000 60650 96020 60850
rect 96090 60650 96100 60850
rect 96000 60620 96100 60650
rect 96400 60850 96600 60880
rect 96400 60650 96410 60850
rect 96480 60650 96520 60850
rect 96590 60650 96600 60850
rect 96400 60620 96600 60650
rect 96900 60850 97100 60880
rect 96900 60650 96910 60850
rect 96980 60650 97020 60850
rect 97090 60650 97100 60850
rect 96900 60620 97100 60650
rect 97400 60850 97600 60880
rect 97400 60650 97410 60850
rect 97480 60650 97520 60850
rect 97590 60650 97600 60850
rect 97400 60620 97600 60650
rect 97900 60850 98100 60880
rect 97900 60650 97910 60850
rect 97980 60650 98020 60850
rect 98090 60650 98100 60850
rect 97900 60620 98100 60650
rect 98400 60850 98600 60880
rect 98400 60650 98410 60850
rect 98480 60650 98520 60850
rect 98590 60650 98600 60850
rect 98400 60620 98600 60650
rect 98900 60850 99100 60880
rect 98900 60650 98910 60850
rect 98980 60650 99020 60850
rect 99090 60650 99100 60850
rect 98900 60620 99100 60650
rect 99400 60850 99600 60880
rect 99400 60650 99410 60850
rect 99480 60650 99520 60850
rect 99590 60650 99600 60850
rect 99400 60620 99600 60650
rect 99900 60850 100000 60880
rect 99900 60650 99910 60850
rect 99980 60650 100000 60850
rect 99900 60620 100000 60650
rect 96000 60600 96120 60620
rect 96380 60600 96620 60620
rect 96880 60600 97120 60620
rect 97380 60600 97620 60620
rect 97880 60600 98120 60620
rect 98380 60600 98620 60620
rect 98880 60600 99120 60620
rect 99380 60600 99620 60620
rect 99880 60600 100000 60620
rect 96000 60590 100000 60600
rect 96000 60520 96150 60590
rect 96350 60520 96650 60590
rect 96850 60520 97150 60590
rect 97350 60520 97650 60590
rect 97850 60520 98150 60590
rect 98350 60520 98650 60590
rect 98850 60520 99150 60590
rect 99350 60520 99650 60590
rect 99850 60520 100000 60590
rect 96000 60480 100000 60520
rect 96000 60410 96150 60480
rect 96350 60410 96650 60480
rect 96850 60410 97150 60480
rect 97350 60410 97650 60480
rect 97850 60410 98150 60480
rect 98350 60410 98650 60480
rect 98850 60410 99150 60480
rect 99350 60410 99650 60480
rect 99850 60410 100000 60480
rect 96000 60400 100000 60410
rect 96000 60380 96120 60400
rect 96380 60380 96620 60400
rect 96880 60380 97120 60400
rect 97380 60380 97620 60400
rect 97880 60380 98120 60400
rect 98380 60380 98620 60400
rect 98880 60380 99120 60400
rect 99380 60380 99620 60400
rect 99880 60380 100000 60400
rect 96000 60350 96100 60380
rect 96000 60150 96020 60350
rect 96090 60150 96100 60350
rect 96000 60120 96100 60150
rect 96400 60350 96600 60380
rect 96400 60150 96410 60350
rect 96480 60150 96520 60350
rect 96590 60150 96600 60350
rect 96400 60120 96600 60150
rect 96900 60350 97100 60380
rect 96900 60150 96910 60350
rect 96980 60150 97020 60350
rect 97090 60150 97100 60350
rect 96900 60120 97100 60150
rect 97400 60350 97600 60380
rect 97400 60150 97410 60350
rect 97480 60150 97520 60350
rect 97590 60150 97600 60350
rect 97400 60120 97600 60150
rect 97900 60350 98100 60380
rect 97900 60150 97910 60350
rect 97980 60150 98020 60350
rect 98090 60150 98100 60350
rect 97900 60120 98100 60150
rect 98400 60350 98600 60380
rect 98400 60150 98410 60350
rect 98480 60150 98520 60350
rect 98590 60150 98600 60350
rect 98400 60120 98600 60150
rect 98900 60350 99100 60380
rect 98900 60150 98910 60350
rect 98980 60150 99020 60350
rect 99090 60150 99100 60350
rect 98900 60120 99100 60150
rect 99400 60350 99600 60380
rect 99400 60150 99410 60350
rect 99480 60150 99520 60350
rect 99590 60150 99600 60350
rect 99400 60120 99600 60150
rect 99900 60350 100000 60380
rect 99900 60150 99910 60350
rect 99980 60150 100000 60350
rect 99900 60120 100000 60150
rect 96000 60100 96120 60120
rect 96380 60100 96620 60120
rect 96880 60100 97120 60120
rect 97380 60100 97620 60120
rect 97880 60100 98120 60120
rect 98380 60100 98620 60120
rect 98880 60100 99120 60120
rect 99380 60100 99620 60120
rect 99880 60100 100000 60120
rect 96000 60090 100000 60100
rect 96000 60020 96150 60090
rect 96350 60020 96650 60090
rect 96850 60020 97150 60090
rect 97350 60020 97650 60090
rect 97850 60020 98150 60090
rect 98350 60020 98650 60090
rect 98850 60020 99150 60090
rect 99350 60020 99650 60090
rect 99850 60020 100000 60090
rect 96000 59980 100000 60020
rect 96000 59910 96150 59980
rect 96350 59910 96650 59980
rect 96850 59910 97150 59980
rect 97350 59910 97650 59980
rect 97850 59910 98150 59980
rect 98350 59910 98650 59980
rect 98850 59910 99150 59980
rect 99350 59910 99650 59980
rect 99850 59910 100000 59980
rect 96000 59900 100000 59910
rect 96000 59880 96120 59900
rect 96380 59880 96620 59900
rect 96880 59880 97120 59900
rect 97380 59880 97620 59900
rect 97880 59880 98120 59900
rect 98380 59880 98620 59900
rect 98880 59880 99120 59900
rect 99380 59880 99620 59900
rect 99880 59880 100000 59900
rect 96000 59850 96100 59880
rect 96000 59650 96020 59850
rect 96090 59650 96100 59850
rect 96000 59620 96100 59650
rect 96400 59850 96600 59880
rect 96400 59650 96410 59850
rect 96480 59650 96520 59850
rect 96590 59650 96600 59850
rect 96400 59620 96600 59650
rect 96900 59850 97100 59880
rect 96900 59650 96910 59850
rect 96980 59650 97020 59850
rect 97090 59650 97100 59850
rect 96900 59620 97100 59650
rect 97400 59850 97600 59880
rect 97400 59650 97410 59850
rect 97480 59650 97520 59850
rect 97590 59650 97600 59850
rect 97400 59620 97600 59650
rect 97900 59850 98100 59880
rect 97900 59650 97910 59850
rect 97980 59650 98020 59850
rect 98090 59650 98100 59850
rect 97900 59620 98100 59650
rect 98400 59850 98600 59880
rect 98400 59650 98410 59850
rect 98480 59650 98520 59850
rect 98590 59650 98600 59850
rect 98400 59620 98600 59650
rect 98900 59850 99100 59880
rect 98900 59650 98910 59850
rect 98980 59650 99020 59850
rect 99090 59650 99100 59850
rect 98900 59620 99100 59650
rect 99400 59850 99600 59880
rect 99400 59650 99410 59850
rect 99480 59650 99520 59850
rect 99590 59650 99600 59850
rect 99400 59620 99600 59650
rect 99900 59850 100000 59880
rect 99900 59650 99910 59850
rect 99980 59650 100000 59850
rect 99900 59620 100000 59650
rect 96000 59600 96120 59620
rect 96380 59600 96620 59620
rect 96880 59600 97120 59620
rect 97380 59600 97620 59620
rect 97880 59600 98120 59620
rect 98380 59600 98620 59620
rect 98880 59600 99120 59620
rect 99380 59600 99620 59620
rect 99880 59600 100000 59620
rect 96000 59590 100000 59600
rect 96000 59520 96150 59590
rect 96350 59520 96650 59590
rect 96850 59520 97150 59590
rect 97350 59520 97650 59590
rect 97850 59520 98150 59590
rect 98350 59520 98650 59590
rect 98850 59520 99150 59590
rect 99350 59520 99650 59590
rect 99850 59520 100000 59590
rect 96000 59480 100000 59520
rect 96000 59410 96150 59480
rect 96350 59410 96650 59480
rect 96850 59410 97150 59480
rect 97350 59410 97650 59480
rect 97850 59410 98150 59480
rect 98350 59410 98650 59480
rect 98850 59410 99150 59480
rect 99350 59410 99650 59480
rect 99850 59410 100000 59480
rect 96000 59400 100000 59410
rect 96000 59380 96120 59400
rect 96380 59380 96620 59400
rect 96880 59380 97120 59400
rect 97380 59380 97620 59400
rect 97880 59380 98120 59400
rect 98380 59380 98620 59400
rect 98880 59380 99120 59400
rect 99380 59380 99620 59400
rect 99880 59380 100000 59400
rect 96000 59350 96100 59380
rect 96000 59150 96020 59350
rect 96090 59150 96100 59350
rect 96000 59120 96100 59150
rect 96400 59350 96600 59380
rect 96400 59150 96410 59350
rect 96480 59150 96520 59350
rect 96590 59150 96600 59350
rect 96400 59120 96600 59150
rect 96900 59350 97100 59380
rect 96900 59150 96910 59350
rect 96980 59150 97020 59350
rect 97090 59150 97100 59350
rect 96900 59120 97100 59150
rect 97400 59350 97600 59380
rect 97400 59150 97410 59350
rect 97480 59150 97520 59350
rect 97590 59150 97600 59350
rect 97400 59120 97600 59150
rect 97900 59350 98100 59380
rect 97900 59150 97910 59350
rect 97980 59150 98020 59350
rect 98090 59150 98100 59350
rect 97900 59120 98100 59150
rect 98400 59350 98600 59380
rect 98400 59150 98410 59350
rect 98480 59150 98520 59350
rect 98590 59150 98600 59350
rect 98400 59120 98600 59150
rect 98900 59350 99100 59380
rect 98900 59150 98910 59350
rect 98980 59150 99020 59350
rect 99090 59150 99100 59350
rect 98900 59120 99100 59150
rect 99400 59350 99600 59380
rect 99400 59150 99410 59350
rect 99480 59150 99520 59350
rect 99590 59150 99600 59350
rect 99400 59120 99600 59150
rect 99900 59350 100000 59380
rect 99900 59150 99910 59350
rect 99980 59150 100000 59350
rect 99900 59120 100000 59150
rect 96000 59100 96120 59120
rect 96380 59100 96620 59120
rect 96880 59100 97120 59120
rect 97380 59100 97620 59120
rect 97880 59100 98120 59120
rect 98380 59100 98620 59120
rect 98880 59100 99120 59120
rect 99380 59100 99620 59120
rect 99880 59100 100000 59120
rect 96000 59090 100000 59100
rect 96000 59020 96150 59090
rect 96350 59020 96650 59090
rect 96850 59020 97150 59090
rect 97350 59020 97650 59090
rect 97850 59020 98150 59090
rect 98350 59020 98650 59090
rect 98850 59020 99150 59090
rect 99350 59020 99650 59090
rect 99850 59020 100000 59090
rect 96000 58980 100000 59020
rect 96000 58910 96150 58980
rect 96350 58910 96650 58980
rect 96850 58910 97150 58980
rect 97350 58910 97650 58980
rect 97850 58910 98150 58980
rect 98350 58910 98650 58980
rect 98850 58910 99150 58980
rect 99350 58910 99650 58980
rect 99850 58910 100000 58980
rect 96000 58900 100000 58910
rect 96000 58880 96120 58900
rect 96380 58880 96620 58900
rect 96880 58880 97120 58900
rect 97380 58880 97620 58900
rect 97880 58880 98120 58900
rect 98380 58880 98620 58900
rect 98880 58880 99120 58900
rect 99380 58880 99620 58900
rect 99880 58880 100000 58900
rect 96000 58850 96100 58880
rect 96000 58650 96020 58850
rect 96090 58650 96100 58850
rect 96000 58620 96100 58650
rect 96400 58850 96600 58880
rect 96400 58650 96410 58850
rect 96480 58650 96520 58850
rect 96590 58650 96600 58850
rect 96400 58620 96600 58650
rect 96900 58850 97100 58880
rect 96900 58650 96910 58850
rect 96980 58650 97020 58850
rect 97090 58650 97100 58850
rect 96900 58620 97100 58650
rect 97400 58850 97600 58880
rect 97400 58650 97410 58850
rect 97480 58650 97520 58850
rect 97590 58650 97600 58850
rect 97400 58620 97600 58650
rect 97900 58850 98100 58880
rect 97900 58650 97910 58850
rect 97980 58650 98020 58850
rect 98090 58650 98100 58850
rect 97900 58620 98100 58650
rect 98400 58850 98600 58880
rect 98400 58650 98410 58850
rect 98480 58650 98520 58850
rect 98590 58650 98600 58850
rect 98400 58620 98600 58650
rect 98900 58850 99100 58880
rect 98900 58650 98910 58850
rect 98980 58650 99020 58850
rect 99090 58650 99100 58850
rect 98900 58620 99100 58650
rect 99400 58850 99600 58880
rect 99400 58650 99410 58850
rect 99480 58650 99520 58850
rect 99590 58650 99600 58850
rect 99400 58620 99600 58650
rect 99900 58850 100000 58880
rect 99900 58650 99910 58850
rect 99980 58650 100000 58850
rect 99900 58620 100000 58650
rect 96000 58600 96120 58620
rect 96380 58600 96620 58620
rect 96880 58600 97120 58620
rect 97380 58600 97620 58620
rect 97880 58600 98120 58620
rect 98380 58600 98620 58620
rect 98880 58600 99120 58620
rect 99380 58600 99620 58620
rect 99880 58600 100000 58620
rect 96000 58590 100000 58600
rect 96000 58520 96150 58590
rect 96350 58520 96650 58590
rect 96850 58520 97150 58590
rect 97350 58520 97650 58590
rect 97850 58520 98150 58590
rect 98350 58520 98650 58590
rect 98850 58520 99150 58590
rect 99350 58520 99650 58590
rect 99850 58520 100000 58590
rect 96000 58480 100000 58520
rect 96000 58410 96150 58480
rect 96350 58410 96650 58480
rect 96850 58410 97150 58480
rect 97350 58410 97650 58480
rect 97850 58410 98150 58480
rect 98350 58410 98650 58480
rect 98850 58410 99150 58480
rect 99350 58410 99650 58480
rect 99850 58410 100000 58480
rect 96000 58400 100000 58410
rect 96000 58380 96120 58400
rect 96380 58380 96620 58400
rect 96880 58380 97120 58400
rect 97380 58380 97620 58400
rect 97880 58380 98120 58400
rect 98380 58380 98620 58400
rect 98880 58380 99120 58400
rect 99380 58380 99620 58400
rect 99880 58380 100000 58400
rect 96000 58350 96100 58380
rect 96000 58150 96020 58350
rect 96090 58150 96100 58350
rect 96000 58120 96100 58150
rect 96400 58350 96600 58380
rect 96400 58150 96410 58350
rect 96480 58150 96520 58350
rect 96590 58150 96600 58350
rect 96400 58120 96600 58150
rect 96900 58350 97100 58380
rect 96900 58150 96910 58350
rect 96980 58150 97020 58350
rect 97090 58150 97100 58350
rect 96900 58120 97100 58150
rect 97400 58350 97600 58380
rect 97400 58150 97410 58350
rect 97480 58150 97520 58350
rect 97590 58150 97600 58350
rect 97400 58120 97600 58150
rect 97900 58350 98100 58380
rect 97900 58150 97910 58350
rect 97980 58150 98020 58350
rect 98090 58150 98100 58350
rect 97900 58120 98100 58150
rect 98400 58350 98600 58380
rect 98400 58150 98410 58350
rect 98480 58150 98520 58350
rect 98590 58150 98600 58350
rect 98400 58120 98600 58150
rect 98900 58350 99100 58380
rect 98900 58150 98910 58350
rect 98980 58150 99020 58350
rect 99090 58150 99100 58350
rect 98900 58120 99100 58150
rect 99400 58350 99600 58380
rect 99400 58150 99410 58350
rect 99480 58150 99520 58350
rect 99590 58150 99600 58350
rect 99400 58120 99600 58150
rect 99900 58350 100000 58380
rect 99900 58150 99910 58350
rect 99980 58150 100000 58350
rect 99900 58120 100000 58150
rect 96000 58100 96120 58120
rect 96380 58100 96620 58120
rect 96880 58100 97120 58120
rect 97380 58100 97620 58120
rect 97880 58100 98120 58120
rect 98380 58100 98620 58120
rect 98880 58100 99120 58120
rect 99380 58100 99620 58120
rect 99880 58100 100000 58120
rect 96000 58090 100000 58100
rect 96000 58020 96150 58090
rect 96350 58020 96650 58090
rect 96850 58020 97150 58090
rect 97350 58020 97650 58090
rect 97850 58020 98150 58090
rect 98350 58020 98650 58090
rect 98850 58020 99150 58090
rect 99350 58020 99650 58090
rect 99850 58020 100000 58090
rect 96000 57980 100000 58020
rect 96000 57910 96150 57980
rect 96350 57910 96650 57980
rect 96850 57910 97150 57980
rect 97350 57910 97650 57980
rect 97850 57910 98150 57980
rect 98350 57910 98650 57980
rect 98850 57910 99150 57980
rect 99350 57910 99650 57980
rect 99850 57910 100000 57980
rect 96000 57900 100000 57910
rect 96000 57880 96120 57900
rect 96380 57880 96620 57900
rect 96880 57880 97120 57900
rect 97380 57880 97620 57900
rect 97880 57880 98120 57900
rect 98380 57880 98620 57900
rect 98880 57880 99120 57900
rect 99380 57880 99620 57900
rect 99880 57880 100000 57900
rect 96000 57850 96100 57880
rect 96000 57650 96020 57850
rect 96090 57650 96100 57850
rect 96000 57620 96100 57650
rect 96400 57850 96600 57880
rect 96400 57650 96410 57850
rect 96480 57650 96520 57850
rect 96590 57650 96600 57850
rect 96400 57620 96600 57650
rect 96900 57850 97100 57880
rect 96900 57650 96910 57850
rect 96980 57650 97020 57850
rect 97090 57650 97100 57850
rect 96900 57620 97100 57650
rect 97400 57850 97600 57880
rect 97400 57650 97410 57850
rect 97480 57650 97520 57850
rect 97590 57650 97600 57850
rect 97400 57620 97600 57650
rect 97900 57850 98100 57880
rect 97900 57650 97910 57850
rect 97980 57650 98020 57850
rect 98090 57650 98100 57850
rect 97900 57620 98100 57650
rect 98400 57850 98600 57880
rect 98400 57650 98410 57850
rect 98480 57650 98520 57850
rect 98590 57650 98600 57850
rect 98400 57620 98600 57650
rect 98900 57850 99100 57880
rect 98900 57650 98910 57850
rect 98980 57650 99020 57850
rect 99090 57650 99100 57850
rect 98900 57620 99100 57650
rect 99400 57850 99600 57880
rect 99400 57650 99410 57850
rect 99480 57650 99520 57850
rect 99590 57650 99600 57850
rect 99400 57620 99600 57650
rect 99900 57850 100000 57880
rect 99900 57650 99910 57850
rect 99980 57650 100000 57850
rect 99900 57620 100000 57650
rect 96000 57600 96120 57620
rect 96380 57600 96620 57620
rect 96880 57600 97120 57620
rect 97380 57600 97620 57620
rect 97880 57600 98120 57620
rect 98380 57600 98620 57620
rect 98880 57600 99120 57620
rect 99380 57600 99620 57620
rect 99880 57600 100000 57620
rect 96000 57590 100000 57600
rect 96000 57520 96150 57590
rect 96350 57520 96650 57590
rect 96850 57520 97150 57590
rect 97350 57520 97650 57590
rect 97850 57520 98150 57590
rect 98350 57520 98650 57590
rect 98850 57520 99150 57590
rect 99350 57520 99650 57590
rect 99850 57520 100000 57590
rect 96000 57480 100000 57520
rect 96000 57410 96150 57480
rect 96350 57410 96650 57480
rect 96850 57410 97150 57480
rect 97350 57410 97650 57480
rect 97850 57410 98150 57480
rect 98350 57410 98650 57480
rect 98850 57410 99150 57480
rect 99350 57410 99650 57480
rect 99850 57410 100000 57480
rect 96000 57400 100000 57410
rect 96000 57380 96120 57400
rect 96380 57380 96620 57400
rect 96880 57380 97120 57400
rect 97380 57380 97620 57400
rect 97880 57380 98120 57400
rect 98380 57380 98620 57400
rect 98880 57380 99120 57400
rect 99380 57380 99620 57400
rect 99880 57380 100000 57400
rect 96000 57350 96100 57380
rect 96000 57150 96020 57350
rect 96090 57150 96100 57350
rect 96000 57120 96100 57150
rect 96400 57350 96600 57380
rect 96400 57150 96410 57350
rect 96480 57150 96520 57350
rect 96590 57150 96600 57350
rect 96400 57120 96600 57150
rect 96900 57350 97100 57380
rect 96900 57150 96910 57350
rect 96980 57150 97020 57350
rect 97090 57150 97100 57350
rect 96900 57120 97100 57150
rect 97400 57350 97600 57380
rect 97400 57150 97410 57350
rect 97480 57150 97520 57350
rect 97590 57150 97600 57350
rect 97400 57120 97600 57150
rect 97900 57350 98100 57380
rect 97900 57150 97910 57350
rect 97980 57150 98020 57350
rect 98090 57150 98100 57350
rect 97900 57120 98100 57150
rect 98400 57350 98600 57380
rect 98400 57150 98410 57350
rect 98480 57150 98520 57350
rect 98590 57150 98600 57350
rect 98400 57120 98600 57150
rect 98900 57350 99100 57380
rect 98900 57150 98910 57350
rect 98980 57150 99020 57350
rect 99090 57150 99100 57350
rect 98900 57120 99100 57150
rect 99400 57350 99600 57380
rect 99400 57150 99410 57350
rect 99480 57150 99520 57350
rect 99590 57150 99600 57350
rect 99400 57120 99600 57150
rect 99900 57350 100000 57380
rect 99900 57150 99910 57350
rect 99980 57150 100000 57350
rect 99900 57120 100000 57150
rect 96000 57100 96120 57120
rect 96380 57100 96620 57120
rect 96880 57100 97120 57120
rect 97380 57100 97620 57120
rect 97880 57100 98120 57120
rect 98380 57100 98620 57120
rect 98880 57100 99120 57120
rect 99380 57100 99620 57120
rect 99880 57100 100000 57120
rect 96000 57090 100000 57100
rect 96000 57020 96150 57090
rect 96350 57020 96650 57090
rect 96850 57020 97150 57090
rect 97350 57020 97650 57090
rect 97850 57020 98150 57090
rect 98350 57020 98650 57090
rect 98850 57020 99150 57090
rect 99350 57020 99650 57090
rect 99850 57020 100000 57090
rect 96000 56980 100000 57020
rect 96000 56910 96150 56980
rect 96350 56910 96650 56980
rect 96850 56910 97150 56980
rect 97350 56910 97650 56980
rect 97850 56910 98150 56980
rect 98350 56910 98650 56980
rect 98850 56910 99150 56980
rect 99350 56910 99650 56980
rect 99850 56910 100000 56980
rect 96000 56900 100000 56910
rect 96000 56880 96120 56900
rect 96380 56880 96620 56900
rect 96880 56880 97120 56900
rect 97380 56880 97620 56900
rect 97880 56880 98120 56900
rect 98380 56880 98620 56900
rect 98880 56880 99120 56900
rect 99380 56880 99620 56900
rect 99880 56880 100000 56900
rect 96000 56850 96100 56880
rect 96000 56650 96020 56850
rect 96090 56650 96100 56850
rect 96000 56620 96100 56650
rect 96400 56850 96600 56880
rect 96400 56650 96410 56850
rect 96480 56650 96520 56850
rect 96590 56650 96600 56850
rect 96400 56620 96600 56650
rect 96900 56850 97100 56880
rect 96900 56650 96910 56850
rect 96980 56650 97020 56850
rect 97090 56650 97100 56850
rect 96900 56620 97100 56650
rect 97400 56850 97600 56880
rect 97400 56650 97410 56850
rect 97480 56650 97520 56850
rect 97590 56650 97600 56850
rect 97400 56620 97600 56650
rect 97900 56850 98100 56880
rect 97900 56650 97910 56850
rect 97980 56650 98020 56850
rect 98090 56650 98100 56850
rect 97900 56620 98100 56650
rect 98400 56850 98600 56880
rect 98400 56650 98410 56850
rect 98480 56650 98520 56850
rect 98590 56650 98600 56850
rect 98400 56620 98600 56650
rect 98900 56850 99100 56880
rect 98900 56650 98910 56850
rect 98980 56650 99020 56850
rect 99090 56650 99100 56850
rect 98900 56620 99100 56650
rect 99400 56850 99600 56880
rect 99400 56650 99410 56850
rect 99480 56650 99520 56850
rect 99590 56650 99600 56850
rect 99400 56620 99600 56650
rect 99900 56850 100000 56880
rect 99900 56650 99910 56850
rect 99980 56650 100000 56850
rect 99900 56620 100000 56650
rect 96000 56600 96120 56620
rect 96380 56600 96620 56620
rect 96880 56600 97120 56620
rect 97380 56600 97620 56620
rect 97880 56600 98120 56620
rect 98380 56600 98620 56620
rect 98880 56600 99120 56620
rect 99380 56600 99620 56620
rect 99880 56600 100000 56620
rect 96000 56590 100000 56600
rect 96000 56520 96150 56590
rect 96350 56520 96650 56590
rect 96850 56520 97150 56590
rect 97350 56520 97650 56590
rect 97850 56520 98150 56590
rect 98350 56520 98650 56590
rect 98850 56520 99150 56590
rect 99350 56520 99650 56590
rect 99850 56520 100000 56590
rect 96000 56480 100000 56520
rect 96000 56410 96150 56480
rect 96350 56410 96650 56480
rect 96850 56410 97150 56480
rect 97350 56410 97650 56480
rect 97850 56410 98150 56480
rect 98350 56410 98650 56480
rect 98850 56410 99150 56480
rect 99350 56410 99650 56480
rect 99850 56410 100000 56480
rect 96000 56400 100000 56410
rect 96000 56380 96120 56400
rect 96380 56380 96620 56400
rect 96880 56380 97120 56400
rect 97380 56380 97620 56400
rect 97880 56380 98120 56400
rect 98380 56380 98620 56400
rect 98880 56380 99120 56400
rect 99380 56380 99620 56400
rect 99880 56380 100000 56400
rect 96000 56350 96100 56380
rect 96000 56150 96020 56350
rect 96090 56150 96100 56350
rect 96000 56120 96100 56150
rect 96400 56350 96600 56380
rect 96400 56150 96410 56350
rect 96480 56150 96520 56350
rect 96590 56150 96600 56350
rect 96400 56120 96600 56150
rect 96900 56350 97100 56380
rect 96900 56150 96910 56350
rect 96980 56150 97020 56350
rect 97090 56150 97100 56350
rect 96900 56120 97100 56150
rect 97400 56350 97600 56380
rect 97400 56150 97410 56350
rect 97480 56150 97520 56350
rect 97590 56150 97600 56350
rect 97400 56120 97600 56150
rect 97900 56350 98100 56380
rect 97900 56150 97910 56350
rect 97980 56150 98020 56350
rect 98090 56150 98100 56350
rect 97900 56120 98100 56150
rect 98400 56350 98600 56380
rect 98400 56150 98410 56350
rect 98480 56150 98520 56350
rect 98590 56150 98600 56350
rect 98400 56120 98600 56150
rect 98900 56350 99100 56380
rect 98900 56150 98910 56350
rect 98980 56150 99020 56350
rect 99090 56150 99100 56350
rect 98900 56120 99100 56150
rect 99400 56350 99600 56380
rect 99400 56150 99410 56350
rect 99480 56150 99520 56350
rect 99590 56150 99600 56350
rect 99400 56120 99600 56150
rect 99900 56350 100000 56380
rect 99900 56150 99910 56350
rect 99980 56150 100000 56350
rect 99900 56120 100000 56150
rect 96000 56100 96120 56120
rect 96380 56100 96620 56120
rect 96880 56100 97120 56120
rect 97380 56100 97620 56120
rect 97880 56100 98120 56120
rect 98380 56100 98620 56120
rect 98880 56100 99120 56120
rect 99380 56100 99620 56120
rect 99880 56100 100000 56120
rect 96000 56090 100000 56100
rect 96000 56020 96150 56090
rect 96350 56020 96650 56090
rect 96850 56020 97150 56090
rect 97350 56020 97650 56090
rect 97850 56020 98150 56090
rect 98350 56020 98650 56090
rect 98850 56020 99150 56090
rect 99350 56020 99650 56090
rect 99850 56020 100000 56090
rect 96000 55980 100000 56020
rect 96000 55910 96150 55980
rect 96350 55910 96650 55980
rect 96850 55910 97150 55980
rect 97350 55910 97650 55980
rect 97850 55910 98150 55980
rect 98350 55910 98650 55980
rect 98850 55910 99150 55980
rect 99350 55910 99650 55980
rect 99850 55910 100000 55980
rect 96000 55900 100000 55910
rect 96000 55880 96120 55900
rect 96380 55880 96620 55900
rect 96880 55880 97120 55900
rect 97380 55880 97620 55900
rect 97880 55880 98120 55900
rect 98380 55880 98620 55900
rect 98880 55880 99120 55900
rect 99380 55880 99620 55900
rect 99880 55880 100000 55900
rect 96000 55850 96100 55880
rect 96000 55650 96020 55850
rect 96090 55650 96100 55850
rect 96000 55620 96100 55650
rect 96400 55850 96600 55880
rect 96400 55650 96410 55850
rect 96480 55650 96520 55850
rect 96590 55650 96600 55850
rect 96400 55620 96600 55650
rect 96900 55850 97100 55880
rect 96900 55650 96910 55850
rect 96980 55650 97020 55850
rect 97090 55650 97100 55850
rect 96900 55620 97100 55650
rect 97400 55850 97600 55880
rect 97400 55650 97410 55850
rect 97480 55650 97520 55850
rect 97590 55650 97600 55850
rect 97400 55620 97600 55650
rect 97900 55850 98100 55880
rect 97900 55650 97910 55850
rect 97980 55650 98020 55850
rect 98090 55650 98100 55850
rect 97900 55620 98100 55650
rect 98400 55850 98600 55880
rect 98400 55650 98410 55850
rect 98480 55650 98520 55850
rect 98590 55650 98600 55850
rect 98400 55620 98600 55650
rect 98900 55850 99100 55880
rect 98900 55650 98910 55850
rect 98980 55650 99020 55850
rect 99090 55650 99100 55850
rect 98900 55620 99100 55650
rect 99400 55850 99600 55880
rect 99400 55650 99410 55850
rect 99480 55650 99520 55850
rect 99590 55650 99600 55850
rect 99400 55620 99600 55650
rect 99900 55850 100000 55880
rect 99900 55650 99910 55850
rect 99980 55650 100000 55850
rect 99900 55620 100000 55650
rect 96000 55600 96120 55620
rect 96380 55600 96620 55620
rect 96880 55600 97120 55620
rect 97380 55600 97620 55620
rect 97880 55600 98120 55620
rect 98380 55600 98620 55620
rect 98880 55600 99120 55620
rect 99380 55600 99620 55620
rect 99880 55600 100000 55620
rect 96000 55590 100000 55600
rect 96000 55520 96150 55590
rect 96350 55520 96650 55590
rect 96850 55520 97150 55590
rect 97350 55520 97650 55590
rect 97850 55520 98150 55590
rect 98350 55520 98650 55590
rect 98850 55520 99150 55590
rect 99350 55520 99650 55590
rect 99850 55520 100000 55590
rect 96000 55480 100000 55520
rect 96000 55410 96150 55480
rect 96350 55410 96650 55480
rect 96850 55410 97150 55480
rect 97350 55410 97650 55480
rect 97850 55410 98150 55480
rect 98350 55410 98650 55480
rect 98850 55410 99150 55480
rect 99350 55410 99650 55480
rect 99850 55410 100000 55480
rect 96000 55400 100000 55410
rect 96000 55380 96120 55400
rect 96380 55380 96620 55400
rect 96880 55380 97120 55400
rect 97380 55380 97620 55400
rect 97880 55380 98120 55400
rect 98380 55380 98620 55400
rect 98880 55380 99120 55400
rect 99380 55380 99620 55400
rect 99880 55380 100000 55400
rect 96000 55350 96100 55380
rect 96000 55150 96020 55350
rect 96090 55150 96100 55350
rect 96000 55120 96100 55150
rect 96400 55350 96600 55380
rect 96400 55150 96410 55350
rect 96480 55150 96520 55350
rect 96590 55150 96600 55350
rect 96400 55120 96600 55150
rect 96900 55350 97100 55380
rect 96900 55150 96910 55350
rect 96980 55150 97020 55350
rect 97090 55150 97100 55350
rect 96900 55120 97100 55150
rect 97400 55350 97600 55380
rect 97400 55150 97410 55350
rect 97480 55150 97520 55350
rect 97590 55150 97600 55350
rect 97400 55120 97600 55150
rect 97900 55350 98100 55380
rect 97900 55150 97910 55350
rect 97980 55150 98020 55350
rect 98090 55150 98100 55350
rect 97900 55120 98100 55150
rect 98400 55350 98600 55380
rect 98400 55150 98410 55350
rect 98480 55150 98520 55350
rect 98590 55150 98600 55350
rect 98400 55120 98600 55150
rect 98900 55350 99100 55380
rect 98900 55150 98910 55350
rect 98980 55150 99020 55350
rect 99090 55150 99100 55350
rect 98900 55120 99100 55150
rect 99400 55350 99600 55380
rect 99400 55150 99410 55350
rect 99480 55150 99520 55350
rect 99590 55150 99600 55350
rect 99400 55120 99600 55150
rect 99900 55350 100000 55380
rect 99900 55150 99910 55350
rect 99980 55150 100000 55350
rect 99900 55120 100000 55150
rect 96000 55100 96120 55120
rect 96380 55100 96620 55120
rect 96880 55100 97120 55120
rect 97380 55100 97620 55120
rect 97880 55100 98120 55120
rect 98380 55100 98620 55120
rect 98880 55100 99120 55120
rect 99380 55100 99620 55120
rect 99880 55100 100000 55120
rect 96000 55090 100000 55100
rect 96000 55020 96150 55090
rect 96350 55020 96650 55090
rect 96850 55020 97150 55090
rect 97350 55020 97650 55090
rect 97850 55020 98150 55090
rect 98350 55020 98650 55090
rect 98850 55020 99150 55090
rect 99350 55020 99650 55090
rect 99850 55020 100000 55090
rect 96000 54980 100000 55020
rect 96000 54910 96150 54980
rect 96350 54910 96650 54980
rect 96850 54910 97150 54980
rect 97350 54910 97650 54980
rect 97850 54910 98150 54980
rect 98350 54910 98650 54980
rect 98850 54910 99150 54980
rect 99350 54910 99650 54980
rect 99850 54910 100000 54980
rect 96000 54900 100000 54910
rect 96000 54880 96120 54900
rect 96380 54880 96620 54900
rect 96880 54880 97120 54900
rect 97380 54880 97620 54900
rect 97880 54880 98120 54900
rect 98380 54880 98620 54900
rect 98880 54880 99120 54900
rect 99380 54880 99620 54900
rect 99880 54880 100000 54900
rect 96000 54850 96100 54880
rect 96000 54650 96020 54850
rect 96090 54650 96100 54850
rect 96000 54620 96100 54650
rect 96400 54850 96600 54880
rect 96400 54650 96410 54850
rect 96480 54650 96520 54850
rect 96590 54650 96600 54850
rect 96400 54620 96600 54650
rect 96900 54850 97100 54880
rect 96900 54650 96910 54850
rect 96980 54650 97020 54850
rect 97090 54650 97100 54850
rect 96900 54620 97100 54650
rect 97400 54850 97600 54880
rect 97400 54650 97410 54850
rect 97480 54650 97520 54850
rect 97590 54650 97600 54850
rect 97400 54620 97600 54650
rect 97900 54850 98100 54880
rect 97900 54650 97910 54850
rect 97980 54650 98020 54850
rect 98090 54650 98100 54850
rect 97900 54620 98100 54650
rect 98400 54850 98600 54880
rect 98400 54650 98410 54850
rect 98480 54650 98520 54850
rect 98590 54650 98600 54850
rect 98400 54620 98600 54650
rect 98900 54850 99100 54880
rect 98900 54650 98910 54850
rect 98980 54650 99020 54850
rect 99090 54650 99100 54850
rect 98900 54620 99100 54650
rect 99400 54850 99600 54880
rect 99400 54650 99410 54850
rect 99480 54650 99520 54850
rect 99590 54650 99600 54850
rect 99400 54620 99600 54650
rect 99900 54850 100000 54880
rect 99900 54650 99910 54850
rect 99980 54650 100000 54850
rect 99900 54620 100000 54650
rect 96000 54600 96120 54620
rect 96380 54600 96620 54620
rect 96880 54600 97120 54620
rect 97380 54600 97620 54620
rect 97880 54600 98120 54620
rect 98380 54600 98620 54620
rect 98880 54600 99120 54620
rect 99380 54600 99620 54620
rect 99880 54600 100000 54620
rect 96000 54590 100000 54600
rect 96000 54520 96150 54590
rect 96350 54520 96650 54590
rect 96850 54520 97150 54590
rect 97350 54520 97650 54590
rect 97850 54520 98150 54590
rect 98350 54520 98650 54590
rect 98850 54520 99150 54590
rect 99350 54520 99650 54590
rect 99850 54520 100000 54590
rect 96000 54480 100000 54520
rect 96000 54410 96150 54480
rect 96350 54410 96650 54480
rect 96850 54410 97150 54480
rect 97350 54410 97650 54480
rect 97850 54410 98150 54480
rect 98350 54410 98650 54480
rect 98850 54410 99150 54480
rect 99350 54410 99650 54480
rect 99850 54410 100000 54480
rect 96000 54400 100000 54410
rect 96000 54380 96120 54400
rect 96380 54380 96620 54400
rect 96880 54380 97120 54400
rect 97380 54380 97620 54400
rect 97880 54380 98120 54400
rect 98380 54380 98620 54400
rect 98880 54380 99120 54400
rect 99380 54380 99620 54400
rect 99880 54380 100000 54400
rect 96000 54350 96100 54380
rect 96000 54150 96020 54350
rect 96090 54150 96100 54350
rect 96000 54120 96100 54150
rect 96400 54350 96600 54380
rect 96400 54150 96410 54350
rect 96480 54150 96520 54350
rect 96590 54150 96600 54350
rect 96400 54120 96600 54150
rect 96900 54350 97100 54380
rect 96900 54150 96910 54350
rect 96980 54150 97020 54350
rect 97090 54150 97100 54350
rect 96900 54120 97100 54150
rect 97400 54350 97600 54380
rect 97400 54150 97410 54350
rect 97480 54150 97520 54350
rect 97590 54150 97600 54350
rect 97400 54120 97600 54150
rect 97900 54350 98100 54380
rect 97900 54150 97910 54350
rect 97980 54150 98020 54350
rect 98090 54150 98100 54350
rect 97900 54120 98100 54150
rect 98400 54350 98600 54380
rect 98400 54150 98410 54350
rect 98480 54150 98520 54350
rect 98590 54150 98600 54350
rect 98400 54120 98600 54150
rect 98900 54350 99100 54380
rect 98900 54150 98910 54350
rect 98980 54150 99020 54350
rect 99090 54150 99100 54350
rect 98900 54120 99100 54150
rect 99400 54350 99600 54380
rect 99400 54150 99410 54350
rect 99480 54150 99520 54350
rect 99590 54150 99600 54350
rect 99400 54120 99600 54150
rect 99900 54350 100000 54380
rect 99900 54150 99910 54350
rect 99980 54150 100000 54350
rect 99900 54120 100000 54150
rect 96000 54100 96120 54120
rect 96380 54100 96620 54120
rect 96880 54100 97120 54120
rect 97380 54100 97620 54120
rect 97880 54100 98120 54120
rect 98380 54100 98620 54120
rect 98880 54100 99120 54120
rect 99380 54100 99620 54120
rect 99880 54100 100000 54120
rect 96000 54090 100000 54100
rect 96000 54020 96150 54090
rect 96350 54020 96650 54090
rect 96850 54020 97150 54090
rect 97350 54020 97650 54090
rect 97850 54020 98150 54090
rect 98350 54020 98650 54090
rect 98850 54020 99150 54090
rect 99350 54020 99650 54090
rect 99850 54020 100000 54090
rect 96000 53980 100000 54020
rect 96000 53910 96150 53980
rect 96350 53910 96650 53980
rect 96850 53910 97150 53980
rect 97350 53910 97650 53980
rect 97850 53910 98150 53980
rect 98350 53910 98650 53980
rect 98850 53910 99150 53980
rect 99350 53910 99650 53980
rect 99850 53910 100000 53980
rect 96000 53900 100000 53910
rect 96000 53880 96120 53900
rect 96380 53880 96620 53900
rect 96880 53880 97120 53900
rect 97380 53880 97620 53900
rect 97880 53880 98120 53900
rect 98380 53880 98620 53900
rect 98880 53880 99120 53900
rect 99380 53880 99620 53900
rect 99880 53880 100000 53900
rect 96000 53850 96100 53880
rect 96000 53650 96020 53850
rect 96090 53650 96100 53850
rect 96000 53620 96100 53650
rect 96400 53850 96600 53880
rect 96400 53650 96410 53850
rect 96480 53650 96520 53850
rect 96590 53650 96600 53850
rect 96400 53620 96600 53650
rect 96900 53850 97100 53880
rect 96900 53650 96910 53850
rect 96980 53650 97020 53850
rect 97090 53650 97100 53850
rect 96900 53620 97100 53650
rect 97400 53850 97600 53880
rect 97400 53650 97410 53850
rect 97480 53650 97520 53850
rect 97590 53650 97600 53850
rect 97400 53620 97600 53650
rect 97900 53850 98100 53880
rect 97900 53650 97910 53850
rect 97980 53650 98020 53850
rect 98090 53650 98100 53850
rect 97900 53620 98100 53650
rect 98400 53850 98600 53880
rect 98400 53650 98410 53850
rect 98480 53650 98520 53850
rect 98590 53650 98600 53850
rect 98400 53620 98600 53650
rect 98900 53850 99100 53880
rect 98900 53650 98910 53850
rect 98980 53650 99020 53850
rect 99090 53650 99100 53850
rect 98900 53620 99100 53650
rect 99400 53850 99600 53880
rect 99400 53650 99410 53850
rect 99480 53650 99520 53850
rect 99590 53650 99600 53850
rect 99400 53620 99600 53650
rect 99900 53850 100000 53880
rect 99900 53650 99910 53850
rect 99980 53650 100000 53850
rect 99900 53620 100000 53650
rect 96000 53600 96120 53620
rect 96380 53600 96620 53620
rect 96880 53600 97120 53620
rect 97380 53600 97620 53620
rect 97880 53600 98120 53620
rect 98380 53600 98620 53620
rect 98880 53600 99120 53620
rect 99380 53600 99620 53620
rect 99880 53600 100000 53620
rect 96000 53590 100000 53600
rect 96000 53520 96150 53590
rect 96350 53520 96650 53590
rect 96850 53520 97150 53590
rect 97350 53520 97650 53590
rect 97850 53520 98150 53590
rect 98350 53520 98650 53590
rect 98850 53520 99150 53590
rect 99350 53520 99650 53590
rect 99850 53520 100000 53590
rect 96000 53480 100000 53520
rect 96000 53410 96150 53480
rect 96350 53410 96650 53480
rect 96850 53410 97150 53480
rect 97350 53410 97650 53480
rect 97850 53410 98150 53480
rect 98350 53410 98650 53480
rect 98850 53410 99150 53480
rect 99350 53410 99650 53480
rect 99850 53410 100000 53480
rect 96000 53400 100000 53410
rect 96000 53380 96120 53400
rect 96380 53380 96620 53400
rect 96880 53380 97120 53400
rect 97380 53380 97620 53400
rect 97880 53380 98120 53400
rect 98380 53380 98620 53400
rect 98880 53380 99120 53400
rect 99380 53380 99620 53400
rect 99880 53380 100000 53400
rect 96000 53350 96100 53380
rect 96000 53150 96020 53350
rect 96090 53150 96100 53350
rect 96000 53120 96100 53150
rect 96400 53350 96600 53380
rect 96400 53150 96410 53350
rect 96480 53150 96520 53350
rect 96590 53150 96600 53350
rect 96400 53120 96600 53150
rect 96900 53350 97100 53380
rect 96900 53150 96910 53350
rect 96980 53150 97020 53350
rect 97090 53150 97100 53350
rect 96900 53120 97100 53150
rect 97400 53350 97600 53380
rect 97400 53150 97410 53350
rect 97480 53150 97520 53350
rect 97590 53150 97600 53350
rect 97400 53120 97600 53150
rect 97900 53350 98100 53380
rect 97900 53150 97910 53350
rect 97980 53150 98020 53350
rect 98090 53150 98100 53350
rect 97900 53120 98100 53150
rect 98400 53350 98600 53380
rect 98400 53150 98410 53350
rect 98480 53150 98520 53350
rect 98590 53150 98600 53350
rect 98400 53120 98600 53150
rect 98900 53350 99100 53380
rect 98900 53150 98910 53350
rect 98980 53150 99020 53350
rect 99090 53150 99100 53350
rect 98900 53120 99100 53150
rect 99400 53350 99600 53380
rect 99400 53150 99410 53350
rect 99480 53150 99520 53350
rect 99590 53150 99600 53350
rect 99400 53120 99600 53150
rect 99900 53350 100000 53380
rect 99900 53150 99910 53350
rect 99980 53150 100000 53350
rect 99900 53120 100000 53150
rect 96000 53100 96120 53120
rect 96380 53100 96620 53120
rect 96880 53100 97120 53120
rect 97380 53100 97620 53120
rect 97880 53100 98120 53120
rect 98380 53100 98620 53120
rect 98880 53100 99120 53120
rect 99380 53100 99620 53120
rect 99880 53100 100000 53120
rect 96000 53090 100000 53100
rect 96000 53020 96150 53090
rect 96350 53020 96650 53090
rect 96850 53020 97150 53090
rect 97350 53020 97650 53090
rect 97850 53020 98150 53090
rect 98350 53020 98650 53090
rect 98850 53020 99150 53090
rect 99350 53020 99650 53090
rect 99850 53020 100000 53090
rect 96000 52980 100000 53020
rect 96000 52910 96150 52980
rect 96350 52910 96650 52980
rect 96850 52910 97150 52980
rect 97350 52910 97650 52980
rect 97850 52910 98150 52980
rect 98350 52910 98650 52980
rect 98850 52910 99150 52980
rect 99350 52910 99650 52980
rect 99850 52910 100000 52980
rect 96000 52900 100000 52910
rect 96000 52880 96120 52900
rect 96380 52880 96620 52900
rect 96880 52880 97120 52900
rect 97380 52880 97620 52900
rect 97880 52880 98120 52900
rect 98380 52880 98620 52900
rect 98880 52880 99120 52900
rect 99380 52880 99620 52900
rect 99880 52880 100000 52900
rect 96000 52850 96100 52880
rect 96000 52650 96020 52850
rect 96090 52650 96100 52850
rect 96000 52620 96100 52650
rect 96400 52850 96600 52880
rect 96400 52650 96410 52850
rect 96480 52650 96520 52850
rect 96590 52650 96600 52850
rect 96400 52620 96600 52650
rect 96900 52850 97100 52880
rect 96900 52650 96910 52850
rect 96980 52650 97020 52850
rect 97090 52650 97100 52850
rect 96900 52620 97100 52650
rect 97400 52850 97600 52880
rect 97400 52650 97410 52850
rect 97480 52650 97520 52850
rect 97590 52650 97600 52850
rect 97400 52620 97600 52650
rect 97900 52850 98100 52880
rect 97900 52650 97910 52850
rect 97980 52650 98020 52850
rect 98090 52650 98100 52850
rect 97900 52620 98100 52650
rect 98400 52850 98600 52880
rect 98400 52650 98410 52850
rect 98480 52650 98520 52850
rect 98590 52650 98600 52850
rect 98400 52620 98600 52650
rect 98900 52850 99100 52880
rect 98900 52650 98910 52850
rect 98980 52650 99020 52850
rect 99090 52650 99100 52850
rect 98900 52620 99100 52650
rect 99400 52850 99600 52880
rect 99400 52650 99410 52850
rect 99480 52650 99520 52850
rect 99590 52650 99600 52850
rect 99400 52620 99600 52650
rect 99900 52850 100000 52880
rect 99900 52650 99910 52850
rect 99980 52650 100000 52850
rect 99900 52620 100000 52650
rect 96000 52600 96120 52620
rect 96380 52600 96620 52620
rect 96880 52600 97120 52620
rect 97380 52600 97620 52620
rect 97880 52600 98120 52620
rect 98380 52600 98620 52620
rect 98880 52600 99120 52620
rect 99380 52600 99620 52620
rect 99880 52600 100000 52620
rect 96000 52590 100000 52600
rect 96000 52520 96150 52590
rect 96350 52520 96650 52590
rect 96850 52520 97150 52590
rect 97350 52520 97650 52590
rect 97850 52520 98150 52590
rect 98350 52520 98650 52590
rect 98850 52520 99150 52590
rect 99350 52520 99650 52590
rect 99850 52520 100000 52590
rect 96000 52480 100000 52520
rect 96000 52410 96150 52480
rect 96350 52410 96650 52480
rect 96850 52410 97150 52480
rect 97350 52410 97650 52480
rect 97850 52410 98150 52480
rect 98350 52410 98650 52480
rect 98850 52410 99150 52480
rect 99350 52410 99650 52480
rect 99850 52410 100000 52480
rect 96000 52400 100000 52410
rect 96000 52380 96120 52400
rect 96380 52380 96620 52400
rect 96880 52380 97120 52400
rect 97380 52380 97620 52400
rect 97880 52380 98120 52400
rect 98380 52380 98620 52400
rect 98880 52380 99120 52400
rect 99380 52380 99620 52400
rect 99880 52380 100000 52400
rect 96000 52350 96100 52380
rect 96000 52150 96020 52350
rect 96090 52150 96100 52350
rect 96000 52120 96100 52150
rect 96400 52350 96600 52380
rect 96400 52150 96410 52350
rect 96480 52150 96520 52350
rect 96590 52150 96600 52350
rect 96400 52120 96600 52150
rect 96900 52350 97100 52380
rect 96900 52150 96910 52350
rect 96980 52150 97020 52350
rect 97090 52150 97100 52350
rect 96900 52120 97100 52150
rect 97400 52350 97600 52380
rect 97400 52150 97410 52350
rect 97480 52150 97520 52350
rect 97590 52150 97600 52350
rect 97400 52120 97600 52150
rect 97900 52350 98100 52380
rect 97900 52150 97910 52350
rect 97980 52150 98020 52350
rect 98090 52150 98100 52350
rect 97900 52120 98100 52150
rect 98400 52350 98600 52380
rect 98400 52150 98410 52350
rect 98480 52150 98520 52350
rect 98590 52150 98600 52350
rect 98400 52120 98600 52150
rect 98900 52350 99100 52380
rect 98900 52150 98910 52350
rect 98980 52150 99020 52350
rect 99090 52150 99100 52350
rect 98900 52120 99100 52150
rect 99400 52350 99600 52380
rect 99400 52150 99410 52350
rect 99480 52150 99520 52350
rect 99590 52150 99600 52350
rect 99400 52120 99600 52150
rect 99900 52350 100000 52380
rect 99900 52150 99910 52350
rect 99980 52150 100000 52350
rect 99900 52120 100000 52150
rect 96000 52100 96120 52120
rect 96380 52100 96620 52120
rect 96880 52100 97120 52120
rect 97380 52100 97620 52120
rect 97880 52100 98120 52120
rect 98380 52100 98620 52120
rect 98880 52100 99120 52120
rect 99380 52100 99620 52120
rect 99880 52100 100000 52120
rect 96000 52090 100000 52100
rect 96000 52020 96150 52090
rect 96350 52020 96650 52090
rect 96850 52020 97150 52090
rect 97350 52020 97650 52090
rect 97850 52020 98150 52090
rect 98350 52020 98650 52090
rect 98850 52020 99150 52090
rect 99350 52020 99650 52090
rect 99850 52020 100000 52090
rect 96000 51980 100000 52020
rect 96000 51910 96150 51980
rect 96350 51910 96650 51980
rect 96850 51910 97150 51980
rect 97350 51910 97650 51980
rect 97850 51910 98150 51980
rect 98350 51910 98650 51980
rect 98850 51910 99150 51980
rect 99350 51910 99650 51980
rect 99850 51910 100000 51980
rect 96000 51900 100000 51910
rect 96000 51880 96120 51900
rect 96380 51880 96620 51900
rect 96880 51880 97120 51900
rect 97380 51880 97620 51900
rect 97880 51880 98120 51900
rect 98380 51880 98620 51900
rect 98880 51880 99120 51900
rect 99380 51880 99620 51900
rect 99880 51880 100000 51900
rect 96000 51850 96100 51880
rect 96000 51650 96020 51850
rect 96090 51650 96100 51850
rect 96000 51620 96100 51650
rect 96400 51850 96600 51880
rect 96400 51650 96410 51850
rect 96480 51650 96520 51850
rect 96590 51650 96600 51850
rect 96400 51620 96600 51650
rect 96900 51850 97100 51880
rect 96900 51650 96910 51850
rect 96980 51650 97020 51850
rect 97090 51650 97100 51850
rect 96900 51620 97100 51650
rect 97400 51850 97600 51880
rect 97400 51650 97410 51850
rect 97480 51650 97520 51850
rect 97590 51650 97600 51850
rect 97400 51620 97600 51650
rect 97900 51850 98100 51880
rect 97900 51650 97910 51850
rect 97980 51650 98020 51850
rect 98090 51650 98100 51850
rect 97900 51620 98100 51650
rect 98400 51850 98600 51880
rect 98400 51650 98410 51850
rect 98480 51650 98520 51850
rect 98590 51650 98600 51850
rect 98400 51620 98600 51650
rect 98900 51850 99100 51880
rect 98900 51650 98910 51850
rect 98980 51650 99020 51850
rect 99090 51650 99100 51850
rect 98900 51620 99100 51650
rect 99400 51850 99600 51880
rect 99400 51650 99410 51850
rect 99480 51650 99520 51850
rect 99590 51650 99600 51850
rect 99400 51620 99600 51650
rect 99900 51850 100000 51880
rect 99900 51650 99910 51850
rect 99980 51650 100000 51850
rect 99900 51620 100000 51650
rect 96000 51600 96120 51620
rect 96380 51600 96620 51620
rect 96880 51600 97120 51620
rect 97380 51600 97620 51620
rect 97880 51600 98120 51620
rect 98380 51600 98620 51620
rect 98880 51600 99120 51620
rect 99380 51600 99620 51620
rect 99880 51600 100000 51620
rect 96000 51590 100000 51600
rect 96000 51520 96150 51590
rect 96350 51520 96650 51590
rect 96850 51520 97150 51590
rect 97350 51520 97650 51590
rect 97850 51520 98150 51590
rect 98350 51520 98650 51590
rect 98850 51520 99150 51590
rect 99350 51520 99650 51590
rect 99850 51520 100000 51590
rect 96000 51480 100000 51520
rect 96000 51410 96150 51480
rect 96350 51410 96650 51480
rect 96850 51410 97150 51480
rect 97350 51410 97650 51480
rect 97850 51410 98150 51480
rect 98350 51410 98650 51480
rect 98850 51410 99150 51480
rect 99350 51410 99650 51480
rect 99850 51410 100000 51480
rect 96000 51400 100000 51410
rect 96000 51380 96120 51400
rect 96380 51380 96620 51400
rect 96880 51380 97120 51400
rect 97380 51380 97620 51400
rect 97880 51380 98120 51400
rect 98380 51380 98620 51400
rect 98880 51380 99120 51400
rect 99380 51380 99620 51400
rect 99880 51380 100000 51400
rect 96000 51350 96100 51380
rect 96000 51150 96020 51350
rect 96090 51150 96100 51350
rect 96000 51120 96100 51150
rect 96400 51350 96600 51380
rect 96400 51150 96410 51350
rect 96480 51150 96520 51350
rect 96590 51150 96600 51350
rect 96400 51120 96600 51150
rect 96900 51350 97100 51380
rect 96900 51150 96910 51350
rect 96980 51150 97020 51350
rect 97090 51150 97100 51350
rect 96900 51120 97100 51150
rect 97400 51350 97600 51380
rect 97400 51150 97410 51350
rect 97480 51150 97520 51350
rect 97590 51150 97600 51350
rect 97400 51120 97600 51150
rect 97900 51350 98100 51380
rect 97900 51150 97910 51350
rect 97980 51150 98020 51350
rect 98090 51150 98100 51350
rect 97900 51120 98100 51150
rect 98400 51350 98600 51380
rect 98400 51150 98410 51350
rect 98480 51150 98520 51350
rect 98590 51150 98600 51350
rect 98400 51120 98600 51150
rect 98900 51350 99100 51380
rect 98900 51150 98910 51350
rect 98980 51150 99020 51350
rect 99090 51150 99100 51350
rect 98900 51120 99100 51150
rect 99400 51350 99600 51380
rect 99400 51150 99410 51350
rect 99480 51150 99520 51350
rect 99590 51150 99600 51350
rect 99400 51120 99600 51150
rect 99900 51350 100000 51380
rect 99900 51150 99910 51350
rect 99980 51150 100000 51350
rect 99900 51120 100000 51150
rect 96000 51100 96120 51120
rect 96380 51100 96620 51120
rect 96880 51100 97120 51120
rect 97380 51100 97620 51120
rect 97880 51100 98120 51120
rect 98380 51100 98620 51120
rect 98880 51100 99120 51120
rect 99380 51100 99620 51120
rect 99880 51100 100000 51120
rect 96000 51090 100000 51100
rect 96000 51020 96150 51090
rect 96350 51020 96650 51090
rect 96850 51020 97150 51090
rect 97350 51020 97650 51090
rect 97850 51020 98150 51090
rect 98350 51020 98650 51090
rect 98850 51020 99150 51090
rect 99350 51020 99650 51090
rect 99850 51020 100000 51090
rect 96000 50980 100000 51020
rect 96000 50910 96150 50980
rect 96350 50910 96650 50980
rect 96850 50910 97150 50980
rect 97350 50910 97650 50980
rect 97850 50910 98150 50980
rect 98350 50910 98650 50980
rect 98850 50910 99150 50980
rect 99350 50910 99650 50980
rect 99850 50910 100000 50980
rect 96000 50900 100000 50910
rect 96000 50880 96120 50900
rect 96380 50880 96620 50900
rect 96880 50880 97120 50900
rect 97380 50880 97620 50900
rect 97880 50880 98120 50900
rect 98380 50880 98620 50900
rect 98880 50880 99120 50900
rect 99380 50880 99620 50900
rect 99880 50880 100000 50900
rect 96000 50850 96100 50880
rect 96000 50650 96020 50850
rect 96090 50650 96100 50850
rect 96000 50620 96100 50650
rect 96400 50850 96600 50880
rect 96400 50650 96410 50850
rect 96480 50650 96520 50850
rect 96590 50650 96600 50850
rect 96400 50620 96600 50650
rect 96900 50850 97100 50880
rect 96900 50650 96910 50850
rect 96980 50650 97020 50850
rect 97090 50650 97100 50850
rect 96900 50620 97100 50650
rect 97400 50850 97600 50880
rect 97400 50650 97410 50850
rect 97480 50650 97520 50850
rect 97590 50650 97600 50850
rect 97400 50620 97600 50650
rect 97900 50850 98100 50880
rect 97900 50650 97910 50850
rect 97980 50650 98020 50850
rect 98090 50650 98100 50850
rect 97900 50620 98100 50650
rect 98400 50850 98600 50880
rect 98400 50650 98410 50850
rect 98480 50650 98520 50850
rect 98590 50650 98600 50850
rect 98400 50620 98600 50650
rect 98900 50850 99100 50880
rect 98900 50650 98910 50850
rect 98980 50650 99020 50850
rect 99090 50650 99100 50850
rect 98900 50620 99100 50650
rect 99400 50850 99600 50880
rect 99400 50650 99410 50850
rect 99480 50650 99520 50850
rect 99590 50650 99600 50850
rect 99400 50620 99600 50650
rect 99900 50850 100000 50880
rect 99900 50650 99910 50850
rect 99980 50650 100000 50850
rect 99900 50620 100000 50650
rect 96000 50600 96120 50620
rect 96380 50600 96620 50620
rect 96880 50600 97120 50620
rect 97380 50600 97620 50620
rect 97880 50600 98120 50620
rect 98380 50600 98620 50620
rect 98880 50600 99120 50620
rect 99380 50600 99620 50620
rect 99880 50600 100000 50620
rect 96000 50590 100000 50600
rect 96000 50520 96150 50590
rect 96350 50520 96650 50590
rect 96850 50520 97150 50590
rect 97350 50520 97650 50590
rect 97850 50520 98150 50590
rect 98350 50520 98650 50590
rect 98850 50520 99150 50590
rect 99350 50520 99650 50590
rect 99850 50520 100000 50590
rect 96000 50480 100000 50520
rect 96000 50410 96150 50480
rect 96350 50410 96650 50480
rect 96850 50410 97150 50480
rect 97350 50410 97650 50480
rect 97850 50410 98150 50480
rect 98350 50410 98650 50480
rect 98850 50410 99150 50480
rect 99350 50410 99650 50480
rect 99850 50410 100000 50480
rect 96000 50400 100000 50410
rect 96000 50380 96120 50400
rect 96380 50380 96620 50400
rect 96880 50380 97120 50400
rect 97380 50380 97620 50400
rect 97880 50380 98120 50400
rect 98380 50380 98620 50400
rect 98880 50380 99120 50400
rect 99380 50380 99620 50400
rect 99880 50380 100000 50400
rect 96000 50350 96100 50380
rect 96000 50150 96020 50350
rect 96090 50150 96100 50350
rect 96000 50120 96100 50150
rect 96400 50350 96600 50380
rect 96400 50150 96410 50350
rect 96480 50150 96520 50350
rect 96590 50150 96600 50350
rect 96400 50120 96600 50150
rect 96900 50350 97100 50380
rect 96900 50150 96910 50350
rect 96980 50150 97020 50350
rect 97090 50150 97100 50350
rect 96900 50120 97100 50150
rect 97400 50350 97600 50380
rect 97400 50150 97410 50350
rect 97480 50150 97520 50350
rect 97590 50150 97600 50350
rect 97400 50120 97600 50150
rect 97900 50350 98100 50380
rect 97900 50150 97910 50350
rect 97980 50150 98020 50350
rect 98090 50150 98100 50350
rect 97900 50120 98100 50150
rect 98400 50350 98600 50380
rect 98400 50150 98410 50350
rect 98480 50150 98520 50350
rect 98590 50150 98600 50350
rect 98400 50120 98600 50150
rect 98900 50350 99100 50380
rect 98900 50150 98910 50350
rect 98980 50150 99020 50350
rect 99090 50150 99100 50350
rect 98900 50120 99100 50150
rect 99400 50350 99600 50380
rect 99400 50150 99410 50350
rect 99480 50150 99520 50350
rect 99590 50150 99600 50350
rect 99400 50120 99600 50150
rect 99900 50350 100000 50380
rect 99900 50150 99910 50350
rect 99980 50150 100000 50350
rect 99900 50120 100000 50150
rect 96000 50100 96120 50120
rect 96380 50100 96620 50120
rect 96880 50100 97120 50120
rect 97380 50100 97620 50120
rect 97880 50100 98120 50120
rect 98380 50100 98620 50120
rect 98880 50100 99120 50120
rect 99380 50100 99620 50120
rect 99880 50100 100000 50120
rect 96000 50090 100000 50100
rect 96000 50020 96150 50090
rect 96350 50020 96650 50090
rect 96850 50020 97150 50090
rect 97350 50020 97650 50090
rect 97850 50020 98150 50090
rect 98350 50020 98650 50090
rect 98850 50020 99150 50090
rect 99350 50020 99650 50090
rect 99850 50020 100000 50090
rect 96000 50000 100000 50020
rect -16000 49910 -15850 49980
rect -15650 49910 -15350 49980
rect -15150 49910 -14850 49980
rect -14650 49910 -14350 49980
rect -14150 49910 -13850 49980
rect -13650 49910 -13350 49980
rect -13150 49910 -12850 49980
rect -12650 49910 -12350 49980
rect -12150 49910 -12000 49980
rect -16000 49900 -12000 49910
rect -16000 49880 -15880 49900
rect -15620 49880 -15380 49900
rect -15120 49880 -14880 49900
rect -14620 49880 -14380 49900
rect -14120 49880 -13880 49900
rect -13620 49880 -13380 49900
rect -13120 49880 -12880 49900
rect -12620 49880 -12380 49900
rect -12120 49880 -12000 49900
rect -16000 49850 -15900 49880
rect -16000 49650 -15980 49850
rect -15910 49650 -15900 49850
rect -16000 49620 -15900 49650
rect -15600 49850 -15400 49880
rect -15600 49650 -15590 49850
rect -15520 49650 -15480 49850
rect -15410 49650 -15400 49850
rect -15600 49620 -15400 49650
rect -15100 49850 -14900 49880
rect -15100 49650 -15090 49850
rect -15020 49650 -14980 49850
rect -14910 49650 -14900 49850
rect -15100 49620 -14900 49650
rect -14600 49850 -14400 49880
rect -14600 49650 -14590 49850
rect -14520 49650 -14480 49850
rect -14410 49650 -14400 49850
rect -14600 49620 -14400 49650
rect -14100 49850 -13900 49880
rect -14100 49650 -14090 49850
rect -14020 49650 -13980 49850
rect -13910 49650 -13900 49850
rect -14100 49620 -13900 49650
rect -13600 49850 -13400 49880
rect -13600 49650 -13590 49850
rect -13520 49650 -13480 49850
rect -13410 49650 -13400 49850
rect -13600 49620 -13400 49650
rect -13100 49850 -12900 49880
rect -13100 49650 -13090 49850
rect -13020 49650 -12980 49850
rect -12910 49650 -12900 49850
rect -13100 49620 -12900 49650
rect -12600 49850 -12400 49880
rect -12600 49650 -12590 49850
rect -12520 49650 -12480 49850
rect -12410 49650 -12400 49850
rect -12600 49620 -12400 49650
rect -12100 49850 -12000 49880
rect -12100 49650 -12090 49850
rect -12020 49650 -12000 49850
rect -12100 49620 -12000 49650
rect -16000 49600 -15880 49620
rect -15620 49600 -15380 49620
rect -15120 49600 -14880 49620
rect -14620 49600 -14380 49620
rect -14120 49600 -13880 49620
rect -13620 49600 -13380 49620
rect -13120 49600 -12880 49620
rect -12620 49600 -12380 49620
rect -12120 49600 -12000 49620
rect -16000 49590 -12000 49600
rect -16000 49520 -15850 49590
rect -15650 49520 -15350 49590
rect -15150 49520 -14850 49590
rect -14650 49520 -14350 49590
rect -14150 49520 -13850 49590
rect -13650 49520 -13350 49590
rect -13150 49520 -12850 49590
rect -12650 49520 -12350 49590
rect -12150 49520 -12000 49590
rect -16000 49480 -12000 49520
rect -16000 49410 -15850 49480
rect -15650 49410 -15350 49480
rect -15150 49410 -14850 49480
rect -14650 49410 -14350 49480
rect -14150 49410 -13850 49480
rect -13650 49410 -13350 49480
rect -13150 49410 -12850 49480
rect -12650 49410 -12350 49480
rect -12150 49410 -12000 49480
rect -16000 49400 -12000 49410
rect -16000 49380 -15880 49400
rect -15620 49380 -15380 49400
rect -15120 49380 -14880 49400
rect -14620 49380 -14380 49400
rect -14120 49380 -13880 49400
rect -13620 49380 -13380 49400
rect -13120 49380 -12880 49400
rect -12620 49380 -12380 49400
rect -12120 49380 -12000 49400
rect -16000 49350 -15900 49380
rect -16000 49150 -15980 49350
rect -15910 49150 -15900 49350
rect -16000 49120 -15900 49150
rect -15600 49350 -15400 49380
rect -15600 49150 -15590 49350
rect -15520 49150 -15480 49350
rect -15410 49150 -15400 49350
rect -15600 49120 -15400 49150
rect -15100 49350 -14900 49380
rect -15100 49150 -15090 49350
rect -15020 49150 -14980 49350
rect -14910 49150 -14900 49350
rect -15100 49120 -14900 49150
rect -14600 49350 -14400 49380
rect -14600 49150 -14590 49350
rect -14520 49150 -14480 49350
rect -14410 49150 -14400 49350
rect -14600 49120 -14400 49150
rect -14100 49350 -13900 49380
rect -14100 49150 -14090 49350
rect -14020 49150 -13980 49350
rect -13910 49150 -13900 49350
rect -14100 49120 -13900 49150
rect -13600 49350 -13400 49380
rect -13600 49150 -13590 49350
rect -13520 49150 -13480 49350
rect -13410 49150 -13400 49350
rect -13600 49120 -13400 49150
rect -13100 49350 -12900 49380
rect -13100 49150 -13090 49350
rect -13020 49150 -12980 49350
rect -12910 49150 -12900 49350
rect -13100 49120 -12900 49150
rect -12600 49350 -12400 49380
rect -12600 49150 -12590 49350
rect -12520 49150 -12480 49350
rect -12410 49150 -12400 49350
rect -12600 49120 -12400 49150
rect -12100 49350 -12000 49380
rect -12100 49150 -12090 49350
rect -12020 49150 -12000 49350
rect -12100 49120 -12000 49150
rect -16000 49100 -15880 49120
rect -15620 49100 -15380 49120
rect -15120 49100 -14880 49120
rect -14620 49100 -14380 49120
rect -14120 49100 -13880 49120
rect -13620 49100 -13380 49120
rect -13120 49100 -12880 49120
rect -12620 49100 -12380 49120
rect -12120 49100 -12000 49120
rect -16000 49090 -12000 49100
rect -16000 49020 -15850 49090
rect -15650 49020 -15350 49090
rect -15150 49020 -14850 49090
rect -14650 49020 -14350 49090
rect -14150 49020 -13850 49090
rect -13650 49020 -13350 49090
rect -13150 49020 -12850 49090
rect -12650 49020 -12350 49090
rect -12150 49020 -12000 49090
rect -16000 48980 -12000 49020
rect -16000 48910 -15850 48980
rect -15650 48910 -15350 48980
rect -15150 48910 -14850 48980
rect -14650 48910 -14350 48980
rect -14150 48910 -13850 48980
rect -13650 48910 -13350 48980
rect -13150 48910 -12850 48980
rect -12650 48910 -12350 48980
rect -12150 48910 -12000 48980
rect -16000 48900 -12000 48910
rect -16000 48880 -15880 48900
rect -15620 48880 -15380 48900
rect -15120 48880 -14880 48900
rect -14620 48880 -14380 48900
rect -14120 48880 -13880 48900
rect -13620 48880 -13380 48900
rect -13120 48880 -12880 48900
rect -12620 48880 -12380 48900
rect -12120 48880 -12000 48900
rect -16000 48850 -15900 48880
rect -16000 48650 -15980 48850
rect -15910 48650 -15900 48850
rect -16000 48620 -15900 48650
rect -15600 48850 -15400 48880
rect -15600 48650 -15590 48850
rect -15520 48650 -15480 48850
rect -15410 48650 -15400 48850
rect -15600 48620 -15400 48650
rect -15100 48850 -14900 48880
rect -15100 48650 -15090 48850
rect -15020 48650 -14980 48850
rect -14910 48650 -14900 48850
rect -15100 48620 -14900 48650
rect -14600 48850 -14400 48880
rect -14600 48650 -14590 48850
rect -14520 48650 -14480 48850
rect -14410 48650 -14400 48850
rect -14600 48620 -14400 48650
rect -14100 48850 -13900 48880
rect -14100 48650 -14090 48850
rect -14020 48650 -13980 48850
rect -13910 48650 -13900 48850
rect -14100 48620 -13900 48650
rect -13600 48850 -13400 48880
rect -13600 48650 -13590 48850
rect -13520 48650 -13480 48850
rect -13410 48650 -13400 48850
rect -13600 48620 -13400 48650
rect -13100 48850 -12900 48880
rect -13100 48650 -13090 48850
rect -13020 48650 -12980 48850
rect -12910 48650 -12900 48850
rect -13100 48620 -12900 48650
rect -12600 48850 -12400 48880
rect -12600 48650 -12590 48850
rect -12520 48650 -12480 48850
rect -12410 48650 -12400 48850
rect -12600 48620 -12400 48650
rect -12100 48850 -12000 48880
rect -12100 48650 -12090 48850
rect -12020 48650 -12000 48850
rect -12100 48620 -12000 48650
rect -16000 48600 -15880 48620
rect -15620 48600 -15380 48620
rect -15120 48600 -14880 48620
rect -14620 48600 -14380 48620
rect -14120 48600 -13880 48620
rect -13620 48600 -13380 48620
rect -13120 48600 -12880 48620
rect -12620 48600 -12380 48620
rect -12120 48600 -12000 48620
rect -16000 48590 -12000 48600
rect -16000 48520 -15850 48590
rect -15650 48520 -15350 48590
rect -15150 48520 -14850 48590
rect -14650 48520 -14350 48590
rect -14150 48520 -13850 48590
rect -13650 48520 -13350 48590
rect -13150 48520 -12850 48590
rect -12650 48520 -12350 48590
rect -12150 48520 -12000 48590
rect -16000 48480 -12000 48520
rect -16000 48410 -15850 48480
rect -15650 48410 -15350 48480
rect -15150 48410 -14850 48480
rect -14650 48410 -14350 48480
rect -14150 48410 -13850 48480
rect -13650 48410 -13350 48480
rect -13150 48410 -12850 48480
rect -12650 48410 -12350 48480
rect -12150 48410 -12000 48480
rect -16000 48400 -12000 48410
rect -16000 48380 -15880 48400
rect -15620 48380 -15380 48400
rect -15120 48380 -14880 48400
rect -14620 48380 -14380 48400
rect -14120 48380 -13880 48400
rect -13620 48380 -13380 48400
rect -13120 48380 -12880 48400
rect -12620 48380 -12380 48400
rect -12120 48380 -12000 48400
rect -16000 48350 -15900 48380
rect -16000 48150 -15980 48350
rect -15910 48150 -15900 48350
rect -16000 48120 -15900 48150
rect -15600 48350 -15400 48380
rect -15600 48150 -15590 48350
rect -15520 48150 -15480 48350
rect -15410 48150 -15400 48350
rect -15600 48120 -15400 48150
rect -15100 48350 -14900 48380
rect -15100 48150 -15090 48350
rect -15020 48150 -14980 48350
rect -14910 48150 -14900 48350
rect -15100 48120 -14900 48150
rect -14600 48350 -14400 48380
rect -14600 48150 -14590 48350
rect -14520 48150 -14480 48350
rect -14410 48150 -14400 48350
rect -14600 48120 -14400 48150
rect -14100 48350 -13900 48380
rect -14100 48150 -14090 48350
rect -14020 48150 -13980 48350
rect -13910 48150 -13900 48350
rect -14100 48120 -13900 48150
rect -13600 48350 -13400 48380
rect -13600 48150 -13590 48350
rect -13520 48150 -13480 48350
rect -13410 48150 -13400 48350
rect -13600 48120 -13400 48150
rect -13100 48350 -12900 48380
rect -13100 48150 -13090 48350
rect -13020 48150 -12980 48350
rect -12910 48150 -12900 48350
rect -13100 48120 -12900 48150
rect -12600 48350 -12400 48380
rect -12600 48150 -12590 48350
rect -12520 48150 -12480 48350
rect -12410 48150 -12400 48350
rect -12600 48120 -12400 48150
rect -12100 48350 -12000 48380
rect -12100 48150 -12090 48350
rect -12020 48150 -12000 48350
rect -12100 48120 -12000 48150
rect -16000 48100 -15880 48120
rect -15620 48100 -15380 48120
rect -15120 48100 -14880 48120
rect -14620 48100 -14380 48120
rect -14120 48100 -13880 48120
rect -13620 48100 -13380 48120
rect -13120 48100 -12880 48120
rect -12620 48100 -12380 48120
rect -12120 48100 -12000 48120
rect -16000 48090 -12000 48100
rect -16000 48020 -15850 48090
rect -15650 48020 -15350 48090
rect -15150 48020 -14850 48090
rect -14650 48020 -14350 48090
rect -14150 48020 -13850 48090
rect -13650 48020 -13350 48090
rect -13150 48020 -12850 48090
rect -12650 48020 -12350 48090
rect -12150 48020 -12000 48090
rect -16000 47980 -12000 48020
rect -16000 47910 -15850 47980
rect -15650 47910 -15350 47980
rect -15150 47910 -14850 47980
rect -14650 47910 -14350 47980
rect -14150 47910 -13850 47980
rect -13650 47910 -13350 47980
rect -13150 47910 -12850 47980
rect -12650 47910 -12350 47980
rect -12150 47910 -12000 47980
rect -16000 47900 -12000 47910
rect -16000 47880 -15880 47900
rect -15620 47880 -15380 47900
rect -15120 47880 -14880 47900
rect -14620 47880 -14380 47900
rect -14120 47880 -13880 47900
rect -13620 47880 -13380 47900
rect -13120 47880 -12880 47900
rect -12620 47880 -12380 47900
rect -12120 47880 -12000 47900
rect -16000 47850 -15900 47880
rect -16000 47650 -15980 47850
rect -15910 47650 -15900 47850
rect -16000 47620 -15900 47650
rect -15600 47850 -15400 47880
rect -15600 47650 -15590 47850
rect -15520 47650 -15480 47850
rect -15410 47650 -15400 47850
rect -15600 47620 -15400 47650
rect -15100 47850 -14900 47880
rect -15100 47650 -15090 47850
rect -15020 47650 -14980 47850
rect -14910 47650 -14900 47850
rect -15100 47620 -14900 47650
rect -14600 47850 -14400 47880
rect -14600 47650 -14590 47850
rect -14520 47650 -14480 47850
rect -14410 47650 -14400 47850
rect -14600 47620 -14400 47650
rect -14100 47850 -13900 47880
rect -14100 47650 -14090 47850
rect -14020 47650 -13980 47850
rect -13910 47650 -13900 47850
rect -14100 47620 -13900 47650
rect -13600 47850 -13400 47880
rect -13600 47650 -13590 47850
rect -13520 47650 -13480 47850
rect -13410 47650 -13400 47850
rect -13600 47620 -13400 47650
rect -13100 47850 -12900 47880
rect -13100 47650 -13090 47850
rect -13020 47650 -12980 47850
rect -12910 47650 -12900 47850
rect -13100 47620 -12900 47650
rect -12600 47850 -12400 47880
rect -12600 47650 -12590 47850
rect -12520 47650 -12480 47850
rect -12410 47650 -12400 47850
rect -12600 47620 -12400 47650
rect -12100 47850 -12000 47880
rect -12100 47650 -12090 47850
rect -12020 47650 -12000 47850
rect -12100 47620 -12000 47650
rect -16000 47600 -15880 47620
rect -15620 47600 -15380 47620
rect -15120 47600 -14880 47620
rect -14620 47600 -14380 47620
rect -14120 47600 -13880 47620
rect -13620 47600 -13380 47620
rect -13120 47600 -12880 47620
rect -12620 47600 -12380 47620
rect -12120 47600 -12000 47620
rect -16000 47590 -12000 47600
rect -16000 47520 -15850 47590
rect -15650 47520 -15350 47590
rect -15150 47520 -14850 47590
rect -14650 47520 -14350 47590
rect -14150 47520 -13850 47590
rect -13650 47520 -13350 47590
rect -13150 47520 -12850 47590
rect -12650 47520 -12350 47590
rect -12150 47520 -12000 47590
rect -16000 47480 -12000 47520
rect -16000 47410 -15850 47480
rect -15650 47410 -15350 47480
rect -15150 47410 -14850 47480
rect -14650 47410 -14350 47480
rect -14150 47410 -13850 47480
rect -13650 47410 -13350 47480
rect -13150 47410 -12850 47480
rect -12650 47410 -12350 47480
rect -12150 47410 -12000 47480
rect -16000 47400 -12000 47410
rect -16000 47380 -15880 47400
rect -15620 47380 -15380 47400
rect -15120 47380 -14880 47400
rect -14620 47380 -14380 47400
rect -14120 47380 -13880 47400
rect -13620 47380 -13380 47400
rect -13120 47380 -12880 47400
rect -12620 47380 -12380 47400
rect -12120 47380 -12000 47400
rect -16000 47350 -15900 47380
rect -16000 47150 -15980 47350
rect -15910 47150 -15900 47350
rect -16000 47120 -15900 47150
rect -15600 47350 -15400 47380
rect -15600 47150 -15590 47350
rect -15520 47150 -15480 47350
rect -15410 47150 -15400 47350
rect -15600 47120 -15400 47150
rect -15100 47350 -14900 47380
rect -15100 47150 -15090 47350
rect -15020 47150 -14980 47350
rect -14910 47150 -14900 47350
rect -15100 47120 -14900 47150
rect -14600 47350 -14400 47380
rect -14600 47150 -14590 47350
rect -14520 47150 -14480 47350
rect -14410 47150 -14400 47350
rect -14600 47120 -14400 47150
rect -14100 47350 -13900 47380
rect -14100 47150 -14090 47350
rect -14020 47150 -13980 47350
rect -13910 47150 -13900 47350
rect -14100 47120 -13900 47150
rect -13600 47350 -13400 47380
rect -13600 47150 -13590 47350
rect -13520 47150 -13480 47350
rect -13410 47150 -13400 47350
rect -13600 47120 -13400 47150
rect -13100 47350 -12900 47380
rect -13100 47150 -13090 47350
rect -13020 47150 -12980 47350
rect -12910 47150 -12900 47350
rect -13100 47120 -12900 47150
rect -12600 47350 -12400 47380
rect -12600 47150 -12590 47350
rect -12520 47150 -12480 47350
rect -12410 47150 -12400 47350
rect -12600 47120 -12400 47150
rect -12100 47350 -12000 47380
rect -12100 47150 -12090 47350
rect -12020 47150 -12000 47350
rect -12100 47120 -12000 47150
rect -16000 47100 -15880 47120
rect -15620 47100 -15380 47120
rect -15120 47100 -14880 47120
rect -14620 47100 -14380 47120
rect -14120 47100 -13880 47120
rect -13620 47100 -13380 47120
rect -13120 47100 -12880 47120
rect -12620 47100 -12380 47120
rect -12120 47100 -12000 47120
rect -16000 47090 -12000 47100
rect -16000 47020 -15850 47090
rect -15650 47020 -15350 47090
rect -15150 47020 -14850 47090
rect -14650 47020 -14350 47090
rect -14150 47020 -13850 47090
rect -13650 47020 -13350 47090
rect -13150 47020 -12850 47090
rect -12650 47020 -12350 47090
rect -12150 47020 -12000 47090
rect -16000 46980 -12000 47020
rect -16000 46910 -15850 46980
rect -15650 46910 -15350 46980
rect -15150 46910 -14850 46980
rect -14650 46910 -14350 46980
rect -14150 46910 -13850 46980
rect -13650 46910 -13350 46980
rect -13150 46910 -12850 46980
rect -12650 46910 -12350 46980
rect -12150 46910 -12000 46980
rect -16000 46900 -12000 46910
rect -16000 46880 -15880 46900
rect -15620 46880 -15380 46900
rect -15120 46880 -14880 46900
rect -14620 46880 -14380 46900
rect -14120 46880 -13880 46900
rect -13620 46880 -13380 46900
rect -13120 46880 -12880 46900
rect -12620 46880 -12380 46900
rect -12120 46880 -12000 46900
rect -16000 46850 -15900 46880
rect -16000 46650 -15980 46850
rect -15910 46650 -15900 46850
rect -16000 46620 -15900 46650
rect -15600 46850 -15400 46880
rect -15600 46650 -15590 46850
rect -15520 46650 -15480 46850
rect -15410 46650 -15400 46850
rect -15600 46620 -15400 46650
rect -15100 46850 -14900 46880
rect -15100 46650 -15090 46850
rect -15020 46650 -14980 46850
rect -14910 46650 -14900 46850
rect -15100 46620 -14900 46650
rect -14600 46850 -14400 46880
rect -14600 46650 -14590 46850
rect -14520 46650 -14480 46850
rect -14410 46650 -14400 46850
rect -14600 46620 -14400 46650
rect -14100 46850 -13900 46880
rect -14100 46650 -14090 46850
rect -14020 46650 -13980 46850
rect -13910 46650 -13900 46850
rect -14100 46620 -13900 46650
rect -13600 46850 -13400 46880
rect -13600 46650 -13590 46850
rect -13520 46650 -13480 46850
rect -13410 46650 -13400 46850
rect -13600 46620 -13400 46650
rect -13100 46850 -12900 46880
rect -13100 46650 -13090 46850
rect -13020 46650 -12980 46850
rect -12910 46650 -12900 46850
rect -13100 46620 -12900 46650
rect -12600 46850 -12400 46880
rect -12600 46650 -12590 46850
rect -12520 46650 -12480 46850
rect -12410 46650 -12400 46850
rect -12600 46620 -12400 46650
rect -12100 46850 -12000 46880
rect -12100 46650 -12090 46850
rect -12020 46650 -12000 46850
rect -12100 46620 -12000 46650
rect -16000 46600 -15880 46620
rect -15620 46600 -15380 46620
rect -15120 46600 -14880 46620
rect -14620 46600 -14380 46620
rect -14120 46600 -13880 46620
rect -13620 46600 -13380 46620
rect -13120 46600 -12880 46620
rect -12620 46600 -12380 46620
rect -12120 46600 -12000 46620
rect -16000 46590 -12000 46600
rect -16000 46520 -15850 46590
rect -15650 46520 -15350 46590
rect -15150 46520 -14850 46590
rect -14650 46520 -14350 46590
rect -14150 46520 -13850 46590
rect -13650 46520 -13350 46590
rect -13150 46520 -12850 46590
rect -12650 46520 -12350 46590
rect -12150 46520 -12000 46590
rect -16000 46480 -12000 46520
rect -16000 46410 -15850 46480
rect -15650 46410 -15350 46480
rect -15150 46410 -14850 46480
rect -14650 46410 -14350 46480
rect -14150 46410 -13850 46480
rect -13650 46410 -13350 46480
rect -13150 46410 -12850 46480
rect -12650 46410 -12350 46480
rect -12150 46410 -12000 46480
rect -16000 46400 -12000 46410
rect -16000 46380 -15880 46400
rect -15620 46380 -15380 46400
rect -15120 46380 -14880 46400
rect -14620 46380 -14380 46400
rect -14120 46380 -13880 46400
rect -13620 46380 -13380 46400
rect -13120 46380 -12880 46400
rect -12620 46380 -12380 46400
rect -12120 46380 -12000 46400
rect -16000 46350 -15900 46380
rect -16000 46150 -15980 46350
rect -15910 46150 -15900 46350
rect -16000 46120 -15900 46150
rect -15600 46350 -15400 46380
rect -15600 46150 -15590 46350
rect -15520 46150 -15480 46350
rect -15410 46150 -15400 46350
rect -15600 46120 -15400 46150
rect -15100 46350 -14900 46380
rect -15100 46150 -15090 46350
rect -15020 46150 -14980 46350
rect -14910 46150 -14900 46350
rect -15100 46120 -14900 46150
rect -14600 46350 -14400 46380
rect -14600 46150 -14590 46350
rect -14520 46150 -14480 46350
rect -14410 46150 -14400 46350
rect -14600 46120 -14400 46150
rect -14100 46350 -13900 46380
rect -14100 46150 -14090 46350
rect -14020 46150 -13980 46350
rect -13910 46150 -13900 46350
rect -14100 46120 -13900 46150
rect -13600 46350 -13400 46380
rect -13600 46150 -13590 46350
rect -13520 46150 -13480 46350
rect -13410 46150 -13400 46350
rect -13600 46120 -13400 46150
rect -13100 46350 -12900 46380
rect -13100 46150 -13090 46350
rect -13020 46150 -12980 46350
rect -12910 46150 -12900 46350
rect -13100 46120 -12900 46150
rect -12600 46350 -12400 46380
rect -12600 46150 -12590 46350
rect -12520 46150 -12480 46350
rect -12410 46150 -12400 46350
rect -12600 46120 -12400 46150
rect -12100 46350 -12000 46380
rect -12100 46150 -12090 46350
rect -12020 46150 -12000 46350
rect -12100 46120 -12000 46150
rect -16000 46100 -15880 46120
rect -15620 46100 -15380 46120
rect -15120 46100 -14880 46120
rect -14620 46100 -14380 46120
rect -14120 46100 -13880 46120
rect -13620 46100 -13380 46120
rect -13120 46100 -12880 46120
rect -12620 46100 -12380 46120
rect -12120 46100 -12000 46120
rect -16000 46090 -12000 46100
rect -16000 46020 -15850 46090
rect -15650 46020 -15350 46090
rect -15150 46020 -14850 46090
rect -14650 46020 -14350 46090
rect -14150 46020 -13850 46090
rect -13650 46020 -13350 46090
rect -13150 46020 -12850 46090
rect -12650 46020 -12350 46090
rect -12150 46020 -12000 46090
rect -16000 45980 -12000 46020
rect -16000 45910 -15850 45980
rect -15650 45910 -15350 45980
rect -15150 45910 -14850 45980
rect -14650 45910 -14350 45980
rect -14150 45910 -13850 45980
rect -13650 45910 -13350 45980
rect -13150 45910 -12850 45980
rect -12650 45910 -12350 45980
rect -12150 45910 -12000 45980
rect -16000 45900 -12000 45910
rect -16000 45880 -15880 45900
rect -15620 45880 -15380 45900
rect -15120 45880 -14880 45900
rect -14620 45880 -14380 45900
rect -14120 45880 -13880 45900
rect -13620 45880 -13380 45900
rect -13120 45880 -12880 45900
rect -12620 45880 -12380 45900
rect -12120 45880 -12000 45900
rect -16000 45850 -15900 45880
rect -16000 45650 -15980 45850
rect -15910 45650 -15900 45850
rect -16000 45620 -15900 45650
rect -15600 45850 -15400 45880
rect -15600 45650 -15590 45850
rect -15520 45650 -15480 45850
rect -15410 45650 -15400 45850
rect -15600 45620 -15400 45650
rect -15100 45850 -14900 45880
rect -15100 45650 -15090 45850
rect -15020 45650 -14980 45850
rect -14910 45650 -14900 45850
rect -15100 45620 -14900 45650
rect -14600 45850 -14400 45880
rect -14600 45650 -14590 45850
rect -14520 45650 -14480 45850
rect -14410 45650 -14400 45850
rect -14600 45620 -14400 45650
rect -14100 45850 -13900 45880
rect -14100 45650 -14090 45850
rect -14020 45650 -13980 45850
rect -13910 45650 -13900 45850
rect -14100 45620 -13900 45650
rect -13600 45850 -13400 45880
rect -13600 45650 -13590 45850
rect -13520 45650 -13480 45850
rect -13410 45650 -13400 45850
rect -13600 45620 -13400 45650
rect -13100 45850 -12900 45880
rect -13100 45650 -13090 45850
rect -13020 45650 -12980 45850
rect -12910 45650 -12900 45850
rect -13100 45620 -12900 45650
rect -12600 45850 -12400 45880
rect -12600 45650 -12590 45850
rect -12520 45650 -12480 45850
rect -12410 45650 -12400 45850
rect -12600 45620 -12400 45650
rect -12100 45850 -12000 45880
rect -12100 45650 -12090 45850
rect -12020 45650 -12000 45850
rect -12100 45620 -12000 45650
rect -16000 45600 -15880 45620
rect -15620 45600 -15380 45620
rect -15120 45600 -14880 45620
rect -14620 45600 -14380 45620
rect -14120 45600 -13880 45620
rect -13620 45600 -13380 45620
rect -13120 45600 -12880 45620
rect -12620 45600 -12380 45620
rect -12120 45600 -12000 45620
rect -16000 45590 -12000 45600
rect -16000 45520 -15850 45590
rect -15650 45520 -15350 45590
rect -15150 45520 -14850 45590
rect -14650 45520 -14350 45590
rect -14150 45520 -13850 45590
rect -13650 45520 -13350 45590
rect -13150 45520 -12850 45590
rect -12650 45520 -12350 45590
rect -12150 45520 -12000 45590
rect -16000 45480 -12000 45520
rect -16000 45410 -15850 45480
rect -15650 45410 -15350 45480
rect -15150 45410 -14850 45480
rect -14650 45410 -14350 45480
rect -14150 45410 -13850 45480
rect -13650 45410 -13350 45480
rect -13150 45410 -12850 45480
rect -12650 45410 -12350 45480
rect -12150 45410 -12000 45480
rect -16000 45400 -12000 45410
rect -16000 45380 -15880 45400
rect -15620 45380 -15380 45400
rect -15120 45380 -14880 45400
rect -14620 45380 -14380 45400
rect -14120 45380 -13880 45400
rect -13620 45380 -13380 45400
rect -13120 45380 -12880 45400
rect -12620 45380 -12380 45400
rect -12120 45380 -12000 45400
rect -16000 45350 -15900 45380
rect -16000 45150 -15980 45350
rect -15910 45150 -15900 45350
rect -16000 45120 -15900 45150
rect -15600 45350 -15400 45380
rect -15600 45150 -15590 45350
rect -15520 45150 -15480 45350
rect -15410 45150 -15400 45350
rect -15600 45120 -15400 45150
rect -15100 45350 -14900 45380
rect -15100 45150 -15090 45350
rect -15020 45150 -14980 45350
rect -14910 45150 -14900 45350
rect -15100 45120 -14900 45150
rect -14600 45350 -14400 45380
rect -14600 45150 -14590 45350
rect -14520 45150 -14480 45350
rect -14410 45150 -14400 45350
rect -14600 45120 -14400 45150
rect -14100 45350 -13900 45380
rect -14100 45150 -14090 45350
rect -14020 45150 -13980 45350
rect -13910 45150 -13900 45350
rect -14100 45120 -13900 45150
rect -13600 45350 -13400 45380
rect -13600 45150 -13590 45350
rect -13520 45150 -13480 45350
rect -13410 45150 -13400 45350
rect -13600 45120 -13400 45150
rect -13100 45350 -12900 45380
rect -13100 45150 -13090 45350
rect -13020 45150 -12980 45350
rect -12910 45150 -12900 45350
rect -13100 45120 -12900 45150
rect -12600 45350 -12400 45380
rect -12600 45150 -12590 45350
rect -12520 45150 -12480 45350
rect -12410 45150 -12400 45350
rect -12600 45120 -12400 45150
rect -12100 45350 -12000 45380
rect -12100 45150 -12090 45350
rect -12020 45150 -12000 45350
rect -12100 45120 -12000 45150
rect -16000 45100 -15880 45120
rect -15620 45100 -15380 45120
rect -15120 45100 -14880 45120
rect -14620 45100 -14380 45120
rect -14120 45100 -13880 45120
rect -13620 45100 -13380 45120
rect -13120 45100 -12880 45120
rect -12620 45100 -12380 45120
rect -12120 45100 -12000 45120
rect -16000 45090 -12000 45100
rect -16000 45020 -15850 45090
rect -15650 45020 -15350 45090
rect -15150 45020 -14850 45090
rect -14650 45020 -14350 45090
rect -14150 45020 -13850 45090
rect -13650 45020 -13350 45090
rect -13150 45020 -12850 45090
rect -12650 45020 -12350 45090
rect -12150 45020 -12000 45090
rect -16000 44980 -12000 45020
rect -16000 44910 -15850 44980
rect -15650 44910 -15350 44980
rect -15150 44910 -14850 44980
rect -14650 44910 -14350 44980
rect -14150 44910 -13850 44980
rect -13650 44910 -13350 44980
rect -13150 44910 -12850 44980
rect -12650 44910 -12350 44980
rect -12150 44910 -12000 44980
rect -16000 44900 -12000 44910
rect -16000 44880 -15880 44900
rect -15620 44880 -15380 44900
rect -15120 44880 -14880 44900
rect -14620 44880 -14380 44900
rect -14120 44880 -13880 44900
rect -13620 44880 -13380 44900
rect -13120 44880 -12880 44900
rect -12620 44880 -12380 44900
rect -12120 44880 -12000 44900
rect -16000 44850 -15900 44880
rect -16000 44650 -15980 44850
rect -15910 44650 -15900 44850
rect -16000 44620 -15900 44650
rect -15600 44850 -15400 44880
rect -15600 44650 -15590 44850
rect -15520 44650 -15480 44850
rect -15410 44650 -15400 44850
rect -15600 44620 -15400 44650
rect -15100 44850 -14900 44880
rect -15100 44650 -15090 44850
rect -15020 44650 -14980 44850
rect -14910 44650 -14900 44850
rect -15100 44620 -14900 44650
rect -14600 44850 -14400 44880
rect -14600 44650 -14590 44850
rect -14520 44650 -14480 44850
rect -14410 44650 -14400 44850
rect -14600 44620 -14400 44650
rect -14100 44850 -13900 44880
rect -14100 44650 -14090 44850
rect -14020 44650 -13980 44850
rect -13910 44650 -13900 44850
rect -14100 44620 -13900 44650
rect -13600 44850 -13400 44880
rect -13600 44650 -13590 44850
rect -13520 44650 -13480 44850
rect -13410 44650 -13400 44850
rect -13600 44620 -13400 44650
rect -13100 44850 -12900 44880
rect -13100 44650 -13090 44850
rect -13020 44650 -12980 44850
rect -12910 44650 -12900 44850
rect -13100 44620 -12900 44650
rect -12600 44850 -12400 44880
rect -12600 44650 -12590 44850
rect -12520 44650 -12480 44850
rect -12410 44650 -12400 44850
rect -12600 44620 -12400 44650
rect -12100 44850 -12000 44880
rect -12100 44650 -12090 44850
rect -12020 44650 -12000 44850
rect -12100 44620 -12000 44650
rect -16000 44600 -15880 44620
rect -15620 44600 -15380 44620
rect -15120 44600 -14880 44620
rect -14620 44600 -14380 44620
rect -14120 44600 -13880 44620
rect -13620 44600 -13380 44620
rect -13120 44600 -12880 44620
rect -12620 44600 -12380 44620
rect -12120 44600 -12000 44620
rect -16000 44590 -12000 44600
rect -16000 44520 -15850 44590
rect -15650 44520 -15350 44590
rect -15150 44520 -14850 44590
rect -14650 44520 -14350 44590
rect -14150 44520 -13850 44590
rect -13650 44520 -13350 44590
rect -13150 44520 -12850 44590
rect -12650 44520 -12350 44590
rect -12150 44520 -12000 44590
rect -16000 44480 -12000 44520
rect -16000 44410 -15850 44480
rect -15650 44410 -15350 44480
rect -15150 44410 -14850 44480
rect -14650 44410 -14350 44480
rect -14150 44410 -13850 44480
rect -13650 44410 -13350 44480
rect -13150 44410 -12850 44480
rect -12650 44410 -12350 44480
rect -12150 44410 -12000 44480
rect -16000 44400 -12000 44410
rect -16000 44380 -15880 44400
rect -15620 44380 -15380 44400
rect -15120 44380 -14880 44400
rect -14620 44380 -14380 44400
rect -14120 44380 -13880 44400
rect -13620 44380 -13380 44400
rect -13120 44380 -12880 44400
rect -12620 44380 -12380 44400
rect -12120 44380 -12000 44400
rect -16000 44350 -15900 44380
rect -16000 44150 -15980 44350
rect -15910 44150 -15900 44350
rect -16000 44120 -15900 44150
rect -15600 44350 -15400 44380
rect -15600 44150 -15590 44350
rect -15520 44150 -15480 44350
rect -15410 44150 -15400 44350
rect -15600 44120 -15400 44150
rect -15100 44350 -14900 44380
rect -15100 44150 -15090 44350
rect -15020 44150 -14980 44350
rect -14910 44150 -14900 44350
rect -15100 44120 -14900 44150
rect -14600 44350 -14400 44380
rect -14600 44150 -14590 44350
rect -14520 44150 -14480 44350
rect -14410 44150 -14400 44350
rect -14600 44120 -14400 44150
rect -14100 44350 -13900 44380
rect -14100 44150 -14090 44350
rect -14020 44150 -13980 44350
rect -13910 44150 -13900 44350
rect -14100 44120 -13900 44150
rect -13600 44350 -13400 44380
rect -13600 44150 -13590 44350
rect -13520 44150 -13480 44350
rect -13410 44150 -13400 44350
rect -13600 44120 -13400 44150
rect -13100 44350 -12900 44380
rect -13100 44150 -13090 44350
rect -13020 44150 -12980 44350
rect -12910 44150 -12900 44350
rect -13100 44120 -12900 44150
rect -12600 44350 -12400 44380
rect -12600 44150 -12590 44350
rect -12520 44150 -12480 44350
rect -12410 44150 -12400 44350
rect -12600 44120 -12400 44150
rect -12100 44350 -12000 44380
rect -12100 44150 -12090 44350
rect -12020 44150 -12000 44350
rect -12100 44120 -12000 44150
rect -16000 44100 -15880 44120
rect -15620 44100 -15380 44120
rect -15120 44100 -14880 44120
rect -14620 44100 -14380 44120
rect -14120 44100 -13880 44120
rect -13620 44100 -13380 44120
rect -13120 44100 -12880 44120
rect -12620 44100 -12380 44120
rect -12120 44100 -12000 44120
rect -16000 44090 -12000 44100
rect -16000 44020 -15850 44090
rect -15650 44020 -15350 44090
rect -15150 44020 -14850 44090
rect -14650 44020 -14350 44090
rect -14150 44020 -13850 44090
rect -13650 44020 -13350 44090
rect -13150 44020 -12850 44090
rect -12650 44020 -12350 44090
rect -12150 44020 -12000 44090
rect -16000 43980 -12000 44020
rect -16000 43910 -15850 43980
rect -15650 43910 -15350 43980
rect -15150 43910 -14850 43980
rect -14650 43910 -14350 43980
rect -14150 43910 -13850 43980
rect -13650 43910 -13350 43980
rect -13150 43910 -12850 43980
rect -12650 43910 -12350 43980
rect -12150 43910 -12000 43980
rect -16000 43900 -12000 43910
rect -16000 43880 -15880 43900
rect -15620 43880 -15380 43900
rect -15120 43880 -14880 43900
rect -14620 43880 -14380 43900
rect -14120 43880 -13880 43900
rect -13620 43880 -13380 43900
rect -13120 43880 -12880 43900
rect -12620 43880 -12380 43900
rect -12120 43880 -12000 43900
rect -16000 43850 -15900 43880
rect -16000 43650 -15980 43850
rect -15910 43650 -15900 43850
rect -16000 43620 -15900 43650
rect -15600 43850 -15400 43880
rect -15600 43650 -15590 43850
rect -15520 43650 -15480 43850
rect -15410 43650 -15400 43850
rect -15600 43620 -15400 43650
rect -15100 43850 -14900 43880
rect -15100 43650 -15090 43850
rect -15020 43650 -14980 43850
rect -14910 43650 -14900 43850
rect -15100 43620 -14900 43650
rect -14600 43850 -14400 43880
rect -14600 43650 -14590 43850
rect -14520 43650 -14480 43850
rect -14410 43650 -14400 43850
rect -14600 43620 -14400 43650
rect -14100 43850 -13900 43880
rect -14100 43650 -14090 43850
rect -14020 43650 -13980 43850
rect -13910 43650 -13900 43850
rect -14100 43620 -13900 43650
rect -13600 43850 -13400 43880
rect -13600 43650 -13590 43850
rect -13520 43650 -13480 43850
rect -13410 43650 -13400 43850
rect -13600 43620 -13400 43650
rect -13100 43850 -12900 43880
rect -13100 43650 -13090 43850
rect -13020 43650 -12980 43850
rect -12910 43650 -12900 43850
rect -13100 43620 -12900 43650
rect -12600 43850 -12400 43880
rect -12600 43650 -12590 43850
rect -12520 43650 -12480 43850
rect -12410 43650 -12400 43850
rect -12600 43620 -12400 43650
rect -12100 43850 -12000 43880
rect -12100 43650 -12090 43850
rect -12020 43650 -12000 43850
rect -12100 43620 -12000 43650
rect -16000 43600 -15880 43620
rect -15620 43600 -15380 43620
rect -15120 43600 -14880 43620
rect -14620 43600 -14380 43620
rect -14120 43600 -13880 43620
rect -13620 43600 -13380 43620
rect -13120 43600 -12880 43620
rect -12620 43600 -12380 43620
rect -12120 43600 -12000 43620
rect -16000 43590 -12000 43600
rect -16000 43520 -15850 43590
rect -15650 43520 -15350 43590
rect -15150 43520 -14850 43590
rect -14650 43520 -14350 43590
rect -14150 43520 -13850 43590
rect -13650 43520 -13350 43590
rect -13150 43520 -12850 43590
rect -12650 43520 -12350 43590
rect -12150 43520 -12000 43590
rect -16000 43480 -12000 43520
rect -16000 43410 -15850 43480
rect -15650 43410 -15350 43480
rect -15150 43410 -14850 43480
rect -14650 43410 -14350 43480
rect -14150 43410 -13850 43480
rect -13650 43410 -13350 43480
rect -13150 43410 -12850 43480
rect -12650 43410 -12350 43480
rect -12150 43410 -12000 43480
rect -16000 43400 -12000 43410
rect -16000 43380 -15880 43400
rect -15620 43380 -15380 43400
rect -15120 43380 -14880 43400
rect -14620 43380 -14380 43400
rect -14120 43380 -13880 43400
rect -13620 43380 -13380 43400
rect -13120 43380 -12880 43400
rect -12620 43380 -12380 43400
rect -12120 43380 -12000 43400
rect -16000 43350 -15900 43380
rect -16000 43150 -15980 43350
rect -15910 43150 -15900 43350
rect -16000 43120 -15900 43150
rect -15600 43350 -15400 43380
rect -15600 43150 -15590 43350
rect -15520 43150 -15480 43350
rect -15410 43150 -15400 43350
rect -15600 43120 -15400 43150
rect -15100 43350 -14900 43380
rect -15100 43150 -15090 43350
rect -15020 43150 -14980 43350
rect -14910 43150 -14900 43350
rect -15100 43120 -14900 43150
rect -14600 43350 -14400 43380
rect -14600 43150 -14590 43350
rect -14520 43150 -14480 43350
rect -14410 43150 -14400 43350
rect -14600 43120 -14400 43150
rect -14100 43350 -13900 43380
rect -14100 43150 -14090 43350
rect -14020 43150 -13980 43350
rect -13910 43150 -13900 43350
rect -14100 43120 -13900 43150
rect -13600 43350 -13400 43380
rect -13600 43150 -13590 43350
rect -13520 43150 -13480 43350
rect -13410 43150 -13400 43350
rect -13600 43120 -13400 43150
rect -13100 43350 -12900 43380
rect -13100 43150 -13090 43350
rect -13020 43150 -12980 43350
rect -12910 43150 -12900 43350
rect -13100 43120 -12900 43150
rect -12600 43350 -12400 43380
rect -12600 43150 -12590 43350
rect -12520 43150 -12480 43350
rect -12410 43150 -12400 43350
rect -12600 43120 -12400 43150
rect -12100 43350 -12000 43380
rect -12100 43150 -12090 43350
rect -12020 43150 -12000 43350
rect -12100 43120 -12000 43150
rect -16000 43100 -15880 43120
rect -15620 43100 -15380 43120
rect -15120 43100 -14880 43120
rect -14620 43100 -14380 43120
rect -14120 43100 -13880 43120
rect -13620 43100 -13380 43120
rect -13120 43100 -12880 43120
rect -12620 43100 -12380 43120
rect -12120 43100 -12000 43120
rect -16000 43090 -12000 43100
rect -16000 43020 -15850 43090
rect -15650 43020 -15350 43090
rect -15150 43020 -14850 43090
rect -14650 43020 -14350 43090
rect -14150 43020 -13850 43090
rect -13650 43020 -13350 43090
rect -13150 43020 -12850 43090
rect -12650 43020 -12350 43090
rect -12150 43020 -12000 43090
rect -16000 42980 -12000 43020
rect -16000 42910 -15850 42980
rect -15650 42910 -15350 42980
rect -15150 42910 -14850 42980
rect -14650 42910 -14350 42980
rect -14150 42910 -13850 42980
rect -13650 42910 -13350 42980
rect -13150 42910 -12850 42980
rect -12650 42910 -12350 42980
rect -12150 42910 -12000 42980
rect -16000 42900 -12000 42910
rect -16000 42880 -15880 42900
rect -15620 42880 -15380 42900
rect -15120 42880 -14880 42900
rect -14620 42880 -14380 42900
rect -14120 42880 -13880 42900
rect -13620 42880 -13380 42900
rect -13120 42880 -12880 42900
rect -12620 42880 -12380 42900
rect -12120 42880 -12000 42900
rect -16000 42850 -15900 42880
rect -16000 42650 -15980 42850
rect -15910 42650 -15900 42850
rect -16000 42620 -15900 42650
rect -15600 42850 -15400 42880
rect -15600 42650 -15590 42850
rect -15520 42650 -15480 42850
rect -15410 42650 -15400 42850
rect -15600 42620 -15400 42650
rect -15100 42850 -14900 42880
rect -15100 42650 -15090 42850
rect -15020 42650 -14980 42850
rect -14910 42650 -14900 42850
rect -15100 42620 -14900 42650
rect -14600 42850 -14400 42880
rect -14600 42650 -14590 42850
rect -14520 42650 -14480 42850
rect -14410 42650 -14400 42850
rect -14600 42620 -14400 42650
rect -14100 42850 -13900 42880
rect -14100 42650 -14090 42850
rect -14020 42650 -13980 42850
rect -13910 42650 -13900 42850
rect -14100 42620 -13900 42650
rect -13600 42850 -13400 42880
rect -13600 42650 -13590 42850
rect -13520 42650 -13480 42850
rect -13410 42650 -13400 42850
rect -13600 42620 -13400 42650
rect -13100 42850 -12900 42880
rect -13100 42650 -13090 42850
rect -13020 42650 -12980 42850
rect -12910 42650 -12900 42850
rect -13100 42620 -12900 42650
rect -12600 42850 -12400 42880
rect -12600 42650 -12590 42850
rect -12520 42650 -12480 42850
rect -12410 42650 -12400 42850
rect -12600 42620 -12400 42650
rect -12100 42850 -12000 42880
rect -12100 42650 -12090 42850
rect -12020 42650 -12000 42850
rect -12100 42620 -12000 42650
rect -16000 42600 -15880 42620
rect -15620 42600 -15380 42620
rect -15120 42600 -14880 42620
rect -14620 42600 -14380 42620
rect -14120 42600 -13880 42620
rect -13620 42600 -13380 42620
rect -13120 42600 -12880 42620
rect -12620 42600 -12380 42620
rect -12120 42600 -12000 42620
rect -16000 42590 -12000 42600
rect -16000 42520 -15850 42590
rect -15650 42520 -15350 42590
rect -15150 42520 -14850 42590
rect -14650 42520 -14350 42590
rect -14150 42520 -13850 42590
rect -13650 42520 -13350 42590
rect -13150 42520 -12850 42590
rect -12650 42520 -12350 42590
rect -12150 42520 -12000 42590
rect -16000 42480 -12000 42520
rect -16000 42410 -15850 42480
rect -15650 42410 -15350 42480
rect -15150 42410 -14850 42480
rect -14650 42410 -14350 42480
rect -14150 42410 -13850 42480
rect -13650 42410 -13350 42480
rect -13150 42410 -12850 42480
rect -12650 42410 -12350 42480
rect -12150 42410 -12000 42480
rect -16000 42400 -12000 42410
rect -16000 42380 -15880 42400
rect -15620 42380 -15380 42400
rect -15120 42380 -14880 42400
rect -14620 42380 -14380 42400
rect -14120 42380 -13880 42400
rect -13620 42380 -13380 42400
rect -13120 42380 -12880 42400
rect -12620 42380 -12380 42400
rect -12120 42380 -12000 42400
rect -16000 42350 -15900 42380
rect -16000 42150 -15980 42350
rect -15910 42150 -15900 42350
rect -16000 42120 -15900 42150
rect -15600 42350 -15400 42380
rect -15600 42150 -15590 42350
rect -15520 42150 -15480 42350
rect -15410 42150 -15400 42350
rect -15600 42120 -15400 42150
rect -15100 42350 -14900 42380
rect -15100 42150 -15090 42350
rect -15020 42150 -14980 42350
rect -14910 42150 -14900 42350
rect -15100 42120 -14900 42150
rect -14600 42350 -14400 42380
rect -14600 42150 -14590 42350
rect -14520 42150 -14480 42350
rect -14410 42150 -14400 42350
rect -14600 42120 -14400 42150
rect -14100 42350 -13900 42380
rect -14100 42150 -14090 42350
rect -14020 42150 -13980 42350
rect -13910 42150 -13900 42350
rect -14100 42120 -13900 42150
rect -13600 42350 -13400 42380
rect -13600 42150 -13590 42350
rect -13520 42150 -13480 42350
rect -13410 42150 -13400 42350
rect -13600 42120 -13400 42150
rect -13100 42350 -12900 42380
rect -13100 42150 -13090 42350
rect -13020 42150 -12980 42350
rect -12910 42150 -12900 42350
rect -13100 42120 -12900 42150
rect -12600 42350 -12400 42380
rect -12600 42150 -12590 42350
rect -12520 42150 -12480 42350
rect -12410 42150 -12400 42350
rect -12600 42120 -12400 42150
rect -12100 42350 -12000 42380
rect -12100 42150 -12090 42350
rect -12020 42150 -12000 42350
rect -12100 42120 -12000 42150
rect -16000 42100 -15880 42120
rect -15620 42100 -15380 42120
rect -15120 42100 -14880 42120
rect -14620 42100 -14380 42120
rect -14120 42100 -13880 42120
rect -13620 42100 -13380 42120
rect -13120 42100 -12880 42120
rect -12620 42100 -12380 42120
rect -12120 42100 -12000 42120
rect -16000 42090 -12000 42100
rect -16000 42020 -15850 42090
rect -15650 42020 -15350 42090
rect -15150 42020 -14850 42090
rect -14650 42020 -14350 42090
rect -14150 42020 -13850 42090
rect -13650 42020 -13350 42090
rect -13150 42020 -12850 42090
rect -12650 42020 -12350 42090
rect -12150 42020 -12000 42090
rect -16000 42000 -12000 42020
rect -16000 41980 4000 42000
rect -16000 41910 -15850 41980
rect -15650 41910 -15350 41980
rect -15150 41910 -14850 41980
rect -14650 41910 -14350 41980
rect -14150 41910 -13850 41980
rect -13650 41910 -13350 41980
rect -13150 41910 -12850 41980
rect -12650 41910 -12350 41980
rect -12150 41910 -11850 41980
rect -11650 41910 -11350 41980
rect -11150 41910 -10850 41980
rect -10650 41910 -10350 41980
rect -10150 41910 -9850 41980
rect -9650 41910 -9350 41980
rect -9150 41910 -8850 41980
rect -8650 41910 -8350 41980
rect -8150 41910 -7850 41980
rect -7650 41910 -7350 41980
rect -7150 41910 -6850 41980
rect -6650 41910 -6350 41980
rect -6150 41910 -5850 41980
rect -5650 41910 -5350 41980
rect -5150 41910 -4850 41980
rect -4650 41910 -4350 41980
rect -4150 41910 -3850 41980
rect -3650 41910 -3350 41980
rect -3150 41910 -2850 41980
rect -2650 41910 -2350 41980
rect -2150 41910 -1850 41980
rect -1650 41910 -1350 41980
rect -1150 41910 -850 41980
rect -650 41910 -350 41980
rect -150 41910 150 41980
rect 350 41910 650 41980
rect 850 41910 1150 41980
rect 1350 41910 1650 41980
rect 1850 41910 2150 41980
rect 2350 41910 2650 41980
rect 2850 41910 3150 41980
rect 3350 41910 3650 41980
rect 3850 41910 4000 41980
rect -16000 41900 4000 41910
rect -16000 41880 -15880 41900
rect -15620 41880 -15380 41900
rect -15120 41880 -14880 41900
rect -14620 41880 -14380 41900
rect -14120 41880 -13880 41900
rect -13620 41880 -13380 41900
rect -13120 41880 -12880 41900
rect -12620 41880 -12380 41900
rect -12120 41880 -11880 41900
rect -11620 41880 -11380 41900
rect -11120 41880 -10880 41900
rect -10620 41880 -10380 41900
rect -10120 41880 -9880 41900
rect -9620 41880 -9380 41900
rect -9120 41880 -8880 41900
rect -8620 41880 -8380 41900
rect -8120 41880 -7880 41900
rect -7620 41880 -7380 41900
rect -7120 41880 -6880 41900
rect -6620 41880 -6380 41900
rect -6120 41880 -5880 41900
rect -5620 41880 -5380 41900
rect -5120 41880 -4880 41900
rect -4620 41880 -4380 41900
rect -4120 41880 -3880 41900
rect -3620 41880 -3380 41900
rect -3120 41880 -2880 41900
rect -2620 41880 -2380 41900
rect -2120 41880 -1880 41900
rect -1620 41880 -1380 41900
rect -1120 41880 -880 41900
rect -620 41880 -380 41900
rect -120 41880 120 41900
rect 380 41880 620 41900
rect 880 41880 1120 41900
rect 1380 41880 1620 41900
rect 1880 41880 2120 41900
rect 2380 41880 2620 41900
rect 2880 41880 3120 41900
rect 3380 41880 3620 41900
rect 3880 41880 4000 41900
rect -16000 41850 -15900 41880
rect -16000 41650 -15980 41850
rect -15910 41650 -15900 41850
rect -16000 41620 -15900 41650
rect -15600 41850 -15400 41880
rect -15600 41650 -15590 41850
rect -15520 41650 -15480 41850
rect -15410 41650 -15400 41850
rect -15600 41620 -15400 41650
rect -15100 41850 -14900 41880
rect -15100 41650 -15090 41850
rect -15020 41650 -14980 41850
rect -14910 41650 -14900 41850
rect -15100 41620 -14900 41650
rect -14600 41850 -14400 41880
rect -14600 41650 -14590 41850
rect -14520 41650 -14480 41850
rect -14410 41650 -14400 41850
rect -14600 41620 -14400 41650
rect -14100 41850 -13900 41880
rect -14100 41650 -14090 41850
rect -14020 41650 -13980 41850
rect -13910 41650 -13900 41850
rect -14100 41620 -13900 41650
rect -13600 41850 -13400 41880
rect -13600 41650 -13590 41850
rect -13520 41650 -13480 41850
rect -13410 41650 -13400 41850
rect -13600 41620 -13400 41650
rect -13100 41850 -12900 41880
rect -13100 41650 -13090 41850
rect -13020 41650 -12980 41850
rect -12910 41650 -12900 41850
rect -13100 41620 -12900 41650
rect -12600 41850 -12400 41880
rect -12600 41650 -12590 41850
rect -12520 41650 -12480 41850
rect -12410 41650 -12400 41850
rect -12600 41620 -12400 41650
rect -12100 41850 -11900 41880
rect -12100 41650 -12090 41850
rect -12020 41650 -11980 41850
rect -11910 41650 -11900 41850
rect -12100 41620 -11900 41650
rect -11600 41850 -11400 41880
rect -11600 41650 -11590 41850
rect -11520 41650 -11480 41850
rect -11410 41650 -11400 41850
rect -11600 41620 -11400 41650
rect -11100 41850 -10900 41880
rect -11100 41650 -11090 41850
rect -11020 41650 -10980 41850
rect -10910 41650 -10900 41850
rect -11100 41620 -10900 41650
rect -10600 41850 -10400 41880
rect -10600 41650 -10590 41850
rect -10520 41650 -10480 41850
rect -10410 41650 -10400 41850
rect -10600 41620 -10400 41650
rect -10100 41850 -9900 41880
rect -10100 41650 -10090 41850
rect -10020 41650 -9980 41850
rect -9910 41650 -9900 41850
rect -10100 41620 -9900 41650
rect -9600 41850 -9400 41880
rect -9600 41650 -9590 41850
rect -9520 41650 -9480 41850
rect -9410 41650 -9400 41850
rect -9600 41620 -9400 41650
rect -9100 41850 -8900 41880
rect -9100 41650 -9090 41850
rect -9020 41650 -8980 41850
rect -8910 41650 -8900 41850
rect -9100 41620 -8900 41650
rect -8600 41850 -8400 41880
rect -8600 41650 -8590 41850
rect -8520 41650 -8480 41850
rect -8410 41650 -8400 41850
rect -8600 41620 -8400 41650
rect -8100 41850 -7900 41880
rect -8100 41650 -8090 41850
rect -8020 41650 -7980 41850
rect -7910 41650 -7900 41850
rect -8100 41620 -7900 41650
rect -7600 41850 -7400 41880
rect -7600 41650 -7590 41850
rect -7520 41650 -7480 41850
rect -7410 41650 -7400 41850
rect -7600 41620 -7400 41650
rect -7100 41850 -6900 41880
rect -7100 41650 -7090 41850
rect -7020 41650 -6980 41850
rect -6910 41650 -6900 41850
rect -7100 41620 -6900 41650
rect -6600 41850 -6400 41880
rect -6600 41650 -6590 41850
rect -6520 41650 -6480 41850
rect -6410 41650 -6400 41850
rect -6600 41620 -6400 41650
rect -6100 41850 -5900 41880
rect -6100 41650 -6090 41850
rect -6020 41650 -5980 41850
rect -5910 41650 -5900 41850
rect -6100 41620 -5900 41650
rect -5600 41850 -5400 41880
rect -5600 41650 -5590 41850
rect -5520 41650 -5480 41850
rect -5410 41650 -5400 41850
rect -5600 41620 -5400 41650
rect -5100 41850 -4900 41880
rect -5100 41650 -5090 41850
rect -5020 41650 -4980 41850
rect -4910 41650 -4900 41850
rect -5100 41620 -4900 41650
rect -4600 41850 -4400 41880
rect -4600 41650 -4590 41850
rect -4520 41650 -4480 41850
rect -4410 41650 -4400 41850
rect -4600 41620 -4400 41650
rect -4100 41850 -3900 41880
rect -4100 41650 -4090 41850
rect -4020 41650 -3980 41850
rect -3910 41650 -3900 41850
rect -4100 41620 -3900 41650
rect -3600 41850 -3400 41880
rect -3600 41650 -3590 41850
rect -3520 41650 -3480 41850
rect -3410 41650 -3400 41850
rect -3600 41620 -3400 41650
rect -3100 41850 -2900 41880
rect -3100 41650 -3090 41850
rect -3020 41650 -2980 41850
rect -2910 41650 -2900 41850
rect -3100 41620 -2900 41650
rect -2600 41850 -2400 41880
rect -2600 41650 -2590 41850
rect -2520 41650 -2480 41850
rect -2410 41650 -2400 41850
rect -2600 41620 -2400 41650
rect -2100 41850 -1900 41880
rect -2100 41650 -2090 41850
rect -2020 41650 -1980 41850
rect -1910 41650 -1900 41850
rect -2100 41620 -1900 41650
rect -1600 41850 -1400 41880
rect -1600 41650 -1590 41850
rect -1520 41650 -1480 41850
rect -1410 41650 -1400 41850
rect -1600 41620 -1400 41650
rect -1100 41850 -900 41880
rect -1100 41650 -1090 41850
rect -1020 41650 -980 41850
rect -910 41650 -900 41850
rect -1100 41620 -900 41650
rect -600 41850 -400 41880
rect -600 41650 -590 41850
rect -520 41650 -480 41850
rect -410 41650 -400 41850
rect -600 41620 -400 41650
rect -100 41850 100 41880
rect -100 41650 -90 41850
rect -20 41650 20 41850
rect 90 41650 100 41850
rect -100 41620 100 41650
rect 400 41850 600 41880
rect 400 41650 410 41850
rect 480 41650 520 41850
rect 590 41650 600 41850
rect 400 41620 600 41650
rect 900 41850 1100 41880
rect 900 41650 910 41850
rect 980 41650 1020 41850
rect 1090 41650 1100 41850
rect 900 41620 1100 41650
rect 1400 41850 1600 41880
rect 1400 41650 1410 41850
rect 1480 41650 1520 41850
rect 1590 41650 1600 41850
rect 1400 41620 1600 41650
rect 1900 41850 2100 41880
rect 1900 41650 1910 41850
rect 1980 41650 2020 41850
rect 2090 41650 2100 41850
rect 1900 41620 2100 41650
rect 2400 41850 2600 41880
rect 2400 41650 2410 41850
rect 2480 41650 2520 41850
rect 2590 41650 2600 41850
rect 2400 41620 2600 41650
rect 2900 41850 3100 41880
rect 2900 41650 2910 41850
rect 2980 41650 3020 41850
rect 3090 41650 3100 41850
rect 2900 41620 3100 41650
rect 3400 41850 3600 41880
rect 3400 41650 3410 41850
rect 3480 41650 3520 41850
rect 3590 41650 3600 41850
rect 3400 41620 3600 41650
rect 3900 41850 4000 41880
rect 3900 41650 3910 41850
rect 3980 41650 4000 41850
rect 3900 41620 4000 41650
rect -16000 41600 -15880 41620
rect -15620 41600 -15380 41620
rect -15120 41600 -14880 41620
rect -14620 41600 -14380 41620
rect -14120 41600 -13880 41620
rect -13620 41600 -13380 41620
rect -13120 41600 -12880 41620
rect -12620 41600 -12380 41620
rect -12120 41600 -11880 41620
rect -11620 41600 -11380 41620
rect -11120 41600 -10880 41620
rect -10620 41600 -10380 41620
rect -10120 41600 -9880 41620
rect -9620 41600 -9380 41620
rect -9120 41600 -8880 41620
rect -8620 41600 -8380 41620
rect -8120 41600 -7880 41620
rect -7620 41600 -7380 41620
rect -7120 41600 -6880 41620
rect -6620 41600 -6380 41620
rect -6120 41600 -5880 41620
rect -5620 41600 -5380 41620
rect -5120 41600 -4880 41620
rect -4620 41600 -4380 41620
rect -4120 41600 -3880 41620
rect -3620 41600 -3380 41620
rect -3120 41600 -2880 41620
rect -2620 41600 -2380 41620
rect -2120 41600 -1880 41620
rect -1620 41600 -1380 41620
rect -1120 41600 -880 41620
rect -620 41600 -380 41620
rect -120 41600 120 41620
rect 380 41600 620 41620
rect 880 41600 1120 41620
rect 1380 41600 1620 41620
rect 1880 41600 2120 41620
rect 2380 41600 2620 41620
rect 2880 41600 3120 41620
rect 3380 41600 3620 41620
rect 3880 41600 4000 41620
rect -16000 41590 4000 41600
rect -16000 41520 -15850 41590
rect -15650 41520 -15350 41590
rect -15150 41520 -14850 41590
rect -14650 41520 -14350 41590
rect -14150 41520 -13850 41590
rect -13650 41520 -13350 41590
rect -13150 41520 -12850 41590
rect -12650 41520 -12350 41590
rect -12150 41520 -11850 41590
rect -11650 41520 -11350 41590
rect -11150 41520 -10850 41590
rect -10650 41520 -10350 41590
rect -10150 41520 -9850 41590
rect -9650 41520 -9350 41590
rect -9150 41520 -8850 41590
rect -8650 41520 -8350 41590
rect -8150 41520 -7850 41590
rect -7650 41520 -7350 41590
rect -7150 41520 -6850 41590
rect -6650 41520 -6350 41590
rect -6150 41520 -5850 41590
rect -5650 41520 -5350 41590
rect -5150 41520 -4850 41590
rect -4650 41520 -4350 41590
rect -4150 41520 -3850 41590
rect -3650 41520 -3350 41590
rect -3150 41520 -2850 41590
rect -2650 41520 -2350 41590
rect -2150 41520 -1850 41590
rect -1650 41520 -1350 41590
rect -1150 41520 -850 41590
rect -650 41520 -350 41590
rect -150 41520 150 41590
rect 350 41520 650 41590
rect 850 41520 1150 41590
rect 1350 41520 1650 41590
rect 1850 41520 2150 41590
rect 2350 41520 2650 41590
rect 2850 41520 3150 41590
rect 3350 41520 3650 41590
rect 3850 41520 4000 41590
rect -16000 41480 4000 41520
rect -16000 41410 -15850 41480
rect -15650 41410 -15350 41480
rect -15150 41410 -14850 41480
rect -14650 41410 -14350 41480
rect -14150 41410 -13850 41480
rect -13650 41410 -13350 41480
rect -13150 41410 -12850 41480
rect -12650 41410 -12350 41480
rect -12150 41410 -11850 41480
rect -11650 41410 -11350 41480
rect -11150 41410 -10850 41480
rect -10650 41410 -10350 41480
rect -10150 41410 -9850 41480
rect -9650 41410 -9350 41480
rect -9150 41410 -8850 41480
rect -8650 41410 -8350 41480
rect -8150 41410 -7850 41480
rect -7650 41410 -7350 41480
rect -7150 41410 -6850 41480
rect -6650 41410 -6350 41480
rect -6150 41410 -5850 41480
rect -5650 41410 -5350 41480
rect -5150 41410 -4850 41480
rect -4650 41410 -4350 41480
rect -4150 41410 -3850 41480
rect -3650 41410 -3350 41480
rect -3150 41410 -2850 41480
rect -2650 41410 -2350 41480
rect -2150 41410 -1850 41480
rect -1650 41410 -1350 41480
rect -1150 41410 -850 41480
rect -650 41410 -350 41480
rect -150 41410 150 41480
rect 350 41410 650 41480
rect 850 41410 1150 41480
rect 1350 41410 1650 41480
rect 1850 41410 2150 41480
rect 2350 41410 2650 41480
rect 2850 41410 3150 41480
rect 3350 41410 3650 41480
rect 3850 41410 4000 41480
rect -16000 41400 4000 41410
rect -16000 41380 -15880 41400
rect -15620 41380 -15380 41400
rect -15120 41380 -14880 41400
rect -14620 41380 -14380 41400
rect -14120 41380 -13880 41400
rect -13620 41380 -13380 41400
rect -13120 41380 -12880 41400
rect -12620 41380 -12380 41400
rect -12120 41380 -11880 41400
rect -11620 41380 -11380 41400
rect -11120 41380 -10880 41400
rect -10620 41380 -10380 41400
rect -10120 41380 -9880 41400
rect -9620 41380 -9380 41400
rect -9120 41380 -8880 41400
rect -8620 41380 -8380 41400
rect -8120 41380 -7880 41400
rect -7620 41380 -7380 41400
rect -7120 41380 -6880 41400
rect -6620 41380 -6380 41400
rect -6120 41380 -5880 41400
rect -5620 41380 -5380 41400
rect -5120 41380 -4880 41400
rect -4620 41380 -4380 41400
rect -4120 41380 -3880 41400
rect -3620 41380 -3380 41400
rect -3120 41380 -2880 41400
rect -2620 41380 -2380 41400
rect -2120 41380 -1880 41400
rect -1620 41380 -1380 41400
rect -1120 41380 -880 41400
rect -620 41380 -380 41400
rect -120 41380 120 41400
rect 380 41380 620 41400
rect 880 41380 1120 41400
rect 1380 41380 1620 41400
rect 1880 41380 2120 41400
rect 2380 41380 2620 41400
rect 2880 41380 3120 41400
rect 3380 41380 3620 41400
rect 3880 41380 4000 41400
rect -16000 41350 -15900 41380
rect -16000 41150 -15980 41350
rect -15910 41150 -15900 41350
rect -16000 41120 -15900 41150
rect -15600 41350 -15400 41380
rect -15600 41150 -15590 41350
rect -15520 41150 -15480 41350
rect -15410 41150 -15400 41350
rect -15600 41120 -15400 41150
rect -15100 41350 -14900 41380
rect -15100 41150 -15090 41350
rect -15020 41150 -14980 41350
rect -14910 41150 -14900 41350
rect -15100 41120 -14900 41150
rect -14600 41350 -14400 41380
rect -14600 41150 -14590 41350
rect -14520 41150 -14480 41350
rect -14410 41150 -14400 41350
rect -14600 41120 -14400 41150
rect -14100 41350 -13900 41380
rect -14100 41150 -14090 41350
rect -14020 41150 -13980 41350
rect -13910 41150 -13900 41350
rect -14100 41120 -13900 41150
rect -13600 41350 -13400 41380
rect -13600 41150 -13590 41350
rect -13520 41150 -13480 41350
rect -13410 41150 -13400 41350
rect -13600 41120 -13400 41150
rect -13100 41350 -12900 41380
rect -13100 41150 -13090 41350
rect -13020 41150 -12980 41350
rect -12910 41150 -12900 41350
rect -13100 41120 -12900 41150
rect -12600 41350 -12400 41380
rect -12600 41150 -12590 41350
rect -12520 41150 -12480 41350
rect -12410 41150 -12400 41350
rect -12600 41120 -12400 41150
rect -12100 41350 -11900 41380
rect -12100 41150 -12090 41350
rect -12020 41150 -11980 41350
rect -11910 41150 -11900 41350
rect -12100 41120 -11900 41150
rect -11600 41350 -11400 41380
rect -11600 41150 -11590 41350
rect -11520 41150 -11480 41350
rect -11410 41150 -11400 41350
rect -11600 41120 -11400 41150
rect -11100 41350 -10900 41380
rect -11100 41150 -11090 41350
rect -11020 41150 -10980 41350
rect -10910 41150 -10900 41350
rect -11100 41120 -10900 41150
rect -10600 41350 -10400 41380
rect -10600 41150 -10590 41350
rect -10520 41150 -10480 41350
rect -10410 41150 -10400 41350
rect -10600 41120 -10400 41150
rect -10100 41350 -9900 41380
rect -10100 41150 -10090 41350
rect -10020 41150 -9980 41350
rect -9910 41150 -9900 41350
rect -10100 41120 -9900 41150
rect -9600 41350 -9400 41380
rect -9600 41150 -9590 41350
rect -9520 41150 -9480 41350
rect -9410 41150 -9400 41350
rect -9600 41120 -9400 41150
rect -9100 41350 -8900 41380
rect -9100 41150 -9090 41350
rect -9020 41150 -8980 41350
rect -8910 41150 -8900 41350
rect -9100 41120 -8900 41150
rect -8600 41350 -8400 41380
rect -8600 41150 -8590 41350
rect -8520 41150 -8480 41350
rect -8410 41150 -8400 41350
rect -8600 41120 -8400 41150
rect -8100 41350 -7900 41380
rect -8100 41150 -8090 41350
rect -8020 41150 -7980 41350
rect -7910 41150 -7900 41350
rect -8100 41120 -7900 41150
rect -7600 41350 -7400 41380
rect -7600 41150 -7590 41350
rect -7520 41150 -7480 41350
rect -7410 41150 -7400 41350
rect -7600 41120 -7400 41150
rect -7100 41350 -6900 41380
rect -7100 41150 -7090 41350
rect -7020 41150 -6980 41350
rect -6910 41150 -6900 41350
rect -7100 41120 -6900 41150
rect -6600 41350 -6400 41380
rect -6600 41150 -6590 41350
rect -6520 41150 -6480 41350
rect -6410 41150 -6400 41350
rect -6600 41120 -6400 41150
rect -6100 41350 -5900 41380
rect -6100 41150 -6090 41350
rect -6020 41150 -5980 41350
rect -5910 41150 -5900 41350
rect -6100 41120 -5900 41150
rect -5600 41350 -5400 41380
rect -5600 41150 -5590 41350
rect -5520 41150 -5480 41350
rect -5410 41150 -5400 41350
rect -5600 41120 -5400 41150
rect -5100 41350 -4900 41380
rect -5100 41150 -5090 41350
rect -5020 41150 -4980 41350
rect -4910 41150 -4900 41350
rect -5100 41120 -4900 41150
rect -4600 41350 -4400 41380
rect -4600 41150 -4590 41350
rect -4520 41150 -4480 41350
rect -4410 41150 -4400 41350
rect -4600 41120 -4400 41150
rect -4100 41350 -3900 41380
rect -4100 41150 -4090 41350
rect -4020 41150 -3980 41350
rect -3910 41150 -3900 41350
rect -4100 41120 -3900 41150
rect -3600 41350 -3400 41380
rect -3600 41150 -3590 41350
rect -3520 41150 -3480 41350
rect -3410 41150 -3400 41350
rect -3600 41120 -3400 41150
rect -3100 41350 -2900 41380
rect -3100 41150 -3090 41350
rect -3020 41150 -2980 41350
rect -2910 41150 -2900 41350
rect -3100 41120 -2900 41150
rect -2600 41350 -2400 41380
rect -2600 41150 -2590 41350
rect -2520 41150 -2480 41350
rect -2410 41150 -2400 41350
rect -2600 41120 -2400 41150
rect -2100 41350 -1900 41380
rect -2100 41150 -2090 41350
rect -2020 41150 -1980 41350
rect -1910 41150 -1900 41350
rect -2100 41120 -1900 41150
rect -1600 41350 -1400 41380
rect -1600 41150 -1590 41350
rect -1520 41150 -1480 41350
rect -1410 41150 -1400 41350
rect -1600 41120 -1400 41150
rect -1100 41350 -900 41380
rect -1100 41150 -1090 41350
rect -1020 41150 -980 41350
rect -910 41150 -900 41350
rect -1100 41120 -900 41150
rect -600 41350 -400 41380
rect -600 41150 -590 41350
rect -520 41150 -480 41350
rect -410 41150 -400 41350
rect -600 41120 -400 41150
rect -100 41350 100 41380
rect -100 41150 -90 41350
rect -20 41150 20 41350
rect 90 41150 100 41350
rect -100 41120 100 41150
rect 400 41350 600 41380
rect 400 41150 410 41350
rect 480 41150 520 41350
rect 590 41150 600 41350
rect 400 41120 600 41150
rect 900 41350 1100 41380
rect 900 41150 910 41350
rect 980 41150 1020 41350
rect 1090 41150 1100 41350
rect 900 41120 1100 41150
rect 1400 41350 1600 41380
rect 1400 41150 1410 41350
rect 1480 41150 1520 41350
rect 1590 41150 1600 41350
rect 1400 41120 1600 41150
rect 1900 41350 2100 41380
rect 1900 41150 1910 41350
rect 1980 41150 2020 41350
rect 2090 41150 2100 41350
rect 1900 41120 2100 41150
rect 2400 41350 2600 41380
rect 2400 41150 2410 41350
rect 2480 41150 2520 41350
rect 2590 41150 2600 41350
rect 2400 41120 2600 41150
rect 2900 41350 3100 41380
rect 2900 41150 2910 41350
rect 2980 41150 3020 41350
rect 3090 41150 3100 41350
rect 2900 41120 3100 41150
rect 3400 41350 3600 41380
rect 3400 41150 3410 41350
rect 3480 41150 3520 41350
rect 3590 41150 3600 41350
rect 3400 41120 3600 41150
rect 3900 41350 4000 41380
rect 3900 41150 3910 41350
rect 3980 41150 4000 41350
rect 3900 41120 4000 41150
rect -16000 41100 -15880 41120
rect -15620 41100 -15380 41120
rect -15120 41100 -14880 41120
rect -14620 41100 -14380 41120
rect -14120 41100 -13880 41120
rect -13620 41100 -13380 41120
rect -13120 41100 -12880 41120
rect -12620 41100 -12380 41120
rect -12120 41100 -11880 41120
rect -11620 41100 -11380 41120
rect -11120 41100 -10880 41120
rect -10620 41100 -10380 41120
rect -10120 41100 -9880 41120
rect -9620 41100 -9380 41120
rect -9120 41100 -8880 41120
rect -8620 41100 -8380 41120
rect -8120 41100 -7880 41120
rect -7620 41100 -7380 41120
rect -7120 41100 -6880 41120
rect -6620 41100 -6380 41120
rect -6120 41100 -5880 41120
rect -5620 41100 -5380 41120
rect -5120 41100 -4880 41120
rect -4620 41100 -4380 41120
rect -4120 41100 -3880 41120
rect -3620 41100 -3380 41120
rect -3120 41100 -2880 41120
rect -2620 41100 -2380 41120
rect -2120 41100 -1880 41120
rect -1620 41100 -1380 41120
rect -1120 41100 -880 41120
rect -620 41100 -380 41120
rect -120 41100 120 41120
rect 380 41100 620 41120
rect 880 41100 1120 41120
rect 1380 41100 1620 41120
rect 1880 41100 2120 41120
rect 2380 41100 2620 41120
rect 2880 41100 3120 41120
rect 3380 41100 3620 41120
rect 3880 41100 4000 41120
rect -16000 41090 4000 41100
rect -16000 41020 -15850 41090
rect -15650 41020 -15350 41090
rect -15150 41020 -14850 41090
rect -14650 41020 -14350 41090
rect -14150 41020 -13850 41090
rect -13650 41020 -13350 41090
rect -13150 41020 -12850 41090
rect -12650 41020 -12350 41090
rect -12150 41020 -11850 41090
rect -11650 41020 -11350 41090
rect -11150 41020 -10850 41090
rect -10650 41020 -10350 41090
rect -10150 41020 -9850 41090
rect -9650 41020 -9350 41090
rect -9150 41020 -8850 41090
rect -8650 41020 -8350 41090
rect -8150 41020 -7850 41090
rect -7650 41020 -7350 41090
rect -7150 41020 -6850 41090
rect -6650 41020 -6350 41090
rect -6150 41020 -5850 41090
rect -5650 41020 -5350 41090
rect -5150 41020 -4850 41090
rect -4650 41020 -4350 41090
rect -4150 41020 -3850 41090
rect -3650 41020 -3350 41090
rect -3150 41020 -2850 41090
rect -2650 41020 -2350 41090
rect -2150 41020 -1850 41090
rect -1650 41020 -1350 41090
rect -1150 41020 -850 41090
rect -650 41020 -350 41090
rect -150 41020 150 41090
rect 350 41020 650 41090
rect 850 41020 1150 41090
rect 1350 41020 1650 41090
rect 1850 41020 2150 41090
rect 2350 41020 2650 41090
rect 2850 41020 3150 41090
rect 3350 41020 3650 41090
rect 3850 41020 4000 41090
rect -16000 40980 4000 41020
rect -16000 40910 -15850 40980
rect -15650 40910 -15350 40980
rect -15150 40910 -14850 40980
rect -14650 40910 -14350 40980
rect -14150 40910 -13850 40980
rect -13650 40910 -13350 40980
rect -13150 40910 -12850 40980
rect -12650 40910 -12350 40980
rect -12150 40910 -11850 40980
rect -11650 40910 -11350 40980
rect -11150 40910 -10850 40980
rect -10650 40910 -10350 40980
rect -10150 40910 -9850 40980
rect -9650 40910 -9350 40980
rect -9150 40910 -8850 40980
rect -8650 40910 -8350 40980
rect -8150 40910 -7850 40980
rect -7650 40910 -7350 40980
rect -7150 40910 -6850 40980
rect -6650 40910 -6350 40980
rect -6150 40910 -5850 40980
rect -5650 40910 -5350 40980
rect -5150 40910 -4850 40980
rect -4650 40910 -4350 40980
rect -4150 40910 -3850 40980
rect -3650 40910 -3350 40980
rect -3150 40910 -2850 40980
rect -2650 40910 -2350 40980
rect -2150 40910 -1850 40980
rect -1650 40910 -1350 40980
rect -1150 40910 -850 40980
rect -650 40910 -350 40980
rect -150 40910 150 40980
rect 350 40910 650 40980
rect 850 40910 1150 40980
rect 1350 40910 1650 40980
rect 1850 40910 2150 40980
rect 2350 40910 2650 40980
rect 2850 40910 3150 40980
rect 3350 40910 3650 40980
rect 3850 40910 4000 40980
rect -16000 40900 4000 40910
rect -16000 40880 -15880 40900
rect -15620 40880 -15380 40900
rect -15120 40880 -14880 40900
rect -14620 40880 -14380 40900
rect -14120 40880 -13880 40900
rect -13620 40880 -13380 40900
rect -13120 40880 -12880 40900
rect -12620 40880 -12380 40900
rect -12120 40880 -11880 40900
rect -11620 40880 -11380 40900
rect -11120 40880 -10880 40900
rect -10620 40880 -10380 40900
rect -10120 40880 -9880 40900
rect -9620 40880 -9380 40900
rect -9120 40880 -8880 40900
rect -8620 40880 -8380 40900
rect -8120 40880 -7880 40900
rect -7620 40880 -7380 40900
rect -7120 40880 -6880 40900
rect -6620 40880 -6380 40900
rect -6120 40880 -5880 40900
rect -5620 40880 -5380 40900
rect -5120 40880 -4880 40900
rect -4620 40880 -4380 40900
rect -4120 40880 -3880 40900
rect -3620 40880 -3380 40900
rect -3120 40880 -2880 40900
rect -2620 40880 -2380 40900
rect -2120 40880 -1880 40900
rect -1620 40880 -1380 40900
rect -1120 40880 -880 40900
rect -620 40880 -380 40900
rect -120 40880 120 40900
rect 380 40880 620 40900
rect 880 40880 1120 40900
rect 1380 40880 1620 40900
rect 1880 40880 2120 40900
rect 2380 40880 2620 40900
rect 2880 40880 3120 40900
rect 3380 40880 3620 40900
rect 3880 40880 4000 40900
rect -16000 40850 -15900 40880
rect -16000 40650 -15980 40850
rect -15910 40650 -15900 40850
rect -16000 40620 -15900 40650
rect -15600 40850 -15400 40880
rect -15600 40650 -15590 40850
rect -15520 40650 -15480 40850
rect -15410 40650 -15400 40850
rect -15600 40620 -15400 40650
rect -15100 40850 -14900 40880
rect -15100 40650 -15090 40850
rect -15020 40650 -14980 40850
rect -14910 40650 -14900 40850
rect -15100 40620 -14900 40650
rect -14600 40850 -14400 40880
rect -14600 40650 -14590 40850
rect -14520 40650 -14480 40850
rect -14410 40650 -14400 40850
rect -14600 40620 -14400 40650
rect -14100 40850 -13900 40880
rect -14100 40650 -14090 40850
rect -14020 40650 -13980 40850
rect -13910 40650 -13900 40850
rect -14100 40620 -13900 40650
rect -13600 40850 -13400 40880
rect -13600 40650 -13590 40850
rect -13520 40650 -13480 40850
rect -13410 40650 -13400 40850
rect -13600 40620 -13400 40650
rect -13100 40850 -12900 40880
rect -13100 40650 -13090 40850
rect -13020 40650 -12980 40850
rect -12910 40650 -12900 40850
rect -13100 40620 -12900 40650
rect -12600 40850 -12400 40880
rect -12600 40650 -12590 40850
rect -12520 40650 -12480 40850
rect -12410 40650 -12400 40850
rect -12600 40620 -12400 40650
rect -12100 40850 -11900 40880
rect -12100 40650 -12090 40850
rect -12020 40650 -11980 40850
rect -11910 40650 -11900 40850
rect -12100 40620 -11900 40650
rect -11600 40850 -11400 40880
rect -11600 40650 -11590 40850
rect -11520 40650 -11480 40850
rect -11410 40650 -11400 40850
rect -11600 40620 -11400 40650
rect -11100 40850 -10900 40880
rect -11100 40650 -11090 40850
rect -11020 40650 -10980 40850
rect -10910 40650 -10900 40850
rect -11100 40620 -10900 40650
rect -10600 40850 -10400 40880
rect -10600 40650 -10590 40850
rect -10520 40650 -10480 40850
rect -10410 40650 -10400 40850
rect -10600 40620 -10400 40650
rect -10100 40850 -9900 40880
rect -10100 40650 -10090 40850
rect -10020 40650 -9980 40850
rect -9910 40650 -9900 40850
rect -10100 40620 -9900 40650
rect -9600 40850 -9400 40880
rect -9600 40650 -9590 40850
rect -9520 40650 -9480 40850
rect -9410 40650 -9400 40850
rect -9600 40620 -9400 40650
rect -9100 40850 -8900 40880
rect -9100 40650 -9090 40850
rect -9020 40650 -8980 40850
rect -8910 40650 -8900 40850
rect -9100 40620 -8900 40650
rect -8600 40850 -8400 40880
rect -8600 40650 -8590 40850
rect -8520 40650 -8480 40850
rect -8410 40650 -8400 40850
rect -8600 40620 -8400 40650
rect -8100 40850 -7900 40880
rect -8100 40650 -8090 40850
rect -8020 40650 -7980 40850
rect -7910 40650 -7900 40850
rect -8100 40620 -7900 40650
rect -7600 40850 -7400 40880
rect -7600 40650 -7590 40850
rect -7520 40650 -7480 40850
rect -7410 40650 -7400 40850
rect -7600 40620 -7400 40650
rect -7100 40850 -6900 40880
rect -7100 40650 -7090 40850
rect -7020 40650 -6980 40850
rect -6910 40650 -6900 40850
rect -7100 40620 -6900 40650
rect -6600 40850 -6400 40880
rect -6600 40650 -6590 40850
rect -6520 40650 -6480 40850
rect -6410 40650 -6400 40850
rect -6600 40620 -6400 40650
rect -6100 40850 -5900 40880
rect -6100 40650 -6090 40850
rect -6020 40650 -5980 40850
rect -5910 40650 -5900 40850
rect -6100 40620 -5900 40650
rect -5600 40850 -5400 40880
rect -5600 40650 -5590 40850
rect -5520 40650 -5480 40850
rect -5410 40650 -5400 40850
rect -5600 40620 -5400 40650
rect -5100 40850 -4900 40880
rect -5100 40650 -5090 40850
rect -5020 40650 -4980 40850
rect -4910 40650 -4900 40850
rect -5100 40620 -4900 40650
rect -4600 40850 -4400 40880
rect -4600 40650 -4590 40850
rect -4520 40650 -4480 40850
rect -4410 40650 -4400 40850
rect -4600 40620 -4400 40650
rect -4100 40850 -3900 40880
rect -4100 40650 -4090 40850
rect -4020 40650 -3980 40850
rect -3910 40650 -3900 40850
rect -4100 40620 -3900 40650
rect -3600 40850 -3400 40880
rect -3600 40650 -3590 40850
rect -3520 40650 -3480 40850
rect -3410 40650 -3400 40850
rect -3600 40620 -3400 40650
rect -3100 40850 -2900 40880
rect -3100 40650 -3090 40850
rect -3020 40650 -2980 40850
rect -2910 40650 -2900 40850
rect -3100 40620 -2900 40650
rect -2600 40850 -2400 40880
rect -2600 40650 -2590 40850
rect -2520 40650 -2480 40850
rect -2410 40650 -2400 40850
rect -2600 40620 -2400 40650
rect -2100 40850 -1900 40880
rect -2100 40650 -2090 40850
rect -2020 40650 -1980 40850
rect -1910 40650 -1900 40850
rect -2100 40620 -1900 40650
rect -1600 40850 -1400 40880
rect -1600 40650 -1590 40850
rect -1520 40650 -1480 40850
rect -1410 40650 -1400 40850
rect -1600 40620 -1400 40650
rect -1100 40850 -900 40880
rect -1100 40650 -1090 40850
rect -1020 40650 -980 40850
rect -910 40650 -900 40850
rect -1100 40620 -900 40650
rect -600 40850 -400 40880
rect -600 40650 -590 40850
rect -520 40650 -480 40850
rect -410 40650 -400 40850
rect -600 40620 -400 40650
rect -100 40850 100 40880
rect -100 40650 -90 40850
rect -20 40650 20 40850
rect 90 40650 100 40850
rect -100 40620 100 40650
rect 400 40850 600 40880
rect 400 40650 410 40850
rect 480 40650 520 40850
rect 590 40650 600 40850
rect 400 40620 600 40650
rect 900 40850 1100 40880
rect 900 40650 910 40850
rect 980 40650 1020 40850
rect 1090 40650 1100 40850
rect 900 40620 1100 40650
rect 1400 40850 1600 40880
rect 1400 40650 1410 40850
rect 1480 40650 1520 40850
rect 1590 40650 1600 40850
rect 1400 40620 1600 40650
rect 1900 40850 2100 40880
rect 1900 40650 1910 40850
rect 1980 40650 2020 40850
rect 2090 40650 2100 40850
rect 1900 40620 2100 40650
rect 2400 40850 2600 40880
rect 2400 40650 2410 40850
rect 2480 40650 2520 40850
rect 2590 40650 2600 40850
rect 2400 40620 2600 40650
rect 2900 40850 3100 40880
rect 2900 40650 2910 40850
rect 2980 40650 3020 40850
rect 3090 40650 3100 40850
rect 2900 40620 3100 40650
rect 3400 40850 3600 40880
rect 3400 40650 3410 40850
rect 3480 40650 3520 40850
rect 3590 40650 3600 40850
rect 3400 40620 3600 40650
rect 3900 40850 4000 40880
rect 3900 40650 3910 40850
rect 3980 40650 4000 40850
rect 3900 40620 4000 40650
rect -16000 40600 -15880 40620
rect -15620 40600 -15380 40620
rect -15120 40600 -14880 40620
rect -14620 40600 -14380 40620
rect -14120 40600 -13880 40620
rect -13620 40600 -13380 40620
rect -13120 40600 -12880 40620
rect -12620 40600 -12380 40620
rect -12120 40600 -11880 40620
rect -11620 40600 -11380 40620
rect -11120 40600 -10880 40620
rect -10620 40600 -10380 40620
rect -10120 40600 -9880 40620
rect -9620 40600 -9380 40620
rect -9120 40600 -8880 40620
rect -8620 40600 -8380 40620
rect -8120 40600 -7880 40620
rect -7620 40600 -7380 40620
rect -7120 40600 -6880 40620
rect -6620 40600 -6380 40620
rect -6120 40600 -5880 40620
rect -5620 40600 -5380 40620
rect -5120 40600 -4880 40620
rect -4620 40600 -4380 40620
rect -4120 40600 -3880 40620
rect -3620 40600 -3380 40620
rect -3120 40600 -2880 40620
rect -2620 40600 -2380 40620
rect -2120 40600 -1880 40620
rect -1620 40600 -1380 40620
rect -1120 40600 -880 40620
rect -620 40600 -380 40620
rect -120 40600 120 40620
rect 380 40600 620 40620
rect 880 40600 1120 40620
rect 1380 40600 1620 40620
rect 1880 40600 2120 40620
rect 2380 40600 2620 40620
rect 2880 40600 3120 40620
rect 3380 40600 3620 40620
rect 3880 40600 4000 40620
rect -16000 40590 4000 40600
rect -16000 40520 -15850 40590
rect -15650 40520 -15350 40590
rect -15150 40520 -14850 40590
rect -14650 40520 -14350 40590
rect -14150 40520 -13850 40590
rect -13650 40520 -13350 40590
rect -13150 40520 -12850 40590
rect -12650 40520 -12350 40590
rect -12150 40520 -11850 40590
rect -11650 40520 -11350 40590
rect -11150 40520 -10850 40590
rect -10650 40520 -10350 40590
rect -10150 40520 -9850 40590
rect -9650 40520 -9350 40590
rect -9150 40520 -8850 40590
rect -8650 40520 -8350 40590
rect -8150 40520 -7850 40590
rect -7650 40520 -7350 40590
rect -7150 40520 -6850 40590
rect -6650 40520 -6350 40590
rect -6150 40520 -5850 40590
rect -5650 40520 -5350 40590
rect -5150 40520 -4850 40590
rect -4650 40520 -4350 40590
rect -4150 40520 -3850 40590
rect -3650 40520 -3350 40590
rect -3150 40520 -2850 40590
rect -2650 40520 -2350 40590
rect -2150 40520 -1850 40590
rect -1650 40520 -1350 40590
rect -1150 40520 -850 40590
rect -650 40520 -350 40590
rect -150 40520 150 40590
rect 350 40520 650 40590
rect 850 40520 1150 40590
rect 1350 40520 1650 40590
rect 1850 40520 2150 40590
rect 2350 40520 2650 40590
rect 2850 40520 3150 40590
rect 3350 40520 3650 40590
rect 3850 40520 4000 40590
rect -16000 40480 4000 40520
rect -16000 40410 -15850 40480
rect -15650 40410 -15350 40480
rect -15150 40410 -14850 40480
rect -14650 40410 -14350 40480
rect -14150 40410 -13850 40480
rect -13650 40410 -13350 40480
rect -13150 40410 -12850 40480
rect -12650 40410 -12350 40480
rect -12150 40410 -11850 40480
rect -11650 40410 -11350 40480
rect -11150 40410 -10850 40480
rect -10650 40410 -10350 40480
rect -10150 40410 -9850 40480
rect -9650 40410 -9350 40480
rect -9150 40410 -8850 40480
rect -8650 40410 -8350 40480
rect -8150 40410 -7850 40480
rect -7650 40410 -7350 40480
rect -7150 40410 -6850 40480
rect -6650 40410 -6350 40480
rect -6150 40410 -5850 40480
rect -5650 40410 -5350 40480
rect -5150 40410 -4850 40480
rect -4650 40410 -4350 40480
rect -4150 40410 -3850 40480
rect -3650 40410 -3350 40480
rect -3150 40410 -2850 40480
rect -2650 40410 -2350 40480
rect -2150 40410 -1850 40480
rect -1650 40410 -1350 40480
rect -1150 40410 -850 40480
rect -650 40410 -350 40480
rect -150 40410 150 40480
rect 350 40410 650 40480
rect 850 40410 1150 40480
rect 1350 40410 1650 40480
rect 1850 40410 2150 40480
rect 2350 40410 2650 40480
rect 2850 40410 3150 40480
rect 3350 40410 3650 40480
rect 3850 40410 4000 40480
rect -16000 40400 4000 40410
rect -16000 40380 -15880 40400
rect -15620 40380 -15380 40400
rect -15120 40380 -14880 40400
rect -14620 40380 -14380 40400
rect -14120 40380 -13880 40400
rect -13620 40380 -13380 40400
rect -13120 40380 -12880 40400
rect -12620 40380 -12380 40400
rect -12120 40380 -11880 40400
rect -11620 40380 -11380 40400
rect -11120 40380 -10880 40400
rect -10620 40380 -10380 40400
rect -10120 40380 -9880 40400
rect -9620 40380 -9380 40400
rect -9120 40380 -8880 40400
rect -8620 40380 -8380 40400
rect -8120 40380 -7880 40400
rect -7620 40380 -7380 40400
rect -7120 40380 -6880 40400
rect -6620 40380 -6380 40400
rect -6120 40380 -5880 40400
rect -5620 40380 -5380 40400
rect -5120 40380 -4880 40400
rect -4620 40380 -4380 40400
rect -4120 40380 -3880 40400
rect -3620 40380 -3380 40400
rect -3120 40380 -2880 40400
rect -2620 40380 -2380 40400
rect -2120 40380 -1880 40400
rect -1620 40380 -1380 40400
rect -1120 40380 -880 40400
rect -620 40380 -380 40400
rect -120 40380 120 40400
rect 380 40380 620 40400
rect 880 40380 1120 40400
rect 1380 40380 1620 40400
rect 1880 40380 2120 40400
rect 2380 40380 2620 40400
rect 2880 40380 3120 40400
rect 3380 40380 3620 40400
rect 3880 40380 4000 40400
rect -16000 40350 -15900 40380
rect -16000 40150 -15980 40350
rect -15910 40150 -15900 40350
rect -16000 40120 -15900 40150
rect -15600 40350 -15400 40380
rect -15600 40150 -15590 40350
rect -15520 40150 -15480 40350
rect -15410 40150 -15400 40350
rect -15600 40120 -15400 40150
rect -15100 40350 -14900 40380
rect -15100 40150 -15090 40350
rect -15020 40150 -14980 40350
rect -14910 40150 -14900 40350
rect -15100 40120 -14900 40150
rect -14600 40350 -14400 40380
rect -14600 40150 -14590 40350
rect -14520 40150 -14480 40350
rect -14410 40150 -14400 40350
rect -14600 40120 -14400 40150
rect -14100 40350 -13900 40380
rect -14100 40150 -14090 40350
rect -14020 40150 -13980 40350
rect -13910 40150 -13900 40350
rect -14100 40120 -13900 40150
rect -13600 40350 -13400 40380
rect -13600 40150 -13590 40350
rect -13520 40150 -13480 40350
rect -13410 40150 -13400 40350
rect -13600 40120 -13400 40150
rect -13100 40350 -12900 40380
rect -13100 40150 -13090 40350
rect -13020 40150 -12980 40350
rect -12910 40150 -12900 40350
rect -13100 40120 -12900 40150
rect -12600 40350 -12400 40380
rect -12600 40150 -12590 40350
rect -12520 40150 -12480 40350
rect -12410 40150 -12400 40350
rect -12600 40120 -12400 40150
rect -12100 40350 -11900 40380
rect -12100 40150 -12090 40350
rect -12020 40150 -11980 40350
rect -11910 40150 -11900 40350
rect -12100 40120 -11900 40150
rect -11600 40350 -11400 40380
rect -11600 40150 -11590 40350
rect -11520 40150 -11480 40350
rect -11410 40150 -11400 40350
rect -11600 40120 -11400 40150
rect -11100 40350 -10900 40380
rect -11100 40150 -11090 40350
rect -11020 40150 -10980 40350
rect -10910 40150 -10900 40350
rect -11100 40120 -10900 40150
rect -10600 40350 -10400 40380
rect -10600 40150 -10590 40350
rect -10520 40150 -10480 40350
rect -10410 40150 -10400 40350
rect -10600 40120 -10400 40150
rect -10100 40350 -9900 40380
rect -10100 40150 -10090 40350
rect -10020 40150 -9980 40350
rect -9910 40150 -9900 40350
rect -10100 40120 -9900 40150
rect -9600 40350 -9400 40380
rect -9600 40150 -9590 40350
rect -9520 40150 -9480 40350
rect -9410 40150 -9400 40350
rect -9600 40120 -9400 40150
rect -9100 40350 -8900 40380
rect -9100 40150 -9090 40350
rect -9020 40150 -8980 40350
rect -8910 40150 -8900 40350
rect -9100 40120 -8900 40150
rect -8600 40350 -8400 40380
rect -8600 40150 -8590 40350
rect -8520 40150 -8480 40350
rect -8410 40150 -8400 40350
rect -8600 40120 -8400 40150
rect -8100 40350 -7900 40380
rect -8100 40150 -8090 40350
rect -8020 40150 -7980 40350
rect -7910 40150 -7900 40350
rect -8100 40120 -7900 40150
rect -7600 40350 -7400 40380
rect -7600 40150 -7590 40350
rect -7520 40150 -7480 40350
rect -7410 40150 -7400 40350
rect -7600 40120 -7400 40150
rect -7100 40350 -6900 40380
rect -7100 40150 -7090 40350
rect -7020 40150 -6980 40350
rect -6910 40150 -6900 40350
rect -7100 40120 -6900 40150
rect -6600 40350 -6400 40380
rect -6600 40150 -6590 40350
rect -6520 40150 -6480 40350
rect -6410 40150 -6400 40350
rect -6600 40120 -6400 40150
rect -6100 40350 -5900 40380
rect -6100 40150 -6090 40350
rect -6020 40150 -5980 40350
rect -5910 40150 -5900 40350
rect -6100 40120 -5900 40150
rect -5600 40350 -5400 40380
rect -5600 40150 -5590 40350
rect -5520 40150 -5480 40350
rect -5410 40150 -5400 40350
rect -5600 40120 -5400 40150
rect -5100 40350 -4900 40380
rect -5100 40150 -5090 40350
rect -5020 40150 -4980 40350
rect -4910 40150 -4900 40350
rect -5100 40120 -4900 40150
rect -4600 40350 -4400 40380
rect -4600 40150 -4590 40350
rect -4520 40150 -4480 40350
rect -4410 40150 -4400 40350
rect -4600 40120 -4400 40150
rect -4100 40350 -3900 40380
rect -4100 40150 -4090 40350
rect -4020 40150 -3980 40350
rect -3910 40150 -3900 40350
rect -4100 40120 -3900 40150
rect -3600 40350 -3400 40380
rect -3600 40150 -3590 40350
rect -3520 40150 -3480 40350
rect -3410 40150 -3400 40350
rect -3600 40120 -3400 40150
rect -3100 40350 -2900 40380
rect -3100 40150 -3090 40350
rect -3020 40150 -2980 40350
rect -2910 40150 -2900 40350
rect -3100 40120 -2900 40150
rect -2600 40350 -2400 40380
rect -2600 40150 -2590 40350
rect -2520 40150 -2480 40350
rect -2410 40150 -2400 40350
rect -2600 40120 -2400 40150
rect -2100 40350 -1900 40380
rect -2100 40150 -2090 40350
rect -2020 40150 -1980 40350
rect -1910 40150 -1900 40350
rect -2100 40120 -1900 40150
rect -1600 40350 -1400 40380
rect -1600 40150 -1590 40350
rect -1520 40150 -1480 40350
rect -1410 40150 -1400 40350
rect -1600 40120 -1400 40150
rect -1100 40350 -900 40380
rect -1100 40150 -1090 40350
rect -1020 40150 -980 40350
rect -910 40150 -900 40350
rect -1100 40120 -900 40150
rect -600 40350 -400 40380
rect -600 40150 -590 40350
rect -520 40150 -480 40350
rect -410 40150 -400 40350
rect -600 40120 -400 40150
rect -100 40350 100 40380
rect -100 40150 -90 40350
rect -20 40150 20 40350
rect 90 40150 100 40350
rect -100 40120 100 40150
rect 400 40350 600 40380
rect 400 40150 410 40350
rect 480 40150 520 40350
rect 590 40150 600 40350
rect 400 40120 600 40150
rect 900 40350 1100 40380
rect 900 40150 910 40350
rect 980 40150 1020 40350
rect 1090 40150 1100 40350
rect 900 40120 1100 40150
rect 1400 40350 1600 40380
rect 1400 40150 1410 40350
rect 1480 40150 1520 40350
rect 1590 40150 1600 40350
rect 1400 40120 1600 40150
rect 1900 40350 2100 40380
rect 1900 40150 1910 40350
rect 1980 40150 2020 40350
rect 2090 40150 2100 40350
rect 1900 40120 2100 40150
rect 2400 40350 2600 40380
rect 2400 40150 2410 40350
rect 2480 40150 2520 40350
rect 2590 40150 2600 40350
rect 2400 40120 2600 40150
rect 2900 40350 3100 40380
rect 2900 40150 2910 40350
rect 2980 40150 3020 40350
rect 3090 40150 3100 40350
rect 2900 40120 3100 40150
rect 3400 40350 3600 40380
rect 3400 40150 3410 40350
rect 3480 40150 3520 40350
rect 3590 40150 3600 40350
rect 3400 40120 3600 40150
rect 3900 40350 4000 40380
rect 3900 40150 3910 40350
rect 3980 40150 4000 40350
rect 3900 40120 4000 40150
rect -16000 40100 -15880 40120
rect -15620 40100 -15380 40120
rect -15120 40100 -14880 40120
rect -14620 40100 -14380 40120
rect -14120 40100 -13880 40120
rect -13620 40100 -13380 40120
rect -13120 40100 -12880 40120
rect -12620 40100 -12380 40120
rect -12120 40100 -11880 40120
rect -11620 40100 -11380 40120
rect -11120 40100 -10880 40120
rect -10620 40100 -10380 40120
rect -10120 40100 -9880 40120
rect -9620 40100 -9380 40120
rect -9120 40100 -8880 40120
rect -8620 40100 -8380 40120
rect -8120 40100 -7880 40120
rect -7620 40100 -7380 40120
rect -7120 40100 -6880 40120
rect -6620 40100 -6380 40120
rect -6120 40100 -5880 40120
rect -5620 40100 -5380 40120
rect -5120 40100 -4880 40120
rect -4620 40100 -4380 40120
rect -4120 40100 -3880 40120
rect -3620 40100 -3380 40120
rect -3120 40100 -2880 40120
rect -2620 40100 -2380 40120
rect -2120 40100 -1880 40120
rect -1620 40100 -1380 40120
rect -1120 40100 -880 40120
rect -620 40100 -380 40120
rect -120 40100 120 40120
rect 380 40100 620 40120
rect 880 40100 1120 40120
rect 1380 40100 1620 40120
rect 1880 40100 2120 40120
rect 2380 40100 2620 40120
rect 2880 40100 3120 40120
rect 3380 40100 3620 40120
rect 3880 40100 4000 40120
rect -16000 40090 4000 40100
rect -16000 40020 -15850 40090
rect -15650 40020 -15350 40090
rect -15150 40020 -14850 40090
rect -14650 40020 -14350 40090
rect -14150 40020 -13850 40090
rect -13650 40020 -13350 40090
rect -13150 40020 -12850 40090
rect -12650 40020 -12350 40090
rect -12150 40020 -11850 40090
rect -11650 40020 -11350 40090
rect -11150 40020 -10850 40090
rect -10650 40020 -10350 40090
rect -10150 40020 -9850 40090
rect -9650 40020 -9350 40090
rect -9150 40020 -8850 40090
rect -8650 40020 -8350 40090
rect -8150 40020 -7850 40090
rect -7650 40020 -7350 40090
rect -7150 40020 -6850 40090
rect -6650 40020 -6350 40090
rect -6150 40020 -5850 40090
rect -5650 40020 -5350 40090
rect -5150 40020 -4850 40090
rect -4650 40020 -4350 40090
rect -4150 40020 -3850 40090
rect -3650 40020 -3350 40090
rect -3150 40020 -2850 40090
rect -2650 40020 -2350 40090
rect -2150 40020 -1850 40090
rect -1650 40020 -1350 40090
rect -1150 40020 -850 40090
rect -650 40020 -350 40090
rect -150 40020 150 40090
rect 350 40020 650 40090
rect 850 40020 1150 40090
rect 1350 40020 1650 40090
rect 1850 40020 2150 40090
rect 2350 40020 2650 40090
rect 2850 40020 3150 40090
rect 3350 40020 3650 40090
rect 3850 40020 4000 40090
rect -16000 40000 4000 40020
rect -28000 39980 4000 40000
rect -28000 39910 -27850 39980
rect -27650 39910 -27350 39980
rect -27150 39910 -26850 39980
rect -26650 39910 -26350 39980
rect -26150 39910 -25850 39980
rect -25650 39910 -25350 39980
rect -25150 39910 -24850 39980
rect -24650 39910 -24350 39980
rect -24150 39910 -23850 39980
rect -23650 39910 -23350 39980
rect -23150 39910 -22850 39980
rect -22650 39910 -22350 39980
rect -22150 39910 -21850 39980
rect -21650 39910 -21350 39980
rect -21150 39910 -20850 39980
rect -20650 39910 -20350 39980
rect -20150 39910 -19850 39980
rect -19650 39910 -19350 39980
rect -19150 39910 -18850 39980
rect -18650 39910 -18350 39980
rect -18150 39910 -17850 39980
rect -17650 39910 -17350 39980
rect -17150 39910 -16850 39980
rect -16650 39910 -16350 39980
rect -16150 39910 -15850 39980
rect -15650 39910 -15350 39980
rect -15150 39910 -14850 39980
rect -14650 39910 -14350 39980
rect -14150 39910 -13850 39980
rect -13650 39910 -13350 39980
rect -13150 39910 -12850 39980
rect -12650 39910 -12350 39980
rect -12150 39910 -11850 39980
rect -11650 39910 -11350 39980
rect -11150 39910 -10850 39980
rect -10650 39910 -10350 39980
rect -10150 39910 -9850 39980
rect -9650 39910 -9350 39980
rect -9150 39910 -8850 39980
rect -8650 39910 -8350 39980
rect -8150 39910 -7850 39980
rect -7650 39910 -7350 39980
rect -7150 39910 -6850 39980
rect -6650 39910 -6350 39980
rect -6150 39910 -5850 39980
rect -5650 39910 -5350 39980
rect -5150 39910 -4850 39980
rect -4650 39910 -4350 39980
rect -4150 39910 -3850 39980
rect -3650 39910 -3350 39980
rect -3150 39910 -2850 39980
rect -2650 39910 -2350 39980
rect -2150 39910 -1850 39980
rect -1650 39910 -1350 39980
rect -1150 39910 -850 39980
rect -650 39910 -350 39980
rect -150 39910 150 39980
rect 350 39910 650 39980
rect 850 39910 1150 39980
rect 1350 39910 1650 39980
rect 1850 39910 2150 39980
rect 2350 39910 2650 39980
rect 2850 39910 3150 39980
rect 3350 39910 3650 39980
rect 3850 39910 4000 39980
rect -28000 39900 4000 39910
rect -28000 39880 -27880 39900
rect -27620 39880 -27380 39900
rect -27120 39880 -26880 39900
rect -26620 39880 -26380 39900
rect -26120 39880 -25880 39900
rect -25620 39880 -25380 39900
rect -25120 39880 -24880 39900
rect -24620 39880 -24380 39900
rect -24120 39880 -23880 39900
rect -23620 39880 -23380 39900
rect -23120 39880 -22880 39900
rect -22620 39880 -22380 39900
rect -22120 39880 -21880 39900
rect -21620 39880 -21380 39900
rect -21120 39880 -20880 39900
rect -20620 39880 -20380 39900
rect -20120 39880 -19880 39900
rect -19620 39880 -19380 39900
rect -19120 39880 -18880 39900
rect -18620 39880 -18380 39900
rect -18120 39880 -17880 39900
rect -17620 39880 -17380 39900
rect -17120 39880 -16880 39900
rect -16620 39880 -16380 39900
rect -16120 39880 -15880 39900
rect -15620 39880 -15380 39900
rect -15120 39880 -14880 39900
rect -14620 39880 -14380 39900
rect -14120 39880 -13880 39900
rect -13620 39880 -13380 39900
rect -13120 39880 -12880 39900
rect -12620 39880 -12380 39900
rect -12120 39880 -11880 39900
rect -11620 39880 -11380 39900
rect -11120 39880 -10880 39900
rect -10620 39880 -10380 39900
rect -10120 39880 -9880 39900
rect -9620 39880 -9380 39900
rect -9120 39880 -8880 39900
rect -8620 39880 -8380 39900
rect -8120 39880 -7880 39900
rect -7620 39880 -7380 39900
rect -7120 39880 -6880 39900
rect -6620 39880 -6380 39900
rect -6120 39880 -5880 39900
rect -5620 39880 -5380 39900
rect -5120 39880 -4880 39900
rect -4620 39880 -4380 39900
rect -4120 39880 -3880 39900
rect -3620 39880 -3380 39900
rect -3120 39880 -2880 39900
rect -2620 39880 -2380 39900
rect -2120 39880 -1880 39900
rect -1620 39880 -1380 39900
rect -1120 39880 -880 39900
rect -620 39880 -380 39900
rect -120 39880 120 39900
rect 380 39880 620 39900
rect 880 39880 1120 39900
rect 1380 39880 1620 39900
rect 1880 39880 2120 39900
rect 2380 39880 2620 39900
rect 2880 39880 3120 39900
rect 3380 39880 3620 39900
rect 3880 39880 4000 39900
rect -28000 39850 -27900 39880
rect -28000 39650 -27980 39850
rect -27910 39650 -27900 39850
rect -28000 39620 -27900 39650
rect -27600 39850 -27400 39880
rect -27600 39650 -27590 39850
rect -27520 39650 -27480 39850
rect -27410 39650 -27400 39850
rect -27600 39620 -27400 39650
rect -27100 39850 -26900 39880
rect -27100 39650 -27090 39850
rect -27020 39650 -26980 39850
rect -26910 39650 -26900 39850
rect -27100 39620 -26900 39650
rect -26600 39850 -26400 39880
rect -26600 39650 -26590 39850
rect -26520 39650 -26480 39850
rect -26410 39650 -26400 39850
rect -26600 39620 -26400 39650
rect -26100 39850 -25900 39880
rect -26100 39650 -26090 39850
rect -26020 39650 -25980 39850
rect -25910 39650 -25900 39850
rect -26100 39620 -25900 39650
rect -25600 39850 -25400 39880
rect -25600 39650 -25590 39850
rect -25520 39650 -25480 39850
rect -25410 39650 -25400 39850
rect -25600 39620 -25400 39650
rect -25100 39850 -24900 39880
rect -25100 39650 -25090 39850
rect -25020 39650 -24980 39850
rect -24910 39650 -24900 39850
rect -25100 39620 -24900 39650
rect -24600 39850 -24400 39880
rect -24600 39650 -24590 39850
rect -24520 39650 -24480 39850
rect -24410 39650 -24400 39850
rect -24600 39620 -24400 39650
rect -24100 39850 -23900 39880
rect -24100 39650 -24090 39850
rect -24020 39650 -23980 39850
rect -23910 39650 -23900 39850
rect -24100 39620 -23900 39650
rect -23600 39850 -23400 39880
rect -23600 39650 -23590 39850
rect -23520 39650 -23480 39850
rect -23410 39650 -23400 39850
rect -23600 39620 -23400 39650
rect -23100 39850 -22900 39880
rect -23100 39650 -23090 39850
rect -23020 39650 -22980 39850
rect -22910 39650 -22900 39850
rect -23100 39620 -22900 39650
rect -22600 39850 -22400 39880
rect -22600 39650 -22590 39850
rect -22520 39650 -22480 39850
rect -22410 39650 -22400 39850
rect -22600 39620 -22400 39650
rect -22100 39850 -21900 39880
rect -22100 39650 -22090 39850
rect -22020 39650 -21980 39850
rect -21910 39650 -21900 39850
rect -22100 39620 -21900 39650
rect -21600 39850 -21400 39880
rect -21600 39650 -21590 39850
rect -21520 39650 -21480 39850
rect -21410 39650 -21400 39850
rect -21600 39620 -21400 39650
rect -21100 39850 -20900 39880
rect -21100 39650 -21090 39850
rect -21020 39650 -20980 39850
rect -20910 39650 -20900 39850
rect -21100 39620 -20900 39650
rect -20600 39850 -20400 39880
rect -20600 39650 -20590 39850
rect -20520 39650 -20480 39850
rect -20410 39650 -20400 39850
rect -20600 39620 -20400 39650
rect -20100 39850 -19900 39880
rect -20100 39650 -20090 39850
rect -20020 39650 -19980 39850
rect -19910 39650 -19900 39850
rect -20100 39620 -19900 39650
rect -19600 39850 -19400 39880
rect -19600 39650 -19590 39850
rect -19520 39650 -19480 39850
rect -19410 39650 -19400 39850
rect -19600 39620 -19400 39650
rect -19100 39850 -18900 39880
rect -19100 39650 -19090 39850
rect -19020 39650 -18980 39850
rect -18910 39650 -18900 39850
rect -19100 39620 -18900 39650
rect -18600 39850 -18400 39880
rect -18600 39650 -18590 39850
rect -18520 39650 -18480 39850
rect -18410 39650 -18400 39850
rect -18600 39620 -18400 39650
rect -18100 39850 -17900 39880
rect -18100 39650 -18090 39850
rect -18020 39650 -17980 39850
rect -17910 39650 -17900 39850
rect -18100 39620 -17900 39650
rect -17600 39850 -17400 39880
rect -17600 39650 -17590 39850
rect -17520 39650 -17480 39850
rect -17410 39650 -17400 39850
rect -17600 39620 -17400 39650
rect -17100 39850 -16900 39880
rect -17100 39650 -17090 39850
rect -17020 39650 -16980 39850
rect -16910 39650 -16900 39850
rect -17100 39620 -16900 39650
rect -16600 39850 -16400 39880
rect -16600 39650 -16590 39850
rect -16520 39650 -16480 39850
rect -16410 39650 -16400 39850
rect -16600 39620 -16400 39650
rect -16100 39850 -15900 39880
rect -16100 39650 -16090 39850
rect -16020 39650 -15980 39850
rect -15910 39650 -15900 39850
rect -16100 39620 -15900 39650
rect -15600 39850 -15400 39880
rect -15600 39650 -15590 39850
rect -15520 39650 -15480 39850
rect -15410 39650 -15400 39850
rect -15600 39620 -15400 39650
rect -15100 39850 -14900 39880
rect -15100 39650 -15090 39850
rect -15020 39650 -14980 39850
rect -14910 39650 -14900 39850
rect -15100 39620 -14900 39650
rect -14600 39850 -14400 39880
rect -14600 39650 -14590 39850
rect -14520 39650 -14480 39850
rect -14410 39650 -14400 39850
rect -14600 39620 -14400 39650
rect -14100 39850 -13900 39880
rect -14100 39650 -14090 39850
rect -14020 39650 -13980 39850
rect -13910 39650 -13900 39850
rect -14100 39620 -13900 39650
rect -13600 39850 -13400 39880
rect -13600 39650 -13590 39850
rect -13520 39650 -13480 39850
rect -13410 39650 -13400 39850
rect -13600 39620 -13400 39650
rect -13100 39850 -12900 39880
rect -13100 39650 -13090 39850
rect -13020 39650 -12980 39850
rect -12910 39650 -12900 39850
rect -13100 39620 -12900 39650
rect -12600 39850 -12400 39880
rect -12600 39650 -12590 39850
rect -12520 39650 -12480 39850
rect -12410 39650 -12400 39850
rect -12600 39620 -12400 39650
rect -12100 39850 -11900 39880
rect -12100 39650 -12090 39850
rect -12020 39650 -11980 39850
rect -11910 39650 -11900 39850
rect -12100 39620 -11900 39650
rect -11600 39850 -11400 39880
rect -11600 39650 -11590 39850
rect -11520 39650 -11480 39850
rect -11410 39650 -11400 39850
rect -11600 39620 -11400 39650
rect -11100 39850 -10900 39880
rect -11100 39650 -11090 39850
rect -11020 39650 -10980 39850
rect -10910 39650 -10900 39850
rect -11100 39620 -10900 39650
rect -10600 39850 -10400 39880
rect -10600 39650 -10590 39850
rect -10520 39650 -10480 39850
rect -10410 39650 -10400 39850
rect -10600 39620 -10400 39650
rect -10100 39850 -9900 39880
rect -10100 39650 -10090 39850
rect -10020 39650 -9980 39850
rect -9910 39650 -9900 39850
rect -10100 39620 -9900 39650
rect -9600 39850 -9400 39880
rect -9600 39650 -9590 39850
rect -9520 39650 -9480 39850
rect -9410 39650 -9400 39850
rect -9600 39620 -9400 39650
rect -9100 39850 -8900 39880
rect -9100 39650 -9090 39850
rect -9020 39650 -8980 39850
rect -8910 39650 -8900 39850
rect -9100 39620 -8900 39650
rect -8600 39850 -8400 39880
rect -8600 39650 -8590 39850
rect -8520 39650 -8480 39850
rect -8410 39650 -8400 39850
rect -8600 39620 -8400 39650
rect -8100 39850 -7900 39880
rect -8100 39650 -8090 39850
rect -8020 39650 -7980 39850
rect -7910 39650 -7900 39850
rect -8100 39620 -7900 39650
rect -7600 39850 -7400 39880
rect -7600 39650 -7590 39850
rect -7520 39650 -7480 39850
rect -7410 39650 -7400 39850
rect -7600 39620 -7400 39650
rect -7100 39850 -6900 39880
rect -7100 39650 -7090 39850
rect -7020 39650 -6980 39850
rect -6910 39650 -6900 39850
rect -7100 39620 -6900 39650
rect -6600 39850 -6400 39880
rect -6600 39650 -6590 39850
rect -6520 39650 -6480 39850
rect -6410 39650 -6400 39850
rect -6600 39620 -6400 39650
rect -6100 39850 -5900 39880
rect -6100 39650 -6090 39850
rect -6020 39650 -5980 39850
rect -5910 39650 -5900 39850
rect -6100 39620 -5900 39650
rect -5600 39850 -5400 39880
rect -5600 39650 -5590 39850
rect -5520 39650 -5480 39850
rect -5410 39650 -5400 39850
rect -5600 39620 -5400 39650
rect -5100 39850 -4900 39880
rect -5100 39650 -5090 39850
rect -5020 39650 -4980 39850
rect -4910 39650 -4900 39850
rect -5100 39620 -4900 39650
rect -4600 39850 -4400 39880
rect -4600 39650 -4590 39850
rect -4520 39650 -4480 39850
rect -4410 39650 -4400 39850
rect -4600 39620 -4400 39650
rect -4100 39850 -3900 39880
rect -4100 39650 -4090 39850
rect -4020 39650 -3980 39850
rect -3910 39650 -3900 39850
rect -4100 39620 -3900 39650
rect -3600 39850 -3400 39880
rect -3600 39650 -3590 39850
rect -3520 39650 -3480 39850
rect -3410 39650 -3400 39850
rect -3600 39620 -3400 39650
rect -3100 39850 -2900 39880
rect -3100 39650 -3090 39850
rect -3020 39650 -2980 39850
rect -2910 39650 -2900 39850
rect -3100 39620 -2900 39650
rect -2600 39850 -2400 39880
rect -2600 39650 -2590 39850
rect -2520 39650 -2480 39850
rect -2410 39650 -2400 39850
rect -2600 39620 -2400 39650
rect -2100 39850 -1900 39880
rect -2100 39650 -2090 39850
rect -2020 39650 -1980 39850
rect -1910 39650 -1900 39850
rect -2100 39620 -1900 39650
rect -1600 39850 -1400 39880
rect -1600 39650 -1590 39850
rect -1520 39650 -1480 39850
rect -1410 39650 -1400 39850
rect -1600 39620 -1400 39650
rect -1100 39850 -900 39880
rect -1100 39650 -1090 39850
rect -1020 39650 -980 39850
rect -910 39650 -900 39850
rect -1100 39620 -900 39650
rect -600 39850 -400 39880
rect -600 39650 -590 39850
rect -520 39650 -480 39850
rect -410 39650 -400 39850
rect -600 39620 -400 39650
rect -100 39850 100 39880
rect -100 39650 -90 39850
rect -20 39650 20 39850
rect 90 39650 100 39850
rect -100 39620 100 39650
rect 400 39850 600 39880
rect 400 39650 410 39850
rect 480 39650 520 39850
rect 590 39650 600 39850
rect 400 39620 600 39650
rect 900 39850 1100 39880
rect 900 39650 910 39850
rect 980 39650 1020 39850
rect 1090 39650 1100 39850
rect 900 39620 1100 39650
rect 1400 39850 1600 39880
rect 1400 39650 1410 39850
rect 1480 39650 1520 39850
rect 1590 39650 1600 39850
rect 1400 39620 1600 39650
rect 1900 39850 2100 39880
rect 1900 39650 1910 39850
rect 1980 39650 2020 39850
rect 2090 39650 2100 39850
rect 1900 39620 2100 39650
rect 2400 39850 2600 39880
rect 2400 39650 2410 39850
rect 2480 39650 2520 39850
rect 2590 39650 2600 39850
rect 2400 39620 2600 39650
rect 2900 39850 3100 39880
rect 2900 39650 2910 39850
rect 2980 39650 3020 39850
rect 3090 39650 3100 39850
rect 2900 39620 3100 39650
rect 3400 39850 3600 39880
rect 3400 39650 3410 39850
rect 3480 39650 3520 39850
rect 3590 39650 3600 39850
rect 3400 39620 3600 39650
rect 3900 39850 4000 39880
rect 3900 39650 3910 39850
rect 3980 39650 4000 39850
rect 3900 39620 4000 39650
rect -28000 39600 -27880 39620
rect -27620 39600 -27380 39620
rect -27120 39600 -26880 39620
rect -26620 39600 -26380 39620
rect -26120 39600 -25880 39620
rect -25620 39600 -25380 39620
rect -25120 39600 -24880 39620
rect -24620 39600 -24380 39620
rect -24120 39600 -23880 39620
rect -23620 39600 -23380 39620
rect -23120 39600 -22880 39620
rect -22620 39600 -22380 39620
rect -22120 39600 -21880 39620
rect -21620 39600 -21380 39620
rect -21120 39600 -20880 39620
rect -20620 39600 -20380 39620
rect -20120 39600 -19880 39620
rect -19620 39600 -19380 39620
rect -19120 39600 -18880 39620
rect -18620 39600 -18380 39620
rect -18120 39600 -17880 39620
rect -17620 39600 -17380 39620
rect -17120 39600 -16880 39620
rect -16620 39600 -16380 39620
rect -16120 39600 -15880 39620
rect -15620 39600 -15380 39620
rect -15120 39600 -14880 39620
rect -14620 39600 -14380 39620
rect -14120 39600 -13880 39620
rect -13620 39600 -13380 39620
rect -13120 39600 -12880 39620
rect -12620 39600 -12380 39620
rect -12120 39600 -11880 39620
rect -11620 39600 -11380 39620
rect -11120 39600 -10880 39620
rect -10620 39600 -10380 39620
rect -10120 39600 -9880 39620
rect -9620 39600 -9380 39620
rect -9120 39600 -8880 39620
rect -8620 39600 -8380 39620
rect -8120 39600 -7880 39620
rect -7620 39600 -7380 39620
rect -7120 39600 -6880 39620
rect -6620 39600 -6380 39620
rect -6120 39600 -5880 39620
rect -5620 39600 -5380 39620
rect -5120 39600 -4880 39620
rect -4620 39600 -4380 39620
rect -4120 39600 -3880 39620
rect -3620 39600 -3380 39620
rect -3120 39600 -2880 39620
rect -2620 39600 -2380 39620
rect -2120 39600 -1880 39620
rect -1620 39600 -1380 39620
rect -1120 39600 -880 39620
rect -620 39600 -380 39620
rect -120 39600 120 39620
rect 380 39600 620 39620
rect 880 39600 1120 39620
rect 1380 39600 1620 39620
rect 1880 39600 2120 39620
rect 2380 39600 2620 39620
rect 2880 39600 3120 39620
rect 3380 39600 3620 39620
rect 3880 39600 4000 39620
rect -28000 39590 4000 39600
rect -28000 39520 -27850 39590
rect -27650 39520 -27350 39590
rect -27150 39520 -26850 39590
rect -26650 39520 -26350 39590
rect -26150 39520 -25850 39590
rect -25650 39520 -25350 39590
rect -25150 39520 -24850 39590
rect -24650 39520 -24350 39590
rect -24150 39520 -23850 39590
rect -23650 39520 -23350 39590
rect -23150 39520 -22850 39590
rect -22650 39520 -22350 39590
rect -22150 39520 -21850 39590
rect -21650 39520 -21350 39590
rect -21150 39520 -20850 39590
rect -20650 39520 -20350 39590
rect -20150 39520 -19850 39590
rect -19650 39520 -19350 39590
rect -19150 39520 -18850 39590
rect -18650 39520 -18350 39590
rect -18150 39520 -17850 39590
rect -17650 39520 -17350 39590
rect -17150 39520 -16850 39590
rect -16650 39520 -16350 39590
rect -16150 39520 -15850 39590
rect -15650 39520 -15350 39590
rect -15150 39520 -14850 39590
rect -14650 39520 -14350 39590
rect -14150 39520 -13850 39590
rect -13650 39520 -13350 39590
rect -13150 39520 -12850 39590
rect -12650 39520 -12350 39590
rect -12150 39520 -11850 39590
rect -11650 39520 -11350 39590
rect -11150 39520 -10850 39590
rect -10650 39520 -10350 39590
rect -10150 39520 -9850 39590
rect -9650 39520 -9350 39590
rect -9150 39520 -8850 39590
rect -8650 39520 -8350 39590
rect -8150 39520 -7850 39590
rect -7650 39520 -7350 39590
rect -7150 39520 -6850 39590
rect -6650 39520 -6350 39590
rect -6150 39520 -5850 39590
rect -5650 39520 -5350 39590
rect -5150 39520 -4850 39590
rect -4650 39520 -4350 39590
rect -4150 39520 -3850 39590
rect -3650 39520 -3350 39590
rect -3150 39520 -2850 39590
rect -2650 39520 -2350 39590
rect -2150 39520 -1850 39590
rect -1650 39520 -1350 39590
rect -1150 39520 -850 39590
rect -650 39520 -350 39590
rect -150 39520 150 39590
rect 350 39520 650 39590
rect 850 39520 1150 39590
rect 1350 39520 1650 39590
rect 1850 39520 2150 39590
rect 2350 39520 2650 39590
rect 2850 39520 3150 39590
rect 3350 39520 3650 39590
rect 3850 39520 4000 39590
rect -28000 39480 4000 39520
rect -28000 39410 -27850 39480
rect -27650 39410 -27350 39480
rect -27150 39410 -26850 39480
rect -26650 39410 -26350 39480
rect -26150 39410 -25850 39480
rect -25650 39410 -25350 39480
rect -25150 39410 -24850 39480
rect -24650 39410 -24350 39480
rect -24150 39410 -23850 39480
rect -23650 39410 -23350 39480
rect -23150 39410 -22850 39480
rect -22650 39410 -22350 39480
rect -22150 39410 -21850 39480
rect -21650 39410 -21350 39480
rect -21150 39410 -20850 39480
rect -20650 39410 -20350 39480
rect -20150 39410 -19850 39480
rect -19650 39410 -19350 39480
rect -19150 39410 -18850 39480
rect -18650 39410 -18350 39480
rect -18150 39410 -17850 39480
rect -17650 39410 -17350 39480
rect -17150 39410 -16850 39480
rect -16650 39410 -16350 39480
rect -16150 39410 -15850 39480
rect -15650 39410 -15350 39480
rect -15150 39410 -14850 39480
rect -14650 39410 -14350 39480
rect -14150 39410 -13850 39480
rect -13650 39410 -13350 39480
rect -13150 39410 -12850 39480
rect -12650 39410 -12350 39480
rect -12150 39410 -11850 39480
rect -11650 39410 -11350 39480
rect -11150 39410 -10850 39480
rect -10650 39410 -10350 39480
rect -10150 39410 -9850 39480
rect -9650 39410 -9350 39480
rect -9150 39410 -8850 39480
rect -8650 39410 -8350 39480
rect -8150 39410 -7850 39480
rect -7650 39410 -7350 39480
rect -7150 39410 -6850 39480
rect -6650 39410 -6350 39480
rect -6150 39410 -5850 39480
rect -5650 39410 -5350 39480
rect -5150 39410 -4850 39480
rect -4650 39410 -4350 39480
rect -4150 39410 -3850 39480
rect -3650 39410 -3350 39480
rect -3150 39410 -2850 39480
rect -2650 39410 -2350 39480
rect -2150 39410 -1850 39480
rect -1650 39410 -1350 39480
rect -1150 39410 -850 39480
rect -650 39410 -350 39480
rect -150 39410 150 39480
rect 350 39410 650 39480
rect 850 39410 1150 39480
rect 1350 39410 1650 39480
rect 1850 39410 2150 39480
rect 2350 39410 2650 39480
rect 2850 39410 3150 39480
rect 3350 39410 3650 39480
rect 3850 39410 4000 39480
rect -28000 39400 4000 39410
rect -28000 39380 -27880 39400
rect -27620 39380 -27380 39400
rect -27120 39380 -26880 39400
rect -26620 39380 -26380 39400
rect -26120 39380 -25880 39400
rect -25620 39380 -25380 39400
rect -25120 39380 -24880 39400
rect -24620 39380 -24380 39400
rect -24120 39380 -23880 39400
rect -23620 39380 -23380 39400
rect -23120 39380 -22880 39400
rect -22620 39380 -22380 39400
rect -22120 39380 -21880 39400
rect -21620 39380 -21380 39400
rect -21120 39380 -20880 39400
rect -20620 39380 -20380 39400
rect -20120 39380 -19880 39400
rect -19620 39380 -19380 39400
rect -19120 39380 -18880 39400
rect -18620 39380 -18380 39400
rect -18120 39380 -17880 39400
rect -17620 39380 -17380 39400
rect -17120 39380 -16880 39400
rect -16620 39380 -16380 39400
rect -16120 39380 -15880 39400
rect -15620 39380 -15380 39400
rect -15120 39380 -14880 39400
rect -14620 39380 -14380 39400
rect -14120 39380 -13880 39400
rect -13620 39380 -13380 39400
rect -13120 39380 -12880 39400
rect -12620 39380 -12380 39400
rect -12120 39380 -11880 39400
rect -11620 39380 -11380 39400
rect -11120 39380 -10880 39400
rect -10620 39380 -10380 39400
rect -10120 39380 -9880 39400
rect -9620 39380 -9380 39400
rect -9120 39380 -8880 39400
rect -8620 39380 -8380 39400
rect -8120 39380 -7880 39400
rect -7620 39380 -7380 39400
rect -7120 39380 -6880 39400
rect -6620 39380 -6380 39400
rect -6120 39380 -5880 39400
rect -5620 39380 -5380 39400
rect -5120 39380 -4880 39400
rect -4620 39380 -4380 39400
rect -4120 39380 -3880 39400
rect -3620 39380 -3380 39400
rect -3120 39380 -2880 39400
rect -2620 39380 -2380 39400
rect -2120 39380 -1880 39400
rect -1620 39380 -1380 39400
rect -1120 39380 -880 39400
rect -620 39380 -380 39400
rect -120 39380 120 39400
rect 380 39380 620 39400
rect 880 39380 1120 39400
rect 1380 39380 1620 39400
rect 1880 39380 2120 39400
rect 2380 39380 2620 39400
rect 2880 39380 3120 39400
rect 3380 39380 3620 39400
rect 3880 39380 4000 39400
rect -28000 39350 -27900 39380
rect -28000 39150 -27980 39350
rect -27910 39150 -27900 39350
rect -28000 39120 -27900 39150
rect -27600 39350 -27400 39380
rect -27600 39150 -27590 39350
rect -27520 39150 -27480 39350
rect -27410 39150 -27400 39350
rect -27600 39120 -27400 39150
rect -27100 39350 -26900 39380
rect -27100 39150 -27090 39350
rect -27020 39150 -26980 39350
rect -26910 39150 -26900 39350
rect -27100 39120 -26900 39150
rect -26600 39350 -26400 39380
rect -26600 39150 -26590 39350
rect -26520 39150 -26480 39350
rect -26410 39150 -26400 39350
rect -26600 39120 -26400 39150
rect -26100 39350 -25900 39380
rect -26100 39150 -26090 39350
rect -26020 39150 -25980 39350
rect -25910 39150 -25900 39350
rect -26100 39120 -25900 39150
rect -25600 39350 -25400 39380
rect -25600 39150 -25590 39350
rect -25520 39150 -25480 39350
rect -25410 39150 -25400 39350
rect -25600 39120 -25400 39150
rect -25100 39350 -24900 39380
rect -25100 39150 -25090 39350
rect -25020 39150 -24980 39350
rect -24910 39150 -24900 39350
rect -25100 39120 -24900 39150
rect -24600 39350 -24400 39380
rect -24600 39150 -24590 39350
rect -24520 39150 -24480 39350
rect -24410 39150 -24400 39350
rect -24600 39120 -24400 39150
rect -24100 39350 -23900 39380
rect -24100 39150 -24090 39350
rect -24020 39150 -23980 39350
rect -23910 39150 -23900 39350
rect -24100 39120 -23900 39150
rect -23600 39350 -23400 39380
rect -23600 39150 -23590 39350
rect -23520 39150 -23480 39350
rect -23410 39150 -23400 39350
rect -23600 39120 -23400 39150
rect -23100 39350 -22900 39380
rect -23100 39150 -23090 39350
rect -23020 39150 -22980 39350
rect -22910 39150 -22900 39350
rect -23100 39120 -22900 39150
rect -22600 39350 -22400 39380
rect -22600 39150 -22590 39350
rect -22520 39150 -22480 39350
rect -22410 39150 -22400 39350
rect -22600 39120 -22400 39150
rect -22100 39350 -21900 39380
rect -22100 39150 -22090 39350
rect -22020 39150 -21980 39350
rect -21910 39150 -21900 39350
rect -22100 39120 -21900 39150
rect -21600 39350 -21400 39380
rect -21600 39150 -21590 39350
rect -21520 39150 -21480 39350
rect -21410 39150 -21400 39350
rect -21600 39120 -21400 39150
rect -21100 39350 -20900 39380
rect -21100 39150 -21090 39350
rect -21020 39150 -20980 39350
rect -20910 39150 -20900 39350
rect -21100 39120 -20900 39150
rect -20600 39350 -20400 39380
rect -20600 39150 -20590 39350
rect -20520 39150 -20480 39350
rect -20410 39150 -20400 39350
rect -20600 39120 -20400 39150
rect -20100 39350 -19900 39380
rect -20100 39150 -20090 39350
rect -20020 39150 -19980 39350
rect -19910 39150 -19900 39350
rect -20100 39120 -19900 39150
rect -19600 39350 -19400 39380
rect -19600 39150 -19590 39350
rect -19520 39150 -19480 39350
rect -19410 39150 -19400 39350
rect -19600 39120 -19400 39150
rect -19100 39350 -18900 39380
rect -19100 39150 -19090 39350
rect -19020 39150 -18980 39350
rect -18910 39150 -18900 39350
rect -19100 39120 -18900 39150
rect -18600 39350 -18400 39380
rect -18600 39150 -18590 39350
rect -18520 39150 -18480 39350
rect -18410 39150 -18400 39350
rect -18600 39120 -18400 39150
rect -18100 39350 -17900 39380
rect -18100 39150 -18090 39350
rect -18020 39150 -17980 39350
rect -17910 39150 -17900 39350
rect -18100 39120 -17900 39150
rect -17600 39350 -17400 39380
rect -17600 39150 -17590 39350
rect -17520 39150 -17480 39350
rect -17410 39150 -17400 39350
rect -17600 39120 -17400 39150
rect -17100 39350 -16900 39380
rect -17100 39150 -17090 39350
rect -17020 39150 -16980 39350
rect -16910 39150 -16900 39350
rect -17100 39120 -16900 39150
rect -16600 39350 -16400 39380
rect -16600 39150 -16590 39350
rect -16520 39150 -16480 39350
rect -16410 39150 -16400 39350
rect -16600 39120 -16400 39150
rect -16100 39350 -15900 39380
rect -16100 39150 -16090 39350
rect -16020 39150 -15980 39350
rect -15910 39150 -15900 39350
rect -16100 39120 -15900 39150
rect -15600 39350 -15400 39380
rect -15600 39150 -15590 39350
rect -15520 39150 -15480 39350
rect -15410 39150 -15400 39350
rect -15600 39120 -15400 39150
rect -15100 39350 -14900 39380
rect -15100 39150 -15090 39350
rect -15020 39150 -14980 39350
rect -14910 39150 -14900 39350
rect -15100 39120 -14900 39150
rect -14600 39350 -14400 39380
rect -14600 39150 -14590 39350
rect -14520 39150 -14480 39350
rect -14410 39150 -14400 39350
rect -14600 39120 -14400 39150
rect -14100 39350 -13900 39380
rect -14100 39150 -14090 39350
rect -14020 39150 -13980 39350
rect -13910 39150 -13900 39350
rect -14100 39120 -13900 39150
rect -13600 39350 -13400 39380
rect -13600 39150 -13590 39350
rect -13520 39150 -13480 39350
rect -13410 39150 -13400 39350
rect -13600 39120 -13400 39150
rect -13100 39350 -12900 39380
rect -13100 39150 -13090 39350
rect -13020 39150 -12980 39350
rect -12910 39150 -12900 39350
rect -13100 39120 -12900 39150
rect -12600 39350 -12400 39380
rect -12600 39150 -12590 39350
rect -12520 39150 -12480 39350
rect -12410 39150 -12400 39350
rect -12600 39120 -12400 39150
rect -12100 39350 -11900 39380
rect -12100 39150 -12090 39350
rect -12020 39150 -11980 39350
rect -11910 39150 -11900 39350
rect -12100 39120 -11900 39150
rect -11600 39350 -11400 39380
rect -11600 39150 -11590 39350
rect -11520 39150 -11480 39350
rect -11410 39150 -11400 39350
rect -11600 39120 -11400 39150
rect -11100 39350 -10900 39380
rect -11100 39150 -11090 39350
rect -11020 39150 -10980 39350
rect -10910 39150 -10900 39350
rect -11100 39120 -10900 39150
rect -10600 39350 -10400 39380
rect -10600 39150 -10590 39350
rect -10520 39150 -10480 39350
rect -10410 39150 -10400 39350
rect -10600 39120 -10400 39150
rect -10100 39350 -9900 39380
rect -10100 39150 -10090 39350
rect -10020 39150 -9980 39350
rect -9910 39150 -9900 39350
rect -10100 39120 -9900 39150
rect -9600 39350 -9400 39380
rect -9600 39150 -9590 39350
rect -9520 39150 -9480 39350
rect -9410 39150 -9400 39350
rect -9600 39120 -9400 39150
rect -9100 39350 -8900 39380
rect -9100 39150 -9090 39350
rect -9020 39150 -8980 39350
rect -8910 39150 -8900 39350
rect -9100 39120 -8900 39150
rect -8600 39350 -8400 39380
rect -8600 39150 -8590 39350
rect -8520 39150 -8480 39350
rect -8410 39150 -8400 39350
rect -8600 39120 -8400 39150
rect -8100 39350 -7900 39380
rect -8100 39150 -8090 39350
rect -8020 39150 -7980 39350
rect -7910 39150 -7900 39350
rect -8100 39120 -7900 39150
rect -7600 39350 -7400 39380
rect -7600 39150 -7590 39350
rect -7520 39150 -7480 39350
rect -7410 39150 -7400 39350
rect -7600 39120 -7400 39150
rect -7100 39350 -6900 39380
rect -7100 39150 -7090 39350
rect -7020 39150 -6980 39350
rect -6910 39150 -6900 39350
rect -7100 39120 -6900 39150
rect -6600 39350 -6400 39380
rect -6600 39150 -6590 39350
rect -6520 39150 -6480 39350
rect -6410 39150 -6400 39350
rect -6600 39120 -6400 39150
rect -6100 39350 -5900 39380
rect -6100 39150 -6090 39350
rect -6020 39150 -5980 39350
rect -5910 39150 -5900 39350
rect -6100 39120 -5900 39150
rect -5600 39350 -5400 39380
rect -5600 39150 -5590 39350
rect -5520 39150 -5480 39350
rect -5410 39150 -5400 39350
rect -5600 39120 -5400 39150
rect -5100 39350 -4900 39380
rect -5100 39150 -5090 39350
rect -5020 39150 -4980 39350
rect -4910 39150 -4900 39350
rect -5100 39120 -4900 39150
rect -4600 39350 -4400 39380
rect -4600 39150 -4590 39350
rect -4520 39150 -4480 39350
rect -4410 39150 -4400 39350
rect -4600 39120 -4400 39150
rect -4100 39350 -3900 39380
rect -4100 39150 -4090 39350
rect -4020 39150 -3980 39350
rect -3910 39150 -3900 39350
rect -4100 39120 -3900 39150
rect -3600 39350 -3400 39380
rect -3600 39150 -3590 39350
rect -3520 39150 -3480 39350
rect -3410 39150 -3400 39350
rect -3600 39120 -3400 39150
rect -3100 39350 -2900 39380
rect -3100 39150 -3090 39350
rect -3020 39150 -2980 39350
rect -2910 39150 -2900 39350
rect -3100 39120 -2900 39150
rect -2600 39350 -2400 39380
rect -2600 39150 -2590 39350
rect -2520 39150 -2480 39350
rect -2410 39150 -2400 39350
rect -2600 39120 -2400 39150
rect -2100 39350 -1900 39380
rect -2100 39150 -2090 39350
rect -2020 39150 -1980 39350
rect -1910 39150 -1900 39350
rect -2100 39120 -1900 39150
rect -1600 39350 -1400 39380
rect -1600 39150 -1590 39350
rect -1520 39150 -1480 39350
rect -1410 39150 -1400 39350
rect -1600 39120 -1400 39150
rect -1100 39350 -900 39380
rect -1100 39150 -1090 39350
rect -1020 39150 -980 39350
rect -910 39150 -900 39350
rect -1100 39120 -900 39150
rect -600 39350 -400 39380
rect -600 39150 -590 39350
rect -520 39150 -480 39350
rect -410 39150 -400 39350
rect -600 39120 -400 39150
rect -100 39350 100 39380
rect -100 39150 -90 39350
rect -20 39150 20 39350
rect 90 39150 100 39350
rect -100 39120 100 39150
rect 400 39350 600 39380
rect 400 39150 410 39350
rect 480 39150 520 39350
rect 590 39150 600 39350
rect 400 39120 600 39150
rect 900 39350 1100 39380
rect 900 39150 910 39350
rect 980 39150 1020 39350
rect 1090 39150 1100 39350
rect 900 39120 1100 39150
rect 1400 39350 1600 39380
rect 1400 39150 1410 39350
rect 1480 39150 1520 39350
rect 1590 39150 1600 39350
rect 1400 39120 1600 39150
rect 1900 39350 2100 39380
rect 1900 39150 1910 39350
rect 1980 39150 2020 39350
rect 2090 39150 2100 39350
rect 1900 39120 2100 39150
rect 2400 39350 2600 39380
rect 2400 39150 2410 39350
rect 2480 39150 2520 39350
rect 2590 39150 2600 39350
rect 2400 39120 2600 39150
rect 2900 39350 3100 39380
rect 2900 39150 2910 39350
rect 2980 39150 3020 39350
rect 3090 39150 3100 39350
rect 2900 39120 3100 39150
rect 3400 39350 3600 39380
rect 3400 39150 3410 39350
rect 3480 39150 3520 39350
rect 3590 39150 3600 39350
rect 3400 39120 3600 39150
rect 3900 39350 4000 39380
rect 3900 39150 3910 39350
rect 3980 39150 4000 39350
rect 3900 39120 4000 39150
rect -28000 39100 -27880 39120
rect -27620 39100 -27380 39120
rect -27120 39100 -26880 39120
rect -26620 39100 -26380 39120
rect -26120 39100 -25880 39120
rect -25620 39100 -25380 39120
rect -25120 39100 -24880 39120
rect -24620 39100 -24380 39120
rect -24120 39100 -23880 39120
rect -23620 39100 -23380 39120
rect -23120 39100 -22880 39120
rect -22620 39100 -22380 39120
rect -22120 39100 -21880 39120
rect -21620 39100 -21380 39120
rect -21120 39100 -20880 39120
rect -20620 39100 -20380 39120
rect -20120 39100 -19880 39120
rect -19620 39100 -19380 39120
rect -19120 39100 -18880 39120
rect -18620 39100 -18380 39120
rect -18120 39100 -17880 39120
rect -17620 39100 -17380 39120
rect -17120 39100 -16880 39120
rect -16620 39100 -16380 39120
rect -16120 39100 -15880 39120
rect -15620 39100 -15380 39120
rect -15120 39100 -14880 39120
rect -14620 39100 -14380 39120
rect -14120 39100 -13880 39120
rect -13620 39100 -13380 39120
rect -13120 39100 -12880 39120
rect -12620 39100 -12380 39120
rect -12120 39100 -11880 39120
rect -11620 39100 -11380 39120
rect -11120 39100 -10880 39120
rect -10620 39100 -10380 39120
rect -10120 39100 -9880 39120
rect -9620 39100 -9380 39120
rect -9120 39100 -8880 39120
rect -8620 39100 -8380 39120
rect -8120 39100 -7880 39120
rect -7620 39100 -7380 39120
rect -7120 39100 -6880 39120
rect -6620 39100 -6380 39120
rect -6120 39100 -5880 39120
rect -5620 39100 -5380 39120
rect -5120 39100 -4880 39120
rect -4620 39100 -4380 39120
rect -4120 39100 -3880 39120
rect -3620 39100 -3380 39120
rect -3120 39100 -2880 39120
rect -2620 39100 -2380 39120
rect -2120 39100 -1880 39120
rect -1620 39100 -1380 39120
rect -1120 39100 -880 39120
rect -620 39100 -380 39120
rect -120 39100 120 39120
rect 380 39100 620 39120
rect 880 39100 1120 39120
rect 1380 39100 1620 39120
rect 1880 39100 2120 39120
rect 2380 39100 2620 39120
rect 2880 39100 3120 39120
rect 3380 39100 3620 39120
rect 3880 39100 4000 39120
rect -28000 39090 4000 39100
rect -28000 39020 -27850 39090
rect -27650 39020 -27350 39090
rect -27150 39020 -26850 39090
rect -26650 39020 -26350 39090
rect -26150 39020 -25850 39090
rect -25650 39020 -25350 39090
rect -25150 39020 -24850 39090
rect -24650 39020 -24350 39090
rect -24150 39020 -23850 39090
rect -23650 39020 -23350 39090
rect -23150 39020 -22850 39090
rect -22650 39020 -22350 39090
rect -22150 39020 -21850 39090
rect -21650 39020 -21350 39090
rect -21150 39020 -20850 39090
rect -20650 39020 -20350 39090
rect -20150 39020 -19850 39090
rect -19650 39020 -19350 39090
rect -19150 39020 -18850 39090
rect -18650 39020 -18350 39090
rect -18150 39020 -17850 39090
rect -17650 39020 -17350 39090
rect -17150 39020 -16850 39090
rect -16650 39020 -16350 39090
rect -16150 39020 -15850 39090
rect -15650 39020 -15350 39090
rect -15150 39020 -14850 39090
rect -14650 39020 -14350 39090
rect -14150 39020 -13850 39090
rect -13650 39020 -13350 39090
rect -13150 39020 -12850 39090
rect -12650 39020 -12350 39090
rect -12150 39020 -11850 39090
rect -11650 39020 -11350 39090
rect -11150 39020 -10850 39090
rect -10650 39020 -10350 39090
rect -10150 39020 -9850 39090
rect -9650 39020 -9350 39090
rect -9150 39020 -8850 39090
rect -8650 39020 -8350 39090
rect -8150 39020 -7850 39090
rect -7650 39020 -7350 39090
rect -7150 39020 -6850 39090
rect -6650 39020 -6350 39090
rect -6150 39020 -5850 39090
rect -5650 39020 -5350 39090
rect -5150 39020 -4850 39090
rect -4650 39020 -4350 39090
rect -4150 39020 -3850 39090
rect -3650 39020 -3350 39090
rect -3150 39020 -2850 39090
rect -2650 39020 -2350 39090
rect -2150 39020 -1850 39090
rect -1650 39020 -1350 39090
rect -1150 39020 -850 39090
rect -650 39020 -350 39090
rect -150 39020 150 39090
rect 350 39020 650 39090
rect 850 39020 1150 39090
rect 1350 39020 1650 39090
rect 1850 39020 2150 39090
rect 2350 39020 2650 39090
rect 2850 39020 3150 39090
rect 3350 39020 3650 39090
rect 3850 39020 4000 39090
rect -28000 38980 4000 39020
rect -28000 38910 -27850 38980
rect -27650 38910 -27350 38980
rect -27150 38910 -26850 38980
rect -26650 38910 -26350 38980
rect -26150 38910 -25850 38980
rect -25650 38910 -25350 38980
rect -25150 38910 -24850 38980
rect -24650 38910 -24350 38980
rect -24150 38910 -23850 38980
rect -23650 38910 -23350 38980
rect -23150 38910 -22850 38980
rect -22650 38910 -22350 38980
rect -22150 38910 -21850 38980
rect -21650 38910 -21350 38980
rect -21150 38910 -20850 38980
rect -20650 38910 -20350 38980
rect -20150 38910 -19850 38980
rect -19650 38910 -19350 38980
rect -19150 38910 -18850 38980
rect -18650 38910 -18350 38980
rect -18150 38910 -17850 38980
rect -17650 38910 -17350 38980
rect -17150 38910 -16850 38980
rect -16650 38910 -16350 38980
rect -16150 38910 -15850 38980
rect -15650 38910 -15350 38980
rect -15150 38910 -14850 38980
rect -14650 38910 -14350 38980
rect -14150 38910 -13850 38980
rect -13650 38910 -13350 38980
rect -13150 38910 -12850 38980
rect -12650 38910 -12350 38980
rect -12150 38910 -11850 38980
rect -11650 38910 -11350 38980
rect -11150 38910 -10850 38980
rect -10650 38910 -10350 38980
rect -10150 38910 -9850 38980
rect -9650 38910 -9350 38980
rect -9150 38910 -8850 38980
rect -8650 38910 -8350 38980
rect -8150 38910 -7850 38980
rect -7650 38910 -7350 38980
rect -7150 38910 -6850 38980
rect -6650 38910 -6350 38980
rect -6150 38910 -5850 38980
rect -5650 38910 -5350 38980
rect -5150 38910 -4850 38980
rect -4650 38910 -4350 38980
rect -4150 38910 -3850 38980
rect -3650 38910 -3350 38980
rect -3150 38910 -2850 38980
rect -2650 38910 -2350 38980
rect -2150 38910 -1850 38980
rect -1650 38910 -1350 38980
rect -1150 38910 -850 38980
rect -650 38910 -350 38980
rect -150 38910 150 38980
rect 350 38910 650 38980
rect 850 38910 1150 38980
rect 1350 38910 1650 38980
rect 1850 38910 2150 38980
rect 2350 38910 2650 38980
rect 2850 38910 3150 38980
rect 3350 38910 3650 38980
rect 3850 38910 4000 38980
rect -28000 38900 4000 38910
rect -28000 38880 -27880 38900
rect -27620 38880 -27380 38900
rect -27120 38880 -26880 38900
rect -26620 38880 -26380 38900
rect -26120 38880 -25880 38900
rect -25620 38880 -25380 38900
rect -25120 38880 -24880 38900
rect -24620 38880 -24380 38900
rect -24120 38880 -23880 38900
rect -23620 38880 -23380 38900
rect -23120 38880 -22880 38900
rect -22620 38880 -22380 38900
rect -22120 38880 -21880 38900
rect -21620 38880 -21380 38900
rect -21120 38880 -20880 38900
rect -20620 38880 -20380 38900
rect -20120 38880 -19880 38900
rect -19620 38880 -19380 38900
rect -19120 38880 -18880 38900
rect -18620 38880 -18380 38900
rect -18120 38880 -17880 38900
rect -17620 38880 -17380 38900
rect -17120 38880 -16880 38900
rect -16620 38880 -16380 38900
rect -16120 38880 -15880 38900
rect -15620 38880 -15380 38900
rect -15120 38880 -14880 38900
rect -14620 38880 -14380 38900
rect -14120 38880 -13880 38900
rect -13620 38880 -13380 38900
rect -13120 38880 -12880 38900
rect -12620 38880 -12380 38900
rect -12120 38880 -11880 38900
rect -11620 38880 -11380 38900
rect -11120 38880 -10880 38900
rect -10620 38880 -10380 38900
rect -10120 38880 -9880 38900
rect -9620 38880 -9380 38900
rect -9120 38880 -8880 38900
rect -8620 38880 -8380 38900
rect -8120 38880 -7880 38900
rect -7620 38880 -7380 38900
rect -7120 38880 -6880 38900
rect -6620 38880 -6380 38900
rect -6120 38880 -5880 38900
rect -5620 38880 -5380 38900
rect -5120 38880 -4880 38900
rect -4620 38880 -4380 38900
rect -4120 38880 -3880 38900
rect -3620 38880 -3380 38900
rect -3120 38880 -2880 38900
rect -2620 38880 -2380 38900
rect -2120 38880 -1880 38900
rect -1620 38880 -1380 38900
rect -1120 38880 -880 38900
rect -620 38880 -380 38900
rect -120 38880 120 38900
rect 380 38880 620 38900
rect 880 38880 1120 38900
rect 1380 38880 1620 38900
rect 1880 38880 2120 38900
rect 2380 38880 2620 38900
rect 2880 38880 3120 38900
rect 3380 38880 3620 38900
rect 3880 38880 4000 38900
rect -28000 38850 -27900 38880
rect -28000 38650 -27980 38850
rect -27910 38650 -27900 38850
rect -28000 38620 -27900 38650
rect -27600 38850 -27400 38880
rect -27600 38650 -27590 38850
rect -27520 38650 -27480 38850
rect -27410 38650 -27400 38850
rect -27600 38620 -27400 38650
rect -27100 38850 -26900 38880
rect -27100 38650 -27090 38850
rect -27020 38650 -26980 38850
rect -26910 38650 -26900 38850
rect -27100 38620 -26900 38650
rect -26600 38850 -26400 38880
rect -26600 38650 -26590 38850
rect -26520 38650 -26480 38850
rect -26410 38650 -26400 38850
rect -26600 38620 -26400 38650
rect -26100 38850 -25900 38880
rect -26100 38650 -26090 38850
rect -26020 38650 -25980 38850
rect -25910 38650 -25900 38850
rect -26100 38620 -25900 38650
rect -25600 38850 -25400 38880
rect -25600 38650 -25590 38850
rect -25520 38650 -25480 38850
rect -25410 38650 -25400 38850
rect -25600 38620 -25400 38650
rect -25100 38850 -24900 38880
rect -25100 38650 -25090 38850
rect -25020 38650 -24980 38850
rect -24910 38650 -24900 38850
rect -25100 38620 -24900 38650
rect -24600 38850 -24400 38880
rect -24600 38650 -24590 38850
rect -24520 38650 -24480 38850
rect -24410 38650 -24400 38850
rect -24600 38620 -24400 38650
rect -24100 38850 -23900 38880
rect -24100 38650 -24090 38850
rect -24020 38650 -23980 38850
rect -23910 38650 -23900 38850
rect -24100 38620 -23900 38650
rect -23600 38850 -23400 38880
rect -23600 38650 -23590 38850
rect -23520 38650 -23480 38850
rect -23410 38650 -23400 38850
rect -23600 38620 -23400 38650
rect -23100 38850 -22900 38880
rect -23100 38650 -23090 38850
rect -23020 38650 -22980 38850
rect -22910 38650 -22900 38850
rect -23100 38620 -22900 38650
rect -22600 38850 -22400 38880
rect -22600 38650 -22590 38850
rect -22520 38650 -22480 38850
rect -22410 38650 -22400 38850
rect -22600 38620 -22400 38650
rect -22100 38850 -21900 38880
rect -22100 38650 -22090 38850
rect -22020 38650 -21980 38850
rect -21910 38650 -21900 38850
rect -22100 38620 -21900 38650
rect -21600 38850 -21400 38880
rect -21600 38650 -21590 38850
rect -21520 38650 -21480 38850
rect -21410 38650 -21400 38850
rect -21600 38620 -21400 38650
rect -21100 38850 -20900 38880
rect -21100 38650 -21090 38850
rect -21020 38650 -20980 38850
rect -20910 38650 -20900 38850
rect -21100 38620 -20900 38650
rect -20600 38850 -20400 38880
rect -20600 38650 -20590 38850
rect -20520 38650 -20480 38850
rect -20410 38650 -20400 38850
rect -20600 38620 -20400 38650
rect -20100 38850 -19900 38880
rect -20100 38650 -20090 38850
rect -20020 38650 -19980 38850
rect -19910 38650 -19900 38850
rect -20100 38620 -19900 38650
rect -19600 38850 -19400 38880
rect -19600 38650 -19590 38850
rect -19520 38650 -19480 38850
rect -19410 38650 -19400 38850
rect -19600 38620 -19400 38650
rect -19100 38850 -18900 38880
rect -19100 38650 -19090 38850
rect -19020 38650 -18980 38850
rect -18910 38650 -18900 38850
rect -19100 38620 -18900 38650
rect -18600 38850 -18400 38880
rect -18600 38650 -18590 38850
rect -18520 38650 -18480 38850
rect -18410 38650 -18400 38850
rect -18600 38620 -18400 38650
rect -18100 38850 -17900 38880
rect -18100 38650 -18090 38850
rect -18020 38650 -17980 38850
rect -17910 38650 -17900 38850
rect -18100 38620 -17900 38650
rect -17600 38850 -17400 38880
rect -17600 38650 -17590 38850
rect -17520 38650 -17480 38850
rect -17410 38650 -17400 38850
rect -17600 38620 -17400 38650
rect -17100 38850 -16900 38880
rect -17100 38650 -17090 38850
rect -17020 38650 -16980 38850
rect -16910 38650 -16900 38850
rect -17100 38620 -16900 38650
rect -16600 38850 -16400 38880
rect -16600 38650 -16590 38850
rect -16520 38650 -16480 38850
rect -16410 38650 -16400 38850
rect -16600 38620 -16400 38650
rect -16100 38850 -15900 38880
rect -16100 38650 -16090 38850
rect -16020 38650 -15980 38850
rect -15910 38650 -15900 38850
rect -16100 38620 -15900 38650
rect -15600 38850 -15400 38880
rect -15600 38650 -15590 38850
rect -15520 38650 -15480 38850
rect -15410 38650 -15400 38850
rect -15600 38620 -15400 38650
rect -15100 38850 -14900 38880
rect -15100 38650 -15090 38850
rect -15020 38650 -14980 38850
rect -14910 38650 -14900 38850
rect -15100 38620 -14900 38650
rect -14600 38850 -14400 38880
rect -14600 38650 -14590 38850
rect -14520 38650 -14480 38850
rect -14410 38650 -14400 38850
rect -14600 38620 -14400 38650
rect -14100 38850 -13900 38880
rect -14100 38650 -14090 38850
rect -14020 38650 -13980 38850
rect -13910 38650 -13900 38850
rect -14100 38620 -13900 38650
rect -13600 38850 -13400 38880
rect -13600 38650 -13590 38850
rect -13520 38650 -13480 38850
rect -13410 38650 -13400 38850
rect -13600 38620 -13400 38650
rect -13100 38850 -12900 38880
rect -13100 38650 -13090 38850
rect -13020 38650 -12980 38850
rect -12910 38650 -12900 38850
rect -13100 38620 -12900 38650
rect -12600 38850 -12400 38880
rect -12600 38650 -12590 38850
rect -12520 38650 -12480 38850
rect -12410 38650 -12400 38850
rect -12600 38620 -12400 38650
rect -12100 38850 -11900 38880
rect -12100 38650 -12090 38850
rect -12020 38650 -11980 38850
rect -11910 38650 -11900 38850
rect -12100 38620 -11900 38650
rect -11600 38850 -11400 38880
rect -11600 38650 -11590 38850
rect -11520 38650 -11480 38850
rect -11410 38650 -11400 38850
rect -11600 38620 -11400 38650
rect -11100 38850 -10900 38880
rect -11100 38650 -11090 38850
rect -11020 38650 -10980 38850
rect -10910 38650 -10900 38850
rect -11100 38620 -10900 38650
rect -10600 38850 -10400 38880
rect -10600 38650 -10590 38850
rect -10520 38650 -10480 38850
rect -10410 38650 -10400 38850
rect -10600 38620 -10400 38650
rect -10100 38850 -9900 38880
rect -10100 38650 -10090 38850
rect -10020 38650 -9980 38850
rect -9910 38650 -9900 38850
rect -10100 38620 -9900 38650
rect -9600 38850 -9400 38880
rect -9600 38650 -9590 38850
rect -9520 38650 -9480 38850
rect -9410 38650 -9400 38850
rect -9600 38620 -9400 38650
rect -9100 38850 -8900 38880
rect -9100 38650 -9090 38850
rect -9020 38650 -8980 38850
rect -8910 38650 -8900 38850
rect -9100 38620 -8900 38650
rect -8600 38850 -8400 38880
rect -8600 38650 -8590 38850
rect -8520 38650 -8480 38850
rect -8410 38650 -8400 38850
rect -8600 38620 -8400 38650
rect -8100 38850 -7900 38880
rect -8100 38650 -8090 38850
rect -8020 38650 -7980 38850
rect -7910 38650 -7900 38850
rect -8100 38620 -7900 38650
rect -7600 38850 -7400 38880
rect -7600 38650 -7590 38850
rect -7520 38650 -7480 38850
rect -7410 38650 -7400 38850
rect -7600 38620 -7400 38650
rect -7100 38850 -6900 38880
rect -7100 38650 -7090 38850
rect -7020 38650 -6980 38850
rect -6910 38650 -6900 38850
rect -7100 38620 -6900 38650
rect -6600 38850 -6400 38880
rect -6600 38650 -6590 38850
rect -6520 38650 -6480 38850
rect -6410 38650 -6400 38850
rect -6600 38620 -6400 38650
rect -6100 38850 -5900 38880
rect -6100 38650 -6090 38850
rect -6020 38650 -5980 38850
rect -5910 38650 -5900 38850
rect -6100 38620 -5900 38650
rect -5600 38850 -5400 38880
rect -5600 38650 -5590 38850
rect -5520 38650 -5480 38850
rect -5410 38650 -5400 38850
rect -5600 38620 -5400 38650
rect -5100 38850 -4900 38880
rect -5100 38650 -5090 38850
rect -5020 38650 -4980 38850
rect -4910 38650 -4900 38850
rect -5100 38620 -4900 38650
rect -4600 38850 -4400 38880
rect -4600 38650 -4590 38850
rect -4520 38650 -4480 38850
rect -4410 38650 -4400 38850
rect -4600 38620 -4400 38650
rect -4100 38850 -3900 38880
rect -4100 38650 -4090 38850
rect -4020 38650 -3980 38850
rect -3910 38650 -3900 38850
rect -4100 38620 -3900 38650
rect -3600 38850 -3400 38880
rect -3600 38650 -3590 38850
rect -3520 38650 -3480 38850
rect -3410 38650 -3400 38850
rect -3600 38620 -3400 38650
rect -3100 38850 -2900 38880
rect -3100 38650 -3090 38850
rect -3020 38650 -2980 38850
rect -2910 38650 -2900 38850
rect -3100 38620 -2900 38650
rect -2600 38850 -2400 38880
rect -2600 38650 -2590 38850
rect -2520 38650 -2480 38850
rect -2410 38650 -2400 38850
rect -2600 38620 -2400 38650
rect -2100 38850 -1900 38880
rect -2100 38650 -2090 38850
rect -2020 38650 -1980 38850
rect -1910 38650 -1900 38850
rect -2100 38620 -1900 38650
rect -1600 38850 -1400 38880
rect -1600 38650 -1590 38850
rect -1520 38650 -1480 38850
rect -1410 38650 -1400 38850
rect -1600 38620 -1400 38650
rect -1100 38850 -900 38880
rect -1100 38650 -1090 38850
rect -1020 38650 -980 38850
rect -910 38650 -900 38850
rect -1100 38620 -900 38650
rect -600 38850 -400 38880
rect -600 38650 -590 38850
rect -520 38650 -480 38850
rect -410 38650 -400 38850
rect -600 38620 -400 38650
rect -100 38850 100 38880
rect -100 38650 -90 38850
rect -20 38650 20 38850
rect 90 38650 100 38850
rect -100 38620 100 38650
rect 400 38850 600 38880
rect 400 38650 410 38850
rect 480 38650 520 38850
rect 590 38650 600 38850
rect 400 38620 600 38650
rect 900 38850 1100 38880
rect 900 38650 910 38850
rect 980 38650 1020 38850
rect 1090 38650 1100 38850
rect 900 38620 1100 38650
rect 1400 38850 1600 38880
rect 1400 38650 1410 38850
rect 1480 38650 1520 38850
rect 1590 38650 1600 38850
rect 1400 38620 1600 38650
rect 1900 38850 2100 38880
rect 1900 38650 1910 38850
rect 1980 38650 2020 38850
rect 2090 38650 2100 38850
rect 1900 38620 2100 38650
rect 2400 38850 2600 38880
rect 2400 38650 2410 38850
rect 2480 38650 2520 38850
rect 2590 38650 2600 38850
rect 2400 38620 2600 38650
rect 2900 38850 3100 38880
rect 2900 38650 2910 38850
rect 2980 38650 3020 38850
rect 3090 38650 3100 38850
rect 2900 38620 3100 38650
rect 3400 38850 3600 38880
rect 3400 38650 3410 38850
rect 3480 38650 3520 38850
rect 3590 38650 3600 38850
rect 3400 38620 3600 38650
rect 3900 38850 4000 38880
rect 3900 38650 3910 38850
rect 3980 38650 4000 38850
rect 3900 38620 4000 38650
rect -28000 38600 -27880 38620
rect -27620 38600 -27380 38620
rect -27120 38600 -26880 38620
rect -26620 38600 -26380 38620
rect -26120 38600 -25880 38620
rect -25620 38600 -25380 38620
rect -25120 38600 -24880 38620
rect -24620 38600 -24380 38620
rect -24120 38600 -23880 38620
rect -23620 38600 -23380 38620
rect -23120 38600 -22880 38620
rect -22620 38600 -22380 38620
rect -22120 38600 -21880 38620
rect -21620 38600 -21380 38620
rect -21120 38600 -20880 38620
rect -20620 38600 -20380 38620
rect -20120 38600 -19880 38620
rect -19620 38600 -19380 38620
rect -19120 38600 -18880 38620
rect -18620 38600 -18380 38620
rect -18120 38600 -17880 38620
rect -17620 38600 -17380 38620
rect -17120 38600 -16880 38620
rect -16620 38600 -16380 38620
rect -16120 38600 -15880 38620
rect -15620 38600 -15380 38620
rect -15120 38600 -14880 38620
rect -14620 38600 -14380 38620
rect -14120 38600 -13880 38620
rect -13620 38600 -13380 38620
rect -13120 38600 -12880 38620
rect -12620 38600 -12380 38620
rect -12120 38600 -11880 38620
rect -11620 38600 -11380 38620
rect -11120 38600 -10880 38620
rect -10620 38600 -10380 38620
rect -10120 38600 -9880 38620
rect -9620 38600 -9380 38620
rect -9120 38600 -8880 38620
rect -8620 38600 -8380 38620
rect -8120 38600 -7880 38620
rect -7620 38600 -7380 38620
rect -7120 38600 -6880 38620
rect -6620 38600 -6380 38620
rect -6120 38600 -5880 38620
rect -5620 38600 -5380 38620
rect -5120 38600 -4880 38620
rect -4620 38600 -4380 38620
rect -4120 38600 -3880 38620
rect -3620 38600 -3380 38620
rect -3120 38600 -2880 38620
rect -2620 38600 -2380 38620
rect -2120 38600 -1880 38620
rect -1620 38600 -1380 38620
rect -1120 38600 -880 38620
rect -620 38600 -380 38620
rect -120 38600 120 38620
rect 380 38600 620 38620
rect 880 38600 1120 38620
rect 1380 38600 1620 38620
rect 1880 38600 2120 38620
rect 2380 38600 2620 38620
rect 2880 38600 3120 38620
rect 3380 38600 3620 38620
rect 3880 38600 4000 38620
rect -28000 38590 4000 38600
rect -28000 38520 -27850 38590
rect -27650 38520 -27350 38590
rect -27150 38520 -26850 38590
rect -26650 38520 -26350 38590
rect -26150 38520 -25850 38590
rect -25650 38520 -25350 38590
rect -25150 38520 -24850 38590
rect -24650 38520 -24350 38590
rect -24150 38520 -23850 38590
rect -23650 38520 -23350 38590
rect -23150 38520 -22850 38590
rect -22650 38520 -22350 38590
rect -22150 38520 -21850 38590
rect -21650 38520 -21350 38590
rect -21150 38520 -20850 38590
rect -20650 38520 -20350 38590
rect -20150 38520 -19850 38590
rect -19650 38520 -19350 38590
rect -19150 38520 -18850 38590
rect -18650 38520 -18350 38590
rect -18150 38520 -17850 38590
rect -17650 38520 -17350 38590
rect -17150 38520 -16850 38590
rect -16650 38520 -16350 38590
rect -16150 38520 -15850 38590
rect -15650 38520 -15350 38590
rect -15150 38520 -14850 38590
rect -14650 38520 -14350 38590
rect -14150 38520 -13850 38590
rect -13650 38520 -13350 38590
rect -13150 38520 -12850 38590
rect -12650 38520 -12350 38590
rect -12150 38520 -11850 38590
rect -11650 38520 -11350 38590
rect -11150 38520 -10850 38590
rect -10650 38520 -10350 38590
rect -10150 38520 -9850 38590
rect -9650 38520 -9350 38590
rect -9150 38520 -8850 38590
rect -8650 38520 -8350 38590
rect -8150 38520 -7850 38590
rect -7650 38520 -7350 38590
rect -7150 38520 -6850 38590
rect -6650 38520 -6350 38590
rect -6150 38520 -5850 38590
rect -5650 38520 -5350 38590
rect -5150 38520 -4850 38590
rect -4650 38520 -4350 38590
rect -4150 38520 -3850 38590
rect -3650 38520 -3350 38590
rect -3150 38520 -2850 38590
rect -2650 38520 -2350 38590
rect -2150 38520 -1850 38590
rect -1650 38520 -1350 38590
rect -1150 38520 -850 38590
rect -650 38520 -350 38590
rect -150 38520 150 38590
rect 350 38520 650 38590
rect 850 38520 1150 38590
rect 1350 38520 1650 38590
rect 1850 38520 2150 38590
rect 2350 38520 2650 38590
rect 2850 38520 3150 38590
rect 3350 38520 3650 38590
rect 3850 38520 4000 38590
rect -28000 38480 4000 38520
rect -28000 38410 -27850 38480
rect -27650 38410 -27350 38480
rect -27150 38410 -26850 38480
rect -26650 38410 -26350 38480
rect -26150 38410 -25850 38480
rect -25650 38410 -25350 38480
rect -25150 38410 -24850 38480
rect -24650 38410 -24350 38480
rect -24150 38410 -23850 38480
rect -23650 38410 -23350 38480
rect -23150 38410 -22850 38480
rect -22650 38410 -22350 38480
rect -22150 38410 -21850 38480
rect -21650 38410 -21350 38480
rect -21150 38410 -20850 38480
rect -20650 38410 -20350 38480
rect -20150 38410 -19850 38480
rect -19650 38410 -19350 38480
rect -19150 38410 -18850 38480
rect -18650 38410 -18350 38480
rect -18150 38410 -17850 38480
rect -17650 38410 -17350 38480
rect -17150 38410 -16850 38480
rect -16650 38410 -16350 38480
rect -16150 38410 -15850 38480
rect -15650 38410 -15350 38480
rect -15150 38410 -14850 38480
rect -14650 38410 -14350 38480
rect -14150 38410 -13850 38480
rect -13650 38410 -13350 38480
rect -13150 38410 -12850 38480
rect -12650 38410 -12350 38480
rect -12150 38410 -11850 38480
rect -11650 38410 -11350 38480
rect -11150 38410 -10850 38480
rect -10650 38410 -10350 38480
rect -10150 38410 -9850 38480
rect -9650 38410 -9350 38480
rect -9150 38410 -8850 38480
rect -8650 38410 -8350 38480
rect -8150 38410 -7850 38480
rect -7650 38410 -7350 38480
rect -7150 38410 -6850 38480
rect -6650 38410 -6350 38480
rect -6150 38410 -5850 38480
rect -5650 38410 -5350 38480
rect -5150 38410 -4850 38480
rect -4650 38410 -4350 38480
rect -4150 38410 -3850 38480
rect -3650 38410 -3350 38480
rect -3150 38410 -2850 38480
rect -2650 38410 -2350 38480
rect -2150 38410 -1850 38480
rect -1650 38410 -1350 38480
rect -1150 38410 -850 38480
rect -650 38410 -350 38480
rect -150 38410 150 38480
rect 350 38410 650 38480
rect 850 38410 1150 38480
rect 1350 38410 1650 38480
rect 1850 38410 2150 38480
rect 2350 38410 2650 38480
rect 2850 38410 3150 38480
rect 3350 38410 3650 38480
rect 3850 38410 4000 38480
rect -28000 38400 4000 38410
rect -28000 38380 -27880 38400
rect -27620 38380 -27380 38400
rect -27120 38380 -26880 38400
rect -26620 38380 -26380 38400
rect -26120 38380 -25880 38400
rect -25620 38380 -25380 38400
rect -25120 38380 -24880 38400
rect -24620 38380 -24380 38400
rect -24120 38380 -23880 38400
rect -23620 38380 -23380 38400
rect -23120 38380 -22880 38400
rect -22620 38380 -22380 38400
rect -22120 38380 -21880 38400
rect -21620 38380 -21380 38400
rect -21120 38380 -20880 38400
rect -20620 38380 -20380 38400
rect -20120 38380 -19880 38400
rect -19620 38380 -19380 38400
rect -19120 38380 -18880 38400
rect -18620 38380 -18380 38400
rect -18120 38380 -17880 38400
rect -17620 38380 -17380 38400
rect -17120 38380 -16880 38400
rect -16620 38380 -16380 38400
rect -16120 38380 -15880 38400
rect -15620 38380 -15380 38400
rect -15120 38380 -14880 38400
rect -14620 38380 -14380 38400
rect -14120 38380 -13880 38400
rect -13620 38380 -13380 38400
rect -13120 38380 -12880 38400
rect -12620 38380 -12380 38400
rect -12120 38380 -11880 38400
rect -11620 38380 -11380 38400
rect -11120 38380 -10880 38400
rect -10620 38380 -10380 38400
rect -10120 38380 -9880 38400
rect -9620 38380 -9380 38400
rect -9120 38380 -8880 38400
rect -8620 38380 -8380 38400
rect -8120 38380 -7880 38400
rect -7620 38380 -7380 38400
rect -7120 38380 -6880 38400
rect -6620 38380 -6380 38400
rect -6120 38380 -5880 38400
rect -5620 38380 -5380 38400
rect -5120 38380 -4880 38400
rect -4620 38380 -4380 38400
rect -4120 38380 -3880 38400
rect -3620 38380 -3380 38400
rect -3120 38380 -2880 38400
rect -2620 38380 -2380 38400
rect -2120 38380 -1880 38400
rect -1620 38380 -1380 38400
rect -1120 38380 -880 38400
rect -620 38380 -380 38400
rect -120 38380 120 38400
rect 380 38380 620 38400
rect 880 38380 1120 38400
rect 1380 38380 1620 38400
rect 1880 38380 2120 38400
rect 2380 38380 2620 38400
rect 2880 38380 3120 38400
rect 3380 38380 3620 38400
rect 3880 38380 4000 38400
rect -28000 38350 -27900 38380
rect -28000 38150 -27980 38350
rect -27910 38150 -27900 38350
rect -28000 38120 -27900 38150
rect -27600 38350 -27400 38380
rect -27600 38150 -27590 38350
rect -27520 38150 -27480 38350
rect -27410 38150 -27400 38350
rect -27600 38120 -27400 38150
rect -27100 38350 -26900 38380
rect -27100 38150 -27090 38350
rect -27020 38150 -26980 38350
rect -26910 38150 -26900 38350
rect -27100 38120 -26900 38150
rect -26600 38350 -26400 38380
rect -26600 38150 -26590 38350
rect -26520 38150 -26480 38350
rect -26410 38150 -26400 38350
rect -26600 38120 -26400 38150
rect -26100 38350 -25900 38380
rect -26100 38150 -26090 38350
rect -26020 38150 -25980 38350
rect -25910 38150 -25900 38350
rect -26100 38120 -25900 38150
rect -25600 38350 -25400 38380
rect -25600 38150 -25590 38350
rect -25520 38150 -25480 38350
rect -25410 38150 -25400 38350
rect -25600 38120 -25400 38150
rect -25100 38350 -24900 38380
rect -25100 38150 -25090 38350
rect -25020 38150 -24980 38350
rect -24910 38150 -24900 38350
rect -25100 38120 -24900 38150
rect -24600 38350 -24400 38380
rect -24600 38150 -24590 38350
rect -24520 38150 -24480 38350
rect -24410 38150 -24400 38350
rect -24600 38120 -24400 38150
rect -24100 38350 -23900 38380
rect -24100 38150 -24090 38350
rect -24020 38150 -23980 38350
rect -23910 38150 -23900 38350
rect -24100 38120 -23900 38150
rect -23600 38350 -23400 38380
rect -23600 38150 -23590 38350
rect -23520 38150 -23480 38350
rect -23410 38150 -23400 38350
rect -23600 38120 -23400 38150
rect -23100 38350 -22900 38380
rect -23100 38150 -23090 38350
rect -23020 38150 -22980 38350
rect -22910 38150 -22900 38350
rect -23100 38120 -22900 38150
rect -22600 38350 -22400 38380
rect -22600 38150 -22590 38350
rect -22520 38150 -22480 38350
rect -22410 38150 -22400 38350
rect -22600 38120 -22400 38150
rect -22100 38350 -21900 38380
rect -22100 38150 -22090 38350
rect -22020 38150 -21980 38350
rect -21910 38150 -21900 38350
rect -22100 38120 -21900 38150
rect -21600 38350 -21400 38380
rect -21600 38150 -21590 38350
rect -21520 38150 -21480 38350
rect -21410 38150 -21400 38350
rect -21600 38120 -21400 38150
rect -21100 38350 -20900 38380
rect -21100 38150 -21090 38350
rect -21020 38150 -20980 38350
rect -20910 38150 -20900 38350
rect -21100 38120 -20900 38150
rect -20600 38350 -20400 38380
rect -20600 38150 -20590 38350
rect -20520 38150 -20480 38350
rect -20410 38150 -20400 38350
rect -20600 38120 -20400 38150
rect -20100 38350 -19900 38380
rect -20100 38150 -20090 38350
rect -20020 38150 -19980 38350
rect -19910 38150 -19900 38350
rect -20100 38120 -19900 38150
rect -19600 38350 -19400 38380
rect -19600 38150 -19590 38350
rect -19520 38150 -19480 38350
rect -19410 38150 -19400 38350
rect -19600 38120 -19400 38150
rect -19100 38350 -18900 38380
rect -19100 38150 -19090 38350
rect -19020 38150 -18980 38350
rect -18910 38150 -18900 38350
rect -19100 38120 -18900 38150
rect -18600 38350 -18400 38380
rect -18600 38150 -18590 38350
rect -18520 38150 -18480 38350
rect -18410 38150 -18400 38350
rect -18600 38120 -18400 38150
rect -18100 38350 -17900 38380
rect -18100 38150 -18090 38350
rect -18020 38150 -17980 38350
rect -17910 38150 -17900 38350
rect -18100 38120 -17900 38150
rect -17600 38350 -17400 38380
rect -17600 38150 -17590 38350
rect -17520 38150 -17480 38350
rect -17410 38150 -17400 38350
rect -17600 38120 -17400 38150
rect -17100 38350 -16900 38380
rect -17100 38150 -17090 38350
rect -17020 38150 -16980 38350
rect -16910 38150 -16900 38350
rect -17100 38120 -16900 38150
rect -16600 38350 -16400 38380
rect -16600 38150 -16590 38350
rect -16520 38150 -16480 38350
rect -16410 38150 -16400 38350
rect -16600 38120 -16400 38150
rect -16100 38350 -15900 38380
rect -16100 38150 -16090 38350
rect -16020 38150 -15980 38350
rect -15910 38150 -15900 38350
rect -16100 38120 -15900 38150
rect -15600 38350 -15400 38380
rect -15600 38150 -15590 38350
rect -15520 38150 -15480 38350
rect -15410 38150 -15400 38350
rect -15600 38120 -15400 38150
rect -15100 38350 -14900 38380
rect -15100 38150 -15090 38350
rect -15020 38150 -14980 38350
rect -14910 38150 -14900 38350
rect -15100 38120 -14900 38150
rect -14600 38350 -14400 38380
rect -14600 38150 -14590 38350
rect -14520 38150 -14480 38350
rect -14410 38150 -14400 38350
rect -14600 38120 -14400 38150
rect -14100 38350 -13900 38380
rect -14100 38150 -14090 38350
rect -14020 38150 -13980 38350
rect -13910 38150 -13900 38350
rect -14100 38120 -13900 38150
rect -13600 38350 -13400 38380
rect -13600 38150 -13590 38350
rect -13520 38150 -13480 38350
rect -13410 38150 -13400 38350
rect -13600 38120 -13400 38150
rect -13100 38350 -12900 38380
rect -13100 38150 -13090 38350
rect -13020 38150 -12980 38350
rect -12910 38150 -12900 38350
rect -13100 38120 -12900 38150
rect -12600 38350 -12400 38380
rect -12600 38150 -12590 38350
rect -12520 38150 -12480 38350
rect -12410 38150 -12400 38350
rect -12600 38120 -12400 38150
rect -12100 38350 -11900 38380
rect -12100 38150 -12090 38350
rect -12020 38150 -11980 38350
rect -11910 38150 -11900 38350
rect -12100 38120 -11900 38150
rect -11600 38350 -11400 38380
rect -11600 38150 -11590 38350
rect -11520 38150 -11480 38350
rect -11410 38150 -11400 38350
rect -11600 38120 -11400 38150
rect -11100 38350 -10900 38380
rect -11100 38150 -11090 38350
rect -11020 38150 -10980 38350
rect -10910 38150 -10900 38350
rect -11100 38120 -10900 38150
rect -10600 38350 -10400 38380
rect -10600 38150 -10590 38350
rect -10520 38150 -10480 38350
rect -10410 38150 -10400 38350
rect -10600 38120 -10400 38150
rect -10100 38350 -9900 38380
rect -10100 38150 -10090 38350
rect -10020 38150 -9980 38350
rect -9910 38150 -9900 38350
rect -10100 38120 -9900 38150
rect -9600 38350 -9400 38380
rect -9600 38150 -9590 38350
rect -9520 38150 -9480 38350
rect -9410 38150 -9400 38350
rect -9600 38120 -9400 38150
rect -9100 38350 -8900 38380
rect -9100 38150 -9090 38350
rect -9020 38150 -8980 38350
rect -8910 38150 -8900 38350
rect -9100 38120 -8900 38150
rect -8600 38350 -8400 38380
rect -8600 38150 -8590 38350
rect -8520 38150 -8480 38350
rect -8410 38150 -8400 38350
rect -8600 38120 -8400 38150
rect -8100 38350 -7900 38380
rect -8100 38150 -8090 38350
rect -8020 38150 -7980 38350
rect -7910 38150 -7900 38350
rect -8100 38120 -7900 38150
rect -7600 38350 -7400 38380
rect -7600 38150 -7590 38350
rect -7520 38150 -7480 38350
rect -7410 38150 -7400 38350
rect -7600 38120 -7400 38150
rect -7100 38350 -6900 38380
rect -7100 38150 -7090 38350
rect -7020 38150 -6980 38350
rect -6910 38150 -6900 38350
rect -7100 38120 -6900 38150
rect -6600 38350 -6400 38380
rect -6600 38150 -6590 38350
rect -6520 38150 -6480 38350
rect -6410 38150 -6400 38350
rect -6600 38120 -6400 38150
rect -6100 38350 -5900 38380
rect -6100 38150 -6090 38350
rect -6020 38150 -5980 38350
rect -5910 38150 -5900 38350
rect -6100 38120 -5900 38150
rect -5600 38350 -5400 38380
rect -5600 38150 -5590 38350
rect -5520 38150 -5480 38350
rect -5410 38150 -5400 38350
rect -5600 38120 -5400 38150
rect -5100 38350 -4900 38380
rect -5100 38150 -5090 38350
rect -5020 38150 -4980 38350
rect -4910 38150 -4900 38350
rect -5100 38120 -4900 38150
rect -4600 38350 -4400 38380
rect -4600 38150 -4590 38350
rect -4520 38150 -4480 38350
rect -4410 38150 -4400 38350
rect -4600 38120 -4400 38150
rect -4100 38350 -3900 38380
rect -4100 38150 -4090 38350
rect -4020 38150 -3980 38350
rect -3910 38150 -3900 38350
rect -4100 38120 -3900 38150
rect -3600 38350 -3400 38380
rect -3600 38150 -3590 38350
rect -3520 38150 -3480 38350
rect -3410 38150 -3400 38350
rect -3600 38120 -3400 38150
rect -3100 38350 -2900 38380
rect -3100 38150 -3090 38350
rect -3020 38150 -2980 38350
rect -2910 38150 -2900 38350
rect -3100 38120 -2900 38150
rect -2600 38350 -2400 38380
rect -2600 38150 -2590 38350
rect -2520 38150 -2480 38350
rect -2410 38150 -2400 38350
rect -2600 38120 -2400 38150
rect -2100 38350 -1900 38380
rect -2100 38150 -2090 38350
rect -2020 38150 -1980 38350
rect -1910 38150 -1900 38350
rect -2100 38120 -1900 38150
rect -1600 38350 -1400 38380
rect -1600 38150 -1590 38350
rect -1520 38150 -1480 38350
rect -1410 38150 -1400 38350
rect -1600 38120 -1400 38150
rect -1100 38350 -900 38380
rect -1100 38150 -1090 38350
rect -1020 38150 -980 38350
rect -910 38150 -900 38350
rect -1100 38120 -900 38150
rect -600 38350 -400 38380
rect -600 38150 -590 38350
rect -520 38150 -480 38350
rect -410 38150 -400 38350
rect -600 38120 -400 38150
rect -100 38350 100 38380
rect -100 38150 -90 38350
rect -20 38150 20 38350
rect 90 38150 100 38350
rect -100 38120 100 38150
rect 400 38350 600 38380
rect 400 38150 410 38350
rect 480 38150 520 38350
rect 590 38150 600 38350
rect 400 38120 600 38150
rect 900 38350 1100 38380
rect 900 38150 910 38350
rect 980 38150 1020 38350
rect 1090 38150 1100 38350
rect 900 38120 1100 38150
rect 1400 38350 1600 38380
rect 1400 38150 1410 38350
rect 1480 38150 1520 38350
rect 1590 38150 1600 38350
rect 1400 38120 1600 38150
rect 1900 38350 2100 38380
rect 1900 38150 1910 38350
rect 1980 38150 2020 38350
rect 2090 38150 2100 38350
rect 1900 38120 2100 38150
rect 2400 38350 2600 38380
rect 2400 38150 2410 38350
rect 2480 38150 2520 38350
rect 2590 38150 2600 38350
rect 2400 38120 2600 38150
rect 2900 38350 3100 38380
rect 2900 38150 2910 38350
rect 2980 38150 3020 38350
rect 3090 38150 3100 38350
rect 2900 38120 3100 38150
rect 3400 38350 3600 38380
rect 3400 38150 3410 38350
rect 3480 38150 3520 38350
rect 3590 38150 3600 38350
rect 3400 38120 3600 38150
rect 3900 38350 4000 38380
rect 3900 38150 3910 38350
rect 3980 38150 4000 38350
rect 3900 38120 4000 38150
rect -28000 38100 -27880 38120
rect -27620 38100 -27380 38120
rect -27120 38100 -26880 38120
rect -26620 38100 -26380 38120
rect -26120 38100 -25880 38120
rect -25620 38100 -25380 38120
rect -25120 38100 -24880 38120
rect -24620 38100 -24380 38120
rect -24120 38100 -23880 38120
rect -23620 38100 -23380 38120
rect -23120 38100 -22880 38120
rect -22620 38100 -22380 38120
rect -22120 38100 -21880 38120
rect -21620 38100 -21380 38120
rect -21120 38100 -20880 38120
rect -20620 38100 -20380 38120
rect -20120 38100 -19880 38120
rect -19620 38100 -19380 38120
rect -19120 38100 -18880 38120
rect -18620 38100 -18380 38120
rect -18120 38100 -17880 38120
rect -17620 38100 -17380 38120
rect -17120 38100 -16880 38120
rect -16620 38100 -16380 38120
rect -16120 38100 -15880 38120
rect -15620 38100 -15380 38120
rect -15120 38100 -14880 38120
rect -14620 38100 -14380 38120
rect -14120 38100 -13880 38120
rect -13620 38100 -13380 38120
rect -13120 38100 -12880 38120
rect -12620 38100 -12380 38120
rect -12120 38100 -11880 38120
rect -11620 38100 -11380 38120
rect -11120 38100 -10880 38120
rect -10620 38100 -10380 38120
rect -10120 38100 -9880 38120
rect -9620 38100 -9380 38120
rect -9120 38100 -8880 38120
rect -8620 38100 -8380 38120
rect -8120 38100 -7880 38120
rect -7620 38100 -7380 38120
rect -7120 38100 -6880 38120
rect -6620 38100 -6380 38120
rect -6120 38100 -5880 38120
rect -5620 38100 -5380 38120
rect -5120 38100 -4880 38120
rect -4620 38100 -4380 38120
rect -4120 38100 -3880 38120
rect -3620 38100 -3380 38120
rect -3120 38100 -2880 38120
rect -2620 38100 -2380 38120
rect -2120 38100 -1880 38120
rect -1620 38100 -1380 38120
rect -1120 38100 -880 38120
rect -620 38100 -380 38120
rect -120 38100 120 38120
rect 380 38100 620 38120
rect 880 38100 1120 38120
rect 1380 38100 1620 38120
rect 1880 38100 2120 38120
rect 2380 38100 2620 38120
rect 2880 38100 3120 38120
rect 3380 38100 3620 38120
rect 3880 38100 4000 38120
rect -28000 38090 4000 38100
rect -28000 38020 -27850 38090
rect -27650 38020 -27350 38090
rect -27150 38020 -26850 38090
rect -26650 38020 -26350 38090
rect -26150 38020 -25850 38090
rect -25650 38020 -25350 38090
rect -25150 38020 -24850 38090
rect -24650 38020 -24350 38090
rect -24150 38020 -23850 38090
rect -23650 38020 -23350 38090
rect -23150 38020 -22850 38090
rect -22650 38020 -22350 38090
rect -22150 38020 -21850 38090
rect -21650 38020 -21350 38090
rect -21150 38020 -20850 38090
rect -20650 38020 -20350 38090
rect -20150 38020 -19850 38090
rect -19650 38020 -19350 38090
rect -19150 38020 -18850 38090
rect -18650 38020 -18350 38090
rect -18150 38020 -17850 38090
rect -17650 38020 -17350 38090
rect -17150 38020 -16850 38090
rect -16650 38020 -16350 38090
rect -16150 38020 -15850 38090
rect -15650 38020 -15350 38090
rect -15150 38020 -14850 38090
rect -14650 38020 -14350 38090
rect -14150 38020 -13850 38090
rect -13650 38020 -13350 38090
rect -13150 38020 -12850 38090
rect -12650 38020 -12350 38090
rect -12150 38020 -11850 38090
rect -11650 38020 -11350 38090
rect -11150 38020 -10850 38090
rect -10650 38020 -10350 38090
rect -10150 38020 -9850 38090
rect -9650 38020 -9350 38090
rect -9150 38020 -8850 38090
rect -8650 38020 -8350 38090
rect -8150 38020 -7850 38090
rect -7650 38020 -7350 38090
rect -7150 38020 -6850 38090
rect -6650 38020 -6350 38090
rect -6150 38020 -5850 38090
rect -5650 38020 -5350 38090
rect -5150 38020 -4850 38090
rect -4650 38020 -4350 38090
rect -4150 38020 -3850 38090
rect -3650 38020 -3350 38090
rect -3150 38020 -2850 38090
rect -2650 38020 -2350 38090
rect -2150 38020 -1850 38090
rect -1650 38020 -1350 38090
rect -1150 38020 -850 38090
rect -650 38020 -350 38090
rect -150 38020 150 38090
rect 350 38020 650 38090
rect 850 38020 1150 38090
rect 1350 38020 1650 38090
rect 1850 38020 2150 38090
rect 2350 38020 2650 38090
rect 2850 38020 3150 38090
rect 3350 38020 3650 38090
rect 3850 38020 4000 38090
rect -28000 38000 4000 38020
rect 92000 37900 96000 38000
rect 92000 37880 92120 37900
rect 92380 37880 92620 37900
rect 92880 37880 93120 37900
rect 93380 37880 93620 37900
rect 93880 37880 94120 37900
rect 94380 37880 94620 37900
rect 94880 37880 95120 37900
rect 95380 37880 95620 37900
rect 95880 37880 96000 37900
rect 92000 37620 92100 37880
rect 92400 37620 92600 37880
rect 92900 37620 93100 37880
rect 93400 37620 93600 37880
rect 93900 37620 94100 37880
rect 94400 37620 94600 37880
rect 94900 37620 95100 37880
rect 95400 37620 95600 37880
rect 95900 37620 96000 37880
rect 92000 37600 92120 37620
rect 92380 37600 92620 37620
rect 92880 37600 93120 37620
rect 93380 37600 93620 37620
rect 93880 37600 94120 37620
rect 94380 37600 94620 37620
rect 94880 37600 95120 37620
rect 95380 37600 95620 37620
rect 95880 37600 96000 37620
rect 92000 37400 96000 37600
rect 92000 37380 92120 37400
rect 92380 37380 92620 37400
rect 92880 37380 93120 37400
rect 93380 37380 93620 37400
rect 93880 37380 94120 37400
rect 94380 37380 94620 37400
rect 94880 37380 95120 37400
rect 95380 37380 95620 37400
rect 95880 37380 96000 37400
rect 92000 37120 92100 37380
rect 92400 37120 92600 37380
rect 92900 37120 93100 37380
rect 93400 37120 93600 37380
rect 93900 37120 94100 37380
rect 94400 37120 94600 37380
rect 94900 37120 95100 37380
rect 95400 37120 95600 37380
rect 95900 37120 96000 37380
rect 92000 37100 92120 37120
rect 92380 37100 92620 37120
rect 92880 37100 93120 37120
rect 93380 37100 93620 37120
rect 93880 37100 94120 37120
rect 94380 37100 94620 37120
rect 94880 37100 95120 37120
rect 95380 37100 95620 37120
rect 95880 37100 96000 37120
rect 92000 36900 96000 37100
rect 92000 36880 92120 36900
rect 92380 36880 92620 36900
rect 92880 36880 93120 36900
rect 93380 36880 93620 36900
rect 93880 36880 94120 36900
rect 94380 36880 94620 36900
rect 94880 36880 95120 36900
rect 95380 36880 95620 36900
rect 95880 36880 96000 36900
rect 92000 36620 92100 36880
rect 92400 36620 92600 36880
rect 92900 36620 93100 36880
rect 93400 36620 93600 36880
rect 93900 36620 94100 36880
rect 94400 36620 94600 36880
rect 94900 36620 95100 36880
rect 95400 36620 95600 36880
rect 95900 36620 96000 36880
rect 92000 36600 92120 36620
rect 92380 36600 92620 36620
rect 92880 36600 93120 36620
rect 93380 36600 93620 36620
rect 93880 36600 94120 36620
rect 94380 36600 94620 36620
rect 94880 36600 95120 36620
rect 95380 36600 95620 36620
rect 95880 36600 96000 36620
rect 92000 36400 96000 36600
rect 92000 36380 92120 36400
rect 92380 36380 92620 36400
rect 92880 36380 93120 36400
rect 93380 36380 93620 36400
rect 93880 36380 94120 36400
rect 94380 36380 94620 36400
rect 94880 36380 95120 36400
rect 95380 36380 95620 36400
rect 95880 36380 96000 36400
rect 92000 36120 92100 36380
rect 92400 36120 92600 36380
rect 92900 36120 93100 36380
rect 93400 36120 93600 36380
rect 93900 36120 94100 36380
rect 94400 36120 94600 36380
rect 94900 36120 95100 36380
rect 95400 36120 95600 36380
rect 95900 36120 96000 36380
rect 92000 36100 92120 36120
rect 92380 36100 92620 36120
rect 92880 36100 93120 36120
rect 93380 36100 93620 36120
rect 93880 36100 94120 36120
rect 94380 36100 94620 36120
rect 94880 36100 95120 36120
rect 95380 36100 95620 36120
rect 95880 36100 96000 36120
rect 92000 35900 96000 36100
rect 92000 35880 92120 35900
rect 92380 35880 92620 35900
rect 92880 35880 93120 35900
rect 93380 35880 93620 35900
rect 93880 35880 94120 35900
rect 94380 35880 94620 35900
rect 94880 35880 95120 35900
rect 95380 35880 95620 35900
rect 95880 35880 96000 35900
rect 92000 35620 92100 35880
rect 92400 35620 92600 35880
rect 92900 35620 93100 35880
rect 93400 35620 93600 35880
rect 93900 35620 94100 35880
rect 94400 35620 94600 35880
rect 94900 35620 95100 35880
rect 95400 35620 95600 35880
rect 95900 35620 96000 35880
rect 92000 35600 92120 35620
rect 92380 35600 92620 35620
rect 92880 35600 93120 35620
rect 93380 35600 93620 35620
rect 93880 35600 94120 35620
rect 94380 35600 94620 35620
rect 94880 35600 95120 35620
rect 95380 35600 95620 35620
rect 95880 35600 96000 35620
rect 92000 35400 96000 35600
rect 92000 35380 92120 35400
rect 92380 35380 92620 35400
rect 92880 35380 93120 35400
rect 93380 35380 93620 35400
rect 93880 35380 94120 35400
rect 94380 35380 94620 35400
rect 94880 35380 95120 35400
rect 95380 35380 95620 35400
rect 95880 35380 96000 35400
rect 92000 35120 92100 35380
rect 92400 35120 92600 35380
rect 92900 35120 93100 35380
rect 93400 35120 93600 35380
rect 93900 35120 94100 35380
rect 94400 35120 94600 35380
rect 94900 35120 95100 35380
rect 95400 35120 95600 35380
rect 95900 35120 96000 35380
rect 92000 35100 92120 35120
rect 92380 35100 92620 35120
rect 92880 35100 93120 35120
rect 93380 35100 93620 35120
rect 93880 35100 94120 35120
rect 94380 35100 94620 35120
rect 94880 35100 95120 35120
rect 95380 35100 95620 35120
rect 95880 35100 96000 35120
rect 92000 34900 96000 35100
rect 92000 34880 92120 34900
rect 92380 34880 92620 34900
rect 92880 34880 93120 34900
rect 93380 34880 93620 34900
rect 93880 34880 94120 34900
rect 94380 34880 94620 34900
rect 94880 34880 95120 34900
rect 95380 34880 95620 34900
rect 95880 34880 96000 34900
rect 92000 34620 92100 34880
rect 92400 34620 92600 34880
rect 92900 34620 93100 34880
rect 93400 34620 93600 34880
rect 93900 34620 94100 34880
rect 94400 34620 94600 34880
rect 94900 34620 95100 34880
rect 95400 34620 95600 34880
rect 95900 34620 96000 34880
rect 92000 34600 92120 34620
rect 92380 34600 92620 34620
rect 92880 34600 93120 34620
rect 93380 34600 93620 34620
rect 93880 34600 94120 34620
rect 94380 34600 94620 34620
rect 94880 34600 95120 34620
rect 95380 34600 95620 34620
rect 95880 34600 96000 34620
rect 92000 34400 96000 34600
rect 92000 34380 92120 34400
rect 92380 34380 92620 34400
rect 92880 34380 93120 34400
rect 93380 34380 93620 34400
rect 93880 34380 94120 34400
rect 94380 34380 94620 34400
rect 94880 34380 95120 34400
rect 95380 34380 95620 34400
rect 95880 34380 96000 34400
rect 92000 34120 92100 34380
rect 92400 34120 92600 34380
rect 92900 34120 93100 34380
rect 93400 34120 93600 34380
rect 93900 34120 94100 34380
rect 94400 34120 94600 34380
rect 94900 34120 95100 34380
rect 95400 34120 95600 34380
rect 95900 34120 96000 34380
rect 92000 34100 92120 34120
rect 92380 34100 92620 34120
rect 92880 34100 93120 34120
rect 93380 34100 93620 34120
rect 93880 34100 94120 34120
rect 94380 34100 94620 34120
rect 94880 34100 95120 34120
rect 95380 34100 95620 34120
rect 95880 34100 96000 34120
rect 92000 33900 96000 34100
rect 92000 33880 92120 33900
rect 92380 33880 92620 33900
rect 92880 33880 93120 33900
rect 93380 33880 93620 33900
rect 93880 33880 94120 33900
rect 94380 33880 94620 33900
rect 94880 33880 95120 33900
rect 95380 33880 95620 33900
rect 95880 33880 96000 33900
rect 92000 33620 92100 33880
rect 92400 33620 92600 33880
rect 92900 33620 93100 33880
rect 93400 33620 93600 33880
rect 93900 33620 94100 33880
rect 94400 33620 94600 33880
rect 94900 33620 95100 33880
rect 95400 33620 95600 33880
rect 95900 33620 96000 33880
rect 92000 33600 92120 33620
rect 92380 33600 92620 33620
rect 92880 33600 93120 33620
rect 93380 33600 93620 33620
rect 93880 33600 94120 33620
rect 94380 33600 94620 33620
rect 94880 33600 95120 33620
rect 95380 33600 95620 33620
rect 95880 33600 96000 33620
rect 92000 33400 96000 33600
rect 92000 33380 92120 33400
rect 92380 33380 92620 33400
rect 92880 33380 93120 33400
rect 93380 33380 93620 33400
rect 93880 33380 94120 33400
rect 94380 33380 94620 33400
rect 94880 33380 95120 33400
rect 95380 33380 95620 33400
rect 95880 33380 96000 33400
rect 92000 33120 92100 33380
rect 92400 33120 92600 33380
rect 92900 33120 93100 33380
rect 93400 33120 93600 33380
rect 93900 33120 94100 33380
rect 94400 33120 94600 33380
rect 94900 33120 95100 33380
rect 95400 33120 95600 33380
rect 95900 33120 96000 33380
rect 92000 33100 92120 33120
rect 92380 33100 92620 33120
rect 92880 33100 93120 33120
rect 93380 33100 93620 33120
rect 93880 33100 94120 33120
rect 94380 33100 94620 33120
rect 94880 33100 95120 33120
rect 95380 33100 95620 33120
rect 95880 33100 96000 33120
rect 92000 32900 96000 33100
rect 92000 32880 92120 32900
rect 92380 32880 92620 32900
rect 92880 32880 93120 32900
rect 93380 32880 93620 32900
rect 93880 32880 94120 32900
rect 94380 32880 94620 32900
rect 94880 32880 95120 32900
rect 95380 32880 95620 32900
rect 95880 32880 96000 32900
rect 92000 32620 92100 32880
rect 92400 32620 92600 32880
rect 92900 32620 93100 32880
rect 93400 32620 93600 32880
rect 93900 32620 94100 32880
rect 94400 32620 94600 32880
rect 94900 32620 95100 32880
rect 95400 32620 95600 32880
rect 95900 32620 96000 32880
rect 92000 32600 92120 32620
rect 92380 32600 92620 32620
rect 92880 32600 93120 32620
rect 93380 32600 93620 32620
rect 93880 32600 94120 32620
rect 94380 32600 94620 32620
rect 94880 32600 95120 32620
rect 95380 32600 95620 32620
rect 95880 32600 96000 32620
rect 92000 32400 96000 32600
rect 92000 32380 92120 32400
rect 92380 32380 92620 32400
rect 92880 32380 93120 32400
rect 93380 32380 93620 32400
rect 93880 32380 94120 32400
rect 94380 32380 94620 32400
rect 94880 32380 95120 32400
rect 95380 32380 95620 32400
rect 95880 32380 96000 32400
rect 92000 32120 92100 32380
rect 92400 32120 92600 32380
rect 92900 32120 93100 32380
rect 93400 32120 93600 32380
rect 93900 32120 94100 32380
rect 94400 32120 94600 32380
rect 94900 32120 95100 32380
rect 95400 32120 95600 32380
rect 95900 32120 96000 32380
rect 92000 32100 92120 32120
rect 92380 32100 92620 32120
rect 92880 32100 93120 32120
rect 93380 32100 93620 32120
rect 93880 32100 94120 32120
rect 94380 32100 94620 32120
rect 94880 32100 95120 32120
rect 95380 32100 95620 32120
rect 95880 32100 96000 32120
rect 92000 31900 96000 32100
rect 92000 31880 92120 31900
rect 92380 31880 92620 31900
rect 92880 31880 93120 31900
rect 93380 31880 93620 31900
rect 93880 31880 94120 31900
rect 94380 31880 94620 31900
rect 94880 31880 95120 31900
rect 95380 31880 95620 31900
rect 95880 31880 96000 31900
rect 92000 31620 92100 31880
rect 92400 31620 92600 31880
rect 92900 31620 93100 31880
rect 93400 31620 93600 31880
rect 93900 31620 94100 31880
rect 94400 31620 94600 31880
rect 94900 31620 95100 31880
rect 95400 31620 95600 31880
rect 95900 31620 96000 31880
rect 92000 31600 92120 31620
rect 92380 31600 92620 31620
rect 92880 31600 93120 31620
rect 93380 31600 93620 31620
rect 93880 31600 94120 31620
rect 94380 31600 94620 31620
rect 94880 31600 95120 31620
rect 95380 31600 95620 31620
rect 95880 31600 96000 31620
rect 92000 31400 96000 31600
rect 92000 31380 92120 31400
rect 92380 31380 92620 31400
rect 92880 31380 93120 31400
rect 93380 31380 93620 31400
rect 93880 31380 94120 31400
rect 94380 31380 94620 31400
rect 94880 31380 95120 31400
rect 95380 31380 95620 31400
rect 95880 31380 96000 31400
rect 92000 31120 92100 31380
rect 92400 31120 92600 31380
rect 92900 31120 93100 31380
rect 93400 31120 93600 31380
rect 93900 31120 94100 31380
rect 94400 31120 94600 31380
rect 94900 31120 95100 31380
rect 95400 31120 95600 31380
rect 95900 31120 96000 31380
rect 92000 31100 92120 31120
rect 92380 31100 92620 31120
rect 92880 31100 93120 31120
rect 93380 31100 93620 31120
rect 93880 31100 94120 31120
rect 94380 31100 94620 31120
rect 94880 31100 95120 31120
rect 95380 31100 95620 31120
rect 95880 31100 96000 31120
rect 92000 30900 96000 31100
rect 92000 30880 92120 30900
rect 92380 30880 92620 30900
rect 92880 30880 93120 30900
rect 93380 30880 93620 30900
rect 93880 30880 94120 30900
rect 94380 30880 94620 30900
rect 94880 30880 95120 30900
rect 95380 30880 95620 30900
rect 95880 30880 96000 30900
rect 92000 30620 92100 30880
rect 92400 30620 92600 30880
rect 92900 30620 93100 30880
rect 93400 30620 93600 30880
rect 93900 30620 94100 30880
rect 94400 30620 94600 30880
rect 94900 30620 95100 30880
rect 95400 30620 95600 30880
rect 95900 30620 96000 30880
rect 92000 30600 92120 30620
rect 92380 30600 92620 30620
rect 92880 30600 93120 30620
rect 93380 30600 93620 30620
rect 93880 30600 94120 30620
rect 94380 30600 94620 30620
rect 94880 30600 95120 30620
rect 95380 30600 95620 30620
rect 95880 30600 96000 30620
rect 92000 30400 96000 30600
rect 92000 30380 92120 30400
rect 92380 30380 92620 30400
rect 92880 30380 93120 30400
rect 93380 30380 93620 30400
rect 93880 30380 94120 30400
rect 94380 30380 94620 30400
rect 94880 30380 95120 30400
rect 95380 30380 95620 30400
rect 95880 30380 96000 30400
rect 92000 30120 92100 30380
rect 92400 30120 92600 30380
rect 92900 30120 93100 30380
rect 93400 30120 93600 30380
rect 93900 30120 94100 30380
rect 94400 30120 94600 30380
rect 94900 30120 95100 30380
rect 95400 30120 95600 30380
rect 95900 30120 96000 30380
rect 92000 30100 92120 30120
rect 92380 30100 92620 30120
rect 92880 30100 93120 30120
rect 93380 30100 93620 30120
rect 93880 30100 94120 30120
rect 94380 30100 94620 30120
rect 94880 30100 95120 30120
rect 95380 30100 95620 30120
rect 95880 30100 96000 30120
rect 92000 29900 96000 30100
rect 92000 29880 92120 29900
rect 92380 29880 92620 29900
rect 92880 29880 93120 29900
rect 93380 29880 93620 29900
rect 93880 29880 94120 29900
rect 94380 29880 94620 29900
rect 94880 29880 95120 29900
rect 95380 29880 95620 29900
rect 95880 29880 96000 29900
rect 92000 29620 92100 29880
rect 92400 29620 92600 29880
rect 92900 29620 93100 29880
rect 93400 29620 93600 29880
rect 93900 29620 94100 29880
rect 94400 29620 94600 29880
rect 94900 29620 95100 29880
rect 95400 29620 95600 29880
rect 95900 29620 96000 29880
rect 92000 29600 92120 29620
rect 92380 29600 92620 29620
rect 92880 29600 93120 29620
rect 93380 29600 93620 29620
rect 93880 29600 94120 29620
rect 94380 29600 94620 29620
rect 94880 29600 95120 29620
rect 95380 29600 95620 29620
rect 95880 29600 96000 29620
rect 92000 29400 96000 29600
rect 92000 29380 92120 29400
rect 92380 29380 92620 29400
rect 92880 29380 93120 29400
rect 93380 29380 93620 29400
rect 93880 29380 94120 29400
rect 94380 29380 94620 29400
rect 94880 29380 95120 29400
rect 95380 29380 95620 29400
rect 95880 29380 96000 29400
rect 92000 29120 92100 29380
rect 92400 29120 92600 29380
rect 92900 29120 93100 29380
rect 93400 29120 93600 29380
rect 93900 29120 94100 29380
rect 94400 29120 94600 29380
rect 94900 29120 95100 29380
rect 95400 29120 95600 29380
rect 95900 29120 96000 29380
rect 92000 29100 92120 29120
rect 92380 29100 92620 29120
rect 92880 29100 93120 29120
rect 93380 29100 93620 29120
rect 93880 29100 94120 29120
rect 94380 29100 94620 29120
rect 94880 29100 95120 29120
rect 95380 29100 95620 29120
rect 95880 29100 96000 29120
rect 92000 28900 96000 29100
rect 92000 28880 92120 28900
rect 92380 28880 92620 28900
rect 92880 28880 93120 28900
rect 93380 28880 93620 28900
rect 93880 28880 94120 28900
rect 94380 28880 94620 28900
rect 94880 28880 95120 28900
rect 95380 28880 95620 28900
rect 95880 28880 96000 28900
rect 92000 28620 92100 28880
rect 92400 28620 92600 28880
rect 92900 28620 93100 28880
rect 93400 28620 93600 28880
rect 93900 28620 94100 28880
rect 94400 28620 94600 28880
rect 94900 28620 95100 28880
rect 95400 28620 95600 28880
rect 95900 28620 96000 28880
rect 92000 28600 92120 28620
rect 92380 28600 92620 28620
rect 92880 28600 93120 28620
rect 93380 28600 93620 28620
rect 93880 28600 94120 28620
rect 94380 28600 94620 28620
rect 94880 28600 95120 28620
rect 95380 28600 95620 28620
rect 95880 28600 96000 28620
rect 92000 28400 96000 28600
rect 92000 28380 92120 28400
rect 92380 28380 92620 28400
rect 92880 28380 93120 28400
rect 93380 28380 93620 28400
rect 93880 28380 94120 28400
rect 94380 28380 94620 28400
rect 94880 28380 95120 28400
rect 95380 28380 95620 28400
rect 95880 28380 96000 28400
rect 92000 28120 92100 28380
rect 92400 28120 92600 28380
rect 92900 28120 93100 28380
rect 93400 28120 93600 28380
rect 93900 28120 94100 28380
rect 94400 28120 94600 28380
rect 94900 28120 95100 28380
rect 95400 28120 95600 28380
rect 95900 28120 96000 28380
rect 92000 28100 92120 28120
rect 92380 28100 92620 28120
rect 92880 28100 93120 28120
rect 93380 28100 93620 28120
rect 93880 28100 94120 28120
rect 94380 28100 94620 28120
rect 94880 28100 95120 28120
rect 95380 28100 95620 28120
rect 95880 28100 96000 28120
rect 92000 28000 96000 28100
rect 88000 27900 96000 28000
rect 88000 27880 88120 27900
rect 88380 27880 88620 27900
rect 88880 27880 89120 27900
rect 89380 27880 89620 27900
rect 89880 27880 90120 27900
rect 90380 27880 90620 27900
rect 90880 27880 91120 27900
rect 91380 27880 91620 27900
rect 91880 27880 92120 27900
rect 92380 27880 92620 27900
rect 92880 27880 93120 27900
rect 93380 27880 93620 27900
rect 93880 27880 94120 27900
rect 94380 27880 94620 27900
rect 94880 27880 95120 27900
rect 95380 27880 95620 27900
rect 95880 27880 96000 27900
rect 88000 27620 88100 27880
rect 88400 27620 88600 27880
rect 88900 27620 89100 27880
rect 89400 27620 89600 27880
rect 89900 27620 90100 27880
rect 90400 27620 90600 27880
rect 90900 27620 91100 27880
rect 91400 27620 91600 27880
rect 91900 27620 92100 27880
rect 92400 27620 92600 27880
rect 92900 27620 93100 27880
rect 93400 27620 93600 27880
rect 93900 27620 94100 27880
rect 94400 27620 94600 27880
rect 94900 27620 95100 27880
rect 95400 27620 95600 27880
rect 95900 27620 96000 27880
rect 88000 27600 88120 27620
rect 88380 27600 88620 27620
rect 88880 27600 89120 27620
rect 89380 27600 89620 27620
rect 89880 27600 90120 27620
rect 90380 27600 90620 27620
rect 90880 27600 91120 27620
rect 91380 27600 91620 27620
rect 91880 27600 92120 27620
rect 92380 27600 92620 27620
rect 92880 27600 93120 27620
rect 93380 27600 93620 27620
rect 93880 27600 94120 27620
rect 94380 27600 94620 27620
rect 94880 27600 95120 27620
rect 95380 27600 95620 27620
rect 95880 27600 96000 27620
rect 88000 27400 96000 27600
rect 88000 27380 88120 27400
rect 88380 27380 88620 27400
rect 88880 27380 89120 27400
rect 89380 27380 89620 27400
rect 89880 27380 90120 27400
rect 90380 27380 90620 27400
rect 90880 27380 91120 27400
rect 91380 27380 91620 27400
rect 91880 27380 92120 27400
rect 92380 27380 92620 27400
rect 92880 27380 93120 27400
rect 93380 27380 93620 27400
rect 93880 27380 94120 27400
rect 94380 27380 94620 27400
rect 94880 27380 95120 27400
rect 95380 27380 95620 27400
rect 95880 27380 96000 27400
rect 88000 27120 88100 27380
rect 88400 27120 88600 27380
rect 88900 27120 89100 27380
rect 89400 27120 89600 27380
rect 89900 27120 90100 27380
rect 90400 27120 90600 27380
rect 90900 27120 91100 27380
rect 91400 27120 91600 27380
rect 91900 27120 92100 27380
rect 92400 27120 92600 27380
rect 92900 27120 93100 27380
rect 93400 27120 93600 27380
rect 93900 27120 94100 27380
rect 94400 27120 94600 27380
rect 94900 27120 95100 27380
rect 95400 27120 95600 27380
rect 95900 27120 96000 27380
rect 88000 27100 88120 27120
rect 88380 27100 88620 27120
rect 88880 27100 89120 27120
rect 89380 27100 89620 27120
rect 89880 27100 90120 27120
rect 90380 27100 90620 27120
rect 90880 27100 91120 27120
rect 91380 27100 91620 27120
rect 91880 27100 92120 27120
rect 92380 27100 92620 27120
rect 92880 27100 93120 27120
rect 93380 27100 93620 27120
rect 93880 27100 94120 27120
rect 94380 27100 94620 27120
rect 94880 27100 95120 27120
rect 95380 27100 95620 27120
rect 95880 27100 96000 27120
rect 88000 26900 96000 27100
rect 88000 26880 88120 26900
rect 88380 26880 88620 26900
rect 88880 26880 89120 26900
rect 89380 26880 89620 26900
rect 89880 26880 90120 26900
rect 90380 26880 90620 26900
rect 90880 26880 91120 26900
rect 91380 26880 91620 26900
rect 91880 26880 92120 26900
rect 92380 26880 92620 26900
rect 92880 26880 93120 26900
rect 93380 26880 93620 26900
rect 93880 26880 94120 26900
rect 94380 26880 94620 26900
rect 94880 26880 95120 26900
rect 95380 26880 95620 26900
rect 95880 26880 96000 26900
rect 88000 26620 88100 26880
rect 88400 26620 88600 26880
rect 88900 26620 89100 26880
rect 89400 26620 89600 26880
rect 89900 26620 90100 26880
rect 90400 26620 90600 26880
rect 90900 26620 91100 26880
rect 91400 26620 91600 26880
rect 91900 26620 92100 26880
rect 92400 26620 92600 26880
rect 92900 26620 93100 26880
rect 93400 26620 93600 26880
rect 93900 26620 94100 26880
rect 94400 26620 94600 26880
rect 94900 26620 95100 26880
rect 95400 26620 95600 26880
rect 95900 26620 96000 26880
rect 88000 26600 88120 26620
rect 88380 26600 88620 26620
rect 88880 26600 89120 26620
rect 89380 26600 89620 26620
rect 89880 26600 90120 26620
rect 90380 26600 90620 26620
rect 90880 26600 91120 26620
rect 91380 26600 91620 26620
rect 91880 26600 92120 26620
rect 92380 26600 92620 26620
rect 92880 26600 93120 26620
rect 93380 26600 93620 26620
rect 93880 26600 94120 26620
rect 94380 26600 94620 26620
rect 94880 26600 95120 26620
rect 95380 26600 95620 26620
rect 95880 26600 96000 26620
rect 88000 26400 96000 26600
rect 88000 26380 88120 26400
rect 88380 26380 88620 26400
rect 88880 26380 89120 26400
rect 89380 26380 89620 26400
rect 89880 26380 90120 26400
rect 90380 26380 90620 26400
rect 90880 26380 91120 26400
rect 91380 26380 91620 26400
rect 91880 26380 92120 26400
rect 92380 26380 92620 26400
rect 92880 26380 93120 26400
rect 93380 26380 93620 26400
rect 93880 26380 94120 26400
rect 94380 26380 94620 26400
rect 94880 26380 95120 26400
rect 95380 26380 95620 26400
rect 95880 26380 96000 26400
rect 88000 26120 88100 26380
rect 88400 26120 88600 26380
rect 88900 26120 89100 26380
rect 89400 26120 89600 26380
rect 89900 26120 90100 26380
rect 90400 26120 90600 26380
rect 90900 26120 91100 26380
rect 91400 26120 91600 26380
rect 91900 26120 92100 26380
rect 92400 26120 92600 26380
rect 92900 26120 93100 26380
rect 93400 26120 93600 26380
rect 93900 26120 94100 26380
rect 94400 26120 94600 26380
rect 94900 26120 95100 26380
rect 95400 26120 95600 26380
rect 95900 26120 96000 26380
rect 88000 26100 88120 26120
rect 88380 26100 88620 26120
rect 88880 26100 89120 26120
rect 89380 26100 89620 26120
rect 89880 26100 90120 26120
rect 90380 26100 90620 26120
rect 90880 26100 91120 26120
rect 91380 26100 91620 26120
rect 91880 26100 92120 26120
rect 92380 26100 92620 26120
rect 92880 26100 93120 26120
rect 93380 26100 93620 26120
rect 93880 26100 94120 26120
rect 94380 26100 94620 26120
rect 94880 26100 95120 26120
rect 95380 26100 95620 26120
rect 95880 26100 96000 26120
rect 88000 26000 96000 26100
rect 88000 25900 100000 26000
rect 88000 25880 88120 25900
rect 88380 25880 88620 25900
rect 88880 25880 89120 25900
rect 89380 25880 89620 25900
rect 89880 25880 90120 25900
rect 90380 25880 90620 25900
rect 90880 25880 91120 25900
rect 91380 25880 91620 25900
rect 91880 25880 92120 25900
rect 92380 25880 92620 25900
rect 92880 25880 93120 25900
rect 93380 25880 93620 25900
rect 93880 25880 94120 25900
rect 94380 25880 94620 25900
rect 94880 25880 95120 25900
rect 95380 25880 95620 25900
rect 95880 25880 96120 25900
rect 96380 25880 96620 25900
rect 96880 25880 97120 25900
rect 97380 25880 97620 25900
rect 97880 25880 98120 25900
rect 98380 25880 98620 25900
rect 98880 25880 99120 25900
rect 99380 25880 99620 25900
rect 99880 25880 100000 25900
rect 88000 25620 88100 25880
rect 88400 25620 88600 25880
rect 88900 25620 89100 25880
rect 89400 25620 89600 25880
rect 89900 25620 90100 25880
rect 90400 25620 90600 25880
rect 90900 25620 91100 25880
rect 91400 25620 91600 25880
rect 91900 25620 92100 25880
rect 92400 25620 92600 25880
rect 92900 25620 93100 25880
rect 93400 25620 93600 25880
rect 93900 25620 94100 25880
rect 94400 25620 94600 25880
rect 94900 25620 95100 25880
rect 95400 25620 95600 25880
rect 95900 25620 96100 25880
rect 96400 25620 96600 25880
rect 96900 25620 97100 25880
rect 97400 25620 97600 25880
rect 97900 25620 98100 25880
rect 98400 25620 98600 25880
rect 98900 25620 99100 25880
rect 99400 25620 99600 25880
rect 99900 25620 100000 25880
rect 88000 25600 88120 25620
rect 88380 25600 88620 25620
rect 88880 25600 89120 25620
rect 89380 25600 89620 25620
rect 89880 25600 90120 25620
rect 90380 25600 90620 25620
rect 90880 25600 91120 25620
rect 91380 25600 91620 25620
rect 91880 25600 92120 25620
rect 92380 25600 92620 25620
rect 92880 25600 93120 25620
rect 93380 25600 93620 25620
rect 93880 25600 94120 25620
rect 94380 25600 94620 25620
rect 94880 25600 95120 25620
rect 95380 25600 95620 25620
rect 95880 25600 96120 25620
rect 96380 25600 96620 25620
rect 96880 25600 97120 25620
rect 97380 25600 97620 25620
rect 97880 25600 98120 25620
rect 98380 25600 98620 25620
rect 98880 25600 99120 25620
rect 99380 25600 99620 25620
rect 99880 25600 100000 25620
rect 88000 25400 100000 25600
rect 88000 25380 88120 25400
rect 88380 25380 88620 25400
rect 88880 25380 89120 25400
rect 89380 25380 89620 25400
rect 89880 25380 90120 25400
rect 90380 25380 90620 25400
rect 90880 25380 91120 25400
rect 91380 25380 91620 25400
rect 91880 25380 92120 25400
rect 92380 25380 92620 25400
rect 92880 25380 93120 25400
rect 93380 25380 93620 25400
rect 93880 25380 94120 25400
rect 94380 25380 94620 25400
rect 94880 25380 95120 25400
rect 95380 25380 95620 25400
rect 95880 25380 96120 25400
rect 96380 25380 96620 25400
rect 96880 25380 97120 25400
rect 97380 25380 97620 25400
rect 97880 25380 98120 25400
rect 98380 25380 98620 25400
rect 98880 25380 99120 25400
rect 99380 25380 99620 25400
rect 99880 25380 100000 25400
rect 88000 25120 88100 25380
rect 88400 25120 88600 25380
rect 88900 25120 89100 25380
rect 89400 25120 89600 25380
rect 89900 25120 90100 25380
rect 90400 25120 90600 25380
rect 90900 25120 91100 25380
rect 91400 25120 91600 25380
rect 91900 25120 92100 25380
rect 92400 25120 92600 25380
rect 92900 25120 93100 25380
rect 93400 25120 93600 25380
rect 93900 25120 94100 25380
rect 94400 25120 94600 25380
rect 94900 25120 95100 25380
rect 95400 25120 95600 25380
rect 95900 25120 96100 25380
rect 96400 25120 96600 25380
rect 96900 25120 97100 25380
rect 97400 25120 97600 25380
rect 97900 25120 98100 25380
rect 98400 25120 98600 25380
rect 98900 25120 99100 25380
rect 99400 25120 99600 25380
rect 99900 25120 100000 25380
rect 88000 25100 88120 25120
rect 88380 25100 88620 25120
rect 88880 25100 89120 25120
rect 89380 25100 89620 25120
rect 89880 25100 90120 25120
rect 90380 25100 90620 25120
rect 90880 25100 91120 25120
rect 91380 25100 91620 25120
rect 91880 25100 92120 25120
rect 92380 25100 92620 25120
rect 92880 25100 93120 25120
rect 93380 25100 93620 25120
rect 93880 25100 94120 25120
rect 94380 25100 94620 25120
rect 94880 25100 95120 25120
rect 95380 25100 95620 25120
rect 95880 25100 96120 25120
rect 96380 25100 96620 25120
rect 96880 25100 97120 25120
rect 97380 25100 97620 25120
rect 97880 25100 98120 25120
rect 98380 25100 98620 25120
rect 98880 25100 99120 25120
rect 99380 25100 99620 25120
rect 99880 25100 100000 25120
rect 88000 24900 100000 25100
rect 88000 24880 88120 24900
rect 88380 24880 88620 24900
rect 88880 24880 89120 24900
rect 89380 24880 89620 24900
rect 89880 24880 90120 24900
rect 90380 24880 90620 24900
rect 90880 24880 91120 24900
rect 91380 24880 91620 24900
rect 91880 24880 92120 24900
rect 92380 24880 92620 24900
rect 92880 24880 93120 24900
rect 93380 24880 93620 24900
rect 93880 24880 94120 24900
rect 94380 24880 94620 24900
rect 94880 24880 95120 24900
rect 95380 24880 95620 24900
rect 95880 24880 96120 24900
rect 96380 24880 96620 24900
rect 96880 24880 97120 24900
rect 97380 24880 97620 24900
rect 97880 24880 98120 24900
rect 98380 24880 98620 24900
rect 98880 24880 99120 24900
rect 99380 24880 99620 24900
rect 99880 24880 100000 24900
rect 88000 24620 88100 24880
rect 88400 24620 88600 24880
rect 88900 24620 89100 24880
rect 89400 24620 89600 24880
rect 89900 24620 90100 24880
rect 90400 24620 90600 24880
rect 90900 24620 91100 24880
rect 91400 24620 91600 24880
rect 91900 24620 92100 24880
rect 92400 24620 92600 24880
rect 92900 24620 93100 24880
rect 93400 24620 93600 24880
rect 93900 24620 94100 24880
rect 94400 24620 94600 24880
rect 94900 24620 95100 24880
rect 95400 24620 95600 24880
rect 95900 24620 96100 24880
rect 96400 24620 96600 24880
rect 96900 24620 97100 24880
rect 97400 24620 97600 24880
rect 97900 24620 98100 24880
rect 98400 24620 98600 24880
rect 98900 24620 99100 24880
rect 99400 24620 99600 24880
rect 99900 24620 100000 24880
rect 88000 24600 88120 24620
rect 88380 24600 88620 24620
rect 88880 24600 89120 24620
rect 89380 24600 89620 24620
rect 89880 24600 90120 24620
rect 90380 24600 90620 24620
rect 90880 24600 91120 24620
rect 91380 24600 91620 24620
rect 91880 24600 92120 24620
rect 92380 24600 92620 24620
rect 92880 24600 93120 24620
rect 93380 24600 93620 24620
rect 93880 24600 94120 24620
rect 94380 24600 94620 24620
rect 94880 24600 95120 24620
rect 95380 24600 95620 24620
rect 95880 24600 96120 24620
rect 96380 24600 96620 24620
rect 96880 24600 97120 24620
rect 97380 24600 97620 24620
rect 97880 24600 98120 24620
rect 98380 24600 98620 24620
rect 98880 24600 99120 24620
rect 99380 24600 99620 24620
rect 99880 24600 100000 24620
rect 88000 24400 100000 24600
rect 88000 24380 88120 24400
rect 88380 24380 88620 24400
rect 88880 24380 89120 24400
rect 89380 24380 89620 24400
rect 89880 24380 90120 24400
rect 90380 24380 90620 24400
rect 90880 24380 91120 24400
rect 91380 24380 91620 24400
rect 91880 24380 92120 24400
rect 92380 24380 92620 24400
rect 92880 24380 93120 24400
rect 93380 24380 93620 24400
rect 93880 24380 94120 24400
rect 94380 24380 94620 24400
rect 94880 24380 95120 24400
rect 95380 24380 95620 24400
rect 95880 24380 96120 24400
rect 96380 24380 96620 24400
rect 96880 24380 97120 24400
rect 97380 24380 97620 24400
rect 97880 24380 98120 24400
rect 98380 24380 98620 24400
rect 98880 24380 99120 24400
rect 99380 24380 99620 24400
rect 99880 24380 100000 24400
rect 88000 24120 88100 24380
rect 88400 24120 88600 24380
rect 88900 24120 89100 24380
rect 89400 24120 89600 24380
rect 89900 24120 90100 24380
rect 90400 24120 90600 24380
rect 90900 24120 91100 24380
rect 91400 24120 91600 24380
rect 91900 24120 92100 24380
rect 92400 24120 92600 24380
rect 92900 24120 93100 24380
rect 93400 24120 93600 24380
rect 93900 24120 94100 24380
rect 94400 24120 94600 24380
rect 94900 24120 95100 24380
rect 95400 24120 95600 24380
rect 95900 24120 96100 24380
rect 96400 24120 96600 24380
rect 96900 24120 97100 24380
rect 97400 24120 97600 24380
rect 97900 24120 98100 24380
rect 98400 24120 98600 24380
rect 98900 24120 99100 24380
rect 99400 24120 99600 24380
rect 99900 24120 100000 24380
rect 88000 24100 88120 24120
rect 88380 24100 88620 24120
rect 88880 24100 89120 24120
rect 89380 24100 89620 24120
rect 89880 24100 90120 24120
rect 90380 24100 90620 24120
rect 90880 24100 91120 24120
rect 91380 24100 91620 24120
rect 91880 24100 92120 24120
rect 92380 24100 92620 24120
rect 92880 24100 93120 24120
rect 93380 24100 93620 24120
rect 93880 24100 94120 24120
rect 94380 24100 94620 24120
rect 94880 24100 95120 24120
rect 95380 24100 95620 24120
rect 95880 24100 96120 24120
rect 96380 24100 96620 24120
rect 96880 24100 97120 24120
rect 97380 24100 97620 24120
rect 97880 24100 98120 24120
rect 98380 24100 98620 24120
rect 98880 24100 99120 24120
rect 99380 24100 99620 24120
rect 99880 24100 100000 24120
rect 88000 24000 100000 24100
rect 96000 23900 100000 24000
rect 96000 23880 96120 23900
rect 96380 23880 96620 23900
rect 96880 23880 97120 23900
rect 97380 23880 97620 23900
rect 97880 23880 98120 23900
rect 98380 23880 98620 23900
rect 98880 23880 99120 23900
rect 99380 23880 99620 23900
rect 99880 23880 100000 23900
rect 96000 23620 96100 23880
rect 96400 23620 96600 23880
rect 96900 23620 97100 23880
rect 97400 23620 97600 23880
rect 97900 23620 98100 23880
rect 98400 23620 98600 23880
rect 98900 23620 99100 23880
rect 99400 23620 99600 23880
rect 99900 23620 100000 23880
rect 96000 23600 96120 23620
rect 96380 23600 96620 23620
rect 96880 23600 97120 23620
rect 97380 23600 97620 23620
rect 97880 23600 98120 23620
rect 98380 23600 98620 23620
rect 98880 23600 99120 23620
rect 99380 23600 99620 23620
rect 99880 23600 100000 23620
rect 96000 23400 100000 23600
rect 96000 23380 96120 23400
rect 96380 23380 96620 23400
rect 96880 23380 97120 23400
rect 97380 23380 97620 23400
rect 97880 23380 98120 23400
rect 98380 23380 98620 23400
rect 98880 23380 99120 23400
rect 99380 23380 99620 23400
rect 99880 23380 100000 23400
rect 96000 23120 96100 23380
rect 96400 23120 96600 23380
rect 96900 23120 97100 23380
rect 97400 23120 97600 23380
rect 97900 23120 98100 23380
rect 98400 23120 98600 23380
rect 98900 23120 99100 23380
rect 99400 23120 99600 23380
rect 99900 23120 100000 23380
rect 96000 23100 96120 23120
rect 96380 23100 96620 23120
rect 96880 23100 97120 23120
rect 97380 23100 97620 23120
rect 97880 23100 98120 23120
rect 98380 23100 98620 23120
rect 98880 23100 99120 23120
rect 99380 23100 99620 23120
rect 99880 23100 100000 23120
rect 96000 22900 100000 23100
rect 96000 22880 96120 22900
rect 96380 22880 96620 22900
rect 96880 22880 97120 22900
rect 97380 22880 97620 22900
rect 97880 22880 98120 22900
rect 98380 22880 98620 22900
rect 98880 22880 99120 22900
rect 99380 22880 99620 22900
rect 99880 22880 100000 22900
rect 96000 22620 96100 22880
rect 96400 22620 96600 22880
rect 96900 22620 97100 22880
rect 97400 22620 97600 22880
rect 97900 22620 98100 22880
rect 98400 22620 98600 22880
rect 98900 22620 99100 22880
rect 99400 22620 99600 22880
rect 99900 22620 100000 22880
rect 96000 22600 96120 22620
rect 96380 22600 96620 22620
rect 96880 22600 97120 22620
rect 97380 22600 97620 22620
rect 97880 22600 98120 22620
rect 98380 22600 98620 22620
rect 98880 22600 99120 22620
rect 99380 22600 99620 22620
rect 99880 22600 100000 22620
rect 96000 22400 100000 22600
rect 96000 22380 96120 22400
rect 96380 22380 96620 22400
rect 96880 22380 97120 22400
rect 97380 22380 97620 22400
rect 97880 22380 98120 22400
rect 98380 22380 98620 22400
rect 98880 22380 99120 22400
rect 99380 22380 99620 22400
rect 99880 22380 100000 22400
rect 96000 22120 96100 22380
rect 96400 22120 96600 22380
rect 96900 22120 97100 22380
rect 97400 22120 97600 22380
rect 97900 22120 98100 22380
rect 98400 22120 98600 22380
rect 98900 22120 99100 22380
rect 99400 22120 99600 22380
rect 99900 22120 100000 22380
rect 96000 22100 96120 22120
rect 96380 22100 96620 22120
rect 96880 22100 97120 22120
rect 97380 22100 97620 22120
rect 97880 22100 98120 22120
rect 98380 22100 98620 22120
rect 98880 22100 99120 22120
rect 99380 22100 99620 22120
rect 99880 22100 100000 22120
rect 96000 22000 100000 22100
rect 104000 13900 127000 14000
rect 104000 13880 104120 13900
rect 104380 13880 104620 13900
rect 104880 13880 105120 13900
rect 105380 13880 105620 13900
rect 105880 13880 106120 13900
rect 106380 13880 106620 13900
rect 106880 13880 107120 13900
rect 107380 13880 107620 13900
rect 107880 13880 108120 13900
rect 108380 13880 108620 13900
rect 108880 13880 109120 13900
rect 109380 13880 109620 13900
rect 109880 13880 110120 13900
rect 110380 13880 110620 13900
rect 110880 13880 111120 13900
rect 111380 13880 111620 13900
rect 111880 13880 112120 13900
rect 112380 13880 112620 13900
rect 112880 13880 113120 13900
rect 113380 13880 113620 13900
rect 113880 13880 114120 13900
rect 114380 13880 114620 13900
rect 114880 13880 115120 13900
rect 115380 13880 115620 13900
rect 115880 13880 116120 13900
rect 116380 13880 116620 13900
rect 116880 13880 117120 13900
rect 117380 13880 117620 13900
rect 117880 13880 118120 13900
rect 118380 13880 118620 13900
rect 118880 13880 119120 13900
rect 119380 13880 119620 13900
rect 119880 13880 120120 13900
rect 120380 13880 120620 13900
rect 120880 13880 121120 13900
rect 121380 13880 121620 13900
rect 121880 13880 122120 13900
rect 122380 13880 122620 13900
rect 122880 13880 123120 13900
rect 123380 13880 123620 13900
rect 123880 13880 124120 13900
rect 124380 13880 124620 13900
rect 124880 13880 125120 13900
rect 125380 13880 125620 13900
rect 125880 13880 126120 13900
rect 126380 13880 126620 13900
rect 126880 13880 127000 13900
rect 104000 13620 104100 13880
rect 104400 13620 104600 13880
rect 104900 13620 105100 13880
rect 105400 13620 105600 13880
rect 105900 13620 106100 13880
rect 106400 13620 106600 13880
rect 106900 13620 107100 13880
rect 107400 13620 107600 13880
rect 107900 13620 108100 13880
rect 108400 13620 108600 13880
rect 108900 13620 109100 13880
rect 109400 13620 109600 13880
rect 109900 13620 110100 13880
rect 110400 13620 110600 13880
rect 110900 13620 111100 13880
rect 111400 13620 111600 13880
rect 111900 13620 112100 13880
rect 112400 13620 112600 13880
rect 112900 13620 113100 13880
rect 113400 13620 113600 13880
rect 113900 13620 114100 13880
rect 114400 13620 114600 13880
rect 114900 13620 115100 13880
rect 115400 13620 115600 13880
rect 115900 13620 116100 13880
rect 116400 13620 116600 13880
rect 116900 13620 117100 13880
rect 117400 13620 117600 13880
rect 117900 13620 118100 13880
rect 118400 13620 118600 13880
rect 118900 13620 119100 13880
rect 119400 13620 119600 13880
rect 119900 13620 120100 13880
rect 120400 13620 120600 13880
rect 120900 13620 121100 13880
rect 121400 13620 121600 13880
rect 121900 13620 122100 13880
rect 122400 13620 122600 13880
rect 122900 13620 123100 13880
rect 123400 13620 123600 13880
rect 123900 13620 124100 13880
rect 124400 13620 124600 13880
rect 124900 13620 125100 13880
rect 125400 13620 125600 13880
rect 125900 13620 126100 13880
rect 126400 13620 126600 13880
rect 126900 13620 127000 13880
rect 104000 13600 104120 13620
rect 104380 13600 104620 13620
rect 104880 13600 105120 13620
rect 105380 13600 105620 13620
rect 105880 13600 106120 13620
rect 106380 13600 106620 13620
rect 106880 13600 107120 13620
rect 107380 13600 107620 13620
rect 107880 13600 108120 13620
rect 108380 13600 108620 13620
rect 108880 13600 109120 13620
rect 109380 13600 109620 13620
rect 109880 13600 110120 13620
rect 110380 13600 110620 13620
rect 110880 13600 111120 13620
rect 111380 13600 111620 13620
rect 111880 13600 112120 13620
rect 112380 13600 112620 13620
rect 112880 13600 113120 13620
rect 113380 13600 113620 13620
rect 113880 13600 114120 13620
rect 114380 13600 114620 13620
rect 114880 13600 115120 13620
rect 115380 13600 115620 13620
rect 115880 13600 116120 13620
rect 116380 13600 116620 13620
rect 116880 13600 117120 13620
rect 117380 13600 117620 13620
rect 117880 13600 118120 13620
rect 118380 13600 118620 13620
rect 118880 13600 119120 13620
rect 119380 13600 119620 13620
rect 119880 13600 120120 13620
rect 120380 13600 120620 13620
rect 120880 13600 121120 13620
rect 121380 13600 121620 13620
rect 121880 13600 122120 13620
rect 122380 13600 122620 13620
rect 122880 13600 123120 13620
rect 123380 13600 123620 13620
rect 123880 13600 124120 13620
rect 124380 13600 124620 13620
rect 124880 13600 125120 13620
rect 125380 13600 125620 13620
rect 125880 13600 126120 13620
rect 126380 13600 126620 13620
rect 126880 13600 127000 13620
rect 104000 13400 127000 13600
rect 104000 13380 104120 13400
rect 104380 13380 104620 13400
rect 104880 13380 105120 13400
rect 105380 13380 105620 13400
rect 105880 13380 106120 13400
rect 106380 13380 106620 13400
rect 106880 13380 107120 13400
rect 107380 13380 107620 13400
rect 107880 13380 108120 13400
rect 108380 13380 108620 13400
rect 108880 13380 109120 13400
rect 109380 13380 109620 13400
rect 109880 13380 110120 13400
rect 110380 13380 110620 13400
rect 110880 13380 111120 13400
rect 111380 13380 111620 13400
rect 111880 13380 112120 13400
rect 112380 13380 112620 13400
rect 112880 13380 113120 13400
rect 113380 13380 113620 13400
rect 113880 13380 114120 13400
rect 114380 13380 114620 13400
rect 114880 13380 115120 13400
rect 115380 13380 115620 13400
rect 115880 13380 116120 13400
rect 116380 13380 116620 13400
rect 116880 13380 117120 13400
rect 117380 13380 117620 13400
rect 117880 13380 118120 13400
rect 118380 13380 118620 13400
rect 118880 13380 119120 13400
rect 119380 13380 119620 13400
rect 119880 13380 120120 13400
rect 120380 13380 120620 13400
rect 120880 13380 121120 13400
rect 121380 13380 121620 13400
rect 121880 13380 122120 13400
rect 122380 13380 122620 13400
rect 122880 13380 123120 13400
rect 123380 13380 123620 13400
rect 123880 13380 124120 13400
rect 124380 13380 124620 13400
rect 124880 13380 125120 13400
rect 125380 13380 125620 13400
rect 125880 13380 126120 13400
rect 126380 13380 126620 13400
rect 126880 13380 127000 13400
rect 104000 13120 104100 13380
rect 104400 13120 104600 13380
rect 104900 13120 105100 13380
rect 105400 13120 105600 13380
rect 105900 13120 106100 13380
rect 106400 13120 106600 13380
rect 106900 13120 107100 13380
rect 107400 13120 107600 13380
rect 107900 13120 108100 13380
rect 108400 13120 108600 13380
rect 108900 13120 109100 13380
rect 109400 13120 109600 13380
rect 109900 13120 110100 13380
rect 110400 13120 110600 13380
rect 110900 13120 111100 13380
rect 111400 13120 111600 13380
rect 111900 13120 112100 13380
rect 112400 13120 112600 13380
rect 112900 13120 113100 13380
rect 113400 13120 113600 13380
rect 113900 13120 114100 13380
rect 114400 13120 114600 13380
rect 114900 13120 115100 13380
rect 115400 13120 115600 13380
rect 115900 13120 116100 13380
rect 116400 13120 116600 13380
rect 116900 13120 117100 13380
rect 117400 13120 117600 13380
rect 117900 13120 118100 13380
rect 118400 13120 118600 13380
rect 118900 13120 119100 13380
rect 119400 13120 119600 13380
rect 119900 13120 120100 13380
rect 120400 13120 120600 13380
rect 120900 13120 121100 13380
rect 121400 13120 121600 13380
rect 121900 13120 122100 13380
rect 122400 13120 122600 13380
rect 122900 13120 123100 13380
rect 123400 13120 123600 13380
rect 123900 13120 124100 13380
rect 124400 13120 124600 13380
rect 124900 13120 125100 13380
rect 125400 13120 125600 13380
rect 125900 13120 126100 13380
rect 126400 13120 126600 13380
rect 126900 13120 127000 13380
rect 104000 13100 104120 13120
rect 104380 13100 104620 13120
rect 104880 13100 105120 13120
rect 105380 13100 105620 13120
rect 105880 13100 106120 13120
rect 106380 13100 106620 13120
rect 106880 13100 107120 13120
rect 107380 13100 107620 13120
rect 107880 13100 108120 13120
rect 108380 13100 108620 13120
rect 108880 13100 109120 13120
rect 109380 13100 109620 13120
rect 109880 13100 110120 13120
rect 110380 13100 110620 13120
rect 110880 13100 111120 13120
rect 111380 13100 111620 13120
rect 111880 13100 112120 13120
rect 112380 13100 112620 13120
rect 112880 13100 113120 13120
rect 113380 13100 113620 13120
rect 113880 13100 114120 13120
rect 114380 13100 114620 13120
rect 114880 13100 115120 13120
rect 115380 13100 115620 13120
rect 115880 13100 116120 13120
rect 116380 13100 116620 13120
rect 116880 13100 117120 13120
rect 117380 13100 117620 13120
rect 117880 13100 118120 13120
rect 118380 13100 118620 13120
rect 118880 13100 119120 13120
rect 119380 13100 119620 13120
rect 119880 13100 120120 13120
rect 120380 13100 120620 13120
rect 120880 13100 121120 13120
rect 121380 13100 121620 13120
rect 121880 13100 122120 13120
rect 122380 13100 122620 13120
rect 122880 13100 123120 13120
rect 123380 13100 123620 13120
rect 123880 13100 124120 13120
rect 124380 13100 124620 13120
rect 124880 13100 125120 13120
rect 125380 13100 125620 13120
rect 125880 13100 126120 13120
rect 126380 13100 126620 13120
rect 126880 13100 127000 13120
rect 104000 12900 127000 13100
rect 104000 12880 104120 12900
rect 104380 12880 104620 12900
rect 104880 12880 105120 12900
rect 105380 12880 105620 12900
rect 105880 12880 106120 12900
rect 106380 12880 106620 12900
rect 106880 12880 107120 12900
rect 107380 12880 107620 12900
rect 107880 12880 108120 12900
rect 108380 12880 108620 12900
rect 108880 12880 109120 12900
rect 109380 12880 109620 12900
rect 109880 12880 110120 12900
rect 110380 12880 110620 12900
rect 110880 12880 111120 12900
rect 111380 12880 111620 12900
rect 111880 12880 112120 12900
rect 112380 12880 112620 12900
rect 112880 12880 113120 12900
rect 113380 12880 113620 12900
rect 113880 12880 114120 12900
rect 114380 12880 114620 12900
rect 114880 12880 115120 12900
rect 115380 12880 115620 12900
rect 115880 12880 116120 12900
rect 116380 12880 116620 12900
rect 116880 12880 117120 12900
rect 117380 12880 117620 12900
rect 117880 12880 118120 12900
rect 118380 12880 118620 12900
rect 118880 12880 119120 12900
rect 119380 12880 119620 12900
rect 119880 12880 120120 12900
rect 120380 12880 120620 12900
rect 120880 12880 121120 12900
rect 121380 12880 121620 12900
rect 121880 12880 122120 12900
rect 122380 12880 122620 12900
rect 122880 12880 123120 12900
rect 123380 12880 123620 12900
rect 123880 12880 124120 12900
rect 124380 12880 124620 12900
rect 124880 12880 125120 12900
rect 125380 12880 125620 12900
rect 125880 12880 126120 12900
rect 126380 12880 126620 12900
rect 126880 12880 127000 12900
rect 104000 12620 104100 12880
rect 104400 12620 104600 12880
rect 104900 12620 105100 12880
rect 105400 12620 105600 12880
rect 105900 12620 106100 12880
rect 106400 12620 106600 12880
rect 106900 12620 107100 12880
rect 107400 12620 107600 12880
rect 107900 12620 108100 12880
rect 108400 12620 108600 12880
rect 108900 12620 109100 12880
rect 109400 12620 109600 12880
rect 109900 12620 110100 12880
rect 110400 12620 110600 12880
rect 110900 12620 111100 12880
rect 111400 12620 111600 12880
rect 111900 12620 112100 12880
rect 112400 12620 112600 12880
rect 112900 12620 113100 12880
rect 113400 12620 113600 12880
rect 113900 12620 114100 12880
rect 114400 12620 114600 12880
rect 114900 12620 115100 12880
rect 115400 12620 115600 12880
rect 115900 12620 116100 12880
rect 116400 12620 116600 12880
rect 116900 12620 117100 12880
rect 117400 12620 117600 12880
rect 117900 12620 118100 12880
rect 118400 12620 118600 12880
rect 118900 12620 119100 12880
rect 119400 12620 119600 12880
rect 119900 12620 120100 12880
rect 120400 12620 120600 12880
rect 120900 12620 121100 12880
rect 121400 12620 121600 12880
rect 121900 12620 122100 12880
rect 122400 12620 122600 12880
rect 122900 12620 123100 12880
rect 123400 12620 123600 12880
rect 123900 12620 124100 12880
rect 124400 12620 124600 12880
rect 124900 12620 125100 12880
rect 125400 12620 125600 12880
rect 125900 12620 126100 12880
rect 126400 12620 126600 12880
rect 126900 12620 127000 12880
rect 104000 12600 104120 12620
rect 104380 12600 104620 12620
rect 104880 12600 105120 12620
rect 105380 12600 105620 12620
rect 105880 12600 106120 12620
rect 106380 12600 106620 12620
rect 106880 12600 107120 12620
rect 107380 12600 107620 12620
rect 107880 12600 108120 12620
rect 108380 12600 108620 12620
rect 108880 12600 109120 12620
rect 109380 12600 109620 12620
rect 109880 12600 110120 12620
rect 110380 12600 110620 12620
rect 110880 12600 111120 12620
rect 111380 12600 111620 12620
rect 111880 12600 112120 12620
rect 112380 12600 112620 12620
rect 112880 12600 113120 12620
rect 113380 12600 113620 12620
rect 113880 12600 114120 12620
rect 114380 12600 114620 12620
rect 114880 12600 115120 12620
rect 115380 12600 115620 12620
rect 115880 12600 116120 12620
rect 116380 12600 116620 12620
rect 116880 12600 117120 12620
rect 117380 12600 117620 12620
rect 117880 12600 118120 12620
rect 118380 12600 118620 12620
rect 118880 12600 119120 12620
rect 119380 12600 119620 12620
rect 119880 12600 120120 12620
rect 120380 12600 120620 12620
rect 120880 12600 121120 12620
rect 121380 12600 121620 12620
rect 121880 12600 122120 12620
rect 122380 12600 122620 12620
rect 122880 12600 123120 12620
rect 123380 12600 123620 12620
rect 123880 12600 124120 12620
rect 124380 12600 124620 12620
rect 124880 12600 125120 12620
rect 125380 12600 125620 12620
rect 125880 12600 126120 12620
rect 126380 12600 126620 12620
rect 126880 12600 127000 12620
rect 104000 12400 127000 12600
rect 104000 12380 104120 12400
rect 104380 12380 104620 12400
rect 104880 12380 105120 12400
rect 105380 12380 105620 12400
rect 105880 12380 106120 12400
rect 106380 12380 106620 12400
rect 106880 12380 107120 12400
rect 107380 12380 107620 12400
rect 107880 12380 108120 12400
rect 108380 12380 108620 12400
rect 108880 12380 109120 12400
rect 109380 12380 109620 12400
rect 109880 12380 110120 12400
rect 110380 12380 110620 12400
rect 110880 12380 111120 12400
rect 111380 12380 111620 12400
rect 111880 12380 112120 12400
rect 112380 12380 112620 12400
rect 112880 12380 113120 12400
rect 113380 12380 113620 12400
rect 113880 12380 114120 12400
rect 114380 12380 114620 12400
rect 114880 12380 115120 12400
rect 115380 12380 115620 12400
rect 115880 12380 116120 12400
rect 116380 12380 116620 12400
rect 116880 12380 117120 12400
rect 117380 12380 117620 12400
rect 117880 12380 118120 12400
rect 118380 12380 118620 12400
rect 118880 12380 119120 12400
rect 119380 12380 119620 12400
rect 119880 12380 120120 12400
rect 120380 12380 120620 12400
rect 120880 12380 121120 12400
rect 121380 12380 121620 12400
rect 121880 12380 122120 12400
rect 122380 12380 122620 12400
rect 122880 12380 123120 12400
rect 123380 12380 123620 12400
rect 123880 12380 124120 12400
rect 124380 12380 124620 12400
rect 124880 12380 125120 12400
rect 125380 12380 125620 12400
rect 125880 12380 126120 12400
rect 126380 12380 126620 12400
rect 126880 12380 127000 12400
rect 104000 12120 104100 12380
rect 104400 12120 104600 12380
rect 104900 12120 105100 12380
rect 105400 12120 105600 12380
rect 105900 12120 106100 12380
rect 106400 12120 106600 12380
rect 106900 12120 107100 12380
rect 107400 12120 107600 12380
rect 107900 12120 108100 12380
rect 108400 12120 108600 12380
rect 108900 12120 109100 12380
rect 109400 12120 109600 12380
rect 109900 12120 110100 12380
rect 110400 12120 110600 12380
rect 110900 12120 111100 12380
rect 111400 12120 111600 12380
rect 111900 12120 112100 12380
rect 112400 12120 112600 12380
rect 112900 12120 113100 12380
rect 113400 12120 113600 12380
rect 113900 12120 114100 12380
rect 114400 12120 114600 12380
rect 114900 12120 115100 12380
rect 115400 12120 115600 12380
rect 115900 12120 116100 12380
rect 116400 12120 116600 12380
rect 116900 12120 117100 12380
rect 117400 12120 117600 12380
rect 117900 12120 118100 12380
rect 118400 12120 118600 12380
rect 118900 12120 119100 12380
rect 119400 12120 119600 12380
rect 119900 12120 120100 12380
rect 120400 12120 120600 12380
rect 120900 12120 121100 12380
rect 121400 12120 121600 12380
rect 121900 12120 122100 12380
rect 122400 12120 122600 12380
rect 122900 12120 123100 12380
rect 123400 12120 123600 12380
rect 123900 12120 124100 12380
rect 124400 12120 124600 12380
rect 124900 12120 125100 12380
rect 125400 12120 125600 12380
rect 125900 12120 126100 12380
rect 126400 12120 126600 12380
rect 126900 12120 127000 12380
rect 104000 12100 104120 12120
rect 104380 12100 104620 12120
rect 104880 12100 105120 12120
rect 105380 12100 105620 12120
rect 105880 12100 106120 12120
rect 106380 12100 106620 12120
rect 106880 12100 107120 12120
rect 107380 12100 107620 12120
rect 107880 12100 108120 12120
rect 108380 12100 108620 12120
rect 108880 12100 109120 12120
rect 109380 12100 109620 12120
rect 109880 12100 110120 12120
rect 110380 12100 110620 12120
rect 110880 12100 111120 12120
rect 111380 12100 111620 12120
rect 111880 12100 112120 12120
rect 112380 12100 112620 12120
rect 112880 12100 113120 12120
rect 113380 12100 113620 12120
rect 113880 12100 114120 12120
rect 114380 12100 114620 12120
rect 114880 12100 115120 12120
rect 115380 12100 115620 12120
rect 115880 12100 116120 12120
rect 116380 12100 116620 12120
rect 116880 12100 117120 12120
rect 117380 12100 117620 12120
rect 117880 12100 118120 12120
rect 118380 12100 118620 12120
rect 118880 12100 119120 12120
rect 119380 12100 119620 12120
rect 119880 12100 120120 12120
rect 120380 12100 120620 12120
rect 120880 12100 121120 12120
rect 121380 12100 121620 12120
rect 121880 12100 122120 12120
rect 122380 12100 122620 12120
rect 122880 12100 123120 12120
rect 123380 12100 123620 12120
rect 123880 12100 124120 12120
rect 124380 12100 124620 12120
rect 124880 12100 125120 12120
rect 125380 12100 125620 12120
rect 125880 12100 126120 12120
rect 126380 12100 126620 12120
rect 126880 12100 127000 12120
rect 104000 11900 127000 12100
rect 104000 11880 104120 11900
rect 104380 11880 104620 11900
rect 104880 11880 105120 11900
rect 105380 11880 105620 11900
rect 105880 11880 106120 11900
rect 106380 11880 106620 11900
rect 106880 11880 107120 11900
rect 107380 11880 107620 11900
rect 107880 11880 108120 11900
rect 108380 11880 108620 11900
rect 108880 11880 109120 11900
rect 109380 11880 109620 11900
rect 109880 11880 110120 11900
rect 110380 11880 110620 11900
rect 110880 11880 111120 11900
rect 111380 11880 111620 11900
rect 111880 11880 112120 11900
rect 112380 11880 112620 11900
rect 112880 11880 113120 11900
rect 113380 11880 113620 11900
rect 113880 11880 114120 11900
rect 114380 11880 114620 11900
rect 114880 11880 115120 11900
rect 115380 11880 115620 11900
rect 115880 11880 116120 11900
rect 116380 11880 116620 11900
rect 116880 11880 117120 11900
rect 117380 11880 117620 11900
rect 117880 11880 118120 11900
rect 118380 11880 118620 11900
rect 118880 11880 119120 11900
rect 119380 11880 119620 11900
rect 119880 11880 120120 11900
rect 120380 11880 120620 11900
rect 120880 11880 121120 11900
rect 121380 11880 121620 11900
rect 121880 11880 122120 11900
rect 122380 11880 122620 11900
rect 122880 11880 123120 11900
rect 123380 11880 123620 11900
rect 123880 11880 124120 11900
rect 124380 11880 124620 11900
rect 124880 11880 125120 11900
rect 125380 11880 125620 11900
rect 125880 11880 126120 11900
rect 126380 11880 126620 11900
rect 126880 11880 127000 11900
rect 104000 11620 104100 11880
rect 104400 11620 104600 11880
rect 104900 11620 105100 11880
rect 105400 11620 105600 11880
rect 105900 11620 106100 11880
rect 106400 11620 106600 11880
rect 106900 11620 107100 11880
rect 107400 11620 107600 11880
rect 107900 11620 108100 11880
rect 108400 11620 108600 11880
rect 108900 11620 109100 11880
rect 109400 11620 109600 11880
rect 109900 11620 110100 11880
rect 110400 11620 110600 11880
rect 110900 11620 111100 11880
rect 111400 11620 111600 11880
rect 111900 11620 112100 11880
rect 112400 11620 112600 11880
rect 112900 11620 113100 11880
rect 113400 11620 113600 11880
rect 113900 11620 114100 11880
rect 114400 11620 114600 11880
rect 114900 11620 115100 11880
rect 115400 11620 115600 11880
rect 115900 11620 116100 11880
rect 116400 11620 116600 11880
rect 116900 11620 117100 11880
rect 117400 11620 117600 11880
rect 117900 11620 118100 11880
rect 118400 11620 118600 11880
rect 118900 11620 119100 11880
rect 119400 11620 119600 11880
rect 119900 11620 120100 11880
rect 120400 11620 120600 11880
rect 120900 11620 121100 11880
rect 121400 11620 121600 11880
rect 121900 11620 122100 11880
rect 122400 11620 122600 11880
rect 122900 11620 123100 11880
rect 123400 11620 123600 11880
rect 123900 11620 124100 11880
rect 124400 11620 124600 11880
rect 124900 11620 125100 11880
rect 125400 11620 125600 11880
rect 125900 11620 126100 11880
rect 126400 11620 126600 11880
rect 126900 11620 127000 11880
rect 104000 11600 104120 11620
rect 104380 11600 104620 11620
rect 104880 11600 105120 11620
rect 105380 11600 105620 11620
rect 105880 11600 106120 11620
rect 106380 11600 106620 11620
rect 106880 11600 107120 11620
rect 107380 11600 107620 11620
rect 107880 11600 108120 11620
rect 108380 11600 108620 11620
rect 108880 11600 109120 11620
rect 109380 11600 109620 11620
rect 109880 11600 110120 11620
rect 110380 11600 110620 11620
rect 110880 11600 111120 11620
rect 111380 11600 111620 11620
rect 111880 11600 112120 11620
rect 112380 11600 112620 11620
rect 112880 11600 113120 11620
rect 113380 11600 113620 11620
rect 113880 11600 114120 11620
rect 114380 11600 114620 11620
rect 114880 11600 115120 11620
rect 115380 11600 115620 11620
rect 115880 11600 116120 11620
rect 116380 11600 116620 11620
rect 116880 11600 117120 11620
rect 117380 11600 117620 11620
rect 117880 11600 118120 11620
rect 118380 11600 118620 11620
rect 118880 11600 119120 11620
rect 119380 11600 119620 11620
rect 119880 11600 120120 11620
rect 120380 11600 120620 11620
rect 120880 11600 121120 11620
rect 121380 11600 121620 11620
rect 121880 11600 122120 11620
rect 122380 11600 122620 11620
rect 122880 11600 123120 11620
rect 123380 11600 123620 11620
rect 123880 11600 124120 11620
rect 124380 11600 124620 11620
rect 124880 11600 125120 11620
rect 125380 11600 125620 11620
rect 125880 11600 126120 11620
rect 126380 11600 126620 11620
rect 126880 11600 127000 11620
rect 104000 11400 127000 11600
rect 104000 11380 104120 11400
rect 104380 11380 104620 11400
rect 104880 11380 105120 11400
rect 105380 11380 105620 11400
rect 105880 11380 106120 11400
rect 106380 11380 106620 11400
rect 106880 11380 107120 11400
rect 107380 11380 107620 11400
rect 107880 11380 108120 11400
rect 108380 11380 108620 11400
rect 108880 11380 109120 11400
rect 109380 11380 109620 11400
rect 109880 11380 110120 11400
rect 110380 11380 110620 11400
rect 110880 11380 111120 11400
rect 111380 11380 111620 11400
rect 111880 11380 112120 11400
rect 112380 11380 112620 11400
rect 112880 11380 113120 11400
rect 113380 11380 113620 11400
rect 113880 11380 114120 11400
rect 114380 11380 114620 11400
rect 114880 11380 115120 11400
rect 115380 11380 115620 11400
rect 115880 11380 116120 11400
rect 116380 11380 116620 11400
rect 116880 11380 117120 11400
rect 117380 11380 117620 11400
rect 117880 11380 118120 11400
rect 118380 11380 118620 11400
rect 118880 11380 119120 11400
rect 119380 11380 119620 11400
rect 119880 11380 120120 11400
rect 120380 11380 120620 11400
rect 120880 11380 121120 11400
rect 121380 11380 121620 11400
rect 121880 11380 122120 11400
rect 122380 11380 122620 11400
rect 122880 11380 123120 11400
rect 123380 11380 123620 11400
rect 123880 11380 124120 11400
rect 124380 11380 124620 11400
rect 124880 11380 125120 11400
rect 125380 11380 125620 11400
rect 125880 11380 126120 11400
rect 126380 11380 126620 11400
rect 126880 11380 127000 11400
rect 104000 11120 104100 11380
rect 104400 11120 104600 11380
rect 104900 11120 105100 11380
rect 105400 11120 105600 11380
rect 105900 11120 106100 11380
rect 106400 11120 106600 11380
rect 106900 11120 107100 11380
rect 107400 11120 107600 11380
rect 107900 11120 108100 11380
rect 108400 11120 108600 11380
rect 108900 11120 109100 11380
rect 109400 11120 109600 11380
rect 109900 11120 110100 11380
rect 110400 11120 110600 11380
rect 110900 11120 111100 11380
rect 111400 11120 111600 11380
rect 111900 11120 112100 11380
rect 112400 11120 112600 11380
rect 112900 11120 113100 11380
rect 113400 11120 113600 11380
rect 113900 11120 114100 11380
rect 114400 11120 114600 11380
rect 114900 11120 115100 11380
rect 115400 11120 115600 11380
rect 115900 11120 116100 11380
rect 116400 11120 116600 11380
rect 116900 11120 117100 11380
rect 117400 11120 117600 11380
rect 117900 11120 118100 11380
rect 118400 11120 118600 11380
rect 118900 11120 119100 11380
rect 119400 11120 119600 11380
rect 119900 11120 120100 11380
rect 120400 11120 120600 11380
rect 120900 11120 121100 11380
rect 121400 11120 121600 11380
rect 121900 11120 122100 11380
rect 122400 11120 122600 11380
rect 122900 11120 123100 11380
rect 123400 11120 123600 11380
rect 123900 11120 124100 11380
rect 124400 11120 124600 11380
rect 124900 11120 125100 11380
rect 125400 11120 125600 11380
rect 125900 11120 126100 11380
rect 126400 11120 126600 11380
rect 126900 11120 127000 11380
rect 104000 11100 104120 11120
rect 104380 11100 104620 11120
rect 104880 11100 105120 11120
rect 105380 11100 105620 11120
rect 105880 11100 106120 11120
rect 106380 11100 106620 11120
rect 106880 11100 107120 11120
rect 107380 11100 107620 11120
rect 107880 11100 108120 11120
rect 108380 11100 108620 11120
rect 108880 11100 109120 11120
rect 109380 11100 109620 11120
rect 109880 11100 110120 11120
rect 110380 11100 110620 11120
rect 110880 11100 111120 11120
rect 111380 11100 111620 11120
rect 111880 11100 112120 11120
rect 112380 11100 112620 11120
rect 112880 11100 113120 11120
rect 113380 11100 113620 11120
rect 113880 11100 114120 11120
rect 114380 11100 114620 11120
rect 114880 11100 115120 11120
rect 115380 11100 115620 11120
rect 115880 11100 116120 11120
rect 116380 11100 116620 11120
rect 116880 11100 117120 11120
rect 117380 11100 117620 11120
rect 117880 11100 118120 11120
rect 118380 11100 118620 11120
rect 118880 11100 119120 11120
rect 119380 11100 119620 11120
rect 119880 11100 120120 11120
rect 120380 11100 120620 11120
rect 120880 11100 121120 11120
rect 121380 11100 121620 11120
rect 121880 11100 122120 11120
rect 122380 11100 122620 11120
rect 122880 11100 123120 11120
rect 123380 11100 123620 11120
rect 123880 11100 124120 11120
rect 124380 11100 124620 11120
rect 124880 11100 125120 11120
rect 125380 11100 125620 11120
rect 125880 11100 126120 11120
rect 126380 11100 126620 11120
rect 126880 11100 127000 11120
rect 104000 11000 127000 11100
rect 104000 10980 140000 11000
rect 104000 10910 128150 10980
rect 128350 10910 128650 10980
rect 128850 10910 129150 10980
rect 129350 10910 129650 10980
rect 129850 10910 130150 10980
rect 130350 10910 130650 10980
rect 130850 10910 131150 10980
rect 131350 10910 131650 10980
rect 131850 10910 132150 10980
rect 132350 10910 132650 10980
rect 132850 10910 133150 10980
rect 133350 10910 133650 10980
rect 133850 10910 134150 10980
rect 134350 10910 134650 10980
rect 134850 10910 135150 10980
rect 135350 10910 135650 10980
rect 135850 10910 136150 10980
rect 136350 10910 136650 10980
rect 136850 10910 137150 10980
rect 137350 10910 137650 10980
rect 137850 10910 138150 10980
rect 138350 10910 138650 10980
rect 138850 10910 139150 10980
rect 139350 10910 139650 10980
rect 139850 10910 140000 10980
rect 104000 10900 140000 10910
rect 104000 10880 104120 10900
rect 104380 10880 104620 10900
rect 104880 10880 105120 10900
rect 105380 10880 105620 10900
rect 105880 10880 106120 10900
rect 106380 10880 106620 10900
rect 106880 10880 107120 10900
rect 107380 10880 107620 10900
rect 107880 10880 108120 10900
rect 108380 10880 108620 10900
rect 108880 10880 109120 10900
rect 109380 10880 109620 10900
rect 109880 10880 110120 10900
rect 110380 10880 110620 10900
rect 110880 10880 111120 10900
rect 111380 10880 111620 10900
rect 111880 10880 112120 10900
rect 112380 10880 112620 10900
rect 112880 10880 113120 10900
rect 113380 10880 113620 10900
rect 113880 10880 114120 10900
rect 114380 10880 114620 10900
rect 114880 10880 115120 10900
rect 115380 10880 115620 10900
rect 115880 10880 116120 10900
rect 116380 10880 116620 10900
rect 116880 10880 117120 10900
rect 117380 10880 117620 10900
rect 117880 10880 118120 10900
rect 118380 10880 118620 10900
rect 118880 10880 119120 10900
rect 119380 10880 119620 10900
rect 119880 10880 120120 10900
rect 120380 10880 120620 10900
rect 120880 10880 121120 10900
rect 121380 10880 121620 10900
rect 121880 10880 122120 10900
rect 122380 10880 122620 10900
rect 122880 10880 123120 10900
rect 123380 10880 123620 10900
rect 123880 10880 124120 10900
rect 124380 10880 124620 10900
rect 124880 10880 125120 10900
rect 125380 10880 125620 10900
rect 125880 10880 126120 10900
rect 126380 10880 126620 10900
rect 126880 10880 127120 10900
rect 127380 10880 127620 10900
rect 127880 10880 128120 10900
rect 128380 10880 128620 10900
rect 128880 10880 129120 10900
rect 129380 10880 129620 10900
rect 129880 10880 130120 10900
rect 130380 10880 130620 10900
rect 130880 10880 131120 10900
rect 131380 10880 131620 10900
rect 131880 10880 132120 10900
rect 132380 10880 132620 10900
rect 132880 10880 133120 10900
rect 133380 10880 133620 10900
rect 133880 10880 134120 10900
rect 134380 10880 134620 10900
rect 134880 10880 135120 10900
rect 135380 10880 135620 10900
rect 135880 10880 136120 10900
rect 136380 10880 136620 10900
rect 136880 10880 137120 10900
rect 137380 10880 137620 10900
rect 137880 10880 138120 10900
rect 138380 10880 138620 10900
rect 138880 10880 139120 10900
rect 139380 10880 139620 10900
rect 139880 10880 140000 10900
rect 104000 10620 104100 10880
rect 104400 10620 104600 10880
rect 104900 10620 105100 10880
rect 105400 10620 105600 10880
rect 105900 10620 106100 10880
rect 106400 10620 106600 10880
rect 106900 10620 107100 10880
rect 107400 10620 107600 10880
rect 107900 10620 108100 10880
rect 108400 10620 108600 10880
rect 108900 10620 109100 10880
rect 109400 10620 109600 10880
rect 109900 10620 110100 10880
rect 110400 10620 110600 10880
rect 110900 10620 111100 10880
rect 111400 10620 111600 10880
rect 111900 10620 112100 10880
rect 112400 10620 112600 10880
rect 112900 10620 113100 10880
rect 113400 10620 113600 10880
rect 113900 10620 114100 10880
rect 114400 10620 114600 10880
rect 114900 10620 115100 10880
rect 115400 10620 115600 10880
rect 115900 10620 116100 10880
rect 116400 10620 116600 10880
rect 116900 10620 117100 10880
rect 117400 10620 117600 10880
rect 117900 10620 118100 10880
rect 118400 10620 118600 10880
rect 118900 10620 119100 10880
rect 119400 10620 119600 10880
rect 119900 10620 120100 10880
rect 120400 10620 120600 10880
rect 120900 10620 121100 10880
rect 121400 10620 121600 10880
rect 121900 10620 122100 10880
rect 122400 10620 122600 10880
rect 122900 10620 123100 10880
rect 123400 10620 123600 10880
rect 123900 10620 124100 10880
rect 124400 10620 124600 10880
rect 124900 10620 125100 10880
rect 125400 10620 125600 10880
rect 125900 10620 126100 10880
rect 126400 10620 126600 10880
rect 126900 10620 127100 10880
rect 127400 10620 127600 10880
rect 127900 10850 128100 10880
rect 127900 10650 128020 10850
rect 128090 10650 128100 10850
rect 127900 10620 128100 10650
rect 128400 10850 128600 10880
rect 128400 10650 128410 10850
rect 128480 10650 128520 10850
rect 128590 10650 128600 10850
rect 128400 10620 128600 10650
rect 128900 10850 129100 10880
rect 128900 10650 128910 10850
rect 128980 10650 129020 10850
rect 129090 10650 129100 10850
rect 128900 10620 129100 10650
rect 129400 10850 129600 10880
rect 129400 10650 129410 10850
rect 129480 10650 129520 10850
rect 129590 10650 129600 10850
rect 129400 10620 129600 10650
rect 129900 10850 130100 10880
rect 129900 10650 129910 10850
rect 129980 10650 130020 10850
rect 130090 10650 130100 10850
rect 129900 10620 130100 10650
rect 130400 10850 130600 10880
rect 130400 10650 130410 10850
rect 130480 10650 130520 10850
rect 130590 10650 130600 10850
rect 130400 10620 130600 10650
rect 130900 10850 131100 10880
rect 130900 10650 130910 10850
rect 130980 10650 131020 10850
rect 131090 10650 131100 10850
rect 130900 10620 131100 10650
rect 131400 10850 131600 10880
rect 131400 10650 131410 10850
rect 131480 10650 131520 10850
rect 131590 10650 131600 10850
rect 131400 10620 131600 10650
rect 131900 10850 132100 10880
rect 131900 10650 131910 10850
rect 131980 10650 132020 10850
rect 132090 10650 132100 10850
rect 131900 10620 132100 10650
rect 132400 10850 132600 10880
rect 132400 10650 132410 10850
rect 132480 10650 132520 10850
rect 132590 10650 132600 10850
rect 132400 10620 132600 10650
rect 132900 10850 133100 10880
rect 132900 10650 132910 10850
rect 132980 10650 133020 10850
rect 133090 10650 133100 10850
rect 132900 10620 133100 10650
rect 133400 10850 133600 10880
rect 133400 10650 133410 10850
rect 133480 10650 133520 10850
rect 133590 10650 133600 10850
rect 133400 10620 133600 10650
rect 133900 10850 134100 10880
rect 133900 10650 133910 10850
rect 133980 10650 134020 10850
rect 134090 10650 134100 10850
rect 133900 10620 134100 10650
rect 134400 10850 134600 10880
rect 134400 10650 134410 10850
rect 134480 10650 134520 10850
rect 134590 10650 134600 10850
rect 134400 10620 134600 10650
rect 134900 10850 135100 10880
rect 134900 10650 134910 10850
rect 134980 10650 135020 10850
rect 135090 10650 135100 10850
rect 134900 10620 135100 10650
rect 135400 10850 135600 10880
rect 135400 10650 135410 10850
rect 135480 10650 135520 10850
rect 135590 10650 135600 10850
rect 135400 10620 135600 10650
rect 135900 10850 136100 10880
rect 135900 10650 135910 10850
rect 135980 10650 136020 10850
rect 136090 10650 136100 10850
rect 135900 10620 136100 10650
rect 136400 10850 136600 10880
rect 136400 10650 136410 10850
rect 136480 10650 136520 10850
rect 136590 10650 136600 10850
rect 136400 10620 136600 10650
rect 136900 10850 137100 10880
rect 136900 10650 136910 10850
rect 136980 10650 137020 10850
rect 137090 10650 137100 10850
rect 136900 10620 137100 10650
rect 137400 10850 137600 10880
rect 137400 10650 137410 10850
rect 137480 10650 137520 10850
rect 137590 10650 137600 10850
rect 137400 10620 137600 10650
rect 137900 10850 138100 10880
rect 137900 10650 137910 10850
rect 137980 10650 138020 10850
rect 138090 10650 138100 10850
rect 137900 10620 138100 10650
rect 138400 10850 138600 10880
rect 138400 10650 138410 10850
rect 138480 10650 138520 10850
rect 138590 10650 138600 10850
rect 138400 10620 138600 10650
rect 138900 10850 139100 10880
rect 138900 10650 138910 10850
rect 138980 10650 139020 10850
rect 139090 10650 139100 10850
rect 138900 10620 139100 10650
rect 139400 10850 139600 10880
rect 139400 10650 139410 10850
rect 139480 10650 139520 10850
rect 139590 10650 139600 10850
rect 139400 10620 139600 10650
rect 139900 10850 140000 10880
rect 139900 10650 139910 10850
rect 139980 10650 140000 10850
rect 139900 10620 140000 10650
rect 104000 10600 104120 10620
rect 104380 10600 104620 10620
rect 104880 10600 105120 10620
rect 105380 10600 105620 10620
rect 105880 10600 106120 10620
rect 106380 10600 106620 10620
rect 106880 10600 107120 10620
rect 107380 10600 107620 10620
rect 107880 10600 108120 10620
rect 108380 10600 108620 10620
rect 108880 10600 109120 10620
rect 109380 10600 109620 10620
rect 109880 10600 110120 10620
rect 110380 10600 110620 10620
rect 110880 10600 111120 10620
rect 111380 10600 111620 10620
rect 111880 10600 112120 10620
rect 112380 10600 112620 10620
rect 112880 10600 113120 10620
rect 113380 10600 113620 10620
rect 113880 10600 114120 10620
rect 114380 10600 114620 10620
rect 114880 10600 115120 10620
rect 115380 10600 115620 10620
rect 115880 10600 116120 10620
rect 116380 10600 116620 10620
rect 116880 10600 117120 10620
rect 117380 10600 117620 10620
rect 117880 10600 118120 10620
rect 118380 10600 118620 10620
rect 118880 10600 119120 10620
rect 119380 10600 119620 10620
rect 119880 10600 120120 10620
rect 120380 10600 120620 10620
rect 120880 10600 121120 10620
rect 121380 10600 121620 10620
rect 121880 10600 122120 10620
rect 122380 10600 122620 10620
rect 122880 10600 123120 10620
rect 123380 10600 123620 10620
rect 123880 10600 124120 10620
rect 124380 10600 124620 10620
rect 124880 10600 125120 10620
rect 125380 10600 125620 10620
rect 125880 10600 126120 10620
rect 126380 10600 126620 10620
rect 126880 10600 127120 10620
rect 127380 10600 127620 10620
rect 127880 10600 128120 10620
rect 128380 10600 128620 10620
rect 128880 10600 129120 10620
rect 129380 10600 129620 10620
rect 129880 10600 130120 10620
rect 130380 10600 130620 10620
rect 130880 10600 131120 10620
rect 131380 10600 131620 10620
rect 131880 10600 132120 10620
rect 132380 10600 132620 10620
rect 132880 10600 133120 10620
rect 133380 10600 133620 10620
rect 133880 10600 134120 10620
rect 134380 10600 134620 10620
rect 134880 10600 135120 10620
rect 135380 10600 135620 10620
rect 135880 10600 136120 10620
rect 136380 10600 136620 10620
rect 136880 10600 137120 10620
rect 137380 10600 137620 10620
rect 137880 10600 138120 10620
rect 138380 10600 138620 10620
rect 138880 10600 139120 10620
rect 139380 10600 139620 10620
rect 139880 10600 140000 10620
rect 104000 10590 140000 10600
rect 104000 10520 128150 10590
rect 128350 10520 128650 10590
rect 128850 10520 129150 10590
rect 129350 10520 129650 10590
rect 129850 10520 130150 10590
rect 130350 10520 130650 10590
rect 130850 10520 131150 10590
rect 131350 10520 131650 10590
rect 131850 10520 132150 10590
rect 132350 10520 132650 10590
rect 132850 10520 133150 10590
rect 133350 10520 133650 10590
rect 133850 10520 134150 10590
rect 134350 10520 134650 10590
rect 134850 10520 135150 10590
rect 135350 10520 135650 10590
rect 135850 10520 136150 10590
rect 136350 10520 136650 10590
rect 136850 10520 137150 10590
rect 137350 10520 137650 10590
rect 137850 10520 138150 10590
rect 138350 10520 138650 10590
rect 138850 10520 139150 10590
rect 139350 10520 139650 10590
rect 139850 10520 140000 10590
rect 104000 10480 140000 10520
rect 104000 10410 128150 10480
rect 128350 10410 128650 10480
rect 128850 10410 129150 10480
rect 129350 10410 129650 10480
rect 129850 10410 130150 10480
rect 130350 10410 130650 10480
rect 130850 10410 131150 10480
rect 131350 10410 131650 10480
rect 131850 10410 132150 10480
rect 132350 10410 132650 10480
rect 132850 10410 133150 10480
rect 133350 10410 133650 10480
rect 133850 10410 134150 10480
rect 134350 10410 134650 10480
rect 134850 10410 135150 10480
rect 135350 10410 135650 10480
rect 135850 10410 136150 10480
rect 136350 10410 136650 10480
rect 136850 10410 137150 10480
rect 137350 10410 137650 10480
rect 137850 10410 138150 10480
rect 138350 10410 138650 10480
rect 138850 10410 139150 10480
rect 139350 10410 139650 10480
rect 139850 10410 140000 10480
rect 104000 10400 140000 10410
rect 104000 10380 104120 10400
rect 104380 10380 104620 10400
rect 104880 10380 105120 10400
rect 105380 10380 105620 10400
rect 105880 10380 106120 10400
rect 106380 10380 106620 10400
rect 106880 10380 107120 10400
rect 107380 10380 107620 10400
rect 107880 10380 108120 10400
rect 108380 10380 108620 10400
rect 108880 10380 109120 10400
rect 109380 10380 109620 10400
rect 109880 10380 110120 10400
rect 110380 10380 110620 10400
rect 110880 10380 111120 10400
rect 111380 10380 111620 10400
rect 111880 10380 112120 10400
rect 112380 10380 112620 10400
rect 112880 10380 113120 10400
rect 113380 10380 113620 10400
rect 113880 10380 114120 10400
rect 114380 10380 114620 10400
rect 114880 10380 115120 10400
rect 115380 10380 115620 10400
rect 115880 10380 116120 10400
rect 116380 10380 116620 10400
rect 116880 10380 117120 10400
rect 117380 10380 117620 10400
rect 117880 10380 118120 10400
rect 118380 10380 118620 10400
rect 118880 10380 119120 10400
rect 119380 10380 119620 10400
rect 119880 10380 120120 10400
rect 120380 10380 120620 10400
rect 120880 10380 121120 10400
rect 121380 10380 121620 10400
rect 121880 10380 122120 10400
rect 122380 10380 122620 10400
rect 122880 10380 123120 10400
rect 123380 10380 123620 10400
rect 123880 10380 124120 10400
rect 124380 10380 124620 10400
rect 124880 10380 125120 10400
rect 125380 10380 125620 10400
rect 125880 10380 126120 10400
rect 126380 10380 126620 10400
rect 126880 10380 127120 10400
rect 127380 10380 127620 10400
rect 127880 10380 128120 10400
rect 128380 10380 128620 10400
rect 128880 10380 129120 10400
rect 129380 10380 129620 10400
rect 129880 10380 130120 10400
rect 130380 10380 130620 10400
rect 130880 10380 131120 10400
rect 131380 10380 131620 10400
rect 131880 10380 132120 10400
rect 132380 10380 132620 10400
rect 132880 10380 133120 10400
rect 133380 10380 133620 10400
rect 133880 10380 134120 10400
rect 134380 10380 134620 10400
rect 134880 10380 135120 10400
rect 135380 10380 135620 10400
rect 135880 10380 136120 10400
rect 136380 10380 136620 10400
rect 136880 10380 137120 10400
rect 137380 10380 137620 10400
rect 137880 10380 138120 10400
rect 138380 10380 138620 10400
rect 138880 10380 139120 10400
rect 139380 10380 139620 10400
rect 139880 10380 140000 10400
rect 104000 10120 104100 10380
rect 104400 10120 104600 10380
rect 104900 10120 105100 10380
rect 105400 10120 105600 10380
rect 105900 10120 106100 10380
rect 106400 10120 106600 10380
rect 106900 10120 107100 10380
rect 107400 10120 107600 10380
rect 107900 10120 108100 10380
rect 108400 10120 108600 10380
rect 108900 10120 109100 10380
rect 109400 10120 109600 10380
rect 109900 10120 110100 10380
rect 110400 10120 110600 10380
rect 110900 10120 111100 10380
rect 111400 10120 111600 10380
rect 111900 10120 112100 10380
rect 112400 10120 112600 10380
rect 112900 10120 113100 10380
rect 113400 10120 113600 10380
rect 113900 10120 114100 10380
rect 114400 10120 114600 10380
rect 114900 10120 115100 10380
rect 115400 10120 115600 10380
rect 115900 10120 116100 10380
rect 116400 10120 116600 10380
rect 116900 10120 117100 10380
rect 117400 10120 117600 10380
rect 117900 10120 118100 10380
rect 118400 10120 118600 10380
rect 118900 10120 119100 10380
rect 119400 10120 119600 10380
rect 119900 10120 120100 10380
rect 120400 10120 120600 10380
rect 120900 10120 121100 10380
rect 121400 10120 121600 10380
rect 121900 10120 122100 10380
rect 122400 10120 122600 10380
rect 122900 10120 123100 10380
rect 123400 10120 123600 10380
rect 123900 10120 124100 10380
rect 124400 10120 124600 10380
rect 124900 10120 125100 10380
rect 125400 10120 125600 10380
rect 125900 10120 126100 10380
rect 126400 10120 126600 10380
rect 126900 10120 127100 10380
rect 127400 10120 127600 10380
rect 127900 10350 128100 10380
rect 127900 10150 128020 10350
rect 128090 10150 128100 10350
rect 127900 10120 128100 10150
rect 128400 10350 128600 10380
rect 128400 10150 128410 10350
rect 128480 10150 128520 10350
rect 128590 10150 128600 10350
rect 128400 10120 128600 10150
rect 128900 10350 129100 10380
rect 128900 10150 128910 10350
rect 128980 10150 129020 10350
rect 129090 10150 129100 10350
rect 128900 10120 129100 10150
rect 129400 10350 129600 10380
rect 129400 10150 129410 10350
rect 129480 10150 129520 10350
rect 129590 10150 129600 10350
rect 129400 10120 129600 10150
rect 129900 10350 130100 10380
rect 129900 10150 129910 10350
rect 129980 10150 130020 10350
rect 130090 10150 130100 10350
rect 129900 10120 130100 10150
rect 130400 10350 130600 10380
rect 130400 10150 130410 10350
rect 130480 10150 130520 10350
rect 130590 10150 130600 10350
rect 130400 10120 130600 10150
rect 130900 10350 131100 10380
rect 130900 10150 130910 10350
rect 130980 10150 131020 10350
rect 131090 10150 131100 10350
rect 130900 10120 131100 10150
rect 131400 10350 131600 10380
rect 131400 10150 131410 10350
rect 131480 10150 131520 10350
rect 131590 10150 131600 10350
rect 131400 10120 131600 10150
rect 131900 10350 132100 10380
rect 131900 10150 131910 10350
rect 131980 10150 132020 10350
rect 132090 10150 132100 10350
rect 131900 10120 132100 10150
rect 132400 10350 132600 10380
rect 132400 10150 132410 10350
rect 132480 10150 132520 10350
rect 132590 10150 132600 10350
rect 132400 10120 132600 10150
rect 132900 10350 133100 10380
rect 132900 10150 132910 10350
rect 132980 10150 133020 10350
rect 133090 10150 133100 10350
rect 132900 10120 133100 10150
rect 133400 10350 133600 10380
rect 133400 10150 133410 10350
rect 133480 10150 133520 10350
rect 133590 10150 133600 10350
rect 133400 10120 133600 10150
rect 133900 10350 134100 10380
rect 133900 10150 133910 10350
rect 133980 10150 134020 10350
rect 134090 10150 134100 10350
rect 133900 10120 134100 10150
rect 134400 10350 134600 10380
rect 134400 10150 134410 10350
rect 134480 10150 134520 10350
rect 134590 10150 134600 10350
rect 134400 10120 134600 10150
rect 134900 10350 135100 10380
rect 134900 10150 134910 10350
rect 134980 10150 135020 10350
rect 135090 10150 135100 10350
rect 134900 10120 135100 10150
rect 135400 10350 135600 10380
rect 135400 10150 135410 10350
rect 135480 10150 135520 10350
rect 135590 10150 135600 10350
rect 135400 10120 135600 10150
rect 135900 10350 136100 10380
rect 135900 10150 135910 10350
rect 135980 10150 136020 10350
rect 136090 10150 136100 10350
rect 135900 10120 136100 10150
rect 136400 10350 136600 10380
rect 136400 10150 136410 10350
rect 136480 10150 136520 10350
rect 136590 10150 136600 10350
rect 136400 10120 136600 10150
rect 136900 10350 137100 10380
rect 136900 10150 136910 10350
rect 136980 10150 137020 10350
rect 137090 10150 137100 10350
rect 136900 10120 137100 10150
rect 137400 10350 137600 10380
rect 137400 10150 137410 10350
rect 137480 10150 137520 10350
rect 137590 10150 137600 10350
rect 137400 10120 137600 10150
rect 137900 10350 138100 10380
rect 137900 10150 137910 10350
rect 137980 10150 138020 10350
rect 138090 10150 138100 10350
rect 137900 10120 138100 10150
rect 138400 10350 138600 10380
rect 138400 10150 138410 10350
rect 138480 10150 138520 10350
rect 138590 10150 138600 10350
rect 138400 10120 138600 10150
rect 138900 10350 139100 10380
rect 138900 10150 138910 10350
rect 138980 10150 139020 10350
rect 139090 10150 139100 10350
rect 138900 10120 139100 10150
rect 139400 10350 139600 10380
rect 139400 10150 139410 10350
rect 139480 10150 139520 10350
rect 139590 10150 139600 10350
rect 139400 10120 139600 10150
rect 139900 10350 140000 10380
rect 139900 10150 139910 10350
rect 139980 10150 140000 10350
rect 139900 10120 140000 10150
rect 104000 10100 104120 10120
rect 104380 10100 104620 10120
rect 104880 10100 105120 10120
rect 105380 10100 105620 10120
rect 105880 10100 106120 10120
rect 106380 10100 106620 10120
rect 106880 10100 107120 10120
rect 107380 10100 107620 10120
rect 107880 10100 108120 10120
rect 108380 10100 108620 10120
rect 108880 10100 109120 10120
rect 109380 10100 109620 10120
rect 109880 10100 110120 10120
rect 110380 10100 110620 10120
rect 110880 10100 111120 10120
rect 111380 10100 111620 10120
rect 111880 10100 112120 10120
rect 112380 10100 112620 10120
rect 112880 10100 113120 10120
rect 113380 10100 113620 10120
rect 113880 10100 114120 10120
rect 114380 10100 114620 10120
rect 114880 10100 115120 10120
rect 115380 10100 115620 10120
rect 115880 10100 116120 10120
rect 116380 10100 116620 10120
rect 116880 10100 117120 10120
rect 117380 10100 117620 10120
rect 117880 10100 118120 10120
rect 118380 10100 118620 10120
rect 118880 10100 119120 10120
rect 119380 10100 119620 10120
rect 119880 10100 120120 10120
rect 120380 10100 120620 10120
rect 120880 10100 121120 10120
rect 121380 10100 121620 10120
rect 121880 10100 122120 10120
rect 122380 10100 122620 10120
rect 122880 10100 123120 10120
rect 123380 10100 123620 10120
rect 123880 10100 124120 10120
rect 124380 10100 124620 10120
rect 124880 10100 125120 10120
rect 125380 10100 125620 10120
rect 125880 10100 126120 10120
rect 126380 10100 126620 10120
rect 126880 10100 127120 10120
rect 127380 10100 127620 10120
rect 127880 10100 128120 10120
rect 128380 10100 128620 10120
rect 128880 10100 129120 10120
rect 129380 10100 129620 10120
rect 129880 10100 130120 10120
rect 130380 10100 130620 10120
rect 130880 10100 131120 10120
rect 131380 10100 131620 10120
rect 131880 10100 132120 10120
rect 132380 10100 132620 10120
rect 132880 10100 133120 10120
rect 133380 10100 133620 10120
rect 133880 10100 134120 10120
rect 134380 10100 134620 10120
rect 134880 10100 135120 10120
rect 135380 10100 135620 10120
rect 135880 10100 136120 10120
rect 136380 10100 136620 10120
rect 136880 10100 137120 10120
rect 137380 10100 137620 10120
rect 137880 10100 138120 10120
rect 138380 10100 138620 10120
rect 138880 10100 139120 10120
rect 139380 10100 139620 10120
rect 139880 10100 140000 10120
rect 104000 10090 140000 10100
rect 104000 10020 128150 10090
rect 128350 10020 128650 10090
rect 128850 10020 129150 10090
rect 129350 10020 129650 10090
rect 129850 10020 130150 10090
rect 130350 10020 130650 10090
rect 130850 10020 131150 10090
rect 131350 10020 131650 10090
rect 131850 10020 132150 10090
rect 132350 10020 132650 10090
rect 132850 10020 133150 10090
rect 133350 10020 133650 10090
rect 133850 10020 134150 10090
rect 134350 10020 134650 10090
rect 134850 10020 135150 10090
rect 135350 10020 135650 10090
rect 135850 10020 136150 10090
rect 136350 10020 136650 10090
rect 136850 10020 137150 10090
rect 137350 10020 137650 10090
rect 137850 10020 138150 10090
rect 138350 10020 138650 10090
rect 138850 10020 139150 10090
rect 139350 10020 139650 10090
rect 139850 10020 140000 10090
rect 104000 9980 140000 10020
rect 104000 9910 128150 9980
rect 128350 9910 128650 9980
rect 128850 9910 129150 9980
rect 129350 9910 129650 9980
rect 129850 9910 130150 9980
rect 130350 9910 130650 9980
rect 130850 9910 131150 9980
rect 131350 9910 131650 9980
rect 131850 9910 132150 9980
rect 132350 9910 132650 9980
rect 132850 9910 133150 9980
rect 133350 9910 133650 9980
rect 133850 9910 134150 9980
rect 134350 9910 134650 9980
rect 134850 9910 135150 9980
rect 135350 9910 135650 9980
rect 135850 9910 136150 9980
rect 136350 9910 136650 9980
rect 136850 9910 137150 9980
rect 137350 9910 137650 9980
rect 137850 9910 138150 9980
rect 138350 9910 138650 9980
rect 138850 9910 139150 9980
rect 139350 9910 139650 9980
rect 139850 9910 140000 9980
rect 104000 9900 140000 9910
rect 104000 9880 104120 9900
rect 104380 9880 104620 9900
rect 104880 9880 105120 9900
rect 105380 9880 105620 9900
rect 105880 9880 106120 9900
rect 106380 9880 106620 9900
rect 106880 9880 107120 9900
rect 107380 9880 107620 9900
rect 107880 9880 108120 9900
rect 108380 9880 108620 9900
rect 108880 9880 109120 9900
rect 109380 9880 109620 9900
rect 109880 9880 110120 9900
rect 110380 9880 110620 9900
rect 110880 9880 111120 9900
rect 111380 9880 111620 9900
rect 111880 9880 112120 9900
rect 112380 9880 112620 9900
rect 112880 9880 113120 9900
rect 113380 9880 113620 9900
rect 113880 9880 114120 9900
rect 114380 9880 114620 9900
rect 114880 9880 115120 9900
rect 115380 9880 115620 9900
rect 115880 9880 116120 9900
rect 116380 9880 116620 9900
rect 116880 9880 117120 9900
rect 117380 9880 117620 9900
rect 117880 9880 118120 9900
rect 118380 9880 118620 9900
rect 118880 9880 119120 9900
rect 119380 9880 119620 9900
rect 119880 9880 120120 9900
rect 120380 9880 120620 9900
rect 120880 9880 121120 9900
rect 121380 9880 121620 9900
rect 121880 9880 122120 9900
rect 122380 9880 122620 9900
rect 122880 9880 123120 9900
rect 123380 9880 123620 9900
rect 123880 9880 124120 9900
rect 124380 9880 124620 9900
rect 124880 9880 125120 9900
rect 125380 9880 125620 9900
rect 125880 9880 126120 9900
rect 126380 9880 126620 9900
rect 126880 9880 127120 9900
rect 127380 9880 127620 9900
rect 127880 9880 128120 9900
rect 128380 9880 128620 9900
rect 128880 9880 129120 9900
rect 129380 9880 129620 9900
rect 129880 9880 130120 9900
rect 130380 9880 130620 9900
rect 130880 9880 131120 9900
rect 131380 9880 131620 9900
rect 131880 9880 132120 9900
rect 132380 9880 132620 9900
rect 132880 9880 133120 9900
rect 133380 9880 133620 9900
rect 133880 9880 134120 9900
rect 134380 9880 134620 9900
rect 134880 9880 135120 9900
rect 135380 9880 135620 9900
rect 135880 9880 136120 9900
rect 136380 9880 136620 9900
rect 136880 9880 137120 9900
rect 137380 9880 137620 9900
rect 137880 9880 138120 9900
rect 138380 9880 138620 9900
rect 138880 9880 139120 9900
rect 139380 9880 139620 9900
rect 139880 9880 140000 9900
rect 104000 9620 104100 9880
rect 104400 9620 104600 9880
rect 104900 9620 105100 9880
rect 105400 9620 105600 9880
rect 105900 9620 106100 9880
rect 106400 9620 106600 9880
rect 106900 9620 107100 9880
rect 107400 9620 107600 9880
rect 107900 9620 108100 9880
rect 108400 9620 108600 9880
rect 108900 9620 109100 9880
rect 109400 9620 109600 9880
rect 109900 9620 110100 9880
rect 110400 9620 110600 9880
rect 110900 9620 111100 9880
rect 111400 9620 111600 9880
rect 111900 9620 112100 9880
rect 112400 9620 112600 9880
rect 112900 9620 113100 9880
rect 113400 9620 113600 9880
rect 113900 9620 114100 9880
rect 114400 9620 114600 9880
rect 114900 9620 115100 9880
rect 115400 9620 115600 9880
rect 115900 9620 116100 9880
rect 116400 9620 116600 9880
rect 116900 9620 117100 9880
rect 117400 9620 117600 9880
rect 117900 9620 118100 9880
rect 118400 9620 118600 9880
rect 118900 9620 119100 9880
rect 119400 9620 119600 9880
rect 119900 9620 120100 9880
rect 120400 9620 120600 9880
rect 120900 9620 121100 9880
rect 121400 9620 121600 9880
rect 121900 9620 122100 9880
rect 122400 9620 122600 9880
rect 122900 9620 123100 9880
rect 123400 9620 123600 9880
rect 123900 9620 124100 9880
rect 124400 9620 124600 9880
rect 124900 9620 125100 9880
rect 125400 9620 125600 9880
rect 125900 9620 126100 9880
rect 126400 9620 126600 9880
rect 126900 9620 127100 9880
rect 127400 9620 127600 9880
rect 127900 9850 128100 9880
rect 127900 9650 128020 9850
rect 128090 9650 128100 9850
rect 127900 9620 128100 9650
rect 128400 9850 128600 9880
rect 128400 9650 128410 9850
rect 128480 9650 128520 9850
rect 128590 9650 128600 9850
rect 128400 9620 128600 9650
rect 128900 9850 129100 9880
rect 128900 9650 128910 9850
rect 128980 9650 129020 9850
rect 129090 9650 129100 9850
rect 128900 9620 129100 9650
rect 129400 9850 129600 9880
rect 129400 9650 129410 9850
rect 129480 9650 129520 9850
rect 129590 9650 129600 9850
rect 129400 9620 129600 9650
rect 129900 9850 130100 9880
rect 129900 9650 129910 9850
rect 129980 9650 130020 9850
rect 130090 9650 130100 9850
rect 129900 9620 130100 9650
rect 130400 9850 130600 9880
rect 130400 9650 130410 9850
rect 130480 9650 130520 9850
rect 130590 9650 130600 9850
rect 130400 9620 130600 9650
rect 130900 9850 131100 9880
rect 130900 9650 130910 9850
rect 130980 9650 131020 9850
rect 131090 9650 131100 9850
rect 130900 9620 131100 9650
rect 131400 9850 131600 9880
rect 131400 9650 131410 9850
rect 131480 9650 131520 9850
rect 131590 9650 131600 9850
rect 131400 9620 131600 9650
rect 131900 9850 132100 9880
rect 131900 9650 131910 9850
rect 131980 9650 132020 9850
rect 132090 9650 132100 9850
rect 131900 9620 132100 9650
rect 132400 9850 132600 9880
rect 132400 9650 132410 9850
rect 132480 9650 132520 9850
rect 132590 9650 132600 9850
rect 132400 9620 132600 9650
rect 132900 9850 133100 9880
rect 132900 9650 132910 9850
rect 132980 9650 133020 9850
rect 133090 9650 133100 9850
rect 132900 9620 133100 9650
rect 133400 9850 133600 9880
rect 133400 9650 133410 9850
rect 133480 9650 133520 9850
rect 133590 9650 133600 9850
rect 133400 9620 133600 9650
rect 133900 9850 134100 9880
rect 133900 9650 133910 9850
rect 133980 9650 134020 9850
rect 134090 9650 134100 9850
rect 133900 9620 134100 9650
rect 134400 9850 134600 9880
rect 134400 9650 134410 9850
rect 134480 9650 134520 9850
rect 134590 9650 134600 9850
rect 134400 9620 134600 9650
rect 134900 9850 135100 9880
rect 134900 9650 134910 9850
rect 134980 9650 135020 9850
rect 135090 9650 135100 9850
rect 134900 9620 135100 9650
rect 135400 9850 135600 9880
rect 135400 9650 135410 9850
rect 135480 9650 135520 9850
rect 135590 9650 135600 9850
rect 135400 9620 135600 9650
rect 135900 9850 136100 9880
rect 135900 9650 135910 9850
rect 135980 9650 136020 9850
rect 136090 9650 136100 9850
rect 135900 9620 136100 9650
rect 136400 9850 136600 9880
rect 136400 9650 136410 9850
rect 136480 9650 136520 9850
rect 136590 9650 136600 9850
rect 136400 9620 136600 9650
rect 136900 9850 137100 9880
rect 136900 9650 136910 9850
rect 136980 9650 137020 9850
rect 137090 9650 137100 9850
rect 136900 9620 137100 9650
rect 137400 9850 137600 9880
rect 137400 9650 137410 9850
rect 137480 9650 137520 9850
rect 137590 9650 137600 9850
rect 137400 9620 137600 9650
rect 137900 9850 138100 9880
rect 137900 9650 137910 9850
rect 137980 9650 138020 9850
rect 138090 9650 138100 9850
rect 137900 9620 138100 9650
rect 138400 9850 138600 9880
rect 138400 9650 138410 9850
rect 138480 9650 138520 9850
rect 138590 9650 138600 9850
rect 138400 9620 138600 9650
rect 138900 9850 139100 9880
rect 138900 9650 138910 9850
rect 138980 9650 139020 9850
rect 139090 9650 139100 9850
rect 138900 9620 139100 9650
rect 139400 9850 139600 9880
rect 139400 9650 139410 9850
rect 139480 9650 139520 9850
rect 139590 9650 139600 9850
rect 139400 9620 139600 9650
rect 139900 9850 140000 9880
rect 139900 9650 139910 9850
rect 139980 9650 140000 9850
rect 139900 9620 140000 9650
rect 104000 9600 104120 9620
rect 104380 9600 104620 9620
rect 104880 9600 105120 9620
rect 105380 9600 105620 9620
rect 105880 9600 106120 9620
rect 106380 9600 106620 9620
rect 106880 9600 107120 9620
rect 107380 9600 107620 9620
rect 107880 9600 108120 9620
rect 108380 9600 108620 9620
rect 108880 9600 109120 9620
rect 109380 9600 109620 9620
rect 109880 9600 110120 9620
rect 110380 9600 110620 9620
rect 110880 9600 111120 9620
rect 111380 9600 111620 9620
rect 111880 9600 112120 9620
rect 112380 9600 112620 9620
rect 112880 9600 113120 9620
rect 113380 9600 113620 9620
rect 113880 9600 114120 9620
rect 114380 9600 114620 9620
rect 114880 9600 115120 9620
rect 115380 9600 115620 9620
rect 115880 9600 116120 9620
rect 116380 9600 116620 9620
rect 116880 9600 117120 9620
rect 117380 9600 117620 9620
rect 117880 9600 118120 9620
rect 118380 9600 118620 9620
rect 118880 9600 119120 9620
rect 119380 9600 119620 9620
rect 119880 9600 120120 9620
rect 120380 9600 120620 9620
rect 120880 9600 121120 9620
rect 121380 9600 121620 9620
rect 121880 9600 122120 9620
rect 122380 9600 122620 9620
rect 122880 9600 123120 9620
rect 123380 9600 123620 9620
rect 123880 9600 124120 9620
rect 124380 9600 124620 9620
rect 124880 9600 125120 9620
rect 125380 9600 125620 9620
rect 125880 9600 126120 9620
rect 126380 9600 126620 9620
rect 126880 9600 127120 9620
rect 127380 9600 127620 9620
rect 127880 9600 128120 9620
rect 128380 9600 128620 9620
rect 128880 9600 129120 9620
rect 129380 9600 129620 9620
rect 129880 9600 130120 9620
rect 130380 9600 130620 9620
rect 130880 9600 131120 9620
rect 131380 9600 131620 9620
rect 131880 9600 132120 9620
rect 132380 9600 132620 9620
rect 132880 9600 133120 9620
rect 133380 9600 133620 9620
rect 133880 9600 134120 9620
rect 134380 9600 134620 9620
rect 134880 9600 135120 9620
rect 135380 9600 135620 9620
rect 135880 9600 136120 9620
rect 136380 9600 136620 9620
rect 136880 9600 137120 9620
rect 137380 9600 137620 9620
rect 137880 9600 138120 9620
rect 138380 9600 138620 9620
rect 138880 9600 139120 9620
rect 139380 9600 139620 9620
rect 139880 9600 140000 9620
rect 104000 9590 140000 9600
rect 104000 9520 128150 9590
rect 128350 9520 128650 9590
rect 128850 9520 129150 9590
rect 129350 9520 129650 9590
rect 129850 9520 130150 9590
rect 130350 9520 130650 9590
rect 130850 9520 131150 9590
rect 131350 9520 131650 9590
rect 131850 9520 132150 9590
rect 132350 9520 132650 9590
rect 132850 9520 133150 9590
rect 133350 9520 133650 9590
rect 133850 9520 134150 9590
rect 134350 9520 134650 9590
rect 134850 9520 135150 9590
rect 135350 9520 135650 9590
rect 135850 9520 136150 9590
rect 136350 9520 136650 9590
rect 136850 9520 137150 9590
rect 137350 9520 137650 9590
rect 137850 9520 138150 9590
rect 138350 9520 138650 9590
rect 138850 9520 139150 9590
rect 139350 9520 139650 9590
rect 139850 9520 140000 9590
rect 104000 9480 140000 9520
rect 104000 9410 128150 9480
rect 128350 9410 128650 9480
rect 128850 9410 129150 9480
rect 129350 9410 129650 9480
rect 129850 9410 130150 9480
rect 130350 9410 130650 9480
rect 130850 9410 131150 9480
rect 131350 9410 131650 9480
rect 131850 9410 132150 9480
rect 132350 9410 132650 9480
rect 132850 9410 133150 9480
rect 133350 9410 133650 9480
rect 133850 9410 134150 9480
rect 134350 9410 134650 9480
rect 134850 9410 135150 9480
rect 135350 9410 135650 9480
rect 135850 9410 136150 9480
rect 136350 9410 136650 9480
rect 136850 9410 137150 9480
rect 137350 9410 137650 9480
rect 137850 9410 138150 9480
rect 138350 9410 138650 9480
rect 138850 9410 139150 9480
rect 139350 9410 139650 9480
rect 139850 9410 140000 9480
rect 104000 9400 140000 9410
rect 104000 9380 104120 9400
rect 104380 9380 104620 9400
rect 104880 9380 105120 9400
rect 105380 9380 105620 9400
rect 105880 9380 106120 9400
rect 106380 9380 106620 9400
rect 106880 9380 107120 9400
rect 107380 9380 107620 9400
rect 107880 9380 108120 9400
rect 108380 9380 108620 9400
rect 108880 9380 109120 9400
rect 109380 9380 109620 9400
rect 109880 9380 110120 9400
rect 110380 9380 110620 9400
rect 110880 9380 111120 9400
rect 111380 9380 111620 9400
rect 111880 9380 112120 9400
rect 112380 9380 112620 9400
rect 112880 9380 113120 9400
rect 113380 9380 113620 9400
rect 113880 9380 114120 9400
rect 114380 9380 114620 9400
rect 114880 9380 115120 9400
rect 115380 9380 115620 9400
rect 115880 9380 116120 9400
rect 116380 9380 116620 9400
rect 116880 9380 117120 9400
rect 117380 9380 117620 9400
rect 117880 9380 118120 9400
rect 118380 9380 118620 9400
rect 118880 9380 119120 9400
rect 119380 9380 119620 9400
rect 119880 9380 120120 9400
rect 120380 9380 120620 9400
rect 120880 9380 121120 9400
rect 121380 9380 121620 9400
rect 121880 9380 122120 9400
rect 122380 9380 122620 9400
rect 122880 9380 123120 9400
rect 123380 9380 123620 9400
rect 123880 9380 124120 9400
rect 124380 9380 124620 9400
rect 124880 9380 125120 9400
rect 125380 9380 125620 9400
rect 125880 9380 126120 9400
rect 126380 9380 126620 9400
rect 126880 9380 127120 9400
rect 127380 9380 127620 9400
rect 127880 9380 128120 9400
rect 128380 9380 128620 9400
rect 128880 9380 129120 9400
rect 129380 9380 129620 9400
rect 129880 9380 130120 9400
rect 130380 9380 130620 9400
rect 130880 9380 131120 9400
rect 131380 9380 131620 9400
rect 131880 9380 132120 9400
rect 132380 9380 132620 9400
rect 132880 9380 133120 9400
rect 133380 9380 133620 9400
rect 133880 9380 134120 9400
rect 134380 9380 134620 9400
rect 134880 9380 135120 9400
rect 135380 9380 135620 9400
rect 135880 9380 136120 9400
rect 136380 9380 136620 9400
rect 136880 9380 137120 9400
rect 137380 9380 137620 9400
rect 137880 9380 138120 9400
rect 138380 9380 138620 9400
rect 138880 9380 139120 9400
rect 139380 9380 139620 9400
rect 139880 9380 140000 9400
rect 104000 9120 104100 9380
rect 104400 9120 104600 9380
rect 104900 9120 105100 9380
rect 105400 9120 105600 9380
rect 105900 9120 106100 9380
rect 106400 9120 106600 9380
rect 106900 9120 107100 9380
rect 107400 9120 107600 9380
rect 107900 9120 108100 9380
rect 108400 9120 108600 9380
rect 108900 9120 109100 9380
rect 109400 9120 109600 9380
rect 109900 9120 110100 9380
rect 110400 9120 110600 9380
rect 110900 9120 111100 9380
rect 111400 9120 111600 9380
rect 111900 9120 112100 9380
rect 112400 9120 112600 9380
rect 112900 9120 113100 9380
rect 113400 9120 113600 9380
rect 113900 9120 114100 9380
rect 114400 9120 114600 9380
rect 114900 9120 115100 9380
rect 115400 9120 115600 9380
rect 115900 9120 116100 9380
rect 116400 9120 116600 9380
rect 116900 9120 117100 9380
rect 117400 9120 117600 9380
rect 117900 9120 118100 9380
rect 118400 9120 118600 9380
rect 118900 9120 119100 9380
rect 119400 9120 119600 9380
rect 119900 9120 120100 9380
rect 120400 9120 120600 9380
rect 120900 9120 121100 9380
rect 121400 9120 121600 9380
rect 121900 9120 122100 9380
rect 122400 9120 122600 9380
rect 122900 9120 123100 9380
rect 123400 9120 123600 9380
rect 123900 9120 124100 9380
rect 124400 9120 124600 9380
rect 124900 9120 125100 9380
rect 125400 9120 125600 9380
rect 125900 9120 126100 9380
rect 126400 9120 126600 9380
rect 126900 9120 127100 9380
rect 127400 9120 127600 9380
rect 127900 9350 128100 9380
rect 127900 9150 128020 9350
rect 128090 9150 128100 9350
rect 127900 9120 128100 9150
rect 128400 9350 128600 9380
rect 128400 9150 128410 9350
rect 128480 9150 128520 9350
rect 128590 9150 128600 9350
rect 128400 9120 128600 9150
rect 128900 9350 129100 9380
rect 128900 9150 128910 9350
rect 128980 9150 129020 9350
rect 129090 9150 129100 9350
rect 128900 9120 129100 9150
rect 129400 9350 129600 9380
rect 129400 9150 129410 9350
rect 129480 9150 129520 9350
rect 129590 9150 129600 9350
rect 129400 9120 129600 9150
rect 129900 9350 130100 9380
rect 129900 9150 129910 9350
rect 129980 9150 130020 9350
rect 130090 9150 130100 9350
rect 129900 9120 130100 9150
rect 130400 9350 130600 9380
rect 130400 9150 130410 9350
rect 130480 9150 130520 9350
rect 130590 9150 130600 9350
rect 130400 9120 130600 9150
rect 130900 9350 131100 9380
rect 130900 9150 130910 9350
rect 130980 9150 131020 9350
rect 131090 9150 131100 9350
rect 130900 9120 131100 9150
rect 131400 9350 131600 9380
rect 131400 9150 131410 9350
rect 131480 9150 131520 9350
rect 131590 9150 131600 9350
rect 131400 9120 131600 9150
rect 131900 9350 132100 9380
rect 131900 9150 131910 9350
rect 131980 9150 132020 9350
rect 132090 9150 132100 9350
rect 131900 9120 132100 9150
rect 132400 9350 132600 9380
rect 132400 9150 132410 9350
rect 132480 9150 132520 9350
rect 132590 9150 132600 9350
rect 132400 9120 132600 9150
rect 132900 9350 133100 9380
rect 132900 9150 132910 9350
rect 132980 9150 133020 9350
rect 133090 9150 133100 9350
rect 132900 9120 133100 9150
rect 133400 9350 133600 9380
rect 133400 9150 133410 9350
rect 133480 9150 133520 9350
rect 133590 9150 133600 9350
rect 133400 9120 133600 9150
rect 133900 9350 134100 9380
rect 133900 9150 133910 9350
rect 133980 9150 134020 9350
rect 134090 9150 134100 9350
rect 133900 9120 134100 9150
rect 134400 9350 134600 9380
rect 134400 9150 134410 9350
rect 134480 9150 134520 9350
rect 134590 9150 134600 9350
rect 134400 9120 134600 9150
rect 134900 9350 135100 9380
rect 134900 9150 134910 9350
rect 134980 9150 135020 9350
rect 135090 9150 135100 9350
rect 134900 9120 135100 9150
rect 135400 9350 135600 9380
rect 135400 9150 135410 9350
rect 135480 9150 135520 9350
rect 135590 9150 135600 9350
rect 135400 9120 135600 9150
rect 135900 9350 136100 9380
rect 135900 9150 135910 9350
rect 135980 9150 136020 9350
rect 136090 9150 136100 9350
rect 135900 9120 136100 9150
rect 136400 9350 136600 9380
rect 136400 9150 136410 9350
rect 136480 9150 136520 9350
rect 136590 9150 136600 9350
rect 136400 9120 136600 9150
rect 136900 9350 137100 9380
rect 136900 9150 136910 9350
rect 136980 9150 137020 9350
rect 137090 9150 137100 9350
rect 136900 9120 137100 9150
rect 137400 9350 137600 9380
rect 137400 9150 137410 9350
rect 137480 9150 137520 9350
rect 137590 9150 137600 9350
rect 137400 9120 137600 9150
rect 137900 9350 138100 9380
rect 137900 9150 137910 9350
rect 137980 9150 138020 9350
rect 138090 9150 138100 9350
rect 137900 9120 138100 9150
rect 138400 9350 138600 9380
rect 138400 9150 138410 9350
rect 138480 9150 138520 9350
rect 138590 9150 138600 9350
rect 138400 9120 138600 9150
rect 138900 9350 139100 9380
rect 138900 9150 138910 9350
rect 138980 9150 139020 9350
rect 139090 9150 139100 9350
rect 138900 9120 139100 9150
rect 139400 9350 139600 9380
rect 139400 9150 139410 9350
rect 139480 9150 139520 9350
rect 139590 9150 139600 9350
rect 139400 9120 139600 9150
rect 139900 9350 140000 9380
rect 139900 9150 139910 9350
rect 139980 9150 140000 9350
rect 139900 9120 140000 9150
rect 104000 9100 104120 9120
rect 104380 9100 104620 9120
rect 104880 9100 105120 9120
rect 105380 9100 105620 9120
rect 105880 9100 106120 9120
rect 106380 9100 106620 9120
rect 106880 9100 107120 9120
rect 107380 9100 107620 9120
rect 107880 9100 108120 9120
rect 108380 9100 108620 9120
rect 108880 9100 109120 9120
rect 109380 9100 109620 9120
rect 109880 9100 110120 9120
rect 110380 9100 110620 9120
rect 110880 9100 111120 9120
rect 111380 9100 111620 9120
rect 111880 9100 112120 9120
rect 112380 9100 112620 9120
rect 112880 9100 113120 9120
rect 113380 9100 113620 9120
rect 113880 9100 114120 9120
rect 114380 9100 114620 9120
rect 114880 9100 115120 9120
rect 115380 9100 115620 9120
rect 115880 9100 116120 9120
rect 116380 9100 116620 9120
rect 116880 9100 117120 9120
rect 117380 9100 117620 9120
rect 117880 9100 118120 9120
rect 118380 9100 118620 9120
rect 118880 9100 119120 9120
rect 119380 9100 119620 9120
rect 119880 9100 120120 9120
rect 120380 9100 120620 9120
rect 120880 9100 121120 9120
rect 121380 9100 121620 9120
rect 121880 9100 122120 9120
rect 122380 9100 122620 9120
rect 122880 9100 123120 9120
rect 123380 9100 123620 9120
rect 123880 9100 124120 9120
rect 124380 9100 124620 9120
rect 124880 9100 125120 9120
rect 125380 9100 125620 9120
rect 125880 9100 126120 9120
rect 126380 9100 126620 9120
rect 126880 9100 127120 9120
rect 127380 9100 127620 9120
rect 127880 9100 128120 9120
rect 128380 9100 128620 9120
rect 128880 9100 129120 9120
rect 129380 9100 129620 9120
rect 129880 9100 130120 9120
rect 130380 9100 130620 9120
rect 130880 9100 131120 9120
rect 131380 9100 131620 9120
rect 131880 9100 132120 9120
rect 132380 9100 132620 9120
rect 132880 9100 133120 9120
rect 133380 9100 133620 9120
rect 133880 9100 134120 9120
rect 134380 9100 134620 9120
rect 134880 9100 135120 9120
rect 135380 9100 135620 9120
rect 135880 9100 136120 9120
rect 136380 9100 136620 9120
rect 136880 9100 137120 9120
rect 137380 9100 137620 9120
rect 137880 9100 138120 9120
rect 138380 9100 138620 9120
rect 138880 9100 139120 9120
rect 139380 9100 139620 9120
rect 139880 9100 140000 9120
rect 104000 9090 140000 9100
rect 104000 9020 128150 9090
rect 128350 9020 128650 9090
rect 128850 9020 129150 9090
rect 129350 9020 129650 9090
rect 129850 9020 130150 9090
rect 130350 9020 130650 9090
rect 130850 9020 131150 9090
rect 131350 9020 131650 9090
rect 131850 9020 132150 9090
rect 132350 9020 132650 9090
rect 132850 9020 133150 9090
rect 133350 9020 133650 9090
rect 133850 9020 134150 9090
rect 134350 9020 134650 9090
rect 134850 9020 135150 9090
rect 135350 9020 135650 9090
rect 135850 9020 136150 9090
rect 136350 9020 136650 9090
rect 136850 9020 137150 9090
rect 137350 9020 137650 9090
rect 137850 9020 138150 9090
rect 138350 9020 138650 9090
rect 138850 9020 139150 9090
rect 139350 9020 139650 9090
rect 139850 9020 140000 9090
rect 104000 8980 140000 9020
rect 104000 8910 128150 8980
rect 128350 8910 128650 8980
rect 128850 8910 129150 8980
rect 129350 8910 129650 8980
rect 129850 8910 130150 8980
rect 130350 8910 130650 8980
rect 130850 8910 131150 8980
rect 131350 8910 131650 8980
rect 131850 8910 132150 8980
rect 132350 8910 132650 8980
rect 132850 8910 133150 8980
rect 133350 8910 133650 8980
rect 133850 8910 134150 8980
rect 134350 8910 134650 8980
rect 134850 8910 135150 8980
rect 135350 8910 135650 8980
rect 135850 8910 136150 8980
rect 136350 8910 136650 8980
rect 136850 8910 137150 8980
rect 137350 8910 137650 8980
rect 137850 8910 138150 8980
rect 138350 8910 138650 8980
rect 138850 8910 139150 8980
rect 139350 8910 139650 8980
rect 139850 8910 140000 8980
rect 104000 8900 140000 8910
rect 104000 8880 104120 8900
rect 104380 8880 104620 8900
rect 104880 8880 105120 8900
rect 105380 8880 105620 8900
rect 105880 8880 106120 8900
rect 106380 8880 106620 8900
rect 106880 8880 107120 8900
rect 107380 8880 107620 8900
rect 107880 8880 108120 8900
rect 108380 8880 108620 8900
rect 108880 8880 109120 8900
rect 109380 8880 109620 8900
rect 109880 8880 110120 8900
rect 110380 8880 110620 8900
rect 110880 8880 111120 8900
rect 111380 8880 111620 8900
rect 111880 8880 112120 8900
rect 112380 8880 112620 8900
rect 112880 8880 113120 8900
rect 113380 8880 113620 8900
rect 113880 8880 114120 8900
rect 114380 8880 114620 8900
rect 114880 8880 115120 8900
rect 115380 8880 115620 8900
rect 115880 8880 116120 8900
rect 116380 8880 116620 8900
rect 116880 8880 117120 8900
rect 117380 8880 117620 8900
rect 117880 8880 118120 8900
rect 118380 8880 118620 8900
rect 118880 8880 119120 8900
rect 119380 8880 119620 8900
rect 119880 8880 120120 8900
rect 120380 8880 120620 8900
rect 120880 8880 121120 8900
rect 121380 8880 121620 8900
rect 121880 8880 122120 8900
rect 122380 8880 122620 8900
rect 122880 8880 123120 8900
rect 123380 8880 123620 8900
rect 123880 8880 124120 8900
rect 124380 8880 124620 8900
rect 124880 8880 125120 8900
rect 125380 8880 125620 8900
rect 125880 8880 126120 8900
rect 126380 8880 126620 8900
rect 126880 8880 127120 8900
rect 127380 8880 127620 8900
rect 127880 8880 128120 8900
rect 128380 8880 128620 8900
rect 128880 8880 129120 8900
rect 129380 8880 129620 8900
rect 129880 8880 130120 8900
rect 130380 8880 130620 8900
rect 130880 8880 131120 8900
rect 131380 8880 131620 8900
rect 131880 8880 132120 8900
rect 132380 8880 132620 8900
rect 132880 8880 133120 8900
rect 133380 8880 133620 8900
rect 133880 8880 134120 8900
rect 134380 8880 134620 8900
rect 134880 8880 135120 8900
rect 135380 8880 135620 8900
rect 135880 8880 136120 8900
rect 136380 8880 136620 8900
rect 136880 8880 137120 8900
rect 137380 8880 137620 8900
rect 137880 8880 138120 8900
rect 138380 8880 138620 8900
rect 138880 8880 139120 8900
rect 139380 8880 139620 8900
rect 139880 8880 140000 8900
rect 104000 8620 104100 8880
rect 104400 8620 104600 8880
rect 104900 8620 105100 8880
rect 105400 8620 105600 8880
rect 105900 8620 106100 8880
rect 106400 8620 106600 8880
rect 106900 8620 107100 8880
rect 107400 8620 107600 8880
rect 107900 8620 108100 8880
rect 108400 8620 108600 8880
rect 108900 8620 109100 8880
rect 109400 8620 109600 8880
rect 109900 8620 110100 8880
rect 110400 8620 110600 8880
rect 110900 8620 111100 8880
rect 111400 8620 111600 8880
rect 111900 8620 112100 8880
rect 112400 8620 112600 8880
rect 112900 8620 113100 8880
rect 113400 8620 113600 8880
rect 113900 8620 114100 8880
rect 114400 8620 114600 8880
rect 114900 8620 115100 8880
rect 115400 8620 115600 8880
rect 115900 8620 116100 8880
rect 116400 8620 116600 8880
rect 116900 8620 117100 8880
rect 117400 8620 117600 8880
rect 117900 8620 118100 8880
rect 118400 8620 118600 8880
rect 118900 8620 119100 8880
rect 119400 8620 119600 8880
rect 119900 8620 120100 8880
rect 120400 8620 120600 8880
rect 120900 8620 121100 8880
rect 121400 8620 121600 8880
rect 121900 8620 122100 8880
rect 122400 8620 122600 8880
rect 122900 8620 123100 8880
rect 123400 8620 123600 8880
rect 123900 8620 124100 8880
rect 124400 8620 124600 8880
rect 124900 8620 125100 8880
rect 125400 8620 125600 8880
rect 125900 8620 126100 8880
rect 126400 8620 126600 8880
rect 126900 8620 127100 8880
rect 127400 8620 127600 8880
rect 127900 8850 128100 8880
rect 127900 8650 128020 8850
rect 128090 8650 128100 8850
rect 127900 8620 128100 8650
rect 128400 8850 128600 8880
rect 128400 8650 128410 8850
rect 128480 8650 128520 8850
rect 128590 8650 128600 8850
rect 128400 8620 128600 8650
rect 128900 8850 129100 8880
rect 128900 8650 128910 8850
rect 128980 8650 129020 8850
rect 129090 8650 129100 8850
rect 128900 8620 129100 8650
rect 129400 8850 129600 8880
rect 129400 8650 129410 8850
rect 129480 8650 129520 8850
rect 129590 8650 129600 8850
rect 129400 8620 129600 8650
rect 129900 8850 130100 8880
rect 129900 8650 129910 8850
rect 129980 8650 130020 8850
rect 130090 8650 130100 8850
rect 129900 8620 130100 8650
rect 130400 8850 130600 8880
rect 130400 8650 130410 8850
rect 130480 8650 130520 8850
rect 130590 8650 130600 8850
rect 130400 8620 130600 8650
rect 130900 8850 131100 8880
rect 130900 8650 130910 8850
rect 130980 8650 131020 8850
rect 131090 8650 131100 8850
rect 130900 8620 131100 8650
rect 131400 8850 131600 8880
rect 131400 8650 131410 8850
rect 131480 8650 131520 8850
rect 131590 8650 131600 8850
rect 131400 8620 131600 8650
rect 131900 8850 132100 8880
rect 131900 8650 131910 8850
rect 131980 8650 132020 8850
rect 132090 8650 132100 8850
rect 131900 8620 132100 8650
rect 132400 8850 132600 8880
rect 132400 8650 132410 8850
rect 132480 8650 132520 8850
rect 132590 8650 132600 8850
rect 132400 8620 132600 8650
rect 132900 8850 133100 8880
rect 132900 8650 132910 8850
rect 132980 8650 133020 8850
rect 133090 8650 133100 8850
rect 132900 8620 133100 8650
rect 133400 8850 133600 8880
rect 133400 8650 133410 8850
rect 133480 8650 133520 8850
rect 133590 8650 133600 8850
rect 133400 8620 133600 8650
rect 133900 8850 134100 8880
rect 133900 8650 133910 8850
rect 133980 8650 134020 8850
rect 134090 8650 134100 8850
rect 133900 8620 134100 8650
rect 134400 8850 134600 8880
rect 134400 8650 134410 8850
rect 134480 8650 134520 8850
rect 134590 8650 134600 8850
rect 134400 8620 134600 8650
rect 134900 8850 135100 8880
rect 134900 8650 134910 8850
rect 134980 8650 135020 8850
rect 135090 8650 135100 8850
rect 134900 8620 135100 8650
rect 135400 8850 135600 8880
rect 135400 8650 135410 8850
rect 135480 8650 135520 8850
rect 135590 8650 135600 8850
rect 135400 8620 135600 8650
rect 135900 8850 136100 8880
rect 135900 8650 135910 8850
rect 135980 8650 136020 8850
rect 136090 8650 136100 8850
rect 135900 8620 136100 8650
rect 136400 8850 136600 8880
rect 136400 8650 136410 8850
rect 136480 8650 136520 8850
rect 136590 8650 136600 8850
rect 136400 8620 136600 8650
rect 136900 8850 137100 8880
rect 136900 8650 136910 8850
rect 136980 8650 137020 8850
rect 137090 8650 137100 8850
rect 136900 8620 137100 8650
rect 137400 8850 137600 8880
rect 137400 8650 137410 8850
rect 137480 8650 137520 8850
rect 137590 8650 137600 8850
rect 137400 8620 137600 8650
rect 137900 8850 138100 8880
rect 137900 8650 137910 8850
rect 137980 8650 138020 8850
rect 138090 8650 138100 8850
rect 137900 8620 138100 8650
rect 138400 8850 138600 8880
rect 138400 8650 138410 8850
rect 138480 8650 138520 8850
rect 138590 8650 138600 8850
rect 138400 8620 138600 8650
rect 138900 8850 139100 8880
rect 138900 8650 138910 8850
rect 138980 8650 139020 8850
rect 139090 8650 139100 8850
rect 138900 8620 139100 8650
rect 139400 8850 139600 8880
rect 139400 8650 139410 8850
rect 139480 8650 139520 8850
rect 139590 8650 139600 8850
rect 139400 8620 139600 8650
rect 139900 8850 140000 8880
rect 139900 8650 139910 8850
rect 139980 8650 140000 8850
rect 139900 8620 140000 8650
rect 104000 8600 104120 8620
rect 104380 8600 104620 8620
rect 104880 8600 105120 8620
rect 105380 8600 105620 8620
rect 105880 8600 106120 8620
rect 106380 8600 106620 8620
rect 106880 8600 107120 8620
rect 107380 8600 107620 8620
rect 107880 8600 108120 8620
rect 108380 8600 108620 8620
rect 108880 8600 109120 8620
rect 109380 8600 109620 8620
rect 109880 8600 110120 8620
rect 110380 8600 110620 8620
rect 110880 8600 111120 8620
rect 111380 8600 111620 8620
rect 111880 8600 112120 8620
rect 112380 8600 112620 8620
rect 112880 8600 113120 8620
rect 113380 8600 113620 8620
rect 113880 8600 114120 8620
rect 114380 8600 114620 8620
rect 114880 8600 115120 8620
rect 115380 8600 115620 8620
rect 115880 8600 116120 8620
rect 116380 8600 116620 8620
rect 116880 8600 117120 8620
rect 117380 8600 117620 8620
rect 117880 8600 118120 8620
rect 118380 8600 118620 8620
rect 118880 8600 119120 8620
rect 119380 8600 119620 8620
rect 119880 8600 120120 8620
rect 120380 8600 120620 8620
rect 120880 8600 121120 8620
rect 121380 8600 121620 8620
rect 121880 8600 122120 8620
rect 122380 8600 122620 8620
rect 122880 8600 123120 8620
rect 123380 8600 123620 8620
rect 123880 8600 124120 8620
rect 124380 8600 124620 8620
rect 124880 8600 125120 8620
rect 125380 8600 125620 8620
rect 125880 8600 126120 8620
rect 126380 8600 126620 8620
rect 126880 8600 127120 8620
rect 127380 8600 127620 8620
rect 127880 8600 128120 8620
rect 128380 8600 128620 8620
rect 128880 8600 129120 8620
rect 129380 8600 129620 8620
rect 129880 8600 130120 8620
rect 130380 8600 130620 8620
rect 130880 8600 131120 8620
rect 131380 8600 131620 8620
rect 131880 8600 132120 8620
rect 132380 8600 132620 8620
rect 132880 8600 133120 8620
rect 133380 8600 133620 8620
rect 133880 8600 134120 8620
rect 134380 8600 134620 8620
rect 134880 8600 135120 8620
rect 135380 8600 135620 8620
rect 135880 8600 136120 8620
rect 136380 8600 136620 8620
rect 136880 8600 137120 8620
rect 137380 8600 137620 8620
rect 137880 8600 138120 8620
rect 138380 8600 138620 8620
rect 138880 8600 139120 8620
rect 139380 8600 139620 8620
rect 139880 8600 140000 8620
rect 104000 8590 140000 8600
rect 104000 8520 128150 8590
rect 128350 8520 128650 8590
rect 128850 8520 129150 8590
rect 129350 8520 129650 8590
rect 129850 8520 130150 8590
rect 130350 8520 130650 8590
rect 130850 8520 131150 8590
rect 131350 8520 131650 8590
rect 131850 8520 132150 8590
rect 132350 8520 132650 8590
rect 132850 8520 133150 8590
rect 133350 8520 133650 8590
rect 133850 8520 134150 8590
rect 134350 8520 134650 8590
rect 134850 8520 135150 8590
rect 135350 8520 135650 8590
rect 135850 8520 136150 8590
rect 136350 8520 136650 8590
rect 136850 8520 137150 8590
rect 137350 8520 137650 8590
rect 137850 8520 138150 8590
rect 138350 8520 138650 8590
rect 138850 8520 139150 8590
rect 139350 8520 139650 8590
rect 139850 8520 140000 8590
rect 104000 8480 140000 8520
rect 104000 8410 128150 8480
rect 128350 8410 128650 8480
rect 128850 8410 129150 8480
rect 129350 8410 129650 8480
rect 129850 8410 130150 8480
rect 130350 8410 130650 8480
rect 130850 8410 131150 8480
rect 131350 8410 131650 8480
rect 131850 8410 132150 8480
rect 132350 8410 132650 8480
rect 132850 8410 133150 8480
rect 133350 8410 133650 8480
rect 133850 8410 134150 8480
rect 134350 8410 134650 8480
rect 134850 8410 135150 8480
rect 135350 8410 135650 8480
rect 135850 8410 136150 8480
rect 136350 8410 136650 8480
rect 136850 8410 137150 8480
rect 137350 8410 137650 8480
rect 137850 8410 138150 8480
rect 138350 8410 138650 8480
rect 138850 8410 139150 8480
rect 139350 8410 139650 8480
rect 139850 8410 140000 8480
rect 104000 8400 140000 8410
rect 104000 8380 104120 8400
rect 104380 8380 104620 8400
rect 104880 8380 105120 8400
rect 105380 8380 105620 8400
rect 105880 8380 106120 8400
rect 106380 8380 106620 8400
rect 106880 8380 107120 8400
rect 107380 8380 107620 8400
rect 107880 8380 108120 8400
rect 108380 8380 108620 8400
rect 108880 8380 109120 8400
rect 109380 8380 109620 8400
rect 109880 8380 110120 8400
rect 110380 8380 110620 8400
rect 110880 8380 111120 8400
rect 111380 8380 111620 8400
rect 111880 8380 112120 8400
rect 112380 8380 112620 8400
rect 112880 8380 113120 8400
rect 113380 8380 113620 8400
rect 113880 8380 114120 8400
rect 114380 8380 114620 8400
rect 114880 8380 115120 8400
rect 115380 8380 115620 8400
rect 115880 8380 116120 8400
rect 116380 8380 116620 8400
rect 116880 8380 117120 8400
rect 117380 8380 117620 8400
rect 117880 8380 118120 8400
rect 118380 8380 118620 8400
rect 118880 8380 119120 8400
rect 119380 8380 119620 8400
rect 119880 8380 120120 8400
rect 120380 8380 120620 8400
rect 120880 8380 121120 8400
rect 121380 8380 121620 8400
rect 121880 8380 122120 8400
rect 122380 8380 122620 8400
rect 122880 8380 123120 8400
rect 123380 8380 123620 8400
rect 123880 8380 124120 8400
rect 124380 8380 124620 8400
rect 124880 8380 125120 8400
rect 125380 8380 125620 8400
rect 125880 8380 126120 8400
rect 126380 8380 126620 8400
rect 126880 8380 127120 8400
rect 127380 8380 127620 8400
rect 127880 8380 128120 8400
rect 128380 8380 128620 8400
rect 128880 8380 129120 8400
rect 129380 8380 129620 8400
rect 129880 8380 130120 8400
rect 130380 8380 130620 8400
rect 130880 8380 131120 8400
rect 131380 8380 131620 8400
rect 131880 8380 132120 8400
rect 132380 8380 132620 8400
rect 132880 8380 133120 8400
rect 133380 8380 133620 8400
rect 133880 8380 134120 8400
rect 134380 8380 134620 8400
rect 134880 8380 135120 8400
rect 135380 8380 135620 8400
rect 135880 8380 136120 8400
rect 136380 8380 136620 8400
rect 136880 8380 137120 8400
rect 137380 8380 137620 8400
rect 137880 8380 138120 8400
rect 138380 8380 138620 8400
rect 138880 8380 139120 8400
rect 139380 8380 139620 8400
rect 139880 8380 140000 8400
rect 104000 8120 104100 8380
rect 104400 8120 104600 8380
rect 104900 8120 105100 8380
rect 105400 8120 105600 8380
rect 105900 8120 106100 8380
rect 106400 8120 106600 8380
rect 106900 8120 107100 8380
rect 107400 8120 107600 8380
rect 107900 8120 108100 8380
rect 108400 8120 108600 8380
rect 108900 8120 109100 8380
rect 109400 8120 109600 8380
rect 109900 8120 110100 8380
rect 110400 8120 110600 8380
rect 110900 8120 111100 8380
rect 111400 8120 111600 8380
rect 111900 8120 112100 8380
rect 112400 8120 112600 8380
rect 112900 8120 113100 8380
rect 113400 8120 113600 8380
rect 113900 8120 114100 8380
rect 114400 8120 114600 8380
rect 114900 8120 115100 8380
rect 115400 8120 115600 8380
rect 115900 8120 116100 8380
rect 116400 8120 116600 8380
rect 116900 8120 117100 8380
rect 117400 8120 117600 8380
rect 117900 8120 118100 8380
rect 118400 8120 118600 8380
rect 118900 8120 119100 8380
rect 119400 8120 119600 8380
rect 119900 8120 120100 8380
rect 120400 8120 120600 8380
rect 120900 8120 121100 8380
rect 121400 8120 121600 8380
rect 121900 8120 122100 8380
rect 122400 8120 122600 8380
rect 122900 8120 123100 8380
rect 123400 8120 123600 8380
rect 123900 8120 124100 8380
rect 124400 8120 124600 8380
rect 124900 8120 125100 8380
rect 125400 8120 125600 8380
rect 125900 8120 126100 8380
rect 126400 8120 126600 8380
rect 126900 8120 127100 8380
rect 127400 8120 127600 8380
rect 127900 8350 128100 8380
rect 127900 8150 128020 8350
rect 128090 8150 128100 8350
rect 127900 8120 128100 8150
rect 128400 8350 128600 8380
rect 128400 8150 128410 8350
rect 128480 8150 128520 8350
rect 128590 8150 128600 8350
rect 128400 8120 128600 8150
rect 128900 8350 129100 8380
rect 128900 8150 128910 8350
rect 128980 8150 129020 8350
rect 129090 8150 129100 8350
rect 128900 8120 129100 8150
rect 129400 8350 129600 8380
rect 129400 8150 129410 8350
rect 129480 8150 129520 8350
rect 129590 8150 129600 8350
rect 129400 8120 129600 8150
rect 129900 8350 130100 8380
rect 129900 8150 129910 8350
rect 129980 8150 130020 8350
rect 130090 8150 130100 8350
rect 129900 8120 130100 8150
rect 130400 8350 130600 8380
rect 130400 8150 130410 8350
rect 130480 8150 130520 8350
rect 130590 8150 130600 8350
rect 130400 8120 130600 8150
rect 130900 8350 131100 8380
rect 130900 8150 130910 8350
rect 130980 8150 131020 8350
rect 131090 8150 131100 8350
rect 130900 8120 131100 8150
rect 131400 8350 131600 8380
rect 131400 8150 131410 8350
rect 131480 8150 131520 8350
rect 131590 8150 131600 8350
rect 131400 8120 131600 8150
rect 131900 8350 132100 8380
rect 131900 8150 131910 8350
rect 131980 8150 132020 8350
rect 132090 8150 132100 8350
rect 131900 8120 132100 8150
rect 132400 8350 132600 8380
rect 132400 8150 132410 8350
rect 132480 8150 132520 8350
rect 132590 8150 132600 8350
rect 132400 8120 132600 8150
rect 132900 8350 133100 8380
rect 132900 8150 132910 8350
rect 132980 8150 133020 8350
rect 133090 8150 133100 8350
rect 132900 8120 133100 8150
rect 133400 8350 133600 8380
rect 133400 8150 133410 8350
rect 133480 8150 133520 8350
rect 133590 8150 133600 8350
rect 133400 8120 133600 8150
rect 133900 8350 134100 8380
rect 133900 8150 133910 8350
rect 133980 8150 134020 8350
rect 134090 8150 134100 8350
rect 133900 8120 134100 8150
rect 134400 8350 134600 8380
rect 134400 8150 134410 8350
rect 134480 8150 134520 8350
rect 134590 8150 134600 8350
rect 134400 8120 134600 8150
rect 134900 8350 135100 8380
rect 134900 8150 134910 8350
rect 134980 8150 135020 8350
rect 135090 8150 135100 8350
rect 134900 8120 135100 8150
rect 135400 8350 135600 8380
rect 135400 8150 135410 8350
rect 135480 8150 135520 8350
rect 135590 8150 135600 8350
rect 135400 8120 135600 8150
rect 135900 8350 136100 8380
rect 135900 8150 135910 8350
rect 135980 8150 136020 8350
rect 136090 8150 136100 8350
rect 135900 8120 136100 8150
rect 136400 8350 136600 8380
rect 136400 8150 136410 8350
rect 136480 8150 136520 8350
rect 136590 8150 136600 8350
rect 136400 8120 136600 8150
rect 136900 8350 137100 8380
rect 136900 8150 136910 8350
rect 136980 8150 137020 8350
rect 137090 8150 137100 8350
rect 136900 8120 137100 8150
rect 137400 8350 137600 8380
rect 137400 8150 137410 8350
rect 137480 8150 137520 8350
rect 137590 8150 137600 8350
rect 137400 8120 137600 8150
rect 137900 8350 138100 8380
rect 137900 8150 137910 8350
rect 137980 8150 138020 8350
rect 138090 8150 138100 8350
rect 137900 8120 138100 8150
rect 138400 8350 138600 8380
rect 138400 8150 138410 8350
rect 138480 8150 138520 8350
rect 138590 8150 138600 8350
rect 138400 8120 138600 8150
rect 138900 8350 139100 8380
rect 138900 8150 138910 8350
rect 138980 8150 139020 8350
rect 139090 8150 139100 8350
rect 138900 8120 139100 8150
rect 139400 8350 139600 8380
rect 139400 8150 139410 8350
rect 139480 8150 139520 8350
rect 139590 8150 139600 8350
rect 139400 8120 139600 8150
rect 139900 8350 140000 8380
rect 139900 8150 139910 8350
rect 139980 8150 140000 8350
rect 139900 8120 140000 8150
rect 104000 8100 104120 8120
rect 104380 8100 104620 8120
rect 104880 8100 105120 8120
rect 105380 8100 105620 8120
rect 105880 8100 106120 8120
rect 106380 8100 106620 8120
rect 106880 8100 107120 8120
rect 107380 8100 107620 8120
rect 107880 8100 108120 8120
rect 108380 8100 108620 8120
rect 108880 8100 109120 8120
rect 109380 8100 109620 8120
rect 109880 8100 110120 8120
rect 110380 8100 110620 8120
rect 110880 8100 111120 8120
rect 111380 8100 111620 8120
rect 111880 8100 112120 8120
rect 112380 8100 112620 8120
rect 112880 8100 113120 8120
rect 113380 8100 113620 8120
rect 113880 8100 114120 8120
rect 114380 8100 114620 8120
rect 114880 8100 115120 8120
rect 115380 8100 115620 8120
rect 115880 8100 116120 8120
rect 116380 8100 116620 8120
rect 116880 8100 117120 8120
rect 117380 8100 117620 8120
rect 117880 8100 118120 8120
rect 118380 8100 118620 8120
rect 118880 8100 119120 8120
rect 119380 8100 119620 8120
rect 119880 8100 120120 8120
rect 120380 8100 120620 8120
rect 120880 8100 121120 8120
rect 121380 8100 121620 8120
rect 121880 8100 122120 8120
rect 122380 8100 122620 8120
rect 122880 8100 123120 8120
rect 123380 8100 123620 8120
rect 123880 8100 124120 8120
rect 124380 8100 124620 8120
rect 124880 8100 125120 8120
rect 125380 8100 125620 8120
rect 125880 8100 126120 8120
rect 126380 8100 126620 8120
rect 126880 8100 127120 8120
rect 127380 8100 127620 8120
rect 127880 8100 128120 8120
rect 128380 8100 128620 8120
rect 128880 8100 129120 8120
rect 129380 8100 129620 8120
rect 129880 8100 130120 8120
rect 130380 8100 130620 8120
rect 130880 8100 131120 8120
rect 131380 8100 131620 8120
rect 131880 8100 132120 8120
rect 132380 8100 132620 8120
rect 132880 8100 133120 8120
rect 133380 8100 133620 8120
rect 133880 8100 134120 8120
rect 134380 8100 134620 8120
rect 134880 8100 135120 8120
rect 135380 8100 135620 8120
rect 135880 8100 136120 8120
rect 136380 8100 136620 8120
rect 136880 8100 137120 8120
rect 137380 8100 137620 8120
rect 137880 8100 138120 8120
rect 138380 8100 138620 8120
rect 138880 8100 139120 8120
rect 139380 8100 139620 8120
rect 139880 8100 140000 8120
rect 104000 8090 140000 8100
rect 104000 8020 128150 8090
rect 128350 8020 128650 8090
rect 128850 8020 129150 8090
rect 129350 8020 129650 8090
rect 129850 8020 130150 8090
rect 130350 8020 130650 8090
rect 130850 8020 131150 8090
rect 131350 8020 131650 8090
rect 131850 8020 132150 8090
rect 132350 8020 132650 8090
rect 132850 8020 133150 8090
rect 133350 8020 133650 8090
rect 133850 8020 134150 8090
rect 134350 8020 134650 8090
rect 134850 8020 135150 8090
rect 135350 8020 135650 8090
rect 135850 8020 136150 8090
rect 136350 8020 136650 8090
rect 136850 8020 137150 8090
rect 137350 8020 137650 8090
rect 137850 8020 138150 8090
rect 138350 8020 138650 8090
rect 138850 8020 139150 8090
rect 139350 8020 139650 8090
rect 139850 8020 140000 8090
rect 104000 7980 140000 8020
rect 104000 7910 128150 7980
rect 128350 7910 128650 7980
rect 128850 7910 129150 7980
rect 129350 7910 129650 7980
rect 129850 7910 130150 7980
rect 130350 7910 130650 7980
rect 130850 7910 131150 7980
rect 131350 7910 131650 7980
rect 131850 7910 132150 7980
rect 132350 7910 132650 7980
rect 132850 7910 133150 7980
rect 133350 7910 133650 7980
rect 133850 7910 134150 7980
rect 134350 7910 134650 7980
rect 134850 7910 135150 7980
rect 135350 7910 135650 7980
rect 135850 7910 136150 7980
rect 136350 7910 136650 7980
rect 136850 7910 137150 7980
rect 137350 7910 137650 7980
rect 137850 7910 138150 7980
rect 138350 7910 138650 7980
rect 138850 7910 139150 7980
rect 139350 7910 139650 7980
rect 139850 7910 140000 7980
rect 104000 7900 140000 7910
rect 104000 7880 104120 7900
rect 104380 7880 104620 7900
rect 104880 7880 105120 7900
rect 105380 7880 105620 7900
rect 105880 7880 106120 7900
rect 106380 7880 106620 7900
rect 106880 7880 107120 7900
rect 107380 7880 107620 7900
rect 107880 7880 108120 7900
rect 108380 7880 108620 7900
rect 108880 7880 109120 7900
rect 109380 7880 109620 7900
rect 109880 7880 110120 7900
rect 110380 7880 110620 7900
rect 110880 7880 111120 7900
rect 111380 7880 111620 7900
rect 111880 7880 112120 7900
rect 112380 7880 112620 7900
rect 112880 7880 113120 7900
rect 113380 7880 113620 7900
rect 113880 7880 114120 7900
rect 114380 7880 114620 7900
rect 114880 7880 115120 7900
rect 115380 7880 115620 7900
rect 115880 7880 116120 7900
rect 116380 7880 116620 7900
rect 116880 7880 117120 7900
rect 117380 7880 117620 7900
rect 117880 7880 118120 7900
rect 118380 7880 118620 7900
rect 118880 7880 119120 7900
rect 119380 7880 119620 7900
rect 119880 7880 120120 7900
rect 120380 7880 120620 7900
rect 120880 7880 121120 7900
rect 121380 7880 121620 7900
rect 121880 7880 122120 7900
rect 122380 7880 122620 7900
rect 122880 7880 123120 7900
rect 123380 7880 123620 7900
rect 123880 7880 124120 7900
rect 124380 7880 124620 7900
rect 124880 7880 125120 7900
rect 125380 7880 125620 7900
rect 125880 7880 126120 7900
rect 126380 7880 126620 7900
rect 126880 7880 127120 7900
rect 127380 7880 127620 7900
rect 127880 7880 128120 7900
rect 128380 7880 128620 7900
rect 128880 7880 129120 7900
rect 129380 7880 129620 7900
rect 129880 7880 130120 7900
rect 130380 7880 130620 7900
rect 130880 7880 131120 7900
rect 131380 7880 131620 7900
rect 131880 7880 132120 7900
rect 132380 7880 132620 7900
rect 132880 7880 133120 7900
rect 133380 7880 133620 7900
rect 133880 7880 134120 7900
rect 134380 7880 134620 7900
rect 134880 7880 135120 7900
rect 135380 7880 135620 7900
rect 135880 7880 136120 7900
rect 136380 7880 136620 7900
rect 136880 7880 137120 7900
rect 137380 7880 137620 7900
rect 137880 7880 138120 7900
rect 138380 7880 138620 7900
rect 138880 7880 139120 7900
rect 139380 7880 139620 7900
rect 139880 7880 140000 7900
rect 104000 7620 104100 7880
rect 104400 7620 104600 7880
rect 104900 7620 105100 7880
rect 105400 7620 105600 7880
rect 105900 7620 106100 7880
rect 106400 7620 106600 7880
rect 106900 7620 107100 7880
rect 107400 7620 107600 7880
rect 107900 7620 108100 7880
rect 108400 7620 108600 7880
rect 108900 7620 109100 7880
rect 109400 7620 109600 7880
rect 109900 7620 110100 7880
rect 110400 7620 110600 7880
rect 110900 7620 111100 7880
rect 111400 7620 111600 7880
rect 111900 7620 112100 7880
rect 112400 7620 112600 7880
rect 112900 7620 113100 7880
rect 113400 7620 113600 7880
rect 113900 7620 114100 7880
rect 114400 7620 114600 7880
rect 114900 7620 115100 7880
rect 115400 7620 115600 7880
rect 115900 7620 116100 7880
rect 116400 7620 116600 7880
rect 116900 7620 117100 7880
rect 117400 7620 117600 7880
rect 117900 7620 118100 7880
rect 118400 7620 118600 7880
rect 118900 7620 119100 7880
rect 119400 7620 119600 7880
rect 119900 7620 120100 7880
rect 120400 7620 120600 7880
rect 120900 7620 121100 7880
rect 121400 7620 121600 7880
rect 121900 7620 122100 7880
rect 122400 7620 122600 7880
rect 122900 7620 123100 7880
rect 123400 7620 123600 7880
rect 123900 7620 124100 7880
rect 124400 7620 124600 7880
rect 124900 7620 125100 7880
rect 125400 7620 125600 7880
rect 125900 7620 126100 7880
rect 126400 7620 126600 7880
rect 126900 7620 127100 7880
rect 127400 7620 127600 7880
rect 127900 7850 128100 7880
rect 127900 7650 128020 7850
rect 128090 7650 128100 7850
rect 127900 7620 128100 7650
rect 128400 7850 128600 7880
rect 128400 7650 128410 7850
rect 128480 7650 128520 7850
rect 128590 7650 128600 7850
rect 128400 7620 128600 7650
rect 128900 7850 129100 7880
rect 128900 7650 128910 7850
rect 128980 7650 129020 7850
rect 129090 7650 129100 7850
rect 128900 7620 129100 7650
rect 129400 7850 129600 7880
rect 129400 7650 129410 7850
rect 129480 7650 129520 7850
rect 129590 7650 129600 7850
rect 129400 7620 129600 7650
rect 129900 7850 130100 7880
rect 129900 7650 129910 7850
rect 129980 7650 130020 7850
rect 130090 7650 130100 7850
rect 129900 7620 130100 7650
rect 130400 7850 130600 7880
rect 130400 7650 130410 7850
rect 130480 7650 130520 7850
rect 130590 7650 130600 7850
rect 130400 7620 130600 7650
rect 130900 7850 131100 7880
rect 130900 7650 130910 7850
rect 130980 7650 131020 7850
rect 131090 7650 131100 7850
rect 130900 7620 131100 7650
rect 131400 7850 131600 7880
rect 131400 7650 131410 7850
rect 131480 7650 131520 7850
rect 131590 7650 131600 7850
rect 131400 7620 131600 7650
rect 131900 7850 132100 7880
rect 131900 7650 131910 7850
rect 131980 7650 132020 7850
rect 132090 7650 132100 7850
rect 131900 7620 132100 7650
rect 132400 7850 132600 7880
rect 132400 7650 132410 7850
rect 132480 7650 132520 7850
rect 132590 7650 132600 7850
rect 132400 7620 132600 7650
rect 132900 7850 133100 7880
rect 132900 7650 132910 7850
rect 132980 7650 133020 7850
rect 133090 7650 133100 7850
rect 132900 7620 133100 7650
rect 133400 7850 133600 7880
rect 133400 7650 133410 7850
rect 133480 7650 133520 7850
rect 133590 7650 133600 7850
rect 133400 7620 133600 7650
rect 133900 7850 134100 7880
rect 133900 7650 133910 7850
rect 133980 7650 134020 7850
rect 134090 7650 134100 7850
rect 133900 7620 134100 7650
rect 134400 7850 134600 7880
rect 134400 7650 134410 7850
rect 134480 7650 134520 7850
rect 134590 7650 134600 7850
rect 134400 7620 134600 7650
rect 134900 7850 135100 7880
rect 134900 7650 134910 7850
rect 134980 7650 135020 7850
rect 135090 7650 135100 7850
rect 134900 7620 135100 7650
rect 135400 7850 135600 7880
rect 135400 7650 135410 7850
rect 135480 7650 135520 7850
rect 135590 7650 135600 7850
rect 135400 7620 135600 7650
rect 135900 7850 136100 7880
rect 135900 7650 135910 7850
rect 135980 7650 136020 7850
rect 136090 7650 136100 7850
rect 135900 7620 136100 7650
rect 136400 7850 136600 7880
rect 136400 7650 136410 7850
rect 136480 7650 136520 7850
rect 136590 7650 136600 7850
rect 136400 7620 136600 7650
rect 136900 7850 137100 7880
rect 136900 7650 136910 7850
rect 136980 7650 137020 7850
rect 137090 7650 137100 7850
rect 136900 7620 137100 7650
rect 137400 7850 137600 7880
rect 137400 7650 137410 7850
rect 137480 7650 137520 7850
rect 137590 7650 137600 7850
rect 137400 7620 137600 7650
rect 137900 7850 138100 7880
rect 137900 7650 137910 7850
rect 137980 7650 138020 7850
rect 138090 7650 138100 7850
rect 137900 7620 138100 7650
rect 138400 7850 138600 7880
rect 138400 7650 138410 7850
rect 138480 7650 138520 7850
rect 138590 7650 138600 7850
rect 138400 7620 138600 7650
rect 138900 7850 139100 7880
rect 138900 7650 138910 7850
rect 138980 7650 139020 7850
rect 139090 7650 139100 7850
rect 138900 7620 139100 7650
rect 139400 7850 139600 7880
rect 139400 7650 139410 7850
rect 139480 7650 139520 7850
rect 139590 7650 139600 7850
rect 139400 7620 139600 7650
rect 139900 7850 140000 7880
rect 139900 7650 139910 7850
rect 139980 7650 140000 7850
rect 139900 7620 140000 7650
rect 104000 7600 104120 7620
rect 104380 7600 104620 7620
rect 104880 7600 105120 7620
rect 105380 7600 105620 7620
rect 105880 7600 106120 7620
rect 106380 7600 106620 7620
rect 106880 7600 107120 7620
rect 107380 7600 107620 7620
rect 107880 7600 108120 7620
rect 108380 7600 108620 7620
rect 108880 7600 109120 7620
rect 109380 7600 109620 7620
rect 109880 7600 110120 7620
rect 110380 7600 110620 7620
rect 110880 7600 111120 7620
rect 111380 7600 111620 7620
rect 111880 7600 112120 7620
rect 112380 7600 112620 7620
rect 112880 7600 113120 7620
rect 113380 7600 113620 7620
rect 113880 7600 114120 7620
rect 114380 7600 114620 7620
rect 114880 7600 115120 7620
rect 115380 7600 115620 7620
rect 115880 7600 116120 7620
rect 116380 7600 116620 7620
rect 116880 7600 117120 7620
rect 117380 7600 117620 7620
rect 117880 7600 118120 7620
rect 118380 7600 118620 7620
rect 118880 7600 119120 7620
rect 119380 7600 119620 7620
rect 119880 7600 120120 7620
rect 120380 7600 120620 7620
rect 120880 7600 121120 7620
rect 121380 7600 121620 7620
rect 121880 7600 122120 7620
rect 122380 7600 122620 7620
rect 122880 7600 123120 7620
rect 123380 7600 123620 7620
rect 123880 7600 124120 7620
rect 124380 7600 124620 7620
rect 124880 7600 125120 7620
rect 125380 7600 125620 7620
rect 125880 7600 126120 7620
rect 126380 7600 126620 7620
rect 126880 7600 127120 7620
rect 127380 7600 127620 7620
rect 127880 7600 128120 7620
rect 128380 7600 128620 7620
rect 128880 7600 129120 7620
rect 129380 7600 129620 7620
rect 129880 7600 130120 7620
rect 130380 7600 130620 7620
rect 130880 7600 131120 7620
rect 131380 7600 131620 7620
rect 131880 7600 132120 7620
rect 132380 7600 132620 7620
rect 132880 7600 133120 7620
rect 133380 7600 133620 7620
rect 133880 7600 134120 7620
rect 134380 7600 134620 7620
rect 134880 7600 135120 7620
rect 135380 7600 135620 7620
rect 135880 7600 136120 7620
rect 136380 7600 136620 7620
rect 136880 7600 137120 7620
rect 137380 7600 137620 7620
rect 137880 7600 138120 7620
rect 138380 7600 138620 7620
rect 138880 7600 139120 7620
rect 139380 7600 139620 7620
rect 139880 7600 140000 7620
rect 104000 7590 140000 7600
rect 104000 7520 128150 7590
rect 128350 7520 128650 7590
rect 128850 7520 129150 7590
rect 129350 7520 129650 7590
rect 129850 7520 130150 7590
rect 130350 7520 130650 7590
rect 130850 7520 131150 7590
rect 131350 7520 131650 7590
rect 131850 7520 132150 7590
rect 132350 7520 132650 7590
rect 132850 7520 133150 7590
rect 133350 7520 133650 7590
rect 133850 7520 134150 7590
rect 134350 7520 134650 7590
rect 134850 7520 135150 7590
rect 135350 7520 135650 7590
rect 135850 7520 136150 7590
rect 136350 7520 136650 7590
rect 136850 7520 137150 7590
rect 137350 7520 137650 7590
rect 137850 7520 138150 7590
rect 138350 7520 138650 7590
rect 138850 7520 139150 7590
rect 139350 7520 139650 7590
rect 139850 7520 140000 7590
rect 104000 7480 140000 7520
rect 104000 7410 128150 7480
rect 128350 7410 128650 7480
rect 128850 7410 129150 7480
rect 129350 7410 129650 7480
rect 129850 7410 130150 7480
rect 130350 7410 130650 7480
rect 130850 7410 131150 7480
rect 131350 7410 131650 7480
rect 131850 7410 132150 7480
rect 132350 7410 132650 7480
rect 132850 7410 133150 7480
rect 133350 7410 133650 7480
rect 133850 7410 134150 7480
rect 134350 7410 134650 7480
rect 134850 7410 135150 7480
rect 135350 7410 135650 7480
rect 135850 7410 136150 7480
rect 136350 7410 136650 7480
rect 136850 7410 137150 7480
rect 137350 7410 137650 7480
rect 137850 7410 138150 7480
rect 138350 7410 138650 7480
rect 138850 7410 139150 7480
rect 139350 7410 139650 7480
rect 139850 7410 140000 7480
rect 104000 7400 140000 7410
rect 104000 7380 104120 7400
rect 104380 7380 104620 7400
rect 104880 7380 105120 7400
rect 105380 7380 105620 7400
rect 105880 7380 106120 7400
rect 106380 7380 106620 7400
rect 106880 7380 107120 7400
rect 107380 7380 107620 7400
rect 107880 7380 108120 7400
rect 108380 7380 108620 7400
rect 108880 7380 109120 7400
rect 109380 7380 109620 7400
rect 109880 7380 110120 7400
rect 110380 7380 110620 7400
rect 110880 7380 111120 7400
rect 111380 7380 111620 7400
rect 111880 7380 112120 7400
rect 112380 7380 112620 7400
rect 112880 7380 113120 7400
rect 113380 7380 113620 7400
rect 113880 7380 114120 7400
rect 114380 7380 114620 7400
rect 114880 7380 115120 7400
rect 115380 7380 115620 7400
rect 115880 7380 116120 7400
rect 116380 7380 116620 7400
rect 116880 7380 117120 7400
rect 117380 7380 117620 7400
rect 117880 7380 118120 7400
rect 118380 7380 118620 7400
rect 118880 7380 119120 7400
rect 119380 7380 119620 7400
rect 119880 7380 120120 7400
rect 120380 7380 120620 7400
rect 120880 7380 121120 7400
rect 121380 7380 121620 7400
rect 121880 7380 122120 7400
rect 122380 7380 122620 7400
rect 122880 7380 123120 7400
rect 123380 7380 123620 7400
rect 123880 7380 124120 7400
rect 124380 7380 124620 7400
rect 124880 7380 125120 7400
rect 125380 7380 125620 7400
rect 125880 7380 126120 7400
rect 126380 7380 126620 7400
rect 126880 7380 127120 7400
rect 127380 7380 127620 7400
rect 127880 7380 128120 7400
rect 128380 7380 128620 7400
rect 128880 7380 129120 7400
rect 129380 7380 129620 7400
rect 129880 7380 130120 7400
rect 130380 7380 130620 7400
rect 130880 7380 131120 7400
rect 131380 7380 131620 7400
rect 131880 7380 132120 7400
rect 132380 7380 132620 7400
rect 132880 7380 133120 7400
rect 133380 7380 133620 7400
rect 133880 7380 134120 7400
rect 134380 7380 134620 7400
rect 134880 7380 135120 7400
rect 135380 7380 135620 7400
rect 135880 7380 136120 7400
rect 136380 7380 136620 7400
rect 136880 7380 137120 7400
rect 137380 7380 137620 7400
rect 137880 7380 138120 7400
rect 138380 7380 138620 7400
rect 138880 7380 139120 7400
rect 139380 7380 139620 7400
rect 139880 7380 140000 7400
rect 104000 7120 104100 7380
rect 104400 7120 104600 7380
rect 104900 7120 105100 7380
rect 105400 7120 105600 7380
rect 105900 7120 106100 7380
rect 106400 7120 106600 7380
rect 106900 7120 107100 7380
rect 107400 7120 107600 7380
rect 107900 7120 108100 7380
rect 108400 7120 108600 7380
rect 108900 7120 109100 7380
rect 109400 7120 109600 7380
rect 109900 7120 110100 7380
rect 110400 7120 110600 7380
rect 110900 7120 111100 7380
rect 111400 7120 111600 7380
rect 111900 7120 112100 7380
rect 112400 7120 112600 7380
rect 112900 7120 113100 7380
rect 113400 7120 113600 7380
rect 113900 7120 114100 7380
rect 114400 7120 114600 7380
rect 114900 7120 115100 7380
rect 115400 7120 115600 7380
rect 115900 7120 116100 7380
rect 116400 7120 116600 7380
rect 116900 7120 117100 7380
rect 117400 7120 117600 7380
rect 117900 7120 118100 7380
rect 118400 7120 118600 7380
rect 118900 7120 119100 7380
rect 119400 7120 119600 7380
rect 119900 7120 120100 7380
rect 120400 7120 120600 7380
rect 120900 7120 121100 7380
rect 121400 7120 121600 7380
rect 121900 7120 122100 7380
rect 122400 7120 122600 7380
rect 122900 7120 123100 7380
rect 123400 7120 123600 7380
rect 123900 7120 124100 7380
rect 124400 7120 124600 7380
rect 124900 7120 125100 7380
rect 125400 7120 125600 7380
rect 125900 7120 126100 7380
rect 126400 7120 126600 7380
rect 126900 7120 127100 7380
rect 127400 7120 127600 7380
rect 127900 7350 128100 7380
rect 127900 7150 128020 7350
rect 128090 7150 128100 7350
rect 127900 7120 128100 7150
rect 128400 7350 128600 7380
rect 128400 7150 128410 7350
rect 128480 7150 128520 7350
rect 128590 7150 128600 7350
rect 128400 7120 128600 7150
rect 128900 7350 129100 7380
rect 128900 7150 128910 7350
rect 128980 7150 129020 7350
rect 129090 7150 129100 7350
rect 128900 7120 129100 7150
rect 129400 7350 129600 7380
rect 129400 7150 129410 7350
rect 129480 7150 129520 7350
rect 129590 7150 129600 7350
rect 129400 7120 129600 7150
rect 129900 7350 130100 7380
rect 129900 7150 129910 7350
rect 129980 7150 130020 7350
rect 130090 7150 130100 7350
rect 129900 7120 130100 7150
rect 130400 7350 130600 7380
rect 130400 7150 130410 7350
rect 130480 7150 130520 7350
rect 130590 7150 130600 7350
rect 130400 7120 130600 7150
rect 130900 7350 131100 7380
rect 130900 7150 130910 7350
rect 130980 7150 131020 7350
rect 131090 7150 131100 7350
rect 130900 7120 131100 7150
rect 131400 7350 131600 7380
rect 131400 7150 131410 7350
rect 131480 7150 131520 7350
rect 131590 7150 131600 7350
rect 131400 7120 131600 7150
rect 131900 7350 132100 7380
rect 131900 7150 131910 7350
rect 131980 7150 132020 7350
rect 132090 7150 132100 7350
rect 131900 7120 132100 7150
rect 132400 7350 132600 7380
rect 132400 7150 132410 7350
rect 132480 7150 132520 7350
rect 132590 7150 132600 7350
rect 132400 7120 132600 7150
rect 132900 7350 133100 7380
rect 132900 7150 132910 7350
rect 132980 7150 133020 7350
rect 133090 7150 133100 7350
rect 132900 7120 133100 7150
rect 133400 7350 133600 7380
rect 133400 7150 133410 7350
rect 133480 7150 133520 7350
rect 133590 7150 133600 7350
rect 133400 7120 133600 7150
rect 133900 7350 134100 7380
rect 133900 7150 133910 7350
rect 133980 7150 134020 7350
rect 134090 7150 134100 7350
rect 133900 7120 134100 7150
rect 134400 7350 134600 7380
rect 134400 7150 134410 7350
rect 134480 7150 134520 7350
rect 134590 7150 134600 7350
rect 134400 7120 134600 7150
rect 134900 7350 135100 7380
rect 134900 7150 134910 7350
rect 134980 7150 135020 7350
rect 135090 7150 135100 7350
rect 134900 7120 135100 7150
rect 135400 7350 135600 7380
rect 135400 7150 135410 7350
rect 135480 7150 135520 7350
rect 135590 7150 135600 7350
rect 135400 7120 135600 7150
rect 135900 7350 136100 7380
rect 135900 7150 135910 7350
rect 135980 7150 136020 7350
rect 136090 7150 136100 7350
rect 135900 7120 136100 7150
rect 136400 7350 136600 7380
rect 136400 7150 136410 7350
rect 136480 7150 136520 7350
rect 136590 7150 136600 7350
rect 136400 7120 136600 7150
rect 136900 7350 137100 7380
rect 136900 7150 136910 7350
rect 136980 7150 137020 7350
rect 137090 7150 137100 7350
rect 136900 7120 137100 7150
rect 137400 7350 137600 7380
rect 137400 7150 137410 7350
rect 137480 7150 137520 7350
rect 137590 7150 137600 7350
rect 137400 7120 137600 7150
rect 137900 7350 138100 7380
rect 137900 7150 137910 7350
rect 137980 7150 138020 7350
rect 138090 7150 138100 7350
rect 137900 7120 138100 7150
rect 138400 7350 138600 7380
rect 138400 7150 138410 7350
rect 138480 7150 138520 7350
rect 138590 7150 138600 7350
rect 138400 7120 138600 7150
rect 138900 7350 139100 7380
rect 138900 7150 138910 7350
rect 138980 7150 139020 7350
rect 139090 7150 139100 7350
rect 138900 7120 139100 7150
rect 139400 7350 139600 7380
rect 139400 7150 139410 7350
rect 139480 7150 139520 7350
rect 139590 7150 139600 7350
rect 139400 7120 139600 7150
rect 139900 7350 140000 7380
rect 139900 7150 139910 7350
rect 139980 7150 140000 7350
rect 139900 7120 140000 7150
rect 104000 7100 104120 7120
rect 104380 7100 104620 7120
rect 104880 7100 105120 7120
rect 105380 7100 105620 7120
rect 105880 7100 106120 7120
rect 106380 7100 106620 7120
rect 106880 7100 107120 7120
rect 107380 7100 107620 7120
rect 107880 7100 108120 7120
rect 108380 7100 108620 7120
rect 108880 7100 109120 7120
rect 109380 7100 109620 7120
rect 109880 7100 110120 7120
rect 110380 7100 110620 7120
rect 110880 7100 111120 7120
rect 111380 7100 111620 7120
rect 111880 7100 112120 7120
rect 112380 7100 112620 7120
rect 112880 7100 113120 7120
rect 113380 7100 113620 7120
rect 113880 7100 114120 7120
rect 114380 7100 114620 7120
rect 114880 7100 115120 7120
rect 115380 7100 115620 7120
rect 115880 7100 116120 7120
rect 116380 7100 116620 7120
rect 116880 7100 117120 7120
rect 117380 7100 117620 7120
rect 117880 7100 118120 7120
rect 118380 7100 118620 7120
rect 118880 7100 119120 7120
rect 119380 7100 119620 7120
rect 119880 7100 120120 7120
rect 120380 7100 120620 7120
rect 120880 7100 121120 7120
rect 121380 7100 121620 7120
rect 121880 7100 122120 7120
rect 122380 7100 122620 7120
rect 122880 7100 123120 7120
rect 123380 7100 123620 7120
rect 123880 7100 124120 7120
rect 124380 7100 124620 7120
rect 124880 7100 125120 7120
rect 125380 7100 125620 7120
rect 125880 7100 126120 7120
rect 126380 7100 126620 7120
rect 126880 7100 127120 7120
rect 127380 7100 127620 7120
rect 127880 7100 128120 7120
rect 128380 7100 128620 7120
rect 128880 7100 129120 7120
rect 129380 7100 129620 7120
rect 129880 7100 130120 7120
rect 130380 7100 130620 7120
rect 130880 7100 131120 7120
rect 131380 7100 131620 7120
rect 131880 7100 132120 7120
rect 132380 7100 132620 7120
rect 132880 7100 133120 7120
rect 133380 7100 133620 7120
rect 133880 7100 134120 7120
rect 134380 7100 134620 7120
rect 134880 7100 135120 7120
rect 135380 7100 135620 7120
rect 135880 7100 136120 7120
rect 136380 7100 136620 7120
rect 136880 7100 137120 7120
rect 137380 7100 137620 7120
rect 137880 7100 138120 7120
rect 138380 7100 138620 7120
rect 138880 7100 139120 7120
rect 139380 7100 139620 7120
rect 139880 7100 140000 7120
rect 104000 7090 140000 7100
rect 104000 7020 128150 7090
rect 128350 7020 128650 7090
rect 128850 7020 129150 7090
rect 129350 7020 129650 7090
rect 129850 7020 130150 7090
rect 130350 7020 130650 7090
rect 130850 7020 131150 7090
rect 131350 7020 131650 7090
rect 131850 7020 132150 7090
rect 132350 7020 132650 7090
rect 132850 7020 133150 7090
rect 133350 7020 133650 7090
rect 133850 7020 134150 7090
rect 134350 7020 134650 7090
rect 134850 7020 135150 7090
rect 135350 7020 135650 7090
rect 135850 7020 136150 7090
rect 136350 7020 136650 7090
rect 136850 7020 137150 7090
rect 137350 7020 137650 7090
rect 137850 7020 138150 7090
rect 138350 7020 138650 7090
rect 138850 7020 139150 7090
rect 139350 7020 139650 7090
rect 139850 7020 140000 7090
rect 104000 6980 140000 7020
rect 104000 6910 128150 6980
rect 128350 6910 128650 6980
rect 128850 6910 129150 6980
rect 129350 6910 129650 6980
rect 129850 6910 130150 6980
rect 130350 6910 130650 6980
rect 130850 6910 131150 6980
rect 131350 6910 131650 6980
rect 131850 6910 132150 6980
rect 132350 6910 132650 6980
rect 132850 6910 133150 6980
rect 133350 6910 133650 6980
rect 133850 6910 134150 6980
rect 134350 6910 134650 6980
rect 134850 6910 135150 6980
rect 135350 6910 135650 6980
rect 135850 6910 136150 6980
rect 136350 6910 136650 6980
rect 136850 6910 137150 6980
rect 137350 6910 137650 6980
rect 137850 6910 138150 6980
rect 138350 6910 138650 6980
rect 138850 6910 139150 6980
rect 139350 6910 139650 6980
rect 139850 6910 140000 6980
rect 104000 6900 140000 6910
rect 104000 6880 104120 6900
rect 104380 6880 104620 6900
rect 104880 6880 105120 6900
rect 105380 6880 105620 6900
rect 105880 6880 106120 6900
rect 106380 6880 106620 6900
rect 106880 6880 107120 6900
rect 107380 6880 107620 6900
rect 107880 6880 108120 6900
rect 108380 6880 108620 6900
rect 108880 6880 109120 6900
rect 109380 6880 109620 6900
rect 109880 6880 110120 6900
rect 110380 6880 110620 6900
rect 110880 6880 111120 6900
rect 111380 6880 111620 6900
rect 111880 6880 112120 6900
rect 112380 6880 112620 6900
rect 112880 6880 113120 6900
rect 113380 6880 113620 6900
rect 113880 6880 114120 6900
rect 114380 6880 114620 6900
rect 114880 6880 115120 6900
rect 115380 6880 115620 6900
rect 115880 6880 116120 6900
rect 116380 6880 116620 6900
rect 116880 6880 117120 6900
rect 117380 6880 117620 6900
rect 117880 6880 118120 6900
rect 118380 6880 118620 6900
rect 118880 6880 119120 6900
rect 119380 6880 119620 6900
rect 119880 6880 120120 6900
rect 120380 6880 120620 6900
rect 120880 6880 121120 6900
rect 121380 6880 121620 6900
rect 121880 6880 122120 6900
rect 122380 6880 122620 6900
rect 122880 6880 123120 6900
rect 123380 6880 123620 6900
rect 123880 6880 124120 6900
rect 124380 6880 124620 6900
rect 124880 6880 125120 6900
rect 125380 6880 125620 6900
rect 125880 6880 126120 6900
rect 126380 6880 126620 6900
rect 126880 6880 127120 6900
rect 127380 6880 127620 6900
rect 127880 6880 128120 6900
rect 128380 6880 128620 6900
rect 128880 6880 129120 6900
rect 129380 6880 129620 6900
rect 129880 6880 130120 6900
rect 130380 6880 130620 6900
rect 130880 6880 131120 6900
rect 131380 6880 131620 6900
rect 131880 6880 132120 6900
rect 132380 6880 132620 6900
rect 132880 6880 133120 6900
rect 133380 6880 133620 6900
rect 133880 6880 134120 6900
rect 134380 6880 134620 6900
rect 134880 6880 135120 6900
rect 135380 6880 135620 6900
rect 135880 6880 136120 6900
rect 136380 6880 136620 6900
rect 136880 6880 137120 6900
rect 137380 6880 137620 6900
rect 137880 6880 138120 6900
rect 138380 6880 138620 6900
rect 138880 6880 139120 6900
rect 139380 6880 139620 6900
rect 139880 6880 140000 6900
rect 104000 6620 104100 6880
rect 104400 6620 104600 6880
rect 104900 6620 105100 6880
rect 105400 6620 105600 6880
rect 105900 6620 106100 6880
rect 106400 6620 106600 6880
rect 106900 6620 107100 6880
rect 107400 6620 107600 6880
rect 107900 6620 108100 6880
rect 108400 6620 108600 6880
rect 108900 6620 109100 6880
rect 109400 6620 109600 6880
rect 109900 6620 110100 6880
rect 110400 6620 110600 6880
rect 110900 6620 111100 6880
rect 111400 6620 111600 6880
rect 111900 6620 112100 6880
rect 112400 6620 112600 6880
rect 112900 6620 113100 6880
rect 113400 6620 113600 6880
rect 113900 6620 114100 6880
rect 114400 6620 114600 6880
rect 114900 6620 115100 6880
rect 115400 6620 115600 6880
rect 115900 6620 116100 6880
rect 116400 6620 116600 6880
rect 116900 6620 117100 6880
rect 117400 6620 117600 6880
rect 117900 6620 118100 6880
rect 118400 6620 118600 6880
rect 118900 6620 119100 6880
rect 119400 6620 119600 6880
rect 119900 6620 120100 6880
rect 120400 6620 120600 6880
rect 120900 6620 121100 6880
rect 121400 6620 121600 6880
rect 121900 6620 122100 6880
rect 122400 6620 122600 6880
rect 122900 6620 123100 6880
rect 123400 6620 123600 6880
rect 123900 6620 124100 6880
rect 124400 6620 124600 6880
rect 124900 6620 125100 6880
rect 125400 6620 125600 6880
rect 125900 6620 126100 6880
rect 126400 6620 126600 6880
rect 126900 6620 127100 6880
rect 127400 6620 127600 6880
rect 127900 6850 128100 6880
rect 127900 6650 128020 6850
rect 128090 6650 128100 6850
rect 127900 6620 128100 6650
rect 128400 6850 128600 6880
rect 128400 6650 128410 6850
rect 128480 6650 128520 6850
rect 128590 6650 128600 6850
rect 128400 6620 128600 6650
rect 128900 6850 129100 6880
rect 128900 6650 128910 6850
rect 128980 6650 129020 6850
rect 129090 6650 129100 6850
rect 128900 6620 129100 6650
rect 129400 6850 129600 6880
rect 129400 6650 129410 6850
rect 129480 6650 129520 6850
rect 129590 6650 129600 6850
rect 129400 6620 129600 6650
rect 129900 6850 130100 6880
rect 129900 6650 129910 6850
rect 129980 6650 130020 6850
rect 130090 6650 130100 6850
rect 129900 6620 130100 6650
rect 130400 6850 130600 6880
rect 130400 6650 130410 6850
rect 130480 6650 130520 6850
rect 130590 6650 130600 6850
rect 130400 6620 130600 6650
rect 130900 6850 131100 6880
rect 130900 6650 130910 6850
rect 130980 6650 131020 6850
rect 131090 6650 131100 6850
rect 130900 6620 131100 6650
rect 131400 6850 131600 6880
rect 131400 6650 131410 6850
rect 131480 6650 131520 6850
rect 131590 6650 131600 6850
rect 131400 6620 131600 6650
rect 131900 6850 132100 6880
rect 131900 6650 131910 6850
rect 131980 6650 132020 6850
rect 132090 6650 132100 6850
rect 131900 6620 132100 6650
rect 132400 6850 132600 6880
rect 132400 6650 132410 6850
rect 132480 6650 132520 6850
rect 132590 6650 132600 6850
rect 132400 6620 132600 6650
rect 132900 6850 133100 6880
rect 132900 6650 132910 6850
rect 132980 6650 133020 6850
rect 133090 6650 133100 6850
rect 132900 6620 133100 6650
rect 133400 6850 133600 6880
rect 133400 6650 133410 6850
rect 133480 6650 133520 6850
rect 133590 6650 133600 6850
rect 133400 6620 133600 6650
rect 133900 6850 134100 6880
rect 133900 6650 133910 6850
rect 133980 6650 134020 6850
rect 134090 6650 134100 6850
rect 133900 6620 134100 6650
rect 134400 6850 134600 6880
rect 134400 6650 134410 6850
rect 134480 6650 134520 6850
rect 134590 6650 134600 6850
rect 134400 6620 134600 6650
rect 134900 6850 135100 6880
rect 134900 6650 134910 6850
rect 134980 6650 135020 6850
rect 135090 6650 135100 6850
rect 134900 6620 135100 6650
rect 135400 6850 135600 6880
rect 135400 6650 135410 6850
rect 135480 6650 135520 6850
rect 135590 6650 135600 6850
rect 135400 6620 135600 6650
rect 135900 6850 136100 6880
rect 135900 6650 135910 6850
rect 135980 6650 136020 6850
rect 136090 6650 136100 6850
rect 135900 6620 136100 6650
rect 136400 6850 136600 6880
rect 136400 6650 136410 6850
rect 136480 6650 136520 6850
rect 136590 6650 136600 6850
rect 136400 6620 136600 6650
rect 136900 6850 137100 6880
rect 136900 6650 136910 6850
rect 136980 6650 137020 6850
rect 137090 6650 137100 6850
rect 136900 6620 137100 6650
rect 137400 6850 137600 6880
rect 137400 6650 137410 6850
rect 137480 6650 137520 6850
rect 137590 6650 137600 6850
rect 137400 6620 137600 6650
rect 137900 6850 138100 6880
rect 137900 6650 137910 6850
rect 137980 6650 138020 6850
rect 138090 6650 138100 6850
rect 137900 6620 138100 6650
rect 138400 6850 138600 6880
rect 138400 6650 138410 6850
rect 138480 6650 138520 6850
rect 138590 6650 138600 6850
rect 138400 6620 138600 6650
rect 138900 6850 139100 6880
rect 138900 6650 138910 6850
rect 138980 6650 139020 6850
rect 139090 6650 139100 6850
rect 138900 6620 139100 6650
rect 139400 6850 139600 6880
rect 139400 6650 139410 6850
rect 139480 6650 139520 6850
rect 139590 6650 139600 6850
rect 139400 6620 139600 6650
rect 139900 6850 140000 6880
rect 139900 6650 139910 6850
rect 139980 6650 140000 6850
rect 139900 6620 140000 6650
rect 104000 6600 104120 6620
rect 104380 6600 104620 6620
rect 104880 6600 105120 6620
rect 105380 6600 105620 6620
rect 105880 6600 106120 6620
rect 106380 6600 106620 6620
rect 106880 6600 107120 6620
rect 107380 6600 107620 6620
rect 107880 6600 108120 6620
rect 108380 6600 108620 6620
rect 108880 6600 109120 6620
rect 109380 6600 109620 6620
rect 109880 6600 110120 6620
rect 110380 6600 110620 6620
rect 110880 6600 111120 6620
rect 111380 6600 111620 6620
rect 111880 6600 112120 6620
rect 112380 6600 112620 6620
rect 112880 6600 113120 6620
rect 113380 6600 113620 6620
rect 113880 6600 114120 6620
rect 114380 6600 114620 6620
rect 114880 6600 115120 6620
rect 115380 6600 115620 6620
rect 115880 6600 116120 6620
rect 116380 6600 116620 6620
rect 116880 6600 117120 6620
rect 117380 6600 117620 6620
rect 117880 6600 118120 6620
rect 118380 6600 118620 6620
rect 118880 6600 119120 6620
rect 119380 6600 119620 6620
rect 119880 6600 120120 6620
rect 120380 6600 120620 6620
rect 120880 6600 121120 6620
rect 121380 6600 121620 6620
rect 121880 6600 122120 6620
rect 122380 6600 122620 6620
rect 122880 6600 123120 6620
rect 123380 6600 123620 6620
rect 123880 6600 124120 6620
rect 124380 6600 124620 6620
rect 124880 6600 125120 6620
rect 125380 6600 125620 6620
rect 125880 6600 126120 6620
rect 126380 6600 126620 6620
rect 126880 6600 127120 6620
rect 127380 6600 127620 6620
rect 127880 6600 128120 6620
rect 128380 6600 128620 6620
rect 128880 6600 129120 6620
rect 129380 6600 129620 6620
rect 129880 6600 130120 6620
rect 130380 6600 130620 6620
rect 130880 6600 131120 6620
rect 131380 6600 131620 6620
rect 131880 6600 132120 6620
rect 132380 6600 132620 6620
rect 132880 6600 133120 6620
rect 133380 6600 133620 6620
rect 133880 6600 134120 6620
rect 134380 6600 134620 6620
rect 134880 6600 135120 6620
rect 135380 6600 135620 6620
rect 135880 6600 136120 6620
rect 136380 6600 136620 6620
rect 136880 6600 137120 6620
rect 137380 6600 137620 6620
rect 137880 6600 138120 6620
rect 138380 6600 138620 6620
rect 138880 6600 139120 6620
rect 139380 6600 139620 6620
rect 139880 6600 140000 6620
rect 104000 6590 140000 6600
rect 104000 6520 128150 6590
rect 128350 6520 128650 6590
rect 128850 6520 129150 6590
rect 129350 6520 129650 6590
rect 129850 6520 130150 6590
rect 130350 6520 130650 6590
rect 130850 6520 131150 6590
rect 131350 6520 131650 6590
rect 131850 6520 132150 6590
rect 132350 6520 132650 6590
rect 132850 6520 133150 6590
rect 133350 6520 133650 6590
rect 133850 6520 134150 6590
rect 134350 6520 134650 6590
rect 134850 6520 135150 6590
rect 135350 6520 135650 6590
rect 135850 6520 136150 6590
rect 136350 6520 136650 6590
rect 136850 6520 137150 6590
rect 137350 6520 137650 6590
rect 137850 6520 138150 6590
rect 138350 6520 138650 6590
rect 138850 6520 139150 6590
rect 139350 6520 139650 6590
rect 139850 6520 140000 6590
rect 104000 6480 140000 6520
rect 104000 6410 128150 6480
rect 128350 6410 128650 6480
rect 128850 6410 129150 6480
rect 129350 6410 129650 6480
rect 129850 6410 130150 6480
rect 130350 6410 130650 6480
rect 130850 6410 131150 6480
rect 131350 6410 131650 6480
rect 131850 6410 132150 6480
rect 132350 6410 132650 6480
rect 132850 6410 133150 6480
rect 133350 6410 133650 6480
rect 133850 6410 134150 6480
rect 134350 6410 134650 6480
rect 134850 6410 135150 6480
rect 135350 6410 135650 6480
rect 135850 6410 136150 6480
rect 136350 6410 136650 6480
rect 136850 6410 137150 6480
rect 137350 6410 137650 6480
rect 137850 6410 138150 6480
rect 138350 6410 138650 6480
rect 138850 6410 139150 6480
rect 139350 6410 139650 6480
rect 139850 6410 140000 6480
rect 104000 6400 140000 6410
rect 104000 6380 104120 6400
rect 104380 6380 104620 6400
rect 104880 6380 105120 6400
rect 105380 6380 105620 6400
rect 105880 6380 106120 6400
rect 106380 6380 106620 6400
rect 106880 6380 107120 6400
rect 107380 6380 107620 6400
rect 107880 6380 108120 6400
rect 108380 6380 108620 6400
rect 108880 6380 109120 6400
rect 109380 6380 109620 6400
rect 109880 6380 110120 6400
rect 110380 6380 110620 6400
rect 110880 6380 111120 6400
rect 111380 6380 111620 6400
rect 111880 6380 112120 6400
rect 112380 6380 112620 6400
rect 112880 6380 113120 6400
rect 113380 6380 113620 6400
rect 113880 6380 114120 6400
rect 114380 6380 114620 6400
rect 114880 6380 115120 6400
rect 115380 6380 115620 6400
rect 115880 6380 116120 6400
rect 116380 6380 116620 6400
rect 116880 6380 117120 6400
rect 117380 6380 117620 6400
rect 117880 6380 118120 6400
rect 118380 6380 118620 6400
rect 118880 6380 119120 6400
rect 119380 6380 119620 6400
rect 119880 6380 120120 6400
rect 120380 6380 120620 6400
rect 120880 6380 121120 6400
rect 121380 6380 121620 6400
rect 121880 6380 122120 6400
rect 122380 6380 122620 6400
rect 122880 6380 123120 6400
rect 123380 6380 123620 6400
rect 123880 6380 124120 6400
rect 124380 6380 124620 6400
rect 124880 6380 125120 6400
rect 125380 6380 125620 6400
rect 125880 6380 126120 6400
rect 126380 6380 126620 6400
rect 126880 6380 127120 6400
rect 127380 6380 127620 6400
rect 127880 6380 128120 6400
rect 128380 6380 128620 6400
rect 128880 6380 129120 6400
rect 129380 6380 129620 6400
rect 129880 6380 130120 6400
rect 130380 6380 130620 6400
rect 130880 6380 131120 6400
rect 131380 6380 131620 6400
rect 131880 6380 132120 6400
rect 132380 6380 132620 6400
rect 132880 6380 133120 6400
rect 133380 6380 133620 6400
rect 133880 6380 134120 6400
rect 134380 6380 134620 6400
rect 134880 6380 135120 6400
rect 135380 6380 135620 6400
rect 135880 6380 136120 6400
rect 136380 6380 136620 6400
rect 136880 6380 137120 6400
rect 137380 6380 137620 6400
rect 137880 6380 138120 6400
rect 138380 6380 138620 6400
rect 138880 6380 139120 6400
rect 139380 6380 139620 6400
rect 139880 6380 140000 6400
rect 104000 6120 104100 6380
rect 104400 6120 104600 6380
rect 104900 6120 105100 6380
rect 105400 6120 105600 6380
rect 105900 6120 106100 6380
rect 106400 6120 106600 6380
rect 106900 6120 107100 6380
rect 107400 6120 107600 6380
rect 107900 6120 108100 6380
rect 108400 6120 108600 6380
rect 108900 6120 109100 6380
rect 109400 6120 109600 6380
rect 109900 6120 110100 6380
rect 110400 6120 110600 6380
rect 110900 6120 111100 6380
rect 111400 6120 111600 6380
rect 111900 6120 112100 6380
rect 112400 6120 112600 6380
rect 112900 6120 113100 6380
rect 113400 6120 113600 6380
rect 113900 6120 114100 6380
rect 114400 6120 114600 6380
rect 114900 6120 115100 6380
rect 115400 6120 115600 6380
rect 115900 6120 116100 6380
rect 116400 6120 116600 6380
rect 116900 6120 117100 6380
rect 117400 6120 117600 6380
rect 117900 6120 118100 6380
rect 118400 6120 118600 6380
rect 118900 6120 119100 6380
rect 119400 6120 119600 6380
rect 119900 6120 120100 6380
rect 120400 6120 120600 6380
rect 120900 6120 121100 6380
rect 121400 6120 121600 6380
rect 121900 6120 122100 6380
rect 122400 6120 122600 6380
rect 122900 6120 123100 6380
rect 123400 6120 123600 6380
rect 123900 6120 124100 6380
rect 124400 6120 124600 6380
rect 124900 6120 125100 6380
rect 125400 6120 125600 6380
rect 125900 6120 126100 6380
rect 126400 6120 126600 6380
rect 126900 6120 127100 6380
rect 127400 6120 127600 6380
rect 127900 6350 128100 6380
rect 127900 6150 128020 6350
rect 128090 6150 128100 6350
rect 127900 6120 128100 6150
rect 128400 6350 128600 6380
rect 128400 6150 128410 6350
rect 128480 6150 128520 6350
rect 128590 6150 128600 6350
rect 128400 6120 128600 6150
rect 128900 6350 129100 6380
rect 128900 6150 128910 6350
rect 128980 6150 129020 6350
rect 129090 6150 129100 6350
rect 128900 6120 129100 6150
rect 129400 6350 129600 6380
rect 129400 6150 129410 6350
rect 129480 6150 129520 6350
rect 129590 6150 129600 6350
rect 129400 6120 129600 6150
rect 129900 6350 130100 6380
rect 129900 6150 129910 6350
rect 129980 6150 130020 6350
rect 130090 6150 130100 6350
rect 129900 6120 130100 6150
rect 130400 6350 130600 6380
rect 130400 6150 130410 6350
rect 130480 6150 130520 6350
rect 130590 6150 130600 6350
rect 130400 6120 130600 6150
rect 130900 6350 131100 6380
rect 130900 6150 130910 6350
rect 130980 6150 131020 6350
rect 131090 6150 131100 6350
rect 130900 6120 131100 6150
rect 131400 6350 131600 6380
rect 131400 6150 131410 6350
rect 131480 6150 131520 6350
rect 131590 6150 131600 6350
rect 131400 6120 131600 6150
rect 131900 6350 132100 6380
rect 131900 6150 131910 6350
rect 131980 6150 132020 6350
rect 132090 6150 132100 6350
rect 131900 6120 132100 6150
rect 132400 6350 132600 6380
rect 132400 6150 132410 6350
rect 132480 6150 132520 6350
rect 132590 6150 132600 6350
rect 132400 6120 132600 6150
rect 132900 6350 133100 6380
rect 132900 6150 132910 6350
rect 132980 6150 133020 6350
rect 133090 6150 133100 6350
rect 132900 6120 133100 6150
rect 133400 6350 133600 6380
rect 133400 6150 133410 6350
rect 133480 6150 133520 6350
rect 133590 6150 133600 6350
rect 133400 6120 133600 6150
rect 133900 6350 134100 6380
rect 133900 6150 133910 6350
rect 133980 6150 134020 6350
rect 134090 6150 134100 6350
rect 133900 6120 134100 6150
rect 134400 6350 134600 6380
rect 134400 6150 134410 6350
rect 134480 6150 134520 6350
rect 134590 6150 134600 6350
rect 134400 6120 134600 6150
rect 134900 6350 135100 6380
rect 134900 6150 134910 6350
rect 134980 6150 135020 6350
rect 135090 6150 135100 6350
rect 134900 6120 135100 6150
rect 135400 6350 135600 6380
rect 135400 6150 135410 6350
rect 135480 6150 135520 6350
rect 135590 6150 135600 6350
rect 135400 6120 135600 6150
rect 135900 6350 136100 6380
rect 135900 6150 135910 6350
rect 135980 6150 136020 6350
rect 136090 6150 136100 6350
rect 135900 6120 136100 6150
rect 136400 6350 136600 6380
rect 136400 6150 136410 6350
rect 136480 6150 136520 6350
rect 136590 6150 136600 6350
rect 136400 6120 136600 6150
rect 136900 6350 137100 6380
rect 136900 6150 136910 6350
rect 136980 6150 137020 6350
rect 137090 6150 137100 6350
rect 136900 6120 137100 6150
rect 137400 6350 137600 6380
rect 137400 6150 137410 6350
rect 137480 6150 137520 6350
rect 137590 6150 137600 6350
rect 137400 6120 137600 6150
rect 137900 6350 138100 6380
rect 137900 6150 137910 6350
rect 137980 6150 138020 6350
rect 138090 6150 138100 6350
rect 137900 6120 138100 6150
rect 138400 6350 138600 6380
rect 138400 6150 138410 6350
rect 138480 6150 138520 6350
rect 138590 6150 138600 6350
rect 138400 6120 138600 6150
rect 138900 6350 139100 6380
rect 138900 6150 138910 6350
rect 138980 6150 139020 6350
rect 139090 6150 139100 6350
rect 138900 6120 139100 6150
rect 139400 6350 139600 6380
rect 139400 6150 139410 6350
rect 139480 6150 139520 6350
rect 139590 6150 139600 6350
rect 139400 6120 139600 6150
rect 139900 6350 140000 6380
rect 139900 6150 139910 6350
rect 139980 6150 140000 6350
rect 139900 6120 140000 6150
rect 104000 6100 104120 6120
rect 104380 6100 104620 6120
rect 104880 6100 105120 6120
rect 105380 6100 105620 6120
rect 105880 6100 106120 6120
rect 106380 6100 106620 6120
rect 106880 6100 107120 6120
rect 107380 6100 107620 6120
rect 107880 6100 108120 6120
rect 108380 6100 108620 6120
rect 108880 6100 109120 6120
rect 109380 6100 109620 6120
rect 109880 6100 110120 6120
rect 110380 6100 110620 6120
rect 110880 6100 111120 6120
rect 111380 6100 111620 6120
rect 111880 6100 112120 6120
rect 112380 6100 112620 6120
rect 112880 6100 113120 6120
rect 113380 6100 113620 6120
rect 113880 6100 114120 6120
rect 114380 6100 114620 6120
rect 114880 6100 115120 6120
rect 115380 6100 115620 6120
rect 115880 6100 116120 6120
rect 116380 6100 116620 6120
rect 116880 6100 117120 6120
rect 117380 6100 117620 6120
rect 117880 6100 118120 6120
rect 118380 6100 118620 6120
rect 118880 6100 119120 6120
rect 119380 6100 119620 6120
rect 119880 6100 120120 6120
rect 120380 6100 120620 6120
rect 120880 6100 121120 6120
rect 121380 6100 121620 6120
rect 121880 6100 122120 6120
rect 122380 6100 122620 6120
rect 122880 6100 123120 6120
rect 123380 6100 123620 6120
rect 123880 6100 124120 6120
rect 124380 6100 124620 6120
rect 124880 6100 125120 6120
rect 125380 6100 125620 6120
rect 125880 6100 126120 6120
rect 126380 6100 126620 6120
rect 126880 6100 127120 6120
rect 127380 6100 127620 6120
rect 127880 6100 128120 6120
rect 128380 6100 128620 6120
rect 128880 6100 129120 6120
rect 129380 6100 129620 6120
rect 129880 6100 130120 6120
rect 130380 6100 130620 6120
rect 130880 6100 131120 6120
rect 131380 6100 131620 6120
rect 131880 6100 132120 6120
rect 132380 6100 132620 6120
rect 132880 6100 133120 6120
rect 133380 6100 133620 6120
rect 133880 6100 134120 6120
rect 134380 6100 134620 6120
rect 134880 6100 135120 6120
rect 135380 6100 135620 6120
rect 135880 6100 136120 6120
rect 136380 6100 136620 6120
rect 136880 6100 137120 6120
rect 137380 6100 137620 6120
rect 137880 6100 138120 6120
rect 138380 6100 138620 6120
rect 138880 6100 139120 6120
rect 139380 6100 139620 6120
rect 139880 6100 140000 6120
rect 104000 6090 140000 6100
rect 104000 6020 128150 6090
rect 128350 6020 128650 6090
rect 128850 6020 129150 6090
rect 129350 6020 129650 6090
rect 129850 6020 130150 6090
rect 130350 6020 130650 6090
rect 130850 6020 131150 6090
rect 131350 6020 131650 6090
rect 131850 6020 132150 6090
rect 132350 6020 132650 6090
rect 132850 6020 133150 6090
rect 133350 6020 133650 6090
rect 133850 6020 134150 6090
rect 134350 6020 134650 6090
rect 134850 6020 135150 6090
rect 135350 6020 135650 6090
rect 135850 6020 136150 6090
rect 136350 6020 136650 6090
rect 136850 6020 137150 6090
rect 137350 6020 137650 6090
rect 137850 6020 138150 6090
rect 138350 6020 138650 6090
rect 138850 6020 139150 6090
rect 139350 6020 139650 6090
rect 139850 6020 140000 6090
rect 104000 6000 140000 6020
rect 104000 5900 128000 6000
rect 104000 5880 104120 5900
rect 104380 5880 104620 5900
rect 104880 5880 105120 5900
rect 105380 5880 105620 5900
rect 105880 5880 106120 5900
rect 106380 5880 106620 5900
rect 106880 5880 107120 5900
rect 107380 5880 107620 5900
rect 107880 5880 108120 5900
rect 108380 5880 108620 5900
rect 108880 5880 109120 5900
rect 109380 5880 109620 5900
rect 109880 5880 110120 5900
rect 110380 5880 110620 5900
rect 110880 5880 111120 5900
rect 111380 5880 111620 5900
rect 111880 5880 112120 5900
rect 112380 5880 112620 5900
rect 112880 5880 113120 5900
rect 113380 5880 113620 5900
rect 113880 5880 114120 5900
rect 114380 5880 114620 5900
rect 114880 5880 115120 5900
rect 115380 5880 115620 5900
rect 115880 5880 116120 5900
rect 116380 5880 116620 5900
rect 116880 5880 117120 5900
rect 117380 5880 117620 5900
rect 117880 5880 118120 5900
rect 118380 5880 118620 5900
rect 118880 5880 119120 5900
rect 119380 5880 119620 5900
rect 119880 5880 120120 5900
rect 120380 5880 120620 5900
rect 120880 5880 121120 5900
rect 121380 5880 121620 5900
rect 121880 5880 122120 5900
rect 122380 5880 122620 5900
rect 122880 5880 123120 5900
rect 123380 5880 123620 5900
rect 123880 5880 124120 5900
rect 124380 5880 124620 5900
rect 124880 5880 125120 5900
rect 125380 5880 125620 5900
rect 125880 5880 126120 5900
rect 126380 5880 126620 5900
rect 126880 5880 127120 5900
rect 127380 5880 127620 5900
rect 127880 5880 128000 5900
rect 104000 5620 104100 5880
rect 104400 5620 104600 5880
rect 104900 5620 105100 5880
rect 105400 5620 105600 5880
rect 105900 5620 106100 5880
rect 106400 5620 106600 5880
rect 106900 5620 107100 5880
rect 107400 5620 107600 5880
rect 107900 5620 108100 5880
rect 108400 5620 108600 5880
rect 108900 5620 109100 5880
rect 109400 5620 109600 5880
rect 109900 5620 110100 5880
rect 110400 5620 110600 5880
rect 110900 5620 111100 5880
rect 111400 5620 111600 5880
rect 111900 5620 112100 5880
rect 112400 5620 112600 5880
rect 112900 5620 113100 5880
rect 113400 5620 113600 5880
rect 113900 5620 114100 5880
rect 114400 5620 114600 5880
rect 114900 5620 115100 5880
rect 115400 5620 115600 5880
rect 115900 5620 116100 5880
rect 116400 5620 116600 5880
rect 116900 5620 117100 5880
rect 117400 5620 117600 5880
rect 117900 5620 118100 5880
rect 118400 5620 118600 5880
rect 118900 5620 119100 5880
rect 119400 5620 119600 5880
rect 119900 5620 120100 5880
rect 120400 5620 120600 5880
rect 120900 5620 121100 5880
rect 121400 5620 121600 5880
rect 121900 5620 122100 5880
rect 122400 5620 122600 5880
rect 122900 5620 123100 5880
rect 123400 5620 123600 5880
rect 123900 5620 124100 5880
rect 124400 5620 124600 5880
rect 124900 5620 125100 5880
rect 125400 5620 125600 5880
rect 125900 5620 126100 5880
rect 126400 5620 126600 5880
rect 126900 5620 127100 5880
rect 127400 5620 127600 5880
rect 127900 5620 128000 5880
rect 104000 5600 104120 5620
rect 104380 5600 104620 5620
rect 104880 5600 105120 5620
rect 105380 5600 105620 5620
rect 105880 5600 106120 5620
rect 106380 5600 106620 5620
rect 106880 5600 107120 5620
rect 107380 5600 107620 5620
rect 107880 5600 108120 5620
rect 108380 5600 108620 5620
rect 108880 5600 109120 5620
rect 109380 5600 109620 5620
rect 109880 5600 110120 5620
rect 110380 5600 110620 5620
rect 110880 5600 111120 5620
rect 111380 5600 111620 5620
rect 111880 5600 112120 5620
rect 112380 5600 112620 5620
rect 112880 5600 113120 5620
rect 113380 5600 113620 5620
rect 113880 5600 114120 5620
rect 114380 5600 114620 5620
rect 114880 5600 115120 5620
rect 115380 5600 115620 5620
rect 115880 5600 116120 5620
rect 116380 5600 116620 5620
rect 116880 5600 117120 5620
rect 117380 5600 117620 5620
rect 117880 5600 118120 5620
rect 118380 5600 118620 5620
rect 118880 5600 119120 5620
rect 119380 5600 119620 5620
rect 119880 5600 120120 5620
rect 120380 5600 120620 5620
rect 120880 5600 121120 5620
rect 121380 5600 121620 5620
rect 121880 5600 122120 5620
rect 122380 5600 122620 5620
rect 122880 5600 123120 5620
rect 123380 5600 123620 5620
rect 123880 5600 124120 5620
rect 124380 5600 124620 5620
rect 124880 5600 125120 5620
rect 125380 5600 125620 5620
rect 125880 5600 126120 5620
rect 126380 5600 126620 5620
rect 126880 5600 127120 5620
rect 127380 5600 127620 5620
rect 127880 5600 128000 5620
rect 104000 5400 128000 5600
rect 104000 5380 104120 5400
rect 104380 5380 104620 5400
rect 104880 5380 105120 5400
rect 105380 5380 105620 5400
rect 105880 5380 106120 5400
rect 106380 5380 106620 5400
rect 106880 5380 107120 5400
rect 107380 5380 107620 5400
rect 107880 5380 108120 5400
rect 108380 5380 108620 5400
rect 108880 5380 109120 5400
rect 109380 5380 109620 5400
rect 109880 5380 110120 5400
rect 110380 5380 110620 5400
rect 110880 5380 111120 5400
rect 111380 5380 111620 5400
rect 111880 5380 112120 5400
rect 112380 5380 112620 5400
rect 112880 5380 113120 5400
rect 113380 5380 113620 5400
rect 113880 5380 114120 5400
rect 114380 5380 114620 5400
rect 114880 5380 115120 5400
rect 115380 5380 115620 5400
rect 115880 5380 116120 5400
rect 116380 5380 116620 5400
rect 116880 5380 117120 5400
rect 117380 5380 117620 5400
rect 117880 5380 118120 5400
rect 118380 5380 118620 5400
rect 118880 5380 119120 5400
rect 119380 5380 119620 5400
rect 119880 5380 120120 5400
rect 120380 5380 120620 5400
rect 120880 5380 121120 5400
rect 121380 5380 121620 5400
rect 121880 5380 122120 5400
rect 122380 5380 122620 5400
rect 122880 5380 123120 5400
rect 123380 5380 123620 5400
rect 123880 5380 124120 5400
rect 124380 5380 124620 5400
rect 124880 5380 125120 5400
rect 125380 5380 125620 5400
rect 125880 5380 126120 5400
rect 126380 5380 126620 5400
rect 126880 5380 127120 5400
rect 127380 5380 127620 5400
rect 127880 5380 128000 5400
rect 104000 5120 104100 5380
rect 104400 5120 104600 5380
rect 104900 5120 105100 5380
rect 105400 5120 105600 5380
rect 105900 5120 106100 5380
rect 106400 5120 106600 5380
rect 106900 5120 107100 5380
rect 107400 5120 107600 5380
rect 107900 5120 108100 5380
rect 108400 5120 108600 5380
rect 108900 5120 109100 5380
rect 109400 5120 109600 5380
rect 109900 5120 110100 5380
rect 110400 5120 110600 5380
rect 110900 5120 111100 5380
rect 111400 5120 111600 5380
rect 111900 5120 112100 5380
rect 112400 5120 112600 5380
rect 112900 5120 113100 5380
rect 113400 5120 113600 5380
rect 113900 5120 114100 5380
rect 114400 5120 114600 5380
rect 114900 5120 115100 5380
rect 115400 5120 115600 5380
rect 115900 5120 116100 5380
rect 116400 5120 116600 5380
rect 116900 5120 117100 5380
rect 117400 5120 117600 5380
rect 117900 5120 118100 5380
rect 118400 5120 118600 5380
rect 118900 5120 119100 5380
rect 119400 5120 119600 5380
rect 119900 5120 120100 5380
rect 120400 5120 120600 5380
rect 120900 5120 121100 5380
rect 121400 5120 121600 5380
rect 121900 5120 122100 5380
rect 122400 5120 122600 5380
rect 122900 5120 123100 5380
rect 123400 5120 123600 5380
rect 123900 5120 124100 5380
rect 124400 5120 124600 5380
rect 124900 5120 125100 5380
rect 125400 5120 125600 5380
rect 125900 5120 126100 5380
rect 126400 5120 126600 5380
rect 126900 5120 127100 5380
rect 127400 5120 127600 5380
rect 127900 5120 128000 5380
rect 104000 5100 104120 5120
rect 104380 5100 104620 5120
rect 104880 5100 105120 5120
rect 105380 5100 105620 5120
rect 105880 5100 106120 5120
rect 106380 5100 106620 5120
rect 106880 5100 107120 5120
rect 107380 5100 107620 5120
rect 107880 5100 108120 5120
rect 108380 5100 108620 5120
rect 108880 5100 109120 5120
rect 109380 5100 109620 5120
rect 109880 5100 110120 5120
rect 110380 5100 110620 5120
rect 110880 5100 111120 5120
rect 111380 5100 111620 5120
rect 111880 5100 112120 5120
rect 112380 5100 112620 5120
rect 112880 5100 113120 5120
rect 113380 5100 113620 5120
rect 113880 5100 114120 5120
rect 114380 5100 114620 5120
rect 114880 5100 115120 5120
rect 115380 5100 115620 5120
rect 115880 5100 116120 5120
rect 116380 5100 116620 5120
rect 116880 5100 117120 5120
rect 117380 5100 117620 5120
rect 117880 5100 118120 5120
rect 118380 5100 118620 5120
rect 118880 5100 119120 5120
rect 119380 5100 119620 5120
rect 119880 5100 120120 5120
rect 120380 5100 120620 5120
rect 120880 5100 121120 5120
rect 121380 5100 121620 5120
rect 121880 5100 122120 5120
rect 122380 5100 122620 5120
rect 122880 5100 123120 5120
rect 123380 5100 123620 5120
rect 123880 5100 124120 5120
rect 124380 5100 124620 5120
rect 124880 5100 125120 5120
rect 125380 5100 125620 5120
rect 125880 5100 126120 5120
rect 126380 5100 126620 5120
rect 126880 5100 127120 5120
rect 127380 5100 127620 5120
rect 127880 5100 128000 5120
rect 104000 4900 128000 5100
rect 104000 4880 104120 4900
rect 104380 4880 104620 4900
rect 104880 4880 105120 4900
rect 105380 4880 105620 4900
rect 105880 4880 106120 4900
rect 106380 4880 106620 4900
rect 106880 4880 107120 4900
rect 107380 4880 107620 4900
rect 107880 4880 108120 4900
rect 108380 4880 108620 4900
rect 108880 4880 109120 4900
rect 109380 4880 109620 4900
rect 109880 4880 110120 4900
rect 110380 4880 110620 4900
rect 110880 4880 111120 4900
rect 111380 4880 111620 4900
rect 111880 4880 112120 4900
rect 112380 4880 112620 4900
rect 112880 4880 113120 4900
rect 113380 4880 113620 4900
rect 113880 4880 114120 4900
rect 114380 4880 114620 4900
rect 114880 4880 115120 4900
rect 115380 4880 115620 4900
rect 115880 4880 116120 4900
rect 116380 4880 116620 4900
rect 116880 4880 117120 4900
rect 117380 4880 117620 4900
rect 117880 4880 118120 4900
rect 118380 4880 118620 4900
rect 118880 4880 119120 4900
rect 119380 4880 119620 4900
rect 119880 4880 120120 4900
rect 120380 4880 120620 4900
rect 120880 4880 121120 4900
rect 121380 4880 121620 4900
rect 121880 4880 122120 4900
rect 122380 4880 122620 4900
rect 122880 4880 123120 4900
rect 123380 4880 123620 4900
rect 123880 4880 124120 4900
rect 124380 4880 124620 4900
rect 124880 4880 125120 4900
rect 125380 4880 125620 4900
rect 125880 4880 126120 4900
rect 126380 4880 126620 4900
rect 126880 4880 127120 4900
rect 127380 4880 127620 4900
rect 127880 4880 128000 4900
rect 104000 4620 104100 4880
rect 104400 4620 104600 4880
rect 104900 4620 105100 4880
rect 105400 4620 105600 4880
rect 105900 4620 106100 4880
rect 106400 4620 106600 4880
rect 106900 4620 107100 4880
rect 107400 4620 107600 4880
rect 107900 4620 108100 4880
rect 108400 4620 108600 4880
rect 108900 4620 109100 4880
rect 109400 4620 109600 4880
rect 109900 4620 110100 4880
rect 110400 4620 110600 4880
rect 110900 4620 111100 4880
rect 111400 4620 111600 4880
rect 111900 4620 112100 4880
rect 112400 4620 112600 4880
rect 112900 4620 113100 4880
rect 113400 4620 113600 4880
rect 113900 4620 114100 4880
rect 114400 4620 114600 4880
rect 114900 4620 115100 4880
rect 115400 4620 115600 4880
rect 115900 4620 116100 4880
rect 116400 4620 116600 4880
rect 116900 4620 117100 4880
rect 117400 4620 117600 4880
rect 117900 4620 118100 4880
rect 118400 4620 118600 4880
rect 118900 4620 119100 4880
rect 119400 4620 119600 4880
rect 119900 4620 120100 4880
rect 120400 4620 120600 4880
rect 120900 4620 121100 4880
rect 121400 4620 121600 4880
rect 121900 4620 122100 4880
rect 122400 4620 122600 4880
rect 122900 4620 123100 4880
rect 123400 4620 123600 4880
rect 123900 4620 124100 4880
rect 124400 4620 124600 4880
rect 124900 4620 125100 4880
rect 125400 4620 125600 4880
rect 125900 4620 126100 4880
rect 126400 4620 126600 4880
rect 126900 4620 127100 4880
rect 127400 4620 127600 4880
rect 127900 4620 128000 4880
rect 104000 4600 104120 4620
rect 104380 4600 104620 4620
rect 104880 4600 105120 4620
rect 105380 4600 105620 4620
rect 105880 4600 106120 4620
rect 106380 4600 106620 4620
rect 106880 4600 107120 4620
rect 107380 4600 107620 4620
rect 107880 4600 108120 4620
rect 108380 4600 108620 4620
rect 108880 4600 109120 4620
rect 109380 4600 109620 4620
rect 109880 4600 110120 4620
rect 110380 4600 110620 4620
rect 110880 4600 111120 4620
rect 111380 4600 111620 4620
rect 111880 4600 112120 4620
rect 112380 4600 112620 4620
rect 112880 4600 113120 4620
rect 113380 4600 113620 4620
rect 113880 4600 114120 4620
rect 114380 4600 114620 4620
rect 114880 4600 115120 4620
rect 115380 4600 115620 4620
rect 115880 4600 116120 4620
rect 116380 4600 116620 4620
rect 116880 4600 117120 4620
rect 117380 4600 117620 4620
rect 117880 4600 118120 4620
rect 118380 4600 118620 4620
rect 118880 4600 119120 4620
rect 119380 4600 119620 4620
rect 119880 4600 120120 4620
rect 120380 4600 120620 4620
rect 120880 4600 121120 4620
rect 121380 4600 121620 4620
rect 121880 4600 122120 4620
rect 122380 4600 122620 4620
rect 122880 4600 123120 4620
rect 123380 4600 123620 4620
rect 123880 4600 124120 4620
rect 124380 4600 124620 4620
rect 124880 4600 125120 4620
rect 125380 4600 125620 4620
rect 125880 4600 126120 4620
rect 126380 4600 126620 4620
rect 126880 4600 127120 4620
rect 127380 4600 127620 4620
rect 127880 4600 128000 4620
rect 104000 4400 128000 4600
rect 104000 4380 104120 4400
rect 104380 4380 104620 4400
rect 104880 4380 105120 4400
rect 105380 4380 105620 4400
rect 105880 4380 106120 4400
rect 106380 4380 106620 4400
rect 106880 4380 107120 4400
rect 107380 4380 107620 4400
rect 107880 4380 108120 4400
rect 108380 4380 108620 4400
rect 108880 4380 109120 4400
rect 109380 4380 109620 4400
rect 109880 4380 110120 4400
rect 110380 4380 110620 4400
rect 110880 4380 111120 4400
rect 111380 4380 111620 4400
rect 111880 4380 112120 4400
rect 112380 4380 112620 4400
rect 112880 4380 113120 4400
rect 113380 4380 113620 4400
rect 113880 4380 114120 4400
rect 114380 4380 114620 4400
rect 114880 4380 115120 4400
rect 115380 4380 115620 4400
rect 115880 4380 116120 4400
rect 116380 4380 116620 4400
rect 116880 4380 117120 4400
rect 117380 4380 117620 4400
rect 117880 4380 118120 4400
rect 118380 4380 118620 4400
rect 118880 4380 119120 4400
rect 119380 4380 119620 4400
rect 119880 4380 120120 4400
rect 120380 4380 120620 4400
rect 120880 4380 121120 4400
rect 121380 4380 121620 4400
rect 121880 4380 122120 4400
rect 122380 4380 122620 4400
rect 122880 4380 123120 4400
rect 123380 4380 123620 4400
rect 123880 4380 124120 4400
rect 124380 4380 124620 4400
rect 124880 4380 125120 4400
rect 125380 4380 125620 4400
rect 125880 4380 126120 4400
rect 126380 4380 126620 4400
rect 126880 4380 127120 4400
rect 127380 4380 127620 4400
rect 127880 4380 128000 4400
rect 104000 4120 104100 4380
rect 104400 4120 104600 4380
rect 104900 4120 105100 4380
rect 105400 4120 105600 4380
rect 105900 4120 106100 4380
rect 106400 4120 106600 4380
rect 106900 4120 107100 4380
rect 107400 4120 107600 4380
rect 107900 4120 108100 4380
rect 108400 4120 108600 4380
rect 108900 4120 109100 4380
rect 109400 4120 109600 4380
rect 109900 4120 110100 4380
rect 110400 4120 110600 4380
rect 110900 4120 111100 4380
rect 111400 4120 111600 4380
rect 111900 4120 112100 4380
rect 112400 4120 112600 4380
rect 112900 4120 113100 4380
rect 113400 4120 113600 4380
rect 113900 4120 114100 4380
rect 114400 4120 114600 4380
rect 114900 4120 115100 4380
rect 115400 4120 115600 4380
rect 115900 4120 116100 4380
rect 116400 4120 116600 4380
rect 116900 4120 117100 4380
rect 117400 4120 117600 4380
rect 117900 4120 118100 4380
rect 118400 4120 118600 4380
rect 118900 4120 119100 4380
rect 119400 4120 119600 4380
rect 119900 4120 120100 4380
rect 120400 4120 120600 4380
rect 120900 4120 121100 4380
rect 121400 4120 121600 4380
rect 121900 4120 122100 4380
rect 122400 4120 122600 4380
rect 122900 4120 123100 4380
rect 123400 4120 123600 4380
rect 123900 4120 124100 4380
rect 124400 4120 124600 4380
rect 124900 4120 125100 4380
rect 125400 4120 125600 4380
rect 125900 4120 126100 4380
rect 126400 4120 126600 4380
rect 126900 4120 127100 4380
rect 127400 4120 127600 4380
rect 127900 4120 128000 4380
rect 104000 4100 104120 4120
rect 104380 4100 104620 4120
rect 104880 4100 105120 4120
rect 105380 4100 105620 4120
rect 105880 4100 106120 4120
rect 106380 4100 106620 4120
rect 106880 4100 107120 4120
rect 107380 4100 107620 4120
rect 107880 4100 108120 4120
rect 108380 4100 108620 4120
rect 108880 4100 109120 4120
rect 109380 4100 109620 4120
rect 109880 4100 110120 4120
rect 110380 4100 110620 4120
rect 110880 4100 111120 4120
rect 111380 4100 111620 4120
rect 111880 4100 112120 4120
rect 112380 4100 112620 4120
rect 112880 4100 113120 4120
rect 113380 4100 113620 4120
rect 113880 4100 114120 4120
rect 114380 4100 114620 4120
rect 114880 4100 115120 4120
rect 115380 4100 115620 4120
rect 115880 4100 116120 4120
rect 116380 4100 116620 4120
rect 116880 4100 117120 4120
rect 117380 4100 117620 4120
rect 117880 4100 118120 4120
rect 118380 4100 118620 4120
rect 118880 4100 119120 4120
rect 119380 4100 119620 4120
rect 119880 4100 120120 4120
rect 120380 4100 120620 4120
rect 120880 4100 121120 4120
rect 121380 4100 121620 4120
rect 121880 4100 122120 4120
rect 122380 4100 122620 4120
rect 122880 4100 123120 4120
rect 123380 4100 123620 4120
rect 123880 4100 124120 4120
rect 124380 4100 124620 4120
rect 124880 4100 125120 4120
rect 125380 4100 125620 4120
rect 125880 4100 126120 4120
rect 126380 4100 126620 4120
rect 126880 4100 127120 4120
rect 127380 4100 127620 4120
rect 127880 4100 128000 4120
rect 104000 3900 128000 4100
rect 104000 3880 104120 3900
rect 104380 3880 104620 3900
rect 104880 3880 105120 3900
rect 105380 3880 105620 3900
rect 105880 3880 106120 3900
rect 106380 3880 106620 3900
rect 106880 3880 107120 3900
rect 107380 3880 107620 3900
rect 107880 3880 108120 3900
rect 108380 3880 108620 3900
rect 108880 3880 109120 3900
rect 109380 3880 109620 3900
rect 109880 3880 110120 3900
rect 110380 3880 110620 3900
rect 110880 3880 111120 3900
rect 111380 3880 111620 3900
rect 111880 3880 112120 3900
rect 112380 3880 112620 3900
rect 112880 3880 113120 3900
rect 113380 3880 113620 3900
rect 113880 3880 114120 3900
rect 114380 3880 114620 3900
rect 114880 3880 115120 3900
rect 115380 3880 115620 3900
rect 115880 3880 116120 3900
rect 116380 3880 116620 3900
rect 116880 3880 117120 3900
rect 117380 3880 117620 3900
rect 117880 3880 118120 3900
rect 118380 3880 118620 3900
rect 118880 3880 119120 3900
rect 119380 3880 119620 3900
rect 119880 3880 120120 3900
rect 120380 3880 120620 3900
rect 120880 3880 121120 3900
rect 121380 3880 121620 3900
rect 121880 3880 122120 3900
rect 122380 3880 122620 3900
rect 122880 3880 123120 3900
rect 123380 3880 123620 3900
rect 123880 3880 124120 3900
rect 124380 3880 124620 3900
rect 124880 3880 125120 3900
rect 125380 3880 125620 3900
rect 125880 3880 126120 3900
rect 126380 3880 126620 3900
rect 126880 3880 127120 3900
rect 127380 3880 127620 3900
rect 127880 3880 128000 3900
rect 104000 3620 104100 3880
rect 104400 3620 104600 3880
rect 104900 3620 105100 3880
rect 105400 3620 105600 3880
rect 105900 3620 106100 3880
rect 106400 3620 106600 3880
rect 106900 3620 107100 3880
rect 107400 3620 107600 3880
rect 107900 3620 108100 3880
rect 108400 3620 108600 3880
rect 108900 3620 109100 3880
rect 109400 3620 109600 3880
rect 109900 3620 110100 3880
rect 110400 3620 110600 3880
rect 110900 3620 111100 3880
rect 111400 3620 111600 3880
rect 111900 3620 112100 3880
rect 112400 3620 112600 3880
rect 112900 3620 113100 3880
rect 113400 3620 113600 3880
rect 113900 3620 114100 3880
rect 114400 3620 114600 3880
rect 114900 3620 115100 3880
rect 115400 3620 115600 3880
rect 115900 3620 116100 3880
rect 116400 3620 116600 3880
rect 116900 3620 117100 3880
rect 117400 3620 117600 3880
rect 117900 3620 118100 3880
rect 118400 3620 118600 3880
rect 118900 3620 119100 3880
rect 119400 3620 119600 3880
rect 119900 3620 120100 3880
rect 120400 3620 120600 3880
rect 120900 3620 121100 3880
rect 121400 3620 121600 3880
rect 121900 3620 122100 3880
rect 122400 3620 122600 3880
rect 122900 3620 123100 3880
rect 123400 3620 123600 3880
rect 123900 3620 124100 3880
rect 124400 3620 124600 3880
rect 124900 3620 125100 3880
rect 125400 3620 125600 3880
rect 125900 3620 126100 3880
rect 126400 3620 126600 3880
rect 126900 3620 127100 3880
rect 127400 3620 127600 3880
rect 127900 3620 128000 3880
rect 104000 3600 104120 3620
rect 104380 3600 104620 3620
rect 104880 3600 105120 3620
rect 105380 3600 105620 3620
rect 105880 3600 106120 3620
rect 106380 3600 106620 3620
rect 106880 3600 107120 3620
rect 107380 3600 107620 3620
rect 107880 3600 108120 3620
rect 108380 3600 108620 3620
rect 108880 3600 109120 3620
rect 109380 3600 109620 3620
rect 109880 3600 110120 3620
rect 110380 3600 110620 3620
rect 110880 3600 111120 3620
rect 111380 3600 111620 3620
rect 111880 3600 112120 3620
rect 112380 3600 112620 3620
rect 112880 3600 113120 3620
rect 113380 3600 113620 3620
rect 113880 3600 114120 3620
rect 114380 3600 114620 3620
rect 114880 3600 115120 3620
rect 115380 3600 115620 3620
rect 115880 3600 116120 3620
rect 116380 3600 116620 3620
rect 116880 3600 117120 3620
rect 117380 3600 117620 3620
rect 117880 3600 118120 3620
rect 118380 3600 118620 3620
rect 118880 3600 119120 3620
rect 119380 3600 119620 3620
rect 119880 3600 120120 3620
rect 120380 3600 120620 3620
rect 120880 3600 121120 3620
rect 121380 3600 121620 3620
rect 121880 3600 122120 3620
rect 122380 3600 122620 3620
rect 122880 3600 123120 3620
rect 123380 3600 123620 3620
rect 123880 3600 124120 3620
rect 124380 3600 124620 3620
rect 124880 3600 125120 3620
rect 125380 3600 125620 3620
rect 125880 3600 126120 3620
rect 126380 3600 126620 3620
rect 126880 3600 127120 3620
rect 127380 3600 127620 3620
rect 127880 3600 128000 3620
rect 104000 3400 128000 3600
rect 104000 3380 104120 3400
rect 104380 3380 104620 3400
rect 104880 3380 105120 3400
rect 105380 3380 105620 3400
rect 105880 3380 106120 3400
rect 106380 3380 106620 3400
rect 106880 3380 107120 3400
rect 107380 3380 107620 3400
rect 107880 3380 108120 3400
rect 108380 3380 108620 3400
rect 108880 3380 109120 3400
rect 109380 3380 109620 3400
rect 109880 3380 110120 3400
rect 110380 3380 110620 3400
rect 110880 3380 111120 3400
rect 111380 3380 111620 3400
rect 111880 3380 112120 3400
rect 112380 3380 112620 3400
rect 112880 3380 113120 3400
rect 113380 3380 113620 3400
rect 113880 3380 114120 3400
rect 114380 3380 114620 3400
rect 114880 3380 115120 3400
rect 115380 3380 115620 3400
rect 115880 3380 116120 3400
rect 116380 3380 116620 3400
rect 116880 3380 117120 3400
rect 117380 3380 117620 3400
rect 117880 3380 118120 3400
rect 118380 3380 118620 3400
rect 118880 3380 119120 3400
rect 119380 3380 119620 3400
rect 119880 3380 120120 3400
rect 120380 3380 120620 3400
rect 120880 3380 121120 3400
rect 121380 3380 121620 3400
rect 121880 3380 122120 3400
rect 122380 3380 122620 3400
rect 122880 3380 123120 3400
rect 123380 3380 123620 3400
rect 123880 3380 124120 3400
rect 124380 3380 124620 3400
rect 124880 3380 125120 3400
rect 125380 3380 125620 3400
rect 125880 3380 126120 3400
rect 126380 3380 126620 3400
rect 126880 3380 127120 3400
rect 127380 3380 127620 3400
rect 127880 3380 128000 3400
rect 104000 3120 104100 3380
rect 104400 3120 104600 3380
rect 104900 3120 105100 3380
rect 105400 3120 105600 3380
rect 105900 3120 106100 3380
rect 106400 3120 106600 3380
rect 106900 3120 107100 3380
rect 107400 3120 107600 3380
rect 107900 3120 108100 3380
rect 108400 3120 108600 3380
rect 108900 3120 109100 3380
rect 109400 3120 109600 3380
rect 109900 3120 110100 3380
rect 110400 3120 110600 3380
rect 110900 3120 111100 3380
rect 111400 3120 111600 3380
rect 111900 3120 112100 3380
rect 112400 3120 112600 3380
rect 112900 3120 113100 3380
rect 113400 3120 113600 3380
rect 113900 3120 114100 3380
rect 114400 3120 114600 3380
rect 114900 3120 115100 3380
rect 115400 3120 115600 3380
rect 115900 3120 116100 3380
rect 116400 3120 116600 3380
rect 116900 3120 117100 3380
rect 117400 3120 117600 3380
rect 117900 3120 118100 3380
rect 118400 3120 118600 3380
rect 118900 3120 119100 3380
rect 119400 3120 119600 3380
rect 119900 3120 120100 3380
rect 120400 3120 120600 3380
rect 120900 3120 121100 3380
rect 121400 3120 121600 3380
rect 121900 3120 122100 3380
rect 122400 3120 122600 3380
rect 122900 3120 123100 3380
rect 123400 3120 123600 3380
rect 123900 3120 124100 3380
rect 124400 3120 124600 3380
rect 124900 3120 125100 3380
rect 125400 3120 125600 3380
rect 125900 3120 126100 3380
rect 126400 3120 126600 3380
rect 126900 3120 127100 3380
rect 127400 3120 127600 3380
rect 127900 3120 128000 3380
rect 104000 3100 104120 3120
rect 104380 3100 104620 3120
rect 104880 3100 105120 3120
rect 105380 3100 105620 3120
rect 105880 3100 106120 3120
rect 106380 3100 106620 3120
rect 106880 3100 107120 3120
rect 107380 3100 107620 3120
rect 107880 3100 108120 3120
rect 108380 3100 108620 3120
rect 108880 3100 109120 3120
rect 109380 3100 109620 3120
rect 109880 3100 110120 3120
rect 110380 3100 110620 3120
rect 110880 3100 111120 3120
rect 111380 3100 111620 3120
rect 111880 3100 112120 3120
rect 112380 3100 112620 3120
rect 112880 3100 113120 3120
rect 113380 3100 113620 3120
rect 113880 3100 114120 3120
rect 114380 3100 114620 3120
rect 114880 3100 115120 3120
rect 115380 3100 115620 3120
rect 115880 3100 116120 3120
rect 116380 3100 116620 3120
rect 116880 3100 117120 3120
rect 117380 3100 117620 3120
rect 117880 3100 118120 3120
rect 118380 3100 118620 3120
rect 118880 3100 119120 3120
rect 119380 3100 119620 3120
rect 119880 3100 120120 3120
rect 120380 3100 120620 3120
rect 120880 3100 121120 3120
rect 121380 3100 121620 3120
rect 121880 3100 122120 3120
rect 122380 3100 122620 3120
rect 122880 3100 123120 3120
rect 123380 3100 123620 3120
rect 123880 3100 124120 3120
rect 124380 3100 124620 3120
rect 124880 3100 125120 3120
rect 125380 3100 125620 3120
rect 125880 3100 126120 3120
rect 126380 3100 126620 3120
rect 126880 3100 127120 3120
rect 127380 3100 127620 3120
rect 127880 3100 128000 3120
rect 104000 2900 128000 3100
rect 104000 2880 104120 2900
rect 104380 2880 104620 2900
rect 104880 2880 105120 2900
rect 105380 2880 105620 2900
rect 105880 2880 106120 2900
rect 106380 2880 106620 2900
rect 106880 2880 107120 2900
rect 107380 2880 107620 2900
rect 107880 2880 108120 2900
rect 108380 2880 108620 2900
rect 108880 2880 109120 2900
rect 109380 2880 109620 2900
rect 109880 2880 110120 2900
rect 110380 2880 110620 2900
rect 110880 2880 111120 2900
rect 111380 2880 111620 2900
rect 111880 2880 112120 2900
rect 112380 2880 112620 2900
rect 112880 2880 113120 2900
rect 113380 2880 113620 2900
rect 113880 2880 114120 2900
rect 114380 2880 114620 2900
rect 114880 2880 115120 2900
rect 115380 2880 115620 2900
rect 115880 2880 116120 2900
rect 116380 2880 116620 2900
rect 116880 2880 117120 2900
rect 117380 2880 117620 2900
rect 117880 2880 118120 2900
rect 118380 2880 118620 2900
rect 118880 2880 119120 2900
rect 119380 2880 119620 2900
rect 119880 2880 120120 2900
rect 120380 2880 120620 2900
rect 120880 2880 121120 2900
rect 121380 2880 121620 2900
rect 121880 2880 122120 2900
rect 122380 2880 122620 2900
rect 122880 2880 123120 2900
rect 123380 2880 123620 2900
rect 123880 2880 124120 2900
rect 124380 2880 124620 2900
rect 124880 2880 125120 2900
rect 125380 2880 125620 2900
rect 125880 2880 126120 2900
rect 126380 2880 126620 2900
rect 126880 2880 127120 2900
rect 127380 2880 127620 2900
rect 127880 2880 128000 2900
rect 104000 2620 104100 2880
rect 104400 2620 104600 2880
rect 104900 2620 105100 2880
rect 105400 2620 105600 2880
rect 105900 2620 106100 2880
rect 106400 2620 106600 2880
rect 106900 2620 107100 2880
rect 107400 2620 107600 2880
rect 107900 2620 108100 2880
rect 108400 2620 108600 2880
rect 108900 2620 109100 2880
rect 109400 2620 109600 2880
rect 109900 2620 110100 2880
rect 110400 2620 110600 2880
rect 110900 2620 111100 2880
rect 111400 2620 111600 2880
rect 111900 2620 112100 2880
rect 112400 2620 112600 2880
rect 112900 2620 113100 2880
rect 113400 2620 113600 2880
rect 113900 2620 114100 2880
rect 114400 2620 114600 2880
rect 114900 2620 115100 2880
rect 115400 2620 115600 2880
rect 115900 2620 116100 2880
rect 116400 2620 116600 2880
rect 116900 2620 117100 2880
rect 117400 2620 117600 2880
rect 117900 2620 118100 2880
rect 118400 2620 118600 2880
rect 118900 2620 119100 2880
rect 119400 2620 119600 2880
rect 119900 2620 120100 2880
rect 120400 2620 120600 2880
rect 120900 2620 121100 2880
rect 121400 2620 121600 2880
rect 121900 2620 122100 2880
rect 122400 2620 122600 2880
rect 122900 2620 123100 2880
rect 123400 2620 123600 2880
rect 123900 2620 124100 2880
rect 124400 2620 124600 2880
rect 124900 2620 125100 2880
rect 125400 2620 125600 2880
rect 125900 2620 126100 2880
rect 126400 2620 126600 2880
rect 126900 2620 127100 2880
rect 127400 2620 127600 2880
rect 127900 2620 128000 2880
rect 104000 2600 104120 2620
rect 104380 2600 104620 2620
rect 104880 2600 105120 2620
rect 105380 2600 105620 2620
rect 105880 2600 106120 2620
rect 106380 2600 106620 2620
rect 106880 2600 107120 2620
rect 107380 2600 107620 2620
rect 107880 2600 108120 2620
rect 108380 2600 108620 2620
rect 108880 2600 109120 2620
rect 109380 2600 109620 2620
rect 109880 2600 110120 2620
rect 110380 2600 110620 2620
rect 110880 2600 111120 2620
rect 111380 2600 111620 2620
rect 111880 2600 112120 2620
rect 112380 2600 112620 2620
rect 112880 2600 113120 2620
rect 113380 2600 113620 2620
rect 113880 2600 114120 2620
rect 114380 2600 114620 2620
rect 114880 2600 115120 2620
rect 115380 2600 115620 2620
rect 115880 2600 116120 2620
rect 116380 2600 116620 2620
rect 116880 2600 117120 2620
rect 117380 2600 117620 2620
rect 117880 2600 118120 2620
rect 118380 2600 118620 2620
rect 118880 2600 119120 2620
rect 119380 2600 119620 2620
rect 119880 2600 120120 2620
rect 120380 2600 120620 2620
rect 120880 2600 121120 2620
rect 121380 2600 121620 2620
rect 121880 2600 122120 2620
rect 122380 2600 122620 2620
rect 122880 2600 123120 2620
rect 123380 2600 123620 2620
rect 123880 2600 124120 2620
rect 124380 2600 124620 2620
rect 124880 2600 125120 2620
rect 125380 2600 125620 2620
rect 125880 2600 126120 2620
rect 126380 2600 126620 2620
rect 126880 2600 127120 2620
rect 127380 2600 127620 2620
rect 127880 2600 128000 2620
rect 104000 2400 128000 2600
rect 104000 2380 104120 2400
rect 104380 2380 104620 2400
rect 104880 2380 105120 2400
rect 105380 2380 105620 2400
rect 105880 2380 106120 2400
rect 106380 2380 106620 2400
rect 106880 2380 107120 2400
rect 107380 2380 107620 2400
rect 107880 2380 108120 2400
rect 108380 2380 108620 2400
rect 108880 2380 109120 2400
rect 109380 2380 109620 2400
rect 109880 2380 110120 2400
rect 110380 2380 110620 2400
rect 110880 2380 111120 2400
rect 111380 2380 111620 2400
rect 111880 2380 112120 2400
rect 112380 2380 112620 2400
rect 112880 2380 113120 2400
rect 113380 2380 113620 2400
rect 113880 2380 114120 2400
rect 114380 2380 114620 2400
rect 114880 2380 115120 2400
rect 115380 2380 115620 2400
rect 115880 2380 116120 2400
rect 116380 2380 116620 2400
rect 116880 2380 117120 2400
rect 117380 2380 117620 2400
rect 117880 2380 118120 2400
rect 118380 2380 118620 2400
rect 118880 2380 119120 2400
rect 119380 2380 119620 2400
rect 119880 2380 120120 2400
rect 120380 2380 120620 2400
rect 120880 2380 121120 2400
rect 121380 2380 121620 2400
rect 121880 2380 122120 2400
rect 122380 2380 122620 2400
rect 122880 2380 123120 2400
rect 123380 2380 123620 2400
rect 123880 2380 124120 2400
rect 124380 2380 124620 2400
rect 124880 2380 125120 2400
rect 125380 2380 125620 2400
rect 125880 2380 126120 2400
rect 126380 2380 126620 2400
rect 126880 2380 127120 2400
rect 127380 2380 127620 2400
rect 127880 2380 128000 2400
rect 104000 2120 104100 2380
rect 104400 2120 104600 2380
rect 104900 2120 105100 2380
rect 105400 2120 105600 2380
rect 105900 2120 106100 2380
rect 106400 2120 106600 2380
rect 106900 2120 107100 2380
rect 107400 2120 107600 2380
rect 107900 2120 108100 2380
rect 108400 2120 108600 2380
rect 108900 2120 109100 2380
rect 109400 2120 109600 2380
rect 109900 2120 110100 2380
rect 110400 2120 110600 2380
rect 110900 2120 111100 2380
rect 111400 2120 111600 2380
rect 111900 2120 112100 2380
rect 112400 2120 112600 2380
rect 112900 2120 113100 2380
rect 113400 2120 113600 2380
rect 113900 2120 114100 2380
rect 114400 2120 114600 2380
rect 114900 2120 115100 2380
rect 115400 2120 115600 2380
rect 115900 2120 116100 2380
rect 116400 2120 116600 2380
rect 116900 2120 117100 2380
rect 117400 2120 117600 2380
rect 117900 2120 118100 2380
rect 118400 2120 118600 2380
rect 118900 2120 119100 2380
rect 119400 2120 119600 2380
rect 119900 2120 120100 2380
rect 120400 2120 120600 2380
rect 120900 2120 121100 2380
rect 121400 2120 121600 2380
rect 121900 2120 122100 2380
rect 122400 2120 122600 2380
rect 122900 2120 123100 2380
rect 123400 2120 123600 2380
rect 123900 2120 124100 2380
rect 124400 2120 124600 2380
rect 124900 2120 125100 2380
rect 125400 2120 125600 2380
rect 125900 2120 126100 2380
rect 126400 2120 126600 2380
rect 126900 2120 127100 2380
rect 127400 2120 127600 2380
rect 127900 2120 128000 2380
rect 104000 2100 104120 2120
rect 104380 2100 104620 2120
rect 104880 2100 105120 2120
rect 105380 2100 105620 2120
rect 105880 2100 106120 2120
rect 106380 2100 106620 2120
rect 106880 2100 107120 2120
rect 107380 2100 107620 2120
rect 107880 2100 108120 2120
rect 108380 2100 108620 2120
rect 108880 2100 109120 2120
rect 109380 2100 109620 2120
rect 109880 2100 110120 2120
rect 110380 2100 110620 2120
rect 110880 2100 111120 2120
rect 111380 2100 111620 2120
rect 111880 2100 112120 2120
rect 112380 2100 112620 2120
rect 112880 2100 113120 2120
rect 113380 2100 113620 2120
rect 113880 2100 114120 2120
rect 114380 2100 114620 2120
rect 114880 2100 115120 2120
rect 115380 2100 115620 2120
rect 115880 2100 116120 2120
rect 116380 2100 116620 2120
rect 116880 2100 117120 2120
rect 117380 2100 117620 2120
rect 117880 2100 118120 2120
rect 118380 2100 118620 2120
rect 118880 2100 119120 2120
rect 119380 2100 119620 2120
rect 119880 2100 120120 2120
rect 120380 2100 120620 2120
rect 120880 2100 121120 2120
rect 121380 2100 121620 2120
rect 121880 2100 122120 2120
rect 122380 2100 122620 2120
rect 122880 2100 123120 2120
rect 123380 2100 123620 2120
rect 123880 2100 124120 2120
rect 124380 2100 124620 2120
rect 124880 2100 125120 2120
rect 125380 2100 125620 2120
rect 125880 2100 126120 2120
rect 126380 2100 126620 2120
rect 126880 2100 127120 2120
rect 127380 2100 127620 2120
rect 127880 2100 128000 2120
rect 104000 2000 128000 2100
rect 136000 5980 140000 6000
rect 136000 5910 136150 5980
rect 136350 5910 136650 5980
rect 136850 5910 137150 5980
rect 137350 5910 137650 5980
rect 137850 5910 138150 5980
rect 138350 5910 138650 5980
rect 138850 5910 139150 5980
rect 139350 5910 139650 5980
rect 139850 5910 140000 5980
rect 136000 5900 140000 5910
rect 136000 5880 136120 5900
rect 136380 5880 136620 5900
rect 136880 5880 137120 5900
rect 137380 5880 137620 5900
rect 137880 5880 138120 5900
rect 138380 5880 138620 5900
rect 138880 5880 139120 5900
rect 139380 5880 139620 5900
rect 139880 5880 140000 5900
rect 136000 5850 136100 5880
rect 136000 5650 136020 5850
rect 136090 5650 136100 5850
rect 136000 5620 136100 5650
rect 136400 5850 136600 5880
rect 136400 5650 136410 5850
rect 136480 5650 136520 5850
rect 136590 5650 136600 5850
rect 136400 5620 136600 5650
rect 136900 5850 137100 5880
rect 136900 5650 136910 5850
rect 136980 5650 137020 5850
rect 137090 5650 137100 5850
rect 136900 5620 137100 5650
rect 137400 5850 137600 5880
rect 137400 5650 137410 5850
rect 137480 5650 137520 5850
rect 137590 5650 137600 5850
rect 137400 5620 137600 5650
rect 137900 5850 138100 5880
rect 137900 5650 137910 5850
rect 137980 5650 138020 5850
rect 138090 5650 138100 5850
rect 137900 5620 138100 5650
rect 138400 5850 138600 5880
rect 138400 5650 138410 5850
rect 138480 5650 138520 5850
rect 138590 5650 138600 5850
rect 138400 5620 138600 5650
rect 138900 5850 139100 5880
rect 138900 5650 138910 5850
rect 138980 5650 139020 5850
rect 139090 5650 139100 5850
rect 138900 5620 139100 5650
rect 139400 5850 139600 5880
rect 139400 5650 139410 5850
rect 139480 5650 139520 5850
rect 139590 5650 139600 5850
rect 139400 5620 139600 5650
rect 139900 5850 140000 5880
rect 139900 5650 139910 5850
rect 139980 5650 140000 5850
rect 139900 5620 140000 5650
rect 136000 5600 136120 5620
rect 136380 5600 136620 5620
rect 136880 5600 137120 5620
rect 137380 5600 137620 5620
rect 137880 5600 138120 5620
rect 138380 5600 138620 5620
rect 138880 5600 139120 5620
rect 139380 5600 139620 5620
rect 139880 5600 140000 5620
rect 136000 5590 140000 5600
rect 136000 5520 136150 5590
rect 136350 5520 136650 5590
rect 136850 5520 137150 5590
rect 137350 5520 137650 5590
rect 137850 5520 138150 5590
rect 138350 5520 138650 5590
rect 138850 5520 139150 5590
rect 139350 5520 139650 5590
rect 139850 5520 140000 5590
rect 136000 5480 140000 5520
rect 136000 5410 136150 5480
rect 136350 5410 136650 5480
rect 136850 5410 137150 5480
rect 137350 5410 137650 5480
rect 137850 5410 138150 5480
rect 138350 5410 138650 5480
rect 138850 5410 139150 5480
rect 139350 5410 139650 5480
rect 139850 5410 140000 5480
rect 136000 5400 140000 5410
rect 136000 5380 136120 5400
rect 136380 5380 136620 5400
rect 136880 5380 137120 5400
rect 137380 5380 137620 5400
rect 137880 5380 138120 5400
rect 138380 5380 138620 5400
rect 138880 5380 139120 5400
rect 139380 5380 139620 5400
rect 139880 5380 140000 5400
rect 136000 5350 136100 5380
rect 136000 5150 136020 5350
rect 136090 5150 136100 5350
rect 136000 5120 136100 5150
rect 136400 5350 136600 5380
rect 136400 5150 136410 5350
rect 136480 5150 136520 5350
rect 136590 5150 136600 5350
rect 136400 5120 136600 5150
rect 136900 5350 137100 5380
rect 136900 5150 136910 5350
rect 136980 5150 137020 5350
rect 137090 5150 137100 5350
rect 136900 5120 137100 5150
rect 137400 5350 137600 5380
rect 137400 5150 137410 5350
rect 137480 5150 137520 5350
rect 137590 5150 137600 5350
rect 137400 5120 137600 5150
rect 137900 5350 138100 5380
rect 137900 5150 137910 5350
rect 137980 5150 138020 5350
rect 138090 5150 138100 5350
rect 137900 5120 138100 5150
rect 138400 5350 138600 5380
rect 138400 5150 138410 5350
rect 138480 5150 138520 5350
rect 138590 5150 138600 5350
rect 138400 5120 138600 5150
rect 138900 5350 139100 5380
rect 138900 5150 138910 5350
rect 138980 5150 139020 5350
rect 139090 5150 139100 5350
rect 138900 5120 139100 5150
rect 139400 5350 139600 5380
rect 139400 5150 139410 5350
rect 139480 5150 139520 5350
rect 139590 5150 139600 5350
rect 139400 5120 139600 5150
rect 139900 5350 140000 5380
rect 139900 5150 139910 5350
rect 139980 5150 140000 5350
rect 139900 5120 140000 5150
rect 136000 5100 136120 5120
rect 136380 5100 136620 5120
rect 136880 5100 137120 5120
rect 137380 5100 137620 5120
rect 137880 5100 138120 5120
rect 138380 5100 138620 5120
rect 138880 5100 139120 5120
rect 139380 5100 139620 5120
rect 139880 5100 140000 5120
rect 136000 5090 140000 5100
rect 136000 5020 136150 5090
rect 136350 5020 136650 5090
rect 136850 5020 137150 5090
rect 137350 5020 137650 5090
rect 137850 5020 138150 5090
rect 138350 5020 138650 5090
rect 138850 5020 139150 5090
rect 139350 5020 139650 5090
rect 139850 5020 140000 5090
rect 136000 4980 140000 5020
rect 136000 4910 136150 4980
rect 136350 4910 136650 4980
rect 136850 4910 137150 4980
rect 137350 4910 137650 4980
rect 137850 4910 138150 4980
rect 138350 4910 138650 4980
rect 138850 4910 139150 4980
rect 139350 4910 139650 4980
rect 139850 4910 140000 4980
rect 136000 4900 140000 4910
rect 136000 4880 136120 4900
rect 136380 4880 136620 4900
rect 136880 4880 137120 4900
rect 137380 4880 137620 4900
rect 137880 4880 138120 4900
rect 138380 4880 138620 4900
rect 138880 4880 139120 4900
rect 139380 4880 139620 4900
rect 139880 4880 140000 4900
rect 136000 4850 136100 4880
rect 136000 4650 136020 4850
rect 136090 4650 136100 4850
rect 136000 4620 136100 4650
rect 136400 4850 136600 4880
rect 136400 4650 136410 4850
rect 136480 4650 136520 4850
rect 136590 4650 136600 4850
rect 136400 4620 136600 4650
rect 136900 4850 137100 4880
rect 136900 4650 136910 4850
rect 136980 4650 137020 4850
rect 137090 4650 137100 4850
rect 136900 4620 137100 4650
rect 137400 4850 137600 4880
rect 137400 4650 137410 4850
rect 137480 4650 137520 4850
rect 137590 4650 137600 4850
rect 137400 4620 137600 4650
rect 137900 4850 138100 4880
rect 137900 4650 137910 4850
rect 137980 4650 138020 4850
rect 138090 4650 138100 4850
rect 137900 4620 138100 4650
rect 138400 4850 138600 4880
rect 138400 4650 138410 4850
rect 138480 4650 138520 4850
rect 138590 4650 138600 4850
rect 138400 4620 138600 4650
rect 138900 4850 139100 4880
rect 138900 4650 138910 4850
rect 138980 4650 139020 4850
rect 139090 4650 139100 4850
rect 138900 4620 139100 4650
rect 139400 4850 139600 4880
rect 139400 4650 139410 4850
rect 139480 4650 139520 4850
rect 139590 4650 139600 4850
rect 139400 4620 139600 4650
rect 139900 4850 140000 4880
rect 139900 4650 139910 4850
rect 139980 4650 140000 4850
rect 139900 4620 140000 4650
rect 136000 4600 136120 4620
rect 136380 4600 136620 4620
rect 136880 4600 137120 4620
rect 137380 4600 137620 4620
rect 137880 4600 138120 4620
rect 138380 4600 138620 4620
rect 138880 4600 139120 4620
rect 139380 4600 139620 4620
rect 139880 4600 140000 4620
rect 136000 4590 140000 4600
rect 136000 4520 136150 4590
rect 136350 4520 136650 4590
rect 136850 4520 137150 4590
rect 137350 4520 137650 4590
rect 137850 4520 138150 4590
rect 138350 4520 138650 4590
rect 138850 4520 139150 4590
rect 139350 4520 139650 4590
rect 139850 4520 140000 4590
rect 136000 4480 140000 4520
rect 136000 4410 136150 4480
rect 136350 4410 136650 4480
rect 136850 4410 137150 4480
rect 137350 4410 137650 4480
rect 137850 4410 138150 4480
rect 138350 4410 138650 4480
rect 138850 4410 139150 4480
rect 139350 4410 139650 4480
rect 139850 4410 140000 4480
rect 136000 4400 140000 4410
rect 136000 4380 136120 4400
rect 136380 4380 136620 4400
rect 136880 4380 137120 4400
rect 137380 4380 137620 4400
rect 137880 4380 138120 4400
rect 138380 4380 138620 4400
rect 138880 4380 139120 4400
rect 139380 4380 139620 4400
rect 139880 4380 140000 4400
rect 136000 4350 136100 4380
rect 136000 4150 136020 4350
rect 136090 4150 136100 4350
rect 136000 4120 136100 4150
rect 136400 4350 136600 4380
rect 136400 4150 136410 4350
rect 136480 4150 136520 4350
rect 136590 4150 136600 4350
rect 136400 4120 136600 4150
rect 136900 4350 137100 4380
rect 136900 4150 136910 4350
rect 136980 4150 137020 4350
rect 137090 4150 137100 4350
rect 136900 4120 137100 4150
rect 137400 4350 137600 4380
rect 137400 4150 137410 4350
rect 137480 4150 137520 4350
rect 137590 4150 137600 4350
rect 137400 4120 137600 4150
rect 137900 4350 138100 4380
rect 137900 4150 137910 4350
rect 137980 4150 138020 4350
rect 138090 4150 138100 4350
rect 137900 4120 138100 4150
rect 138400 4350 138600 4380
rect 138400 4150 138410 4350
rect 138480 4150 138520 4350
rect 138590 4150 138600 4350
rect 138400 4120 138600 4150
rect 138900 4350 139100 4380
rect 138900 4150 138910 4350
rect 138980 4150 139020 4350
rect 139090 4150 139100 4350
rect 138900 4120 139100 4150
rect 139400 4350 139600 4380
rect 139400 4150 139410 4350
rect 139480 4150 139520 4350
rect 139590 4150 139600 4350
rect 139400 4120 139600 4150
rect 139900 4350 140000 4380
rect 139900 4150 139910 4350
rect 139980 4150 140000 4350
rect 139900 4120 140000 4150
rect 136000 4100 136120 4120
rect 136380 4100 136620 4120
rect 136880 4100 137120 4120
rect 137380 4100 137620 4120
rect 137880 4100 138120 4120
rect 138380 4100 138620 4120
rect 138880 4100 139120 4120
rect 139380 4100 139620 4120
rect 139880 4100 140000 4120
rect 136000 4090 140000 4100
rect 136000 4020 136150 4090
rect 136350 4020 136650 4090
rect 136850 4020 137150 4090
rect 137350 4020 137650 4090
rect 137850 4020 138150 4090
rect 138350 4020 138650 4090
rect 138850 4020 139150 4090
rect 139350 4020 139650 4090
rect 139850 4020 140000 4090
rect 136000 3980 140000 4020
rect 136000 3910 136150 3980
rect 136350 3910 136650 3980
rect 136850 3910 137150 3980
rect 137350 3910 137650 3980
rect 137850 3910 138150 3980
rect 138350 3910 138650 3980
rect 138850 3910 139150 3980
rect 139350 3910 139650 3980
rect 139850 3910 140000 3980
rect 136000 3900 140000 3910
rect 136000 3880 136120 3900
rect 136380 3880 136620 3900
rect 136880 3880 137120 3900
rect 137380 3880 137620 3900
rect 137880 3880 138120 3900
rect 138380 3880 138620 3900
rect 138880 3880 139120 3900
rect 139380 3880 139620 3900
rect 139880 3880 140000 3900
rect 136000 3850 136100 3880
rect 136000 3650 136020 3850
rect 136090 3650 136100 3850
rect 136000 3620 136100 3650
rect 136400 3850 136600 3880
rect 136400 3650 136410 3850
rect 136480 3650 136520 3850
rect 136590 3650 136600 3850
rect 136400 3620 136600 3650
rect 136900 3850 137100 3880
rect 136900 3650 136910 3850
rect 136980 3650 137020 3850
rect 137090 3650 137100 3850
rect 136900 3620 137100 3650
rect 137400 3850 137600 3880
rect 137400 3650 137410 3850
rect 137480 3650 137520 3850
rect 137590 3650 137600 3850
rect 137400 3620 137600 3650
rect 137900 3850 138100 3880
rect 137900 3650 137910 3850
rect 137980 3650 138020 3850
rect 138090 3650 138100 3850
rect 137900 3620 138100 3650
rect 138400 3850 138600 3880
rect 138400 3650 138410 3850
rect 138480 3650 138520 3850
rect 138590 3650 138600 3850
rect 138400 3620 138600 3650
rect 138900 3850 139100 3880
rect 138900 3650 138910 3850
rect 138980 3650 139020 3850
rect 139090 3650 139100 3850
rect 138900 3620 139100 3650
rect 139400 3850 139600 3880
rect 139400 3650 139410 3850
rect 139480 3650 139520 3850
rect 139590 3650 139600 3850
rect 139400 3620 139600 3650
rect 139900 3850 140000 3880
rect 139900 3650 139910 3850
rect 139980 3650 140000 3850
rect 139900 3620 140000 3650
rect 136000 3600 136120 3620
rect 136380 3600 136620 3620
rect 136880 3600 137120 3620
rect 137380 3600 137620 3620
rect 137880 3600 138120 3620
rect 138380 3600 138620 3620
rect 138880 3600 139120 3620
rect 139380 3600 139620 3620
rect 139880 3600 140000 3620
rect 136000 3590 140000 3600
rect 136000 3520 136150 3590
rect 136350 3520 136650 3590
rect 136850 3520 137150 3590
rect 137350 3520 137650 3590
rect 137850 3520 138150 3590
rect 138350 3520 138650 3590
rect 138850 3520 139150 3590
rect 139350 3520 139650 3590
rect 139850 3520 140000 3590
rect 136000 3480 140000 3520
rect 136000 3410 136150 3480
rect 136350 3410 136650 3480
rect 136850 3410 137150 3480
rect 137350 3410 137650 3480
rect 137850 3410 138150 3480
rect 138350 3410 138650 3480
rect 138850 3410 139150 3480
rect 139350 3410 139650 3480
rect 139850 3410 140000 3480
rect 136000 3400 140000 3410
rect 136000 3380 136120 3400
rect 136380 3380 136620 3400
rect 136880 3380 137120 3400
rect 137380 3380 137620 3400
rect 137880 3380 138120 3400
rect 138380 3380 138620 3400
rect 138880 3380 139120 3400
rect 139380 3380 139620 3400
rect 139880 3380 140000 3400
rect 136000 3350 136100 3380
rect 136000 3150 136020 3350
rect 136090 3150 136100 3350
rect 136000 3120 136100 3150
rect 136400 3350 136600 3380
rect 136400 3150 136410 3350
rect 136480 3150 136520 3350
rect 136590 3150 136600 3350
rect 136400 3120 136600 3150
rect 136900 3350 137100 3380
rect 136900 3150 136910 3350
rect 136980 3150 137020 3350
rect 137090 3150 137100 3350
rect 136900 3120 137100 3150
rect 137400 3350 137600 3380
rect 137400 3150 137410 3350
rect 137480 3150 137520 3350
rect 137590 3150 137600 3350
rect 137400 3120 137600 3150
rect 137900 3350 138100 3380
rect 137900 3150 137910 3350
rect 137980 3150 138020 3350
rect 138090 3150 138100 3350
rect 137900 3120 138100 3150
rect 138400 3350 138600 3380
rect 138400 3150 138410 3350
rect 138480 3150 138520 3350
rect 138590 3150 138600 3350
rect 138400 3120 138600 3150
rect 138900 3350 139100 3380
rect 138900 3150 138910 3350
rect 138980 3150 139020 3350
rect 139090 3150 139100 3350
rect 138900 3120 139100 3150
rect 139400 3350 139600 3380
rect 139400 3150 139410 3350
rect 139480 3150 139520 3350
rect 139590 3150 139600 3350
rect 139400 3120 139600 3150
rect 139900 3350 140000 3380
rect 139900 3150 139910 3350
rect 139980 3150 140000 3350
rect 139900 3120 140000 3150
rect 136000 3100 136120 3120
rect 136380 3100 136620 3120
rect 136880 3100 137120 3120
rect 137380 3100 137620 3120
rect 137880 3100 138120 3120
rect 138380 3100 138620 3120
rect 138880 3100 139120 3120
rect 139380 3100 139620 3120
rect 139880 3100 140000 3120
rect 136000 3090 140000 3100
rect 136000 3020 136150 3090
rect 136350 3020 136650 3090
rect 136850 3020 137150 3090
rect 137350 3020 137650 3090
rect 137850 3020 138150 3090
rect 138350 3020 138650 3090
rect 138850 3020 139150 3090
rect 139350 3020 139650 3090
rect 139850 3020 140000 3090
rect 136000 2980 140000 3020
rect 136000 2910 136150 2980
rect 136350 2910 136650 2980
rect 136850 2910 137150 2980
rect 137350 2910 137650 2980
rect 137850 2910 138150 2980
rect 138350 2910 138650 2980
rect 138850 2910 139150 2980
rect 139350 2910 139650 2980
rect 139850 2910 140000 2980
rect 136000 2900 140000 2910
rect 136000 2880 136120 2900
rect 136380 2880 136620 2900
rect 136880 2880 137120 2900
rect 137380 2880 137620 2900
rect 137880 2880 138120 2900
rect 138380 2880 138620 2900
rect 138880 2880 139120 2900
rect 139380 2880 139620 2900
rect 139880 2880 140000 2900
rect 136000 2850 136100 2880
rect 136000 2650 136020 2850
rect 136090 2650 136100 2850
rect 136000 2620 136100 2650
rect 136400 2850 136600 2880
rect 136400 2650 136410 2850
rect 136480 2650 136520 2850
rect 136590 2650 136600 2850
rect 136400 2620 136600 2650
rect 136900 2850 137100 2880
rect 136900 2650 136910 2850
rect 136980 2650 137020 2850
rect 137090 2650 137100 2850
rect 136900 2620 137100 2650
rect 137400 2850 137600 2880
rect 137400 2650 137410 2850
rect 137480 2650 137520 2850
rect 137590 2650 137600 2850
rect 137400 2620 137600 2650
rect 137900 2850 138100 2880
rect 137900 2650 137910 2850
rect 137980 2650 138020 2850
rect 138090 2650 138100 2850
rect 137900 2620 138100 2650
rect 138400 2850 138600 2880
rect 138400 2650 138410 2850
rect 138480 2650 138520 2850
rect 138590 2650 138600 2850
rect 138400 2620 138600 2650
rect 138900 2850 139100 2880
rect 138900 2650 138910 2850
rect 138980 2650 139020 2850
rect 139090 2650 139100 2850
rect 138900 2620 139100 2650
rect 139400 2850 139600 2880
rect 139400 2650 139410 2850
rect 139480 2650 139520 2850
rect 139590 2650 139600 2850
rect 139400 2620 139600 2650
rect 139900 2850 140000 2880
rect 139900 2650 139910 2850
rect 139980 2650 140000 2850
rect 139900 2620 140000 2650
rect 136000 2600 136120 2620
rect 136380 2600 136620 2620
rect 136880 2600 137120 2620
rect 137380 2600 137620 2620
rect 137880 2600 138120 2620
rect 138380 2600 138620 2620
rect 138880 2600 139120 2620
rect 139380 2600 139620 2620
rect 139880 2600 140000 2620
rect 136000 2590 140000 2600
rect 136000 2520 136150 2590
rect 136350 2520 136650 2590
rect 136850 2520 137150 2590
rect 137350 2520 137650 2590
rect 137850 2520 138150 2590
rect 138350 2520 138650 2590
rect 138850 2520 139150 2590
rect 139350 2520 139650 2590
rect 139850 2520 140000 2590
rect 136000 2480 140000 2520
rect 136000 2410 136150 2480
rect 136350 2410 136650 2480
rect 136850 2410 137150 2480
rect 137350 2410 137650 2480
rect 137850 2410 138150 2480
rect 138350 2410 138650 2480
rect 138850 2410 139150 2480
rect 139350 2410 139650 2480
rect 139850 2410 140000 2480
rect 136000 2400 140000 2410
rect 136000 2380 136120 2400
rect 136380 2380 136620 2400
rect 136880 2380 137120 2400
rect 137380 2380 137620 2400
rect 137880 2380 138120 2400
rect 138380 2380 138620 2400
rect 138880 2380 139120 2400
rect 139380 2380 139620 2400
rect 139880 2380 140000 2400
rect 136000 2350 136100 2380
rect 136000 2150 136020 2350
rect 136090 2150 136100 2350
rect 136000 2120 136100 2150
rect 136400 2350 136600 2380
rect 136400 2150 136410 2350
rect 136480 2150 136520 2350
rect 136590 2150 136600 2350
rect 136400 2120 136600 2150
rect 136900 2350 137100 2380
rect 136900 2150 136910 2350
rect 136980 2150 137020 2350
rect 137090 2150 137100 2350
rect 136900 2120 137100 2150
rect 137400 2350 137600 2380
rect 137400 2150 137410 2350
rect 137480 2150 137520 2350
rect 137590 2150 137600 2350
rect 137400 2120 137600 2150
rect 137900 2350 138100 2380
rect 137900 2150 137910 2350
rect 137980 2150 138020 2350
rect 138090 2150 138100 2350
rect 137900 2120 138100 2150
rect 138400 2350 138600 2380
rect 138400 2150 138410 2350
rect 138480 2150 138520 2350
rect 138590 2150 138600 2350
rect 138400 2120 138600 2150
rect 138900 2350 139100 2380
rect 138900 2150 138910 2350
rect 138980 2150 139020 2350
rect 139090 2150 139100 2350
rect 138900 2120 139100 2150
rect 139400 2350 139600 2380
rect 139400 2150 139410 2350
rect 139480 2150 139520 2350
rect 139590 2150 139600 2350
rect 139400 2120 139600 2150
rect 139900 2350 140000 2380
rect 139900 2150 139910 2350
rect 139980 2150 140000 2350
rect 139900 2120 140000 2150
rect 136000 2100 136120 2120
rect 136380 2100 136620 2120
rect 136880 2100 137120 2120
rect 137380 2100 137620 2120
rect 137880 2100 138120 2120
rect 138380 2100 138620 2120
rect 138880 2100 139120 2120
rect 139380 2100 139620 2120
rect 139880 2100 140000 2120
rect 136000 2090 140000 2100
rect 136000 2020 136150 2090
rect 136350 2020 136650 2090
rect 136850 2020 137150 2090
rect 137350 2020 137650 2090
rect 137850 2020 138150 2090
rect 138350 2020 138650 2090
rect 138850 2020 139150 2090
rect 139350 2020 139650 2090
rect 139850 2020 140000 2090
rect 136000 2000 140000 2020
rect 88000 1980 140000 2000
rect 88000 1910 136150 1980
rect 136350 1910 136650 1980
rect 136850 1910 137150 1980
rect 137350 1910 137650 1980
rect 137850 1910 138150 1980
rect 138350 1910 138650 1980
rect 138850 1910 139150 1980
rect 139350 1910 139650 1980
rect 139850 1910 140000 1980
rect 88000 1900 140000 1910
rect 88000 1880 88120 1900
rect 88380 1880 88620 1900
rect 88880 1880 89120 1900
rect 89380 1880 89620 1900
rect 89880 1880 90120 1900
rect 90380 1880 90620 1900
rect 90880 1880 91120 1900
rect 91380 1880 91620 1900
rect 91880 1880 92120 1900
rect 92380 1880 92620 1900
rect 92880 1880 93120 1900
rect 93380 1880 93620 1900
rect 93880 1880 94120 1900
rect 94380 1880 94620 1900
rect 94880 1880 95120 1900
rect 95380 1880 95620 1900
rect 95880 1880 96120 1900
rect 96380 1880 96620 1900
rect 96880 1880 97120 1900
rect 97380 1880 97620 1900
rect 97880 1880 98120 1900
rect 98380 1880 98620 1900
rect 98880 1880 99120 1900
rect 99380 1880 99620 1900
rect 99880 1880 100120 1900
rect 100380 1880 100620 1900
rect 100880 1880 101120 1900
rect 101380 1880 101620 1900
rect 101880 1880 102120 1900
rect 102380 1880 102620 1900
rect 102880 1880 103120 1900
rect 103380 1880 103620 1900
rect 103880 1880 104120 1900
rect 104380 1880 104620 1900
rect 104880 1880 105120 1900
rect 105380 1880 105620 1900
rect 105880 1880 106120 1900
rect 106380 1880 106620 1900
rect 106880 1880 107120 1900
rect 107380 1880 107620 1900
rect 107880 1880 108120 1900
rect 108380 1880 108620 1900
rect 108880 1880 109120 1900
rect 109380 1880 109620 1900
rect 109880 1880 110120 1900
rect 110380 1880 110620 1900
rect 110880 1880 111120 1900
rect 111380 1880 111620 1900
rect 111880 1880 112120 1900
rect 112380 1880 112620 1900
rect 112880 1880 113120 1900
rect 113380 1880 113620 1900
rect 113880 1880 114120 1900
rect 114380 1880 114620 1900
rect 114880 1880 115120 1900
rect 115380 1880 115620 1900
rect 115880 1880 116120 1900
rect 116380 1880 116620 1900
rect 116880 1880 117120 1900
rect 117380 1880 117620 1900
rect 117880 1880 118120 1900
rect 118380 1880 118620 1900
rect 118880 1880 119120 1900
rect 119380 1880 119620 1900
rect 119880 1880 120120 1900
rect 120380 1880 120620 1900
rect 120880 1880 121120 1900
rect 121380 1880 121620 1900
rect 121880 1880 122120 1900
rect 122380 1880 122620 1900
rect 122880 1880 123120 1900
rect 123380 1880 123620 1900
rect 123880 1880 124120 1900
rect 124380 1880 124620 1900
rect 124880 1880 125120 1900
rect 125380 1880 125620 1900
rect 125880 1880 126120 1900
rect 126380 1880 126620 1900
rect 126880 1880 127120 1900
rect 127380 1880 127620 1900
rect 127880 1880 128120 1900
rect 128380 1880 128620 1900
rect 128880 1880 129120 1900
rect 129380 1880 129620 1900
rect 129880 1880 130120 1900
rect 130380 1880 130620 1900
rect 130880 1880 131120 1900
rect 131380 1880 131620 1900
rect 131880 1880 132120 1900
rect 132380 1880 132620 1900
rect 132880 1880 133120 1900
rect 133380 1880 133620 1900
rect 133880 1880 134120 1900
rect 134380 1880 134620 1900
rect 134880 1880 135120 1900
rect 135380 1880 135620 1900
rect 135880 1880 136120 1900
rect 136380 1880 136620 1900
rect 136880 1880 137120 1900
rect 137380 1880 137620 1900
rect 137880 1880 138120 1900
rect 138380 1880 138620 1900
rect 138880 1880 139120 1900
rect 139380 1880 139620 1900
rect 139880 1880 140000 1900
rect 88000 1620 88100 1880
rect 88400 1620 88600 1880
rect 88900 1620 89100 1880
rect 89400 1620 89600 1880
rect 89900 1620 90100 1880
rect 90400 1620 90600 1880
rect 90900 1620 91100 1880
rect 91400 1620 91600 1880
rect 91900 1620 92100 1880
rect 92400 1620 92600 1880
rect 92900 1620 93100 1880
rect 93400 1620 93600 1880
rect 93900 1620 94100 1880
rect 94400 1620 94600 1880
rect 94900 1620 95100 1880
rect 95400 1620 95600 1880
rect 95900 1620 96100 1880
rect 96400 1620 96600 1880
rect 96900 1620 97100 1880
rect 97400 1620 97600 1880
rect 97900 1620 98100 1880
rect 98400 1620 98600 1880
rect 98900 1620 99100 1880
rect 99400 1620 99600 1880
rect 99900 1620 100100 1880
rect 100400 1620 100600 1880
rect 100900 1620 101100 1880
rect 101400 1620 101600 1880
rect 101900 1620 102100 1880
rect 102400 1620 102600 1880
rect 102900 1620 103100 1880
rect 103400 1620 103600 1880
rect 103900 1620 104100 1880
rect 104400 1620 104600 1880
rect 104900 1620 105100 1880
rect 105400 1620 105600 1880
rect 105900 1620 106100 1880
rect 106400 1620 106600 1880
rect 106900 1620 107100 1880
rect 107400 1620 107600 1880
rect 107900 1620 108100 1880
rect 108400 1620 108600 1880
rect 108900 1620 109100 1880
rect 109400 1620 109600 1880
rect 109900 1620 110100 1880
rect 110400 1620 110600 1880
rect 110900 1620 111100 1880
rect 111400 1620 111600 1880
rect 111900 1620 112100 1880
rect 112400 1620 112600 1880
rect 112900 1620 113100 1880
rect 113400 1620 113600 1880
rect 113900 1620 114100 1880
rect 114400 1620 114600 1880
rect 114900 1620 115100 1880
rect 115400 1620 115600 1880
rect 115900 1620 116100 1880
rect 116400 1620 116600 1880
rect 116900 1620 117100 1880
rect 117400 1620 117600 1880
rect 117900 1620 118100 1880
rect 118400 1620 118600 1880
rect 118900 1620 119100 1880
rect 119400 1620 119600 1880
rect 119900 1620 120100 1880
rect 120400 1620 120600 1880
rect 120900 1620 121100 1880
rect 121400 1620 121600 1880
rect 121900 1620 122100 1880
rect 122400 1620 122600 1880
rect 122900 1620 123100 1880
rect 123400 1620 123600 1880
rect 123900 1620 124100 1880
rect 124400 1620 124600 1880
rect 124900 1620 125100 1880
rect 125400 1620 125600 1880
rect 125900 1620 126100 1880
rect 126400 1620 126600 1880
rect 126900 1620 127100 1880
rect 127400 1620 127600 1880
rect 127900 1620 128100 1880
rect 128400 1620 128600 1880
rect 128900 1620 129100 1880
rect 129400 1620 129600 1880
rect 129900 1620 130100 1880
rect 130400 1620 130600 1880
rect 130900 1620 131100 1880
rect 131400 1620 131600 1880
rect 131900 1620 132100 1880
rect 132400 1620 132600 1880
rect 132900 1620 133100 1880
rect 133400 1620 133600 1880
rect 133900 1620 134100 1880
rect 134400 1620 134600 1880
rect 134900 1620 135100 1880
rect 135400 1620 135600 1880
rect 135900 1850 136100 1880
rect 135900 1650 136020 1850
rect 136090 1650 136100 1850
rect 135900 1620 136100 1650
rect 136400 1850 136600 1880
rect 136400 1650 136410 1850
rect 136480 1650 136520 1850
rect 136590 1650 136600 1850
rect 136400 1620 136600 1650
rect 136900 1850 137100 1880
rect 136900 1650 136910 1850
rect 136980 1650 137020 1850
rect 137090 1650 137100 1850
rect 136900 1620 137100 1650
rect 137400 1850 137600 1880
rect 137400 1650 137410 1850
rect 137480 1650 137520 1850
rect 137590 1650 137600 1850
rect 137400 1620 137600 1650
rect 137900 1850 138100 1880
rect 137900 1650 137910 1850
rect 137980 1650 138020 1850
rect 138090 1650 138100 1850
rect 137900 1620 138100 1650
rect 138400 1850 138600 1880
rect 138400 1650 138410 1850
rect 138480 1650 138520 1850
rect 138590 1650 138600 1850
rect 138400 1620 138600 1650
rect 138900 1850 139100 1880
rect 138900 1650 138910 1850
rect 138980 1650 139020 1850
rect 139090 1650 139100 1850
rect 138900 1620 139100 1650
rect 139400 1850 139600 1880
rect 139400 1650 139410 1850
rect 139480 1650 139520 1850
rect 139590 1650 139600 1850
rect 139400 1620 139600 1650
rect 139900 1850 140000 1880
rect 139900 1650 139910 1850
rect 139980 1650 140000 1850
rect 139900 1620 140000 1650
rect 88000 1600 88120 1620
rect 88380 1600 88620 1620
rect 88880 1600 89120 1620
rect 89380 1600 89620 1620
rect 89880 1600 90120 1620
rect 90380 1600 90620 1620
rect 90880 1600 91120 1620
rect 91380 1600 91620 1620
rect 91880 1600 92120 1620
rect 92380 1600 92620 1620
rect 92880 1600 93120 1620
rect 93380 1600 93620 1620
rect 93880 1600 94120 1620
rect 94380 1600 94620 1620
rect 94880 1600 95120 1620
rect 95380 1600 95620 1620
rect 95880 1600 96120 1620
rect 96380 1600 96620 1620
rect 96880 1600 97120 1620
rect 97380 1600 97620 1620
rect 97880 1600 98120 1620
rect 98380 1600 98620 1620
rect 98880 1600 99120 1620
rect 99380 1600 99620 1620
rect 99880 1600 100120 1620
rect 100380 1600 100620 1620
rect 100880 1600 101120 1620
rect 101380 1600 101620 1620
rect 101880 1600 102120 1620
rect 102380 1600 102620 1620
rect 102880 1600 103120 1620
rect 103380 1600 103620 1620
rect 103880 1600 104120 1620
rect 104380 1600 104620 1620
rect 104880 1600 105120 1620
rect 105380 1600 105620 1620
rect 105880 1600 106120 1620
rect 106380 1600 106620 1620
rect 106880 1600 107120 1620
rect 107380 1600 107620 1620
rect 107880 1600 108120 1620
rect 108380 1600 108620 1620
rect 108880 1600 109120 1620
rect 109380 1600 109620 1620
rect 109880 1600 110120 1620
rect 110380 1600 110620 1620
rect 110880 1600 111120 1620
rect 111380 1600 111620 1620
rect 111880 1600 112120 1620
rect 112380 1600 112620 1620
rect 112880 1600 113120 1620
rect 113380 1600 113620 1620
rect 113880 1600 114120 1620
rect 114380 1600 114620 1620
rect 114880 1600 115120 1620
rect 115380 1600 115620 1620
rect 115880 1600 116120 1620
rect 116380 1600 116620 1620
rect 116880 1600 117120 1620
rect 117380 1600 117620 1620
rect 117880 1600 118120 1620
rect 118380 1600 118620 1620
rect 118880 1600 119120 1620
rect 119380 1600 119620 1620
rect 119880 1600 120120 1620
rect 120380 1600 120620 1620
rect 120880 1600 121120 1620
rect 121380 1600 121620 1620
rect 121880 1600 122120 1620
rect 122380 1600 122620 1620
rect 122880 1600 123120 1620
rect 123380 1600 123620 1620
rect 123880 1600 124120 1620
rect 124380 1600 124620 1620
rect 124880 1600 125120 1620
rect 125380 1600 125620 1620
rect 125880 1600 126120 1620
rect 126380 1600 126620 1620
rect 126880 1600 127120 1620
rect 127380 1600 127620 1620
rect 127880 1600 128120 1620
rect 128380 1600 128620 1620
rect 128880 1600 129120 1620
rect 129380 1600 129620 1620
rect 129880 1600 130120 1620
rect 130380 1600 130620 1620
rect 130880 1600 131120 1620
rect 131380 1600 131620 1620
rect 131880 1600 132120 1620
rect 132380 1600 132620 1620
rect 132880 1600 133120 1620
rect 133380 1600 133620 1620
rect 133880 1600 134120 1620
rect 134380 1600 134620 1620
rect 134880 1600 135120 1620
rect 135380 1600 135620 1620
rect 135880 1600 136120 1620
rect 136380 1600 136620 1620
rect 136880 1600 137120 1620
rect 137380 1600 137620 1620
rect 137880 1600 138120 1620
rect 138380 1600 138620 1620
rect 138880 1600 139120 1620
rect 139380 1600 139620 1620
rect 139880 1600 140000 1620
rect 88000 1590 140000 1600
rect 88000 1520 136150 1590
rect 136350 1520 136650 1590
rect 136850 1520 137150 1590
rect 137350 1520 137650 1590
rect 137850 1520 138150 1590
rect 138350 1520 138650 1590
rect 138850 1520 139150 1590
rect 139350 1520 139650 1590
rect 139850 1520 140000 1590
rect 88000 1480 140000 1520
rect 88000 1410 136150 1480
rect 136350 1410 136650 1480
rect 136850 1410 137150 1480
rect 137350 1410 137650 1480
rect 137850 1410 138150 1480
rect 138350 1410 138650 1480
rect 138850 1410 139150 1480
rect 139350 1410 139650 1480
rect 139850 1410 140000 1480
rect 88000 1400 140000 1410
rect 88000 1380 88120 1400
rect 88380 1380 88620 1400
rect 88880 1380 89120 1400
rect 89380 1380 89620 1400
rect 89880 1380 90120 1400
rect 90380 1380 90620 1400
rect 90880 1380 91120 1400
rect 91380 1380 91620 1400
rect 91880 1380 92120 1400
rect 92380 1380 92620 1400
rect 92880 1380 93120 1400
rect 93380 1380 93620 1400
rect 93880 1380 94120 1400
rect 94380 1380 94620 1400
rect 94880 1380 95120 1400
rect 95380 1380 95620 1400
rect 95880 1380 96120 1400
rect 96380 1380 96620 1400
rect 96880 1380 97120 1400
rect 97380 1380 97620 1400
rect 97880 1380 98120 1400
rect 98380 1380 98620 1400
rect 98880 1380 99120 1400
rect 99380 1380 99620 1400
rect 99880 1380 100120 1400
rect 100380 1380 100620 1400
rect 100880 1380 101120 1400
rect 101380 1380 101620 1400
rect 101880 1380 102120 1400
rect 102380 1380 102620 1400
rect 102880 1380 103120 1400
rect 103380 1380 103620 1400
rect 103880 1380 104120 1400
rect 104380 1380 104620 1400
rect 104880 1380 105120 1400
rect 105380 1380 105620 1400
rect 105880 1380 106120 1400
rect 106380 1380 106620 1400
rect 106880 1380 107120 1400
rect 107380 1380 107620 1400
rect 107880 1380 108120 1400
rect 108380 1380 108620 1400
rect 108880 1380 109120 1400
rect 109380 1380 109620 1400
rect 109880 1380 110120 1400
rect 110380 1380 110620 1400
rect 110880 1380 111120 1400
rect 111380 1380 111620 1400
rect 111880 1380 112120 1400
rect 112380 1380 112620 1400
rect 112880 1380 113120 1400
rect 113380 1380 113620 1400
rect 113880 1380 114120 1400
rect 114380 1380 114620 1400
rect 114880 1380 115120 1400
rect 115380 1380 115620 1400
rect 115880 1380 116120 1400
rect 116380 1380 116620 1400
rect 116880 1380 117120 1400
rect 117380 1380 117620 1400
rect 117880 1380 118120 1400
rect 118380 1380 118620 1400
rect 118880 1380 119120 1400
rect 119380 1380 119620 1400
rect 119880 1380 120120 1400
rect 120380 1380 120620 1400
rect 120880 1380 121120 1400
rect 121380 1380 121620 1400
rect 121880 1380 122120 1400
rect 122380 1380 122620 1400
rect 122880 1380 123120 1400
rect 123380 1380 123620 1400
rect 123880 1380 124120 1400
rect 124380 1380 124620 1400
rect 124880 1380 125120 1400
rect 125380 1380 125620 1400
rect 125880 1380 126120 1400
rect 126380 1380 126620 1400
rect 126880 1380 127120 1400
rect 127380 1380 127620 1400
rect 127880 1380 128120 1400
rect 128380 1380 128620 1400
rect 128880 1380 129120 1400
rect 129380 1380 129620 1400
rect 129880 1380 130120 1400
rect 130380 1380 130620 1400
rect 130880 1380 131120 1400
rect 131380 1380 131620 1400
rect 131880 1380 132120 1400
rect 132380 1380 132620 1400
rect 132880 1380 133120 1400
rect 133380 1380 133620 1400
rect 133880 1380 134120 1400
rect 134380 1380 134620 1400
rect 134880 1380 135120 1400
rect 135380 1380 135620 1400
rect 135880 1380 136120 1400
rect 136380 1380 136620 1400
rect 136880 1380 137120 1400
rect 137380 1380 137620 1400
rect 137880 1380 138120 1400
rect 138380 1380 138620 1400
rect 138880 1380 139120 1400
rect 139380 1380 139620 1400
rect 139880 1380 140000 1400
rect 88000 1120 88100 1380
rect 88400 1120 88600 1380
rect 88900 1120 89100 1380
rect 89400 1120 89600 1380
rect 89900 1120 90100 1380
rect 90400 1120 90600 1380
rect 90900 1120 91100 1380
rect 91400 1120 91600 1380
rect 91900 1120 92100 1380
rect 92400 1120 92600 1380
rect 92900 1120 93100 1380
rect 93400 1120 93600 1380
rect 93900 1120 94100 1380
rect 94400 1120 94600 1380
rect 94900 1120 95100 1380
rect 95400 1120 95600 1380
rect 95900 1120 96100 1380
rect 96400 1120 96600 1380
rect 96900 1120 97100 1380
rect 97400 1120 97600 1380
rect 97900 1120 98100 1380
rect 98400 1120 98600 1380
rect 98900 1120 99100 1380
rect 99400 1120 99600 1380
rect 99900 1120 100100 1380
rect 100400 1120 100600 1380
rect 100900 1120 101100 1380
rect 101400 1120 101600 1380
rect 101900 1120 102100 1380
rect 102400 1120 102600 1380
rect 102900 1120 103100 1380
rect 103400 1120 103600 1380
rect 103900 1120 104100 1380
rect 104400 1120 104600 1380
rect 104900 1120 105100 1380
rect 105400 1120 105600 1380
rect 105900 1120 106100 1380
rect 106400 1120 106600 1380
rect 106900 1120 107100 1380
rect 107400 1120 107600 1380
rect 107900 1120 108100 1380
rect 108400 1120 108600 1380
rect 108900 1120 109100 1380
rect 109400 1120 109600 1380
rect 109900 1120 110100 1380
rect 110400 1120 110600 1380
rect 110900 1120 111100 1380
rect 111400 1120 111600 1380
rect 111900 1120 112100 1380
rect 112400 1120 112600 1380
rect 112900 1120 113100 1380
rect 113400 1120 113600 1380
rect 113900 1120 114100 1380
rect 114400 1120 114600 1380
rect 114900 1120 115100 1380
rect 115400 1120 115600 1380
rect 115900 1120 116100 1380
rect 116400 1120 116600 1380
rect 116900 1120 117100 1380
rect 117400 1120 117600 1380
rect 117900 1120 118100 1380
rect 118400 1120 118600 1380
rect 118900 1120 119100 1380
rect 119400 1120 119600 1380
rect 119900 1120 120100 1380
rect 120400 1120 120600 1380
rect 120900 1120 121100 1380
rect 121400 1120 121600 1380
rect 121900 1120 122100 1380
rect 122400 1120 122600 1380
rect 122900 1120 123100 1380
rect 123400 1120 123600 1380
rect 123900 1120 124100 1380
rect 124400 1120 124600 1380
rect 124900 1120 125100 1380
rect 125400 1120 125600 1380
rect 125900 1120 126100 1380
rect 126400 1120 126600 1380
rect 126900 1120 127100 1380
rect 127400 1120 127600 1380
rect 127900 1120 128100 1380
rect 128400 1120 128600 1380
rect 128900 1120 129100 1380
rect 129400 1120 129600 1380
rect 129900 1120 130100 1380
rect 130400 1120 130600 1380
rect 130900 1120 131100 1380
rect 131400 1120 131600 1380
rect 131900 1120 132100 1380
rect 132400 1120 132600 1380
rect 132900 1120 133100 1380
rect 133400 1120 133600 1380
rect 133900 1120 134100 1380
rect 134400 1120 134600 1380
rect 134900 1120 135100 1380
rect 135400 1120 135600 1380
rect 135900 1350 136100 1380
rect 135900 1150 136020 1350
rect 136090 1150 136100 1350
rect 135900 1120 136100 1150
rect 136400 1350 136600 1380
rect 136400 1150 136410 1350
rect 136480 1150 136520 1350
rect 136590 1150 136600 1350
rect 136400 1120 136600 1150
rect 136900 1350 137100 1380
rect 136900 1150 136910 1350
rect 136980 1150 137020 1350
rect 137090 1150 137100 1350
rect 136900 1120 137100 1150
rect 137400 1350 137600 1380
rect 137400 1150 137410 1350
rect 137480 1150 137520 1350
rect 137590 1150 137600 1350
rect 137400 1120 137600 1150
rect 137900 1350 138100 1380
rect 137900 1150 137910 1350
rect 137980 1150 138020 1350
rect 138090 1150 138100 1350
rect 137900 1120 138100 1150
rect 138400 1350 138600 1380
rect 138400 1150 138410 1350
rect 138480 1150 138520 1350
rect 138590 1150 138600 1350
rect 138400 1120 138600 1150
rect 138900 1350 139100 1380
rect 138900 1150 138910 1350
rect 138980 1150 139020 1350
rect 139090 1150 139100 1350
rect 138900 1120 139100 1150
rect 139400 1350 139600 1380
rect 139400 1150 139410 1350
rect 139480 1150 139520 1350
rect 139590 1150 139600 1350
rect 139400 1120 139600 1150
rect 139900 1350 140000 1380
rect 139900 1150 139910 1350
rect 139980 1150 140000 1350
rect 139900 1120 140000 1150
rect 88000 1100 88120 1120
rect 88380 1100 88620 1120
rect 88880 1100 89120 1120
rect 89380 1100 89620 1120
rect 89880 1100 90120 1120
rect 90380 1100 90620 1120
rect 90880 1100 91120 1120
rect 91380 1100 91620 1120
rect 91880 1100 92120 1120
rect 92380 1100 92620 1120
rect 92880 1100 93120 1120
rect 93380 1100 93620 1120
rect 93880 1100 94120 1120
rect 94380 1100 94620 1120
rect 94880 1100 95120 1120
rect 95380 1100 95620 1120
rect 95880 1100 96120 1120
rect 96380 1100 96620 1120
rect 96880 1100 97120 1120
rect 97380 1100 97620 1120
rect 97880 1100 98120 1120
rect 98380 1100 98620 1120
rect 98880 1100 99120 1120
rect 99380 1100 99620 1120
rect 99880 1100 100120 1120
rect 100380 1100 100620 1120
rect 100880 1100 101120 1120
rect 101380 1100 101620 1120
rect 101880 1100 102120 1120
rect 102380 1100 102620 1120
rect 102880 1100 103120 1120
rect 103380 1100 103620 1120
rect 103880 1100 104120 1120
rect 104380 1100 104620 1120
rect 104880 1100 105120 1120
rect 105380 1100 105620 1120
rect 105880 1100 106120 1120
rect 106380 1100 106620 1120
rect 106880 1100 107120 1120
rect 107380 1100 107620 1120
rect 107880 1100 108120 1120
rect 108380 1100 108620 1120
rect 108880 1100 109120 1120
rect 109380 1100 109620 1120
rect 109880 1100 110120 1120
rect 110380 1100 110620 1120
rect 110880 1100 111120 1120
rect 111380 1100 111620 1120
rect 111880 1100 112120 1120
rect 112380 1100 112620 1120
rect 112880 1100 113120 1120
rect 113380 1100 113620 1120
rect 113880 1100 114120 1120
rect 114380 1100 114620 1120
rect 114880 1100 115120 1120
rect 115380 1100 115620 1120
rect 115880 1100 116120 1120
rect 116380 1100 116620 1120
rect 116880 1100 117120 1120
rect 117380 1100 117620 1120
rect 117880 1100 118120 1120
rect 118380 1100 118620 1120
rect 118880 1100 119120 1120
rect 119380 1100 119620 1120
rect 119880 1100 120120 1120
rect 120380 1100 120620 1120
rect 120880 1100 121120 1120
rect 121380 1100 121620 1120
rect 121880 1100 122120 1120
rect 122380 1100 122620 1120
rect 122880 1100 123120 1120
rect 123380 1100 123620 1120
rect 123880 1100 124120 1120
rect 124380 1100 124620 1120
rect 124880 1100 125120 1120
rect 125380 1100 125620 1120
rect 125880 1100 126120 1120
rect 126380 1100 126620 1120
rect 126880 1100 127120 1120
rect 127380 1100 127620 1120
rect 127880 1100 128120 1120
rect 128380 1100 128620 1120
rect 128880 1100 129120 1120
rect 129380 1100 129620 1120
rect 129880 1100 130120 1120
rect 130380 1100 130620 1120
rect 130880 1100 131120 1120
rect 131380 1100 131620 1120
rect 131880 1100 132120 1120
rect 132380 1100 132620 1120
rect 132880 1100 133120 1120
rect 133380 1100 133620 1120
rect 133880 1100 134120 1120
rect 134380 1100 134620 1120
rect 134880 1100 135120 1120
rect 135380 1100 135620 1120
rect 135880 1100 136120 1120
rect 136380 1100 136620 1120
rect 136880 1100 137120 1120
rect 137380 1100 137620 1120
rect 137880 1100 138120 1120
rect 138380 1100 138620 1120
rect 138880 1100 139120 1120
rect 139380 1100 139620 1120
rect 139880 1100 140000 1120
rect 88000 1090 140000 1100
rect 88000 1020 136150 1090
rect 136350 1020 136650 1090
rect 136850 1020 137150 1090
rect 137350 1020 137650 1090
rect 137850 1020 138150 1090
rect 138350 1020 138650 1090
rect 138850 1020 139150 1090
rect 139350 1020 139650 1090
rect 139850 1020 140000 1090
rect 88000 980 140000 1020
rect 88000 910 136150 980
rect 136350 910 136650 980
rect 136850 910 137150 980
rect 137350 910 137650 980
rect 137850 910 138150 980
rect 138350 910 138650 980
rect 138850 910 139150 980
rect 139350 910 139650 980
rect 139850 910 140000 980
rect 88000 900 140000 910
rect 88000 880 88120 900
rect 88380 880 88620 900
rect 88880 880 89120 900
rect 89380 880 89620 900
rect 89880 880 90120 900
rect 90380 880 90620 900
rect 90880 880 91120 900
rect 91380 880 91620 900
rect 91880 880 92120 900
rect 92380 880 92620 900
rect 92880 880 93120 900
rect 93380 880 93620 900
rect 93880 880 94120 900
rect 94380 880 94620 900
rect 94880 880 95120 900
rect 95380 880 95620 900
rect 95880 880 96120 900
rect 96380 880 96620 900
rect 96880 880 97120 900
rect 97380 880 97620 900
rect 97880 880 98120 900
rect 98380 880 98620 900
rect 98880 880 99120 900
rect 99380 880 99620 900
rect 99880 880 100120 900
rect 100380 880 100620 900
rect 100880 880 101120 900
rect 101380 880 101620 900
rect 101880 880 102120 900
rect 102380 880 102620 900
rect 102880 880 103120 900
rect 103380 880 103620 900
rect 103880 880 104120 900
rect 104380 880 104620 900
rect 104880 880 105120 900
rect 105380 880 105620 900
rect 105880 880 106120 900
rect 106380 880 106620 900
rect 106880 880 107120 900
rect 107380 880 107620 900
rect 107880 880 108120 900
rect 108380 880 108620 900
rect 108880 880 109120 900
rect 109380 880 109620 900
rect 109880 880 110120 900
rect 110380 880 110620 900
rect 110880 880 111120 900
rect 111380 880 111620 900
rect 111880 880 112120 900
rect 112380 880 112620 900
rect 112880 880 113120 900
rect 113380 880 113620 900
rect 113880 880 114120 900
rect 114380 880 114620 900
rect 114880 880 115120 900
rect 115380 880 115620 900
rect 115880 880 116120 900
rect 116380 880 116620 900
rect 116880 880 117120 900
rect 117380 880 117620 900
rect 117880 880 118120 900
rect 118380 880 118620 900
rect 118880 880 119120 900
rect 119380 880 119620 900
rect 119880 880 120120 900
rect 120380 880 120620 900
rect 120880 880 121120 900
rect 121380 880 121620 900
rect 121880 880 122120 900
rect 122380 880 122620 900
rect 122880 880 123120 900
rect 123380 880 123620 900
rect 123880 880 124120 900
rect 124380 880 124620 900
rect 124880 880 125120 900
rect 125380 880 125620 900
rect 125880 880 126120 900
rect 126380 880 126620 900
rect 126880 880 127120 900
rect 127380 880 127620 900
rect 127880 880 128120 900
rect 128380 880 128620 900
rect 128880 880 129120 900
rect 129380 880 129620 900
rect 129880 880 130120 900
rect 130380 880 130620 900
rect 130880 880 131120 900
rect 131380 880 131620 900
rect 131880 880 132120 900
rect 132380 880 132620 900
rect 132880 880 133120 900
rect 133380 880 133620 900
rect 133880 880 134120 900
rect 134380 880 134620 900
rect 134880 880 135120 900
rect 135380 880 135620 900
rect 135880 880 136120 900
rect 136380 880 136620 900
rect 136880 880 137120 900
rect 137380 880 137620 900
rect 137880 880 138120 900
rect 138380 880 138620 900
rect 138880 880 139120 900
rect 139380 880 139620 900
rect 139880 880 140000 900
rect 88000 620 88100 880
rect 88400 620 88600 880
rect 88900 620 89100 880
rect 89400 620 89600 880
rect 89900 620 90100 880
rect 90400 620 90600 880
rect 90900 620 91100 880
rect 91400 620 91600 880
rect 91900 620 92100 880
rect 92400 620 92600 880
rect 92900 620 93100 880
rect 93400 620 93600 880
rect 93900 620 94100 880
rect 94400 620 94600 880
rect 94900 620 95100 880
rect 95400 620 95600 880
rect 95900 620 96100 880
rect 96400 620 96600 880
rect 96900 620 97100 880
rect 97400 620 97600 880
rect 97900 620 98100 880
rect 98400 620 98600 880
rect 98900 620 99100 880
rect 99400 620 99600 880
rect 99900 620 100100 880
rect 100400 620 100600 880
rect 100900 620 101100 880
rect 101400 620 101600 880
rect 101900 620 102100 880
rect 102400 620 102600 880
rect 102900 620 103100 880
rect 103400 620 103600 880
rect 103900 620 104100 880
rect 104400 620 104600 880
rect 104900 620 105100 880
rect 105400 620 105600 880
rect 105900 620 106100 880
rect 106400 620 106600 880
rect 106900 620 107100 880
rect 107400 620 107600 880
rect 107900 620 108100 880
rect 108400 620 108600 880
rect 108900 620 109100 880
rect 109400 620 109600 880
rect 109900 620 110100 880
rect 110400 620 110600 880
rect 110900 620 111100 880
rect 111400 620 111600 880
rect 111900 620 112100 880
rect 112400 620 112600 880
rect 112900 620 113100 880
rect 113400 620 113600 880
rect 113900 620 114100 880
rect 114400 620 114600 880
rect 114900 620 115100 880
rect 115400 620 115600 880
rect 115900 620 116100 880
rect 116400 620 116600 880
rect 116900 620 117100 880
rect 117400 620 117600 880
rect 117900 620 118100 880
rect 118400 620 118600 880
rect 118900 620 119100 880
rect 119400 620 119600 880
rect 119900 620 120100 880
rect 120400 620 120600 880
rect 120900 620 121100 880
rect 121400 620 121600 880
rect 121900 620 122100 880
rect 122400 620 122600 880
rect 122900 620 123100 880
rect 123400 620 123600 880
rect 123900 620 124100 880
rect 124400 620 124600 880
rect 124900 620 125100 880
rect 125400 620 125600 880
rect 125900 620 126100 880
rect 126400 620 126600 880
rect 126900 620 127100 880
rect 127400 620 127600 880
rect 127900 620 128100 880
rect 128400 620 128600 880
rect 128900 620 129100 880
rect 129400 620 129600 880
rect 129900 620 130100 880
rect 130400 620 130600 880
rect 130900 620 131100 880
rect 131400 620 131600 880
rect 131900 620 132100 880
rect 132400 620 132600 880
rect 132900 620 133100 880
rect 133400 620 133600 880
rect 133900 620 134100 880
rect 134400 620 134600 880
rect 134900 620 135100 880
rect 135400 620 135600 880
rect 135900 850 136100 880
rect 135900 650 136020 850
rect 136090 650 136100 850
rect 135900 620 136100 650
rect 136400 850 136600 880
rect 136400 650 136410 850
rect 136480 650 136520 850
rect 136590 650 136600 850
rect 136400 620 136600 650
rect 136900 850 137100 880
rect 136900 650 136910 850
rect 136980 650 137020 850
rect 137090 650 137100 850
rect 136900 620 137100 650
rect 137400 850 137600 880
rect 137400 650 137410 850
rect 137480 650 137520 850
rect 137590 650 137600 850
rect 137400 620 137600 650
rect 137900 850 138100 880
rect 137900 650 137910 850
rect 137980 650 138020 850
rect 138090 650 138100 850
rect 137900 620 138100 650
rect 138400 850 138600 880
rect 138400 650 138410 850
rect 138480 650 138520 850
rect 138590 650 138600 850
rect 138400 620 138600 650
rect 138900 850 139100 880
rect 138900 650 138910 850
rect 138980 650 139020 850
rect 139090 650 139100 850
rect 138900 620 139100 650
rect 139400 850 139600 880
rect 139400 650 139410 850
rect 139480 650 139520 850
rect 139590 650 139600 850
rect 139400 620 139600 650
rect 139900 850 140000 880
rect 139900 650 139910 850
rect 139980 650 140000 850
rect 139900 620 140000 650
rect 88000 600 88120 620
rect 88380 600 88620 620
rect 88880 600 89120 620
rect 89380 600 89620 620
rect 89880 600 90120 620
rect 90380 600 90620 620
rect 90880 600 91120 620
rect 91380 600 91620 620
rect 91880 600 92120 620
rect 92380 600 92620 620
rect 92880 600 93120 620
rect 93380 600 93620 620
rect 93880 600 94120 620
rect 94380 600 94620 620
rect 94880 600 95120 620
rect 95380 600 95620 620
rect 95880 600 96120 620
rect 96380 600 96620 620
rect 96880 600 97120 620
rect 97380 600 97620 620
rect 97880 600 98120 620
rect 98380 600 98620 620
rect 98880 600 99120 620
rect 99380 600 99620 620
rect 99880 600 100120 620
rect 100380 600 100620 620
rect 100880 600 101120 620
rect 101380 600 101620 620
rect 101880 600 102120 620
rect 102380 600 102620 620
rect 102880 600 103120 620
rect 103380 600 103620 620
rect 103880 600 104120 620
rect 104380 600 104620 620
rect 104880 600 105120 620
rect 105380 600 105620 620
rect 105880 600 106120 620
rect 106380 600 106620 620
rect 106880 600 107120 620
rect 107380 600 107620 620
rect 107880 600 108120 620
rect 108380 600 108620 620
rect 108880 600 109120 620
rect 109380 600 109620 620
rect 109880 600 110120 620
rect 110380 600 110620 620
rect 110880 600 111120 620
rect 111380 600 111620 620
rect 111880 600 112120 620
rect 112380 600 112620 620
rect 112880 600 113120 620
rect 113380 600 113620 620
rect 113880 600 114120 620
rect 114380 600 114620 620
rect 114880 600 115120 620
rect 115380 600 115620 620
rect 115880 600 116120 620
rect 116380 600 116620 620
rect 116880 600 117120 620
rect 117380 600 117620 620
rect 117880 600 118120 620
rect 118380 600 118620 620
rect 118880 600 119120 620
rect 119380 600 119620 620
rect 119880 600 120120 620
rect 120380 600 120620 620
rect 120880 600 121120 620
rect 121380 600 121620 620
rect 121880 600 122120 620
rect 122380 600 122620 620
rect 122880 600 123120 620
rect 123380 600 123620 620
rect 123880 600 124120 620
rect 124380 600 124620 620
rect 124880 600 125120 620
rect 125380 600 125620 620
rect 125880 600 126120 620
rect 126380 600 126620 620
rect 126880 600 127120 620
rect 127380 600 127620 620
rect 127880 600 128120 620
rect 128380 600 128620 620
rect 128880 600 129120 620
rect 129380 600 129620 620
rect 129880 600 130120 620
rect 130380 600 130620 620
rect 130880 600 131120 620
rect 131380 600 131620 620
rect 131880 600 132120 620
rect 132380 600 132620 620
rect 132880 600 133120 620
rect 133380 600 133620 620
rect 133880 600 134120 620
rect 134380 600 134620 620
rect 134880 600 135120 620
rect 135380 600 135620 620
rect 135880 600 136120 620
rect 136380 600 136620 620
rect 136880 600 137120 620
rect 137380 600 137620 620
rect 137880 600 138120 620
rect 138380 600 138620 620
rect 138880 600 139120 620
rect 139380 600 139620 620
rect 139880 600 140000 620
rect 88000 590 140000 600
rect 88000 520 136150 590
rect 136350 520 136650 590
rect 136850 520 137150 590
rect 137350 520 137650 590
rect 137850 520 138150 590
rect 138350 520 138650 590
rect 138850 520 139150 590
rect 139350 520 139650 590
rect 139850 520 140000 590
rect 88000 480 140000 520
rect 88000 410 136150 480
rect 136350 410 136650 480
rect 136850 410 137150 480
rect 137350 410 137650 480
rect 137850 410 138150 480
rect 138350 410 138650 480
rect 138850 410 139150 480
rect 139350 410 139650 480
rect 139850 410 140000 480
rect 88000 400 140000 410
rect 88000 380 88120 400
rect 88380 380 88620 400
rect 88880 380 89120 400
rect 89380 380 89620 400
rect 89880 380 90120 400
rect 90380 380 90620 400
rect 90880 380 91120 400
rect 91380 380 91620 400
rect 91880 380 92120 400
rect 92380 380 92620 400
rect 92880 380 93120 400
rect 93380 380 93620 400
rect 93880 380 94120 400
rect 94380 380 94620 400
rect 94880 380 95120 400
rect 95380 380 95620 400
rect 95880 380 96120 400
rect 96380 380 96620 400
rect 96880 380 97120 400
rect 97380 380 97620 400
rect 97880 380 98120 400
rect 98380 380 98620 400
rect 98880 380 99120 400
rect 99380 380 99620 400
rect 99880 380 100120 400
rect 100380 380 100620 400
rect 100880 380 101120 400
rect 101380 380 101620 400
rect 101880 380 102120 400
rect 102380 380 102620 400
rect 102880 380 103120 400
rect 103380 380 103620 400
rect 103880 380 104120 400
rect 104380 380 104620 400
rect 104880 380 105120 400
rect 105380 380 105620 400
rect 105880 380 106120 400
rect 106380 380 106620 400
rect 106880 380 107120 400
rect 107380 380 107620 400
rect 107880 380 108120 400
rect 108380 380 108620 400
rect 108880 380 109120 400
rect 109380 380 109620 400
rect 109880 380 110120 400
rect 110380 380 110620 400
rect 110880 380 111120 400
rect 111380 380 111620 400
rect 111880 380 112120 400
rect 112380 380 112620 400
rect 112880 380 113120 400
rect 113380 380 113620 400
rect 113880 380 114120 400
rect 114380 380 114620 400
rect 114880 380 115120 400
rect 115380 380 115620 400
rect 115880 380 116120 400
rect 116380 380 116620 400
rect 116880 380 117120 400
rect 117380 380 117620 400
rect 117880 380 118120 400
rect 118380 380 118620 400
rect 118880 380 119120 400
rect 119380 380 119620 400
rect 119880 380 120120 400
rect 120380 380 120620 400
rect 120880 380 121120 400
rect 121380 380 121620 400
rect 121880 380 122120 400
rect 122380 380 122620 400
rect 122880 380 123120 400
rect 123380 380 123620 400
rect 123880 380 124120 400
rect 124380 380 124620 400
rect 124880 380 125120 400
rect 125380 380 125620 400
rect 125880 380 126120 400
rect 126380 380 126620 400
rect 126880 380 127120 400
rect 127380 380 127620 400
rect 127880 380 128120 400
rect 128380 380 128620 400
rect 128880 380 129120 400
rect 129380 380 129620 400
rect 129880 380 130120 400
rect 130380 380 130620 400
rect 130880 380 131120 400
rect 131380 380 131620 400
rect 131880 380 132120 400
rect 132380 380 132620 400
rect 132880 380 133120 400
rect 133380 380 133620 400
rect 133880 380 134120 400
rect 134380 380 134620 400
rect 134880 380 135120 400
rect 135380 380 135620 400
rect 135880 380 136120 400
rect 136380 380 136620 400
rect 136880 380 137120 400
rect 137380 380 137620 400
rect 137880 380 138120 400
rect 138380 380 138620 400
rect 138880 380 139120 400
rect 139380 380 139620 400
rect 139880 380 140000 400
rect 88000 120 88100 380
rect 88400 120 88600 380
rect 88900 120 89100 380
rect 89400 120 89600 380
rect 89900 120 90100 380
rect 90400 120 90600 380
rect 90900 120 91100 380
rect 91400 120 91600 380
rect 91900 120 92100 380
rect 92400 120 92600 380
rect 92900 120 93100 380
rect 93400 120 93600 380
rect 93900 120 94100 380
rect 94400 120 94600 380
rect 94900 120 95100 380
rect 95400 120 95600 380
rect 95900 120 96100 380
rect 96400 120 96600 380
rect 96900 120 97100 380
rect 97400 120 97600 380
rect 97900 120 98100 380
rect 98400 120 98600 380
rect 98900 120 99100 380
rect 99400 120 99600 380
rect 99900 120 100100 380
rect 100400 120 100600 380
rect 100900 120 101100 380
rect 101400 120 101600 380
rect 101900 120 102100 380
rect 102400 120 102600 380
rect 102900 120 103100 380
rect 103400 120 103600 380
rect 103900 120 104100 380
rect 104400 120 104600 380
rect 104900 120 105100 380
rect 105400 120 105600 380
rect 105900 120 106100 380
rect 106400 120 106600 380
rect 106900 120 107100 380
rect 107400 120 107600 380
rect 107900 120 108100 380
rect 108400 120 108600 380
rect 108900 120 109100 380
rect 109400 120 109600 380
rect 109900 120 110100 380
rect 110400 120 110600 380
rect 110900 120 111100 380
rect 111400 120 111600 380
rect 111900 120 112100 380
rect 112400 120 112600 380
rect 112900 120 113100 380
rect 113400 120 113600 380
rect 113900 120 114100 380
rect 114400 120 114600 380
rect 114900 120 115100 380
rect 115400 120 115600 380
rect 115900 120 116100 380
rect 116400 120 116600 380
rect 116900 120 117100 380
rect 117400 120 117600 380
rect 117900 120 118100 380
rect 118400 120 118600 380
rect 118900 120 119100 380
rect 119400 120 119600 380
rect 119900 120 120100 380
rect 120400 120 120600 380
rect 120900 120 121100 380
rect 121400 120 121600 380
rect 121900 120 122100 380
rect 122400 120 122600 380
rect 122900 120 123100 380
rect 123400 120 123600 380
rect 123900 120 124100 380
rect 124400 120 124600 380
rect 124900 120 125100 380
rect 125400 120 125600 380
rect 125900 120 126100 380
rect 126400 120 126600 380
rect 126900 120 127100 380
rect 127400 120 127600 380
rect 127900 120 128100 380
rect 128400 120 128600 380
rect 128900 120 129100 380
rect 129400 120 129600 380
rect 129900 120 130100 380
rect 130400 120 130600 380
rect 130900 120 131100 380
rect 131400 120 131600 380
rect 131900 120 132100 380
rect 132400 120 132600 380
rect 132900 120 133100 380
rect 133400 120 133600 380
rect 133900 120 134100 380
rect 134400 120 134600 380
rect 134900 120 135100 380
rect 135400 120 135600 380
rect 135900 350 136100 380
rect 135900 150 136020 350
rect 136090 150 136100 350
rect 135900 120 136100 150
rect 136400 350 136600 380
rect 136400 150 136410 350
rect 136480 150 136520 350
rect 136590 150 136600 350
rect 136400 120 136600 150
rect 136900 350 137100 380
rect 136900 150 136910 350
rect 136980 150 137020 350
rect 137090 150 137100 350
rect 136900 120 137100 150
rect 137400 350 137600 380
rect 137400 150 137410 350
rect 137480 150 137520 350
rect 137590 150 137600 350
rect 137400 120 137600 150
rect 137900 350 138100 380
rect 137900 150 137910 350
rect 137980 150 138020 350
rect 138090 150 138100 350
rect 137900 120 138100 150
rect 138400 350 138600 380
rect 138400 150 138410 350
rect 138480 150 138520 350
rect 138590 150 138600 350
rect 138400 120 138600 150
rect 138900 350 139100 380
rect 138900 150 138910 350
rect 138980 150 139020 350
rect 139090 150 139100 350
rect 138900 120 139100 150
rect 139400 350 139600 380
rect 139400 150 139410 350
rect 139480 150 139520 350
rect 139590 150 139600 350
rect 139400 120 139600 150
rect 139900 350 140000 380
rect 139900 150 139910 350
rect 139980 150 140000 350
rect 139900 120 140000 150
rect 88000 100 88120 120
rect 88380 100 88620 120
rect 88880 100 89120 120
rect 89380 100 89620 120
rect 89880 100 90120 120
rect 90380 100 90620 120
rect 90880 100 91120 120
rect 91380 100 91620 120
rect 91880 100 92120 120
rect 92380 100 92620 120
rect 92880 100 93120 120
rect 93380 100 93620 120
rect 93880 100 94120 120
rect 94380 100 94620 120
rect 94880 100 95120 120
rect 95380 100 95620 120
rect 95880 100 96120 120
rect 96380 100 96620 120
rect 96880 100 97120 120
rect 97380 100 97620 120
rect 97880 100 98120 120
rect 98380 100 98620 120
rect 98880 100 99120 120
rect 99380 100 99620 120
rect 99880 100 100120 120
rect 100380 100 100620 120
rect 100880 100 101120 120
rect 101380 100 101620 120
rect 101880 100 102120 120
rect 102380 100 102620 120
rect 102880 100 103120 120
rect 103380 100 103620 120
rect 103880 100 104120 120
rect 104380 100 104620 120
rect 104880 100 105120 120
rect 105380 100 105620 120
rect 105880 100 106120 120
rect 106380 100 106620 120
rect 106880 100 107120 120
rect 107380 100 107620 120
rect 107880 100 108120 120
rect 108380 100 108620 120
rect 108880 100 109120 120
rect 109380 100 109620 120
rect 109880 100 110120 120
rect 110380 100 110620 120
rect 110880 100 111120 120
rect 111380 100 111620 120
rect 111880 100 112120 120
rect 112380 100 112620 120
rect 112880 100 113120 120
rect 113380 100 113620 120
rect 113880 100 114120 120
rect 114380 100 114620 120
rect 114880 100 115120 120
rect 115380 100 115620 120
rect 115880 100 116120 120
rect 116380 100 116620 120
rect 116880 100 117120 120
rect 117380 100 117620 120
rect 117880 100 118120 120
rect 118380 100 118620 120
rect 118880 100 119120 120
rect 119380 100 119620 120
rect 119880 100 120120 120
rect 120380 100 120620 120
rect 120880 100 121120 120
rect 121380 100 121620 120
rect 121880 100 122120 120
rect 122380 100 122620 120
rect 122880 100 123120 120
rect 123380 100 123620 120
rect 123880 100 124120 120
rect 124380 100 124620 120
rect 124880 100 125120 120
rect 125380 100 125620 120
rect 125880 100 126120 120
rect 126380 100 126620 120
rect 126880 100 127120 120
rect 127380 100 127620 120
rect 127880 100 128120 120
rect 128380 100 128620 120
rect 128880 100 129120 120
rect 129380 100 129620 120
rect 129880 100 130120 120
rect 130380 100 130620 120
rect 130880 100 131120 120
rect 131380 100 131620 120
rect 131880 100 132120 120
rect 132380 100 132620 120
rect 132880 100 133120 120
rect 133380 100 133620 120
rect 133880 100 134120 120
rect 134380 100 134620 120
rect 134880 100 135120 120
rect 135380 100 135620 120
rect 135880 100 136120 120
rect 136380 100 136620 120
rect 136880 100 137120 120
rect 137380 100 137620 120
rect 137880 100 138120 120
rect 138380 100 138620 120
rect 138880 100 139120 120
rect 139380 100 139620 120
rect 139880 100 140000 120
rect 88000 90 140000 100
rect 88000 20 136150 90
rect 136350 20 136650 90
rect 136850 20 137150 90
rect 137350 20 137650 90
rect 137850 20 138150 90
rect 138350 20 138650 90
rect 138850 20 139150 90
rect 139350 20 139650 90
rect 139850 20 140000 90
rect 88000 -20 140000 20
rect 88000 -90 136150 -20
rect 136350 -90 136650 -20
rect 136850 -90 137150 -20
rect 137350 -90 137650 -20
rect 137850 -90 138150 -20
rect 138350 -90 138650 -20
rect 138850 -90 139150 -20
rect 139350 -90 139650 -20
rect 139850 -90 140000 -20
rect 88000 -100 140000 -90
rect 88000 -120 88120 -100
rect 88380 -120 88620 -100
rect 88880 -120 89120 -100
rect 89380 -120 89620 -100
rect 89880 -120 90120 -100
rect 90380 -120 90620 -100
rect 90880 -120 91120 -100
rect 91380 -120 91620 -100
rect 91880 -120 92120 -100
rect 92380 -120 92620 -100
rect 92880 -120 93120 -100
rect 93380 -120 93620 -100
rect 93880 -120 94120 -100
rect 94380 -120 94620 -100
rect 94880 -120 95120 -100
rect 95380 -120 95620 -100
rect 95880 -120 96120 -100
rect 96380 -120 96620 -100
rect 96880 -120 97120 -100
rect 97380 -120 97620 -100
rect 97880 -120 98120 -100
rect 98380 -120 98620 -100
rect 98880 -120 99120 -100
rect 99380 -120 99620 -100
rect 99880 -120 100120 -100
rect 100380 -120 100620 -100
rect 100880 -120 101120 -100
rect 101380 -120 101620 -100
rect 101880 -120 102120 -100
rect 102380 -120 102620 -100
rect 102880 -120 103120 -100
rect 103380 -120 103620 -100
rect 103880 -120 104120 -100
rect 104380 -120 104620 -100
rect 104880 -120 105120 -100
rect 105380 -120 105620 -100
rect 105880 -120 106120 -100
rect 106380 -120 106620 -100
rect 106880 -120 107120 -100
rect 107380 -120 107620 -100
rect 107880 -120 108120 -100
rect 108380 -120 108620 -100
rect 108880 -120 109120 -100
rect 109380 -120 109620 -100
rect 109880 -120 110120 -100
rect 110380 -120 110620 -100
rect 110880 -120 111120 -100
rect 111380 -120 111620 -100
rect 111880 -120 112120 -100
rect 112380 -120 112620 -100
rect 112880 -120 113120 -100
rect 113380 -120 113620 -100
rect 113880 -120 114120 -100
rect 114380 -120 114620 -100
rect 114880 -120 115120 -100
rect 115380 -120 115620 -100
rect 115880 -120 116120 -100
rect 116380 -120 116620 -100
rect 116880 -120 117120 -100
rect 117380 -120 117620 -100
rect 117880 -120 118120 -100
rect 118380 -120 118620 -100
rect 118880 -120 119120 -100
rect 119380 -120 119620 -100
rect 119880 -120 120120 -100
rect 120380 -120 120620 -100
rect 120880 -120 121120 -100
rect 121380 -120 121620 -100
rect 121880 -120 122120 -100
rect 122380 -120 122620 -100
rect 122880 -120 123120 -100
rect 123380 -120 123620 -100
rect 123880 -120 124120 -100
rect 124380 -120 124620 -100
rect 124880 -120 125120 -100
rect 125380 -120 125620 -100
rect 125880 -120 126120 -100
rect 126380 -120 126620 -100
rect 126880 -120 127120 -100
rect 127380 -120 127620 -100
rect 127880 -120 128120 -100
rect 128380 -120 128620 -100
rect 128880 -120 129120 -100
rect 129380 -120 129620 -100
rect 129880 -120 130120 -100
rect 130380 -120 130620 -100
rect 130880 -120 131120 -100
rect 131380 -120 131620 -100
rect 131880 -120 132120 -100
rect 132380 -120 132620 -100
rect 132880 -120 133120 -100
rect 133380 -120 133620 -100
rect 133880 -120 134120 -100
rect 134380 -120 134620 -100
rect 134880 -120 135120 -100
rect 135380 -120 135620 -100
rect 135880 -120 136120 -100
rect 136380 -120 136620 -100
rect 136880 -120 137120 -100
rect 137380 -120 137620 -100
rect 137880 -120 138120 -100
rect 138380 -120 138620 -100
rect 138880 -120 139120 -100
rect 139380 -120 139620 -100
rect 139880 -120 140000 -100
rect 88000 -380 88100 -120
rect 88400 -380 88600 -120
rect 88900 -380 89100 -120
rect 89400 -380 89600 -120
rect 89900 -380 90100 -120
rect 90400 -380 90600 -120
rect 90900 -380 91100 -120
rect 91400 -380 91600 -120
rect 91900 -380 92100 -120
rect 92400 -380 92600 -120
rect 92900 -380 93100 -120
rect 93400 -380 93600 -120
rect 93900 -380 94100 -120
rect 94400 -380 94600 -120
rect 94900 -380 95100 -120
rect 95400 -380 95600 -120
rect 95900 -380 96100 -120
rect 96400 -380 96600 -120
rect 96900 -380 97100 -120
rect 97400 -380 97600 -120
rect 97900 -380 98100 -120
rect 98400 -380 98600 -120
rect 98900 -380 99100 -120
rect 99400 -380 99600 -120
rect 99900 -380 100100 -120
rect 100400 -380 100600 -120
rect 100900 -380 101100 -120
rect 101400 -380 101600 -120
rect 101900 -380 102100 -120
rect 102400 -380 102600 -120
rect 102900 -380 103100 -120
rect 103400 -380 103600 -120
rect 103900 -380 104100 -120
rect 104400 -380 104600 -120
rect 104900 -380 105100 -120
rect 105400 -380 105600 -120
rect 105900 -380 106100 -120
rect 106400 -380 106600 -120
rect 106900 -380 107100 -120
rect 107400 -380 107600 -120
rect 107900 -380 108100 -120
rect 108400 -380 108600 -120
rect 108900 -380 109100 -120
rect 109400 -380 109600 -120
rect 109900 -380 110100 -120
rect 110400 -380 110600 -120
rect 110900 -380 111100 -120
rect 111400 -380 111600 -120
rect 111900 -380 112100 -120
rect 112400 -380 112600 -120
rect 112900 -380 113100 -120
rect 113400 -380 113600 -120
rect 113900 -380 114100 -120
rect 114400 -380 114600 -120
rect 114900 -380 115100 -120
rect 115400 -380 115600 -120
rect 115900 -380 116100 -120
rect 116400 -380 116600 -120
rect 116900 -380 117100 -120
rect 117400 -380 117600 -120
rect 117900 -380 118100 -120
rect 118400 -380 118600 -120
rect 118900 -380 119100 -120
rect 119400 -380 119600 -120
rect 119900 -380 120100 -120
rect 120400 -380 120600 -120
rect 120900 -380 121100 -120
rect 121400 -380 121600 -120
rect 121900 -380 122100 -120
rect 122400 -380 122600 -120
rect 122900 -380 123100 -120
rect 123400 -380 123600 -120
rect 123900 -380 124100 -120
rect 124400 -380 124600 -120
rect 124900 -380 125100 -120
rect 125400 -380 125600 -120
rect 125900 -380 126100 -120
rect 126400 -380 126600 -120
rect 126900 -380 127100 -120
rect 127400 -380 127600 -120
rect 127900 -380 128100 -120
rect 128400 -380 128600 -120
rect 128900 -380 129100 -120
rect 129400 -380 129600 -120
rect 129900 -380 130100 -120
rect 130400 -380 130600 -120
rect 130900 -380 131100 -120
rect 131400 -380 131600 -120
rect 131900 -380 132100 -120
rect 132400 -380 132600 -120
rect 132900 -380 133100 -120
rect 133400 -380 133600 -120
rect 133900 -380 134100 -120
rect 134400 -380 134600 -120
rect 134900 -380 135100 -120
rect 135400 -380 135600 -120
rect 135900 -150 136100 -120
rect 135900 -350 136020 -150
rect 136090 -350 136100 -150
rect 135900 -380 136100 -350
rect 136400 -150 136600 -120
rect 136400 -350 136410 -150
rect 136480 -350 136520 -150
rect 136590 -350 136600 -150
rect 136400 -380 136600 -350
rect 136900 -150 137100 -120
rect 136900 -350 136910 -150
rect 136980 -350 137020 -150
rect 137090 -350 137100 -150
rect 136900 -380 137100 -350
rect 137400 -150 137600 -120
rect 137400 -350 137410 -150
rect 137480 -350 137520 -150
rect 137590 -350 137600 -150
rect 137400 -380 137600 -350
rect 137900 -150 138100 -120
rect 137900 -350 137910 -150
rect 137980 -350 138020 -150
rect 138090 -350 138100 -150
rect 137900 -380 138100 -350
rect 138400 -150 138600 -120
rect 138400 -350 138410 -150
rect 138480 -350 138520 -150
rect 138590 -350 138600 -150
rect 138400 -380 138600 -350
rect 138900 -150 139100 -120
rect 138900 -350 138910 -150
rect 138980 -350 139020 -150
rect 139090 -350 139100 -150
rect 138900 -380 139100 -350
rect 139400 -150 139600 -120
rect 139400 -350 139410 -150
rect 139480 -350 139520 -150
rect 139590 -350 139600 -150
rect 139400 -380 139600 -350
rect 139900 -150 140000 -120
rect 139900 -350 139910 -150
rect 139980 -350 140000 -150
rect 139900 -380 140000 -350
rect 88000 -400 88120 -380
rect 88380 -400 88620 -380
rect 88880 -400 89120 -380
rect 89380 -400 89620 -380
rect 89880 -400 90120 -380
rect 90380 -400 90620 -380
rect 90880 -400 91120 -380
rect 91380 -400 91620 -380
rect 91880 -400 92120 -380
rect 92380 -400 92620 -380
rect 92880 -400 93120 -380
rect 93380 -400 93620 -380
rect 93880 -400 94120 -380
rect 94380 -400 94620 -380
rect 94880 -400 95120 -380
rect 95380 -400 95620 -380
rect 95880 -400 96120 -380
rect 96380 -400 96620 -380
rect 96880 -400 97120 -380
rect 97380 -400 97620 -380
rect 97880 -400 98120 -380
rect 98380 -400 98620 -380
rect 98880 -400 99120 -380
rect 99380 -400 99620 -380
rect 99880 -400 100120 -380
rect 100380 -400 100620 -380
rect 100880 -400 101120 -380
rect 101380 -400 101620 -380
rect 101880 -400 102120 -380
rect 102380 -400 102620 -380
rect 102880 -400 103120 -380
rect 103380 -400 103620 -380
rect 103880 -400 104120 -380
rect 104380 -400 104620 -380
rect 104880 -400 105120 -380
rect 105380 -400 105620 -380
rect 105880 -400 106120 -380
rect 106380 -400 106620 -380
rect 106880 -400 107120 -380
rect 107380 -400 107620 -380
rect 107880 -400 108120 -380
rect 108380 -400 108620 -380
rect 108880 -400 109120 -380
rect 109380 -400 109620 -380
rect 109880 -400 110120 -380
rect 110380 -400 110620 -380
rect 110880 -400 111120 -380
rect 111380 -400 111620 -380
rect 111880 -400 112120 -380
rect 112380 -400 112620 -380
rect 112880 -400 113120 -380
rect 113380 -400 113620 -380
rect 113880 -400 114120 -380
rect 114380 -400 114620 -380
rect 114880 -400 115120 -380
rect 115380 -400 115620 -380
rect 115880 -400 116120 -380
rect 116380 -400 116620 -380
rect 116880 -400 117120 -380
rect 117380 -400 117620 -380
rect 117880 -400 118120 -380
rect 118380 -400 118620 -380
rect 118880 -400 119120 -380
rect 119380 -400 119620 -380
rect 119880 -400 120120 -380
rect 120380 -400 120620 -380
rect 120880 -400 121120 -380
rect 121380 -400 121620 -380
rect 121880 -400 122120 -380
rect 122380 -400 122620 -380
rect 122880 -400 123120 -380
rect 123380 -400 123620 -380
rect 123880 -400 124120 -380
rect 124380 -400 124620 -380
rect 124880 -400 125120 -380
rect 125380 -400 125620 -380
rect 125880 -400 126120 -380
rect 126380 -400 126620 -380
rect 126880 -400 127120 -380
rect 127380 -400 127620 -380
rect 127880 -400 128120 -380
rect 128380 -400 128620 -380
rect 128880 -400 129120 -380
rect 129380 -400 129620 -380
rect 129880 -400 130120 -380
rect 130380 -400 130620 -380
rect 130880 -400 131120 -380
rect 131380 -400 131620 -380
rect 131880 -400 132120 -380
rect 132380 -400 132620 -380
rect 132880 -400 133120 -380
rect 133380 -400 133620 -380
rect 133880 -400 134120 -380
rect 134380 -400 134620 -380
rect 134880 -400 135120 -380
rect 135380 -400 135620 -380
rect 135880 -400 136120 -380
rect 136380 -400 136620 -380
rect 136880 -400 137120 -380
rect 137380 -400 137620 -380
rect 137880 -400 138120 -380
rect 138380 -400 138620 -380
rect 138880 -400 139120 -380
rect 139380 -400 139620 -380
rect 139880 -400 140000 -380
rect 88000 -410 140000 -400
rect 88000 -480 136150 -410
rect 136350 -480 136650 -410
rect 136850 -480 137150 -410
rect 137350 -480 137650 -410
rect 137850 -480 138150 -410
rect 138350 -480 138650 -410
rect 138850 -480 139150 -410
rect 139350 -480 139650 -410
rect 139850 -480 140000 -410
rect 88000 -520 140000 -480
rect 88000 -590 136150 -520
rect 136350 -590 136650 -520
rect 136850 -590 137150 -520
rect 137350 -590 137650 -520
rect 137850 -590 138150 -520
rect 138350 -590 138650 -520
rect 138850 -590 139150 -520
rect 139350 -590 139650 -520
rect 139850 -590 140000 -520
rect 88000 -600 140000 -590
rect 88000 -620 88120 -600
rect 88380 -620 88620 -600
rect 88880 -620 89120 -600
rect 89380 -620 89620 -600
rect 89880 -620 90120 -600
rect 90380 -620 90620 -600
rect 90880 -620 91120 -600
rect 91380 -620 91620 -600
rect 91880 -620 92120 -600
rect 92380 -620 92620 -600
rect 92880 -620 93120 -600
rect 93380 -620 93620 -600
rect 93880 -620 94120 -600
rect 94380 -620 94620 -600
rect 94880 -620 95120 -600
rect 95380 -620 95620 -600
rect 95880 -620 96120 -600
rect 96380 -620 96620 -600
rect 96880 -620 97120 -600
rect 97380 -620 97620 -600
rect 97880 -620 98120 -600
rect 98380 -620 98620 -600
rect 98880 -620 99120 -600
rect 99380 -620 99620 -600
rect 99880 -620 100120 -600
rect 100380 -620 100620 -600
rect 100880 -620 101120 -600
rect 101380 -620 101620 -600
rect 101880 -620 102120 -600
rect 102380 -620 102620 -600
rect 102880 -620 103120 -600
rect 103380 -620 103620 -600
rect 103880 -620 104120 -600
rect 104380 -620 104620 -600
rect 104880 -620 105120 -600
rect 105380 -620 105620 -600
rect 105880 -620 106120 -600
rect 106380 -620 106620 -600
rect 106880 -620 107120 -600
rect 107380 -620 107620 -600
rect 107880 -620 108120 -600
rect 108380 -620 108620 -600
rect 108880 -620 109120 -600
rect 109380 -620 109620 -600
rect 109880 -620 110120 -600
rect 110380 -620 110620 -600
rect 110880 -620 111120 -600
rect 111380 -620 111620 -600
rect 111880 -620 112120 -600
rect 112380 -620 112620 -600
rect 112880 -620 113120 -600
rect 113380 -620 113620 -600
rect 113880 -620 114120 -600
rect 114380 -620 114620 -600
rect 114880 -620 115120 -600
rect 115380 -620 115620 -600
rect 115880 -620 116120 -600
rect 116380 -620 116620 -600
rect 116880 -620 117120 -600
rect 117380 -620 117620 -600
rect 117880 -620 118120 -600
rect 118380 -620 118620 -600
rect 118880 -620 119120 -600
rect 119380 -620 119620 -600
rect 119880 -620 120120 -600
rect 120380 -620 120620 -600
rect 120880 -620 121120 -600
rect 121380 -620 121620 -600
rect 121880 -620 122120 -600
rect 122380 -620 122620 -600
rect 122880 -620 123120 -600
rect 123380 -620 123620 -600
rect 123880 -620 124120 -600
rect 124380 -620 124620 -600
rect 124880 -620 125120 -600
rect 125380 -620 125620 -600
rect 125880 -620 126120 -600
rect 126380 -620 126620 -600
rect 126880 -620 127120 -600
rect 127380 -620 127620 -600
rect 127880 -620 128120 -600
rect 128380 -620 128620 -600
rect 128880 -620 129120 -600
rect 129380 -620 129620 -600
rect 129880 -620 130120 -600
rect 130380 -620 130620 -600
rect 130880 -620 131120 -600
rect 131380 -620 131620 -600
rect 131880 -620 132120 -600
rect 132380 -620 132620 -600
rect 132880 -620 133120 -600
rect 133380 -620 133620 -600
rect 133880 -620 134120 -600
rect 134380 -620 134620 -600
rect 134880 -620 135120 -600
rect 135380 -620 135620 -600
rect 135880 -620 136120 -600
rect 136380 -620 136620 -600
rect 136880 -620 137120 -600
rect 137380 -620 137620 -600
rect 137880 -620 138120 -600
rect 138380 -620 138620 -600
rect 138880 -620 139120 -600
rect 139380 -620 139620 -600
rect 139880 -620 140000 -600
rect 88000 -880 88100 -620
rect 88400 -880 88600 -620
rect 88900 -880 89100 -620
rect 89400 -880 89600 -620
rect 89900 -880 90100 -620
rect 90400 -880 90600 -620
rect 90900 -880 91100 -620
rect 91400 -880 91600 -620
rect 91900 -880 92100 -620
rect 92400 -880 92600 -620
rect 92900 -880 93100 -620
rect 93400 -880 93600 -620
rect 93900 -880 94100 -620
rect 94400 -880 94600 -620
rect 94900 -880 95100 -620
rect 95400 -880 95600 -620
rect 95900 -880 96100 -620
rect 96400 -880 96600 -620
rect 96900 -880 97100 -620
rect 97400 -880 97600 -620
rect 97900 -880 98100 -620
rect 98400 -880 98600 -620
rect 98900 -880 99100 -620
rect 99400 -880 99600 -620
rect 99900 -880 100100 -620
rect 100400 -880 100600 -620
rect 100900 -880 101100 -620
rect 101400 -880 101600 -620
rect 101900 -880 102100 -620
rect 102400 -880 102600 -620
rect 102900 -880 103100 -620
rect 103400 -880 103600 -620
rect 103900 -880 104100 -620
rect 104400 -880 104600 -620
rect 104900 -880 105100 -620
rect 105400 -880 105600 -620
rect 105900 -880 106100 -620
rect 106400 -880 106600 -620
rect 106900 -880 107100 -620
rect 107400 -880 107600 -620
rect 107900 -880 108100 -620
rect 108400 -880 108600 -620
rect 108900 -880 109100 -620
rect 109400 -880 109600 -620
rect 109900 -880 110100 -620
rect 110400 -880 110600 -620
rect 110900 -880 111100 -620
rect 111400 -880 111600 -620
rect 111900 -880 112100 -620
rect 112400 -880 112600 -620
rect 112900 -880 113100 -620
rect 113400 -880 113600 -620
rect 113900 -880 114100 -620
rect 114400 -880 114600 -620
rect 114900 -880 115100 -620
rect 115400 -880 115600 -620
rect 115900 -880 116100 -620
rect 116400 -880 116600 -620
rect 116900 -880 117100 -620
rect 117400 -880 117600 -620
rect 117900 -880 118100 -620
rect 118400 -880 118600 -620
rect 118900 -880 119100 -620
rect 119400 -880 119600 -620
rect 119900 -880 120100 -620
rect 120400 -880 120600 -620
rect 120900 -880 121100 -620
rect 121400 -880 121600 -620
rect 121900 -880 122100 -620
rect 122400 -880 122600 -620
rect 122900 -880 123100 -620
rect 123400 -880 123600 -620
rect 123900 -880 124100 -620
rect 124400 -880 124600 -620
rect 124900 -880 125100 -620
rect 125400 -880 125600 -620
rect 125900 -880 126100 -620
rect 126400 -880 126600 -620
rect 126900 -880 127100 -620
rect 127400 -880 127600 -620
rect 127900 -880 128100 -620
rect 128400 -880 128600 -620
rect 128900 -880 129100 -620
rect 129400 -880 129600 -620
rect 129900 -880 130100 -620
rect 130400 -880 130600 -620
rect 130900 -880 131100 -620
rect 131400 -880 131600 -620
rect 131900 -880 132100 -620
rect 132400 -880 132600 -620
rect 132900 -880 133100 -620
rect 133400 -880 133600 -620
rect 133900 -880 134100 -620
rect 134400 -880 134600 -620
rect 134900 -880 135100 -620
rect 135400 -880 135600 -620
rect 135900 -650 136100 -620
rect 135900 -850 136020 -650
rect 136090 -850 136100 -650
rect 135900 -880 136100 -850
rect 136400 -650 136600 -620
rect 136400 -850 136410 -650
rect 136480 -850 136520 -650
rect 136590 -850 136600 -650
rect 136400 -880 136600 -850
rect 136900 -650 137100 -620
rect 136900 -850 136910 -650
rect 136980 -850 137020 -650
rect 137090 -850 137100 -650
rect 136900 -880 137100 -850
rect 137400 -650 137600 -620
rect 137400 -850 137410 -650
rect 137480 -850 137520 -650
rect 137590 -850 137600 -650
rect 137400 -880 137600 -850
rect 137900 -650 138100 -620
rect 137900 -850 137910 -650
rect 137980 -850 138020 -650
rect 138090 -850 138100 -650
rect 137900 -880 138100 -850
rect 138400 -650 138600 -620
rect 138400 -850 138410 -650
rect 138480 -850 138520 -650
rect 138590 -850 138600 -650
rect 138400 -880 138600 -850
rect 138900 -650 139100 -620
rect 138900 -850 138910 -650
rect 138980 -850 139020 -650
rect 139090 -850 139100 -650
rect 138900 -880 139100 -850
rect 139400 -650 139600 -620
rect 139400 -850 139410 -650
rect 139480 -850 139520 -650
rect 139590 -850 139600 -650
rect 139400 -880 139600 -850
rect 139900 -650 140000 -620
rect 139900 -850 139910 -650
rect 139980 -850 140000 -650
rect 139900 -880 140000 -850
rect 88000 -900 88120 -880
rect 88380 -900 88620 -880
rect 88880 -900 89120 -880
rect 89380 -900 89620 -880
rect 89880 -900 90120 -880
rect 90380 -900 90620 -880
rect 90880 -900 91120 -880
rect 91380 -900 91620 -880
rect 91880 -900 92120 -880
rect 92380 -900 92620 -880
rect 92880 -900 93120 -880
rect 93380 -900 93620 -880
rect 93880 -900 94120 -880
rect 94380 -900 94620 -880
rect 94880 -900 95120 -880
rect 95380 -900 95620 -880
rect 95880 -900 96120 -880
rect 96380 -900 96620 -880
rect 96880 -900 97120 -880
rect 97380 -900 97620 -880
rect 97880 -900 98120 -880
rect 98380 -900 98620 -880
rect 98880 -900 99120 -880
rect 99380 -900 99620 -880
rect 99880 -900 100120 -880
rect 100380 -900 100620 -880
rect 100880 -900 101120 -880
rect 101380 -900 101620 -880
rect 101880 -900 102120 -880
rect 102380 -900 102620 -880
rect 102880 -900 103120 -880
rect 103380 -900 103620 -880
rect 103880 -900 104120 -880
rect 104380 -900 104620 -880
rect 104880 -900 105120 -880
rect 105380 -900 105620 -880
rect 105880 -900 106120 -880
rect 106380 -900 106620 -880
rect 106880 -900 107120 -880
rect 107380 -900 107620 -880
rect 107880 -900 108120 -880
rect 108380 -900 108620 -880
rect 108880 -900 109120 -880
rect 109380 -900 109620 -880
rect 109880 -900 110120 -880
rect 110380 -900 110620 -880
rect 110880 -900 111120 -880
rect 111380 -900 111620 -880
rect 111880 -900 112120 -880
rect 112380 -900 112620 -880
rect 112880 -900 113120 -880
rect 113380 -900 113620 -880
rect 113880 -900 114120 -880
rect 114380 -900 114620 -880
rect 114880 -900 115120 -880
rect 115380 -900 115620 -880
rect 115880 -900 116120 -880
rect 116380 -900 116620 -880
rect 116880 -900 117120 -880
rect 117380 -900 117620 -880
rect 117880 -900 118120 -880
rect 118380 -900 118620 -880
rect 118880 -900 119120 -880
rect 119380 -900 119620 -880
rect 119880 -900 120120 -880
rect 120380 -900 120620 -880
rect 120880 -900 121120 -880
rect 121380 -900 121620 -880
rect 121880 -900 122120 -880
rect 122380 -900 122620 -880
rect 122880 -900 123120 -880
rect 123380 -900 123620 -880
rect 123880 -900 124120 -880
rect 124380 -900 124620 -880
rect 124880 -900 125120 -880
rect 125380 -900 125620 -880
rect 125880 -900 126120 -880
rect 126380 -900 126620 -880
rect 126880 -900 127120 -880
rect 127380 -900 127620 -880
rect 127880 -900 128120 -880
rect 128380 -900 128620 -880
rect 128880 -900 129120 -880
rect 129380 -900 129620 -880
rect 129880 -900 130120 -880
rect 130380 -900 130620 -880
rect 130880 -900 131120 -880
rect 131380 -900 131620 -880
rect 131880 -900 132120 -880
rect 132380 -900 132620 -880
rect 132880 -900 133120 -880
rect 133380 -900 133620 -880
rect 133880 -900 134120 -880
rect 134380 -900 134620 -880
rect 134880 -900 135120 -880
rect 135380 -900 135620 -880
rect 135880 -900 136120 -880
rect 136380 -900 136620 -880
rect 136880 -900 137120 -880
rect 137380 -900 137620 -880
rect 137880 -900 138120 -880
rect 138380 -900 138620 -880
rect 138880 -900 139120 -880
rect 139380 -900 139620 -880
rect 139880 -900 140000 -880
rect 88000 -910 140000 -900
rect 88000 -980 136150 -910
rect 136350 -980 136650 -910
rect 136850 -980 137150 -910
rect 137350 -980 137650 -910
rect 137850 -980 138150 -910
rect 138350 -980 138650 -910
rect 138850 -980 139150 -910
rect 139350 -980 139650 -910
rect 139850 -980 140000 -910
rect 88000 -1020 140000 -980
rect 88000 -1090 136150 -1020
rect 136350 -1090 136650 -1020
rect 136850 -1090 137150 -1020
rect 137350 -1090 137650 -1020
rect 137850 -1090 138150 -1020
rect 138350 -1090 138650 -1020
rect 138850 -1090 139150 -1020
rect 139350 -1090 139650 -1020
rect 139850 -1090 140000 -1020
rect 88000 -1100 140000 -1090
rect 88000 -1120 88120 -1100
rect 88380 -1120 88620 -1100
rect 88880 -1120 89120 -1100
rect 89380 -1120 89620 -1100
rect 89880 -1120 90120 -1100
rect 90380 -1120 90620 -1100
rect 90880 -1120 91120 -1100
rect 91380 -1120 91620 -1100
rect 91880 -1120 92120 -1100
rect 92380 -1120 92620 -1100
rect 92880 -1120 93120 -1100
rect 93380 -1120 93620 -1100
rect 93880 -1120 94120 -1100
rect 94380 -1120 94620 -1100
rect 94880 -1120 95120 -1100
rect 95380 -1120 95620 -1100
rect 95880 -1120 96120 -1100
rect 96380 -1120 96620 -1100
rect 96880 -1120 97120 -1100
rect 97380 -1120 97620 -1100
rect 97880 -1120 98120 -1100
rect 98380 -1120 98620 -1100
rect 98880 -1120 99120 -1100
rect 99380 -1120 99620 -1100
rect 99880 -1120 100120 -1100
rect 100380 -1120 100620 -1100
rect 100880 -1120 101120 -1100
rect 101380 -1120 101620 -1100
rect 101880 -1120 102120 -1100
rect 102380 -1120 102620 -1100
rect 102880 -1120 103120 -1100
rect 103380 -1120 103620 -1100
rect 103880 -1120 104120 -1100
rect 104380 -1120 104620 -1100
rect 104880 -1120 105120 -1100
rect 105380 -1120 105620 -1100
rect 105880 -1120 106120 -1100
rect 106380 -1120 106620 -1100
rect 106880 -1120 107120 -1100
rect 107380 -1120 107620 -1100
rect 107880 -1120 108120 -1100
rect 108380 -1120 108620 -1100
rect 108880 -1120 109120 -1100
rect 109380 -1120 109620 -1100
rect 109880 -1120 110120 -1100
rect 110380 -1120 110620 -1100
rect 110880 -1120 111120 -1100
rect 111380 -1120 111620 -1100
rect 111880 -1120 112120 -1100
rect 112380 -1120 112620 -1100
rect 112880 -1120 113120 -1100
rect 113380 -1120 113620 -1100
rect 113880 -1120 114120 -1100
rect 114380 -1120 114620 -1100
rect 114880 -1120 115120 -1100
rect 115380 -1120 115620 -1100
rect 115880 -1120 116120 -1100
rect 116380 -1120 116620 -1100
rect 116880 -1120 117120 -1100
rect 117380 -1120 117620 -1100
rect 117880 -1120 118120 -1100
rect 118380 -1120 118620 -1100
rect 118880 -1120 119120 -1100
rect 119380 -1120 119620 -1100
rect 119880 -1120 120120 -1100
rect 120380 -1120 120620 -1100
rect 120880 -1120 121120 -1100
rect 121380 -1120 121620 -1100
rect 121880 -1120 122120 -1100
rect 122380 -1120 122620 -1100
rect 122880 -1120 123120 -1100
rect 123380 -1120 123620 -1100
rect 123880 -1120 124120 -1100
rect 124380 -1120 124620 -1100
rect 124880 -1120 125120 -1100
rect 125380 -1120 125620 -1100
rect 125880 -1120 126120 -1100
rect 126380 -1120 126620 -1100
rect 126880 -1120 127120 -1100
rect 127380 -1120 127620 -1100
rect 127880 -1120 128120 -1100
rect 128380 -1120 128620 -1100
rect 128880 -1120 129120 -1100
rect 129380 -1120 129620 -1100
rect 129880 -1120 130120 -1100
rect 130380 -1120 130620 -1100
rect 130880 -1120 131120 -1100
rect 131380 -1120 131620 -1100
rect 131880 -1120 132120 -1100
rect 132380 -1120 132620 -1100
rect 132880 -1120 133120 -1100
rect 133380 -1120 133620 -1100
rect 133880 -1120 134120 -1100
rect 134380 -1120 134620 -1100
rect 134880 -1120 135120 -1100
rect 135380 -1120 135620 -1100
rect 135880 -1120 136120 -1100
rect 136380 -1120 136620 -1100
rect 136880 -1120 137120 -1100
rect 137380 -1120 137620 -1100
rect 137880 -1120 138120 -1100
rect 138380 -1120 138620 -1100
rect 138880 -1120 139120 -1100
rect 139380 -1120 139620 -1100
rect 139880 -1120 140000 -1100
rect 88000 -1380 88100 -1120
rect 88400 -1380 88600 -1120
rect 88900 -1380 89100 -1120
rect 89400 -1380 89600 -1120
rect 89900 -1380 90100 -1120
rect 90400 -1380 90600 -1120
rect 90900 -1380 91100 -1120
rect 91400 -1380 91600 -1120
rect 91900 -1380 92100 -1120
rect 92400 -1380 92600 -1120
rect 92900 -1380 93100 -1120
rect 93400 -1380 93600 -1120
rect 93900 -1380 94100 -1120
rect 94400 -1380 94600 -1120
rect 94900 -1380 95100 -1120
rect 95400 -1380 95600 -1120
rect 95900 -1380 96100 -1120
rect 96400 -1380 96600 -1120
rect 96900 -1380 97100 -1120
rect 97400 -1380 97600 -1120
rect 97900 -1380 98100 -1120
rect 98400 -1380 98600 -1120
rect 98900 -1380 99100 -1120
rect 99400 -1380 99600 -1120
rect 99900 -1380 100100 -1120
rect 100400 -1380 100600 -1120
rect 100900 -1380 101100 -1120
rect 101400 -1380 101600 -1120
rect 101900 -1380 102100 -1120
rect 102400 -1380 102600 -1120
rect 102900 -1380 103100 -1120
rect 103400 -1380 103600 -1120
rect 103900 -1380 104100 -1120
rect 104400 -1380 104600 -1120
rect 104900 -1380 105100 -1120
rect 105400 -1380 105600 -1120
rect 105900 -1380 106100 -1120
rect 106400 -1380 106600 -1120
rect 106900 -1380 107100 -1120
rect 107400 -1380 107600 -1120
rect 107900 -1380 108100 -1120
rect 108400 -1380 108600 -1120
rect 108900 -1380 109100 -1120
rect 109400 -1380 109600 -1120
rect 109900 -1380 110100 -1120
rect 110400 -1380 110600 -1120
rect 110900 -1380 111100 -1120
rect 111400 -1380 111600 -1120
rect 111900 -1380 112100 -1120
rect 112400 -1380 112600 -1120
rect 112900 -1380 113100 -1120
rect 113400 -1380 113600 -1120
rect 113900 -1380 114100 -1120
rect 114400 -1380 114600 -1120
rect 114900 -1380 115100 -1120
rect 115400 -1380 115600 -1120
rect 115900 -1380 116100 -1120
rect 116400 -1380 116600 -1120
rect 116900 -1380 117100 -1120
rect 117400 -1380 117600 -1120
rect 117900 -1380 118100 -1120
rect 118400 -1380 118600 -1120
rect 118900 -1380 119100 -1120
rect 119400 -1380 119600 -1120
rect 119900 -1380 120100 -1120
rect 120400 -1380 120600 -1120
rect 120900 -1380 121100 -1120
rect 121400 -1380 121600 -1120
rect 121900 -1380 122100 -1120
rect 122400 -1380 122600 -1120
rect 122900 -1380 123100 -1120
rect 123400 -1380 123600 -1120
rect 123900 -1380 124100 -1120
rect 124400 -1380 124600 -1120
rect 124900 -1380 125100 -1120
rect 125400 -1380 125600 -1120
rect 125900 -1380 126100 -1120
rect 126400 -1380 126600 -1120
rect 126900 -1380 127100 -1120
rect 127400 -1380 127600 -1120
rect 127900 -1380 128100 -1120
rect 128400 -1380 128600 -1120
rect 128900 -1380 129100 -1120
rect 129400 -1380 129600 -1120
rect 129900 -1380 130100 -1120
rect 130400 -1380 130600 -1120
rect 130900 -1380 131100 -1120
rect 131400 -1380 131600 -1120
rect 131900 -1380 132100 -1120
rect 132400 -1380 132600 -1120
rect 132900 -1380 133100 -1120
rect 133400 -1380 133600 -1120
rect 133900 -1380 134100 -1120
rect 134400 -1380 134600 -1120
rect 134900 -1380 135100 -1120
rect 135400 -1380 135600 -1120
rect 135900 -1150 136100 -1120
rect 135900 -1350 136020 -1150
rect 136090 -1350 136100 -1150
rect 135900 -1380 136100 -1350
rect 136400 -1150 136600 -1120
rect 136400 -1350 136410 -1150
rect 136480 -1350 136520 -1150
rect 136590 -1350 136600 -1150
rect 136400 -1380 136600 -1350
rect 136900 -1150 137100 -1120
rect 136900 -1350 136910 -1150
rect 136980 -1350 137020 -1150
rect 137090 -1350 137100 -1150
rect 136900 -1380 137100 -1350
rect 137400 -1150 137600 -1120
rect 137400 -1350 137410 -1150
rect 137480 -1350 137520 -1150
rect 137590 -1350 137600 -1150
rect 137400 -1380 137600 -1350
rect 137900 -1150 138100 -1120
rect 137900 -1350 137910 -1150
rect 137980 -1350 138020 -1150
rect 138090 -1350 138100 -1150
rect 137900 -1380 138100 -1350
rect 138400 -1150 138600 -1120
rect 138400 -1350 138410 -1150
rect 138480 -1350 138520 -1150
rect 138590 -1350 138600 -1150
rect 138400 -1380 138600 -1350
rect 138900 -1150 139100 -1120
rect 138900 -1350 138910 -1150
rect 138980 -1350 139020 -1150
rect 139090 -1350 139100 -1150
rect 138900 -1380 139100 -1350
rect 139400 -1150 139600 -1120
rect 139400 -1350 139410 -1150
rect 139480 -1350 139520 -1150
rect 139590 -1350 139600 -1150
rect 139400 -1380 139600 -1350
rect 139900 -1150 140000 -1120
rect 139900 -1350 139910 -1150
rect 139980 -1350 140000 -1150
rect 139900 -1380 140000 -1350
rect 88000 -1400 88120 -1380
rect 88380 -1400 88620 -1380
rect 88880 -1400 89120 -1380
rect 89380 -1400 89620 -1380
rect 89880 -1400 90120 -1380
rect 90380 -1400 90620 -1380
rect 90880 -1400 91120 -1380
rect 91380 -1400 91620 -1380
rect 91880 -1400 92120 -1380
rect 92380 -1400 92620 -1380
rect 92880 -1400 93120 -1380
rect 93380 -1400 93620 -1380
rect 93880 -1400 94120 -1380
rect 94380 -1400 94620 -1380
rect 94880 -1400 95120 -1380
rect 95380 -1400 95620 -1380
rect 95880 -1400 96120 -1380
rect 96380 -1400 96620 -1380
rect 96880 -1400 97120 -1380
rect 97380 -1400 97620 -1380
rect 97880 -1400 98120 -1380
rect 98380 -1400 98620 -1380
rect 98880 -1400 99120 -1380
rect 99380 -1400 99620 -1380
rect 99880 -1400 100120 -1380
rect 100380 -1400 100620 -1380
rect 100880 -1400 101120 -1380
rect 101380 -1400 101620 -1380
rect 101880 -1400 102120 -1380
rect 102380 -1400 102620 -1380
rect 102880 -1400 103120 -1380
rect 103380 -1400 103620 -1380
rect 103880 -1400 104120 -1380
rect 104380 -1400 104620 -1380
rect 104880 -1400 105120 -1380
rect 105380 -1400 105620 -1380
rect 105880 -1400 106120 -1380
rect 106380 -1400 106620 -1380
rect 106880 -1400 107120 -1380
rect 107380 -1400 107620 -1380
rect 107880 -1400 108120 -1380
rect 108380 -1400 108620 -1380
rect 108880 -1400 109120 -1380
rect 109380 -1400 109620 -1380
rect 109880 -1400 110120 -1380
rect 110380 -1400 110620 -1380
rect 110880 -1400 111120 -1380
rect 111380 -1400 111620 -1380
rect 111880 -1400 112120 -1380
rect 112380 -1400 112620 -1380
rect 112880 -1400 113120 -1380
rect 113380 -1400 113620 -1380
rect 113880 -1400 114120 -1380
rect 114380 -1400 114620 -1380
rect 114880 -1400 115120 -1380
rect 115380 -1400 115620 -1380
rect 115880 -1400 116120 -1380
rect 116380 -1400 116620 -1380
rect 116880 -1400 117120 -1380
rect 117380 -1400 117620 -1380
rect 117880 -1400 118120 -1380
rect 118380 -1400 118620 -1380
rect 118880 -1400 119120 -1380
rect 119380 -1400 119620 -1380
rect 119880 -1400 120120 -1380
rect 120380 -1400 120620 -1380
rect 120880 -1400 121120 -1380
rect 121380 -1400 121620 -1380
rect 121880 -1400 122120 -1380
rect 122380 -1400 122620 -1380
rect 122880 -1400 123120 -1380
rect 123380 -1400 123620 -1380
rect 123880 -1400 124120 -1380
rect 124380 -1400 124620 -1380
rect 124880 -1400 125120 -1380
rect 125380 -1400 125620 -1380
rect 125880 -1400 126120 -1380
rect 126380 -1400 126620 -1380
rect 126880 -1400 127120 -1380
rect 127380 -1400 127620 -1380
rect 127880 -1400 128120 -1380
rect 128380 -1400 128620 -1380
rect 128880 -1400 129120 -1380
rect 129380 -1400 129620 -1380
rect 129880 -1400 130120 -1380
rect 130380 -1400 130620 -1380
rect 130880 -1400 131120 -1380
rect 131380 -1400 131620 -1380
rect 131880 -1400 132120 -1380
rect 132380 -1400 132620 -1380
rect 132880 -1400 133120 -1380
rect 133380 -1400 133620 -1380
rect 133880 -1400 134120 -1380
rect 134380 -1400 134620 -1380
rect 134880 -1400 135120 -1380
rect 135380 -1400 135620 -1380
rect 135880 -1400 136120 -1380
rect 136380 -1400 136620 -1380
rect 136880 -1400 137120 -1380
rect 137380 -1400 137620 -1380
rect 137880 -1400 138120 -1380
rect 138380 -1400 138620 -1380
rect 138880 -1400 139120 -1380
rect 139380 -1400 139620 -1380
rect 139880 -1400 140000 -1380
rect 88000 -1410 140000 -1400
rect 88000 -1480 136150 -1410
rect 136350 -1480 136650 -1410
rect 136850 -1480 137150 -1410
rect 137350 -1480 137650 -1410
rect 137850 -1480 138150 -1410
rect 138350 -1480 138650 -1410
rect 138850 -1480 139150 -1410
rect 139350 -1480 139650 -1410
rect 139850 -1480 140000 -1410
rect 88000 -1520 140000 -1480
rect 88000 -1590 136150 -1520
rect 136350 -1590 136650 -1520
rect 136850 -1590 137150 -1520
rect 137350 -1590 137650 -1520
rect 137850 -1590 138150 -1520
rect 138350 -1590 138650 -1520
rect 138850 -1590 139150 -1520
rect 139350 -1590 139650 -1520
rect 139850 -1590 140000 -1520
rect 88000 -1600 140000 -1590
rect 88000 -1620 88120 -1600
rect 88380 -1620 88620 -1600
rect 88880 -1620 89120 -1600
rect 89380 -1620 89620 -1600
rect 89880 -1620 90120 -1600
rect 90380 -1620 90620 -1600
rect 90880 -1620 91120 -1600
rect 91380 -1620 91620 -1600
rect 91880 -1620 92120 -1600
rect 92380 -1620 92620 -1600
rect 92880 -1620 93120 -1600
rect 93380 -1620 93620 -1600
rect 93880 -1620 94120 -1600
rect 94380 -1620 94620 -1600
rect 94880 -1620 95120 -1600
rect 95380 -1620 95620 -1600
rect 95880 -1620 96120 -1600
rect 96380 -1620 96620 -1600
rect 96880 -1620 97120 -1600
rect 97380 -1620 97620 -1600
rect 97880 -1620 98120 -1600
rect 98380 -1620 98620 -1600
rect 98880 -1620 99120 -1600
rect 99380 -1620 99620 -1600
rect 99880 -1620 100120 -1600
rect 100380 -1620 100620 -1600
rect 100880 -1620 101120 -1600
rect 101380 -1620 101620 -1600
rect 101880 -1620 102120 -1600
rect 102380 -1620 102620 -1600
rect 102880 -1620 103120 -1600
rect 103380 -1620 103620 -1600
rect 103880 -1620 104120 -1600
rect 104380 -1620 104620 -1600
rect 104880 -1620 105120 -1600
rect 105380 -1620 105620 -1600
rect 105880 -1620 106120 -1600
rect 106380 -1620 106620 -1600
rect 106880 -1620 107120 -1600
rect 107380 -1620 107620 -1600
rect 107880 -1620 108120 -1600
rect 108380 -1620 108620 -1600
rect 108880 -1620 109120 -1600
rect 109380 -1620 109620 -1600
rect 109880 -1620 110120 -1600
rect 110380 -1620 110620 -1600
rect 110880 -1620 111120 -1600
rect 111380 -1620 111620 -1600
rect 111880 -1620 112120 -1600
rect 112380 -1620 112620 -1600
rect 112880 -1620 113120 -1600
rect 113380 -1620 113620 -1600
rect 113880 -1620 114120 -1600
rect 114380 -1620 114620 -1600
rect 114880 -1620 115120 -1600
rect 115380 -1620 115620 -1600
rect 115880 -1620 116120 -1600
rect 116380 -1620 116620 -1600
rect 116880 -1620 117120 -1600
rect 117380 -1620 117620 -1600
rect 117880 -1620 118120 -1600
rect 118380 -1620 118620 -1600
rect 118880 -1620 119120 -1600
rect 119380 -1620 119620 -1600
rect 119880 -1620 120120 -1600
rect 120380 -1620 120620 -1600
rect 120880 -1620 121120 -1600
rect 121380 -1620 121620 -1600
rect 121880 -1620 122120 -1600
rect 122380 -1620 122620 -1600
rect 122880 -1620 123120 -1600
rect 123380 -1620 123620 -1600
rect 123880 -1620 124120 -1600
rect 124380 -1620 124620 -1600
rect 124880 -1620 125120 -1600
rect 125380 -1620 125620 -1600
rect 125880 -1620 126120 -1600
rect 126380 -1620 126620 -1600
rect 126880 -1620 127120 -1600
rect 127380 -1620 127620 -1600
rect 127880 -1620 128120 -1600
rect 128380 -1620 128620 -1600
rect 128880 -1620 129120 -1600
rect 129380 -1620 129620 -1600
rect 129880 -1620 130120 -1600
rect 130380 -1620 130620 -1600
rect 130880 -1620 131120 -1600
rect 131380 -1620 131620 -1600
rect 131880 -1620 132120 -1600
rect 132380 -1620 132620 -1600
rect 132880 -1620 133120 -1600
rect 133380 -1620 133620 -1600
rect 133880 -1620 134120 -1600
rect 134380 -1620 134620 -1600
rect 134880 -1620 135120 -1600
rect 135380 -1620 135620 -1600
rect 135880 -1620 136120 -1600
rect 136380 -1620 136620 -1600
rect 136880 -1620 137120 -1600
rect 137380 -1620 137620 -1600
rect 137880 -1620 138120 -1600
rect 138380 -1620 138620 -1600
rect 138880 -1620 139120 -1600
rect 139380 -1620 139620 -1600
rect 139880 -1620 140000 -1600
rect 88000 -1880 88100 -1620
rect 88400 -1880 88600 -1620
rect 88900 -1880 89100 -1620
rect 89400 -1880 89600 -1620
rect 89900 -1880 90100 -1620
rect 90400 -1880 90600 -1620
rect 90900 -1880 91100 -1620
rect 91400 -1880 91600 -1620
rect 91900 -1880 92100 -1620
rect 92400 -1880 92600 -1620
rect 92900 -1880 93100 -1620
rect 93400 -1880 93600 -1620
rect 93900 -1880 94100 -1620
rect 94400 -1880 94600 -1620
rect 94900 -1880 95100 -1620
rect 95400 -1880 95600 -1620
rect 95900 -1880 96100 -1620
rect 96400 -1880 96600 -1620
rect 96900 -1880 97100 -1620
rect 97400 -1880 97600 -1620
rect 97900 -1880 98100 -1620
rect 98400 -1880 98600 -1620
rect 98900 -1880 99100 -1620
rect 99400 -1880 99600 -1620
rect 99900 -1880 100100 -1620
rect 100400 -1880 100600 -1620
rect 100900 -1880 101100 -1620
rect 101400 -1880 101600 -1620
rect 101900 -1880 102100 -1620
rect 102400 -1880 102600 -1620
rect 102900 -1880 103100 -1620
rect 103400 -1880 103600 -1620
rect 103900 -1880 104100 -1620
rect 104400 -1880 104600 -1620
rect 104900 -1880 105100 -1620
rect 105400 -1880 105600 -1620
rect 105900 -1880 106100 -1620
rect 106400 -1880 106600 -1620
rect 106900 -1880 107100 -1620
rect 107400 -1880 107600 -1620
rect 107900 -1880 108100 -1620
rect 108400 -1880 108600 -1620
rect 108900 -1880 109100 -1620
rect 109400 -1880 109600 -1620
rect 109900 -1880 110100 -1620
rect 110400 -1880 110600 -1620
rect 110900 -1880 111100 -1620
rect 111400 -1880 111600 -1620
rect 111900 -1880 112100 -1620
rect 112400 -1880 112600 -1620
rect 112900 -1880 113100 -1620
rect 113400 -1880 113600 -1620
rect 113900 -1880 114100 -1620
rect 114400 -1880 114600 -1620
rect 114900 -1880 115100 -1620
rect 115400 -1880 115600 -1620
rect 115900 -1880 116100 -1620
rect 116400 -1880 116600 -1620
rect 116900 -1880 117100 -1620
rect 117400 -1880 117600 -1620
rect 117900 -1880 118100 -1620
rect 118400 -1880 118600 -1620
rect 118900 -1880 119100 -1620
rect 119400 -1880 119600 -1620
rect 119900 -1880 120100 -1620
rect 120400 -1880 120600 -1620
rect 120900 -1880 121100 -1620
rect 121400 -1880 121600 -1620
rect 121900 -1880 122100 -1620
rect 122400 -1880 122600 -1620
rect 122900 -1880 123100 -1620
rect 123400 -1880 123600 -1620
rect 123900 -1880 124100 -1620
rect 124400 -1880 124600 -1620
rect 124900 -1880 125100 -1620
rect 125400 -1880 125600 -1620
rect 125900 -1880 126100 -1620
rect 126400 -1880 126600 -1620
rect 126900 -1880 127100 -1620
rect 127400 -1880 127600 -1620
rect 127900 -1880 128100 -1620
rect 128400 -1880 128600 -1620
rect 128900 -1880 129100 -1620
rect 129400 -1880 129600 -1620
rect 129900 -1880 130100 -1620
rect 130400 -1880 130600 -1620
rect 130900 -1880 131100 -1620
rect 131400 -1880 131600 -1620
rect 131900 -1880 132100 -1620
rect 132400 -1880 132600 -1620
rect 132900 -1880 133100 -1620
rect 133400 -1880 133600 -1620
rect 133900 -1880 134100 -1620
rect 134400 -1880 134600 -1620
rect 134900 -1880 135100 -1620
rect 135400 -1880 135600 -1620
rect 135900 -1650 136100 -1620
rect 135900 -1850 136020 -1650
rect 136090 -1850 136100 -1650
rect 135900 -1880 136100 -1850
rect 136400 -1650 136600 -1620
rect 136400 -1850 136410 -1650
rect 136480 -1850 136520 -1650
rect 136590 -1850 136600 -1650
rect 136400 -1880 136600 -1850
rect 136900 -1650 137100 -1620
rect 136900 -1850 136910 -1650
rect 136980 -1850 137020 -1650
rect 137090 -1850 137100 -1650
rect 136900 -1880 137100 -1850
rect 137400 -1650 137600 -1620
rect 137400 -1850 137410 -1650
rect 137480 -1850 137520 -1650
rect 137590 -1850 137600 -1650
rect 137400 -1880 137600 -1850
rect 137900 -1650 138100 -1620
rect 137900 -1850 137910 -1650
rect 137980 -1850 138020 -1650
rect 138090 -1850 138100 -1650
rect 137900 -1880 138100 -1850
rect 138400 -1650 138600 -1620
rect 138400 -1850 138410 -1650
rect 138480 -1850 138520 -1650
rect 138590 -1850 138600 -1650
rect 138400 -1880 138600 -1850
rect 138900 -1650 139100 -1620
rect 138900 -1850 138910 -1650
rect 138980 -1850 139020 -1650
rect 139090 -1850 139100 -1650
rect 138900 -1880 139100 -1850
rect 139400 -1650 139600 -1620
rect 139400 -1850 139410 -1650
rect 139480 -1850 139520 -1650
rect 139590 -1850 139600 -1650
rect 139400 -1880 139600 -1850
rect 139900 -1650 140000 -1620
rect 139900 -1850 139910 -1650
rect 139980 -1850 140000 -1650
rect 139900 -1880 140000 -1850
rect 88000 -1900 88120 -1880
rect 88380 -1900 88620 -1880
rect 88880 -1900 89120 -1880
rect 89380 -1900 89620 -1880
rect 89880 -1900 90120 -1880
rect 90380 -1900 90620 -1880
rect 90880 -1900 91120 -1880
rect 91380 -1900 91620 -1880
rect 91880 -1900 92120 -1880
rect 92380 -1900 92620 -1880
rect 92880 -1900 93120 -1880
rect 93380 -1900 93620 -1880
rect 93880 -1900 94120 -1880
rect 94380 -1900 94620 -1880
rect 94880 -1900 95120 -1880
rect 95380 -1900 95620 -1880
rect 95880 -1900 96120 -1880
rect 96380 -1900 96620 -1880
rect 96880 -1900 97120 -1880
rect 97380 -1900 97620 -1880
rect 97880 -1900 98120 -1880
rect 98380 -1900 98620 -1880
rect 98880 -1900 99120 -1880
rect 99380 -1900 99620 -1880
rect 99880 -1900 100120 -1880
rect 100380 -1900 100620 -1880
rect 100880 -1900 101120 -1880
rect 101380 -1900 101620 -1880
rect 101880 -1900 102120 -1880
rect 102380 -1900 102620 -1880
rect 102880 -1900 103120 -1880
rect 103380 -1900 103620 -1880
rect 103880 -1900 104120 -1880
rect 104380 -1900 104620 -1880
rect 104880 -1900 105120 -1880
rect 105380 -1900 105620 -1880
rect 105880 -1900 106120 -1880
rect 106380 -1900 106620 -1880
rect 106880 -1900 107120 -1880
rect 107380 -1900 107620 -1880
rect 107880 -1900 108120 -1880
rect 108380 -1900 108620 -1880
rect 108880 -1900 109120 -1880
rect 109380 -1900 109620 -1880
rect 109880 -1900 110120 -1880
rect 110380 -1900 110620 -1880
rect 110880 -1900 111120 -1880
rect 111380 -1900 111620 -1880
rect 111880 -1900 112120 -1880
rect 112380 -1900 112620 -1880
rect 112880 -1900 113120 -1880
rect 113380 -1900 113620 -1880
rect 113880 -1900 114120 -1880
rect 114380 -1900 114620 -1880
rect 114880 -1900 115120 -1880
rect 115380 -1900 115620 -1880
rect 115880 -1900 116120 -1880
rect 116380 -1900 116620 -1880
rect 116880 -1900 117120 -1880
rect 117380 -1900 117620 -1880
rect 117880 -1900 118120 -1880
rect 118380 -1900 118620 -1880
rect 118880 -1900 119120 -1880
rect 119380 -1900 119620 -1880
rect 119880 -1900 120120 -1880
rect 120380 -1900 120620 -1880
rect 120880 -1900 121120 -1880
rect 121380 -1900 121620 -1880
rect 121880 -1900 122120 -1880
rect 122380 -1900 122620 -1880
rect 122880 -1900 123120 -1880
rect 123380 -1900 123620 -1880
rect 123880 -1900 124120 -1880
rect 124380 -1900 124620 -1880
rect 124880 -1900 125120 -1880
rect 125380 -1900 125620 -1880
rect 125880 -1900 126120 -1880
rect 126380 -1900 126620 -1880
rect 126880 -1900 127120 -1880
rect 127380 -1900 127620 -1880
rect 127880 -1900 128120 -1880
rect 128380 -1900 128620 -1880
rect 128880 -1900 129120 -1880
rect 129380 -1900 129620 -1880
rect 129880 -1900 130120 -1880
rect 130380 -1900 130620 -1880
rect 130880 -1900 131120 -1880
rect 131380 -1900 131620 -1880
rect 131880 -1900 132120 -1880
rect 132380 -1900 132620 -1880
rect 132880 -1900 133120 -1880
rect 133380 -1900 133620 -1880
rect 133880 -1900 134120 -1880
rect 134380 -1900 134620 -1880
rect 134880 -1900 135120 -1880
rect 135380 -1900 135620 -1880
rect 135880 -1900 136120 -1880
rect 136380 -1900 136620 -1880
rect 136880 -1900 137120 -1880
rect 137380 -1900 137620 -1880
rect 137880 -1900 138120 -1880
rect 138380 -1900 138620 -1880
rect 138880 -1900 139120 -1880
rect 139380 -1900 139620 -1880
rect 139880 -1900 140000 -1880
rect 88000 -1910 140000 -1900
rect 88000 -1980 136150 -1910
rect 136350 -1980 136650 -1910
rect 136850 -1980 137150 -1910
rect 137350 -1980 137650 -1910
rect 137850 -1980 138150 -1910
rect 138350 -1980 138650 -1910
rect 138850 -1980 139150 -1910
rect 139350 -1980 139650 -1910
rect 139850 -1980 140000 -1910
rect 12000 -2100 20000 -2000
rect 12000 -2120 12120 -2100
rect 12380 -2120 12620 -2100
rect 12880 -2120 13120 -2100
rect 13380 -2120 13620 -2100
rect 13880 -2120 14120 -2100
rect 14380 -2120 14620 -2100
rect 14880 -2120 15120 -2100
rect 15380 -2120 15620 -2100
rect 15880 -2120 16120 -2100
rect 16380 -2120 16620 -2100
rect 16880 -2120 17120 -2100
rect 17380 -2120 17620 -2100
rect 17880 -2120 18120 -2100
rect 18380 -2120 18620 -2100
rect 18880 -2120 19120 -2100
rect 19380 -2120 19620 -2100
rect 19880 -2120 20000 -2100
rect 12000 -2380 12100 -2120
rect 12400 -2380 12600 -2120
rect 12900 -2380 13100 -2120
rect 13400 -2380 13600 -2120
rect 13900 -2380 14100 -2120
rect 14400 -2380 14600 -2120
rect 14900 -2380 15100 -2120
rect 15400 -2380 15600 -2120
rect 15900 -2380 16100 -2120
rect 16400 -2380 16600 -2120
rect 16900 -2380 17100 -2120
rect 17400 -2380 17600 -2120
rect 17900 -2380 18100 -2120
rect 18400 -2380 18600 -2120
rect 18900 -2380 19100 -2120
rect 19400 -2380 19600 -2120
rect 19900 -2380 20000 -2120
rect 12000 -2400 12120 -2380
rect 12380 -2400 12620 -2380
rect 12880 -2400 13120 -2380
rect 13380 -2400 13620 -2380
rect 13880 -2400 14120 -2380
rect 14380 -2400 14620 -2380
rect 14880 -2400 15120 -2380
rect 15380 -2400 15620 -2380
rect 15880 -2400 16120 -2380
rect 16380 -2400 16620 -2380
rect 16880 -2400 17120 -2380
rect 17380 -2400 17620 -2380
rect 17880 -2400 18120 -2380
rect 18380 -2400 18620 -2380
rect 18880 -2400 19120 -2380
rect 19380 -2400 19620 -2380
rect 19880 -2400 20000 -2380
rect 12000 -2600 20000 -2400
rect 12000 -2620 12120 -2600
rect 12380 -2620 12620 -2600
rect 12880 -2620 13120 -2600
rect 13380 -2620 13620 -2600
rect 13880 -2620 14120 -2600
rect 14380 -2620 14620 -2600
rect 14880 -2620 15120 -2600
rect 15380 -2620 15620 -2600
rect 15880 -2620 16120 -2600
rect 16380 -2620 16620 -2600
rect 16880 -2620 17120 -2600
rect 17380 -2620 17620 -2600
rect 17880 -2620 18120 -2600
rect 18380 -2620 18620 -2600
rect 18880 -2620 19120 -2600
rect 19380 -2620 19620 -2600
rect 19880 -2620 20000 -2600
rect 12000 -2880 12100 -2620
rect 12400 -2880 12600 -2620
rect 12900 -2880 13100 -2620
rect 13400 -2880 13600 -2620
rect 13900 -2880 14100 -2620
rect 14400 -2880 14600 -2620
rect 14900 -2880 15100 -2620
rect 15400 -2880 15600 -2620
rect 15900 -2880 16100 -2620
rect 16400 -2880 16600 -2620
rect 16900 -2880 17100 -2620
rect 17400 -2880 17600 -2620
rect 17900 -2880 18100 -2620
rect 18400 -2880 18600 -2620
rect 18900 -2880 19100 -2620
rect 19400 -2880 19600 -2620
rect 19900 -2880 20000 -2620
rect 12000 -2900 12120 -2880
rect 12380 -2900 12620 -2880
rect 12880 -2900 13120 -2880
rect 13380 -2900 13620 -2880
rect 13880 -2900 14120 -2880
rect 14380 -2900 14620 -2880
rect 14880 -2900 15120 -2880
rect 15380 -2900 15620 -2880
rect 15880 -2900 16120 -2880
rect 16380 -2900 16620 -2880
rect 16880 -2900 17120 -2880
rect 17380 -2900 17620 -2880
rect 17880 -2900 18120 -2880
rect 18380 -2900 18620 -2880
rect 18880 -2900 19120 -2880
rect 19380 -2900 19620 -2880
rect 19880 -2900 20000 -2880
rect 12000 -3100 20000 -2900
rect 12000 -3120 12120 -3100
rect 12380 -3120 12620 -3100
rect 12880 -3120 13120 -3100
rect 13380 -3120 13620 -3100
rect 13880 -3120 14120 -3100
rect 14380 -3120 14620 -3100
rect 14880 -3120 15120 -3100
rect 15380 -3120 15620 -3100
rect 15880 -3120 16120 -3100
rect 16380 -3120 16620 -3100
rect 16880 -3120 17120 -3100
rect 17380 -3120 17620 -3100
rect 17880 -3120 18120 -3100
rect 18380 -3120 18620 -3100
rect 18880 -3120 19120 -3100
rect 19380 -3120 19620 -3100
rect 19880 -3120 20000 -3100
rect 12000 -3380 12100 -3120
rect 12400 -3380 12600 -3120
rect 12900 -3380 13100 -3120
rect 13400 -3380 13600 -3120
rect 13900 -3380 14100 -3120
rect 14400 -3380 14600 -3120
rect 14900 -3380 15100 -3120
rect 15400 -3380 15600 -3120
rect 15900 -3380 16100 -3120
rect 16400 -3380 16600 -3120
rect 16900 -3380 17100 -3120
rect 17400 -3380 17600 -3120
rect 17900 -3380 18100 -3120
rect 18400 -3380 18600 -3120
rect 18900 -3380 19100 -3120
rect 19400 -3380 19600 -3120
rect 19900 -3380 20000 -3120
rect 12000 -3400 12120 -3380
rect 12380 -3400 12620 -3380
rect 12880 -3400 13120 -3380
rect 13380 -3400 13620 -3380
rect 13880 -3400 14120 -3380
rect 14380 -3400 14620 -3380
rect 14880 -3400 15120 -3380
rect 15380 -3400 15620 -3380
rect 15880 -3400 16120 -3380
rect 16380 -3400 16620 -3380
rect 16880 -3400 17120 -3380
rect 17380 -3400 17620 -3380
rect 17880 -3400 18120 -3380
rect 18380 -3400 18620 -3380
rect 18880 -3400 19120 -3380
rect 19380 -3400 19620 -3380
rect 19880 -3400 20000 -3380
rect 12000 -3600 20000 -3400
rect 12000 -3620 12120 -3600
rect 12380 -3620 12620 -3600
rect 12880 -3620 13120 -3600
rect 13380 -3620 13620 -3600
rect 13880 -3620 14120 -3600
rect 14380 -3620 14620 -3600
rect 14880 -3620 15120 -3600
rect 15380 -3620 15620 -3600
rect 15880 -3620 16120 -3600
rect 16380 -3620 16620 -3600
rect 16880 -3620 17120 -3600
rect 17380 -3620 17620 -3600
rect 17880 -3620 18120 -3600
rect 18380 -3620 18620 -3600
rect 18880 -3620 19120 -3600
rect 19380 -3620 19620 -3600
rect 19880 -3620 20000 -3600
rect 12000 -3880 12100 -3620
rect 12400 -3880 12600 -3620
rect 12900 -3880 13100 -3620
rect 13400 -3880 13600 -3620
rect 13900 -3880 14100 -3620
rect 14400 -3880 14600 -3620
rect 14900 -3880 15100 -3620
rect 15400 -3880 15600 -3620
rect 15900 -3880 16100 -3620
rect 16400 -3880 16600 -3620
rect 16900 -3880 17100 -3620
rect 17400 -3880 17600 -3620
rect 17900 -3880 18100 -3620
rect 18400 -3880 18600 -3620
rect 18900 -3880 19100 -3620
rect 19400 -3880 19600 -3620
rect 19900 -3880 20000 -3620
rect 12000 -3900 12120 -3880
rect 12380 -3900 12620 -3880
rect 12880 -3900 13120 -3880
rect 13380 -3900 13620 -3880
rect 13880 -3900 14120 -3880
rect 14380 -3900 14620 -3880
rect 14880 -3900 15120 -3880
rect 15380 -3900 15620 -3880
rect 15880 -3900 16120 -3880
rect 16380 -3900 16620 -3880
rect 16880 -3900 17120 -3880
rect 17380 -3900 17620 -3880
rect 17880 -3900 18120 -3880
rect 18380 -3900 18620 -3880
rect 18880 -3900 19120 -3880
rect 19380 -3900 19620 -3880
rect 19880 -3900 20000 -3880
rect 12000 -4100 20000 -3900
rect 12000 -4120 12120 -4100
rect 12380 -4120 12620 -4100
rect 12880 -4120 13120 -4100
rect 13380 -4120 13620 -4100
rect 13880 -4120 14120 -4100
rect 14380 -4120 14620 -4100
rect 14880 -4120 15120 -4100
rect 15380 -4120 15620 -4100
rect 15880 -4120 16120 -4100
rect 16380 -4120 16620 -4100
rect 16880 -4120 17120 -4100
rect 17380 -4120 17620 -4100
rect 17880 -4120 18120 -4100
rect 18380 -4120 18620 -4100
rect 18880 -4120 19120 -4100
rect 19380 -4120 19620 -4100
rect 19880 -4120 20000 -4100
rect 12000 -4380 12100 -4120
rect 12400 -4380 12600 -4120
rect 12900 -4380 13100 -4120
rect 13400 -4380 13600 -4120
rect 13900 -4380 14100 -4120
rect 14400 -4380 14600 -4120
rect 14900 -4380 15100 -4120
rect 15400 -4380 15600 -4120
rect 15900 -4380 16100 -4120
rect 16400 -4380 16600 -4120
rect 16900 -4380 17100 -4120
rect 17400 -4380 17600 -4120
rect 17900 -4380 18100 -4120
rect 18400 -4380 18600 -4120
rect 18900 -4380 19100 -4120
rect 19400 -4380 19600 -4120
rect 19900 -4380 20000 -4120
rect 12000 -4400 12120 -4380
rect 12380 -4400 12620 -4380
rect 12880 -4400 13120 -4380
rect 13380 -4400 13620 -4380
rect 13880 -4400 14120 -4380
rect 14380 -4400 14620 -4380
rect 14880 -4400 15120 -4380
rect 15380 -4400 15620 -4380
rect 15880 -4400 16120 -4380
rect 16380 -4400 16620 -4380
rect 16880 -4400 17120 -4380
rect 17380 -4400 17620 -4380
rect 17880 -4400 18120 -4380
rect 18380 -4400 18620 -4380
rect 18880 -4400 19120 -4380
rect 19380 -4400 19620 -4380
rect 19880 -4400 20000 -4380
rect 12000 -4600 20000 -4400
rect 12000 -4620 12120 -4600
rect 12380 -4620 12620 -4600
rect 12880 -4620 13120 -4600
rect 13380 -4620 13620 -4600
rect 13880 -4620 14120 -4600
rect 14380 -4620 14620 -4600
rect 14880 -4620 15120 -4600
rect 15380 -4620 15620 -4600
rect 15880 -4620 16120 -4600
rect 16380 -4620 16620 -4600
rect 16880 -4620 17120 -4600
rect 17380 -4620 17620 -4600
rect 17880 -4620 18120 -4600
rect 18380 -4620 18620 -4600
rect 18880 -4620 19120 -4600
rect 19380 -4620 19620 -4600
rect 19880 -4620 20000 -4600
rect 12000 -4880 12100 -4620
rect 12400 -4880 12600 -4620
rect 12900 -4880 13100 -4620
rect 13400 -4880 13600 -4620
rect 13900 -4880 14100 -4620
rect 14400 -4880 14600 -4620
rect 14900 -4880 15100 -4620
rect 15400 -4880 15600 -4620
rect 15900 -4880 16100 -4620
rect 16400 -4880 16600 -4620
rect 16900 -4880 17100 -4620
rect 17400 -4880 17600 -4620
rect 17900 -4880 18100 -4620
rect 18400 -4880 18600 -4620
rect 18900 -4880 19100 -4620
rect 19400 -4880 19600 -4620
rect 19900 -4880 20000 -4620
rect 12000 -4900 12120 -4880
rect 12380 -4900 12620 -4880
rect 12880 -4900 13120 -4880
rect 13380 -4900 13620 -4880
rect 13880 -4900 14120 -4880
rect 14380 -4900 14620 -4880
rect 14880 -4900 15120 -4880
rect 15380 -4900 15620 -4880
rect 15880 -4900 16120 -4880
rect 16380 -4900 16620 -4880
rect 16880 -4900 17120 -4880
rect 17380 -4900 17620 -4880
rect 17880 -4900 18120 -4880
rect 18380 -4900 18620 -4880
rect 18880 -4900 19120 -4880
rect 19380 -4900 19620 -4880
rect 19880 -4900 20000 -4880
rect 12000 -5100 20000 -4900
rect 12000 -5120 12120 -5100
rect 12380 -5120 12620 -5100
rect 12880 -5120 13120 -5100
rect 13380 -5120 13620 -5100
rect 13880 -5120 14120 -5100
rect 14380 -5120 14620 -5100
rect 14880 -5120 15120 -5100
rect 15380 -5120 15620 -5100
rect 15880 -5120 16120 -5100
rect 16380 -5120 16620 -5100
rect 16880 -5120 17120 -5100
rect 17380 -5120 17620 -5100
rect 17880 -5120 18120 -5100
rect 18380 -5120 18620 -5100
rect 18880 -5120 19120 -5100
rect 19380 -5120 19620 -5100
rect 19880 -5120 20000 -5100
rect 12000 -5380 12100 -5120
rect 12400 -5380 12600 -5120
rect 12900 -5380 13100 -5120
rect 13400 -5380 13600 -5120
rect 13900 -5380 14100 -5120
rect 14400 -5380 14600 -5120
rect 14900 -5380 15100 -5120
rect 15400 -5380 15600 -5120
rect 15900 -5380 16100 -5120
rect 16400 -5380 16600 -5120
rect 16900 -5380 17100 -5120
rect 17400 -5380 17600 -5120
rect 17900 -5380 18100 -5120
rect 18400 -5380 18600 -5120
rect 18900 -5380 19100 -5120
rect 19400 -5380 19600 -5120
rect 19900 -5380 20000 -5120
rect 12000 -5400 12120 -5380
rect 12380 -5400 12620 -5380
rect 12880 -5400 13120 -5380
rect 13380 -5400 13620 -5380
rect 13880 -5400 14120 -5380
rect 14380 -5400 14620 -5380
rect 14880 -5400 15120 -5380
rect 15380 -5400 15620 -5380
rect 15880 -5400 16120 -5380
rect 16380 -5400 16620 -5380
rect 16880 -5400 17120 -5380
rect 17380 -5400 17620 -5380
rect 17880 -5400 18120 -5380
rect 18380 -5400 18620 -5380
rect 18880 -5400 19120 -5380
rect 19380 -5400 19620 -5380
rect 19880 -5400 20000 -5380
rect 12000 -5600 20000 -5400
rect 12000 -5620 12120 -5600
rect 12380 -5620 12620 -5600
rect 12880 -5620 13120 -5600
rect 13380 -5620 13620 -5600
rect 13880 -5620 14120 -5600
rect 14380 -5620 14620 -5600
rect 14880 -5620 15120 -5600
rect 15380 -5620 15620 -5600
rect 15880 -5620 16120 -5600
rect 16380 -5620 16620 -5600
rect 16880 -5620 17120 -5600
rect 17380 -5620 17620 -5600
rect 17880 -5620 18120 -5600
rect 18380 -5620 18620 -5600
rect 18880 -5620 19120 -5600
rect 19380 -5620 19620 -5600
rect 19880 -5620 20000 -5600
rect 12000 -5880 12100 -5620
rect 12400 -5880 12600 -5620
rect 12900 -5880 13100 -5620
rect 13400 -5880 13600 -5620
rect 13900 -5880 14100 -5620
rect 14400 -5880 14600 -5620
rect 14900 -5880 15100 -5620
rect 15400 -5880 15600 -5620
rect 15900 -5880 16100 -5620
rect 16400 -5880 16600 -5620
rect 16900 -5880 17100 -5620
rect 17400 -5880 17600 -5620
rect 17900 -5880 18100 -5620
rect 18400 -5880 18600 -5620
rect 18900 -5880 19100 -5620
rect 19400 -5880 19600 -5620
rect 19900 -5880 20000 -5620
rect 12000 -5900 12120 -5880
rect 12380 -5900 12620 -5880
rect 12880 -5900 13120 -5880
rect 13380 -5900 13620 -5880
rect 13880 -5900 14120 -5880
rect 14380 -5900 14620 -5880
rect 14880 -5900 15120 -5880
rect 15380 -5900 15620 -5880
rect 15880 -5900 16120 -5880
rect 16380 -5900 16620 -5880
rect 16880 -5900 17120 -5880
rect 17380 -5900 17620 -5880
rect 17880 -5900 18120 -5880
rect 18380 -5900 18620 -5880
rect 18880 -5900 19120 -5880
rect 19380 -5900 19620 -5880
rect 19880 -5900 20000 -5880
rect 12000 -6100 20000 -5900
rect 12000 -6120 12120 -6100
rect 12380 -6120 12620 -6100
rect 12880 -6120 13120 -6100
rect 13380 -6120 13620 -6100
rect 13880 -6120 14120 -6100
rect 14380 -6120 14620 -6100
rect 14880 -6120 15120 -6100
rect 15380 -6120 15620 -6100
rect 15880 -6120 16120 -6100
rect 16380 -6120 16620 -6100
rect 16880 -6120 17120 -6100
rect 17380 -6120 17620 -6100
rect 17880 -6120 18120 -6100
rect 18380 -6120 18620 -6100
rect 18880 -6120 19120 -6100
rect 19380 -6120 19620 -6100
rect 19880 -6120 20000 -6100
rect 12000 -6380 12100 -6120
rect 12400 -6380 12600 -6120
rect 12900 -6380 13100 -6120
rect 13400 -6380 13600 -6120
rect 13900 -6380 14100 -6120
rect 14400 -6380 14600 -6120
rect 14900 -6380 15100 -6120
rect 15400 -6380 15600 -6120
rect 15900 -6380 16100 -6120
rect 16400 -6380 16600 -6120
rect 16900 -6380 17100 -6120
rect 17400 -6380 17600 -6120
rect 17900 -6380 18100 -6120
rect 18400 -6380 18600 -6120
rect 18900 -6380 19100 -6120
rect 19400 -6380 19600 -6120
rect 19900 -6380 20000 -6120
rect 12000 -6400 12120 -6380
rect 12380 -6400 12620 -6380
rect 12880 -6400 13120 -6380
rect 13380 -6400 13620 -6380
rect 13880 -6400 14120 -6380
rect 14380 -6400 14620 -6380
rect 14880 -6400 15120 -6380
rect 15380 -6400 15620 -6380
rect 15880 -6400 16120 -6380
rect 16380 -6400 16620 -6380
rect 16880 -6400 17120 -6380
rect 17380 -6400 17620 -6380
rect 17880 -6400 18120 -6380
rect 18380 -6400 18620 -6380
rect 18880 -6400 19120 -6380
rect 19380 -6400 19620 -6380
rect 19880 -6400 20000 -6380
rect 12000 -6600 20000 -6400
rect 12000 -6620 12120 -6600
rect 12380 -6620 12620 -6600
rect 12880 -6620 13120 -6600
rect 13380 -6620 13620 -6600
rect 13880 -6620 14120 -6600
rect 14380 -6620 14620 -6600
rect 14880 -6620 15120 -6600
rect 15380 -6620 15620 -6600
rect 15880 -6620 16120 -6600
rect 16380 -6620 16620 -6600
rect 16880 -6620 17120 -6600
rect 17380 -6620 17620 -6600
rect 17880 -6620 18120 -6600
rect 18380 -6620 18620 -6600
rect 18880 -6620 19120 -6600
rect 19380 -6620 19620 -6600
rect 19880 -6620 20000 -6600
rect 12000 -6880 12100 -6620
rect 12400 -6880 12600 -6620
rect 12900 -6880 13100 -6620
rect 13400 -6880 13600 -6620
rect 13900 -6880 14100 -6620
rect 14400 -6880 14600 -6620
rect 14900 -6880 15100 -6620
rect 15400 -6880 15600 -6620
rect 15900 -6880 16100 -6620
rect 16400 -6880 16600 -6620
rect 16900 -6880 17100 -6620
rect 17400 -6880 17600 -6620
rect 17900 -6880 18100 -6620
rect 18400 -6880 18600 -6620
rect 18900 -6880 19100 -6620
rect 19400 -6880 19600 -6620
rect 19900 -6880 20000 -6620
rect 12000 -6900 12120 -6880
rect 12380 -6900 12620 -6880
rect 12880 -6900 13120 -6880
rect 13380 -6900 13620 -6880
rect 13880 -6900 14120 -6880
rect 14380 -6900 14620 -6880
rect 14880 -6900 15120 -6880
rect 15380 -6900 15620 -6880
rect 15880 -6900 16120 -6880
rect 16380 -6900 16620 -6880
rect 16880 -6900 17120 -6880
rect 17380 -6900 17620 -6880
rect 17880 -6900 18120 -6880
rect 18380 -6900 18620 -6880
rect 18880 -6900 19120 -6880
rect 19380 -6900 19620 -6880
rect 19880 -6900 20000 -6880
rect 12000 -7100 20000 -6900
rect 12000 -7120 12120 -7100
rect 12380 -7120 12620 -7100
rect 12880 -7120 13120 -7100
rect 13380 -7120 13620 -7100
rect 13880 -7120 14120 -7100
rect 14380 -7120 14620 -7100
rect 14880 -7120 15120 -7100
rect 15380 -7120 15620 -7100
rect 15880 -7120 16120 -7100
rect 16380 -7120 16620 -7100
rect 16880 -7120 17120 -7100
rect 17380 -7120 17620 -7100
rect 17880 -7120 18120 -7100
rect 18380 -7120 18620 -7100
rect 18880 -7120 19120 -7100
rect 19380 -7120 19620 -7100
rect 19880 -7120 20000 -7100
rect 12000 -7380 12100 -7120
rect 12400 -7380 12600 -7120
rect 12900 -7380 13100 -7120
rect 13400 -7380 13600 -7120
rect 13900 -7380 14100 -7120
rect 14400 -7380 14600 -7120
rect 14900 -7380 15100 -7120
rect 15400 -7380 15600 -7120
rect 15900 -7380 16100 -7120
rect 16400 -7380 16600 -7120
rect 16900 -7380 17100 -7120
rect 17400 -7380 17600 -7120
rect 17900 -7380 18100 -7120
rect 18400 -7380 18600 -7120
rect 18900 -7380 19100 -7120
rect 19400 -7380 19600 -7120
rect 19900 -7380 20000 -7120
rect 12000 -7400 12120 -7380
rect 12380 -7400 12620 -7380
rect 12880 -7400 13120 -7380
rect 13380 -7400 13620 -7380
rect 13880 -7400 14120 -7380
rect 14380 -7400 14620 -7380
rect 14880 -7400 15120 -7380
rect 15380 -7400 15620 -7380
rect 15880 -7400 16120 -7380
rect 16380 -7400 16620 -7380
rect 16880 -7400 17120 -7380
rect 17380 -7400 17620 -7380
rect 17880 -7400 18120 -7380
rect 18380 -7400 18620 -7380
rect 18880 -7400 19120 -7380
rect 19380 -7400 19620 -7380
rect 19880 -7400 20000 -7380
rect 12000 -7600 20000 -7400
rect 12000 -7620 12120 -7600
rect 12380 -7620 12620 -7600
rect 12880 -7620 13120 -7600
rect 13380 -7620 13620 -7600
rect 13880 -7620 14120 -7600
rect 14380 -7620 14620 -7600
rect 14880 -7620 15120 -7600
rect 15380 -7620 15620 -7600
rect 15880 -7620 16120 -7600
rect 16380 -7620 16620 -7600
rect 16880 -7620 17120 -7600
rect 17380 -7620 17620 -7600
rect 17880 -7620 18120 -7600
rect 18380 -7620 18620 -7600
rect 18880 -7620 19120 -7600
rect 19380 -7620 19620 -7600
rect 19880 -7620 20000 -7600
rect 12000 -7880 12100 -7620
rect 12400 -7880 12600 -7620
rect 12900 -7880 13100 -7620
rect 13400 -7880 13600 -7620
rect 13900 -7880 14100 -7620
rect 14400 -7880 14600 -7620
rect 14900 -7880 15100 -7620
rect 15400 -7880 15600 -7620
rect 15900 -7880 16100 -7620
rect 16400 -7880 16600 -7620
rect 16900 -7880 17100 -7620
rect 17400 -7880 17600 -7620
rect 17900 -7880 18100 -7620
rect 18400 -7880 18600 -7620
rect 18900 -7880 19100 -7620
rect 19400 -7880 19600 -7620
rect 19900 -7880 20000 -7620
rect 12000 -7900 12120 -7880
rect 12380 -7900 12620 -7880
rect 12880 -7900 13120 -7880
rect 13380 -7900 13620 -7880
rect 13880 -7900 14120 -7880
rect 14380 -7900 14620 -7880
rect 14880 -7900 15120 -7880
rect 15380 -7900 15620 -7880
rect 15880 -7900 16120 -7880
rect 16380 -7900 16620 -7880
rect 16880 -7900 17120 -7880
rect 17380 -7900 17620 -7880
rect 17880 -7900 18120 -7880
rect 18380 -7900 18620 -7880
rect 18880 -7900 19120 -7880
rect 19380 -7900 19620 -7880
rect 19880 -7900 20000 -7880
rect 12000 -8100 20000 -7900
rect 12000 -8120 12120 -8100
rect 12380 -8120 12620 -8100
rect 12880 -8120 13120 -8100
rect 13380 -8120 13620 -8100
rect 13880 -8120 14120 -8100
rect 14380 -8120 14620 -8100
rect 14880 -8120 15120 -8100
rect 15380 -8120 15620 -8100
rect 15880 -8120 16120 -8100
rect 16380 -8120 16620 -8100
rect 16880 -8120 17120 -8100
rect 17380 -8120 17620 -8100
rect 17880 -8120 18120 -8100
rect 18380 -8120 18620 -8100
rect 18880 -8120 19120 -8100
rect 19380 -8120 19620 -8100
rect 19880 -8120 20000 -8100
rect 12000 -8380 12100 -8120
rect 12400 -8380 12600 -8120
rect 12900 -8380 13100 -8120
rect 13400 -8380 13600 -8120
rect 13900 -8380 14100 -8120
rect 14400 -8380 14600 -8120
rect 14900 -8380 15100 -8120
rect 15400 -8380 15600 -8120
rect 15900 -8380 16100 -8120
rect 16400 -8380 16600 -8120
rect 16900 -8380 17100 -8120
rect 17400 -8380 17600 -8120
rect 17900 -8380 18100 -8120
rect 18400 -8380 18600 -8120
rect 18900 -8380 19100 -8120
rect 19400 -8380 19600 -8120
rect 19900 -8380 20000 -8120
rect 12000 -8400 12120 -8380
rect 12380 -8400 12620 -8380
rect 12880 -8400 13120 -8380
rect 13380 -8400 13620 -8380
rect 13880 -8400 14120 -8380
rect 14380 -8400 14620 -8380
rect 14880 -8400 15120 -8380
rect 15380 -8400 15620 -8380
rect 15880 -8400 16120 -8380
rect 16380 -8400 16620 -8380
rect 16880 -8400 17120 -8380
rect 17380 -8400 17620 -8380
rect 17880 -8400 18120 -8380
rect 18380 -8400 18620 -8380
rect 18880 -8400 19120 -8380
rect 19380 -8400 19620 -8380
rect 19880 -8400 20000 -8380
rect 12000 -8600 20000 -8400
rect 12000 -8620 12120 -8600
rect 12380 -8620 12620 -8600
rect 12880 -8620 13120 -8600
rect 13380 -8620 13620 -8600
rect 13880 -8620 14120 -8600
rect 14380 -8620 14620 -8600
rect 14880 -8620 15120 -8600
rect 15380 -8620 15620 -8600
rect 15880 -8620 16120 -8600
rect 16380 -8620 16620 -8600
rect 16880 -8620 17120 -8600
rect 17380 -8620 17620 -8600
rect 17880 -8620 18120 -8600
rect 18380 -8620 18620 -8600
rect 18880 -8620 19120 -8600
rect 19380 -8620 19620 -8600
rect 19880 -8620 20000 -8600
rect 12000 -8880 12100 -8620
rect 12400 -8880 12600 -8620
rect 12900 -8880 13100 -8620
rect 13400 -8880 13600 -8620
rect 13900 -8880 14100 -8620
rect 14400 -8880 14600 -8620
rect 14900 -8880 15100 -8620
rect 15400 -8880 15600 -8620
rect 15900 -8880 16100 -8620
rect 16400 -8880 16600 -8620
rect 16900 -8880 17100 -8620
rect 17400 -8880 17600 -8620
rect 17900 -8880 18100 -8620
rect 18400 -8880 18600 -8620
rect 18900 -8880 19100 -8620
rect 19400 -8880 19600 -8620
rect 19900 -8880 20000 -8620
rect 12000 -8900 12120 -8880
rect 12380 -8900 12620 -8880
rect 12880 -8900 13120 -8880
rect 13380 -8900 13620 -8880
rect 13880 -8900 14120 -8880
rect 14380 -8900 14620 -8880
rect 14880 -8900 15120 -8880
rect 15380 -8900 15620 -8880
rect 15880 -8900 16120 -8880
rect 16380 -8900 16620 -8880
rect 16880 -8900 17120 -8880
rect 17380 -8900 17620 -8880
rect 17880 -8900 18120 -8880
rect 18380 -8900 18620 -8880
rect 18880 -8900 19120 -8880
rect 19380 -8900 19620 -8880
rect 19880 -8900 20000 -8880
rect 12000 -9100 20000 -8900
rect 12000 -9120 12120 -9100
rect 12380 -9120 12620 -9100
rect 12880 -9120 13120 -9100
rect 13380 -9120 13620 -9100
rect 13880 -9120 14120 -9100
rect 14380 -9120 14620 -9100
rect 14880 -9120 15120 -9100
rect 15380 -9120 15620 -9100
rect 15880 -9120 16120 -9100
rect 16380 -9120 16620 -9100
rect 16880 -9120 17120 -9100
rect 17380 -9120 17620 -9100
rect 17880 -9120 18120 -9100
rect 18380 -9120 18620 -9100
rect 18880 -9120 19120 -9100
rect 19380 -9120 19620 -9100
rect 19880 -9120 20000 -9100
rect 12000 -9380 12100 -9120
rect 12400 -9380 12600 -9120
rect 12900 -9380 13100 -9120
rect 13400 -9380 13600 -9120
rect 13900 -9380 14100 -9120
rect 14400 -9380 14600 -9120
rect 14900 -9380 15100 -9120
rect 15400 -9380 15600 -9120
rect 15900 -9380 16100 -9120
rect 16400 -9380 16600 -9120
rect 16900 -9380 17100 -9120
rect 17400 -9380 17600 -9120
rect 17900 -9380 18100 -9120
rect 18400 -9380 18600 -9120
rect 18900 -9380 19100 -9120
rect 19400 -9380 19600 -9120
rect 19900 -9380 20000 -9120
rect 12000 -9400 12120 -9380
rect 12380 -9400 12620 -9380
rect 12880 -9400 13120 -9380
rect 13380 -9400 13620 -9380
rect 13880 -9400 14120 -9380
rect 14380 -9400 14620 -9380
rect 14880 -9400 15120 -9380
rect 15380 -9400 15620 -9380
rect 15880 -9400 16120 -9380
rect 16380 -9400 16620 -9380
rect 16880 -9400 17120 -9380
rect 17380 -9400 17620 -9380
rect 17880 -9400 18120 -9380
rect 18380 -9400 18620 -9380
rect 18880 -9400 19120 -9380
rect 19380 -9400 19620 -9380
rect 19880 -9400 20000 -9380
rect 12000 -9600 20000 -9400
rect 12000 -9620 12120 -9600
rect 12380 -9620 12620 -9600
rect 12880 -9620 13120 -9600
rect 13380 -9620 13620 -9600
rect 13880 -9620 14120 -9600
rect 14380 -9620 14620 -9600
rect 14880 -9620 15120 -9600
rect 15380 -9620 15620 -9600
rect 15880 -9620 16120 -9600
rect 16380 -9620 16620 -9600
rect 16880 -9620 17120 -9600
rect 17380 -9620 17620 -9600
rect 17880 -9620 18120 -9600
rect 18380 -9620 18620 -9600
rect 18880 -9620 19120 -9600
rect 19380 -9620 19620 -9600
rect 19880 -9620 20000 -9600
rect 12000 -9880 12100 -9620
rect 12400 -9880 12600 -9620
rect 12900 -9880 13100 -9620
rect 13400 -9880 13600 -9620
rect 13900 -9880 14100 -9620
rect 14400 -9880 14600 -9620
rect 14900 -9880 15100 -9620
rect 15400 -9880 15600 -9620
rect 15900 -9880 16100 -9620
rect 16400 -9880 16600 -9620
rect 16900 -9880 17100 -9620
rect 17400 -9880 17600 -9620
rect 17900 -9880 18100 -9620
rect 18400 -9880 18600 -9620
rect 18900 -9880 19100 -9620
rect 19400 -9880 19600 -9620
rect 19900 -9880 20000 -9620
rect 12000 -9900 12120 -9880
rect 12380 -9900 12620 -9880
rect 12880 -9900 13120 -9880
rect 13380 -9900 13620 -9880
rect 13880 -9900 14120 -9880
rect 14380 -9900 14620 -9880
rect 14880 -9900 15120 -9880
rect 15380 -9900 15620 -9880
rect 15880 -9900 16120 -9880
rect 16380 -9900 16620 -9880
rect 16880 -9900 17120 -9880
rect 17380 -9900 17620 -9880
rect 17880 -9900 18120 -9880
rect 18380 -9900 18620 -9880
rect 18880 -9900 19120 -9880
rect 19380 -9900 19620 -9880
rect 19880 -9900 20000 -9880
rect 12000 -10100 20000 -9900
rect 12000 -10120 12120 -10100
rect 12380 -10120 12620 -10100
rect 12880 -10120 13120 -10100
rect 13380 -10120 13620 -10100
rect 13880 -10120 14120 -10100
rect 14380 -10120 14620 -10100
rect 14880 -10120 15120 -10100
rect 15380 -10120 15620 -10100
rect 15880 -10120 16120 -10100
rect 16380 -10120 16620 -10100
rect 16880 -10120 17120 -10100
rect 17380 -10120 17620 -10100
rect 17880 -10120 18120 -10100
rect 18380 -10120 18620 -10100
rect 18880 -10120 19120 -10100
rect 19380 -10120 19620 -10100
rect 19880 -10120 20000 -10100
rect 12000 -10380 12100 -10120
rect 12400 -10380 12600 -10120
rect 12900 -10380 13100 -10120
rect 13400 -10380 13600 -10120
rect 13900 -10380 14100 -10120
rect 14400 -10380 14600 -10120
rect 14900 -10380 15100 -10120
rect 15400 -10380 15600 -10120
rect 15900 -10380 16100 -10120
rect 16400 -10380 16600 -10120
rect 16900 -10380 17100 -10120
rect 17400 -10380 17600 -10120
rect 17900 -10380 18100 -10120
rect 18400 -10380 18600 -10120
rect 18900 -10380 19100 -10120
rect 19400 -10380 19600 -10120
rect 19900 -10380 20000 -10120
rect 12000 -10400 12120 -10380
rect 12380 -10400 12620 -10380
rect 12880 -10400 13120 -10380
rect 13380 -10400 13620 -10380
rect 13880 -10400 14120 -10380
rect 14380 -10400 14620 -10380
rect 14880 -10400 15120 -10380
rect 15380 -10400 15620 -10380
rect 15880 -10400 16120 -10380
rect 16380 -10400 16620 -10380
rect 16880 -10400 17120 -10380
rect 17380 -10400 17620 -10380
rect 17880 -10400 18120 -10380
rect 18380 -10400 18620 -10380
rect 18880 -10400 19120 -10380
rect 19380 -10400 19620 -10380
rect 19880 -10400 20000 -10380
rect 12000 -10600 20000 -10400
rect 12000 -10620 12120 -10600
rect 12380 -10620 12620 -10600
rect 12880 -10620 13120 -10600
rect 13380 -10620 13620 -10600
rect 13880 -10620 14120 -10600
rect 14380 -10620 14620 -10600
rect 14880 -10620 15120 -10600
rect 15380 -10620 15620 -10600
rect 15880 -10620 16120 -10600
rect 16380 -10620 16620 -10600
rect 16880 -10620 17120 -10600
rect 17380 -10620 17620 -10600
rect 17880 -10620 18120 -10600
rect 18380 -10620 18620 -10600
rect 18880 -10620 19120 -10600
rect 19380 -10620 19620 -10600
rect 19880 -10620 20000 -10600
rect 12000 -10880 12100 -10620
rect 12400 -10880 12600 -10620
rect 12900 -10880 13100 -10620
rect 13400 -10880 13600 -10620
rect 13900 -10880 14100 -10620
rect 14400 -10880 14600 -10620
rect 14900 -10880 15100 -10620
rect 15400 -10880 15600 -10620
rect 15900 -10880 16100 -10620
rect 16400 -10880 16600 -10620
rect 16900 -10880 17100 -10620
rect 17400 -10880 17600 -10620
rect 17900 -10880 18100 -10620
rect 18400 -10880 18600 -10620
rect 18900 -10880 19100 -10620
rect 19400 -10880 19600 -10620
rect 19900 -10880 20000 -10620
rect 12000 -10900 12120 -10880
rect 12380 -10900 12620 -10880
rect 12880 -10900 13120 -10880
rect 13380 -10900 13620 -10880
rect 13880 -10900 14120 -10880
rect 14380 -10900 14620 -10880
rect 14880 -10900 15120 -10880
rect 15380 -10900 15620 -10880
rect 15880 -10900 16120 -10880
rect 16380 -10900 16620 -10880
rect 16880 -10900 17120 -10880
rect 17380 -10900 17620 -10880
rect 17880 -10900 18120 -10880
rect 18380 -10900 18620 -10880
rect 18880 -10900 19120 -10880
rect 19380 -10900 19620 -10880
rect 19880 -10900 20000 -10880
rect 12000 -11100 20000 -10900
rect 12000 -11120 12120 -11100
rect 12380 -11120 12620 -11100
rect 12880 -11120 13120 -11100
rect 13380 -11120 13620 -11100
rect 13880 -11120 14120 -11100
rect 14380 -11120 14620 -11100
rect 14880 -11120 15120 -11100
rect 15380 -11120 15620 -11100
rect 15880 -11120 16120 -11100
rect 16380 -11120 16620 -11100
rect 16880 -11120 17120 -11100
rect 17380 -11120 17620 -11100
rect 17880 -11120 18120 -11100
rect 18380 -11120 18620 -11100
rect 18880 -11120 19120 -11100
rect 19380 -11120 19620 -11100
rect 19880 -11120 20000 -11100
rect 12000 -11380 12100 -11120
rect 12400 -11380 12600 -11120
rect 12900 -11380 13100 -11120
rect 13400 -11380 13600 -11120
rect 13900 -11380 14100 -11120
rect 14400 -11380 14600 -11120
rect 14900 -11380 15100 -11120
rect 15400 -11380 15600 -11120
rect 15900 -11380 16100 -11120
rect 16400 -11380 16600 -11120
rect 16900 -11380 17100 -11120
rect 17400 -11380 17600 -11120
rect 17900 -11380 18100 -11120
rect 18400 -11380 18600 -11120
rect 18900 -11380 19100 -11120
rect 19400 -11380 19600 -11120
rect 19900 -11380 20000 -11120
rect 12000 -11400 12120 -11380
rect 12380 -11400 12620 -11380
rect 12880 -11400 13120 -11380
rect 13380 -11400 13620 -11380
rect 13880 -11400 14120 -11380
rect 14380 -11400 14620 -11380
rect 14880 -11400 15120 -11380
rect 15380 -11400 15620 -11380
rect 15880 -11400 16120 -11380
rect 16380 -11400 16620 -11380
rect 16880 -11400 17120 -11380
rect 17380 -11400 17620 -11380
rect 17880 -11400 18120 -11380
rect 18380 -11400 18620 -11380
rect 18880 -11400 19120 -11380
rect 19380 -11400 19620 -11380
rect 19880 -11400 20000 -11380
rect 12000 -11600 20000 -11400
rect 12000 -11620 12120 -11600
rect 12380 -11620 12620 -11600
rect 12880 -11620 13120 -11600
rect 13380 -11620 13620 -11600
rect 13880 -11620 14120 -11600
rect 14380 -11620 14620 -11600
rect 14880 -11620 15120 -11600
rect 15380 -11620 15620 -11600
rect 15880 -11620 16120 -11600
rect 16380 -11620 16620 -11600
rect 16880 -11620 17120 -11600
rect 17380 -11620 17620 -11600
rect 17880 -11620 18120 -11600
rect 18380 -11620 18620 -11600
rect 18880 -11620 19120 -11600
rect 19380 -11620 19620 -11600
rect 19880 -11620 20000 -11600
rect 12000 -11880 12100 -11620
rect 12400 -11880 12600 -11620
rect 12900 -11880 13100 -11620
rect 13400 -11880 13600 -11620
rect 13900 -11880 14100 -11620
rect 14400 -11880 14600 -11620
rect 14900 -11880 15100 -11620
rect 15400 -11880 15600 -11620
rect 15900 -11880 16100 -11620
rect 16400 -11880 16600 -11620
rect 16900 -11880 17100 -11620
rect 17400 -11880 17600 -11620
rect 17900 -11880 18100 -11620
rect 18400 -11880 18600 -11620
rect 18900 -11880 19100 -11620
rect 19400 -11880 19600 -11620
rect 19900 -11880 20000 -11620
rect 12000 -11900 12120 -11880
rect 12380 -11900 12620 -11880
rect 12880 -11900 13120 -11880
rect 13380 -11900 13620 -11880
rect 13880 -11900 14120 -11880
rect 14380 -11900 14620 -11880
rect 14880 -11900 15120 -11880
rect 15380 -11900 15620 -11880
rect 15880 -11900 16120 -11880
rect 16380 -11900 16620 -11880
rect 16880 -11900 17120 -11880
rect 17380 -11900 17620 -11880
rect 17880 -11900 18120 -11880
rect 18380 -11900 18620 -11880
rect 18880 -11900 19120 -11880
rect 19380 -11900 19620 -11880
rect 19880 -11900 20000 -11880
rect 12000 -12100 20000 -11900
rect 12000 -12120 12120 -12100
rect 12380 -12120 12620 -12100
rect 12880 -12120 13120 -12100
rect 13380 -12120 13620 -12100
rect 13880 -12120 14120 -12100
rect 14380 -12120 14620 -12100
rect 14880 -12120 15120 -12100
rect 15380 -12120 15620 -12100
rect 15880 -12120 16120 -12100
rect 16380 -12120 16620 -12100
rect 16880 -12120 17120 -12100
rect 17380 -12120 17620 -12100
rect 17880 -12120 18120 -12100
rect 18380 -12120 18620 -12100
rect 18880 -12120 19120 -12100
rect 19380 -12120 19620 -12100
rect 19880 -12120 20000 -12100
rect 12000 -12380 12100 -12120
rect 12400 -12380 12600 -12120
rect 12900 -12380 13100 -12120
rect 13400 -12380 13600 -12120
rect 13900 -12380 14100 -12120
rect 14400 -12380 14600 -12120
rect 14900 -12380 15100 -12120
rect 15400 -12380 15600 -12120
rect 15900 -12380 16100 -12120
rect 16400 -12380 16600 -12120
rect 16900 -12380 17100 -12120
rect 17400 -12380 17600 -12120
rect 17900 -12380 18100 -12120
rect 18400 -12380 18600 -12120
rect 18900 -12380 19100 -12120
rect 19400 -12380 19600 -12120
rect 19900 -12380 20000 -12120
rect 12000 -12400 12120 -12380
rect 12380 -12400 12620 -12380
rect 12880 -12400 13120 -12380
rect 13380 -12400 13620 -12380
rect 13880 -12400 14120 -12380
rect 14380 -12400 14620 -12380
rect 14880 -12400 15120 -12380
rect 15380 -12400 15620 -12380
rect 15880 -12400 16120 -12380
rect 16380 -12400 16620 -12380
rect 16880 -12400 17120 -12380
rect 17380 -12400 17620 -12380
rect 17880 -12400 18120 -12380
rect 18380 -12400 18620 -12380
rect 18880 -12400 19120 -12380
rect 19380 -12400 19620 -12380
rect 19880 -12400 20000 -12380
rect 12000 -12600 20000 -12400
rect 12000 -12620 12120 -12600
rect 12380 -12620 12620 -12600
rect 12880 -12620 13120 -12600
rect 13380 -12620 13620 -12600
rect 13880 -12620 14120 -12600
rect 14380 -12620 14620 -12600
rect 14880 -12620 15120 -12600
rect 15380 -12620 15620 -12600
rect 15880 -12620 16120 -12600
rect 16380 -12620 16620 -12600
rect 16880 -12620 17120 -12600
rect 17380 -12620 17620 -12600
rect 17880 -12620 18120 -12600
rect 18380 -12620 18620 -12600
rect 18880 -12620 19120 -12600
rect 19380 -12620 19620 -12600
rect 19880 -12620 20000 -12600
rect 12000 -12880 12100 -12620
rect 12400 -12880 12600 -12620
rect 12900 -12880 13100 -12620
rect 13400 -12880 13600 -12620
rect 13900 -12880 14100 -12620
rect 14400 -12880 14600 -12620
rect 14900 -12880 15100 -12620
rect 15400 -12880 15600 -12620
rect 15900 -12880 16100 -12620
rect 16400 -12880 16600 -12620
rect 16900 -12880 17100 -12620
rect 17400 -12880 17600 -12620
rect 17900 -12880 18100 -12620
rect 18400 -12880 18600 -12620
rect 18900 -12880 19100 -12620
rect 19400 -12880 19600 -12620
rect 19900 -12880 20000 -12620
rect 12000 -12900 12120 -12880
rect 12380 -12900 12620 -12880
rect 12880 -12900 13120 -12880
rect 13380 -12900 13620 -12880
rect 13880 -12900 14120 -12880
rect 14380 -12900 14620 -12880
rect 14880 -12900 15120 -12880
rect 15380 -12900 15620 -12880
rect 15880 -12900 16120 -12880
rect 16380 -12900 16620 -12880
rect 16880 -12900 17120 -12880
rect 17380 -12900 17620 -12880
rect 17880 -12900 18120 -12880
rect 18380 -12900 18620 -12880
rect 18880 -12900 19120 -12880
rect 19380 -12900 19620 -12880
rect 19880 -12900 20000 -12880
rect 12000 -13100 20000 -12900
rect 12000 -13120 12120 -13100
rect 12380 -13120 12620 -13100
rect 12880 -13120 13120 -13100
rect 13380 -13120 13620 -13100
rect 13880 -13120 14120 -13100
rect 14380 -13120 14620 -13100
rect 14880 -13120 15120 -13100
rect 15380 -13120 15620 -13100
rect 15880 -13120 16120 -13100
rect 16380 -13120 16620 -13100
rect 16880 -13120 17120 -13100
rect 17380 -13120 17620 -13100
rect 17880 -13120 18120 -13100
rect 18380 -13120 18620 -13100
rect 18880 -13120 19120 -13100
rect 19380 -13120 19620 -13100
rect 19880 -13120 20000 -13100
rect 12000 -13380 12100 -13120
rect 12400 -13380 12600 -13120
rect 12900 -13380 13100 -13120
rect 13400 -13380 13600 -13120
rect 13900 -13380 14100 -13120
rect 14400 -13380 14600 -13120
rect 14900 -13380 15100 -13120
rect 15400 -13380 15600 -13120
rect 15900 -13380 16100 -13120
rect 16400 -13380 16600 -13120
rect 16900 -13380 17100 -13120
rect 17400 -13380 17600 -13120
rect 17900 -13380 18100 -13120
rect 18400 -13380 18600 -13120
rect 18900 -13380 19100 -13120
rect 19400 -13380 19600 -13120
rect 19900 -13380 20000 -13120
rect 12000 -13400 12120 -13380
rect 12380 -13400 12620 -13380
rect 12880 -13400 13120 -13380
rect 13380 -13400 13620 -13380
rect 13880 -13400 14120 -13380
rect 14380 -13400 14620 -13380
rect 14880 -13400 15120 -13380
rect 15380 -13400 15620 -13380
rect 15880 -13400 16120 -13380
rect 16380 -13400 16620 -13380
rect 16880 -13400 17120 -13380
rect 17380 -13400 17620 -13380
rect 17880 -13400 18120 -13380
rect 18380 -13400 18620 -13380
rect 18880 -13400 19120 -13380
rect 19380 -13400 19620 -13380
rect 19880 -13400 20000 -13380
rect 12000 -13600 20000 -13400
rect 12000 -13620 12120 -13600
rect 12380 -13620 12620 -13600
rect 12880 -13620 13120 -13600
rect 13380 -13620 13620 -13600
rect 13880 -13620 14120 -13600
rect 14380 -13620 14620 -13600
rect 14880 -13620 15120 -13600
rect 15380 -13620 15620 -13600
rect 15880 -13620 16120 -13600
rect 16380 -13620 16620 -13600
rect 16880 -13620 17120 -13600
rect 17380 -13620 17620 -13600
rect 17880 -13620 18120 -13600
rect 18380 -13620 18620 -13600
rect 18880 -13620 19120 -13600
rect 19380 -13620 19620 -13600
rect 19880 -13620 20000 -13600
rect 12000 -13880 12100 -13620
rect 12400 -13880 12600 -13620
rect 12900 -13880 13100 -13620
rect 13400 -13880 13600 -13620
rect 13900 -13880 14100 -13620
rect 14400 -13880 14600 -13620
rect 14900 -13880 15100 -13620
rect 15400 -13880 15600 -13620
rect 15900 -13880 16100 -13620
rect 16400 -13880 16600 -13620
rect 16900 -13880 17100 -13620
rect 17400 -13880 17600 -13620
rect 17900 -13880 18100 -13620
rect 18400 -13880 18600 -13620
rect 18900 -13880 19100 -13620
rect 19400 -13880 19600 -13620
rect 19900 -13880 20000 -13620
rect 12000 -13900 12120 -13880
rect 12380 -13900 12620 -13880
rect 12880 -13900 13120 -13880
rect 13380 -13900 13620 -13880
rect 13880 -13900 14120 -13880
rect 14380 -13900 14620 -13880
rect 14880 -13900 15120 -13880
rect 15380 -13900 15620 -13880
rect 15880 -13900 16120 -13880
rect 16380 -13900 16620 -13880
rect 16880 -13900 17120 -13880
rect 17380 -13900 17620 -13880
rect 17880 -13900 18120 -13880
rect 18380 -13900 18620 -13880
rect 18880 -13900 19120 -13880
rect 19380 -13900 19620 -13880
rect 19880 -13900 20000 -13880
rect 12000 -14000 20000 -13900
rect 88000 -2100 140000 -1980
rect 88000 -2120 88120 -2100
rect 88380 -2120 88620 -2100
rect 88880 -2120 89120 -2100
rect 89380 -2120 89620 -2100
rect 89880 -2120 90120 -2100
rect 90380 -2120 90620 -2100
rect 90880 -2120 91120 -2100
rect 91380 -2120 91620 -2100
rect 91880 -2120 92120 -2100
rect 92380 -2120 92620 -2100
rect 92880 -2120 93120 -2100
rect 93380 -2120 93620 -2100
rect 93880 -2120 94120 -2100
rect 94380 -2120 94620 -2100
rect 94880 -2120 95120 -2100
rect 95380 -2120 95620 -2100
rect 95880 -2120 96120 -2100
rect 96380 -2120 96620 -2100
rect 96880 -2120 97120 -2100
rect 97380 -2120 97620 -2100
rect 97880 -2120 98120 -2100
rect 98380 -2120 98620 -2100
rect 98880 -2120 99120 -2100
rect 99380 -2120 99620 -2100
rect 99880 -2120 100120 -2100
rect 100380 -2120 100620 -2100
rect 100880 -2120 101120 -2100
rect 101380 -2120 101620 -2100
rect 101880 -2120 102120 -2100
rect 102380 -2120 102620 -2100
rect 102880 -2120 103120 -2100
rect 103380 -2120 103620 -2100
rect 103880 -2120 104120 -2100
rect 104380 -2120 104620 -2100
rect 104880 -2120 105120 -2100
rect 105380 -2120 105620 -2100
rect 105880 -2120 106120 -2100
rect 106380 -2120 106620 -2100
rect 106880 -2120 107120 -2100
rect 107380 -2120 107620 -2100
rect 107880 -2120 108120 -2100
rect 108380 -2120 108620 -2100
rect 108880 -2120 109120 -2100
rect 109380 -2120 109620 -2100
rect 109880 -2120 110120 -2100
rect 110380 -2120 110620 -2100
rect 110880 -2120 111120 -2100
rect 111380 -2120 111620 -2100
rect 111880 -2120 112120 -2100
rect 112380 -2120 112620 -2100
rect 112880 -2120 113120 -2100
rect 113380 -2120 113620 -2100
rect 113880 -2120 114120 -2100
rect 114380 -2120 114620 -2100
rect 114880 -2120 115120 -2100
rect 115380 -2120 115620 -2100
rect 115880 -2120 116120 -2100
rect 116380 -2120 116620 -2100
rect 116880 -2120 117120 -2100
rect 117380 -2120 117620 -2100
rect 117880 -2120 118120 -2100
rect 118380 -2120 118620 -2100
rect 118880 -2120 119120 -2100
rect 119380 -2120 119620 -2100
rect 119880 -2120 120120 -2100
rect 120380 -2120 120620 -2100
rect 120880 -2120 121120 -2100
rect 121380 -2120 121620 -2100
rect 121880 -2120 122120 -2100
rect 122380 -2120 122620 -2100
rect 122880 -2120 123120 -2100
rect 123380 -2120 123620 -2100
rect 123880 -2120 124120 -2100
rect 124380 -2120 124620 -2100
rect 124880 -2120 125120 -2100
rect 125380 -2120 125620 -2100
rect 125880 -2120 126120 -2100
rect 126380 -2120 126620 -2100
rect 126880 -2120 127120 -2100
rect 127380 -2120 127620 -2100
rect 127880 -2120 128120 -2100
rect 128380 -2120 128620 -2100
rect 128880 -2120 129120 -2100
rect 129380 -2120 129620 -2100
rect 129880 -2120 130120 -2100
rect 130380 -2120 130620 -2100
rect 130880 -2120 131120 -2100
rect 131380 -2120 131620 -2100
rect 131880 -2120 132120 -2100
rect 132380 -2120 132620 -2100
rect 132880 -2120 133120 -2100
rect 133380 -2120 133620 -2100
rect 133880 -2120 134120 -2100
rect 134380 -2120 134620 -2100
rect 134880 -2120 135120 -2100
rect 135380 -2120 135620 -2100
rect 135880 -2120 136120 -2100
rect 136380 -2120 136620 -2100
rect 136880 -2120 137120 -2100
rect 137380 -2120 137620 -2100
rect 137880 -2120 138120 -2100
rect 138380 -2120 138620 -2100
rect 138880 -2120 139120 -2100
rect 139380 -2120 139620 -2100
rect 139880 -2120 140000 -2100
rect 88000 -2380 88100 -2120
rect 88400 -2380 88600 -2120
rect 88900 -2380 89100 -2120
rect 89400 -2380 89600 -2120
rect 89900 -2380 90100 -2120
rect 90400 -2380 90600 -2120
rect 90900 -2380 91100 -2120
rect 91400 -2380 91600 -2120
rect 91900 -2380 92100 -2120
rect 92400 -2380 92600 -2120
rect 92900 -2380 93100 -2120
rect 93400 -2380 93600 -2120
rect 93900 -2380 94100 -2120
rect 94400 -2380 94600 -2120
rect 94900 -2380 95100 -2120
rect 95400 -2380 95600 -2120
rect 95900 -2380 96100 -2120
rect 96400 -2380 96600 -2120
rect 96900 -2380 97100 -2120
rect 97400 -2380 97600 -2120
rect 97900 -2380 98100 -2120
rect 98400 -2380 98600 -2120
rect 98900 -2380 99100 -2120
rect 99400 -2380 99600 -2120
rect 99900 -2380 100100 -2120
rect 100400 -2380 100600 -2120
rect 100900 -2380 101100 -2120
rect 101400 -2380 101600 -2120
rect 101900 -2380 102100 -2120
rect 102400 -2380 102600 -2120
rect 102900 -2380 103100 -2120
rect 103400 -2380 103600 -2120
rect 103900 -2380 104100 -2120
rect 104400 -2380 104600 -2120
rect 104900 -2380 105100 -2120
rect 105400 -2380 105600 -2120
rect 105900 -2380 106100 -2120
rect 106400 -2380 106600 -2120
rect 106900 -2380 107100 -2120
rect 107400 -2380 107600 -2120
rect 107900 -2380 108100 -2120
rect 108400 -2380 108600 -2120
rect 108900 -2380 109100 -2120
rect 109400 -2380 109600 -2120
rect 109900 -2380 110100 -2120
rect 110400 -2380 110600 -2120
rect 110900 -2380 111100 -2120
rect 111400 -2380 111600 -2120
rect 111900 -2380 112100 -2120
rect 112400 -2380 112600 -2120
rect 112900 -2380 113100 -2120
rect 113400 -2380 113600 -2120
rect 113900 -2380 114100 -2120
rect 114400 -2380 114600 -2120
rect 114900 -2380 115100 -2120
rect 115400 -2380 115600 -2120
rect 115900 -2380 116100 -2120
rect 116400 -2380 116600 -2120
rect 116900 -2380 117100 -2120
rect 117400 -2380 117600 -2120
rect 117900 -2380 118100 -2120
rect 118400 -2380 118600 -2120
rect 118900 -2380 119100 -2120
rect 119400 -2380 119600 -2120
rect 119900 -2380 120100 -2120
rect 120400 -2380 120600 -2120
rect 120900 -2380 121100 -2120
rect 121400 -2380 121600 -2120
rect 121900 -2380 122100 -2120
rect 122400 -2380 122600 -2120
rect 122900 -2380 123100 -2120
rect 123400 -2380 123600 -2120
rect 123900 -2380 124100 -2120
rect 124400 -2380 124600 -2120
rect 124900 -2380 125100 -2120
rect 125400 -2380 125600 -2120
rect 125900 -2380 126100 -2120
rect 126400 -2380 126600 -2120
rect 126900 -2380 127100 -2120
rect 127400 -2380 127600 -2120
rect 127900 -2380 128100 -2120
rect 128400 -2380 128600 -2120
rect 128900 -2380 129100 -2120
rect 129400 -2380 129600 -2120
rect 129900 -2380 130100 -2120
rect 130400 -2380 130600 -2120
rect 130900 -2380 131100 -2120
rect 131400 -2380 131600 -2120
rect 131900 -2380 132100 -2120
rect 132400 -2380 132600 -2120
rect 132900 -2380 133100 -2120
rect 133400 -2380 133600 -2120
rect 133900 -2380 134100 -2120
rect 134400 -2380 134600 -2120
rect 134900 -2380 135100 -2120
rect 135400 -2380 135600 -2120
rect 135900 -2380 136100 -2120
rect 136400 -2380 136600 -2120
rect 136900 -2380 137100 -2120
rect 137400 -2380 137600 -2120
rect 137900 -2380 138100 -2120
rect 138400 -2380 138600 -2120
rect 138900 -2380 139100 -2120
rect 139400 -2380 139600 -2120
rect 139900 -2380 140000 -2120
rect 88000 -2400 88120 -2380
rect 88380 -2400 88620 -2380
rect 88880 -2400 89120 -2380
rect 89380 -2400 89620 -2380
rect 89880 -2400 90120 -2380
rect 90380 -2400 90620 -2380
rect 90880 -2400 91120 -2380
rect 91380 -2400 91620 -2380
rect 91880 -2400 92120 -2380
rect 92380 -2400 92620 -2380
rect 92880 -2400 93120 -2380
rect 93380 -2400 93620 -2380
rect 93880 -2400 94120 -2380
rect 94380 -2400 94620 -2380
rect 94880 -2400 95120 -2380
rect 95380 -2400 95620 -2380
rect 95880 -2400 96120 -2380
rect 96380 -2400 96620 -2380
rect 96880 -2400 97120 -2380
rect 97380 -2400 97620 -2380
rect 97880 -2400 98120 -2380
rect 98380 -2400 98620 -2380
rect 98880 -2400 99120 -2380
rect 99380 -2400 99620 -2380
rect 99880 -2400 100120 -2380
rect 100380 -2400 100620 -2380
rect 100880 -2400 101120 -2380
rect 101380 -2400 101620 -2380
rect 101880 -2400 102120 -2380
rect 102380 -2400 102620 -2380
rect 102880 -2400 103120 -2380
rect 103380 -2400 103620 -2380
rect 103880 -2400 104120 -2380
rect 104380 -2400 104620 -2380
rect 104880 -2400 105120 -2380
rect 105380 -2400 105620 -2380
rect 105880 -2400 106120 -2380
rect 106380 -2400 106620 -2380
rect 106880 -2400 107120 -2380
rect 107380 -2400 107620 -2380
rect 107880 -2400 108120 -2380
rect 108380 -2400 108620 -2380
rect 108880 -2400 109120 -2380
rect 109380 -2400 109620 -2380
rect 109880 -2400 110120 -2380
rect 110380 -2400 110620 -2380
rect 110880 -2400 111120 -2380
rect 111380 -2400 111620 -2380
rect 111880 -2400 112120 -2380
rect 112380 -2400 112620 -2380
rect 112880 -2400 113120 -2380
rect 113380 -2400 113620 -2380
rect 113880 -2400 114120 -2380
rect 114380 -2400 114620 -2380
rect 114880 -2400 115120 -2380
rect 115380 -2400 115620 -2380
rect 115880 -2400 116120 -2380
rect 116380 -2400 116620 -2380
rect 116880 -2400 117120 -2380
rect 117380 -2400 117620 -2380
rect 117880 -2400 118120 -2380
rect 118380 -2400 118620 -2380
rect 118880 -2400 119120 -2380
rect 119380 -2400 119620 -2380
rect 119880 -2400 120120 -2380
rect 120380 -2400 120620 -2380
rect 120880 -2400 121120 -2380
rect 121380 -2400 121620 -2380
rect 121880 -2400 122120 -2380
rect 122380 -2400 122620 -2380
rect 122880 -2400 123120 -2380
rect 123380 -2400 123620 -2380
rect 123880 -2400 124120 -2380
rect 124380 -2400 124620 -2380
rect 124880 -2400 125120 -2380
rect 125380 -2400 125620 -2380
rect 125880 -2400 126120 -2380
rect 126380 -2400 126620 -2380
rect 126880 -2400 127120 -2380
rect 127380 -2400 127620 -2380
rect 127880 -2400 128120 -2380
rect 128380 -2400 128620 -2380
rect 128880 -2400 129120 -2380
rect 129380 -2400 129620 -2380
rect 129880 -2400 130120 -2380
rect 130380 -2400 130620 -2380
rect 130880 -2400 131120 -2380
rect 131380 -2400 131620 -2380
rect 131880 -2400 132120 -2380
rect 132380 -2400 132620 -2380
rect 132880 -2400 133120 -2380
rect 133380 -2400 133620 -2380
rect 133880 -2400 134120 -2380
rect 134380 -2400 134620 -2380
rect 134880 -2400 135120 -2380
rect 135380 -2400 135620 -2380
rect 135880 -2400 136120 -2380
rect 136380 -2400 136620 -2380
rect 136880 -2400 137120 -2380
rect 137380 -2400 137620 -2380
rect 137880 -2400 138120 -2380
rect 138380 -2400 138620 -2380
rect 138880 -2400 139120 -2380
rect 139380 -2400 139620 -2380
rect 139880 -2400 140000 -2380
rect 88000 -2600 140000 -2400
rect 88000 -2620 88120 -2600
rect 88380 -2620 88620 -2600
rect 88880 -2620 89120 -2600
rect 89380 -2620 89620 -2600
rect 89880 -2620 90120 -2600
rect 90380 -2620 90620 -2600
rect 90880 -2620 91120 -2600
rect 91380 -2620 91620 -2600
rect 91880 -2620 92120 -2600
rect 92380 -2620 92620 -2600
rect 92880 -2620 93120 -2600
rect 93380 -2620 93620 -2600
rect 93880 -2620 94120 -2600
rect 94380 -2620 94620 -2600
rect 94880 -2620 95120 -2600
rect 95380 -2620 95620 -2600
rect 95880 -2620 96120 -2600
rect 96380 -2620 96620 -2600
rect 96880 -2620 97120 -2600
rect 97380 -2620 97620 -2600
rect 97880 -2620 98120 -2600
rect 98380 -2620 98620 -2600
rect 98880 -2620 99120 -2600
rect 99380 -2620 99620 -2600
rect 99880 -2620 100120 -2600
rect 100380 -2620 100620 -2600
rect 100880 -2620 101120 -2600
rect 101380 -2620 101620 -2600
rect 101880 -2620 102120 -2600
rect 102380 -2620 102620 -2600
rect 102880 -2620 103120 -2600
rect 103380 -2620 103620 -2600
rect 103880 -2620 104120 -2600
rect 104380 -2620 104620 -2600
rect 104880 -2620 105120 -2600
rect 105380 -2620 105620 -2600
rect 105880 -2620 106120 -2600
rect 106380 -2620 106620 -2600
rect 106880 -2620 107120 -2600
rect 107380 -2620 107620 -2600
rect 107880 -2620 108120 -2600
rect 108380 -2620 108620 -2600
rect 108880 -2620 109120 -2600
rect 109380 -2620 109620 -2600
rect 109880 -2620 110120 -2600
rect 110380 -2620 110620 -2600
rect 110880 -2620 111120 -2600
rect 111380 -2620 111620 -2600
rect 111880 -2620 112120 -2600
rect 112380 -2620 112620 -2600
rect 112880 -2620 113120 -2600
rect 113380 -2620 113620 -2600
rect 113880 -2620 114120 -2600
rect 114380 -2620 114620 -2600
rect 114880 -2620 115120 -2600
rect 115380 -2620 115620 -2600
rect 115880 -2620 116120 -2600
rect 116380 -2620 116620 -2600
rect 116880 -2620 117120 -2600
rect 117380 -2620 117620 -2600
rect 117880 -2620 118120 -2600
rect 118380 -2620 118620 -2600
rect 118880 -2620 119120 -2600
rect 119380 -2620 119620 -2600
rect 119880 -2620 120120 -2600
rect 120380 -2620 120620 -2600
rect 120880 -2620 121120 -2600
rect 121380 -2620 121620 -2600
rect 121880 -2620 122120 -2600
rect 122380 -2620 122620 -2600
rect 122880 -2620 123120 -2600
rect 123380 -2620 123620 -2600
rect 123880 -2620 124120 -2600
rect 124380 -2620 124620 -2600
rect 124880 -2620 125120 -2600
rect 125380 -2620 125620 -2600
rect 125880 -2620 126120 -2600
rect 126380 -2620 126620 -2600
rect 126880 -2620 127120 -2600
rect 127380 -2620 127620 -2600
rect 127880 -2620 128120 -2600
rect 128380 -2620 128620 -2600
rect 128880 -2620 129120 -2600
rect 129380 -2620 129620 -2600
rect 129880 -2620 130120 -2600
rect 130380 -2620 130620 -2600
rect 130880 -2620 131120 -2600
rect 131380 -2620 131620 -2600
rect 131880 -2620 132120 -2600
rect 132380 -2620 132620 -2600
rect 132880 -2620 133120 -2600
rect 133380 -2620 133620 -2600
rect 133880 -2620 134120 -2600
rect 134380 -2620 134620 -2600
rect 134880 -2620 135120 -2600
rect 135380 -2620 135620 -2600
rect 135880 -2620 136120 -2600
rect 136380 -2620 136620 -2600
rect 136880 -2620 137120 -2600
rect 137380 -2620 137620 -2600
rect 137880 -2620 138120 -2600
rect 138380 -2620 138620 -2600
rect 138880 -2620 139120 -2600
rect 139380 -2620 139620 -2600
rect 139880 -2620 140000 -2600
rect 88000 -2880 88100 -2620
rect 88400 -2880 88600 -2620
rect 88900 -2880 89100 -2620
rect 89400 -2880 89600 -2620
rect 89900 -2880 90100 -2620
rect 90400 -2880 90600 -2620
rect 90900 -2880 91100 -2620
rect 91400 -2880 91600 -2620
rect 91900 -2880 92100 -2620
rect 92400 -2880 92600 -2620
rect 92900 -2880 93100 -2620
rect 93400 -2880 93600 -2620
rect 93900 -2880 94100 -2620
rect 94400 -2880 94600 -2620
rect 94900 -2880 95100 -2620
rect 95400 -2880 95600 -2620
rect 95900 -2880 96100 -2620
rect 96400 -2880 96600 -2620
rect 96900 -2880 97100 -2620
rect 97400 -2880 97600 -2620
rect 97900 -2880 98100 -2620
rect 98400 -2880 98600 -2620
rect 98900 -2880 99100 -2620
rect 99400 -2880 99600 -2620
rect 99900 -2880 100100 -2620
rect 100400 -2880 100600 -2620
rect 100900 -2880 101100 -2620
rect 101400 -2880 101600 -2620
rect 101900 -2880 102100 -2620
rect 102400 -2880 102600 -2620
rect 102900 -2880 103100 -2620
rect 103400 -2880 103600 -2620
rect 103900 -2880 104100 -2620
rect 104400 -2880 104600 -2620
rect 104900 -2880 105100 -2620
rect 105400 -2880 105600 -2620
rect 105900 -2880 106100 -2620
rect 106400 -2880 106600 -2620
rect 106900 -2880 107100 -2620
rect 107400 -2880 107600 -2620
rect 107900 -2880 108100 -2620
rect 108400 -2880 108600 -2620
rect 108900 -2880 109100 -2620
rect 109400 -2880 109600 -2620
rect 109900 -2880 110100 -2620
rect 110400 -2880 110600 -2620
rect 110900 -2880 111100 -2620
rect 111400 -2880 111600 -2620
rect 111900 -2880 112100 -2620
rect 112400 -2880 112600 -2620
rect 112900 -2880 113100 -2620
rect 113400 -2880 113600 -2620
rect 113900 -2880 114100 -2620
rect 114400 -2880 114600 -2620
rect 114900 -2880 115100 -2620
rect 115400 -2880 115600 -2620
rect 115900 -2880 116100 -2620
rect 116400 -2880 116600 -2620
rect 116900 -2880 117100 -2620
rect 117400 -2880 117600 -2620
rect 117900 -2880 118100 -2620
rect 118400 -2880 118600 -2620
rect 118900 -2880 119100 -2620
rect 119400 -2880 119600 -2620
rect 119900 -2880 120100 -2620
rect 120400 -2880 120600 -2620
rect 120900 -2880 121100 -2620
rect 121400 -2880 121600 -2620
rect 121900 -2880 122100 -2620
rect 122400 -2880 122600 -2620
rect 122900 -2880 123100 -2620
rect 123400 -2880 123600 -2620
rect 123900 -2880 124100 -2620
rect 124400 -2880 124600 -2620
rect 124900 -2880 125100 -2620
rect 125400 -2880 125600 -2620
rect 125900 -2880 126100 -2620
rect 126400 -2880 126600 -2620
rect 126900 -2880 127100 -2620
rect 127400 -2880 127600 -2620
rect 127900 -2880 128100 -2620
rect 128400 -2880 128600 -2620
rect 128900 -2880 129100 -2620
rect 129400 -2880 129600 -2620
rect 129900 -2880 130100 -2620
rect 130400 -2880 130600 -2620
rect 130900 -2880 131100 -2620
rect 131400 -2880 131600 -2620
rect 131900 -2880 132100 -2620
rect 132400 -2880 132600 -2620
rect 132900 -2880 133100 -2620
rect 133400 -2880 133600 -2620
rect 133900 -2880 134100 -2620
rect 134400 -2880 134600 -2620
rect 134900 -2880 135100 -2620
rect 135400 -2880 135600 -2620
rect 135900 -2880 136100 -2620
rect 136400 -2880 136600 -2620
rect 136900 -2880 137100 -2620
rect 137400 -2880 137600 -2620
rect 137900 -2880 138100 -2620
rect 138400 -2880 138600 -2620
rect 138900 -2880 139100 -2620
rect 139400 -2880 139600 -2620
rect 139900 -2880 140000 -2620
rect 88000 -2900 88120 -2880
rect 88380 -2900 88620 -2880
rect 88880 -2900 89120 -2880
rect 89380 -2900 89620 -2880
rect 89880 -2900 90120 -2880
rect 90380 -2900 90620 -2880
rect 90880 -2900 91120 -2880
rect 91380 -2900 91620 -2880
rect 91880 -2900 92120 -2880
rect 92380 -2900 92620 -2880
rect 92880 -2900 93120 -2880
rect 93380 -2900 93620 -2880
rect 93880 -2900 94120 -2880
rect 94380 -2900 94620 -2880
rect 94880 -2900 95120 -2880
rect 95380 -2900 95620 -2880
rect 95880 -2900 96120 -2880
rect 96380 -2900 96620 -2880
rect 96880 -2900 97120 -2880
rect 97380 -2900 97620 -2880
rect 97880 -2900 98120 -2880
rect 98380 -2900 98620 -2880
rect 98880 -2900 99120 -2880
rect 99380 -2900 99620 -2880
rect 99880 -2900 100120 -2880
rect 100380 -2900 100620 -2880
rect 100880 -2900 101120 -2880
rect 101380 -2900 101620 -2880
rect 101880 -2900 102120 -2880
rect 102380 -2900 102620 -2880
rect 102880 -2900 103120 -2880
rect 103380 -2900 103620 -2880
rect 103880 -2900 104120 -2880
rect 104380 -2900 104620 -2880
rect 104880 -2900 105120 -2880
rect 105380 -2900 105620 -2880
rect 105880 -2900 106120 -2880
rect 106380 -2900 106620 -2880
rect 106880 -2900 107120 -2880
rect 107380 -2900 107620 -2880
rect 107880 -2900 108120 -2880
rect 108380 -2900 108620 -2880
rect 108880 -2900 109120 -2880
rect 109380 -2900 109620 -2880
rect 109880 -2900 110120 -2880
rect 110380 -2900 110620 -2880
rect 110880 -2900 111120 -2880
rect 111380 -2900 111620 -2880
rect 111880 -2900 112120 -2880
rect 112380 -2900 112620 -2880
rect 112880 -2900 113120 -2880
rect 113380 -2900 113620 -2880
rect 113880 -2900 114120 -2880
rect 114380 -2900 114620 -2880
rect 114880 -2900 115120 -2880
rect 115380 -2900 115620 -2880
rect 115880 -2900 116120 -2880
rect 116380 -2900 116620 -2880
rect 116880 -2900 117120 -2880
rect 117380 -2900 117620 -2880
rect 117880 -2900 118120 -2880
rect 118380 -2900 118620 -2880
rect 118880 -2900 119120 -2880
rect 119380 -2900 119620 -2880
rect 119880 -2900 120120 -2880
rect 120380 -2900 120620 -2880
rect 120880 -2900 121120 -2880
rect 121380 -2900 121620 -2880
rect 121880 -2900 122120 -2880
rect 122380 -2900 122620 -2880
rect 122880 -2900 123120 -2880
rect 123380 -2900 123620 -2880
rect 123880 -2900 124120 -2880
rect 124380 -2900 124620 -2880
rect 124880 -2900 125120 -2880
rect 125380 -2900 125620 -2880
rect 125880 -2900 126120 -2880
rect 126380 -2900 126620 -2880
rect 126880 -2900 127120 -2880
rect 127380 -2900 127620 -2880
rect 127880 -2900 128120 -2880
rect 128380 -2900 128620 -2880
rect 128880 -2900 129120 -2880
rect 129380 -2900 129620 -2880
rect 129880 -2900 130120 -2880
rect 130380 -2900 130620 -2880
rect 130880 -2900 131120 -2880
rect 131380 -2900 131620 -2880
rect 131880 -2900 132120 -2880
rect 132380 -2900 132620 -2880
rect 132880 -2900 133120 -2880
rect 133380 -2900 133620 -2880
rect 133880 -2900 134120 -2880
rect 134380 -2900 134620 -2880
rect 134880 -2900 135120 -2880
rect 135380 -2900 135620 -2880
rect 135880 -2900 136120 -2880
rect 136380 -2900 136620 -2880
rect 136880 -2900 137120 -2880
rect 137380 -2900 137620 -2880
rect 137880 -2900 138120 -2880
rect 138380 -2900 138620 -2880
rect 138880 -2900 139120 -2880
rect 139380 -2900 139620 -2880
rect 139880 -2900 140000 -2880
rect 88000 -3100 140000 -2900
rect 88000 -3120 88120 -3100
rect 88380 -3120 88620 -3100
rect 88880 -3120 89120 -3100
rect 89380 -3120 89620 -3100
rect 89880 -3120 90120 -3100
rect 90380 -3120 90620 -3100
rect 90880 -3120 91120 -3100
rect 91380 -3120 91620 -3100
rect 91880 -3120 92120 -3100
rect 92380 -3120 92620 -3100
rect 92880 -3120 93120 -3100
rect 93380 -3120 93620 -3100
rect 93880 -3120 94120 -3100
rect 94380 -3120 94620 -3100
rect 94880 -3120 95120 -3100
rect 95380 -3120 95620 -3100
rect 95880 -3120 96120 -3100
rect 96380 -3120 96620 -3100
rect 96880 -3120 97120 -3100
rect 97380 -3120 97620 -3100
rect 97880 -3120 98120 -3100
rect 98380 -3120 98620 -3100
rect 98880 -3120 99120 -3100
rect 99380 -3120 99620 -3100
rect 99880 -3120 100120 -3100
rect 100380 -3120 100620 -3100
rect 100880 -3120 101120 -3100
rect 101380 -3120 101620 -3100
rect 101880 -3120 102120 -3100
rect 102380 -3120 102620 -3100
rect 102880 -3120 103120 -3100
rect 103380 -3120 103620 -3100
rect 103880 -3120 104120 -3100
rect 104380 -3120 104620 -3100
rect 104880 -3120 105120 -3100
rect 105380 -3120 105620 -3100
rect 105880 -3120 106120 -3100
rect 106380 -3120 106620 -3100
rect 106880 -3120 107120 -3100
rect 107380 -3120 107620 -3100
rect 107880 -3120 108120 -3100
rect 108380 -3120 108620 -3100
rect 108880 -3120 109120 -3100
rect 109380 -3120 109620 -3100
rect 109880 -3120 110120 -3100
rect 110380 -3120 110620 -3100
rect 110880 -3120 111120 -3100
rect 111380 -3120 111620 -3100
rect 111880 -3120 112120 -3100
rect 112380 -3120 112620 -3100
rect 112880 -3120 113120 -3100
rect 113380 -3120 113620 -3100
rect 113880 -3120 114120 -3100
rect 114380 -3120 114620 -3100
rect 114880 -3120 115120 -3100
rect 115380 -3120 115620 -3100
rect 115880 -3120 116120 -3100
rect 116380 -3120 116620 -3100
rect 116880 -3120 117120 -3100
rect 117380 -3120 117620 -3100
rect 117880 -3120 118120 -3100
rect 118380 -3120 118620 -3100
rect 118880 -3120 119120 -3100
rect 119380 -3120 119620 -3100
rect 119880 -3120 120120 -3100
rect 120380 -3120 120620 -3100
rect 120880 -3120 121120 -3100
rect 121380 -3120 121620 -3100
rect 121880 -3120 122120 -3100
rect 122380 -3120 122620 -3100
rect 122880 -3120 123120 -3100
rect 123380 -3120 123620 -3100
rect 123880 -3120 124120 -3100
rect 124380 -3120 124620 -3100
rect 124880 -3120 125120 -3100
rect 125380 -3120 125620 -3100
rect 125880 -3120 126120 -3100
rect 126380 -3120 126620 -3100
rect 126880 -3120 127120 -3100
rect 127380 -3120 127620 -3100
rect 127880 -3120 128120 -3100
rect 128380 -3120 128620 -3100
rect 128880 -3120 129120 -3100
rect 129380 -3120 129620 -3100
rect 129880 -3120 130120 -3100
rect 130380 -3120 130620 -3100
rect 130880 -3120 131120 -3100
rect 131380 -3120 131620 -3100
rect 131880 -3120 132120 -3100
rect 132380 -3120 132620 -3100
rect 132880 -3120 133120 -3100
rect 133380 -3120 133620 -3100
rect 133880 -3120 134120 -3100
rect 134380 -3120 134620 -3100
rect 134880 -3120 135120 -3100
rect 135380 -3120 135620 -3100
rect 135880 -3120 136120 -3100
rect 136380 -3120 136620 -3100
rect 136880 -3120 137120 -3100
rect 137380 -3120 137620 -3100
rect 137880 -3120 138120 -3100
rect 138380 -3120 138620 -3100
rect 138880 -3120 139120 -3100
rect 139380 -3120 139620 -3100
rect 139880 -3120 140000 -3100
rect 88000 -3380 88100 -3120
rect 88400 -3380 88600 -3120
rect 88900 -3380 89100 -3120
rect 89400 -3380 89600 -3120
rect 89900 -3380 90100 -3120
rect 90400 -3380 90600 -3120
rect 90900 -3380 91100 -3120
rect 91400 -3380 91600 -3120
rect 91900 -3380 92100 -3120
rect 92400 -3380 92600 -3120
rect 92900 -3380 93100 -3120
rect 93400 -3380 93600 -3120
rect 93900 -3380 94100 -3120
rect 94400 -3380 94600 -3120
rect 94900 -3380 95100 -3120
rect 95400 -3380 95600 -3120
rect 95900 -3380 96100 -3120
rect 96400 -3380 96600 -3120
rect 96900 -3380 97100 -3120
rect 97400 -3380 97600 -3120
rect 97900 -3380 98100 -3120
rect 98400 -3380 98600 -3120
rect 98900 -3380 99100 -3120
rect 99400 -3380 99600 -3120
rect 99900 -3380 100100 -3120
rect 100400 -3380 100600 -3120
rect 100900 -3380 101100 -3120
rect 101400 -3380 101600 -3120
rect 101900 -3380 102100 -3120
rect 102400 -3380 102600 -3120
rect 102900 -3380 103100 -3120
rect 103400 -3380 103600 -3120
rect 103900 -3380 104100 -3120
rect 104400 -3380 104600 -3120
rect 104900 -3380 105100 -3120
rect 105400 -3380 105600 -3120
rect 105900 -3380 106100 -3120
rect 106400 -3380 106600 -3120
rect 106900 -3380 107100 -3120
rect 107400 -3380 107600 -3120
rect 107900 -3380 108100 -3120
rect 108400 -3380 108600 -3120
rect 108900 -3380 109100 -3120
rect 109400 -3380 109600 -3120
rect 109900 -3380 110100 -3120
rect 110400 -3380 110600 -3120
rect 110900 -3380 111100 -3120
rect 111400 -3380 111600 -3120
rect 111900 -3380 112100 -3120
rect 112400 -3380 112600 -3120
rect 112900 -3380 113100 -3120
rect 113400 -3380 113600 -3120
rect 113900 -3380 114100 -3120
rect 114400 -3380 114600 -3120
rect 114900 -3380 115100 -3120
rect 115400 -3380 115600 -3120
rect 115900 -3380 116100 -3120
rect 116400 -3380 116600 -3120
rect 116900 -3380 117100 -3120
rect 117400 -3380 117600 -3120
rect 117900 -3380 118100 -3120
rect 118400 -3380 118600 -3120
rect 118900 -3380 119100 -3120
rect 119400 -3380 119600 -3120
rect 119900 -3380 120100 -3120
rect 120400 -3380 120600 -3120
rect 120900 -3380 121100 -3120
rect 121400 -3380 121600 -3120
rect 121900 -3380 122100 -3120
rect 122400 -3380 122600 -3120
rect 122900 -3380 123100 -3120
rect 123400 -3380 123600 -3120
rect 123900 -3380 124100 -3120
rect 124400 -3380 124600 -3120
rect 124900 -3380 125100 -3120
rect 125400 -3380 125600 -3120
rect 125900 -3380 126100 -3120
rect 126400 -3380 126600 -3120
rect 126900 -3380 127100 -3120
rect 127400 -3380 127600 -3120
rect 127900 -3380 128100 -3120
rect 128400 -3380 128600 -3120
rect 128900 -3380 129100 -3120
rect 129400 -3380 129600 -3120
rect 129900 -3380 130100 -3120
rect 130400 -3380 130600 -3120
rect 130900 -3380 131100 -3120
rect 131400 -3380 131600 -3120
rect 131900 -3380 132100 -3120
rect 132400 -3380 132600 -3120
rect 132900 -3380 133100 -3120
rect 133400 -3380 133600 -3120
rect 133900 -3380 134100 -3120
rect 134400 -3380 134600 -3120
rect 134900 -3380 135100 -3120
rect 135400 -3380 135600 -3120
rect 135900 -3380 136100 -3120
rect 136400 -3380 136600 -3120
rect 136900 -3380 137100 -3120
rect 137400 -3380 137600 -3120
rect 137900 -3380 138100 -3120
rect 138400 -3380 138600 -3120
rect 138900 -3380 139100 -3120
rect 139400 -3380 139600 -3120
rect 139900 -3380 140000 -3120
rect 88000 -3400 88120 -3380
rect 88380 -3400 88620 -3380
rect 88880 -3400 89120 -3380
rect 89380 -3400 89620 -3380
rect 89880 -3400 90120 -3380
rect 90380 -3400 90620 -3380
rect 90880 -3400 91120 -3380
rect 91380 -3400 91620 -3380
rect 91880 -3400 92120 -3380
rect 92380 -3400 92620 -3380
rect 92880 -3400 93120 -3380
rect 93380 -3400 93620 -3380
rect 93880 -3400 94120 -3380
rect 94380 -3400 94620 -3380
rect 94880 -3400 95120 -3380
rect 95380 -3400 95620 -3380
rect 95880 -3400 96120 -3380
rect 96380 -3400 96620 -3380
rect 96880 -3400 97120 -3380
rect 97380 -3400 97620 -3380
rect 97880 -3400 98120 -3380
rect 98380 -3400 98620 -3380
rect 98880 -3400 99120 -3380
rect 99380 -3400 99620 -3380
rect 99880 -3400 100120 -3380
rect 100380 -3400 100620 -3380
rect 100880 -3400 101120 -3380
rect 101380 -3400 101620 -3380
rect 101880 -3400 102120 -3380
rect 102380 -3400 102620 -3380
rect 102880 -3400 103120 -3380
rect 103380 -3400 103620 -3380
rect 103880 -3400 104120 -3380
rect 104380 -3400 104620 -3380
rect 104880 -3400 105120 -3380
rect 105380 -3400 105620 -3380
rect 105880 -3400 106120 -3380
rect 106380 -3400 106620 -3380
rect 106880 -3400 107120 -3380
rect 107380 -3400 107620 -3380
rect 107880 -3400 108120 -3380
rect 108380 -3400 108620 -3380
rect 108880 -3400 109120 -3380
rect 109380 -3400 109620 -3380
rect 109880 -3400 110120 -3380
rect 110380 -3400 110620 -3380
rect 110880 -3400 111120 -3380
rect 111380 -3400 111620 -3380
rect 111880 -3400 112120 -3380
rect 112380 -3400 112620 -3380
rect 112880 -3400 113120 -3380
rect 113380 -3400 113620 -3380
rect 113880 -3400 114120 -3380
rect 114380 -3400 114620 -3380
rect 114880 -3400 115120 -3380
rect 115380 -3400 115620 -3380
rect 115880 -3400 116120 -3380
rect 116380 -3400 116620 -3380
rect 116880 -3400 117120 -3380
rect 117380 -3400 117620 -3380
rect 117880 -3400 118120 -3380
rect 118380 -3400 118620 -3380
rect 118880 -3400 119120 -3380
rect 119380 -3400 119620 -3380
rect 119880 -3400 120120 -3380
rect 120380 -3400 120620 -3380
rect 120880 -3400 121120 -3380
rect 121380 -3400 121620 -3380
rect 121880 -3400 122120 -3380
rect 122380 -3400 122620 -3380
rect 122880 -3400 123120 -3380
rect 123380 -3400 123620 -3380
rect 123880 -3400 124120 -3380
rect 124380 -3400 124620 -3380
rect 124880 -3400 125120 -3380
rect 125380 -3400 125620 -3380
rect 125880 -3400 126120 -3380
rect 126380 -3400 126620 -3380
rect 126880 -3400 127120 -3380
rect 127380 -3400 127620 -3380
rect 127880 -3400 128120 -3380
rect 128380 -3400 128620 -3380
rect 128880 -3400 129120 -3380
rect 129380 -3400 129620 -3380
rect 129880 -3400 130120 -3380
rect 130380 -3400 130620 -3380
rect 130880 -3400 131120 -3380
rect 131380 -3400 131620 -3380
rect 131880 -3400 132120 -3380
rect 132380 -3400 132620 -3380
rect 132880 -3400 133120 -3380
rect 133380 -3400 133620 -3380
rect 133880 -3400 134120 -3380
rect 134380 -3400 134620 -3380
rect 134880 -3400 135120 -3380
rect 135380 -3400 135620 -3380
rect 135880 -3400 136120 -3380
rect 136380 -3400 136620 -3380
rect 136880 -3400 137120 -3380
rect 137380 -3400 137620 -3380
rect 137880 -3400 138120 -3380
rect 138380 -3400 138620 -3380
rect 138880 -3400 139120 -3380
rect 139380 -3400 139620 -3380
rect 139880 -3400 140000 -3380
rect 88000 -3600 140000 -3400
rect 88000 -3620 88120 -3600
rect 88380 -3620 88620 -3600
rect 88880 -3620 89120 -3600
rect 89380 -3620 89620 -3600
rect 89880 -3620 90120 -3600
rect 90380 -3620 90620 -3600
rect 90880 -3620 91120 -3600
rect 91380 -3620 91620 -3600
rect 91880 -3620 92120 -3600
rect 92380 -3620 92620 -3600
rect 92880 -3620 93120 -3600
rect 93380 -3620 93620 -3600
rect 93880 -3620 94120 -3600
rect 94380 -3620 94620 -3600
rect 94880 -3620 95120 -3600
rect 95380 -3620 95620 -3600
rect 95880 -3620 96120 -3600
rect 96380 -3620 96620 -3600
rect 96880 -3620 97120 -3600
rect 97380 -3620 97620 -3600
rect 97880 -3620 98120 -3600
rect 98380 -3620 98620 -3600
rect 98880 -3620 99120 -3600
rect 99380 -3620 99620 -3600
rect 99880 -3620 100120 -3600
rect 100380 -3620 100620 -3600
rect 100880 -3620 101120 -3600
rect 101380 -3620 101620 -3600
rect 101880 -3620 102120 -3600
rect 102380 -3620 102620 -3600
rect 102880 -3620 103120 -3600
rect 103380 -3620 103620 -3600
rect 103880 -3620 104120 -3600
rect 104380 -3620 104620 -3600
rect 104880 -3620 105120 -3600
rect 105380 -3620 105620 -3600
rect 105880 -3620 106120 -3600
rect 106380 -3620 106620 -3600
rect 106880 -3620 107120 -3600
rect 107380 -3620 107620 -3600
rect 107880 -3620 108120 -3600
rect 108380 -3620 108620 -3600
rect 108880 -3620 109120 -3600
rect 109380 -3620 109620 -3600
rect 109880 -3620 110120 -3600
rect 110380 -3620 110620 -3600
rect 110880 -3620 111120 -3600
rect 111380 -3620 111620 -3600
rect 111880 -3620 112120 -3600
rect 112380 -3620 112620 -3600
rect 112880 -3620 113120 -3600
rect 113380 -3620 113620 -3600
rect 113880 -3620 114120 -3600
rect 114380 -3620 114620 -3600
rect 114880 -3620 115120 -3600
rect 115380 -3620 115620 -3600
rect 115880 -3620 116120 -3600
rect 116380 -3620 116620 -3600
rect 116880 -3620 117120 -3600
rect 117380 -3620 117620 -3600
rect 117880 -3620 118120 -3600
rect 118380 -3620 118620 -3600
rect 118880 -3620 119120 -3600
rect 119380 -3620 119620 -3600
rect 119880 -3620 120120 -3600
rect 120380 -3620 120620 -3600
rect 120880 -3620 121120 -3600
rect 121380 -3620 121620 -3600
rect 121880 -3620 122120 -3600
rect 122380 -3620 122620 -3600
rect 122880 -3620 123120 -3600
rect 123380 -3620 123620 -3600
rect 123880 -3620 124120 -3600
rect 124380 -3620 124620 -3600
rect 124880 -3620 125120 -3600
rect 125380 -3620 125620 -3600
rect 125880 -3620 126120 -3600
rect 126380 -3620 126620 -3600
rect 126880 -3620 127120 -3600
rect 127380 -3620 127620 -3600
rect 127880 -3620 128120 -3600
rect 128380 -3620 128620 -3600
rect 128880 -3620 129120 -3600
rect 129380 -3620 129620 -3600
rect 129880 -3620 130120 -3600
rect 130380 -3620 130620 -3600
rect 130880 -3620 131120 -3600
rect 131380 -3620 131620 -3600
rect 131880 -3620 132120 -3600
rect 132380 -3620 132620 -3600
rect 132880 -3620 133120 -3600
rect 133380 -3620 133620 -3600
rect 133880 -3620 134120 -3600
rect 134380 -3620 134620 -3600
rect 134880 -3620 135120 -3600
rect 135380 -3620 135620 -3600
rect 135880 -3620 136120 -3600
rect 136380 -3620 136620 -3600
rect 136880 -3620 137120 -3600
rect 137380 -3620 137620 -3600
rect 137880 -3620 138120 -3600
rect 138380 -3620 138620 -3600
rect 138880 -3620 139120 -3600
rect 139380 -3620 139620 -3600
rect 139880 -3620 140000 -3600
rect 88000 -3880 88100 -3620
rect 88400 -3880 88600 -3620
rect 88900 -3880 89100 -3620
rect 89400 -3880 89600 -3620
rect 89900 -3880 90100 -3620
rect 90400 -3880 90600 -3620
rect 90900 -3880 91100 -3620
rect 91400 -3880 91600 -3620
rect 91900 -3880 92100 -3620
rect 92400 -3880 92600 -3620
rect 92900 -3880 93100 -3620
rect 93400 -3880 93600 -3620
rect 93900 -3880 94100 -3620
rect 94400 -3880 94600 -3620
rect 94900 -3880 95100 -3620
rect 95400 -3880 95600 -3620
rect 95900 -3880 96100 -3620
rect 96400 -3880 96600 -3620
rect 96900 -3880 97100 -3620
rect 97400 -3880 97600 -3620
rect 97900 -3880 98100 -3620
rect 98400 -3880 98600 -3620
rect 98900 -3880 99100 -3620
rect 99400 -3880 99600 -3620
rect 99900 -3880 100100 -3620
rect 100400 -3880 100600 -3620
rect 100900 -3880 101100 -3620
rect 101400 -3880 101600 -3620
rect 101900 -3880 102100 -3620
rect 102400 -3880 102600 -3620
rect 102900 -3880 103100 -3620
rect 103400 -3880 103600 -3620
rect 103900 -3880 104100 -3620
rect 104400 -3880 104600 -3620
rect 104900 -3880 105100 -3620
rect 105400 -3880 105600 -3620
rect 105900 -3880 106100 -3620
rect 106400 -3880 106600 -3620
rect 106900 -3880 107100 -3620
rect 107400 -3880 107600 -3620
rect 107900 -3880 108100 -3620
rect 108400 -3880 108600 -3620
rect 108900 -3880 109100 -3620
rect 109400 -3880 109600 -3620
rect 109900 -3880 110100 -3620
rect 110400 -3880 110600 -3620
rect 110900 -3880 111100 -3620
rect 111400 -3880 111600 -3620
rect 111900 -3880 112100 -3620
rect 112400 -3880 112600 -3620
rect 112900 -3880 113100 -3620
rect 113400 -3880 113600 -3620
rect 113900 -3880 114100 -3620
rect 114400 -3880 114600 -3620
rect 114900 -3880 115100 -3620
rect 115400 -3880 115600 -3620
rect 115900 -3880 116100 -3620
rect 116400 -3880 116600 -3620
rect 116900 -3880 117100 -3620
rect 117400 -3880 117600 -3620
rect 117900 -3880 118100 -3620
rect 118400 -3880 118600 -3620
rect 118900 -3880 119100 -3620
rect 119400 -3880 119600 -3620
rect 119900 -3880 120100 -3620
rect 120400 -3880 120600 -3620
rect 120900 -3880 121100 -3620
rect 121400 -3880 121600 -3620
rect 121900 -3880 122100 -3620
rect 122400 -3880 122600 -3620
rect 122900 -3880 123100 -3620
rect 123400 -3880 123600 -3620
rect 123900 -3880 124100 -3620
rect 124400 -3880 124600 -3620
rect 124900 -3880 125100 -3620
rect 125400 -3880 125600 -3620
rect 125900 -3880 126100 -3620
rect 126400 -3880 126600 -3620
rect 126900 -3880 127100 -3620
rect 127400 -3880 127600 -3620
rect 127900 -3880 128100 -3620
rect 128400 -3880 128600 -3620
rect 128900 -3880 129100 -3620
rect 129400 -3880 129600 -3620
rect 129900 -3880 130100 -3620
rect 130400 -3880 130600 -3620
rect 130900 -3880 131100 -3620
rect 131400 -3880 131600 -3620
rect 131900 -3880 132100 -3620
rect 132400 -3880 132600 -3620
rect 132900 -3880 133100 -3620
rect 133400 -3880 133600 -3620
rect 133900 -3880 134100 -3620
rect 134400 -3880 134600 -3620
rect 134900 -3880 135100 -3620
rect 135400 -3880 135600 -3620
rect 135900 -3880 136100 -3620
rect 136400 -3880 136600 -3620
rect 136900 -3880 137100 -3620
rect 137400 -3880 137600 -3620
rect 137900 -3880 138100 -3620
rect 138400 -3880 138600 -3620
rect 138900 -3880 139100 -3620
rect 139400 -3880 139600 -3620
rect 139900 -3880 140000 -3620
rect 88000 -3900 88120 -3880
rect 88380 -3900 88620 -3880
rect 88880 -3900 89120 -3880
rect 89380 -3900 89620 -3880
rect 89880 -3900 90120 -3880
rect 90380 -3900 90620 -3880
rect 90880 -3900 91120 -3880
rect 91380 -3900 91620 -3880
rect 91880 -3900 92120 -3880
rect 92380 -3900 92620 -3880
rect 92880 -3900 93120 -3880
rect 93380 -3900 93620 -3880
rect 93880 -3900 94120 -3880
rect 94380 -3900 94620 -3880
rect 94880 -3900 95120 -3880
rect 95380 -3900 95620 -3880
rect 95880 -3900 96120 -3880
rect 96380 -3900 96620 -3880
rect 96880 -3900 97120 -3880
rect 97380 -3900 97620 -3880
rect 97880 -3900 98120 -3880
rect 98380 -3900 98620 -3880
rect 98880 -3900 99120 -3880
rect 99380 -3900 99620 -3880
rect 99880 -3900 100120 -3880
rect 100380 -3900 100620 -3880
rect 100880 -3900 101120 -3880
rect 101380 -3900 101620 -3880
rect 101880 -3900 102120 -3880
rect 102380 -3900 102620 -3880
rect 102880 -3900 103120 -3880
rect 103380 -3900 103620 -3880
rect 103880 -3900 104120 -3880
rect 104380 -3900 104620 -3880
rect 104880 -3900 105120 -3880
rect 105380 -3900 105620 -3880
rect 105880 -3900 106120 -3880
rect 106380 -3900 106620 -3880
rect 106880 -3900 107120 -3880
rect 107380 -3900 107620 -3880
rect 107880 -3900 108120 -3880
rect 108380 -3900 108620 -3880
rect 108880 -3900 109120 -3880
rect 109380 -3900 109620 -3880
rect 109880 -3900 110120 -3880
rect 110380 -3900 110620 -3880
rect 110880 -3900 111120 -3880
rect 111380 -3900 111620 -3880
rect 111880 -3900 112120 -3880
rect 112380 -3900 112620 -3880
rect 112880 -3900 113120 -3880
rect 113380 -3900 113620 -3880
rect 113880 -3900 114120 -3880
rect 114380 -3900 114620 -3880
rect 114880 -3900 115120 -3880
rect 115380 -3900 115620 -3880
rect 115880 -3900 116120 -3880
rect 116380 -3900 116620 -3880
rect 116880 -3900 117120 -3880
rect 117380 -3900 117620 -3880
rect 117880 -3900 118120 -3880
rect 118380 -3900 118620 -3880
rect 118880 -3900 119120 -3880
rect 119380 -3900 119620 -3880
rect 119880 -3900 120120 -3880
rect 120380 -3900 120620 -3880
rect 120880 -3900 121120 -3880
rect 121380 -3900 121620 -3880
rect 121880 -3900 122120 -3880
rect 122380 -3900 122620 -3880
rect 122880 -3900 123120 -3880
rect 123380 -3900 123620 -3880
rect 123880 -3900 124120 -3880
rect 124380 -3900 124620 -3880
rect 124880 -3900 125120 -3880
rect 125380 -3900 125620 -3880
rect 125880 -3900 126120 -3880
rect 126380 -3900 126620 -3880
rect 126880 -3900 127120 -3880
rect 127380 -3900 127620 -3880
rect 127880 -3900 128120 -3880
rect 128380 -3900 128620 -3880
rect 128880 -3900 129120 -3880
rect 129380 -3900 129620 -3880
rect 129880 -3900 130120 -3880
rect 130380 -3900 130620 -3880
rect 130880 -3900 131120 -3880
rect 131380 -3900 131620 -3880
rect 131880 -3900 132120 -3880
rect 132380 -3900 132620 -3880
rect 132880 -3900 133120 -3880
rect 133380 -3900 133620 -3880
rect 133880 -3900 134120 -3880
rect 134380 -3900 134620 -3880
rect 134880 -3900 135120 -3880
rect 135380 -3900 135620 -3880
rect 135880 -3900 136120 -3880
rect 136380 -3900 136620 -3880
rect 136880 -3900 137120 -3880
rect 137380 -3900 137620 -3880
rect 137880 -3900 138120 -3880
rect 138380 -3900 138620 -3880
rect 138880 -3900 139120 -3880
rect 139380 -3900 139620 -3880
rect 139880 -3900 140000 -3880
rect 88000 -4100 140000 -3900
rect 88000 -4120 88120 -4100
rect 88380 -4120 88620 -4100
rect 88880 -4120 89120 -4100
rect 89380 -4120 89620 -4100
rect 89880 -4120 90120 -4100
rect 90380 -4120 90620 -4100
rect 90880 -4120 91120 -4100
rect 91380 -4120 91620 -4100
rect 91880 -4120 92120 -4100
rect 92380 -4120 92620 -4100
rect 92880 -4120 93120 -4100
rect 93380 -4120 93620 -4100
rect 93880 -4120 94120 -4100
rect 94380 -4120 94620 -4100
rect 94880 -4120 95120 -4100
rect 95380 -4120 95620 -4100
rect 95880 -4120 96120 -4100
rect 96380 -4120 96620 -4100
rect 96880 -4120 97120 -4100
rect 97380 -4120 97620 -4100
rect 97880 -4120 98120 -4100
rect 98380 -4120 98620 -4100
rect 98880 -4120 99120 -4100
rect 99380 -4120 99620 -4100
rect 99880 -4120 100120 -4100
rect 100380 -4120 100620 -4100
rect 100880 -4120 101120 -4100
rect 101380 -4120 101620 -4100
rect 101880 -4120 102120 -4100
rect 102380 -4120 102620 -4100
rect 102880 -4120 103120 -4100
rect 103380 -4120 103620 -4100
rect 103880 -4120 104120 -4100
rect 104380 -4120 104620 -4100
rect 104880 -4120 105120 -4100
rect 105380 -4120 105620 -4100
rect 105880 -4120 106120 -4100
rect 106380 -4120 106620 -4100
rect 106880 -4120 107120 -4100
rect 107380 -4120 107620 -4100
rect 107880 -4120 108120 -4100
rect 108380 -4120 108620 -4100
rect 108880 -4120 109120 -4100
rect 109380 -4120 109620 -4100
rect 109880 -4120 110120 -4100
rect 110380 -4120 110620 -4100
rect 110880 -4120 111120 -4100
rect 111380 -4120 111620 -4100
rect 111880 -4120 112120 -4100
rect 112380 -4120 112620 -4100
rect 112880 -4120 113120 -4100
rect 113380 -4120 113620 -4100
rect 113880 -4120 114120 -4100
rect 114380 -4120 114620 -4100
rect 114880 -4120 115120 -4100
rect 115380 -4120 115620 -4100
rect 115880 -4120 116120 -4100
rect 116380 -4120 116620 -4100
rect 116880 -4120 117120 -4100
rect 117380 -4120 117620 -4100
rect 117880 -4120 118120 -4100
rect 118380 -4120 118620 -4100
rect 118880 -4120 119120 -4100
rect 119380 -4120 119620 -4100
rect 119880 -4120 120120 -4100
rect 120380 -4120 120620 -4100
rect 120880 -4120 121120 -4100
rect 121380 -4120 121620 -4100
rect 121880 -4120 122120 -4100
rect 122380 -4120 122620 -4100
rect 122880 -4120 123120 -4100
rect 123380 -4120 123620 -4100
rect 123880 -4120 124120 -4100
rect 124380 -4120 124620 -4100
rect 124880 -4120 125120 -4100
rect 125380 -4120 125620 -4100
rect 125880 -4120 126120 -4100
rect 126380 -4120 126620 -4100
rect 126880 -4120 127120 -4100
rect 127380 -4120 127620 -4100
rect 127880 -4120 128120 -4100
rect 128380 -4120 128620 -4100
rect 128880 -4120 129120 -4100
rect 129380 -4120 129620 -4100
rect 129880 -4120 130120 -4100
rect 130380 -4120 130620 -4100
rect 130880 -4120 131120 -4100
rect 131380 -4120 131620 -4100
rect 131880 -4120 132120 -4100
rect 132380 -4120 132620 -4100
rect 132880 -4120 133120 -4100
rect 133380 -4120 133620 -4100
rect 133880 -4120 134120 -4100
rect 134380 -4120 134620 -4100
rect 134880 -4120 135120 -4100
rect 135380 -4120 135620 -4100
rect 135880 -4120 136120 -4100
rect 136380 -4120 136620 -4100
rect 136880 -4120 137120 -4100
rect 137380 -4120 137620 -4100
rect 137880 -4120 138120 -4100
rect 138380 -4120 138620 -4100
rect 138880 -4120 139120 -4100
rect 139380 -4120 139620 -4100
rect 139880 -4120 140000 -4100
rect 88000 -4380 88100 -4120
rect 88400 -4380 88600 -4120
rect 88900 -4380 89100 -4120
rect 89400 -4380 89600 -4120
rect 89900 -4380 90100 -4120
rect 90400 -4380 90600 -4120
rect 90900 -4380 91100 -4120
rect 91400 -4380 91600 -4120
rect 91900 -4380 92100 -4120
rect 92400 -4380 92600 -4120
rect 92900 -4380 93100 -4120
rect 93400 -4380 93600 -4120
rect 93900 -4380 94100 -4120
rect 94400 -4380 94600 -4120
rect 94900 -4380 95100 -4120
rect 95400 -4380 95600 -4120
rect 95900 -4380 96100 -4120
rect 96400 -4380 96600 -4120
rect 96900 -4380 97100 -4120
rect 97400 -4380 97600 -4120
rect 97900 -4380 98100 -4120
rect 98400 -4380 98600 -4120
rect 98900 -4380 99100 -4120
rect 99400 -4380 99600 -4120
rect 99900 -4380 100100 -4120
rect 100400 -4380 100600 -4120
rect 100900 -4380 101100 -4120
rect 101400 -4380 101600 -4120
rect 101900 -4380 102100 -4120
rect 102400 -4380 102600 -4120
rect 102900 -4380 103100 -4120
rect 103400 -4380 103600 -4120
rect 103900 -4380 104100 -4120
rect 104400 -4380 104600 -4120
rect 104900 -4380 105100 -4120
rect 105400 -4380 105600 -4120
rect 105900 -4380 106100 -4120
rect 106400 -4380 106600 -4120
rect 106900 -4380 107100 -4120
rect 107400 -4380 107600 -4120
rect 107900 -4380 108100 -4120
rect 108400 -4380 108600 -4120
rect 108900 -4380 109100 -4120
rect 109400 -4380 109600 -4120
rect 109900 -4380 110100 -4120
rect 110400 -4380 110600 -4120
rect 110900 -4380 111100 -4120
rect 111400 -4380 111600 -4120
rect 111900 -4380 112100 -4120
rect 112400 -4380 112600 -4120
rect 112900 -4380 113100 -4120
rect 113400 -4380 113600 -4120
rect 113900 -4380 114100 -4120
rect 114400 -4380 114600 -4120
rect 114900 -4380 115100 -4120
rect 115400 -4380 115600 -4120
rect 115900 -4380 116100 -4120
rect 116400 -4380 116600 -4120
rect 116900 -4380 117100 -4120
rect 117400 -4380 117600 -4120
rect 117900 -4380 118100 -4120
rect 118400 -4380 118600 -4120
rect 118900 -4380 119100 -4120
rect 119400 -4380 119600 -4120
rect 119900 -4380 120100 -4120
rect 120400 -4380 120600 -4120
rect 120900 -4380 121100 -4120
rect 121400 -4380 121600 -4120
rect 121900 -4380 122100 -4120
rect 122400 -4380 122600 -4120
rect 122900 -4380 123100 -4120
rect 123400 -4380 123600 -4120
rect 123900 -4380 124100 -4120
rect 124400 -4380 124600 -4120
rect 124900 -4380 125100 -4120
rect 125400 -4380 125600 -4120
rect 125900 -4380 126100 -4120
rect 126400 -4380 126600 -4120
rect 126900 -4380 127100 -4120
rect 127400 -4380 127600 -4120
rect 127900 -4380 128100 -4120
rect 128400 -4380 128600 -4120
rect 128900 -4380 129100 -4120
rect 129400 -4380 129600 -4120
rect 129900 -4380 130100 -4120
rect 130400 -4380 130600 -4120
rect 130900 -4380 131100 -4120
rect 131400 -4380 131600 -4120
rect 131900 -4380 132100 -4120
rect 132400 -4380 132600 -4120
rect 132900 -4380 133100 -4120
rect 133400 -4380 133600 -4120
rect 133900 -4380 134100 -4120
rect 134400 -4380 134600 -4120
rect 134900 -4380 135100 -4120
rect 135400 -4380 135600 -4120
rect 135900 -4380 136100 -4120
rect 136400 -4380 136600 -4120
rect 136900 -4380 137100 -4120
rect 137400 -4380 137600 -4120
rect 137900 -4380 138100 -4120
rect 138400 -4380 138600 -4120
rect 138900 -4380 139100 -4120
rect 139400 -4380 139600 -4120
rect 139900 -4380 140000 -4120
rect 88000 -4400 88120 -4380
rect 88380 -4400 88620 -4380
rect 88880 -4400 89120 -4380
rect 89380 -4400 89620 -4380
rect 89880 -4400 90120 -4380
rect 90380 -4400 90620 -4380
rect 90880 -4400 91120 -4380
rect 91380 -4400 91620 -4380
rect 91880 -4400 92120 -4380
rect 92380 -4400 92620 -4380
rect 92880 -4400 93120 -4380
rect 93380 -4400 93620 -4380
rect 93880 -4400 94120 -4380
rect 94380 -4400 94620 -4380
rect 94880 -4400 95120 -4380
rect 95380 -4400 95620 -4380
rect 95880 -4400 96120 -4380
rect 96380 -4400 96620 -4380
rect 96880 -4400 97120 -4380
rect 97380 -4400 97620 -4380
rect 97880 -4400 98120 -4380
rect 98380 -4400 98620 -4380
rect 98880 -4400 99120 -4380
rect 99380 -4400 99620 -4380
rect 99880 -4400 100120 -4380
rect 100380 -4400 100620 -4380
rect 100880 -4400 101120 -4380
rect 101380 -4400 101620 -4380
rect 101880 -4400 102120 -4380
rect 102380 -4400 102620 -4380
rect 102880 -4400 103120 -4380
rect 103380 -4400 103620 -4380
rect 103880 -4400 104120 -4380
rect 104380 -4400 104620 -4380
rect 104880 -4400 105120 -4380
rect 105380 -4400 105620 -4380
rect 105880 -4400 106120 -4380
rect 106380 -4400 106620 -4380
rect 106880 -4400 107120 -4380
rect 107380 -4400 107620 -4380
rect 107880 -4400 108120 -4380
rect 108380 -4400 108620 -4380
rect 108880 -4400 109120 -4380
rect 109380 -4400 109620 -4380
rect 109880 -4400 110120 -4380
rect 110380 -4400 110620 -4380
rect 110880 -4400 111120 -4380
rect 111380 -4400 111620 -4380
rect 111880 -4400 112120 -4380
rect 112380 -4400 112620 -4380
rect 112880 -4400 113120 -4380
rect 113380 -4400 113620 -4380
rect 113880 -4400 114120 -4380
rect 114380 -4400 114620 -4380
rect 114880 -4400 115120 -4380
rect 115380 -4400 115620 -4380
rect 115880 -4400 116120 -4380
rect 116380 -4400 116620 -4380
rect 116880 -4400 117120 -4380
rect 117380 -4400 117620 -4380
rect 117880 -4400 118120 -4380
rect 118380 -4400 118620 -4380
rect 118880 -4400 119120 -4380
rect 119380 -4400 119620 -4380
rect 119880 -4400 120120 -4380
rect 120380 -4400 120620 -4380
rect 120880 -4400 121120 -4380
rect 121380 -4400 121620 -4380
rect 121880 -4400 122120 -4380
rect 122380 -4400 122620 -4380
rect 122880 -4400 123120 -4380
rect 123380 -4400 123620 -4380
rect 123880 -4400 124120 -4380
rect 124380 -4400 124620 -4380
rect 124880 -4400 125120 -4380
rect 125380 -4400 125620 -4380
rect 125880 -4400 126120 -4380
rect 126380 -4400 126620 -4380
rect 126880 -4400 127120 -4380
rect 127380 -4400 127620 -4380
rect 127880 -4400 128120 -4380
rect 128380 -4400 128620 -4380
rect 128880 -4400 129120 -4380
rect 129380 -4400 129620 -4380
rect 129880 -4400 130120 -4380
rect 130380 -4400 130620 -4380
rect 130880 -4400 131120 -4380
rect 131380 -4400 131620 -4380
rect 131880 -4400 132120 -4380
rect 132380 -4400 132620 -4380
rect 132880 -4400 133120 -4380
rect 133380 -4400 133620 -4380
rect 133880 -4400 134120 -4380
rect 134380 -4400 134620 -4380
rect 134880 -4400 135120 -4380
rect 135380 -4400 135620 -4380
rect 135880 -4400 136120 -4380
rect 136380 -4400 136620 -4380
rect 136880 -4400 137120 -4380
rect 137380 -4400 137620 -4380
rect 137880 -4400 138120 -4380
rect 138380 -4400 138620 -4380
rect 138880 -4400 139120 -4380
rect 139380 -4400 139620 -4380
rect 139880 -4400 140000 -4380
rect 88000 -4600 140000 -4400
rect 88000 -4620 88120 -4600
rect 88380 -4620 88620 -4600
rect 88880 -4620 89120 -4600
rect 89380 -4620 89620 -4600
rect 89880 -4620 90120 -4600
rect 90380 -4620 90620 -4600
rect 90880 -4620 91120 -4600
rect 91380 -4620 91620 -4600
rect 91880 -4620 92120 -4600
rect 92380 -4620 92620 -4600
rect 92880 -4620 93120 -4600
rect 93380 -4620 93620 -4600
rect 93880 -4620 94120 -4600
rect 94380 -4620 94620 -4600
rect 94880 -4620 95120 -4600
rect 95380 -4620 95620 -4600
rect 95880 -4620 96120 -4600
rect 96380 -4620 96620 -4600
rect 96880 -4620 97120 -4600
rect 97380 -4620 97620 -4600
rect 97880 -4620 98120 -4600
rect 98380 -4620 98620 -4600
rect 98880 -4620 99120 -4600
rect 99380 -4620 99620 -4600
rect 99880 -4620 100120 -4600
rect 100380 -4620 100620 -4600
rect 100880 -4620 101120 -4600
rect 101380 -4620 101620 -4600
rect 101880 -4620 102120 -4600
rect 102380 -4620 102620 -4600
rect 102880 -4620 103120 -4600
rect 103380 -4620 103620 -4600
rect 103880 -4620 104120 -4600
rect 104380 -4620 104620 -4600
rect 104880 -4620 105120 -4600
rect 105380 -4620 105620 -4600
rect 105880 -4620 106120 -4600
rect 106380 -4620 106620 -4600
rect 106880 -4620 107120 -4600
rect 107380 -4620 107620 -4600
rect 107880 -4620 108120 -4600
rect 108380 -4620 108620 -4600
rect 108880 -4620 109120 -4600
rect 109380 -4620 109620 -4600
rect 109880 -4620 110120 -4600
rect 110380 -4620 110620 -4600
rect 110880 -4620 111120 -4600
rect 111380 -4620 111620 -4600
rect 111880 -4620 112120 -4600
rect 112380 -4620 112620 -4600
rect 112880 -4620 113120 -4600
rect 113380 -4620 113620 -4600
rect 113880 -4620 114120 -4600
rect 114380 -4620 114620 -4600
rect 114880 -4620 115120 -4600
rect 115380 -4620 115620 -4600
rect 115880 -4620 116120 -4600
rect 116380 -4620 116620 -4600
rect 116880 -4620 117120 -4600
rect 117380 -4620 117620 -4600
rect 117880 -4620 118120 -4600
rect 118380 -4620 118620 -4600
rect 118880 -4620 119120 -4600
rect 119380 -4620 119620 -4600
rect 119880 -4620 120120 -4600
rect 120380 -4620 120620 -4600
rect 120880 -4620 121120 -4600
rect 121380 -4620 121620 -4600
rect 121880 -4620 122120 -4600
rect 122380 -4620 122620 -4600
rect 122880 -4620 123120 -4600
rect 123380 -4620 123620 -4600
rect 123880 -4620 124120 -4600
rect 124380 -4620 124620 -4600
rect 124880 -4620 125120 -4600
rect 125380 -4620 125620 -4600
rect 125880 -4620 126120 -4600
rect 126380 -4620 126620 -4600
rect 126880 -4620 127120 -4600
rect 127380 -4620 127620 -4600
rect 127880 -4620 128120 -4600
rect 128380 -4620 128620 -4600
rect 128880 -4620 129120 -4600
rect 129380 -4620 129620 -4600
rect 129880 -4620 130120 -4600
rect 130380 -4620 130620 -4600
rect 130880 -4620 131120 -4600
rect 131380 -4620 131620 -4600
rect 131880 -4620 132120 -4600
rect 132380 -4620 132620 -4600
rect 132880 -4620 133120 -4600
rect 133380 -4620 133620 -4600
rect 133880 -4620 134120 -4600
rect 134380 -4620 134620 -4600
rect 134880 -4620 135120 -4600
rect 135380 -4620 135620 -4600
rect 135880 -4620 136120 -4600
rect 136380 -4620 136620 -4600
rect 136880 -4620 137120 -4600
rect 137380 -4620 137620 -4600
rect 137880 -4620 138120 -4600
rect 138380 -4620 138620 -4600
rect 138880 -4620 139120 -4600
rect 139380 -4620 139620 -4600
rect 139880 -4620 140000 -4600
rect 88000 -4880 88100 -4620
rect 88400 -4880 88600 -4620
rect 88900 -4880 89100 -4620
rect 89400 -4880 89600 -4620
rect 89900 -4880 90100 -4620
rect 90400 -4880 90600 -4620
rect 90900 -4880 91100 -4620
rect 91400 -4880 91600 -4620
rect 91900 -4880 92100 -4620
rect 92400 -4880 92600 -4620
rect 92900 -4880 93100 -4620
rect 93400 -4880 93600 -4620
rect 93900 -4880 94100 -4620
rect 94400 -4880 94600 -4620
rect 94900 -4880 95100 -4620
rect 95400 -4880 95600 -4620
rect 95900 -4880 96100 -4620
rect 96400 -4880 96600 -4620
rect 96900 -4880 97100 -4620
rect 97400 -4880 97600 -4620
rect 97900 -4880 98100 -4620
rect 98400 -4880 98600 -4620
rect 98900 -4880 99100 -4620
rect 99400 -4880 99600 -4620
rect 99900 -4880 100100 -4620
rect 100400 -4880 100600 -4620
rect 100900 -4880 101100 -4620
rect 101400 -4880 101600 -4620
rect 101900 -4880 102100 -4620
rect 102400 -4880 102600 -4620
rect 102900 -4880 103100 -4620
rect 103400 -4880 103600 -4620
rect 103900 -4880 104100 -4620
rect 104400 -4880 104600 -4620
rect 104900 -4880 105100 -4620
rect 105400 -4880 105600 -4620
rect 105900 -4880 106100 -4620
rect 106400 -4880 106600 -4620
rect 106900 -4880 107100 -4620
rect 107400 -4880 107600 -4620
rect 107900 -4880 108100 -4620
rect 108400 -4880 108600 -4620
rect 108900 -4880 109100 -4620
rect 109400 -4880 109600 -4620
rect 109900 -4880 110100 -4620
rect 110400 -4880 110600 -4620
rect 110900 -4880 111100 -4620
rect 111400 -4880 111600 -4620
rect 111900 -4880 112100 -4620
rect 112400 -4880 112600 -4620
rect 112900 -4880 113100 -4620
rect 113400 -4880 113600 -4620
rect 113900 -4880 114100 -4620
rect 114400 -4880 114600 -4620
rect 114900 -4880 115100 -4620
rect 115400 -4880 115600 -4620
rect 115900 -4880 116100 -4620
rect 116400 -4880 116600 -4620
rect 116900 -4880 117100 -4620
rect 117400 -4880 117600 -4620
rect 117900 -4880 118100 -4620
rect 118400 -4880 118600 -4620
rect 118900 -4880 119100 -4620
rect 119400 -4880 119600 -4620
rect 119900 -4880 120100 -4620
rect 120400 -4880 120600 -4620
rect 120900 -4880 121100 -4620
rect 121400 -4880 121600 -4620
rect 121900 -4880 122100 -4620
rect 122400 -4880 122600 -4620
rect 122900 -4880 123100 -4620
rect 123400 -4880 123600 -4620
rect 123900 -4880 124100 -4620
rect 124400 -4880 124600 -4620
rect 124900 -4880 125100 -4620
rect 125400 -4880 125600 -4620
rect 125900 -4880 126100 -4620
rect 126400 -4880 126600 -4620
rect 126900 -4880 127100 -4620
rect 127400 -4880 127600 -4620
rect 127900 -4880 128100 -4620
rect 128400 -4880 128600 -4620
rect 128900 -4880 129100 -4620
rect 129400 -4880 129600 -4620
rect 129900 -4880 130100 -4620
rect 130400 -4880 130600 -4620
rect 130900 -4880 131100 -4620
rect 131400 -4880 131600 -4620
rect 131900 -4880 132100 -4620
rect 132400 -4880 132600 -4620
rect 132900 -4880 133100 -4620
rect 133400 -4880 133600 -4620
rect 133900 -4880 134100 -4620
rect 134400 -4880 134600 -4620
rect 134900 -4880 135100 -4620
rect 135400 -4880 135600 -4620
rect 135900 -4880 136100 -4620
rect 136400 -4880 136600 -4620
rect 136900 -4880 137100 -4620
rect 137400 -4880 137600 -4620
rect 137900 -4880 138100 -4620
rect 138400 -4880 138600 -4620
rect 138900 -4880 139100 -4620
rect 139400 -4880 139600 -4620
rect 139900 -4880 140000 -4620
rect 88000 -4900 88120 -4880
rect 88380 -4900 88620 -4880
rect 88880 -4900 89120 -4880
rect 89380 -4900 89620 -4880
rect 89880 -4900 90120 -4880
rect 90380 -4900 90620 -4880
rect 90880 -4900 91120 -4880
rect 91380 -4900 91620 -4880
rect 91880 -4900 92120 -4880
rect 92380 -4900 92620 -4880
rect 92880 -4900 93120 -4880
rect 93380 -4900 93620 -4880
rect 93880 -4900 94120 -4880
rect 94380 -4900 94620 -4880
rect 94880 -4900 95120 -4880
rect 95380 -4900 95620 -4880
rect 95880 -4900 96120 -4880
rect 96380 -4900 96620 -4880
rect 96880 -4900 97120 -4880
rect 97380 -4900 97620 -4880
rect 97880 -4900 98120 -4880
rect 98380 -4900 98620 -4880
rect 98880 -4900 99120 -4880
rect 99380 -4900 99620 -4880
rect 99880 -4900 100120 -4880
rect 100380 -4900 100620 -4880
rect 100880 -4900 101120 -4880
rect 101380 -4900 101620 -4880
rect 101880 -4900 102120 -4880
rect 102380 -4900 102620 -4880
rect 102880 -4900 103120 -4880
rect 103380 -4900 103620 -4880
rect 103880 -4900 104120 -4880
rect 104380 -4900 104620 -4880
rect 104880 -4900 105120 -4880
rect 105380 -4900 105620 -4880
rect 105880 -4900 106120 -4880
rect 106380 -4900 106620 -4880
rect 106880 -4900 107120 -4880
rect 107380 -4900 107620 -4880
rect 107880 -4900 108120 -4880
rect 108380 -4900 108620 -4880
rect 108880 -4900 109120 -4880
rect 109380 -4900 109620 -4880
rect 109880 -4900 110120 -4880
rect 110380 -4900 110620 -4880
rect 110880 -4900 111120 -4880
rect 111380 -4900 111620 -4880
rect 111880 -4900 112120 -4880
rect 112380 -4900 112620 -4880
rect 112880 -4900 113120 -4880
rect 113380 -4900 113620 -4880
rect 113880 -4900 114120 -4880
rect 114380 -4900 114620 -4880
rect 114880 -4900 115120 -4880
rect 115380 -4900 115620 -4880
rect 115880 -4900 116120 -4880
rect 116380 -4900 116620 -4880
rect 116880 -4900 117120 -4880
rect 117380 -4900 117620 -4880
rect 117880 -4900 118120 -4880
rect 118380 -4900 118620 -4880
rect 118880 -4900 119120 -4880
rect 119380 -4900 119620 -4880
rect 119880 -4900 120120 -4880
rect 120380 -4900 120620 -4880
rect 120880 -4900 121120 -4880
rect 121380 -4900 121620 -4880
rect 121880 -4900 122120 -4880
rect 122380 -4900 122620 -4880
rect 122880 -4900 123120 -4880
rect 123380 -4900 123620 -4880
rect 123880 -4900 124120 -4880
rect 124380 -4900 124620 -4880
rect 124880 -4900 125120 -4880
rect 125380 -4900 125620 -4880
rect 125880 -4900 126120 -4880
rect 126380 -4900 126620 -4880
rect 126880 -4900 127120 -4880
rect 127380 -4900 127620 -4880
rect 127880 -4900 128120 -4880
rect 128380 -4900 128620 -4880
rect 128880 -4900 129120 -4880
rect 129380 -4900 129620 -4880
rect 129880 -4900 130120 -4880
rect 130380 -4900 130620 -4880
rect 130880 -4900 131120 -4880
rect 131380 -4900 131620 -4880
rect 131880 -4900 132120 -4880
rect 132380 -4900 132620 -4880
rect 132880 -4900 133120 -4880
rect 133380 -4900 133620 -4880
rect 133880 -4900 134120 -4880
rect 134380 -4900 134620 -4880
rect 134880 -4900 135120 -4880
rect 135380 -4900 135620 -4880
rect 135880 -4900 136120 -4880
rect 136380 -4900 136620 -4880
rect 136880 -4900 137120 -4880
rect 137380 -4900 137620 -4880
rect 137880 -4900 138120 -4880
rect 138380 -4900 138620 -4880
rect 138880 -4900 139120 -4880
rect 139380 -4900 139620 -4880
rect 139880 -4900 140000 -4880
rect 88000 -5100 140000 -4900
rect 88000 -5120 88120 -5100
rect 88380 -5120 88620 -5100
rect 88880 -5120 89120 -5100
rect 89380 -5120 89620 -5100
rect 89880 -5120 90120 -5100
rect 90380 -5120 90620 -5100
rect 90880 -5120 91120 -5100
rect 91380 -5120 91620 -5100
rect 91880 -5120 92120 -5100
rect 92380 -5120 92620 -5100
rect 92880 -5120 93120 -5100
rect 93380 -5120 93620 -5100
rect 93880 -5120 94120 -5100
rect 94380 -5120 94620 -5100
rect 94880 -5120 95120 -5100
rect 95380 -5120 95620 -5100
rect 95880 -5120 96120 -5100
rect 96380 -5120 96620 -5100
rect 96880 -5120 97120 -5100
rect 97380 -5120 97620 -5100
rect 97880 -5120 98120 -5100
rect 98380 -5120 98620 -5100
rect 98880 -5120 99120 -5100
rect 99380 -5120 99620 -5100
rect 99880 -5120 100120 -5100
rect 100380 -5120 100620 -5100
rect 100880 -5120 101120 -5100
rect 101380 -5120 101620 -5100
rect 101880 -5120 102120 -5100
rect 102380 -5120 102620 -5100
rect 102880 -5120 103120 -5100
rect 103380 -5120 103620 -5100
rect 103880 -5120 104120 -5100
rect 104380 -5120 104620 -5100
rect 104880 -5120 105120 -5100
rect 105380 -5120 105620 -5100
rect 105880 -5120 106120 -5100
rect 106380 -5120 106620 -5100
rect 106880 -5120 107120 -5100
rect 107380 -5120 107620 -5100
rect 107880 -5120 108120 -5100
rect 108380 -5120 108620 -5100
rect 108880 -5120 109120 -5100
rect 109380 -5120 109620 -5100
rect 109880 -5120 110120 -5100
rect 110380 -5120 110620 -5100
rect 110880 -5120 111120 -5100
rect 111380 -5120 111620 -5100
rect 111880 -5120 112120 -5100
rect 112380 -5120 112620 -5100
rect 112880 -5120 113120 -5100
rect 113380 -5120 113620 -5100
rect 113880 -5120 114120 -5100
rect 114380 -5120 114620 -5100
rect 114880 -5120 115120 -5100
rect 115380 -5120 115620 -5100
rect 115880 -5120 116120 -5100
rect 116380 -5120 116620 -5100
rect 116880 -5120 117120 -5100
rect 117380 -5120 117620 -5100
rect 117880 -5120 118120 -5100
rect 118380 -5120 118620 -5100
rect 118880 -5120 119120 -5100
rect 119380 -5120 119620 -5100
rect 119880 -5120 120120 -5100
rect 120380 -5120 120620 -5100
rect 120880 -5120 121120 -5100
rect 121380 -5120 121620 -5100
rect 121880 -5120 122120 -5100
rect 122380 -5120 122620 -5100
rect 122880 -5120 123120 -5100
rect 123380 -5120 123620 -5100
rect 123880 -5120 124120 -5100
rect 124380 -5120 124620 -5100
rect 124880 -5120 125120 -5100
rect 125380 -5120 125620 -5100
rect 125880 -5120 126120 -5100
rect 126380 -5120 126620 -5100
rect 126880 -5120 127120 -5100
rect 127380 -5120 127620 -5100
rect 127880 -5120 128120 -5100
rect 128380 -5120 128620 -5100
rect 128880 -5120 129120 -5100
rect 129380 -5120 129620 -5100
rect 129880 -5120 130120 -5100
rect 130380 -5120 130620 -5100
rect 130880 -5120 131120 -5100
rect 131380 -5120 131620 -5100
rect 131880 -5120 132120 -5100
rect 132380 -5120 132620 -5100
rect 132880 -5120 133120 -5100
rect 133380 -5120 133620 -5100
rect 133880 -5120 134120 -5100
rect 134380 -5120 134620 -5100
rect 134880 -5120 135120 -5100
rect 135380 -5120 135620 -5100
rect 135880 -5120 136120 -5100
rect 136380 -5120 136620 -5100
rect 136880 -5120 137120 -5100
rect 137380 -5120 137620 -5100
rect 137880 -5120 138120 -5100
rect 138380 -5120 138620 -5100
rect 138880 -5120 139120 -5100
rect 139380 -5120 139620 -5100
rect 139880 -5120 140000 -5100
rect 88000 -5380 88100 -5120
rect 88400 -5380 88600 -5120
rect 88900 -5380 89100 -5120
rect 89400 -5380 89600 -5120
rect 89900 -5380 90100 -5120
rect 90400 -5380 90600 -5120
rect 90900 -5380 91100 -5120
rect 91400 -5380 91600 -5120
rect 91900 -5380 92100 -5120
rect 92400 -5380 92600 -5120
rect 92900 -5380 93100 -5120
rect 93400 -5380 93600 -5120
rect 93900 -5380 94100 -5120
rect 94400 -5380 94600 -5120
rect 94900 -5380 95100 -5120
rect 95400 -5380 95600 -5120
rect 95900 -5380 96100 -5120
rect 96400 -5380 96600 -5120
rect 96900 -5380 97100 -5120
rect 97400 -5380 97600 -5120
rect 97900 -5380 98100 -5120
rect 98400 -5380 98600 -5120
rect 98900 -5380 99100 -5120
rect 99400 -5380 99600 -5120
rect 99900 -5380 100100 -5120
rect 100400 -5380 100600 -5120
rect 100900 -5380 101100 -5120
rect 101400 -5380 101600 -5120
rect 101900 -5380 102100 -5120
rect 102400 -5380 102600 -5120
rect 102900 -5380 103100 -5120
rect 103400 -5380 103600 -5120
rect 103900 -5380 104100 -5120
rect 104400 -5380 104600 -5120
rect 104900 -5380 105100 -5120
rect 105400 -5380 105600 -5120
rect 105900 -5380 106100 -5120
rect 106400 -5380 106600 -5120
rect 106900 -5380 107100 -5120
rect 107400 -5380 107600 -5120
rect 107900 -5380 108100 -5120
rect 108400 -5380 108600 -5120
rect 108900 -5380 109100 -5120
rect 109400 -5380 109600 -5120
rect 109900 -5380 110100 -5120
rect 110400 -5380 110600 -5120
rect 110900 -5380 111100 -5120
rect 111400 -5380 111600 -5120
rect 111900 -5380 112100 -5120
rect 112400 -5380 112600 -5120
rect 112900 -5380 113100 -5120
rect 113400 -5380 113600 -5120
rect 113900 -5380 114100 -5120
rect 114400 -5380 114600 -5120
rect 114900 -5380 115100 -5120
rect 115400 -5380 115600 -5120
rect 115900 -5380 116100 -5120
rect 116400 -5380 116600 -5120
rect 116900 -5380 117100 -5120
rect 117400 -5380 117600 -5120
rect 117900 -5380 118100 -5120
rect 118400 -5380 118600 -5120
rect 118900 -5380 119100 -5120
rect 119400 -5380 119600 -5120
rect 119900 -5380 120100 -5120
rect 120400 -5380 120600 -5120
rect 120900 -5380 121100 -5120
rect 121400 -5380 121600 -5120
rect 121900 -5380 122100 -5120
rect 122400 -5380 122600 -5120
rect 122900 -5380 123100 -5120
rect 123400 -5380 123600 -5120
rect 123900 -5380 124100 -5120
rect 124400 -5380 124600 -5120
rect 124900 -5380 125100 -5120
rect 125400 -5380 125600 -5120
rect 125900 -5380 126100 -5120
rect 126400 -5380 126600 -5120
rect 126900 -5380 127100 -5120
rect 127400 -5380 127600 -5120
rect 127900 -5380 128100 -5120
rect 128400 -5380 128600 -5120
rect 128900 -5380 129100 -5120
rect 129400 -5380 129600 -5120
rect 129900 -5380 130100 -5120
rect 130400 -5380 130600 -5120
rect 130900 -5380 131100 -5120
rect 131400 -5380 131600 -5120
rect 131900 -5380 132100 -5120
rect 132400 -5380 132600 -5120
rect 132900 -5380 133100 -5120
rect 133400 -5380 133600 -5120
rect 133900 -5380 134100 -5120
rect 134400 -5380 134600 -5120
rect 134900 -5380 135100 -5120
rect 135400 -5380 135600 -5120
rect 135900 -5380 136100 -5120
rect 136400 -5380 136600 -5120
rect 136900 -5380 137100 -5120
rect 137400 -5380 137600 -5120
rect 137900 -5380 138100 -5120
rect 138400 -5380 138600 -5120
rect 138900 -5380 139100 -5120
rect 139400 -5380 139600 -5120
rect 139900 -5380 140000 -5120
rect 88000 -5400 88120 -5380
rect 88380 -5400 88620 -5380
rect 88880 -5400 89120 -5380
rect 89380 -5400 89620 -5380
rect 89880 -5400 90120 -5380
rect 90380 -5400 90620 -5380
rect 90880 -5400 91120 -5380
rect 91380 -5400 91620 -5380
rect 91880 -5400 92120 -5380
rect 92380 -5400 92620 -5380
rect 92880 -5400 93120 -5380
rect 93380 -5400 93620 -5380
rect 93880 -5400 94120 -5380
rect 94380 -5400 94620 -5380
rect 94880 -5400 95120 -5380
rect 95380 -5400 95620 -5380
rect 95880 -5400 96120 -5380
rect 96380 -5400 96620 -5380
rect 96880 -5400 97120 -5380
rect 97380 -5400 97620 -5380
rect 97880 -5400 98120 -5380
rect 98380 -5400 98620 -5380
rect 98880 -5400 99120 -5380
rect 99380 -5400 99620 -5380
rect 99880 -5400 100120 -5380
rect 100380 -5400 100620 -5380
rect 100880 -5400 101120 -5380
rect 101380 -5400 101620 -5380
rect 101880 -5400 102120 -5380
rect 102380 -5400 102620 -5380
rect 102880 -5400 103120 -5380
rect 103380 -5400 103620 -5380
rect 103880 -5400 104120 -5380
rect 104380 -5400 104620 -5380
rect 104880 -5400 105120 -5380
rect 105380 -5400 105620 -5380
rect 105880 -5400 106120 -5380
rect 106380 -5400 106620 -5380
rect 106880 -5400 107120 -5380
rect 107380 -5400 107620 -5380
rect 107880 -5400 108120 -5380
rect 108380 -5400 108620 -5380
rect 108880 -5400 109120 -5380
rect 109380 -5400 109620 -5380
rect 109880 -5400 110120 -5380
rect 110380 -5400 110620 -5380
rect 110880 -5400 111120 -5380
rect 111380 -5400 111620 -5380
rect 111880 -5400 112120 -5380
rect 112380 -5400 112620 -5380
rect 112880 -5400 113120 -5380
rect 113380 -5400 113620 -5380
rect 113880 -5400 114120 -5380
rect 114380 -5400 114620 -5380
rect 114880 -5400 115120 -5380
rect 115380 -5400 115620 -5380
rect 115880 -5400 116120 -5380
rect 116380 -5400 116620 -5380
rect 116880 -5400 117120 -5380
rect 117380 -5400 117620 -5380
rect 117880 -5400 118120 -5380
rect 118380 -5400 118620 -5380
rect 118880 -5400 119120 -5380
rect 119380 -5400 119620 -5380
rect 119880 -5400 120120 -5380
rect 120380 -5400 120620 -5380
rect 120880 -5400 121120 -5380
rect 121380 -5400 121620 -5380
rect 121880 -5400 122120 -5380
rect 122380 -5400 122620 -5380
rect 122880 -5400 123120 -5380
rect 123380 -5400 123620 -5380
rect 123880 -5400 124120 -5380
rect 124380 -5400 124620 -5380
rect 124880 -5400 125120 -5380
rect 125380 -5400 125620 -5380
rect 125880 -5400 126120 -5380
rect 126380 -5400 126620 -5380
rect 126880 -5400 127120 -5380
rect 127380 -5400 127620 -5380
rect 127880 -5400 128120 -5380
rect 128380 -5400 128620 -5380
rect 128880 -5400 129120 -5380
rect 129380 -5400 129620 -5380
rect 129880 -5400 130120 -5380
rect 130380 -5400 130620 -5380
rect 130880 -5400 131120 -5380
rect 131380 -5400 131620 -5380
rect 131880 -5400 132120 -5380
rect 132380 -5400 132620 -5380
rect 132880 -5400 133120 -5380
rect 133380 -5400 133620 -5380
rect 133880 -5400 134120 -5380
rect 134380 -5400 134620 -5380
rect 134880 -5400 135120 -5380
rect 135380 -5400 135620 -5380
rect 135880 -5400 136120 -5380
rect 136380 -5400 136620 -5380
rect 136880 -5400 137120 -5380
rect 137380 -5400 137620 -5380
rect 137880 -5400 138120 -5380
rect 138380 -5400 138620 -5380
rect 138880 -5400 139120 -5380
rect 139380 -5400 139620 -5380
rect 139880 -5400 140000 -5380
rect 88000 -5600 140000 -5400
rect 88000 -5620 88120 -5600
rect 88380 -5620 88620 -5600
rect 88880 -5620 89120 -5600
rect 89380 -5620 89620 -5600
rect 89880 -5620 90120 -5600
rect 90380 -5620 90620 -5600
rect 90880 -5620 91120 -5600
rect 91380 -5620 91620 -5600
rect 91880 -5620 92120 -5600
rect 92380 -5620 92620 -5600
rect 92880 -5620 93120 -5600
rect 93380 -5620 93620 -5600
rect 93880 -5620 94120 -5600
rect 94380 -5620 94620 -5600
rect 94880 -5620 95120 -5600
rect 95380 -5620 95620 -5600
rect 95880 -5620 96120 -5600
rect 96380 -5620 96620 -5600
rect 96880 -5620 97120 -5600
rect 97380 -5620 97620 -5600
rect 97880 -5620 98120 -5600
rect 98380 -5620 98620 -5600
rect 98880 -5620 99120 -5600
rect 99380 -5620 99620 -5600
rect 99880 -5620 100120 -5600
rect 100380 -5620 100620 -5600
rect 100880 -5620 101120 -5600
rect 101380 -5620 101620 -5600
rect 101880 -5620 102120 -5600
rect 102380 -5620 102620 -5600
rect 102880 -5620 103120 -5600
rect 103380 -5620 103620 -5600
rect 103880 -5620 104120 -5600
rect 104380 -5620 104620 -5600
rect 104880 -5620 105120 -5600
rect 105380 -5620 105620 -5600
rect 105880 -5620 106120 -5600
rect 106380 -5620 106620 -5600
rect 106880 -5620 107120 -5600
rect 107380 -5620 107620 -5600
rect 107880 -5620 108120 -5600
rect 108380 -5620 108620 -5600
rect 108880 -5620 109120 -5600
rect 109380 -5620 109620 -5600
rect 109880 -5620 110120 -5600
rect 110380 -5620 110620 -5600
rect 110880 -5620 111120 -5600
rect 111380 -5620 111620 -5600
rect 111880 -5620 112120 -5600
rect 112380 -5620 112620 -5600
rect 112880 -5620 113120 -5600
rect 113380 -5620 113620 -5600
rect 113880 -5620 114120 -5600
rect 114380 -5620 114620 -5600
rect 114880 -5620 115120 -5600
rect 115380 -5620 115620 -5600
rect 115880 -5620 116120 -5600
rect 116380 -5620 116620 -5600
rect 116880 -5620 117120 -5600
rect 117380 -5620 117620 -5600
rect 117880 -5620 118120 -5600
rect 118380 -5620 118620 -5600
rect 118880 -5620 119120 -5600
rect 119380 -5620 119620 -5600
rect 119880 -5620 120120 -5600
rect 120380 -5620 120620 -5600
rect 120880 -5620 121120 -5600
rect 121380 -5620 121620 -5600
rect 121880 -5620 122120 -5600
rect 122380 -5620 122620 -5600
rect 122880 -5620 123120 -5600
rect 123380 -5620 123620 -5600
rect 123880 -5620 124120 -5600
rect 124380 -5620 124620 -5600
rect 124880 -5620 125120 -5600
rect 125380 -5620 125620 -5600
rect 125880 -5620 126120 -5600
rect 126380 -5620 126620 -5600
rect 126880 -5620 127120 -5600
rect 127380 -5620 127620 -5600
rect 127880 -5620 128120 -5600
rect 128380 -5620 128620 -5600
rect 128880 -5620 129120 -5600
rect 129380 -5620 129620 -5600
rect 129880 -5620 130120 -5600
rect 130380 -5620 130620 -5600
rect 130880 -5620 131120 -5600
rect 131380 -5620 131620 -5600
rect 131880 -5620 132120 -5600
rect 132380 -5620 132620 -5600
rect 132880 -5620 133120 -5600
rect 133380 -5620 133620 -5600
rect 133880 -5620 134120 -5600
rect 134380 -5620 134620 -5600
rect 134880 -5620 135120 -5600
rect 135380 -5620 135620 -5600
rect 135880 -5620 136120 -5600
rect 136380 -5620 136620 -5600
rect 136880 -5620 137120 -5600
rect 137380 -5620 137620 -5600
rect 137880 -5620 138120 -5600
rect 138380 -5620 138620 -5600
rect 138880 -5620 139120 -5600
rect 139380 -5620 139620 -5600
rect 139880 -5620 140000 -5600
rect 88000 -5880 88100 -5620
rect 88400 -5880 88600 -5620
rect 88900 -5880 89100 -5620
rect 89400 -5880 89600 -5620
rect 89900 -5880 90100 -5620
rect 90400 -5880 90600 -5620
rect 90900 -5880 91100 -5620
rect 91400 -5880 91600 -5620
rect 91900 -5880 92100 -5620
rect 92400 -5880 92600 -5620
rect 92900 -5880 93100 -5620
rect 93400 -5880 93600 -5620
rect 93900 -5880 94100 -5620
rect 94400 -5880 94600 -5620
rect 94900 -5880 95100 -5620
rect 95400 -5880 95600 -5620
rect 95900 -5880 96100 -5620
rect 96400 -5880 96600 -5620
rect 96900 -5880 97100 -5620
rect 97400 -5880 97600 -5620
rect 97900 -5880 98100 -5620
rect 98400 -5880 98600 -5620
rect 98900 -5880 99100 -5620
rect 99400 -5880 99600 -5620
rect 99900 -5880 100100 -5620
rect 100400 -5880 100600 -5620
rect 100900 -5880 101100 -5620
rect 101400 -5880 101600 -5620
rect 101900 -5880 102100 -5620
rect 102400 -5880 102600 -5620
rect 102900 -5880 103100 -5620
rect 103400 -5880 103600 -5620
rect 103900 -5880 104100 -5620
rect 104400 -5880 104600 -5620
rect 104900 -5880 105100 -5620
rect 105400 -5880 105600 -5620
rect 105900 -5880 106100 -5620
rect 106400 -5880 106600 -5620
rect 106900 -5880 107100 -5620
rect 107400 -5880 107600 -5620
rect 107900 -5880 108100 -5620
rect 108400 -5880 108600 -5620
rect 108900 -5880 109100 -5620
rect 109400 -5880 109600 -5620
rect 109900 -5880 110100 -5620
rect 110400 -5880 110600 -5620
rect 110900 -5880 111100 -5620
rect 111400 -5880 111600 -5620
rect 111900 -5880 112100 -5620
rect 112400 -5880 112600 -5620
rect 112900 -5880 113100 -5620
rect 113400 -5880 113600 -5620
rect 113900 -5880 114100 -5620
rect 114400 -5880 114600 -5620
rect 114900 -5880 115100 -5620
rect 115400 -5880 115600 -5620
rect 115900 -5880 116100 -5620
rect 116400 -5880 116600 -5620
rect 116900 -5880 117100 -5620
rect 117400 -5880 117600 -5620
rect 117900 -5880 118100 -5620
rect 118400 -5880 118600 -5620
rect 118900 -5880 119100 -5620
rect 119400 -5880 119600 -5620
rect 119900 -5880 120100 -5620
rect 120400 -5880 120600 -5620
rect 120900 -5880 121100 -5620
rect 121400 -5880 121600 -5620
rect 121900 -5880 122100 -5620
rect 122400 -5880 122600 -5620
rect 122900 -5880 123100 -5620
rect 123400 -5880 123600 -5620
rect 123900 -5880 124100 -5620
rect 124400 -5880 124600 -5620
rect 124900 -5880 125100 -5620
rect 125400 -5880 125600 -5620
rect 125900 -5880 126100 -5620
rect 126400 -5880 126600 -5620
rect 126900 -5880 127100 -5620
rect 127400 -5880 127600 -5620
rect 127900 -5880 128100 -5620
rect 128400 -5880 128600 -5620
rect 128900 -5880 129100 -5620
rect 129400 -5880 129600 -5620
rect 129900 -5880 130100 -5620
rect 130400 -5880 130600 -5620
rect 130900 -5880 131100 -5620
rect 131400 -5880 131600 -5620
rect 131900 -5880 132100 -5620
rect 132400 -5880 132600 -5620
rect 132900 -5880 133100 -5620
rect 133400 -5880 133600 -5620
rect 133900 -5880 134100 -5620
rect 134400 -5880 134600 -5620
rect 134900 -5880 135100 -5620
rect 135400 -5880 135600 -5620
rect 135900 -5880 136100 -5620
rect 136400 -5880 136600 -5620
rect 136900 -5880 137100 -5620
rect 137400 -5880 137600 -5620
rect 137900 -5880 138100 -5620
rect 138400 -5880 138600 -5620
rect 138900 -5880 139100 -5620
rect 139400 -5880 139600 -5620
rect 139900 -5880 140000 -5620
rect 88000 -5900 88120 -5880
rect 88380 -5900 88620 -5880
rect 88880 -5900 89120 -5880
rect 89380 -5900 89620 -5880
rect 89880 -5900 90120 -5880
rect 90380 -5900 90620 -5880
rect 90880 -5900 91120 -5880
rect 91380 -5900 91620 -5880
rect 91880 -5900 92120 -5880
rect 92380 -5900 92620 -5880
rect 92880 -5900 93120 -5880
rect 93380 -5900 93620 -5880
rect 93880 -5900 94120 -5880
rect 94380 -5900 94620 -5880
rect 94880 -5900 95120 -5880
rect 95380 -5900 95620 -5880
rect 95880 -5900 96120 -5880
rect 96380 -5900 96620 -5880
rect 96880 -5900 97120 -5880
rect 97380 -5900 97620 -5880
rect 97880 -5900 98120 -5880
rect 98380 -5900 98620 -5880
rect 98880 -5900 99120 -5880
rect 99380 -5900 99620 -5880
rect 99880 -5900 100120 -5880
rect 100380 -5900 100620 -5880
rect 100880 -5900 101120 -5880
rect 101380 -5900 101620 -5880
rect 101880 -5900 102120 -5880
rect 102380 -5900 102620 -5880
rect 102880 -5900 103120 -5880
rect 103380 -5900 103620 -5880
rect 103880 -5900 104120 -5880
rect 104380 -5900 104620 -5880
rect 104880 -5900 105120 -5880
rect 105380 -5900 105620 -5880
rect 105880 -5900 106120 -5880
rect 106380 -5900 106620 -5880
rect 106880 -5900 107120 -5880
rect 107380 -5900 107620 -5880
rect 107880 -5900 108120 -5880
rect 108380 -5900 108620 -5880
rect 108880 -5900 109120 -5880
rect 109380 -5900 109620 -5880
rect 109880 -5900 110120 -5880
rect 110380 -5900 110620 -5880
rect 110880 -5900 111120 -5880
rect 111380 -5900 111620 -5880
rect 111880 -5900 112120 -5880
rect 112380 -5900 112620 -5880
rect 112880 -5900 113120 -5880
rect 113380 -5900 113620 -5880
rect 113880 -5900 114120 -5880
rect 114380 -5900 114620 -5880
rect 114880 -5900 115120 -5880
rect 115380 -5900 115620 -5880
rect 115880 -5900 116120 -5880
rect 116380 -5900 116620 -5880
rect 116880 -5900 117120 -5880
rect 117380 -5900 117620 -5880
rect 117880 -5900 118120 -5880
rect 118380 -5900 118620 -5880
rect 118880 -5900 119120 -5880
rect 119380 -5900 119620 -5880
rect 119880 -5900 120120 -5880
rect 120380 -5900 120620 -5880
rect 120880 -5900 121120 -5880
rect 121380 -5900 121620 -5880
rect 121880 -5900 122120 -5880
rect 122380 -5900 122620 -5880
rect 122880 -5900 123120 -5880
rect 123380 -5900 123620 -5880
rect 123880 -5900 124120 -5880
rect 124380 -5900 124620 -5880
rect 124880 -5900 125120 -5880
rect 125380 -5900 125620 -5880
rect 125880 -5900 126120 -5880
rect 126380 -5900 126620 -5880
rect 126880 -5900 127120 -5880
rect 127380 -5900 127620 -5880
rect 127880 -5900 128120 -5880
rect 128380 -5900 128620 -5880
rect 128880 -5900 129120 -5880
rect 129380 -5900 129620 -5880
rect 129880 -5900 130120 -5880
rect 130380 -5900 130620 -5880
rect 130880 -5900 131120 -5880
rect 131380 -5900 131620 -5880
rect 131880 -5900 132120 -5880
rect 132380 -5900 132620 -5880
rect 132880 -5900 133120 -5880
rect 133380 -5900 133620 -5880
rect 133880 -5900 134120 -5880
rect 134380 -5900 134620 -5880
rect 134880 -5900 135120 -5880
rect 135380 -5900 135620 -5880
rect 135880 -5900 136120 -5880
rect 136380 -5900 136620 -5880
rect 136880 -5900 137120 -5880
rect 137380 -5900 137620 -5880
rect 137880 -5900 138120 -5880
rect 138380 -5900 138620 -5880
rect 138880 -5900 139120 -5880
rect 139380 -5900 139620 -5880
rect 139880 -5900 140000 -5880
rect 88000 -6100 140000 -5900
rect 88000 -6120 88120 -6100
rect 88380 -6120 88620 -6100
rect 88880 -6120 89120 -6100
rect 89380 -6120 89620 -6100
rect 89880 -6120 90120 -6100
rect 90380 -6120 90620 -6100
rect 90880 -6120 91120 -6100
rect 91380 -6120 91620 -6100
rect 91880 -6120 92120 -6100
rect 92380 -6120 92620 -6100
rect 92880 -6120 93120 -6100
rect 93380 -6120 93620 -6100
rect 93880 -6120 94120 -6100
rect 94380 -6120 94620 -6100
rect 94880 -6120 95120 -6100
rect 95380 -6120 95620 -6100
rect 95880 -6120 96120 -6100
rect 96380 -6120 96620 -6100
rect 96880 -6120 97120 -6100
rect 97380 -6120 97620 -6100
rect 97880 -6120 98120 -6100
rect 98380 -6120 98620 -6100
rect 98880 -6120 99120 -6100
rect 99380 -6120 99620 -6100
rect 99880 -6120 100120 -6100
rect 100380 -6120 100620 -6100
rect 100880 -6120 101120 -6100
rect 101380 -6120 101620 -6100
rect 101880 -6120 102120 -6100
rect 102380 -6120 102620 -6100
rect 102880 -6120 103120 -6100
rect 103380 -6120 103620 -6100
rect 103880 -6120 104120 -6100
rect 104380 -6120 104620 -6100
rect 104880 -6120 105120 -6100
rect 105380 -6120 105620 -6100
rect 105880 -6120 106120 -6100
rect 106380 -6120 106620 -6100
rect 106880 -6120 107120 -6100
rect 107380 -6120 107620 -6100
rect 107880 -6120 108120 -6100
rect 108380 -6120 108620 -6100
rect 108880 -6120 109120 -6100
rect 109380 -6120 109620 -6100
rect 109880 -6120 110120 -6100
rect 110380 -6120 110620 -6100
rect 110880 -6120 111120 -6100
rect 111380 -6120 111620 -6100
rect 111880 -6120 112120 -6100
rect 112380 -6120 112620 -6100
rect 112880 -6120 113120 -6100
rect 113380 -6120 113620 -6100
rect 113880 -6120 114120 -6100
rect 114380 -6120 114620 -6100
rect 114880 -6120 115120 -6100
rect 115380 -6120 115620 -6100
rect 115880 -6120 116120 -6100
rect 116380 -6120 116620 -6100
rect 116880 -6120 117120 -6100
rect 117380 -6120 117620 -6100
rect 117880 -6120 118120 -6100
rect 118380 -6120 118620 -6100
rect 118880 -6120 119120 -6100
rect 119380 -6120 119620 -6100
rect 119880 -6120 120120 -6100
rect 120380 -6120 120620 -6100
rect 120880 -6120 121120 -6100
rect 121380 -6120 121620 -6100
rect 121880 -6120 122120 -6100
rect 122380 -6120 122620 -6100
rect 122880 -6120 123120 -6100
rect 123380 -6120 123620 -6100
rect 123880 -6120 124120 -6100
rect 124380 -6120 124620 -6100
rect 124880 -6120 125120 -6100
rect 125380 -6120 125620 -6100
rect 125880 -6120 126120 -6100
rect 126380 -6120 126620 -6100
rect 126880 -6120 127120 -6100
rect 127380 -6120 127620 -6100
rect 127880 -6120 128120 -6100
rect 128380 -6120 128620 -6100
rect 128880 -6120 129120 -6100
rect 129380 -6120 129620 -6100
rect 129880 -6120 130120 -6100
rect 130380 -6120 130620 -6100
rect 130880 -6120 131120 -6100
rect 131380 -6120 131620 -6100
rect 131880 -6120 132120 -6100
rect 132380 -6120 132620 -6100
rect 132880 -6120 133120 -6100
rect 133380 -6120 133620 -6100
rect 133880 -6120 134120 -6100
rect 134380 -6120 134620 -6100
rect 134880 -6120 135120 -6100
rect 135380 -6120 135620 -6100
rect 135880 -6120 136120 -6100
rect 136380 -6120 136620 -6100
rect 136880 -6120 137120 -6100
rect 137380 -6120 137620 -6100
rect 137880 -6120 138120 -6100
rect 138380 -6120 138620 -6100
rect 138880 -6120 139120 -6100
rect 139380 -6120 139620 -6100
rect 139880 -6120 140000 -6100
rect 88000 -6380 88100 -6120
rect 88400 -6380 88600 -6120
rect 88900 -6380 89100 -6120
rect 89400 -6380 89600 -6120
rect 89900 -6380 90100 -6120
rect 90400 -6380 90600 -6120
rect 90900 -6380 91100 -6120
rect 91400 -6380 91600 -6120
rect 91900 -6380 92100 -6120
rect 92400 -6380 92600 -6120
rect 92900 -6380 93100 -6120
rect 93400 -6380 93600 -6120
rect 93900 -6380 94100 -6120
rect 94400 -6380 94600 -6120
rect 94900 -6380 95100 -6120
rect 95400 -6380 95600 -6120
rect 95900 -6380 96100 -6120
rect 96400 -6380 96600 -6120
rect 96900 -6380 97100 -6120
rect 97400 -6380 97600 -6120
rect 97900 -6380 98100 -6120
rect 98400 -6380 98600 -6120
rect 98900 -6380 99100 -6120
rect 99400 -6380 99600 -6120
rect 99900 -6380 100100 -6120
rect 100400 -6380 100600 -6120
rect 100900 -6380 101100 -6120
rect 101400 -6380 101600 -6120
rect 101900 -6380 102100 -6120
rect 102400 -6380 102600 -6120
rect 102900 -6380 103100 -6120
rect 103400 -6380 103600 -6120
rect 103900 -6380 104100 -6120
rect 104400 -6380 104600 -6120
rect 104900 -6380 105100 -6120
rect 105400 -6380 105600 -6120
rect 105900 -6380 106100 -6120
rect 106400 -6380 106600 -6120
rect 106900 -6380 107100 -6120
rect 107400 -6380 107600 -6120
rect 107900 -6380 108100 -6120
rect 108400 -6380 108600 -6120
rect 108900 -6380 109100 -6120
rect 109400 -6380 109600 -6120
rect 109900 -6380 110100 -6120
rect 110400 -6380 110600 -6120
rect 110900 -6380 111100 -6120
rect 111400 -6380 111600 -6120
rect 111900 -6380 112100 -6120
rect 112400 -6380 112600 -6120
rect 112900 -6380 113100 -6120
rect 113400 -6380 113600 -6120
rect 113900 -6380 114100 -6120
rect 114400 -6380 114600 -6120
rect 114900 -6380 115100 -6120
rect 115400 -6380 115600 -6120
rect 115900 -6380 116100 -6120
rect 116400 -6380 116600 -6120
rect 116900 -6380 117100 -6120
rect 117400 -6380 117600 -6120
rect 117900 -6380 118100 -6120
rect 118400 -6380 118600 -6120
rect 118900 -6380 119100 -6120
rect 119400 -6380 119600 -6120
rect 119900 -6380 120100 -6120
rect 120400 -6380 120600 -6120
rect 120900 -6380 121100 -6120
rect 121400 -6380 121600 -6120
rect 121900 -6380 122100 -6120
rect 122400 -6380 122600 -6120
rect 122900 -6380 123100 -6120
rect 123400 -6380 123600 -6120
rect 123900 -6380 124100 -6120
rect 124400 -6380 124600 -6120
rect 124900 -6380 125100 -6120
rect 125400 -6380 125600 -6120
rect 125900 -6380 126100 -6120
rect 126400 -6380 126600 -6120
rect 126900 -6380 127100 -6120
rect 127400 -6380 127600 -6120
rect 127900 -6380 128100 -6120
rect 128400 -6380 128600 -6120
rect 128900 -6380 129100 -6120
rect 129400 -6380 129600 -6120
rect 129900 -6380 130100 -6120
rect 130400 -6380 130600 -6120
rect 130900 -6380 131100 -6120
rect 131400 -6380 131600 -6120
rect 131900 -6380 132100 -6120
rect 132400 -6380 132600 -6120
rect 132900 -6380 133100 -6120
rect 133400 -6380 133600 -6120
rect 133900 -6380 134100 -6120
rect 134400 -6380 134600 -6120
rect 134900 -6380 135100 -6120
rect 135400 -6380 135600 -6120
rect 135900 -6380 136100 -6120
rect 136400 -6380 136600 -6120
rect 136900 -6380 137100 -6120
rect 137400 -6380 137600 -6120
rect 137900 -6380 138100 -6120
rect 138400 -6380 138600 -6120
rect 138900 -6380 139100 -6120
rect 139400 -6380 139600 -6120
rect 139900 -6380 140000 -6120
rect 88000 -6400 88120 -6380
rect 88380 -6400 88620 -6380
rect 88880 -6400 89120 -6380
rect 89380 -6400 89620 -6380
rect 89880 -6400 90120 -6380
rect 90380 -6400 90620 -6380
rect 90880 -6400 91120 -6380
rect 91380 -6400 91620 -6380
rect 91880 -6400 92120 -6380
rect 92380 -6400 92620 -6380
rect 92880 -6400 93120 -6380
rect 93380 -6400 93620 -6380
rect 93880 -6400 94120 -6380
rect 94380 -6400 94620 -6380
rect 94880 -6400 95120 -6380
rect 95380 -6400 95620 -6380
rect 95880 -6400 96120 -6380
rect 96380 -6400 96620 -6380
rect 96880 -6400 97120 -6380
rect 97380 -6400 97620 -6380
rect 97880 -6400 98120 -6380
rect 98380 -6400 98620 -6380
rect 98880 -6400 99120 -6380
rect 99380 -6400 99620 -6380
rect 99880 -6400 100120 -6380
rect 100380 -6400 100620 -6380
rect 100880 -6400 101120 -6380
rect 101380 -6400 101620 -6380
rect 101880 -6400 102120 -6380
rect 102380 -6400 102620 -6380
rect 102880 -6400 103120 -6380
rect 103380 -6400 103620 -6380
rect 103880 -6400 104120 -6380
rect 104380 -6400 104620 -6380
rect 104880 -6400 105120 -6380
rect 105380 -6400 105620 -6380
rect 105880 -6400 106120 -6380
rect 106380 -6400 106620 -6380
rect 106880 -6400 107120 -6380
rect 107380 -6400 107620 -6380
rect 107880 -6400 108120 -6380
rect 108380 -6400 108620 -6380
rect 108880 -6400 109120 -6380
rect 109380 -6400 109620 -6380
rect 109880 -6400 110120 -6380
rect 110380 -6400 110620 -6380
rect 110880 -6400 111120 -6380
rect 111380 -6400 111620 -6380
rect 111880 -6400 112120 -6380
rect 112380 -6400 112620 -6380
rect 112880 -6400 113120 -6380
rect 113380 -6400 113620 -6380
rect 113880 -6400 114120 -6380
rect 114380 -6400 114620 -6380
rect 114880 -6400 115120 -6380
rect 115380 -6400 115620 -6380
rect 115880 -6400 116120 -6380
rect 116380 -6400 116620 -6380
rect 116880 -6400 117120 -6380
rect 117380 -6400 117620 -6380
rect 117880 -6400 118120 -6380
rect 118380 -6400 118620 -6380
rect 118880 -6400 119120 -6380
rect 119380 -6400 119620 -6380
rect 119880 -6400 120120 -6380
rect 120380 -6400 120620 -6380
rect 120880 -6400 121120 -6380
rect 121380 -6400 121620 -6380
rect 121880 -6400 122120 -6380
rect 122380 -6400 122620 -6380
rect 122880 -6400 123120 -6380
rect 123380 -6400 123620 -6380
rect 123880 -6400 124120 -6380
rect 124380 -6400 124620 -6380
rect 124880 -6400 125120 -6380
rect 125380 -6400 125620 -6380
rect 125880 -6400 126120 -6380
rect 126380 -6400 126620 -6380
rect 126880 -6400 127120 -6380
rect 127380 -6400 127620 -6380
rect 127880 -6400 128120 -6380
rect 128380 -6400 128620 -6380
rect 128880 -6400 129120 -6380
rect 129380 -6400 129620 -6380
rect 129880 -6400 130120 -6380
rect 130380 -6400 130620 -6380
rect 130880 -6400 131120 -6380
rect 131380 -6400 131620 -6380
rect 131880 -6400 132120 -6380
rect 132380 -6400 132620 -6380
rect 132880 -6400 133120 -6380
rect 133380 -6400 133620 -6380
rect 133880 -6400 134120 -6380
rect 134380 -6400 134620 -6380
rect 134880 -6400 135120 -6380
rect 135380 -6400 135620 -6380
rect 135880 -6400 136120 -6380
rect 136380 -6400 136620 -6380
rect 136880 -6400 137120 -6380
rect 137380 -6400 137620 -6380
rect 137880 -6400 138120 -6380
rect 138380 -6400 138620 -6380
rect 138880 -6400 139120 -6380
rect 139380 -6400 139620 -6380
rect 139880 -6400 140000 -6380
rect 88000 -6600 140000 -6400
rect 88000 -6620 88120 -6600
rect 88380 -6620 88620 -6600
rect 88880 -6620 89120 -6600
rect 89380 -6620 89620 -6600
rect 89880 -6620 90120 -6600
rect 90380 -6620 90620 -6600
rect 90880 -6620 91120 -6600
rect 91380 -6620 91620 -6600
rect 91880 -6620 92120 -6600
rect 92380 -6620 92620 -6600
rect 92880 -6620 93120 -6600
rect 93380 -6620 93620 -6600
rect 93880 -6620 94120 -6600
rect 94380 -6620 94620 -6600
rect 94880 -6620 95120 -6600
rect 95380 -6620 95620 -6600
rect 95880 -6620 96120 -6600
rect 96380 -6620 96620 -6600
rect 96880 -6620 97120 -6600
rect 97380 -6620 97620 -6600
rect 97880 -6620 98120 -6600
rect 98380 -6620 98620 -6600
rect 98880 -6620 99120 -6600
rect 99380 -6620 99620 -6600
rect 99880 -6620 100120 -6600
rect 100380 -6620 100620 -6600
rect 100880 -6620 101120 -6600
rect 101380 -6620 101620 -6600
rect 101880 -6620 102120 -6600
rect 102380 -6620 102620 -6600
rect 102880 -6620 103120 -6600
rect 103380 -6620 103620 -6600
rect 103880 -6620 104120 -6600
rect 104380 -6620 104620 -6600
rect 104880 -6620 105120 -6600
rect 105380 -6620 105620 -6600
rect 105880 -6620 106120 -6600
rect 106380 -6620 106620 -6600
rect 106880 -6620 107120 -6600
rect 107380 -6620 107620 -6600
rect 107880 -6620 108120 -6600
rect 108380 -6620 108620 -6600
rect 108880 -6620 109120 -6600
rect 109380 -6620 109620 -6600
rect 109880 -6620 110120 -6600
rect 110380 -6620 110620 -6600
rect 110880 -6620 111120 -6600
rect 111380 -6620 111620 -6600
rect 111880 -6620 112120 -6600
rect 112380 -6620 112620 -6600
rect 112880 -6620 113120 -6600
rect 113380 -6620 113620 -6600
rect 113880 -6620 114120 -6600
rect 114380 -6620 114620 -6600
rect 114880 -6620 115120 -6600
rect 115380 -6620 115620 -6600
rect 115880 -6620 116120 -6600
rect 116380 -6620 116620 -6600
rect 116880 -6620 117120 -6600
rect 117380 -6620 117620 -6600
rect 117880 -6620 118120 -6600
rect 118380 -6620 118620 -6600
rect 118880 -6620 119120 -6600
rect 119380 -6620 119620 -6600
rect 119880 -6620 120120 -6600
rect 120380 -6620 120620 -6600
rect 120880 -6620 121120 -6600
rect 121380 -6620 121620 -6600
rect 121880 -6620 122120 -6600
rect 122380 -6620 122620 -6600
rect 122880 -6620 123120 -6600
rect 123380 -6620 123620 -6600
rect 123880 -6620 124120 -6600
rect 124380 -6620 124620 -6600
rect 124880 -6620 125120 -6600
rect 125380 -6620 125620 -6600
rect 125880 -6620 126120 -6600
rect 126380 -6620 126620 -6600
rect 126880 -6620 127120 -6600
rect 127380 -6620 127620 -6600
rect 127880 -6620 128120 -6600
rect 128380 -6620 128620 -6600
rect 128880 -6620 129120 -6600
rect 129380 -6620 129620 -6600
rect 129880 -6620 130120 -6600
rect 130380 -6620 130620 -6600
rect 130880 -6620 131120 -6600
rect 131380 -6620 131620 -6600
rect 131880 -6620 132120 -6600
rect 132380 -6620 132620 -6600
rect 132880 -6620 133120 -6600
rect 133380 -6620 133620 -6600
rect 133880 -6620 134120 -6600
rect 134380 -6620 134620 -6600
rect 134880 -6620 135120 -6600
rect 135380 -6620 135620 -6600
rect 135880 -6620 136120 -6600
rect 136380 -6620 136620 -6600
rect 136880 -6620 137120 -6600
rect 137380 -6620 137620 -6600
rect 137880 -6620 138120 -6600
rect 138380 -6620 138620 -6600
rect 138880 -6620 139120 -6600
rect 139380 -6620 139620 -6600
rect 139880 -6620 140000 -6600
rect 88000 -6880 88100 -6620
rect 88400 -6880 88600 -6620
rect 88900 -6880 89100 -6620
rect 89400 -6880 89600 -6620
rect 89900 -6880 90100 -6620
rect 90400 -6880 90600 -6620
rect 90900 -6880 91100 -6620
rect 91400 -6880 91600 -6620
rect 91900 -6880 92100 -6620
rect 92400 -6880 92600 -6620
rect 92900 -6880 93100 -6620
rect 93400 -6880 93600 -6620
rect 93900 -6880 94100 -6620
rect 94400 -6880 94600 -6620
rect 94900 -6880 95100 -6620
rect 95400 -6880 95600 -6620
rect 95900 -6880 96100 -6620
rect 96400 -6880 96600 -6620
rect 96900 -6880 97100 -6620
rect 97400 -6880 97600 -6620
rect 97900 -6880 98100 -6620
rect 98400 -6880 98600 -6620
rect 98900 -6880 99100 -6620
rect 99400 -6880 99600 -6620
rect 99900 -6880 100100 -6620
rect 100400 -6880 100600 -6620
rect 100900 -6880 101100 -6620
rect 101400 -6880 101600 -6620
rect 101900 -6880 102100 -6620
rect 102400 -6880 102600 -6620
rect 102900 -6880 103100 -6620
rect 103400 -6880 103600 -6620
rect 103900 -6880 104100 -6620
rect 104400 -6880 104600 -6620
rect 104900 -6880 105100 -6620
rect 105400 -6880 105600 -6620
rect 105900 -6880 106100 -6620
rect 106400 -6880 106600 -6620
rect 106900 -6880 107100 -6620
rect 107400 -6880 107600 -6620
rect 107900 -6880 108100 -6620
rect 108400 -6880 108600 -6620
rect 108900 -6880 109100 -6620
rect 109400 -6880 109600 -6620
rect 109900 -6880 110100 -6620
rect 110400 -6880 110600 -6620
rect 110900 -6880 111100 -6620
rect 111400 -6880 111600 -6620
rect 111900 -6880 112100 -6620
rect 112400 -6880 112600 -6620
rect 112900 -6880 113100 -6620
rect 113400 -6880 113600 -6620
rect 113900 -6880 114100 -6620
rect 114400 -6880 114600 -6620
rect 114900 -6880 115100 -6620
rect 115400 -6880 115600 -6620
rect 115900 -6880 116100 -6620
rect 116400 -6880 116600 -6620
rect 116900 -6880 117100 -6620
rect 117400 -6880 117600 -6620
rect 117900 -6880 118100 -6620
rect 118400 -6880 118600 -6620
rect 118900 -6880 119100 -6620
rect 119400 -6880 119600 -6620
rect 119900 -6880 120100 -6620
rect 120400 -6880 120600 -6620
rect 120900 -6880 121100 -6620
rect 121400 -6880 121600 -6620
rect 121900 -6880 122100 -6620
rect 122400 -6880 122600 -6620
rect 122900 -6880 123100 -6620
rect 123400 -6880 123600 -6620
rect 123900 -6880 124100 -6620
rect 124400 -6880 124600 -6620
rect 124900 -6880 125100 -6620
rect 125400 -6880 125600 -6620
rect 125900 -6880 126100 -6620
rect 126400 -6880 126600 -6620
rect 126900 -6880 127100 -6620
rect 127400 -6880 127600 -6620
rect 127900 -6880 128100 -6620
rect 128400 -6880 128600 -6620
rect 128900 -6880 129100 -6620
rect 129400 -6880 129600 -6620
rect 129900 -6880 130100 -6620
rect 130400 -6880 130600 -6620
rect 130900 -6880 131100 -6620
rect 131400 -6880 131600 -6620
rect 131900 -6880 132100 -6620
rect 132400 -6880 132600 -6620
rect 132900 -6880 133100 -6620
rect 133400 -6880 133600 -6620
rect 133900 -6880 134100 -6620
rect 134400 -6880 134600 -6620
rect 134900 -6880 135100 -6620
rect 135400 -6880 135600 -6620
rect 135900 -6880 136100 -6620
rect 136400 -6880 136600 -6620
rect 136900 -6880 137100 -6620
rect 137400 -6880 137600 -6620
rect 137900 -6880 138100 -6620
rect 138400 -6880 138600 -6620
rect 138900 -6880 139100 -6620
rect 139400 -6880 139600 -6620
rect 139900 -6880 140000 -6620
rect 88000 -6900 88120 -6880
rect 88380 -6900 88620 -6880
rect 88880 -6900 89120 -6880
rect 89380 -6900 89620 -6880
rect 89880 -6900 90120 -6880
rect 90380 -6900 90620 -6880
rect 90880 -6900 91120 -6880
rect 91380 -6900 91620 -6880
rect 91880 -6900 92120 -6880
rect 92380 -6900 92620 -6880
rect 92880 -6900 93120 -6880
rect 93380 -6900 93620 -6880
rect 93880 -6900 94120 -6880
rect 94380 -6900 94620 -6880
rect 94880 -6900 95120 -6880
rect 95380 -6900 95620 -6880
rect 95880 -6900 96120 -6880
rect 96380 -6900 96620 -6880
rect 96880 -6900 97120 -6880
rect 97380 -6900 97620 -6880
rect 97880 -6900 98120 -6880
rect 98380 -6900 98620 -6880
rect 98880 -6900 99120 -6880
rect 99380 -6900 99620 -6880
rect 99880 -6900 100120 -6880
rect 100380 -6900 100620 -6880
rect 100880 -6900 101120 -6880
rect 101380 -6900 101620 -6880
rect 101880 -6900 102120 -6880
rect 102380 -6900 102620 -6880
rect 102880 -6900 103120 -6880
rect 103380 -6900 103620 -6880
rect 103880 -6900 104120 -6880
rect 104380 -6900 104620 -6880
rect 104880 -6900 105120 -6880
rect 105380 -6900 105620 -6880
rect 105880 -6900 106120 -6880
rect 106380 -6900 106620 -6880
rect 106880 -6900 107120 -6880
rect 107380 -6900 107620 -6880
rect 107880 -6900 108120 -6880
rect 108380 -6900 108620 -6880
rect 108880 -6900 109120 -6880
rect 109380 -6900 109620 -6880
rect 109880 -6900 110120 -6880
rect 110380 -6900 110620 -6880
rect 110880 -6900 111120 -6880
rect 111380 -6900 111620 -6880
rect 111880 -6900 112120 -6880
rect 112380 -6900 112620 -6880
rect 112880 -6900 113120 -6880
rect 113380 -6900 113620 -6880
rect 113880 -6900 114120 -6880
rect 114380 -6900 114620 -6880
rect 114880 -6900 115120 -6880
rect 115380 -6900 115620 -6880
rect 115880 -6900 116120 -6880
rect 116380 -6900 116620 -6880
rect 116880 -6900 117120 -6880
rect 117380 -6900 117620 -6880
rect 117880 -6900 118120 -6880
rect 118380 -6900 118620 -6880
rect 118880 -6900 119120 -6880
rect 119380 -6900 119620 -6880
rect 119880 -6900 120120 -6880
rect 120380 -6900 120620 -6880
rect 120880 -6900 121120 -6880
rect 121380 -6900 121620 -6880
rect 121880 -6900 122120 -6880
rect 122380 -6900 122620 -6880
rect 122880 -6900 123120 -6880
rect 123380 -6900 123620 -6880
rect 123880 -6900 124120 -6880
rect 124380 -6900 124620 -6880
rect 124880 -6900 125120 -6880
rect 125380 -6900 125620 -6880
rect 125880 -6900 126120 -6880
rect 126380 -6900 126620 -6880
rect 126880 -6900 127120 -6880
rect 127380 -6900 127620 -6880
rect 127880 -6900 128120 -6880
rect 128380 -6900 128620 -6880
rect 128880 -6900 129120 -6880
rect 129380 -6900 129620 -6880
rect 129880 -6900 130120 -6880
rect 130380 -6900 130620 -6880
rect 130880 -6900 131120 -6880
rect 131380 -6900 131620 -6880
rect 131880 -6900 132120 -6880
rect 132380 -6900 132620 -6880
rect 132880 -6900 133120 -6880
rect 133380 -6900 133620 -6880
rect 133880 -6900 134120 -6880
rect 134380 -6900 134620 -6880
rect 134880 -6900 135120 -6880
rect 135380 -6900 135620 -6880
rect 135880 -6900 136120 -6880
rect 136380 -6900 136620 -6880
rect 136880 -6900 137120 -6880
rect 137380 -6900 137620 -6880
rect 137880 -6900 138120 -6880
rect 138380 -6900 138620 -6880
rect 138880 -6900 139120 -6880
rect 139380 -6900 139620 -6880
rect 139880 -6900 140000 -6880
rect 88000 -7100 140000 -6900
rect 88000 -7120 88120 -7100
rect 88380 -7120 88620 -7100
rect 88880 -7120 89120 -7100
rect 89380 -7120 89620 -7100
rect 89880 -7120 90120 -7100
rect 90380 -7120 90620 -7100
rect 90880 -7120 91120 -7100
rect 91380 -7120 91620 -7100
rect 91880 -7120 92120 -7100
rect 92380 -7120 92620 -7100
rect 92880 -7120 93120 -7100
rect 93380 -7120 93620 -7100
rect 93880 -7120 94120 -7100
rect 94380 -7120 94620 -7100
rect 94880 -7120 95120 -7100
rect 95380 -7120 95620 -7100
rect 95880 -7120 96120 -7100
rect 96380 -7120 96620 -7100
rect 96880 -7120 97120 -7100
rect 97380 -7120 97620 -7100
rect 97880 -7120 98120 -7100
rect 98380 -7120 98620 -7100
rect 98880 -7120 99120 -7100
rect 99380 -7120 99620 -7100
rect 99880 -7120 100120 -7100
rect 100380 -7120 100620 -7100
rect 100880 -7120 101120 -7100
rect 101380 -7120 101620 -7100
rect 101880 -7120 102120 -7100
rect 102380 -7120 102620 -7100
rect 102880 -7120 103120 -7100
rect 103380 -7120 103620 -7100
rect 103880 -7120 104120 -7100
rect 104380 -7120 104620 -7100
rect 104880 -7120 105120 -7100
rect 105380 -7120 105620 -7100
rect 105880 -7120 106120 -7100
rect 106380 -7120 106620 -7100
rect 106880 -7120 107120 -7100
rect 107380 -7120 107620 -7100
rect 107880 -7120 108120 -7100
rect 108380 -7120 108620 -7100
rect 108880 -7120 109120 -7100
rect 109380 -7120 109620 -7100
rect 109880 -7120 110120 -7100
rect 110380 -7120 110620 -7100
rect 110880 -7120 111120 -7100
rect 111380 -7120 111620 -7100
rect 111880 -7120 112120 -7100
rect 112380 -7120 112620 -7100
rect 112880 -7120 113120 -7100
rect 113380 -7120 113620 -7100
rect 113880 -7120 114120 -7100
rect 114380 -7120 114620 -7100
rect 114880 -7120 115120 -7100
rect 115380 -7120 115620 -7100
rect 115880 -7120 116120 -7100
rect 116380 -7120 116620 -7100
rect 116880 -7120 117120 -7100
rect 117380 -7120 117620 -7100
rect 117880 -7120 118120 -7100
rect 118380 -7120 118620 -7100
rect 118880 -7120 119120 -7100
rect 119380 -7120 119620 -7100
rect 119880 -7120 120120 -7100
rect 120380 -7120 120620 -7100
rect 120880 -7120 121120 -7100
rect 121380 -7120 121620 -7100
rect 121880 -7120 122120 -7100
rect 122380 -7120 122620 -7100
rect 122880 -7120 123120 -7100
rect 123380 -7120 123620 -7100
rect 123880 -7120 124120 -7100
rect 124380 -7120 124620 -7100
rect 124880 -7120 125120 -7100
rect 125380 -7120 125620 -7100
rect 125880 -7120 126120 -7100
rect 126380 -7120 126620 -7100
rect 126880 -7120 127120 -7100
rect 127380 -7120 127620 -7100
rect 127880 -7120 128120 -7100
rect 128380 -7120 128620 -7100
rect 128880 -7120 129120 -7100
rect 129380 -7120 129620 -7100
rect 129880 -7120 130120 -7100
rect 130380 -7120 130620 -7100
rect 130880 -7120 131120 -7100
rect 131380 -7120 131620 -7100
rect 131880 -7120 132120 -7100
rect 132380 -7120 132620 -7100
rect 132880 -7120 133120 -7100
rect 133380 -7120 133620 -7100
rect 133880 -7120 134120 -7100
rect 134380 -7120 134620 -7100
rect 134880 -7120 135120 -7100
rect 135380 -7120 135620 -7100
rect 135880 -7120 136120 -7100
rect 136380 -7120 136620 -7100
rect 136880 -7120 137120 -7100
rect 137380 -7120 137620 -7100
rect 137880 -7120 138120 -7100
rect 138380 -7120 138620 -7100
rect 138880 -7120 139120 -7100
rect 139380 -7120 139620 -7100
rect 139880 -7120 140000 -7100
rect 88000 -7380 88100 -7120
rect 88400 -7380 88600 -7120
rect 88900 -7380 89100 -7120
rect 89400 -7380 89600 -7120
rect 89900 -7380 90100 -7120
rect 90400 -7380 90600 -7120
rect 90900 -7380 91100 -7120
rect 91400 -7380 91600 -7120
rect 91900 -7380 92100 -7120
rect 92400 -7380 92600 -7120
rect 92900 -7380 93100 -7120
rect 93400 -7380 93600 -7120
rect 93900 -7380 94100 -7120
rect 94400 -7380 94600 -7120
rect 94900 -7380 95100 -7120
rect 95400 -7380 95600 -7120
rect 95900 -7380 96100 -7120
rect 96400 -7380 96600 -7120
rect 96900 -7380 97100 -7120
rect 97400 -7380 97600 -7120
rect 97900 -7380 98100 -7120
rect 98400 -7380 98600 -7120
rect 98900 -7380 99100 -7120
rect 99400 -7380 99600 -7120
rect 99900 -7380 100100 -7120
rect 100400 -7380 100600 -7120
rect 100900 -7380 101100 -7120
rect 101400 -7380 101600 -7120
rect 101900 -7380 102100 -7120
rect 102400 -7380 102600 -7120
rect 102900 -7380 103100 -7120
rect 103400 -7380 103600 -7120
rect 103900 -7380 104100 -7120
rect 104400 -7380 104600 -7120
rect 104900 -7380 105100 -7120
rect 105400 -7380 105600 -7120
rect 105900 -7380 106100 -7120
rect 106400 -7380 106600 -7120
rect 106900 -7380 107100 -7120
rect 107400 -7380 107600 -7120
rect 107900 -7380 108100 -7120
rect 108400 -7380 108600 -7120
rect 108900 -7380 109100 -7120
rect 109400 -7380 109600 -7120
rect 109900 -7380 110100 -7120
rect 110400 -7380 110600 -7120
rect 110900 -7380 111100 -7120
rect 111400 -7380 111600 -7120
rect 111900 -7380 112100 -7120
rect 112400 -7380 112600 -7120
rect 112900 -7380 113100 -7120
rect 113400 -7380 113600 -7120
rect 113900 -7380 114100 -7120
rect 114400 -7380 114600 -7120
rect 114900 -7380 115100 -7120
rect 115400 -7380 115600 -7120
rect 115900 -7380 116100 -7120
rect 116400 -7380 116600 -7120
rect 116900 -7380 117100 -7120
rect 117400 -7380 117600 -7120
rect 117900 -7380 118100 -7120
rect 118400 -7380 118600 -7120
rect 118900 -7380 119100 -7120
rect 119400 -7380 119600 -7120
rect 119900 -7380 120100 -7120
rect 120400 -7380 120600 -7120
rect 120900 -7380 121100 -7120
rect 121400 -7380 121600 -7120
rect 121900 -7380 122100 -7120
rect 122400 -7380 122600 -7120
rect 122900 -7380 123100 -7120
rect 123400 -7380 123600 -7120
rect 123900 -7380 124100 -7120
rect 124400 -7380 124600 -7120
rect 124900 -7380 125100 -7120
rect 125400 -7380 125600 -7120
rect 125900 -7380 126100 -7120
rect 126400 -7380 126600 -7120
rect 126900 -7380 127100 -7120
rect 127400 -7380 127600 -7120
rect 127900 -7380 128100 -7120
rect 128400 -7380 128600 -7120
rect 128900 -7380 129100 -7120
rect 129400 -7380 129600 -7120
rect 129900 -7380 130100 -7120
rect 130400 -7380 130600 -7120
rect 130900 -7380 131100 -7120
rect 131400 -7380 131600 -7120
rect 131900 -7380 132100 -7120
rect 132400 -7380 132600 -7120
rect 132900 -7380 133100 -7120
rect 133400 -7380 133600 -7120
rect 133900 -7380 134100 -7120
rect 134400 -7380 134600 -7120
rect 134900 -7380 135100 -7120
rect 135400 -7380 135600 -7120
rect 135900 -7380 136100 -7120
rect 136400 -7380 136600 -7120
rect 136900 -7380 137100 -7120
rect 137400 -7380 137600 -7120
rect 137900 -7380 138100 -7120
rect 138400 -7380 138600 -7120
rect 138900 -7380 139100 -7120
rect 139400 -7380 139600 -7120
rect 139900 -7380 140000 -7120
rect 88000 -7400 88120 -7380
rect 88380 -7400 88620 -7380
rect 88880 -7400 89120 -7380
rect 89380 -7400 89620 -7380
rect 89880 -7400 90120 -7380
rect 90380 -7400 90620 -7380
rect 90880 -7400 91120 -7380
rect 91380 -7400 91620 -7380
rect 91880 -7400 92120 -7380
rect 92380 -7400 92620 -7380
rect 92880 -7400 93120 -7380
rect 93380 -7400 93620 -7380
rect 93880 -7400 94120 -7380
rect 94380 -7400 94620 -7380
rect 94880 -7400 95120 -7380
rect 95380 -7400 95620 -7380
rect 95880 -7400 96120 -7380
rect 96380 -7400 96620 -7380
rect 96880 -7400 97120 -7380
rect 97380 -7400 97620 -7380
rect 97880 -7400 98120 -7380
rect 98380 -7400 98620 -7380
rect 98880 -7400 99120 -7380
rect 99380 -7400 99620 -7380
rect 99880 -7400 100120 -7380
rect 100380 -7400 100620 -7380
rect 100880 -7400 101120 -7380
rect 101380 -7400 101620 -7380
rect 101880 -7400 102120 -7380
rect 102380 -7400 102620 -7380
rect 102880 -7400 103120 -7380
rect 103380 -7400 103620 -7380
rect 103880 -7400 104120 -7380
rect 104380 -7400 104620 -7380
rect 104880 -7400 105120 -7380
rect 105380 -7400 105620 -7380
rect 105880 -7400 106120 -7380
rect 106380 -7400 106620 -7380
rect 106880 -7400 107120 -7380
rect 107380 -7400 107620 -7380
rect 107880 -7400 108120 -7380
rect 108380 -7400 108620 -7380
rect 108880 -7400 109120 -7380
rect 109380 -7400 109620 -7380
rect 109880 -7400 110120 -7380
rect 110380 -7400 110620 -7380
rect 110880 -7400 111120 -7380
rect 111380 -7400 111620 -7380
rect 111880 -7400 112120 -7380
rect 112380 -7400 112620 -7380
rect 112880 -7400 113120 -7380
rect 113380 -7400 113620 -7380
rect 113880 -7400 114120 -7380
rect 114380 -7400 114620 -7380
rect 114880 -7400 115120 -7380
rect 115380 -7400 115620 -7380
rect 115880 -7400 116120 -7380
rect 116380 -7400 116620 -7380
rect 116880 -7400 117120 -7380
rect 117380 -7400 117620 -7380
rect 117880 -7400 118120 -7380
rect 118380 -7400 118620 -7380
rect 118880 -7400 119120 -7380
rect 119380 -7400 119620 -7380
rect 119880 -7400 120120 -7380
rect 120380 -7400 120620 -7380
rect 120880 -7400 121120 -7380
rect 121380 -7400 121620 -7380
rect 121880 -7400 122120 -7380
rect 122380 -7400 122620 -7380
rect 122880 -7400 123120 -7380
rect 123380 -7400 123620 -7380
rect 123880 -7400 124120 -7380
rect 124380 -7400 124620 -7380
rect 124880 -7400 125120 -7380
rect 125380 -7400 125620 -7380
rect 125880 -7400 126120 -7380
rect 126380 -7400 126620 -7380
rect 126880 -7400 127120 -7380
rect 127380 -7400 127620 -7380
rect 127880 -7400 128120 -7380
rect 128380 -7400 128620 -7380
rect 128880 -7400 129120 -7380
rect 129380 -7400 129620 -7380
rect 129880 -7400 130120 -7380
rect 130380 -7400 130620 -7380
rect 130880 -7400 131120 -7380
rect 131380 -7400 131620 -7380
rect 131880 -7400 132120 -7380
rect 132380 -7400 132620 -7380
rect 132880 -7400 133120 -7380
rect 133380 -7400 133620 -7380
rect 133880 -7400 134120 -7380
rect 134380 -7400 134620 -7380
rect 134880 -7400 135120 -7380
rect 135380 -7400 135620 -7380
rect 135880 -7400 136120 -7380
rect 136380 -7400 136620 -7380
rect 136880 -7400 137120 -7380
rect 137380 -7400 137620 -7380
rect 137880 -7400 138120 -7380
rect 138380 -7400 138620 -7380
rect 138880 -7400 139120 -7380
rect 139380 -7400 139620 -7380
rect 139880 -7400 140000 -7380
rect 88000 -7600 140000 -7400
rect 88000 -7620 88120 -7600
rect 88380 -7620 88620 -7600
rect 88880 -7620 89120 -7600
rect 89380 -7620 89620 -7600
rect 89880 -7620 90120 -7600
rect 90380 -7620 90620 -7600
rect 90880 -7620 91120 -7600
rect 91380 -7620 91620 -7600
rect 91880 -7620 92120 -7600
rect 92380 -7620 92620 -7600
rect 92880 -7620 93120 -7600
rect 93380 -7620 93620 -7600
rect 93880 -7620 94120 -7600
rect 94380 -7620 94620 -7600
rect 94880 -7620 95120 -7600
rect 95380 -7620 95620 -7600
rect 95880 -7620 96120 -7600
rect 96380 -7620 96620 -7600
rect 96880 -7620 97120 -7600
rect 97380 -7620 97620 -7600
rect 97880 -7620 98120 -7600
rect 98380 -7620 98620 -7600
rect 98880 -7620 99120 -7600
rect 99380 -7620 99620 -7600
rect 99880 -7620 100120 -7600
rect 100380 -7620 100620 -7600
rect 100880 -7620 101120 -7600
rect 101380 -7620 101620 -7600
rect 101880 -7620 102120 -7600
rect 102380 -7620 102620 -7600
rect 102880 -7620 103120 -7600
rect 103380 -7620 103620 -7600
rect 103880 -7620 104120 -7600
rect 104380 -7620 104620 -7600
rect 104880 -7620 105120 -7600
rect 105380 -7620 105620 -7600
rect 105880 -7620 106120 -7600
rect 106380 -7620 106620 -7600
rect 106880 -7620 107120 -7600
rect 107380 -7620 107620 -7600
rect 107880 -7620 108120 -7600
rect 108380 -7620 108620 -7600
rect 108880 -7620 109120 -7600
rect 109380 -7620 109620 -7600
rect 109880 -7620 110120 -7600
rect 110380 -7620 110620 -7600
rect 110880 -7620 111120 -7600
rect 111380 -7620 111620 -7600
rect 111880 -7620 112120 -7600
rect 112380 -7620 112620 -7600
rect 112880 -7620 113120 -7600
rect 113380 -7620 113620 -7600
rect 113880 -7620 114120 -7600
rect 114380 -7620 114620 -7600
rect 114880 -7620 115120 -7600
rect 115380 -7620 115620 -7600
rect 115880 -7620 116120 -7600
rect 116380 -7620 116620 -7600
rect 116880 -7620 117120 -7600
rect 117380 -7620 117620 -7600
rect 117880 -7620 118120 -7600
rect 118380 -7620 118620 -7600
rect 118880 -7620 119120 -7600
rect 119380 -7620 119620 -7600
rect 119880 -7620 120120 -7600
rect 120380 -7620 120620 -7600
rect 120880 -7620 121120 -7600
rect 121380 -7620 121620 -7600
rect 121880 -7620 122120 -7600
rect 122380 -7620 122620 -7600
rect 122880 -7620 123120 -7600
rect 123380 -7620 123620 -7600
rect 123880 -7620 124120 -7600
rect 124380 -7620 124620 -7600
rect 124880 -7620 125120 -7600
rect 125380 -7620 125620 -7600
rect 125880 -7620 126120 -7600
rect 126380 -7620 126620 -7600
rect 126880 -7620 127120 -7600
rect 127380 -7620 127620 -7600
rect 127880 -7620 128120 -7600
rect 128380 -7620 128620 -7600
rect 128880 -7620 129120 -7600
rect 129380 -7620 129620 -7600
rect 129880 -7620 130120 -7600
rect 130380 -7620 130620 -7600
rect 130880 -7620 131120 -7600
rect 131380 -7620 131620 -7600
rect 131880 -7620 132120 -7600
rect 132380 -7620 132620 -7600
rect 132880 -7620 133120 -7600
rect 133380 -7620 133620 -7600
rect 133880 -7620 134120 -7600
rect 134380 -7620 134620 -7600
rect 134880 -7620 135120 -7600
rect 135380 -7620 135620 -7600
rect 135880 -7620 136120 -7600
rect 136380 -7620 136620 -7600
rect 136880 -7620 137120 -7600
rect 137380 -7620 137620 -7600
rect 137880 -7620 138120 -7600
rect 138380 -7620 138620 -7600
rect 138880 -7620 139120 -7600
rect 139380 -7620 139620 -7600
rect 139880 -7620 140000 -7600
rect 88000 -7880 88100 -7620
rect 88400 -7880 88600 -7620
rect 88900 -7880 89100 -7620
rect 89400 -7880 89600 -7620
rect 89900 -7880 90100 -7620
rect 90400 -7880 90600 -7620
rect 90900 -7880 91100 -7620
rect 91400 -7880 91600 -7620
rect 91900 -7880 92100 -7620
rect 92400 -7880 92600 -7620
rect 92900 -7880 93100 -7620
rect 93400 -7880 93600 -7620
rect 93900 -7880 94100 -7620
rect 94400 -7880 94600 -7620
rect 94900 -7880 95100 -7620
rect 95400 -7880 95600 -7620
rect 95900 -7880 96100 -7620
rect 96400 -7880 96600 -7620
rect 96900 -7880 97100 -7620
rect 97400 -7880 97600 -7620
rect 97900 -7880 98100 -7620
rect 98400 -7880 98600 -7620
rect 98900 -7880 99100 -7620
rect 99400 -7880 99600 -7620
rect 99900 -7880 100100 -7620
rect 100400 -7880 100600 -7620
rect 100900 -7880 101100 -7620
rect 101400 -7880 101600 -7620
rect 101900 -7880 102100 -7620
rect 102400 -7880 102600 -7620
rect 102900 -7880 103100 -7620
rect 103400 -7880 103600 -7620
rect 103900 -7880 104100 -7620
rect 104400 -7880 104600 -7620
rect 104900 -7880 105100 -7620
rect 105400 -7880 105600 -7620
rect 105900 -7880 106100 -7620
rect 106400 -7880 106600 -7620
rect 106900 -7880 107100 -7620
rect 107400 -7880 107600 -7620
rect 107900 -7880 108100 -7620
rect 108400 -7880 108600 -7620
rect 108900 -7880 109100 -7620
rect 109400 -7880 109600 -7620
rect 109900 -7880 110100 -7620
rect 110400 -7880 110600 -7620
rect 110900 -7880 111100 -7620
rect 111400 -7880 111600 -7620
rect 111900 -7880 112100 -7620
rect 112400 -7880 112600 -7620
rect 112900 -7880 113100 -7620
rect 113400 -7880 113600 -7620
rect 113900 -7880 114100 -7620
rect 114400 -7880 114600 -7620
rect 114900 -7880 115100 -7620
rect 115400 -7880 115600 -7620
rect 115900 -7880 116100 -7620
rect 116400 -7880 116600 -7620
rect 116900 -7880 117100 -7620
rect 117400 -7880 117600 -7620
rect 117900 -7880 118100 -7620
rect 118400 -7880 118600 -7620
rect 118900 -7880 119100 -7620
rect 119400 -7880 119600 -7620
rect 119900 -7880 120100 -7620
rect 120400 -7880 120600 -7620
rect 120900 -7880 121100 -7620
rect 121400 -7880 121600 -7620
rect 121900 -7880 122100 -7620
rect 122400 -7880 122600 -7620
rect 122900 -7880 123100 -7620
rect 123400 -7880 123600 -7620
rect 123900 -7880 124100 -7620
rect 124400 -7880 124600 -7620
rect 124900 -7880 125100 -7620
rect 125400 -7880 125600 -7620
rect 125900 -7880 126100 -7620
rect 126400 -7880 126600 -7620
rect 126900 -7880 127100 -7620
rect 127400 -7880 127600 -7620
rect 127900 -7880 128100 -7620
rect 128400 -7880 128600 -7620
rect 128900 -7880 129100 -7620
rect 129400 -7880 129600 -7620
rect 129900 -7880 130100 -7620
rect 130400 -7880 130600 -7620
rect 130900 -7880 131100 -7620
rect 131400 -7880 131600 -7620
rect 131900 -7880 132100 -7620
rect 132400 -7880 132600 -7620
rect 132900 -7880 133100 -7620
rect 133400 -7880 133600 -7620
rect 133900 -7880 134100 -7620
rect 134400 -7880 134600 -7620
rect 134900 -7880 135100 -7620
rect 135400 -7880 135600 -7620
rect 135900 -7880 136100 -7620
rect 136400 -7880 136600 -7620
rect 136900 -7880 137100 -7620
rect 137400 -7880 137600 -7620
rect 137900 -7880 138100 -7620
rect 138400 -7880 138600 -7620
rect 138900 -7880 139100 -7620
rect 139400 -7880 139600 -7620
rect 139900 -7880 140000 -7620
rect 88000 -7900 88120 -7880
rect 88380 -7900 88620 -7880
rect 88880 -7900 89120 -7880
rect 89380 -7900 89620 -7880
rect 89880 -7900 90120 -7880
rect 90380 -7900 90620 -7880
rect 90880 -7900 91120 -7880
rect 91380 -7900 91620 -7880
rect 91880 -7900 92120 -7880
rect 92380 -7900 92620 -7880
rect 92880 -7900 93120 -7880
rect 93380 -7900 93620 -7880
rect 93880 -7900 94120 -7880
rect 94380 -7900 94620 -7880
rect 94880 -7900 95120 -7880
rect 95380 -7900 95620 -7880
rect 95880 -7900 96120 -7880
rect 96380 -7900 96620 -7880
rect 96880 -7900 97120 -7880
rect 97380 -7900 97620 -7880
rect 97880 -7900 98120 -7880
rect 98380 -7900 98620 -7880
rect 98880 -7900 99120 -7880
rect 99380 -7900 99620 -7880
rect 99880 -7900 100120 -7880
rect 100380 -7900 100620 -7880
rect 100880 -7900 101120 -7880
rect 101380 -7900 101620 -7880
rect 101880 -7900 102120 -7880
rect 102380 -7900 102620 -7880
rect 102880 -7900 103120 -7880
rect 103380 -7900 103620 -7880
rect 103880 -7900 104120 -7880
rect 104380 -7900 104620 -7880
rect 104880 -7900 105120 -7880
rect 105380 -7900 105620 -7880
rect 105880 -7900 106120 -7880
rect 106380 -7900 106620 -7880
rect 106880 -7900 107120 -7880
rect 107380 -7900 107620 -7880
rect 107880 -7900 108120 -7880
rect 108380 -7900 108620 -7880
rect 108880 -7900 109120 -7880
rect 109380 -7900 109620 -7880
rect 109880 -7900 110120 -7880
rect 110380 -7900 110620 -7880
rect 110880 -7900 111120 -7880
rect 111380 -7900 111620 -7880
rect 111880 -7900 112120 -7880
rect 112380 -7900 112620 -7880
rect 112880 -7900 113120 -7880
rect 113380 -7900 113620 -7880
rect 113880 -7900 114120 -7880
rect 114380 -7900 114620 -7880
rect 114880 -7900 115120 -7880
rect 115380 -7900 115620 -7880
rect 115880 -7900 116120 -7880
rect 116380 -7900 116620 -7880
rect 116880 -7900 117120 -7880
rect 117380 -7900 117620 -7880
rect 117880 -7900 118120 -7880
rect 118380 -7900 118620 -7880
rect 118880 -7900 119120 -7880
rect 119380 -7900 119620 -7880
rect 119880 -7900 120120 -7880
rect 120380 -7900 120620 -7880
rect 120880 -7900 121120 -7880
rect 121380 -7900 121620 -7880
rect 121880 -7900 122120 -7880
rect 122380 -7900 122620 -7880
rect 122880 -7900 123120 -7880
rect 123380 -7900 123620 -7880
rect 123880 -7900 124120 -7880
rect 124380 -7900 124620 -7880
rect 124880 -7900 125120 -7880
rect 125380 -7900 125620 -7880
rect 125880 -7900 126120 -7880
rect 126380 -7900 126620 -7880
rect 126880 -7900 127120 -7880
rect 127380 -7900 127620 -7880
rect 127880 -7900 128120 -7880
rect 128380 -7900 128620 -7880
rect 128880 -7900 129120 -7880
rect 129380 -7900 129620 -7880
rect 129880 -7900 130120 -7880
rect 130380 -7900 130620 -7880
rect 130880 -7900 131120 -7880
rect 131380 -7900 131620 -7880
rect 131880 -7900 132120 -7880
rect 132380 -7900 132620 -7880
rect 132880 -7900 133120 -7880
rect 133380 -7900 133620 -7880
rect 133880 -7900 134120 -7880
rect 134380 -7900 134620 -7880
rect 134880 -7900 135120 -7880
rect 135380 -7900 135620 -7880
rect 135880 -7900 136120 -7880
rect 136380 -7900 136620 -7880
rect 136880 -7900 137120 -7880
rect 137380 -7900 137620 -7880
rect 137880 -7900 138120 -7880
rect 138380 -7900 138620 -7880
rect 138880 -7900 139120 -7880
rect 139380 -7900 139620 -7880
rect 139880 -7900 140000 -7880
rect 88000 -8100 140000 -7900
rect 88000 -8120 88120 -8100
rect 88380 -8120 88620 -8100
rect 88880 -8120 89120 -8100
rect 89380 -8120 89620 -8100
rect 89880 -8120 90120 -8100
rect 90380 -8120 90620 -8100
rect 90880 -8120 91120 -8100
rect 91380 -8120 91620 -8100
rect 91880 -8120 92120 -8100
rect 92380 -8120 92620 -8100
rect 92880 -8120 93120 -8100
rect 93380 -8120 93620 -8100
rect 93880 -8120 94120 -8100
rect 94380 -8120 94620 -8100
rect 94880 -8120 95120 -8100
rect 95380 -8120 95620 -8100
rect 95880 -8120 96120 -8100
rect 96380 -8120 96620 -8100
rect 96880 -8120 97120 -8100
rect 97380 -8120 97620 -8100
rect 97880 -8120 98120 -8100
rect 98380 -8120 98620 -8100
rect 98880 -8120 99120 -8100
rect 99380 -8120 99620 -8100
rect 99880 -8120 100120 -8100
rect 100380 -8120 100620 -8100
rect 100880 -8120 101120 -8100
rect 101380 -8120 101620 -8100
rect 101880 -8120 102120 -8100
rect 102380 -8120 102620 -8100
rect 102880 -8120 103120 -8100
rect 103380 -8120 103620 -8100
rect 103880 -8120 104120 -8100
rect 104380 -8120 104620 -8100
rect 104880 -8120 105120 -8100
rect 105380 -8120 105620 -8100
rect 105880 -8120 106120 -8100
rect 106380 -8120 106620 -8100
rect 106880 -8120 107120 -8100
rect 107380 -8120 107620 -8100
rect 107880 -8120 108120 -8100
rect 108380 -8120 108620 -8100
rect 108880 -8120 109120 -8100
rect 109380 -8120 109620 -8100
rect 109880 -8120 110120 -8100
rect 110380 -8120 110620 -8100
rect 110880 -8120 111120 -8100
rect 111380 -8120 111620 -8100
rect 111880 -8120 112120 -8100
rect 112380 -8120 112620 -8100
rect 112880 -8120 113120 -8100
rect 113380 -8120 113620 -8100
rect 113880 -8120 114120 -8100
rect 114380 -8120 114620 -8100
rect 114880 -8120 115120 -8100
rect 115380 -8120 115620 -8100
rect 115880 -8120 116120 -8100
rect 116380 -8120 116620 -8100
rect 116880 -8120 117120 -8100
rect 117380 -8120 117620 -8100
rect 117880 -8120 118120 -8100
rect 118380 -8120 118620 -8100
rect 118880 -8120 119120 -8100
rect 119380 -8120 119620 -8100
rect 119880 -8120 120120 -8100
rect 120380 -8120 120620 -8100
rect 120880 -8120 121120 -8100
rect 121380 -8120 121620 -8100
rect 121880 -8120 122120 -8100
rect 122380 -8120 122620 -8100
rect 122880 -8120 123120 -8100
rect 123380 -8120 123620 -8100
rect 123880 -8120 124120 -8100
rect 124380 -8120 124620 -8100
rect 124880 -8120 125120 -8100
rect 125380 -8120 125620 -8100
rect 125880 -8120 126120 -8100
rect 126380 -8120 126620 -8100
rect 126880 -8120 127120 -8100
rect 127380 -8120 127620 -8100
rect 127880 -8120 128120 -8100
rect 128380 -8120 128620 -8100
rect 128880 -8120 129120 -8100
rect 129380 -8120 129620 -8100
rect 129880 -8120 130120 -8100
rect 130380 -8120 130620 -8100
rect 130880 -8120 131120 -8100
rect 131380 -8120 131620 -8100
rect 131880 -8120 132120 -8100
rect 132380 -8120 132620 -8100
rect 132880 -8120 133120 -8100
rect 133380 -8120 133620 -8100
rect 133880 -8120 134120 -8100
rect 134380 -8120 134620 -8100
rect 134880 -8120 135120 -8100
rect 135380 -8120 135620 -8100
rect 135880 -8120 136120 -8100
rect 136380 -8120 136620 -8100
rect 136880 -8120 137120 -8100
rect 137380 -8120 137620 -8100
rect 137880 -8120 138120 -8100
rect 138380 -8120 138620 -8100
rect 138880 -8120 139120 -8100
rect 139380 -8120 139620 -8100
rect 139880 -8120 140000 -8100
rect 88000 -8380 88100 -8120
rect 88400 -8380 88600 -8120
rect 88900 -8380 89100 -8120
rect 89400 -8380 89600 -8120
rect 89900 -8380 90100 -8120
rect 90400 -8380 90600 -8120
rect 90900 -8380 91100 -8120
rect 91400 -8380 91600 -8120
rect 91900 -8380 92100 -8120
rect 92400 -8380 92600 -8120
rect 92900 -8380 93100 -8120
rect 93400 -8380 93600 -8120
rect 93900 -8380 94100 -8120
rect 94400 -8380 94600 -8120
rect 94900 -8380 95100 -8120
rect 95400 -8380 95600 -8120
rect 95900 -8380 96100 -8120
rect 96400 -8380 96600 -8120
rect 96900 -8380 97100 -8120
rect 97400 -8380 97600 -8120
rect 97900 -8380 98100 -8120
rect 98400 -8380 98600 -8120
rect 98900 -8380 99100 -8120
rect 99400 -8380 99600 -8120
rect 99900 -8380 100100 -8120
rect 100400 -8380 100600 -8120
rect 100900 -8380 101100 -8120
rect 101400 -8380 101600 -8120
rect 101900 -8380 102100 -8120
rect 102400 -8380 102600 -8120
rect 102900 -8380 103100 -8120
rect 103400 -8380 103600 -8120
rect 103900 -8380 104100 -8120
rect 104400 -8380 104600 -8120
rect 104900 -8380 105100 -8120
rect 105400 -8380 105600 -8120
rect 105900 -8380 106100 -8120
rect 106400 -8380 106600 -8120
rect 106900 -8380 107100 -8120
rect 107400 -8380 107600 -8120
rect 107900 -8380 108100 -8120
rect 108400 -8380 108600 -8120
rect 108900 -8380 109100 -8120
rect 109400 -8380 109600 -8120
rect 109900 -8380 110100 -8120
rect 110400 -8380 110600 -8120
rect 110900 -8380 111100 -8120
rect 111400 -8380 111600 -8120
rect 111900 -8380 112100 -8120
rect 112400 -8380 112600 -8120
rect 112900 -8380 113100 -8120
rect 113400 -8380 113600 -8120
rect 113900 -8380 114100 -8120
rect 114400 -8380 114600 -8120
rect 114900 -8380 115100 -8120
rect 115400 -8380 115600 -8120
rect 115900 -8380 116100 -8120
rect 116400 -8380 116600 -8120
rect 116900 -8380 117100 -8120
rect 117400 -8380 117600 -8120
rect 117900 -8380 118100 -8120
rect 118400 -8380 118600 -8120
rect 118900 -8380 119100 -8120
rect 119400 -8380 119600 -8120
rect 119900 -8380 120100 -8120
rect 120400 -8380 120600 -8120
rect 120900 -8380 121100 -8120
rect 121400 -8380 121600 -8120
rect 121900 -8380 122100 -8120
rect 122400 -8380 122600 -8120
rect 122900 -8380 123100 -8120
rect 123400 -8380 123600 -8120
rect 123900 -8380 124100 -8120
rect 124400 -8380 124600 -8120
rect 124900 -8380 125100 -8120
rect 125400 -8380 125600 -8120
rect 125900 -8380 126100 -8120
rect 126400 -8380 126600 -8120
rect 126900 -8380 127100 -8120
rect 127400 -8380 127600 -8120
rect 127900 -8380 128100 -8120
rect 128400 -8380 128600 -8120
rect 128900 -8380 129100 -8120
rect 129400 -8380 129600 -8120
rect 129900 -8380 130100 -8120
rect 130400 -8380 130600 -8120
rect 130900 -8380 131100 -8120
rect 131400 -8380 131600 -8120
rect 131900 -8380 132100 -8120
rect 132400 -8380 132600 -8120
rect 132900 -8380 133100 -8120
rect 133400 -8380 133600 -8120
rect 133900 -8380 134100 -8120
rect 134400 -8380 134600 -8120
rect 134900 -8380 135100 -8120
rect 135400 -8380 135600 -8120
rect 135900 -8380 136100 -8120
rect 136400 -8380 136600 -8120
rect 136900 -8380 137100 -8120
rect 137400 -8380 137600 -8120
rect 137900 -8380 138100 -8120
rect 138400 -8380 138600 -8120
rect 138900 -8380 139100 -8120
rect 139400 -8380 139600 -8120
rect 139900 -8380 140000 -8120
rect 88000 -8400 88120 -8380
rect 88380 -8400 88620 -8380
rect 88880 -8400 89120 -8380
rect 89380 -8400 89620 -8380
rect 89880 -8400 90120 -8380
rect 90380 -8400 90620 -8380
rect 90880 -8400 91120 -8380
rect 91380 -8400 91620 -8380
rect 91880 -8400 92120 -8380
rect 92380 -8400 92620 -8380
rect 92880 -8400 93120 -8380
rect 93380 -8400 93620 -8380
rect 93880 -8400 94120 -8380
rect 94380 -8400 94620 -8380
rect 94880 -8400 95120 -8380
rect 95380 -8400 95620 -8380
rect 95880 -8400 96120 -8380
rect 96380 -8400 96620 -8380
rect 96880 -8400 97120 -8380
rect 97380 -8400 97620 -8380
rect 97880 -8400 98120 -8380
rect 98380 -8400 98620 -8380
rect 98880 -8400 99120 -8380
rect 99380 -8400 99620 -8380
rect 99880 -8400 100120 -8380
rect 100380 -8400 100620 -8380
rect 100880 -8400 101120 -8380
rect 101380 -8400 101620 -8380
rect 101880 -8400 102120 -8380
rect 102380 -8400 102620 -8380
rect 102880 -8400 103120 -8380
rect 103380 -8400 103620 -8380
rect 103880 -8400 104120 -8380
rect 104380 -8400 104620 -8380
rect 104880 -8400 105120 -8380
rect 105380 -8400 105620 -8380
rect 105880 -8400 106120 -8380
rect 106380 -8400 106620 -8380
rect 106880 -8400 107120 -8380
rect 107380 -8400 107620 -8380
rect 107880 -8400 108120 -8380
rect 108380 -8400 108620 -8380
rect 108880 -8400 109120 -8380
rect 109380 -8400 109620 -8380
rect 109880 -8400 110120 -8380
rect 110380 -8400 110620 -8380
rect 110880 -8400 111120 -8380
rect 111380 -8400 111620 -8380
rect 111880 -8400 112120 -8380
rect 112380 -8400 112620 -8380
rect 112880 -8400 113120 -8380
rect 113380 -8400 113620 -8380
rect 113880 -8400 114120 -8380
rect 114380 -8400 114620 -8380
rect 114880 -8400 115120 -8380
rect 115380 -8400 115620 -8380
rect 115880 -8400 116120 -8380
rect 116380 -8400 116620 -8380
rect 116880 -8400 117120 -8380
rect 117380 -8400 117620 -8380
rect 117880 -8400 118120 -8380
rect 118380 -8400 118620 -8380
rect 118880 -8400 119120 -8380
rect 119380 -8400 119620 -8380
rect 119880 -8400 120120 -8380
rect 120380 -8400 120620 -8380
rect 120880 -8400 121120 -8380
rect 121380 -8400 121620 -8380
rect 121880 -8400 122120 -8380
rect 122380 -8400 122620 -8380
rect 122880 -8400 123120 -8380
rect 123380 -8400 123620 -8380
rect 123880 -8400 124120 -8380
rect 124380 -8400 124620 -8380
rect 124880 -8400 125120 -8380
rect 125380 -8400 125620 -8380
rect 125880 -8400 126120 -8380
rect 126380 -8400 126620 -8380
rect 126880 -8400 127120 -8380
rect 127380 -8400 127620 -8380
rect 127880 -8400 128120 -8380
rect 128380 -8400 128620 -8380
rect 128880 -8400 129120 -8380
rect 129380 -8400 129620 -8380
rect 129880 -8400 130120 -8380
rect 130380 -8400 130620 -8380
rect 130880 -8400 131120 -8380
rect 131380 -8400 131620 -8380
rect 131880 -8400 132120 -8380
rect 132380 -8400 132620 -8380
rect 132880 -8400 133120 -8380
rect 133380 -8400 133620 -8380
rect 133880 -8400 134120 -8380
rect 134380 -8400 134620 -8380
rect 134880 -8400 135120 -8380
rect 135380 -8400 135620 -8380
rect 135880 -8400 136120 -8380
rect 136380 -8400 136620 -8380
rect 136880 -8400 137120 -8380
rect 137380 -8400 137620 -8380
rect 137880 -8400 138120 -8380
rect 138380 -8400 138620 -8380
rect 138880 -8400 139120 -8380
rect 139380 -8400 139620 -8380
rect 139880 -8400 140000 -8380
rect 88000 -8600 140000 -8400
rect 88000 -8620 88120 -8600
rect 88380 -8620 88620 -8600
rect 88880 -8620 89120 -8600
rect 89380 -8620 89620 -8600
rect 89880 -8620 90120 -8600
rect 90380 -8620 90620 -8600
rect 90880 -8620 91120 -8600
rect 91380 -8620 91620 -8600
rect 91880 -8620 92120 -8600
rect 92380 -8620 92620 -8600
rect 92880 -8620 93120 -8600
rect 93380 -8620 93620 -8600
rect 93880 -8620 94120 -8600
rect 94380 -8620 94620 -8600
rect 94880 -8620 95120 -8600
rect 95380 -8620 95620 -8600
rect 95880 -8620 96120 -8600
rect 96380 -8620 96620 -8600
rect 96880 -8620 97120 -8600
rect 97380 -8620 97620 -8600
rect 97880 -8620 98120 -8600
rect 98380 -8620 98620 -8600
rect 98880 -8620 99120 -8600
rect 99380 -8620 99620 -8600
rect 99880 -8620 100120 -8600
rect 100380 -8620 100620 -8600
rect 100880 -8620 101120 -8600
rect 101380 -8620 101620 -8600
rect 101880 -8620 102120 -8600
rect 102380 -8620 102620 -8600
rect 102880 -8620 103120 -8600
rect 103380 -8620 103620 -8600
rect 103880 -8620 104120 -8600
rect 104380 -8620 104620 -8600
rect 104880 -8620 105120 -8600
rect 105380 -8620 105620 -8600
rect 105880 -8620 106120 -8600
rect 106380 -8620 106620 -8600
rect 106880 -8620 107120 -8600
rect 107380 -8620 107620 -8600
rect 107880 -8620 108120 -8600
rect 108380 -8620 108620 -8600
rect 108880 -8620 109120 -8600
rect 109380 -8620 109620 -8600
rect 109880 -8620 110120 -8600
rect 110380 -8620 110620 -8600
rect 110880 -8620 111120 -8600
rect 111380 -8620 111620 -8600
rect 111880 -8620 112120 -8600
rect 112380 -8620 112620 -8600
rect 112880 -8620 113120 -8600
rect 113380 -8620 113620 -8600
rect 113880 -8620 114120 -8600
rect 114380 -8620 114620 -8600
rect 114880 -8620 115120 -8600
rect 115380 -8620 115620 -8600
rect 115880 -8620 116120 -8600
rect 116380 -8620 116620 -8600
rect 116880 -8620 117120 -8600
rect 117380 -8620 117620 -8600
rect 117880 -8620 118120 -8600
rect 118380 -8620 118620 -8600
rect 118880 -8620 119120 -8600
rect 119380 -8620 119620 -8600
rect 119880 -8620 120120 -8600
rect 120380 -8620 120620 -8600
rect 120880 -8620 121120 -8600
rect 121380 -8620 121620 -8600
rect 121880 -8620 122120 -8600
rect 122380 -8620 122620 -8600
rect 122880 -8620 123120 -8600
rect 123380 -8620 123620 -8600
rect 123880 -8620 124120 -8600
rect 124380 -8620 124620 -8600
rect 124880 -8620 125120 -8600
rect 125380 -8620 125620 -8600
rect 125880 -8620 126120 -8600
rect 126380 -8620 126620 -8600
rect 126880 -8620 127120 -8600
rect 127380 -8620 127620 -8600
rect 127880 -8620 128120 -8600
rect 128380 -8620 128620 -8600
rect 128880 -8620 129120 -8600
rect 129380 -8620 129620 -8600
rect 129880 -8620 130120 -8600
rect 130380 -8620 130620 -8600
rect 130880 -8620 131120 -8600
rect 131380 -8620 131620 -8600
rect 131880 -8620 132120 -8600
rect 132380 -8620 132620 -8600
rect 132880 -8620 133120 -8600
rect 133380 -8620 133620 -8600
rect 133880 -8620 134120 -8600
rect 134380 -8620 134620 -8600
rect 134880 -8620 135120 -8600
rect 135380 -8620 135620 -8600
rect 135880 -8620 136120 -8600
rect 136380 -8620 136620 -8600
rect 136880 -8620 137120 -8600
rect 137380 -8620 137620 -8600
rect 137880 -8620 138120 -8600
rect 138380 -8620 138620 -8600
rect 138880 -8620 139120 -8600
rect 139380 -8620 139620 -8600
rect 139880 -8620 140000 -8600
rect 88000 -8880 88100 -8620
rect 88400 -8880 88600 -8620
rect 88900 -8880 89100 -8620
rect 89400 -8880 89600 -8620
rect 89900 -8880 90100 -8620
rect 90400 -8880 90600 -8620
rect 90900 -8880 91100 -8620
rect 91400 -8880 91600 -8620
rect 91900 -8880 92100 -8620
rect 92400 -8880 92600 -8620
rect 92900 -8880 93100 -8620
rect 93400 -8880 93600 -8620
rect 93900 -8880 94100 -8620
rect 94400 -8880 94600 -8620
rect 94900 -8880 95100 -8620
rect 95400 -8880 95600 -8620
rect 95900 -8880 96100 -8620
rect 96400 -8880 96600 -8620
rect 96900 -8880 97100 -8620
rect 97400 -8880 97600 -8620
rect 97900 -8880 98100 -8620
rect 98400 -8880 98600 -8620
rect 98900 -8880 99100 -8620
rect 99400 -8880 99600 -8620
rect 99900 -8880 100100 -8620
rect 100400 -8880 100600 -8620
rect 100900 -8880 101100 -8620
rect 101400 -8880 101600 -8620
rect 101900 -8880 102100 -8620
rect 102400 -8880 102600 -8620
rect 102900 -8880 103100 -8620
rect 103400 -8880 103600 -8620
rect 103900 -8880 104100 -8620
rect 104400 -8880 104600 -8620
rect 104900 -8880 105100 -8620
rect 105400 -8880 105600 -8620
rect 105900 -8880 106100 -8620
rect 106400 -8880 106600 -8620
rect 106900 -8880 107100 -8620
rect 107400 -8880 107600 -8620
rect 107900 -8880 108100 -8620
rect 108400 -8880 108600 -8620
rect 108900 -8880 109100 -8620
rect 109400 -8880 109600 -8620
rect 109900 -8880 110100 -8620
rect 110400 -8880 110600 -8620
rect 110900 -8880 111100 -8620
rect 111400 -8880 111600 -8620
rect 111900 -8880 112100 -8620
rect 112400 -8880 112600 -8620
rect 112900 -8880 113100 -8620
rect 113400 -8880 113600 -8620
rect 113900 -8880 114100 -8620
rect 114400 -8880 114600 -8620
rect 114900 -8880 115100 -8620
rect 115400 -8880 115600 -8620
rect 115900 -8880 116100 -8620
rect 116400 -8880 116600 -8620
rect 116900 -8880 117100 -8620
rect 117400 -8880 117600 -8620
rect 117900 -8880 118100 -8620
rect 118400 -8880 118600 -8620
rect 118900 -8880 119100 -8620
rect 119400 -8880 119600 -8620
rect 119900 -8880 120100 -8620
rect 120400 -8880 120600 -8620
rect 120900 -8880 121100 -8620
rect 121400 -8880 121600 -8620
rect 121900 -8880 122100 -8620
rect 122400 -8880 122600 -8620
rect 122900 -8880 123100 -8620
rect 123400 -8880 123600 -8620
rect 123900 -8880 124100 -8620
rect 124400 -8880 124600 -8620
rect 124900 -8880 125100 -8620
rect 125400 -8880 125600 -8620
rect 125900 -8880 126100 -8620
rect 126400 -8880 126600 -8620
rect 126900 -8880 127100 -8620
rect 127400 -8880 127600 -8620
rect 127900 -8880 128100 -8620
rect 128400 -8880 128600 -8620
rect 128900 -8880 129100 -8620
rect 129400 -8880 129600 -8620
rect 129900 -8880 130100 -8620
rect 130400 -8880 130600 -8620
rect 130900 -8880 131100 -8620
rect 131400 -8880 131600 -8620
rect 131900 -8880 132100 -8620
rect 132400 -8880 132600 -8620
rect 132900 -8880 133100 -8620
rect 133400 -8880 133600 -8620
rect 133900 -8880 134100 -8620
rect 134400 -8880 134600 -8620
rect 134900 -8880 135100 -8620
rect 135400 -8880 135600 -8620
rect 135900 -8880 136100 -8620
rect 136400 -8880 136600 -8620
rect 136900 -8880 137100 -8620
rect 137400 -8880 137600 -8620
rect 137900 -8880 138100 -8620
rect 138400 -8880 138600 -8620
rect 138900 -8880 139100 -8620
rect 139400 -8880 139600 -8620
rect 139900 -8880 140000 -8620
rect 88000 -8900 88120 -8880
rect 88380 -8900 88620 -8880
rect 88880 -8900 89120 -8880
rect 89380 -8900 89620 -8880
rect 89880 -8900 90120 -8880
rect 90380 -8900 90620 -8880
rect 90880 -8900 91120 -8880
rect 91380 -8900 91620 -8880
rect 91880 -8900 92120 -8880
rect 92380 -8900 92620 -8880
rect 92880 -8900 93120 -8880
rect 93380 -8900 93620 -8880
rect 93880 -8900 94120 -8880
rect 94380 -8900 94620 -8880
rect 94880 -8900 95120 -8880
rect 95380 -8900 95620 -8880
rect 95880 -8900 96120 -8880
rect 96380 -8900 96620 -8880
rect 96880 -8900 97120 -8880
rect 97380 -8900 97620 -8880
rect 97880 -8900 98120 -8880
rect 98380 -8900 98620 -8880
rect 98880 -8900 99120 -8880
rect 99380 -8900 99620 -8880
rect 99880 -8900 100120 -8880
rect 100380 -8900 100620 -8880
rect 100880 -8900 101120 -8880
rect 101380 -8900 101620 -8880
rect 101880 -8900 102120 -8880
rect 102380 -8900 102620 -8880
rect 102880 -8900 103120 -8880
rect 103380 -8900 103620 -8880
rect 103880 -8900 104120 -8880
rect 104380 -8900 104620 -8880
rect 104880 -8900 105120 -8880
rect 105380 -8900 105620 -8880
rect 105880 -8900 106120 -8880
rect 106380 -8900 106620 -8880
rect 106880 -8900 107120 -8880
rect 107380 -8900 107620 -8880
rect 107880 -8900 108120 -8880
rect 108380 -8900 108620 -8880
rect 108880 -8900 109120 -8880
rect 109380 -8900 109620 -8880
rect 109880 -8900 110120 -8880
rect 110380 -8900 110620 -8880
rect 110880 -8900 111120 -8880
rect 111380 -8900 111620 -8880
rect 111880 -8900 112120 -8880
rect 112380 -8900 112620 -8880
rect 112880 -8900 113120 -8880
rect 113380 -8900 113620 -8880
rect 113880 -8900 114120 -8880
rect 114380 -8900 114620 -8880
rect 114880 -8900 115120 -8880
rect 115380 -8900 115620 -8880
rect 115880 -8900 116120 -8880
rect 116380 -8900 116620 -8880
rect 116880 -8900 117120 -8880
rect 117380 -8900 117620 -8880
rect 117880 -8900 118120 -8880
rect 118380 -8900 118620 -8880
rect 118880 -8900 119120 -8880
rect 119380 -8900 119620 -8880
rect 119880 -8900 120120 -8880
rect 120380 -8900 120620 -8880
rect 120880 -8900 121120 -8880
rect 121380 -8900 121620 -8880
rect 121880 -8900 122120 -8880
rect 122380 -8900 122620 -8880
rect 122880 -8900 123120 -8880
rect 123380 -8900 123620 -8880
rect 123880 -8900 124120 -8880
rect 124380 -8900 124620 -8880
rect 124880 -8900 125120 -8880
rect 125380 -8900 125620 -8880
rect 125880 -8900 126120 -8880
rect 126380 -8900 126620 -8880
rect 126880 -8900 127120 -8880
rect 127380 -8900 127620 -8880
rect 127880 -8900 128120 -8880
rect 128380 -8900 128620 -8880
rect 128880 -8900 129120 -8880
rect 129380 -8900 129620 -8880
rect 129880 -8900 130120 -8880
rect 130380 -8900 130620 -8880
rect 130880 -8900 131120 -8880
rect 131380 -8900 131620 -8880
rect 131880 -8900 132120 -8880
rect 132380 -8900 132620 -8880
rect 132880 -8900 133120 -8880
rect 133380 -8900 133620 -8880
rect 133880 -8900 134120 -8880
rect 134380 -8900 134620 -8880
rect 134880 -8900 135120 -8880
rect 135380 -8900 135620 -8880
rect 135880 -8900 136120 -8880
rect 136380 -8900 136620 -8880
rect 136880 -8900 137120 -8880
rect 137380 -8900 137620 -8880
rect 137880 -8900 138120 -8880
rect 138380 -8900 138620 -8880
rect 138880 -8900 139120 -8880
rect 139380 -8900 139620 -8880
rect 139880 -8900 140000 -8880
rect 88000 -9100 140000 -8900
rect 88000 -9120 88120 -9100
rect 88380 -9120 88620 -9100
rect 88880 -9120 89120 -9100
rect 89380 -9120 89620 -9100
rect 89880 -9120 90120 -9100
rect 90380 -9120 90620 -9100
rect 90880 -9120 91120 -9100
rect 91380 -9120 91620 -9100
rect 91880 -9120 92120 -9100
rect 92380 -9120 92620 -9100
rect 92880 -9120 93120 -9100
rect 93380 -9120 93620 -9100
rect 93880 -9120 94120 -9100
rect 94380 -9120 94620 -9100
rect 94880 -9120 95120 -9100
rect 95380 -9120 95620 -9100
rect 95880 -9120 96120 -9100
rect 96380 -9120 96620 -9100
rect 96880 -9120 97120 -9100
rect 97380 -9120 97620 -9100
rect 97880 -9120 98120 -9100
rect 98380 -9120 98620 -9100
rect 98880 -9120 99120 -9100
rect 99380 -9120 99620 -9100
rect 99880 -9120 100120 -9100
rect 100380 -9120 100620 -9100
rect 100880 -9120 101120 -9100
rect 101380 -9120 101620 -9100
rect 101880 -9120 102120 -9100
rect 102380 -9120 102620 -9100
rect 102880 -9120 103120 -9100
rect 103380 -9120 103620 -9100
rect 103880 -9120 104120 -9100
rect 104380 -9120 104620 -9100
rect 104880 -9120 105120 -9100
rect 105380 -9120 105620 -9100
rect 105880 -9120 106120 -9100
rect 106380 -9120 106620 -9100
rect 106880 -9120 107120 -9100
rect 107380 -9120 107620 -9100
rect 107880 -9120 108120 -9100
rect 108380 -9120 108620 -9100
rect 108880 -9120 109120 -9100
rect 109380 -9120 109620 -9100
rect 109880 -9120 110120 -9100
rect 110380 -9120 110620 -9100
rect 110880 -9120 111120 -9100
rect 111380 -9120 111620 -9100
rect 111880 -9120 112120 -9100
rect 112380 -9120 112620 -9100
rect 112880 -9120 113120 -9100
rect 113380 -9120 113620 -9100
rect 113880 -9120 114120 -9100
rect 114380 -9120 114620 -9100
rect 114880 -9120 115120 -9100
rect 115380 -9120 115620 -9100
rect 115880 -9120 116120 -9100
rect 116380 -9120 116620 -9100
rect 116880 -9120 117120 -9100
rect 117380 -9120 117620 -9100
rect 117880 -9120 118120 -9100
rect 118380 -9120 118620 -9100
rect 118880 -9120 119120 -9100
rect 119380 -9120 119620 -9100
rect 119880 -9120 120120 -9100
rect 120380 -9120 120620 -9100
rect 120880 -9120 121120 -9100
rect 121380 -9120 121620 -9100
rect 121880 -9120 122120 -9100
rect 122380 -9120 122620 -9100
rect 122880 -9120 123120 -9100
rect 123380 -9120 123620 -9100
rect 123880 -9120 124120 -9100
rect 124380 -9120 124620 -9100
rect 124880 -9120 125120 -9100
rect 125380 -9120 125620 -9100
rect 125880 -9120 126120 -9100
rect 126380 -9120 126620 -9100
rect 126880 -9120 127120 -9100
rect 127380 -9120 127620 -9100
rect 127880 -9120 128120 -9100
rect 128380 -9120 128620 -9100
rect 128880 -9120 129120 -9100
rect 129380 -9120 129620 -9100
rect 129880 -9120 130120 -9100
rect 130380 -9120 130620 -9100
rect 130880 -9120 131120 -9100
rect 131380 -9120 131620 -9100
rect 131880 -9120 132120 -9100
rect 132380 -9120 132620 -9100
rect 132880 -9120 133120 -9100
rect 133380 -9120 133620 -9100
rect 133880 -9120 134120 -9100
rect 134380 -9120 134620 -9100
rect 134880 -9120 135120 -9100
rect 135380 -9120 135620 -9100
rect 135880 -9120 136120 -9100
rect 136380 -9120 136620 -9100
rect 136880 -9120 137120 -9100
rect 137380 -9120 137620 -9100
rect 137880 -9120 138120 -9100
rect 138380 -9120 138620 -9100
rect 138880 -9120 139120 -9100
rect 139380 -9120 139620 -9100
rect 139880 -9120 140000 -9100
rect 88000 -9380 88100 -9120
rect 88400 -9380 88600 -9120
rect 88900 -9380 89100 -9120
rect 89400 -9380 89600 -9120
rect 89900 -9380 90100 -9120
rect 90400 -9380 90600 -9120
rect 90900 -9380 91100 -9120
rect 91400 -9380 91600 -9120
rect 91900 -9380 92100 -9120
rect 92400 -9380 92600 -9120
rect 92900 -9380 93100 -9120
rect 93400 -9380 93600 -9120
rect 93900 -9380 94100 -9120
rect 94400 -9380 94600 -9120
rect 94900 -9380 95100 -9120
rect 95400 -9380 95600 -9120
rect 95900 -9380 96100 -9120
rect 96400 -9380 96600 -9120
rect 96900 -9380 97100 -9120
rect 97400 -9380 97600 -9120
rect 97900 -9380 98100 -9120
rect 98400 -9380 98600 -9120
rect 98900 -9380 99100 -9120
rect 99400 -9380 99600 -9120
rect 99900 -9380 100100 -9120
rect 100400 -9380 100600 -9120
rect 100900 -9380 101100 -9120
rect 101400 -9380 101600 -9120
rect 101900 -9380 102100 -9120
rect 102400 -9380 102600 -9120
rect 102900 -9380 103100 -9120
rect 103400 -9380 103600 -9120
rect 103900 -9380 104100 -9120
rect 104400 -9380 104600 -9120
rect 104900 -9380 105100 -9120
rect 105400 -9380 105600 -9120
rect 105900 -9380 106100 -9120
rect 106400 -9380 106600 -9120
rect 106900 -9380 107100 -9120
rect 107400 -9380 107600 -9120
rect 107900 -9380 108100 -9120
rect 108400 -9380 108600 -9120
rect 108900 -9380 109100 -9120
rect 109400 -9380 109600 -9120
rect 109900 -9380 110100 -9120
rect 110400 -9380 110600 -9120
rect 110900 -9380 111100 -9120
rect 111400 -9380 111600 -9120
rect 111900 -9380 112100 -9120
rect 112400 -9380 112600 -9120
rect 112900 -9380 113100 -9120
rect 113400 -9380 113600 -9120
rect 113900 -9380 114100 -9120
rect 114400 -9380 114600 -9120
rect 114900 -9380 115100 -9120
rect 115400 -9380 115600 -9120
rect 115900 -9380 116100 -9120
rect 116400 -9380 116600 -9120
rect 116900 -9380 117100 -9120
rect 117400 -9380 117600 -9120
rect 117900 -9380 118100 -9120
rect 118400 -9380 118600 -9120
rect 118900 -9380 119100 -9120
rect 119400 -9380 119600 -9120
rect 119900 -9380 120100 -9120
rect 120400 -9380 120600 -9120
rect 120900 -9380 121100 -9120
rect 121400 -9380 121600 -9120
rect 121900 -9380 122100 -9120
rect 122400 -9380 122600 -9120
rect 122900 -9380 123100 -9120
rect 123400 -9380 123600 -9120
rect 123900 -9380 124100 -9120
rect 124400 -9380 124600 -9120
rect 124900 -9380 125100 -9120
rect 125400 -9380 125600 -9120
rect 125900 -9380 126100 -9120
rect 126400 -9380 126600 -9120
rect 126900 -9380 127100 -9120
rect 127400 -9380 127600 -9120
rect 127900 -9380 128100 -9120
rect 128400 -9380 128600 -9120
rect 128900 -9380 129100 -9120
rect 129400 -9380 129600 -9120
rect 129900 -9380 130100 -9120
rect 130400 -9380 130600 -9120
rect 130900 -9380 131100 -9120
rect 131400 -9380 131600 -9120
rect 131900 -9380 132100 -9120
rect 132400 -9380 132600 -9120
rect 132900 -9380 133100 -9120
rect 133400 -9380 133600 -9120
rect 133900 -9380 134100 -9120
rect 134400 -9380 134600 -9120
rect 134900 -9380 135100 -9120
rect 135400 -9380 135600 -9120
rect 135900 -9380 136100 -9120
rect 136400 -9380 136600 -9120
rect 136900 -9380 137100 -9120
rect 137400 -9380 137600 -9120
rect 137900 -9380 138100 -9120
rect 138400 -9380 138600 -9120
rect 138900 -9380 139100 -9120
rect 139400 -9380 139600 -9120
rect 139900 -9380 140000 -9120
rect 88000 -9400 88120 -9380
rect 88380 -9400 88620 -9380
rect 88880 -9400 89120 -9380
rect 89380 -9400 89620 -9380
rect 89880 -9400 90120 -9380
rect 90380 -9400 90620 -9380
rect 90880 -9400 91120 -9380
rect 91380 -9400 91620 -9380
rect 91880 -9400 92120 -9380
rect 92380 -9400 92620 -9380
rect 92880 -9400 93120 -9380
rect 93380 -9400 93620 -9380
rect 93880 -9400 94120 -9380
rect 94380 -9400 94620 -9380
rect 94880 -9400 95120 -9380
rect 95380 -9400 95620 -9380
rect 95880 -9400 96120 -9380
rect 96380 -9400 96620 -9380
rect 96880 -9400 97120 -9380
rect 97380 -9400 97620 -9380
rect 97880 -9400 98120 -9380
rect 98380 -9400 98620 -9380
rect 98880 -9400 99120 -9380
rect 99380 -9400 99620 -9380
rect 99880 -9400 100120 -9380
rect 100380 -9400 100620 -9380
rect 100880 -9400 101120 -9380
rect 101380 -9400 101620 -9380
rect 101880 -9400 102120 -9380
rect 102380 -9400 102620 -9380
rect 102880 -9400 103120 -9380
rect 103380 -9400 103620 -9380
rect 103880 -9400 104120 -9380
rect 104380 -9400 104620 -9380
rect 104880 -9400 105120 -9380
rect 105380 -9400 105620 -9380
rect 105880 -9400 106120 -9380
rect 106380 -9400 106620 -9380
rect 106880 -9400 107120 -9380
rect 107380 -9400 107620 -9380
rect 107880 -9400 108120 -9380
rect 108380 -9400 108620 -9380
rect 108880 -9400 109120 -9380
rect 109380 -9400 109620 -9380
rect 109880 -9400 110120 -9380
rect 110380 -9400 110620 -9380
rect 110880 -9400 111120 -9380
rect 111380 -9400 111620 -9380
rect 111880 -9400 112120 -9380
rect 112380 -9400 112620 -9380
rect 112880 -9400 113120 -9380
rect 113380 -9400 113620 -9380
rect 113880 -9400 114120 -9380
rect 114380 -9400 114620 -9380
rect 114880 -9400 115120 -9380
rect 115380 -9400 115620 -9380
rect 115880 -9400 116120 -9380
rect 116380 -9400 116620 -9380
rect 116880 -9400 117120 -9380
rect 117380 -9400 117620 -9380
rect 117880 -9400 118120 -9380
rect 118380 -9400 118620 -9380
rect 118880 -9400 119120 -9380
rect 119380 -9400 119620 -9380
rect 119880 -9400 120120 -9380
rect 120380 -9400 120620 -9380
rect 120880 -9400 121120 -9380
rect 121380 -9400 121620 -9380
rect 121880 -9400 122120 -9380
rect 122380 -9400 122620 -9380
rect 122880 -9400 123120 -9380
rect 123380 -9400 123620 -9380
rect 123880 -9400 124120 -9380
rect 124380 -9400 124620 -9380
rect 124880 -9400 125120 -9380
rect 125380 -9400 125620 -9380
rect 125880 -9400 126120 -9380
rect 126380 -9400 126620 -9380
rect 126880 -9400 127120 -9380
rect 127380 -9400 127620 -9380
rect 127880 -9400 128120 -9380
rect 128380 -9400 128620 -9380
rect 128880 -9400 129120 -9380
rect 129380 -9400 129620 -9380
rect 129880 -9400 130120 -9380
rect 130380 -9400 130620 -9380
rect 130880 -9400 131120 -9380
rect 131380 -9400 131620 -9380
rect 131880 -9400 132120 -9380
rect 132380 -9400 132620 -9380
rect 132880 -9400 133120 -9380
rect 133380 -9400 133620 -9380
rect 133880 -9400 134120 -9380
rect 134380 -9400 134620 -9380
rect 134880 -9400 135120 -9380
rect 135380 -9400 135620 -9380
rect 135880 -9400 136120 -9380
rect 136380 -9400 136620 -9380
rect 136880 -9400 137120 -9380
rect 137380 -9400 137620 -9380
rect 137880 -9400 138120 -9380
rect 138380 -9400 138620 -9380
rect 138880 -9400 139120 -9380
rect 139380 -9400 139620 -9380
rect 139880 -9400 140000 -9380
rect 88000 -9600 140000 -9400
rect 88000 -9620 88120 -9600
rect 88380 -9620 88620 -9600
rect 88880 -9620 89120 -9600
rect 89380 -9620 89620 -9600
rect 89880 -9620 90120 -9600
rect 90380 -9620 90620 -9600
rect 90880 -9620 91120 -9600
rect 91380 -9620 91620 -9600
rect 91880 -9620 92120 -9600
rect 92380 -9620 92620 -9600
rect 92880 -9620 93120 -9600
rect 93380 -9620 93620 -9600
rect 93880 -9620 94120 -9600
rect 94380 -9620 94620 -9600
rect 94880 -9620 95120 -9600
rect 95380 -9620 95620 -9600
rect 95880 -9620 96120 -9600
rect 96380 -9620 96620 -9600
rect 96880 -9620 97120 -9600
rect 97380 -9620 97620 -9600
rect 97880 -9620 98120 -9600
rect 98380 -9620 98620 -9600
rect 98880 -9620 99120 -9600
rect 99380 -9620 99620 -9600
rect 99880 -9620 100120 -9600
rect 100380 -9620 100620 -9600
rect 100880 -9620 101120 -9600
rect 101380 -9620 101620 -9600
rect 101880 -9620 102120 -9600
rect 102380 -9620 102620 -9600
rect 102880 -9620 103120 -9600
rect 103380 -9620 103620 -9600
rect 103880 -9620 104120 -9600
rect 104380 -9620 104620 -9600
rect 104880 -9620 105120 -9600
rect 105380 -9620 105620 -9600
rect 105880 -9620 106120 -9600
rect 106380 -9620 106620 -9600
rect 106880 -9620 107120 -9600
rect 107380 -9620 107620 -9600
rect 107880 -9620 108120 -9600
rect 108380 -9620 108620 -9600
rect 108880 -9620 109120 -9600
rect 109380 -9620 109620 -9600
rect 109880 -9620 110120 -9600
rect 110380 -9620 110620 -9600
rect 110880 -9620 111120 -9600
rect 111380 -9620 111620 -9600
rect 111880 -9620 112120 -9600
rect 112380 -9620 112620 -9600
rect 112880 -9620 113120 -9600
rect 113380 -9620 113620 -9600
rect 113880 -9620 114120 -9600
rect 114380 -9620 114620 -9600
rect 114880 -9620 115120 -9600
rect 115380 -9620 115620 -9600
rect 115880 -9620 116120 -9600
rect 116380 -9620 116620 -9600
rect 116880 -9620 117120 -9600
rect 117380 -9620 117620 -9600
rect 117880 -9620 118120 -9600
rect 118380 -9620 118620 -9600
rect 118880 -9620 119120 -9600
rect 119380 -9620 119620 -9600
rect 119880 -9620 120120 -9600
rect 120380 -9620 120620 -9600
rect 120880 -9620 121120 -9600
rect 121380 -9620 121620 -9600
rect 121880 -9620 122120 -9600
rect 122380 -9620 122620 -9600
rect 122880 -9620 123120 -9600
rect 123380 -9620 123620 -9600
rect 123880 -9620 124120 -9600
rect 124380 -9620 124620 -9600
rect 124880 -9620 125120 -9600
rect 125380 -9620 125620 -9600
rect 125880 -9620 126120 -9600
rect 126380 -9620 126620 -9600
rect 126880 -9620 127120 -9600
rect 127380 -9620 127620 -9600
rect 127880 -9620 128120 -9600
rect 128380 -9620 128620 -9600
rect 128880 -9620 129120 -9600
rect 129380 -9620 129620 -9600
rect 129880 -9620 130120 -9600
rect 130380 -9620 130620 -9600
rect 130880 -9620 131120 -9600
rect 131380 -9620 131620 -9600
rect 131880 -9620 132120 -9600
rect 132380 -9620 132620 -9600
rect 132880 -9620 133120 -9600
rect 133380 -9620 133620 -9600
rect 133880 -9620 134120 -9600
rect 134380 -9620 134620 -9600
rect 134880 -9620 135120 -9600
rect 135380 -9620 135620 -9600
rect 135880 -9620 136120 -9600
rect 136380 -9620 136620 -9600
rect 136880 -9620 137120 -9600
rect 137380 -9620 137620 -9600
rect 137880 -9620 138120 -9600
rect 138380 -9620 138620 -9600
rect 138880 -9620 139120 -9600
rect 139380 -9620 139620 -9600
rect 139880 -9620 140000 -9600
rect 88000 -9880 88100 -9620
rect 88400 -9880 88600 -9620
rect 88900 -9880 89100 -9620
rect 89400 -9880 89600 -9620
rect 89900 -9880 90100 -9620
rect 90400 -9880 90600 -9620
rect 90900 -9880 91100 -9620
rect 91400 -9880 91600 -9620
rect 91900 -9880 92100 -9620
rect 92400 -9880 92600 -9620
rect 92900 -9880 93100 -9620
rect 93400 -9880 93600 -9620
rect 93900 -9880 94100 -9620
rect 94400 -9880 94600 -9620
rect 94900 -9880 95100 -9620
rect 95400 -9880 95600 -9620
rect 95900 -9880 96100 -9620
rect 96400 -9880 96600 -9620
rect 96900 -9880 97100 -9620
rect 97400 -9880 97600 -9620
rect 97900 -9880 98100 -9620
rect 98400 -9880 98600 -9620
rect 98900 -9880 99100 -9620
rect 99400 -9880 99600 -9620
rect 99900 -9880 100100 -9620
rect 100400 -9880 100600 -9620
rect 100900 -9880 101100 -9620
rect 101400 -9880 101600 -9620
rect 101900 -9880 102100 -9620
rect 102400 -9880 102600 -9620
rect 102900 -9880 103100 -9620
rect 103400 -9880 103600 -9620
rect 103900 -9880 104100 -9620
rect 104400 -9880 104600 -9620
rect 104900 -9880 105100 -9620
rect 105400 -9880 105600 -9620
rect 105900 -9880 106100 -9620
rect 106400 -9880 106600 -9620
rect 106900 -9880 107100 -9620
rect 107400 -9880 107600 -9620
rect 107900 -9880 108100 -9620
rect 108400 -9880 108600 -9620
rect 108900 -9880 109100 -9620
rect 109400 -9880 109600 -9620
rect 109900 -9880 110100 -9620
rect 110400 -9880 110600 -9620
rect 110900 -9880 111100 -9620
rect 111400 -9880 111600 -9620
rect 111900 -9880 112100 -9620
rect 112400 -9880 112600 -9620
rect 112900 -9880 113100 -9620
rect 113400 -9880 113600 -9620
rect 113900 -9880 114100 -9620
rect 114400 -9880 114600 -9620
rect 114900 -9880 115100 -9620
rect 115400 -9880 115600 -9620
rect 115900 -9880 116100 -9620
rect 116400 -9880 116600 -9620
rect 116900 -9880 117100 -9620
rect 117400 -9880 117600 -9620
rect 117900 -9880 118100 -9620
rect 118400 -9880 118600 -9620
rect 118900 -9880 119100 -9620
rect 119400 -9880 119600 -9620
rect 119900 -9880 120100 -9620
rect 120400 -9880 120600 -9620
rect 120900 -9880 121100 -9620
rect 121400 -9880 121600 -9620
rect 121900 -9880 122100 -9620
rect 122400 -9880 122600 -9620
rect 122900 -9880 123100 -9620
rect 123400 -9880 123600 -9620
rect 123900 -9880 124100 -9620
rect 124400 -9880 124600 -9620
rect 124900 -9880 125100 -9620
rect 125400 -9880 125600 -9620
rect 125900 -9880 126100 -9620
rect 126400 -9880 126600 -9620
rect 126900 -9880 127100 -9620
rect 127400 -9880 127600 -9620
rect 127900 -9880 128100 -9620
rect 128400 -9880 128600 -9620
rect 128900 -9880 129100 -9620
rect 129400 -9880 129600 -9620
rect 129900 -9880 130100 -9620
rect 130400 -9880 130600 -9620
rect 130900 -9880 131100 -9620
rect 131400 -9880 131600 -9620
rect 131900 -9880 132100 -9620
rect 132400 -9880 132600 -9620
rect 132900 -9880 133100 -9620
rect 133400 -9880 133600 -9620
rect 133900 -9880 134100 -9620
rect 134400 -9880 134600 -9620
rect 134900 -9880 135100 -9620
rect 135400 -9880 135600 -9620
rect 135900 -9880 136100 -9620
rect 136400 -9880 136600 -9620
rect 136900 -9880 137100 -9620
rect 137400 -9880 137600 -9620
rect 137900 -9880 138100 -9620
rect 138400 -9880 138600 -9620
rect 138900 -9880 139100 -9620
rect 139400 -9880 139600 -9620
rect 139900 -9880 140000 -9620
rect 88000 -9900 88120 -9880
rect 88380 -9900 88620 -9880
rect 88880 -9900 89120 -9880
rect 89380 -9900 89620 -9880
rect 89880 -9900 90120 -9880
rect 90380 -9900 90620 -9880
rect 90880 -9900 91120 -9880
rect 91380 -9900 91620 -9880
rect 91880 -9900 92120 -9880
rect 92380 -9900 92620 -9880
rect 92880 -9900 93120 -9880
rect 93380 -9900 93620 -9880
rect 93880 -9900 94120 -9880
rect 94380 -9900 94620 -9880
rect 94880 -9900 95120 -9880
rect 95380 -9900 95620 -9880
rect 95880 -9900 96120 -9880
rect 96380 -9900 96620 -9880
rect 96880 -9900 97120 -9880
rect 97380 -9900 97620 -9880
rect 97880 -9900 98120 -9880
rect 98380 -9900 98620 -9880
rect 98880 -9900 99120 -9880
rect 99380 -9900 99620 -9880
rect 99880 -9900 100120 -9880
rect 100380 -9900 100620 -9880
rect 100880 -9900 101120 -9880
rect 101380 -9900 101620 -9880
rect 101880 -9900 102120 -9880
rect 102380 -9900 102620 -9880
rect 102880 -9900 103120 -9880
rect 103380 -9900 103620 -9880
rect 103880 -9900 104120 -9880
rect 104380 -9900 104620 -9880
rect 104880 -9900 105120 -9880
rect 105380 -9900 105620 -9880
rect 105880 -9900 106120 -9880
rect 106380 -9900 106620 -9880
rect 106880 -9900 107120 -9880
rect 107380 -9900 107620 -9880
rect 107880 -9900 108120 -9880
rect 108380 -9900 108620 -9880
rect 108880 -9900 109120 -9880
rect 109380 -9900 109620 -9880
rect 109880 -9900 110120 -9880
rect 110380 -9900 110620 -9880
rect 110880 -9900 111120 -9880
rect 111380 -9900 111620 -9880
rect 111880 -9900 112120 -9880
rect 112380 -9900 112620 -9880
rect 112880 -9900 113120 -9880
rect 113380 -9900 113620 -9880
rect 113880 -9900 114120 -9880
rect 114380 -9900 114620 -9880
rect 114880 -9900 115120 -9880
rect 115380 -9900 115620 -9880
rect 115880 -9900 116120 -9880
rect 116380 -9900 116620 -9880
rect 116880 -9900 117120 -9880
rect 117380 -9900 117620 -9880
rect 117880 -9900 118120 -9880
rect 118380 -9900 118620 -9880
rect 118880 -9900 119120 -9880
rect 119380 -9900 119620 -9880
rect 119880 -9900 120120 -9880
rect 120380 -9900 120620 -9880
rect 120880 -9900 121120 -9880
rect 121380 -9900 121620 -9880
rect 121880 -9900 122120 -9880
rect 122380 -9900 122620 -9880
rect 122880 -9900 123120 -9880
rect 123380 -9900 123620 -9880
rect 123880 -9900 124120 -9880
rect 124380 -9900 124620 -9880
rect 124880 -9900 125120 -9880
rect 125380 -9900 125620 -9880
rect 125880 -9900 126120 -9880
rect 126380 -9900 126620 -9880
rect 126880 -9900 127120 -9880
rect 127380 -9900 127620 -9880
rect 127880 -9900 128120 -9880
rect 128380 -9900 128620 -9880
rect 128880 -9900 129120 -9880
rect 129380 -9900 129620 -9880
rect 129880 -9900 130120 -9880
rect 130380 -9900 130620 -9880
rect 130880 -9900 131120 -9880
rect 131380 -9900 131620 -9880
rect 131880 -9900 132120 -9880
rect 132380 -9900 132620 -9880
rect 132880 -9900 133120 -9880
rect 133380 -9900 133620 -9880
rect 133880 -9900 134120 -9880
rect 134380 -9900 134620 -9880
rect 134880 -9900 135120 -9880
rect 135380 -9900 135620 -9880
rect 135880 -9900 136120 -9880
rect 136380 -9900 136620 -9880
rect 136880 -9900 137120 -9880
rect 137380 -9900 137620 -9880
rect 137880 -9900 138120 -9880
rect 138380 -9900 138620 -9880
rect 138880 -9900 139120 -9880
rect 139380 -9900 139620 -9880
rect 139880 -9900 140000 -9880
rect 88000 -10000 140000 -9900
rect 88000 -10100 90000 -10000
rect 88000 -10120 88120 -10100
rect 88380 -10120 88620 -10100
rect 88880 -10120 89120 -10100
rect 89380 -10120 89620 -10100
rect 89880 -10120 90000 -10100
rect 88000 -10380 88100 -10120
rect 88400 -10380 88600 -10120
rect 88900 -10380 89100 -10120
rect 89400 -10380 89600 -10120
rect 89900 -10380 90000 -10120
rect 88000 -10400 88120 -10380
rect 88380 -10400 88620 -10380
rect 88880 -10400 89120 -10380
rect 89380 -10400 89620 -10380
rect 89880 -10400 90000 -10380
rect 88000 -10600 90000 -10400
rect 88000 -10620 88120 -10600
rect 88380 -10620 88620 -10600
rect 88880 -10620 89120 -10600
rect 89380 -10620 89620 -10600
rect 89880 -10620 90000 -10600
rect 88000 -10880 88100 -10620
rect 88400 -10880 88600 -10620
rect 88900 -10880 89100 -10620
rect 89400 -10880 89600 -10620
rect 89900 -10880 90000 -10620
rect 88000 -10900 88120 -10880
rect 88380 -10900 88620 -10880
rect 88880 -10900 89120 -10880
rect 89380 -10900 89620 -10880
rect 89880 -10900 90000 -10880
rect 88000 -11100 90000 -10900
rect 88000 -11120 88120 -11100
rect 88380 -11120 88620 -11100
rect 88880 -11120 89120 -11100
rect 89380 -11120 89620 -11100
rect 89880 -11120 90000 -11100
rect 88000 -11380 88100 -11120
rect 88400 -11380 88600 -11120
rect 88900 -11380 89100 -11120
rect 89400 -11380 89600 -11120
rect 89900 -11380 90000 -11120
rect 88000 -11400 88120 -11380
rect 88380 -11400 88620 -11380
rect 88880 -11400 89120 -11380
rect 89380 -11400 89620 -11380
rect 89880 -11400 90000 -11380
rect 88000 -11600 90000 -11400
rect 88000 -11620 88120 -11600
rect 88380 -11620 88620 -11600
rect 88880 -11620 89120 -11600
rect 89380 -11620 89620 -11600
rect 89880 -11620 90000 -11600
rect 88000 -11880 88100 -11620
rect 88400 -11880 88600 -11620
rect 88900 -11880 89100 -11620
rect 89400 -11880 89600 -11620
rect 89900 -11880 90000 -11620
rect 88000 -11900 88120 -11880
rect 88380 -11900 88620 -11880
rect 88880 -11900 89120 -11880
rect 89380 -11900 89620 -11880
rect 89880 -11900 90000 -11880
rect 88000 -12100 90000 -11900
rect 88000 -12120 88120 -12100
rect 88380 -12120 88620 -12100
rect 88880 -12120 89120 -12100
rect 89380 -12120 89620 -12100
rect 89880 -12120 90000 -12100
rect 88000 -12380 88100 -12120
rect 88400 -12380 88600 -12120
rect 88900 -12380 89100 -12120
rect 89400 -12380 89600 -12120
rect 89900 -12380 90000 -12120
rect 88000 -12400 88120 -12380
rect 88380 -12400 88620 -12380
rect 88880 -12400 89120 -12380
rect 89380 -12400 89620 -12380
rect 89880 -12400 90000 -12380
rect 88000 -12600 90000 -12400
rect 88000 -12620 88120 -12600
rect 88380 -12620 88620 -12600
rect 88880 -12620 89120 -12600
rect 89380 -12620 89620 -12600
rect 89880 -12620 90000 -12600
rect 88000 -12880 88100 -12620
rect 88400 -12880 88600 -12620
rect 88900 -12880 89100 -12620
rect 89400 -12880 89600 -12620
rect 89900 -12880 90000 -12620
rect 88000 -12900 88120 -12880
rect 88380 -12900 88620 -12880
rect 88880 -12900 89120 -12880
rect 89380 -12900 89620 -12880
rect 89880 -12900 90000 -12880
rect 88000 -13100 90000 -12900
rect 88000 -13120 88120 -13100
rect 88380 -13120 88620 -13100
rect 88880 -13120 89120 -13100
rect 89380 -13120 89620 -13100
rect 89880 -13120 90000 -13100
rect 88000 -13380 88100 -13120
rect 88400 -13380 88600 -13120
rect 88900 -13380 89100 -13120
rect 89400 -13380 89600 -13120
rect 89900 -13380 90000 -13120
rect 88000 -13400 88120 -13380
rect 88380 -13400 88620 -13380
rect 88880 -13400 89120 -13380
rect 89380 -13400 89620 -13380
rect 89880 -13400 90000 -13380
rect 88000 -13600 90000 -13400
rect 88000 -13620 88120 -13600
rect 88380 -13620 88620 -13600
rect 88880 -13620 89120 -13600
rect 89380 -13620 89620 -13600
rect 89880 -13620 90000 -13600
rect 88000 -13880 88100 -13620
rect 88400 -13880 88600 -13620
rect 88900 -13880 89100 -13620
rect 89400 -13880 89600 -13620
rect 89900 -13880 90000 -13620
rect 88000 -13900 88120 -13880
rect 88380 -13900 88620 -13880
rect 88880 -13900 89120 -13880
rect 89380 -13900 89620 -13880
rect 89880 -13900 90000 -13880
rect 88000 -14000 90000 -13900
rect 92000 -10100 104000 -10000
rect 92000 -10120 92120 -10100
rect 92380 -10120 92620 -10100
rect 92880 -10120 93120 -10100
rect 93380 -10120 93620 -10100
rect 93880 -10120 94120 -10100
rect 94380 -10120 94620 -10100
rect 94880 -10120 95120 -10100
rect 95380 -10120 95620 -10100
rect 95880 -10120 96120 -10100
rect 96380 -10120 96620 -10100
rect 96880 -10120 97120 -10100
rect 97380 -10120 97620 -10100
rect 97880 -10120 98120 -10100
rect 98380 -10120 98620 -10100
rect 98880 -10120 99120 -10100
rect 99380 -10120 99620 -10100
rect 99880 -10120 100120 -10100
rect 100380 -10120 100620 -10100
rect 100880 -10120 101120 -10100
rect 101380 -10120 101620 -10100
rect 101880 -10120 102120 -10100
rect 102380 -10120 102620 -10100
rect 102880 -10120 103120 -10100
rect 103380 -10120 103620 -10100
rect 103880 -10120 104000 -10100
rect 92000 -10380 92100 -10120
rect 92400 -10380 92600 -10120
rect 92900 -10380 93100 -10120
rect 93400 -10380 93600 -10120
rect 93900 -10380 94100 -10120
rect 94400 -10380 94600 -10120
rect 94900 -10380 95100 -10120
rect 95400 -10380 95600 -10120
rect 95900 -10380 96100 -10120
rect 96400 -10380 96600 -10120
rect 96900 -10380 97100 -10120
rect 97400 -10380 97600 -10120
rect 97900 -10380 98100 -10120
rect 98400 -10380 98600 -10120
rect 98900 -10380 99100 -10120
rect 99400 -10380 99600 -10120
rect 99900 -10380 100100 -10120
rect 100400 -10380 100600 -10120
rect 100900 -10380 101100 -10120
rect 101400 -10380 101600 -10120
rect 101900 -10380 102100 -10120
rect 102400 -10380 102600 -10120
rect 102900 -10380 103100 -10120
rect 103400 -10380 103600 -10120
rect 103900 -10380 104000 -10120
rect 92000 -10400 92120 -10380
rect 92380 -10400 92620 -10380
rect 92880 -10400 93120 -10380
rect 93380 -10400 93620 -10380
rect 93880 -10400 94120 -10380
rect 94380 -10400 94620 -10380
rect 94880 -10400 95120 -10380
rect 95380 -10400 95620 -10380
rect 95880 -10400 96120 -10380
rect 96380 -10400 96620 -10380
rect 96880 -10400 97120 -10380
rect 97380 -10400 97620 -10380
rect 97880 -10400 98120 -10380
rect 98380 -10400 98620 -10380
rect 98880 -10400 99120 -10380
rect 99380 -10400 99620 -10380
rect 99880 -10400 100120 -10380
rect 100380 -10400 100620 -10380
rect 100880 -10400 101120 -10380
rect 101380 -10400 101620 -10380
rect 101880 -10400 102120 -10380
rect 102380 -10400 102620 -10380
rect 102880 -10400 103120 -10380
rect 103380 -10400 103620 -10380
rect 103880 -10400 104000 -10380
rect 92000 -10600 104000 -10400
rect 92000 -10620 92120 -10600
rect 92380 -10620 92620 -10600
rect 92880 -10620 93120 -10600
rect 93380 -10620 93620 -10600
rect 93880 -10620 94120 -10600
rect 94380 -10620 94620 -10600
rect 94880 -10620 95120 -10600
rect 95380 -10620 95620 -10600
rect 95880 -10620 96120 -10600
rect 96380 -10620 96620 -10600
rect 96880 -10620 97120 -10600
rect 97380 -10620 97620 -10600
rect 97880 -10620 98120 -10600
rect 98380 -10620 98620 -10600
rect 98880 -10620 99120 -10600
rect 99380 -10620 99620 -10600
rect 99880 -10620 100120 -10600
rect 100380 -10620 100620 -10600
rect 100880 -10620 101120 -10600
rect 101380 -10620 101620 -10600
rect 101880 -10620 102120 -10600
rect 102380 -10620 102620 -10600
rect 102880 -10620 103120 -10600
rect 103380 -10620 103620 -10600
rect 103880 -10620 104000 -10600
rect 92000 -10880 92100 -10620
rect 92400 -10880 92600 -10620
rect 92900 -10880 93100 -10620
rect 93400 -10880 93600 -10620
rect 93900 -10880 94100 -10620
rect 94400 -10880 94600 -10620
rect 94900 -10880 95100 -10620
rect 95400 -10880 95600 -10620
rect 95900 -10880 96100 -10620
rect 96400 -10880 96600 -10620
rect 96900 -10880 97100 -10620
rect 97400 -10880 97600 -10620
rect 97900 -10880 98100 -10620
rect 98400 -10880 98600 -10620
rect 98900 -10880 99100 -10620
rect 99400 -10880 99600 -10620
rect 99900 -10880 100100 -10620
rect 100400 -10880 100600 -10620
rect 100900 -10880 101100 -10620
rect 101400 -10880 101600 -10620
rect 101900 -10880 102100 -10620
rect 102400 -10880 102600 -10620
rect 102900 -10880 103100 -10620
rect 103400 -10880 103600 -10620
rect 103900 -10880 104000 -10620
rect 92000 -10900 92120 -10880
rect 92380 -10900 92620 -10880
rect 92880 -10900 93120 -10880
rect 93380 -10900 93620 -10880
rect 93880 -10900 94120 -10880
rect 94380 -10900 94620 -10880
rect 94880 -10900 95120 -10880
rect 95380 -10900 95620 -10880
rect 95880 -10900 96120 -10880
rect 96380 -10900 96620 -10880
rect 96880 -10900 97120 -10880
rect 97380 -10900 97620 -10880
rect 97880 -10900 98120 -10880
rect 98380 -10900 98620 -10880
rect 98880 -10900 99120 -10880
rect 99380 -10900 99620 -10880
rect 99880 -10900 100120 -10880
rect 100380 -10900 100620 -10880
rect 100880 -10900 101120 -10880
rect 101380 -10900 101620 -10880
rect 101880 -10900 102120 -10880
rect 102380 -10900 102620 -10880
rect 102880 -10900 103120 -10880
rect 103380 -10900 103620 -10880
rect 103880 -10900 104000 -10880
rect 92000 -11100 104000 -10900
rect 92000 -11120 92120 -11100
rect 92380 -11120 92620 -11100
rect 92880 -11120 93120 -11100
rect 93380 -11120 93620 -11100
rect 93880 -11120 94120 -11100
rect 94380 -11120 94620 -11100
rect 94880 -11120 95120 -11100
rect 95380 -11120 95620 -11100
rect 95880 -11120 96120 -11100
rect 96380 -11120 96620 -11100
rect 96880 -11120 97120 -11100
rect 97380 -11120 97620 -11100
rect 97880 -11120 98120 -11100
rect 98380 -11120 98620 -11100
rect 98880 -11120 99120 -11100
rect 99380 -11120 99620 -11100
rect 99880 -11120 100120 -11100
rect 100380 -11120 100620 -11100
rect 100880 -11120 101120 -11100
rect 101380 -11120 101620 -11100
rect 101880 -11120 102120 -11100
rect 102380 -11120 102620 -11100
rect 102880 -11120 103120 -11100
rect 103380 -11120 103620 -11100
rect 103880 -11120 104000 -11100
rect 92000 -11380 92100 -11120
rect 92400 -11380 92600 -11120
rect 92900 -11380 93100 -11120
rect 93400 -11380 93600 -11120
rect 93900 -11380 94100 -11120
rect 94400 -11380 94600 -11120
rect 94900 -11380 95100 -11120
rect 95400 -11380 95600 -11120
rect 95900 -11380 96100 -11120
rect 96400 -11380 96600 -11120
rect 96900 -11380 97100 -11120
rect 97400 -11380 97600 -11120
rect 97900 -11380 98100 -11120
rect 98400 -11380 98600 -11120
rect 98900 -11380 99100 -11120
rect 99400 -11380 99600 -11120
rect 99900 -11380 100100 -11120
rect 100400 -11380 100600 -11120
rect 100900 -11380 101100 -11120
rect 101400 -11380 101600 -11120
rect 101900 -11380 102100 -11120
rect 102400 -11380 102600 -11120
rect 102900 -11380 103100 -11120
rect 103400 -11380 103600 -11120
rect 103900 -11380 104000 -11120
rect 92000 -11400 92120 -11380
rect 92380 -11400 92620 -11380
rect 92880 -11400 93120 -11380
rect 93380 -11400 93620 -11380
rect 93880 -11400 94120 -11380
rect 94380 -11400 94620 -11380
rect 94880 -11400 95120 -11380
rect 95380 -11400 95620 -11380
rect 95880 -11400 96120 -11380
rect 96380 -11400 96620 -11380
rect 96880 -11400 97120 -11380
rect 97380 -11400 97620 -11380
rect 97880 -11400 98120 -11380
rect 98380 -11400 98620 -11380
rect 98880 -11400 99120 -11380
rect 99380 -11400 99620 -11380
rect 99880 -11400 100120 -11380
rect 100380 -11400 100620 -11380
rect 100880 -11400 101120 -11380
rect 101380 -11400 101620 -11380
rect 101880 -11400 102120 -11380
rect 102380 -11400 102620 -11380
rect 102880 -11400 103120 -11380
rect 103380 -11400 103620 -11380
rect 103880 -11400 104000 -11380
rect 92000 -11600 104000 -11400
rect 92000 -11620 92120 -11600
rect 92380 -11620 92620 -11600
rect 92880 -11620 93120 -11600
rect 93380 -11620 93620 -11600
rect 93880 -11620 94120 -11600
rect 94380 -11620 94620 -11600
rect 94880 -11620 95120 -11600
rect 95380 -11620 95620 -11600
rect 95880 -11620 96120 -11600
rect 96380 -11620 96620 -11600
rect 96880 -11620 97120 -11600
rect 97380 -11620 97620 -11600
rect 97880 -11620 98120 -11600
rect 98380 -11620 98620 -11600
rect 98880 -11620 99120 -11600
rect 99380 -11620 99620 -11600
rect 99880 -11620 100120 -11600
rect 100380 -11620 100620 -11600
rect 100880 -11620 101120 -11600
rect 101380 -11620 101620 -11600
rect 101880 -11620 102120 -11600
rect 102380 -11620 102620 -11600
rect 102880 -11620 103120 -11600
rect 103380 -11620 103620 -11600
rect 103880 -11620 104000 -11600
rect 92000 -11880 92100 -11620
rect 92400 -11880 92600 -11620
rect 92900 -11880 93100 -11620
rect 93400 -11880 93600 -11620
rect 93900 -11880 94100 -11620
rect 94400 -11880 94600 -11620
rect 94900 -11880 95100 -11620
rect 95400 -11880 95600 -11620
rect 95900 -11880 96100 -11620
rect 96400 -11880 96600 -11620
rect 96900 -11880 97100 -11620
rect 97400 -11880 97600 -11620
rect 97900 -11880 98100 -11620
rect 98400 -11880 98600 -11620
rect 98900 -11880 99100 -11620
rect 99400 -11880 99600 -11620
rect 99900 -11880 100100 -11620
rect 100400 -11880 100600 -11620
rect 100900 -11880 101100 -11620
rect 101400 -11880 101600 -11620
rect 101900 -11880 102100 -11620
rect 102400 -11880 102600 -11620
rect 102900 -11880 103100 -11620
rect 103400 -11880 103600 -11620
rect 103900 -11880 104000 -11620
rect 92000 -11900 92120 -11880
rect 92380 -11900 92620 -11880
rect 92880 -11900 93120 -11880
rect 93380 -11900 93620 -11880
rect 93880 -11900 94120 -11880
rect 94380 -11900 94620 -11880
rect 94880 -11900 95120 -11880
rect 95380 -11900 95620 -11880
rect 95880 -11900 96120 -11880
rect 96380 -11900 96620 -11880
rect 96880 -11900 97120 -11880
rect 97380 -11900 97620 -11880
rect 97880 -11900 98120 -11880
rect 98380 -11900 98620 -11880
rect 98880 -11900 99120 -11880
rect 99380 -11900 99620 -11880
rect 99880 -11900 100120 -11880
rect 100380 -11900 100620 -11880
rect 100880 -11900 101120 -11880
rect 101380 -11900 101620 -11880
rect 101880 -11900 102120 -11880
rect 102380 -11900 102620 -11880
rect 102880 -11900 103120 -11880
rect 103380 -11900 103620 -11880
rect 103880 -11900 104000 -11880
rect 92000 -12100 104000 -11900
rect 92000 -12120 92120 -12100
rect 92380 -12120 92620 -12100
rect 92880 -12120 93120 -12100
rect 93380 -12120 93620 -12100
rect 93880 -12120 94120 -12100
rect 94380 -12120 94620 -12100
rect 94880 -12120 95120 -12100
rect 95380 -12120 95620 -12100
rect 95880 -12120 96120 -12100
rect 96380 -12120 96620 -12100
rect 96880 -12120 97120 -12100
rect 97380 -12120 97620 -12100
rect 97880 -12120 98120 -12100
rect 98380 -12120 98620 -12100
rect 98880 -12120 99120 -12100
rect 99380 -12120 99620 -12100
rect 99880 -12120 100120 -12100
rect 100380 -12120 100620 -12100
rect 100880 -12120 101120 -12100
rect 101380 -12120 101620 -12100
rect 101880 -12120 102120 -12100
rect 102380 -12120 102620 -12100
rect 102880 -12120 103120 -12100
rect 103380 -12120 103620 -12100
rect 103880 -12120 104000 -12100
rect 92000 -12380 92100 -12120
rect 92400 -12380 92600 -12120
rect 92900 -12380 93100 -12120
rect 93400 -12380 93600 -12120
rect 93900 -12380 94100 -12120
rect 94400 -12380 94600 -12120
rect 94900 -12380 95100 -12120
rect 95400 -12380 95600 -12120
rect 95900 -12380 96100 -12120
rect 96400 -12380 96600 -12120
rect 96900 -12380 97100 -12120
rect 97400 -12380 97600 -12120
rect 97900 -12380 98100 -12120
rect 98400 -12380 98600 -12120
rect 98900 -12380 99100 -12120
rect 99400 -12380 99600 -12120
rect 99900 -12380 100100 -12120
rect 100400 -12380 100600 -12120
rect 100900 -12380 101100 -12120
rect 101400 -12380 101600 -12120
rect 101900 -12380 102100 -12120
rect 102400 -12380 102600 -12120
rect 102900 -12380 103100 -12120
rect 103400 -12380 103600 -12120
rect 103900 -12380 104000 -12120
rect 92000 -12400 92120 -12380
rect 92380 -12400 92620 -12380
rect 92880 -12400 93120 -12380
rect 93380 -12400 93620 -12380
rect 93880 -12400 94120 -12380
rect 94380 -12400 94620 -12380
rect 94880 -12400 95120 -12380
rect 95380 -12400 95620 -12380
rect 95880 -12400 96120 -12380
rect 96380 -12400 96620 -12380
rect 96880 -12400 97120 -12380
rect 97380 -12400 97620 -12380
rect 97880 -12400 98120 -12380
rect 98380 -12400 98620 -12380
rect 98880 -12400 99120 -12380
rect 99380 -12400 99620 -12380
rect 99880 -12400 100120 -12380
rect 100380 -12400 100620 -12380
rect 100880 -12400 101120 -12380
rect 101380 -12400 101620 -12380
rect 101880 -12400 102120 -12380
rect 102380 -12400 102620 -12380
rect 102880 -12400 103120 -12380
rect 103380 -12400 103620 -12380
rect 103880 -12400 104000 -12380
rect 92000 -12600 104000 -12400
rect 92000 -12620 92120 -12600
rect 92380 -12620 92620 -12600
rect 92880 -12620 93120 -12600
rect 93380 -12620 93620 -12600
rect 93880 -12620 94120 -12600
rect 94380 -12620 94620 -12600
rect 94880 -12620 95120 -12600
rect 95380 -12620 95620 -12600
rect 95880 -12620 96120 -12600
rect 96380 -12620 96620 -12600
rect 96880 -12620 97120 -12600
rect 97380 -12620 97620 -12600
rect 97880 -12620 98120 -12600
rect 98380 -12620 98620 -12600
rect 98880 -12620 99120 -12600
rect 99380 -12620 99620 -12600
rect 99880 -12620 100120 -12600
rect 100380 -12620 100620 -12600
rect 100880 -12620 101120 -12600
rect 101380 -12620 101620 -12600
rect 101880 -12620 102120 -12600
rect 102380 -12620 102620 -12600
rect 102880 -12620 103120 -12600
rect 103380 -12620 103620 -12600
rect 103880 -12620 104000 -12600
rect 92000 -12880 92100 -12620
rect 92400 -12880 92600 -12620
rect 92900 -12880 93100 -12620
rect 93400 -12880 93600 -12620
rect 93900 -12880 94100 -12620
rect 94400 -12880 94600 -12620
rect 94900 -12880 95100 -12620
rect 95400 -12880 95600 -12620
rect 95900 -12880 96100 -12620
rect 96400 -12880 96600 -12620
rect 96900 -12880 97100 -12620
rect 97400 -12880 97600 -12620
rect 97900 -12880 98100 -12620
rect 98400 -12880 98600 -12620
rect 98900 -12880 99100 -12620
rect 99400 -12880 99600 -12620
rect 99900 -12880 100100 -12620
rect 100400 -12880 100600 -12620
rect 100900 -12880 101100 -12620
rect 101400 -12880 101600 -12620
rect 101900 -12880 102100 -12620
rect 102400 -12880 102600 -12620
rect 102900 -12880 103100 -12620
rect 103400 -12880 103600 -12620
rect 103900 -12880 104000 -12620
rect 92000 -12900 92120 -12880
rect 92380 -12900 92620 -12880
rect 92880 -12900 93120 -12880
rect 93380 -12900 93620 -12880
rect 93880 -12900 94120 -12880
rect 94380 -12900 94620 -12880
rect 94880 -12900 95120 -12880
rect 95380 -12900 95620 -12880
rect 95880 -12900 96120 -12880
rect 96380 -12900 96620 -12880
rect 96880 -12900 97120 -12880
rect 97380 -12900 97620 -12880
rect 97880 -12900 98120 -12880
rect 98380 -12900 98620 -12880
rect 98880 -12900 99120 -12880
rect 99380 -12900 99620 -12880
rect 99880 -12900 100120 -12880
rect 100380 -12900 100620 -12880
rect 100880 -12900 101120 -12880
rect 101380 -12900 101620 -12880
rect 101880 -12900 102120 -12880
rect 102380 -12900 102620 -12880
rect 102880 -12900 103120 -12880
rect 103380 -12900 103620 -12880
rect 103880 -12900 104000 -12880
rect 92000 -13100 104000 -12900
rect 92000 -13120 92120 -13100
rect 92380 -13120 92620 -13100
rect 92880 -13120 93120 -13100
rect 93380 -13120 93620 -13100
rect 93880 -13120 94120 -13100
rect 94380 -13120 94620 -13100
rect 94880 -13120 95120 -13100
rect 95380 -13120 95620 -13100
rect 95880 -13120 96120 -13100
rect 96380 -13120 96620 -13100
rect 96880 -13120 97120 -13100
rect 97380 -13120 97620 -13100
rect 97880 -13120 98120 -13100
rect 98380 -13120 98620 -13100
rect 98880 -13120 99120 -13100
rect 99380 -13120 99620 -13100
rect 99880 -13120 100120 -13100
rect 100380 -13120 100620 -13100
rect 100880 -13120 101120 -13100
rect 101380 -13120 101620 -13100
rect 101880 -13120 102120 -13100
rect 102380 -13120 102620 -13100
rect 102880 -13120 103120 -13100
rect 103380 -13120 103620 -13100
rect 103880 -13120 104000 -13100
rect 92000 -13380 92100 -13120
rect 92400 -13380 92600 -13120
rect 92900 -13380 93100 -13120
rect 93400 -13380 93600 -13120
rect 93900 -13380 94100 -13120
rect 94400 -13380 94600 -13120
rect 94900 -13380 95100 -13120
rect 95400 -13380 95600 -13120
rect 95900 -13380 96100 -13120
rect 96400 -13380 96600 -13120
rect 96900 -13380 97100 -13120
rect 97400 -13380 97600 -13120
rect 97900 -13380 98100 -13120
rect 98400 -13380 98600 -13120
rect 98900 -13380 99100 -13120
rect 99400 -13380 99600 -13120
rect 99900 -13380 100100 -13120
rect 100400 -13380 100600 -13120
rect 100900 -13380 101100 -13120
rect 101400 -13380 101600 -13120
rect 101900 -13380 102100 -13120
rect 102400 -13380 102600 -13120
rect 102900 -13380 103100 -13120
rect 103400 -13380 103600 -13120
rect 103900 -13380 104000 -13120
rect 92000 -13400 92120 -13380
rect 92380 -13400 92620 -13380
rect 92880 -13400 93120 -13380
rect 93380 -13400 93620 -13380
rect 93880 -13400 94120 -13380
rect 94380 -13400 94620 -13380
rect 94880 -13400 95120 -13380
rect 95380 -13400 95620 -13380
rect 95880 -13400 96120 -13380
rect 96380 -13400 96620 -13380
rect 96880 -13400 97120 -13380
rect 97380 -13400 97620 -13380
rect 97880 -13400 98120 -13380
rect 98380 -13400 98620 -13380
rect 98880 -13400 99120 -13380
rect 99380 -13400 99620 -13380
rect 99880 -13400 100120 -13380
rect 100380 -13400 100620 -13380
rect 100880 -13400 101120 -13380
rect 101380 -13400 101620 -13380
rect 101880 -13400 102120 -13380
rect 102380 -13400 102620 -13380
rect 102880 -13400 103120 -13380
rect 103380 -13400 103620 -13380
rect 103880 -13400 104000 -13380
rect 92000 -13600 104000 -13400
rect 92000 -13620 92120 -13600
rect 92380 -13620 92620 -13600
rect 92880 -13620 93120 -13600
rect 93380 -13620 93620 -13600
rect 93880 -13620 94120 -13600
rect 94380 -13620 94620 -13600
rect 94880 -13620 95120 -13600
rect 95380 -13620 95620 -13600
rect 95880 -13620 96120 -13600
rect 96380 -13620 96620 -13600
rect 96880 -13620 97120 -13600
rect 97380 -13620 97620 -13600
rect 97880 -13620 98120 -13600
rect 98380 -13620 98620 -13600
rect 98880 -13620 99120 -13600
rect 99380 -13620 99620 -13600
rect 99880 -13620 100120 -13600
rect 100380 -13620 100620 -13600
rect 100880 -13620 101120 -13600
rect 101380 -13620 101620 -13600
rect 101880 -13620 102120 -13600
rect 102380 -13620 102620 -13600
rect 102880 -13620 103120 -13600
rect 103380 -13620 103620 -13600
rect 103880 -13620 104000 -13600
rect 92000 -13880 92100 -13620
rect 92400 -13880 92600 -13620
rect 92900 -13880 93100 -13620
rect 93400 -13880 93600 -13620
rect 93900 -13880 94100 -13620
rect 94400 -13880 94600 -13620
rect 94900 -13880 95100 -13620
rect 95400 -13880 95600 -13620
rect 95900 -13880 96100 -13620
rect 96400 -13880 96600 -13620
rect 96900 -13880 97100 -13620
rect 97400 -13880 97600 -13620
rect 97900 -13880 98100 -13620
rect 98400 -13880 98600 -13620
rect 98900 -13880 99100 -13620
rect 99400 -13880 99600 -13620
rect 99900 -13880 100100 -13620
rect 100400 -13880 100600 -13620
rect 100900 -13880 101100 -13620
rect 101400 -13880 101600 -13620
rect 101900 -13880 102100 -13620
rect 102400 -13880 102600 -13620
rect 102900 -13880 103100 -13620
rect 103400 -13880 103600 -13620
rect 103900 -13880 104000 -13620
rect 92000 -13900 92120 -13880
rect 92380 -13900 92620 -13880
rect 92880 -13900 93120 -13880
rect 93380 -13900 93620 -13880
rect 93880 -13900 94120 -13880
rect 94380 -13900 94620 -13880
rect 94880 -13900 95120 -13880
rect 95380 -13900 95620 -13880
rect 95880 -13900 96120 -13880
rect 96380 -13900 96620 -13880
rect 96880 -13900 97120 -13880
rect 97380 -13900 97620 -13880
rect 97880 -13900 98120 -13880
rect 98380 -13900 98620 -13880
rect 98880 -13900 99120 -13880
rect 99380 -13900 99620 -13880
rect 99880 -13900 100120 -13880
rect 100380 -13900 100620 -13880
rect 100880 -13900 101120 -13880
rect 101380 -13900 101620 -13880
rect 101880 -13900 102120 -13880
rect 102380 -13900 102620 -13880
rect 102880 -13900 103120 -13880
rect 103380 -13900 103620 -13880
rect 103880 -13900 104000 -13880
rect 92000 -14000 104000 -13900
rect 112000 -10100 140000 -10000
rect 112000 -10120 112120 -10100
rect 112380 -10120 112620 -10100
rect 112880 -10120 113120 -10100
rect 113380 -10120 113620 -10100
rect 113880 -10120 114120 -10100
rect 114380 -10120 114620 -10100
rect 114880 -10120 115120 -10100
rect 115380 -10120 115620 -10100
rect 115880 -10120 116120 -10100
rect 116380 -10120 116620 -10100
rect 116880 -10120 117120 -10100
rect 117380 -10120 117620 -10100
rect 117880 -10120 118120 -10100
rect 118380 -10120 118620 -10100
rect 118880 -10120 119120 -10100
rect 119380 -10120 119620 -10100
rect 119880 -10120 120120 -10100
rect 120380 -10120 120620 -10100
rect 120880 -10120 121120 -10100
rect 121380 -10120 121620 -10100
rect 121880 -10120 122120 -10100
rect 122380 -10120 122620 -10100
rect 122880 -10120 123120 -10100
rect 123380 -10120 123620 -10100
rect 123880 -10120 124120 -10100
rect 124380 -10120 124620 -10100
rect 124880 -10120 125120 -10100
rect 125380 -10120 125620 -10100
rect 125880 -10120 126120 -10100
rect 126380 -10120 126620 -10100
rect 126880 -10120 127120 -10100
rect 127380 -10120 127620 -10100
rect 127880 -10120 128120 -10100
rect 128380 -10120 128620 -10100
rect 128880 -10120 129120 -10100
rect 129380 -10120 129620 -10100
rect 129880 -10120 130120 -10100
rect 130380 -10120 130620 -10100
rect 130880 -10120 131120 -10100
rect 131380 -10120 131620 -10100
rect 131880 -10120 132120 -10100
rect 132380 -10120 132620 -10100
rect 132880 -10120 133120 -10100
rect 133380 -10120 133620 -10100
rect 133880 -10120 134120 -10100
rect 134380 -10120 134620 -10100
rect 134880 -10120 135120 -10100
rect 135380 -10120 135620 -10100
rect 135880 -10120 136120 -10100
rect 136380 -10120 136620 -10100
rect 136880 -10120 137120 -10100
rect 137380 -10120 137620 -10100
rect 137880 -10120 138120 -10100
rect 138380 -10120 138620 -10100
rect 138880 -10120 139120 -10100
rect 139380 -10120 139620 -10100
rect 139880 -10120 140000 -10100
rect 112000 -10380 112100 -10120
rect 112400 -10380 112600 -10120
rect 112900 -10380 113100 -10120
rect 113400 -10380 113600 -10120
rect 113900 -10380 114100 -10120
rect 114400 -10380 114600 -10120
rect 114900 -10380 115100 -10120
rect 115400 -10380 115600 -10120
rect 115900 -10380 116100 -10120
rect 116400 -10380 116600 -10120
rect 116900 -10380 117100 -10120
rect 117400 -10380 117600 -10120
rect 117900 -10380 118100 -10120
rect 118400 -10380 118600 -10120
rect 118900 -10380 119100 -10120
rect 119400 -10380 119600 -10120
rect 119900 -10380 120100 -10120
rect 120400 -10380 120600 -10120
rect 120900 -10380 121100 -10120
rect 121400 -10380 121600 -10120
rect 121900 -10380 122100 -10120
rect 122400 -10380 122600 -10120
rect 122900 -10380 123100 -10120
rect 123400 -10380 123600 -10120
rect 123900 -10380 124100 -10120
rect 124400 -10380 124600 -10120
rect 124900 -10380 125100 -10120
rect 125400 -10380 125600 -10120
rect 125900 -10380 126100 -10120
rect 126400 -10380 126600 -10120
rect 126900 -10380 127100 -10120
rect 127400 -10380 127600 -10120
rect 127900 -10380 128100 -10120
rect 128400 -10380 128600 -10120
rect 128900 -10380 129100 -10120
rect 129400 -10380 129600 -10120
rect 129900 -10380 130100 -10120
rect 130400 -10380 130600 -10120
rect 130900 -10380 131100 -10120
rect 131400 -10380 131600 -10120
rect 131900 -10380 132100 -10120
rect 132400 -10380 132600 -10120
rect 132900 -10380 133100 -10120
rect 133400 -10380 133600 -10120
rect 133900 -10380 134100 -10120
rect 134400 -10380 134600 -10120
rect 134900 -10380 135100 -10120
rect 135400 -10380 135600 -10120
rect 135900 -10380 136100 -10120
rect 136400 -10380 136600 -10120
rect 136900 -10380 137100 -10120
rect 137400 -10380 137600 -10120
rect 137900 -10380 138100 -10120
rect 138400 -10380 138600 -10120
rect 138900 -10380 139100 -10120
rect 139400 -10380 139600 -10120
rect 139900 -10380 140000 -10120
rect 112000 -10400 112120 -10380
rect 112380 -10400 112620 -10380
rect 112880 -10400 113120 -10380
rect 113380 -10400 113620 -10380
rect 113880 -10400 114120 -10380
rect 114380 -10400 114620 -10380
rect 114880 -10400 115120 -10380
rect 115380 -10400 115620 -10380
rect 115880 -10400 116120 -10380
rect 116380 -10400 116620 -10380
rect 116880 -10400 117120 -10380
rect 117380 -10400 117620 -10380
rect 117880 -10400 118120 -10380
rect 118380 -10400 118620 -10380
rect 118880 -10400 119120 -10380
rect 119380 -10400 119620 -10380
rect 119880 -10400 120120 -10380
rect 120380 -10400 120620 -10380
rect 120880 -10400 121120 -10380
rect 121380 -10400 121620 -10380
rect 121880 -10400 122120 -10380
rect 122380 -10400 122620 -10380
rect 122880 -10400 123120 -10380
rect 123380 -10400 123620 -10380
rect 123880 -10400 124120 -10380
rect 124380 -10400 124620 -10380
rect 124880 -10400 125120 -10380
rect 125380 -10400 125620 -10380
rect 125880 -10400 126120 -10380
rect 126380 -10400 126620 -10380
rect 126880 -10400 127120 -10380
rect 127380 -10400 127620 -10380
rect 127880 -10400 128120 -10380
rect 128380 -10400 128620 -10380
rect 128880 -10400 129120 -10380
rect 129380 -10400 129620 -10380
rect 129880 -10400 130120 -10380
rect 130380 -10400 130620 -10380
rect 130880 -10400 131120 -10380
rect 131380 -10400 131620 -10380
rect 131880 -10400 132120 -10380
rect 132380 -10400 132620 -10380
rect 132880 -10400 133120 -10380
rect 133380 -10400 133620 -10380
rect 133880 -10400 134120 -10380
rect 134380 -10400 134620 -10380
rect 134880 -10400 135120 -10380
rect 135380 -10400 135620 -10380
rect 135880 -10400 136120 -10380
rect 136380 -10400 136620 -10380
rect 136880 -10400 137120 -10380
rect 137380 -10400 137620 -10380
rect 137880 -10400 138120 -10380
rect 138380 -10400 138620 -10380
rect 138880 -10400 139120 -10380
rect 139380 -10400 139620 -10380
rect 139880 -10400 140000 -10380
rect 112000 -10600 140000 -10400
rect 112000 -10620 112120 -10600
rect 112380 -10620 112620 -10600
rect 112880 -10620 113120 -10600
rect 113380 -10620 113620 -10600
rect 113880 -10620 114120 -10600
rect 114380 -10620 114620 -10600
rect 114880 -10620 115120 -10600
rect 115380 -10620 115620 -10600
rect 115880 -10620 116120 -10600
rect 116380 -10620 116620 -10600
rect 116880 -10620 117120 -10600
rect 117380 -10620 117620 -10600
rect 117880 -10620 118120 -10600
rect 118380 -10620 118620 -10600
rect 118880 -10620 119120 -10600
rect 119380 -10620 119620 -10600
rect 119880 -10620 120120 -10600
rect 120380 -10620 120620 -10600
rect 120880 -10620 121120 -10600
rect 121380 -10620 121620 -10600
rect 121880 -10620 122120 -10600
rect 122380 -10620 122620 -10600
rect 122880 -10620 123120 -10600
rect 123380 -10620 123620 -10600
rect 123880 -10620 124120 -10600
rect 124380 -10620 124620 -10600
rect 124880 -10620 125120 -10600
rect 125380 -10620 125620 -10600
rect 125880 -10620 126120 -10600
rect 126380 -10620 126620 -10600
rect 126880 -10620 127120 -10600
rect 127380 -10620 127620 -10600
rect 127880 -10620 128120 -10600
rect 128380 -10620 128620 -10600
rect 128880 -10620 129120 -10600
rect 129380 -10620 129620 -10600
rect 129880 -10620 130120 -10600
rect 130380 -10620 130620 -10600
rect 130880 -10620 131120 -10600
rect 131380 -10620 131620 -10600
rect 131880 -10620 132120 -10600
rect 132380 -10620 132620 -10600
rect 132880 -10620 133120 -10600
rect 133380 -10620 133620 -10600
rect 133880 -10620 134120 -10600
rect 134380 -10620 134620 -10600
rect 134880 -10620 135120 -10600
rect 135380 -10620 135620 -10600
rect 135880 -10620 136120 -10600
rect 136380 -10620 136620 -10600
rect 136880 -10620 137120 -10600
rect 137380 -10620 137620 -10600
rect 137880 -10620 138120 -10600
rect 138380 -10620 138620 -10600
rect 138880 -10620 139120 -10600
rect 139380 -10620 139620 -10600
rect 139880 -10620 140000 -10600
rect 112000 -10880 112100 -10620
rect 112400 -10880 112600 -10620
rect 112900 -10880 113100 -10620
rect 113400 -10880 113600 -10620
rect 113900 -10880 114100 -10620
rect 114400 -10880 114600 -10620
rect 114900 -10880 115100 -10620
rect 115400 -10880 115600 -10620
rect 115900 -10880 116100 -10620
rect 116400 -10880 116600 -10620
rect 116900 -10880 117100 -10620
rect 117400 -10880 117600 -10620
rect 117900 -10880 118100 -10620
rect 118400 -10880 118600 -10620
rect 118900 -10880 119100 -10620
rect 119400 -10880 119600 -10620
rect 119900 -10880 120100 -10620
rect 120400 -10880 120600 -10620
rect 120900 -10880 121100 -10620
rect 121400 -10880 121600 -10620
rect 121900 -10880 122100 -10620
rect 122400 -10880 122600 -10620
rect 122900 -10880 123100 -10620
rect 123400 -10880 123600 -10620
rect 123900 -10880 124100 -10620
rect 124400 -10880 124600 -10620
rect 124900 -10880 125100 -10620
rect 125400 -10880 125600 -10620
rect 125900 -10880 126100 -10620
rect 126400 -10880 126600 -10620
rect 126900 -10880 127100 -10620
rect 127400 -10880 127600 -10620
rect 127900 -10880 128100 -10620
rect 128400 -10880 128600 -10620
rect 128900 -10880 129100 -10620
rect 129400 -10880 129600 -10620
rect 129900 -10880 130100 -10620
rect 130400 -10880 130600 -10620
rect 130900 -10880 131100 -10620
rect 131400 -10880 131600 -10620
rect 131900 -10880 132100 -10620
rect 132400 -10880 132600 -10620
rect 132900 -10880 133100 -10620
rect 133400 -10880 133600 -10620
rect 133900 -10880 134100 -10620
rect 134400 -10880 134600 -10620
rect 134900 -10880 135100 -10620
rect 135400 -10880 135600 -10620
rect 135900 -10880 136100 -10620
rect 136400 -10880 136600 -10620
rect 136900 -10880 137100 -10620
rect 137400 -10880 137600 -10620
rect 137900 -10880 138100 -10620
rect 138400 -10880 138600 -10620
rect 138900 -10880 139100 -10620
rect 139400 -10880 139600 -10620
rect 139900 -10880 140000 -10620
rect 112000 -10900 112120 -10880
rect 112380 -10900 112620 -10880
rect 112880 -10900 113120 -10880
rect 113380 -10900 113620 -10880
rect 113880 -10900 114120 -10880
rect 114380 -10900 114620 -10880
rect 114880 -10900 115120 -10880
rect 115380 -10900 115620 -10880
rect 115880 -10900 116120 -10880
rect 116380 -10900 116620 -10880
rect 116880 -10900 117120 -10880
rect 117380 -10900 117620 -10880
rect 117880 -10900 118120 -10880
rect 118380 -10900 118620 -10880
rect 118880 -10900 119120 -10880
rect 119380 -10900 119620 -10880
rect 119880 -10900 120120 -10880
rect 120380 -10900 120620 -10880
rect 120880 -10900 121120 -10880
rect 121380 -10900 121620 -10880
rect 121880 -10900 122120 -10880
rect 122380 -10900 122620 -10880
rect 122880 -10900 123120 -10880
rect 123380 -10900 123620 -10880
rect 123880 -10900 124120 -10880
rect 124380 -10900 124620 -10880
rect 124880 -10900 125120 -10880
rect 125380 -10900 125620 -10880
rect 125880 -10900 126120 -10880
rect 126380 -10900 126620 -10880
rect 126880 -10900 127120 -10880
rect 127380 -10900 127620 -10880
rect 127880 -10900 128120 -10880
rect 128380 -10900 128620 -10880
rect 128880 -10900 129120 -10880
rect 129380 -10900 129620 -10880
rect 129880 -10900 130120 -10880
rect 130380 -10900 130620 -10880
rect 130880 -10900 131120 -10880
rect 131380 -10900 131620 -10880
rect 131880 -10900 132120 -10880
rect 132380 -10900 132620 -10880
rect 132880 -10900 133120 -10880
rect 133380 -10900 133620 -10880
rect 133880 -10900 134120 -10880
rect 134380 -10900 134620 -10880
rect 134880 -10900 135120 -10880
rect 135380 -10900 135620 -10880
rect 135880 -10900 136120 -10880
rect 136380 -10900 136620 -10880
rect 136880 -10900 137120 -10880
rect 137380 -10900 137620 -10880
rect 137880 -10900 138120 -10880
rect 138380 -10900 138620 -10880
rect 138880 -10900 139120 -10880
rect 139380 -10900 139620 -10880
rect 139880 -10900 140000 -10880
rect 112000 -11100 140000 -10900
rect 112000 -11120 112120 -11100
rect 112380 -11120 112620 -11100
rect 112880 -11120 113120 -11100
rect 113380 -11120 113620 -11100
rect 113880 -11120 114120 -11100
rect 114380 -11120 114620 -11100
rect 114880 -11120 115120 -11100
rect 115380 -11120 115620 -11100
rect 115880 -11120 116120 -11100
rect 116380 -11120 116620 -11100
rect 116880 -11120 117120 -11100
rect 117380 -11120 117620 -11100
rect 117880 -11120 118120 -11100
rect 118380 -11120 118620 -11100
rect 118880 -11120 119120 -11100
rect 119380 -11120 119620 -11100
rect 119880 -11120 120120 -11100
rect 120380 -11120 120620 -11100
rect 120880 -11120 121120 -11100
rect 121380 -11120 121620 -11100
rect 121880 -11120 122120 -11100
rect 122380 -11120 122620 -11100
rect 122880 -11120 123120 -11100
rect 123380 -11120 123620 -11100
rect 123880 -11120 124120 -11100
rect 124380 -11120 124620 -11100
rect 124880 -11120 125120 -11100
rect 125380 -11120 125620 -11100
rect 125880 -11120 126120 -11100
rect 126380 -11120 126620 -11100
rect 126880 -11120 127120 -11100
rect 127380 -11120 127620 -11100
rect 127880 -11120 128120 -11100
rect 128380 -11120 128620 -11100
rect 128880 -11120 129120 -11100
rect 129380 -11120 129620 -11100
rect 129880 -11120 130120 -11100
rect 130380 -11120 130620 -11100
rect 130880 -11120 131120 -11100
rect 131380 -11120 131620 -11100
rect 131880 -11120 132120 -11100
rect 132380 -11120 132620 -11100
rect 132880 -11120 133120 -11100
rect 133380 -11120 133620 -11100
rect 133880 -11120 134120 -11100
rect 134380 -11120 134620 -11100
rect 134880 -11120 135120 -11100
rect 135380 -11120 135620 -11100
rect 135880 -11120 136120 -11100
rect 136380 -11120 136620 -11100
rect 136880 -11120 137120 -11100
rect 137380 -11120 137620 -11100
rect 137880 -11120 138120 -11100
rect 138380 -11120 138620 -11100
rect 138880 -11120 139120 -11100
rect 139380 -11120 139620 -11100
rect 139880 -11120 140000 -11100
rect 112000 -11380 112100 -11120
rect 112400 -11380 112600 -11120
rect 112900 -11380 113100 -11120
rect 113400 -11380 113600 -11120
rect 113900 -11380 114100 -11120
rect 114400 -11380 114600 -11120
rect 114900 -11380 115100 -11120
rect 115400 -11380 115600 -11120
rect 115900 -11380 116100 -11120
rect 116400 -11380 116600 -11120
rect 116900 -11380 117100 -11120
rect 117400 -11380 117600 -11120
rect 117900 -11380 118100 -11120
rect 118400 -11380 118600 -11120
rect 118900 -11380 119100 -11120
rect 119400 -11380 119600 -11120
rect 119900 -11380 120100 -11120
rect 120400 -11380 120600 -11120
rect 120900 -11380 121100 -11120
rect 121400 -11380 121600 -11120
rect 121900 -11380 122100 -11120
rect 122400 -11380 122600 -11120
rect 122900 -11380 123100 -11120
rect 123400 -11380 123600 -11120
rect 123900 -11380 124100 -11120
rect 124400 -11380 124600 -11120
rect 124900 -11380 125100 -11120
rect 125400 -11380 125600 -11120
rect 125900 -11380 126100 -11120
rect 126400 -11380 126600 -11120
rect 126900 -11380 127100 -11120
rect 127400 -11380 127600 -11120
rect 127900 -11380 128100 -11120
rect 128400 -11380 128600 -11120
rect 128900 -11380 129100 -11120
rect 129400 -11380 129600 -11120
rect 129900 -11380 130100 -11120
rect 130400 -11380 130600 -11120
rect 130900 -11380 131100 -11120
rect 131400 -11380 131600 -11120
rect 131900 -11380 132100 -11120
rect 132400 -11380 132600 -11120
rect 132900 -11380 133100 -11120
rect 133400 -11380 133600 -11120
rect 133900 -11380 134100 -11120
rect 134400 -11380 134600 -11120
rect 134900 -11380 135100 -11120
rect 135400 -11380 135600 -11120
rect 135900 -11380 136100 -11120
rect 136400 -11380 136600 -11120
rect 136900 -11380 137100 -11120
rect 137400 -11380 137600 -11120
rect 137900 -11380 138100 -11120
rect 138400 -11380 138600 -11120
rect 138900 -11380 139100 -11120
rect 139400 -11380 139600 -11120
rect 139900 -11380 140000 -11120
rect 112000 -11400 112120 -11380
rect 112380 -11400 112620 -11380
rect 112880 -11400 113120 -11380
rect 113380 -11400 113620 -11380
rect 113880 -11400 114120 -11380
rect 114380 -11400 114620 -11380
rect 114880 -11400 115120 -11380
rect 115380 -11400 115620 -11380
rect 115880 -11400 116120 -11380
rect 116380 -11400 116620 -11380
rect 116880 -11400 117120 -11380
rect 117380 -11400 117620 -11380
rect 117880 -11400 118120 -11380
rect 118380 -11400 118620 -11380
rect 118880 -11400 119120 -11380
rect 119380 -11400 119620 -11380
rect 119880 -11400 120120 -11380
rect 120380 -11400 120620 -11380
rect 120880 -11400 121120 -11380
rect 121380 -11400 121620 -11380
rect 121880 -11400 122120 -11380
rect 122380 -11400 122620 -11380
rect 122880 -11400 123120 -11380
rect 123380 -11400 123620 -11380
rect 123880 -11400 124120 -11380
rect 124380 -11400 124620 -11380
rect 124880 -11400 125120 -11380
rect 125380 -11400 125620 -11380
rect 125880 -11400 126120 -11380
rect 126380 -11400 126620 -11380
rect 126880 -11400 127120 -11380
rect 127380 -11400 127620 -11380
rect 127880 -11400 128120 -11380
rect 128380 -11400 128620 -11380
rect 128880 -11400 129120 -11380
rect 129380 -11400 129620 -11380
rect 129880 -11400 130120 -11380
rect 130380 -11400 130620 -11380
rect 130880 -11400 131120 -11380
rect 131380 -11400 131620 -11380
rect 131880 -11400 132120 -11380
rect 132380 -11400 132620 -11380
rect 132880 -11400 133120 -11380
rect 133380 -11400 133620 -11380
rect 133880 -11400 134120 -11380
rect 134380 -11400 134620 -11380
rect 134880 -11400 135120 -11380
rect 135380 -11400 135620 -11380
rect 135880 -11400 136120 -11380
rect 136380 -11400 136620 -11380
rect 136880 -11400 137120 -11380
rect 137380 -11400 137620 -11380
rect 137880 -11400 138120 -11380
rect 138380 -11400 138620 -11380
rect 138880 -11400 139120 -11380
rect 139380 -11400 139620 -11380
rect 139880 -11400 140000 -11380
rect 112000 -11600 140000 -11400
rect 112000 -11620 112120 -11600
rect 112380 -11620 112620 -11600
rect 112880 -11620 113120 -11600
rect 113380 -11620 113620 -11600
rect 113880 -11620 114120 -11600
rect 114380 -11620 114620 -11600
rect 114880 -11620 115120 -11600
rect 115380 -11620 115620 -11600
rect 115880 -11620 116120 -11600
rect 116380 -11620 116620 -11600
rect 116880 -11620 117120 -11600
rect 117380 -11620 117620 -11600
rect 117880 -11620 118120 -11600
rect 118380 -11620 118620 -11600
rect 118880 -11620 119120 -11600
rect 119380 -11620 119620 -11600
rect 119880 -11620 120120 -11600
rect 120380 -11620 120620 -11600
rect 120880 -11620 121120 -11600
rect 121380 -11620 121620 -11600
rect 121880 -11620 122120 -11600
rect 122380 -11620 122620 -11600
rect 122880 -11620 123120 -11600
rect 123380 -11620 123620 -11600
rect 123880 -11620 124120 -11600
rect 124380 -11620 124620 -11600
rect 124880 -11620 125120 -11600
rect 125380 -11620 125620 -11600
rect 125880 -11620 126120 -11600
rect 126380 -11620 126620 -11600
rect 126880 -11620 127120 -11600
rect 127380 -11620 127620 -11600
rect 127880 -11620 128120 -11600
rect 128380 -11620 128620 -11600
rect 128880 -11620 129120 -11600
rect 129380 -11620 129620 -11600
rect 129880 -11620 130120 -11600
rect 130380 -11620 130620 -11600
rect 130880 -11620 131120 -11600
rect 131380 -11620 131620 -11600
rect 131880 -11620 132120 -11600
rect 132380 -11620 132620 -11600
rect 132880 -11620 133120 -11600
rect 133380 -11620 133620 -11600
rect 133880 -11620 134120 -11600
rect 134380 -11620 134620 -11600
rect 134880 -11620 135120 -11600
rect 135380 -11620 135620 -11600
rect 135880 -11620 136120 -11600
rect 136380 -11620 136620 -11600
rect 136880 -11620 137120 -11600
rect 137380 -11620 137620 -11600
rect 137880 -11620 138120 -11600
rect 138380 -11620 138620 -11600
rect 138880 -11620 139120 -11600
rect 139380 -11620 139620 -11600
rect 139880 -11620 140000 -11600
rect 112000 -11880 112100 -11620
rect 112400 -11880 112600 -11620
rect 112900 -11880 113100 -11620
rect 113400 -11880 113600 -11620
rect 113900 -11880 114100 -11620
rect 114400 -11880 114600 -11620
rect 114900 -11880 115100 -11620
rect 115400 -11880 115600 -11620
rect 115900 -11880 116100 -11620
rect 116400 -11880 116600 -11620
rect 116900 -11880 117100 -11620
rect 117400 -11880 117600 -11620
rect 117900 -11880 118100 -11620
rect 118400 -11880 118600 -11620
rect 118900 -11880 119100 -11620
rect 119400 -11880 119600 -11620
rect 119900 -11880 120100 -11620
rect 120400 -11880 120600 -11620
rect 120900 -11880 121100 -11620
rect 121400 -11880 121600 -11620
rect 121900 -11880 122100 -11620
rect 122400 -11880 122600 -11620
rect 122900 -11880 123100 -11620
rect 123400 -11880 123600 -11620
rect 123900 -11880 124100 -11620
rect 124400 -11880 124600 -11620
rect 124900 -11880 125100 -11620
rect 125400 -11880 125600 -11620
rect 125900 -11880 126100 -11620
rect 126400 -11880 126600 -11620
rect 126900 -11880 127100 -11620
rect 127400 -11880 127600 -11620
rect 127900 -11880 128100 -11620
rect 128400 -11880 128600 -11620
rect 128900 -11880 129100 -11620
rect 129400 -11880 129600 -11620
rect 129900 -11880 130100 -11620
rect 130400 -11880 130600 -11620
rect 130900 -11880 131100 -11620
rect 131400 -11880 131600 -11620
rect 131900 -11880 132100 -11620
rect 132400 -11880 132600 -11620
rect 132900 -11880 133100 -11620
rect 133400 -11880 133600 -11620
rect 133900 -11880 134100 -11620
rect 134400 -11880 134600 -11620
rect 134900 -11880 135100 -11620
rect 135400 -11880 135600 -11620
rect 135900 -11880 136100 -11620
rect 136400 -11880 136600 -11620
rect 136900 -11880 137100 -11620
rect 137400 -11880 137600 -11620
rect 137900 -11880 138100 -11620
rect 138400 -11880 138600 -11620
rect 138900 -11880 139100 -11620
rect 139400 -11880 139600 -11620
rect 139900 -11880 140000 -11620
rect 112000 -11900 112120 -11880
rect 112380 -11900 112620 -11880
rect 112880 -11900 113120 -11880
rect 113380 -11900 113620 -11880
rect 113880 -11900 114120 -11880
rect 114380 -11900 114620 -11880
rect 114880 -11900 115120 -11880
rect 115380 -11900 115620 -11880
rect 115880 -11900 116120 -11880
rect 116380 -11900 116620 -11880
rect 116880 -11900 117120 -11880
rect 117380 -11900 117620 -11880
rect 117880 -11900 118120 -11880
rect 118380 -11900 118620 -11880
rect 118880 -11900 119120 -11880
rect 119380 -11900 119620 -11880
rect 119880 -11900 120120 -11880
rect 120380 -11900 120620 -11880
rect 120880 -11900 121120 -11880
rect 121380 -11900 121620 -11880
rect 121880 -11900 122120 -11880
rect 122380 -11900 122620 -11880
rect 122880 -11900 123120 -11880
rect 123380 -11900 123620 -11880
rect 123880 -11900 124120 -11880
rect 124380 -11900 124620 -11880
rect 124880 -11900 125120 -11880
rect 125380 -11900 125620 -11880
rect 125880 -11900 126120 -11880
rect 126380 -11900 126620 -11880
rect 126880 -11900 127120 -11880
rect 127380 -11900 127620 -11880
rect 127880 -11900 128120 -11880
rect 128380 -11900 128620 -11880
rect 128880 -11900 129120 -11880
rect 129380 -11900 129620 -11880
rect 129880 -11900 130120 -11880
rect 130380 -11900 130620 -11880
rect 130880 -11900 131120 -11880
rect 131380 -11900 131620 -11880
rect 131880 -11900 132120 -11880
rect 132380 -11900 132620 -11880
rect 132880 -11900 133120 -11880
rect 133380 -11900 133620 -11880
rect 133880 -11900 134120 -11880
rect 134380 -11900 134620 -11880
rect 134880 -11900 135120 -11880
rect 135380 -11900 135620 -11880
rect 135880 -11900 136120 -11880
rect 136380 -11900 136620 -11880
rect 136880 -11900 137120 -11880
rect 137380 -11900 137620 -11880
rect 137880 -11900 138120 -11880
rect 138380 -11900 138620 -11880
rect 138880 -11900 139120 -11880
rect 139380 -11900 139620 -11880
rect 139880 -11900 140000 -11880
rect 112000 -12100 140000 -11900
rect 112000 -12120 112120 -12100
rect 112380 -12120 112620 -12100
rect 112880 -12120 113120 -12100
rect 113380 -12120 113620 -12100
rect 113880 -12120 114120 -12100
rect 114380 -12120 114620 -12100
rect 114880 -12120 115120 -12100
rect 115380 -12120 115620 -12100
rect 115880 -12120 116120 -12100
rect 116380 -12120 116620 -12100
rect 116880 -12120 117120 -12100
rect 117380 -12120 117620 -12100
rect 117880 -12120 118120 -12100
rect 118380 -12120 118620 -12100
rect 118880 -12120 119120 -12100
rect 119380 -12120 119620 -12100
rect 119880 -12120 120120 -12100
rect 120380 -12120 120620 -12100
rect 120880 -12120 121120 -12100
rect 121380 -12120 121620 -12100
rect 121880 -12120 122120 -12100
rect 122380 -12120 122620 -12100
rect 122880 -12120 123120 -12100
rect 123380 -12120 123620 -12100
rect 123880 -12120 124120 -12100
rect 124380 -12120 124620 -12100
rect 124880 -12120 125120 -12100
rect 125380 -12120 125620 -12100
rect 125880 -12120 126120 -12100
rect 126380 -12120 126620 -12100
rect 126880 -12120 127120 -12100
rect 127380 -12120 127620 -12100
rect 127880 -12120 128120 -12100
rect 128380 -12120 128620 -12100
rect 128880 -12120 129120 -12100
rect 129380 -12120 129620 -12100
rect 129880 -12120 130120 -12100
rect 130380 -12120 130620 -12100
rect 130880 -12120 131120 -12100
rect 131380 -12120 131620 -12100
rect 131880 -12120 132120 -12100
rect 132380 -12120 132620 -12100
rect 132880 -12120 133120 -12100
rect 133380 -12120 133620 -12100
rect 133880 -12120 134120 -12100
rect 134380 -12120 134620 -12100
rect 134880 -12120 135120 -12100
rect 135380 -12120 135620 -12100
rect 135880 -12120 136120 -12100
rect 136380 -12120 136620 -12100
rect 136880 -12120 137120 -12100
rect 137380 -12120 137620 -12100
rect 137880 -12120 138120 -12100
rect 138380 -12120 138620 -12100
rect 138880 -12120 139120 -12100
rect 139380 -12120 139620 -12100
rect 139880 -12120 140000 -12100
rect 112000 -12380 112100 -12120
rect 112400 -12380 112600 -12120
rect 112900 -12380 113100 -12120
rect 113400 -12380 113600 -12120
rect 113900 -12380 114100 -12120
rect 114400 -12380 114600 -12120
rect 114900 -12380 115100 -12120
rect 115400 -12380 115600 -12120
rect 115900 -12380 116100 -12120
rect 116400 -12380 116600 -12120
rect 116900 -12380 117100 -12120
rect 117400 -12380 117600 -12120
rect 117900 -12380 118100 -12120
rect 118400 -12380 118600 -12120
rect 118900 -12380 119100 -12120
rect 119400 -12380 119600 -12120
rect 119900 -12380 120100 -12120
rect 120400 -12380 120600 -12120
rect 120900 -12380 121100 -12120
rect 121400 -12380 121600 -12120
rect 121900 -12380 122100 -12120
rect 122400 -12380 122600 -12120
rect 122900 -12380 123100 -12120
rect 123400 -12380 123600 -12120
rect 123900 -12380 124100 -12120
rect 124400 -12380 124600 -12120
rect 124900 -12380 125100 -12120
rect 125400 -12380 125600 -12120
rect 125900 -12380 126100 -12120
rect 126400 -12380 126600 -12120
rect 126900 -12380 127100 -12120
rect 127400 -12380 127600 -12120
rect 127900 -12380 128100 -12120
rect 128400 -12380 128600 -12120
rect 128900 -12380 129100 -12120
rect 129400 -12380 129600 -12120
rect 129900 -12380 130100 -12120
rect 130400 -12380 130600 -12120
rect 130900 -12380 131100 -12120
rect 131400 -12380 131600 -12120
rect 131900 -12380 132100 -12120
rect 132400 -12380 132600 -12120
rect 132900 -12380 133100 -12120
rect 133400 -12380 133600 -12120
rect 133900 -12380 134100 -12120
rect 134400 -12380 134600 -12120
rect 134900 -12380 135100 -12120
rect 135400 -12380 135600 -12120
rect 135900 -12380 136100 -12120
rect 136400 -12380 136600 -12120
rect 136900 -12380 137100 -12120
rect 137400 -12380 137600 -12120
rect 137900 -12380 138100 -12120
rect 138400 -12380 138600 -12120
rect 138900 -12380 139100 -12120
rect 139400 -12380 139600 -12120
rect 139900 -12380 140000 -12120
rect 112000 -12400 112120 -12380
rect 112380 -12400 112620 -12380
rect 112880 -12400 113120 -12380
rect 113380 -12400 113620 -12380
rect 113880 -12400 114120 -12380
rect 114380 -12400 114620 -12380
rect 114880 -12400 115120 -12380
rect 115380 -12400 115620 -12380
rect 115880 -12400 116120 -12380
rect 116380 -12400 116620 -12380
rect 116880 -12400 117120 -12380
rect 117380 -12400 117620 -12380
rect 117880 -12400 118120 -12380
rect 118380 -12400 118620 -12380
rect 118880 -12400 119120 -12380
rect 119380 -12400 119620 -12380
rect 119880 -12400 120120 -12380
rect 120380 -12400 120620 -12380
rect 120880 -12400 121120 -12380
rect 121380 -12400 121620 -12380
rect 121880 -12400 122120 -12380
rect 122380 -12400 122620 -12380
rect 122880 -12400 123120 -12380
rect 123380 -12400 123620 -12380
rect 123880 -12400 124120 -12380
rect 124380 -12400 124620 -12380
rect 124880 -12400 125120 -12380
rect 125380 -12400 125620 -12380
rect 125880 -12400 126120 -12380
rect 126380 -12400 126620 -12380
rect 126880 -12400 127120 -12380
rect 127380 -12400 127620 -12380
rect 127880 -12400 128120 -12380
rect 128380 -12400 128620 -12380
rect 128880 -12400 129120 -12380
rect 129380 -12400 129620 -12380
rect 129880 -12400 130120 -12380
rect 130380 -12400 130620 -12380
rect 130880 -12400 131120 -12380
rect 131380 -12400 131620 -12380
rect 131880 -12400 132120 -12380
rect 132380 -12400 132620 -12380
rect 132880 -12400 133120 -12380
rect 133380 -12400 133620 -12380
rect 133880 -12400 134120 -12380
rect 134380 -12400 134620 -12380
rect 134880 -12400 135120 -12380
rect 135380 -12400 135620 -12380
rect 135880 -12400 136120 -12380
rect 136380 -12400 136620 -12380
rect 136880 -12400 137120 -12380
rect 137380 -12400 137620 -12380
rect 137880 -12400 138120 -12380
rect 138380 -12400 138620 -12380
rect 138880 -12400 139120 -12380
rect 139380 -12400 139620 -12380
rect 139880 -12400 140000 -12380
rect 112000 -12600 140000 -12400
rect 112000 -12620 112120 -12600
rect 112380 -12620 112620 -12600
rect 112880 -12620 113120 -12600
rect 113380 -12620 113620 -12600
rect 113880 -12620 114120 -12600
rect 114380 -12620 114620 -12600
rect 114880 -12620 115120 -12600
rect 115380 -12620 115620 -12600
rect 115880 -12620 116120 -12600
rect 116380 -12620 116620 -12600
rect 116880 -12620 117120 -12600
rect 117380 -12620 117620 -12600
rect 117880 -12620 118120 -12600
rect 118380 -12620 118620 -12600
rect 118880 -12620 119120 -12600
rect 119380 -12620 119620 -12600
rect 119880 -12620 120120 -12600
rect 120380 -12620 120620 -12600
rect 120880 -12620 121120 -12600
rect 121380 -12620 121620 -12600
rect 121880 -12620 122120 -12600
rect 122380 -12620 122620 -12600
rect 122880 -12620 123120 -12600
rect 123380 -12620 123620 -12600
rect 123880 -12620 124120 -12600
rect 124380 -12620 124620 -12600
rect 124880 -12620 125120 -12600
rect 125380 -12620 125620 -12600
rect 125880 -12620 126120 -12600
rect 126380 -12620 126620 -12600
rect 126880 -12620 127120 -12600
rect 127380 -12620 127620 -12600
rect 127880 -12620 128120 -12600
rect 128380 -12620 128620 -12600
rect 128880 -12620 129120 -12600
rect 129380 -12620 129620 -12600
rect 129880 -12620 130120 -12600
rect 130380 -12620 130620 -12600
rect 130880 -12620 131120 -12600
rect 131380 -12620 131620 -12600
rect 131880 -12620 132120 -12600
rect 132380 -12620 132620 -12600
rect 132880 -12620 133120 -12600
rect 133380 -12620 133620 -12600
rect 133880 -12620 134120 -12600
rect 134380 -12620 134620 -12600
rect 134880 -12620 135120 -12600
rect 135380 -12620 135620 -12600
rect 135880 -12620 136120 -12600
rect 136380 -12620 136620 -12600
rect 136880 -12620 137120 -12600
rect 137380 -12620 137620 -12600
rect 137880 -12620 138120 -12600
rect 138380 -12620 138620 -12600
rect 138880 -12620 139120 -12600
rect 139380 -12620 139620 -12600
rect 139880 -12620 140000 -12600
rect 112000 -12880 112100 -12620
rect 112400 -12880 112600 -12620
rect 112900 -12880 113100 -12620
rect 113400 -12880 113600 -12620
rect 113900 -12880 114100 -12620
rect 114400 -12880 114600 -12620
rect 114900 -12880 115100 -12620
rect 115400 -12880 115600 -12620
rect 115900 -12880 116100 -12620
rect 116400 -12880 116600 -12620
rect 116900 -12880 117100 -12620
rect 117400 -12880 117600 -12620
rect 117900 -12880 118100 -12620
rect 118400 -12880 118600 -12620
rect 118900 -12880 119100 -12620
rect 119400 -12880 119600 -12620
rect 119900 -12880 120100 -12620
rect 120400 -12880 120600 -12620
rect 120900 -12880 121100 -12620
rect 121400 -12880 121600 -12620
rect 121900 -12880 122100 -12620
rect 122400 -12880 122600 -12620
rect 122900 -12880 123100 -12620
rect 123400 -12880 123600 -12620
rect 123900 -12880 124100 -12620
rect 124400 -12880 124600 -12620
rect 124900 -12880 125100 -12620
rect 125400 -12880 125600 -12620
rect 125900 -12880 126100 -12620
rect 126400 -12880 126600 -12620
rect 126900 -12880 127100 -12620
rect 127400 -12880 127600 -12620
rect 127900 -12880 128100 -12620
rect 128400 -12880 128600 -12620
rect 128900 -12880 129100 -12620
rect 129400 -12880 129600 -12620
rect 129900 -12880 130100 -12620
rect 130400 -12880 130600 -12620
rect 130900 -12880 131100 -12620
rect 131400 -12880 131600 -12620
rect 131900 -12880 132100 -12620
rect 132400 -12880 132600 -12620
rect 132900 -12880 133100 -12620
rect 133400 -12880 133600 -12620
rect 133900 -12880 134100 -12620
rect 134400 -12880 134600 -12620
rect 134900 -12880 135100 -12620
rect 135400 -12880 135600 -12620
rect 135900 -12880 136100 -12620
rect 136400 -12880 136600 -12620
rect 136900 -12880 137100 -12620
rect 137400 -12880 137600 -12620
rect 137900 -12880 138100 -12620
rect 138400 -12880 138600 -12620
rect 138900 -12880 139100 -12620
rect 139400 -12880 139600 -12620
rect 139900 -12880 140000 -12620
rect 112000 -12900 112120 -12880
rect 112380 -12900 112620 -12880
rect 112880 -12900 113120 -12880
rect 113380 -12900 113620 -12880
rect 113880 -12900 114120 -12880
rect 114380 -12900 114620 -12880
rect 114880 -12900 115120 -12880
rect 115380 -12900 115620 -12880
rect 115880 -12900 116120 -12880
rect 116380 -12900 116620 -12880
rect 116880 -12900 117120 -12880
rect 117380 -12900 117620 -12880
rect 117880 -12900 118120 -12880
rect 118380 -12900 118620 -12880
rect 118880 -12900 119120 -12880
rect 119380 -12900 119620 -12880
rect 119880 -12900 120120 -12880
rect 120380 -12900 120620 -12880
rect 120880 -12900 121120 -12880
rect 121380 -12900 121620 -12880
rect 121880 -12900 122120 -12880
rect 122380 -12900 122620 -12880
rect 122880 -12900 123120 -12880
rect 123380 -12900 123620 -12880
rect 123880 -12900 124120 -12880
rect 124380 -12900 124620 -12880
rect 124880 -12900 125120 -12880
rect 125380 -12900 125620 -12880
rect 125880 -12900 126120 -12880
rect 126380 -12900 126620 -12880
rect 126880 -12900 127120 -12880
rect 127380 -12900 127620 -12880
rect 127880 -12900 128120 -12880
rect 128380 -12900 128620 -12880
rect 128880 -12900 129120 -12880
rect 129380 -12900 129620 -12880
rect 129880 -12900 130120 -12880
rect 130380 -12900 130620 -12880
rect 130880 -12900 131120 -12880
rect 131380 -12900 131620 -12880
rect 131880 -12900 132120 -12880
rect 132380 -12900 132620 -12880
rect 132880 -12900 133120 -12880
rect 133380 -12900 133620 -12880
rect 133880 -12900 134120 -12880
rect 134380 -12900 134620 -12880
rect 134880 -12900 135120 -12880
rect 135380 -12900 135620 -12880
rect 135880 -12900 136120 -12880
rect 136380 -12900 136620 -12880
rect 136880 -12900 137120 -12880
rect 137380 -12900 137620 -12880
rect 137880 -12900 138120 -12880
rect 138380 -12900 138620 -12880
rect 138880 -12900 139120 -12880
rect 139380 -12900 139620 -12880
rect 139880 -12900 140000 -12880
rect 112000 -13100 140000 -12900
rect 112000 -13120 112120 -13100
rect 112380 -13120 112620 -13100
rect 112880 -13120 113120 -13100
rect 113380 -13120 113620 -13100
rect 113880 -13120 114120 -13100
rect 114380 -13120 114620 -13100
rect 114880 -13120 115120 -13100
rect 115380 -13120 115620 -13100
rect 115880 -13120 116120 -13100
rect 116380 -13120 116620 -13100
rect 116880 -13120 117120 -13100
rect 117380 -13120 117620 -13100
rect 117880 -13120 118120 -13100
rect 118380 -13120 118620 -13100
rect 118880 -13120 119120 -13100
rect 119380 -13120 119620 -13100
rect 119880 -13120 120120 -13100
rect 120380 -13120 120620 -13100
rect 120880 -13120 121120 -13100
rect 121380 -13120 121620 -13100
rect 121880 -13120 122120 -13100
rect 122380 -13120 122620 -13100
rect 122880 -13120 123120 -13100
rect 123380 -13120 123620 -13100
rect 123880 -13120 124120 -13100
rect 124380 -13120 124620 -13100
rect 124880 -13120 125120 -13100
rect 125380 -13120 125620 -13100
rect 125880 -13120 126120 -13100
rect 126380 -13120 126620 -13100
rect 126880 -13120 127120 -13100
rect 127380 -13120 127620 -13100
rect 127880 -13120 128120 -13100
rect 128380 -13120 128620 -13100
rect 128880 -13120 129120 -13100
rect 129380 -13120 129620 -13100
rect 129880 -13120 130120 -13100
rect 130380 -13120 130620 -13100
rect 130880 -13120 131120 -13100
rect 131380 -13120 131620 -13100
rect 131880 -13120 132120 -13100
rect 132380 -13120 132620 -13100
rect 132880 -13120 133120 -13100
rect 133380 -13120 133620 -13100
rect 133880 -13120 134120 -13100
rect 134380 -13120 134620 -13100
rect 134880 -13120 135120 -13100
rect 135380 -13120 135620 -13100
rect 135880 -13120 136120 -13100
rect 136380 -13120 136620 -13100
rect 136880 -13120 137120 -13100
rect 137380 -13120 137620 -13100
rect 137880 -13120 138120 -13100
rect 138380 -13120 138620 -13100
rect 138880 -13120 139120 -13100
rect 139380 -13120 139620 -13100
rect 139880 -13120 140000 -13100
rect 112000 -13380 112100 -13120
rect 112400 -13380 112600 -13120
rect 112900 -13380 113100 -13120
rect 113400 -13380 113600 -13120
rect 113900 -13380 114100 -13120
rect 114400 -13380 114600 -13120
rect 114900 -13380 115100 -13120
rect 115400 -13380 115600 -13120
rect 115900 -13380 116100 -13120
rect 116400 -13380 116600 -13120
rect 116900 -13380 117100 -13120
rect 117400 -13380 117600 -13120
rect 117900 -13380 118100 -13120
rect 118400 -13380 118600 -13120
rect 118900 -13380 119100 -13120
rect 119400 -13380 119600 -13120
rect 119900 -13380 120100 -13120
rect 120400 -13380 120600 -13120
rect 120900 -13380 121100 -13120
rect 121400 -13380 121600 -13120
rect 121900 -13380 122100 -13120
rect 122400 -13380 122600 -13120
rect 122900 -13380 123100 -13120
rect 123400 -13380 123600 -13120
rect 123900 -13380 124100 -13120
rect 124400 -13380 124600 -13120
rect 124900 -13380 125100 -13120
rect 125400 -13380 125600 -13120
rect 125900 -13380 126100 -13120
rect 126400 -13380 126600 -13120
rect 126900 -13380 127100 -13120
rect 127400 -13380 127600 -13120
rect 127900 -13380 128100 -13120
rect 128400 -13380 128600 -13120
rect 128900 -13380 129100 -13120
rect 129400 -13380 129600 -13120
rect 129900 -13380 130100 -13120
rect 130400 -13380 130600 -13120
rect 130900 -13380 131100 -13120
rect 131400 -13380 131600 -13120
rect 131900 -13380 132100 -13120
rect 132400 -13380 132600 -13120
rect 132900 -13380 133100 -13120
rect 133400 -13380 133600 -13120
rect 133900 -13380 134100 -13120
rect 134400 -13380 134600 -13120
rect 134900 -13380 135100 -13120
rect 135400 -13380 135600 -13120
rect 135900 -13380 136100 -13120
rect 136400 -13380 136600 -13120
rect 136900 -13380 137100 -13120
rect 137400 -13380 137600 -13120
rect 137900 -13380 138100 -13120
rect 138400 -13380 138600 -13120
rect 138900 -13380 139100 -13120
rect 139400 -13380 139600 -13120
rect 139900 -13380 140000 -13120
rect 112000 -13400 112120 -13380
rect 112380 -13400 112620 -13380
rect 112880 -13400 113120 -13380
rect 113380 -13400 113620 -13380
rect 113880 -13400 114120 -13380
rect 114380 -13400 114620 -13380
rect 114880 -13400 115120 -13380
rect 115380 -13400 115620 -13380
rect 115880 -13400 116120 -13380
rect 116380 -13400 116620 -13380
rect 116880 -13400 117120 -13380
rect 117380 -13400 117620 -13380
rect 117880 -13400 118120 -13380
rect 118380 -13400 118620 -13380
rect 118880 -13400 119120 -13380
rect 119380 -13400 119620 -13380
rect 119880 -13400 120120 -13380
rect 120380 -13400 120620 -13380
rect 120880 -13400 121120 -13380
rect 121380 -13400 121620 -13380
rect 121880 -13400 122120 -13380
rect 122380 -13400 122620 -13380
rect 122880 -13400 123120 -13380
rect 123380 -13400 123620 -13380
rect 123880 -13400 124120 -13380
rect 124380 -13400 124620 -13380
rect 124880 -13400 125120 -13380
rect 125380 -13400 125620 -13380
rect 125880 -13400 126120 -13380
rect 126380 -13400 126620 -13380
rect 126880 -13400 127120 -13380
rect 127380 -13400 127620 -13380
rect 127880 -13400 128120 -13380
rect 128380 -13400 128620 -13380
rect 128880 -13400 129120 -13380
rect 129380 -13400 129620 -13380
rect 129880 -13400 130120 -13380
rect 130380 -13400 130620 -13380
rect 130880 -13400 131120 -13380
rect 131380 -13400 131620 -13380
rect 131880 -13400 132120 -13380
rect 132380 -13400 132620 -13380
rect 132880 -13400 133120 -13380
rect 133380 -13400 133620 -13380
rect 133880 -13400 134120 -13380
rect 134380 -13400 134620 -13380
rect 134880 -13400 135120 -13380
rect 135380 -13400 135620 -13380
rect 135880 -13400 136120 -13380
rect 136380 -13400 136620 -13380
rect 136880 -13400 137120 -13380
rect 137380 -13400 137620 -13380
rect 137880 -13400 138120 -13380
rect 138380 -13400 138620 -13380
rect 138880 -13400 139120 -13380
rect 139380 -13400 139620 -13380
rect 139880 -13400 140000 -13380
rect 112000 -13600 140000 -13400
rect 112000 -13620 112120 -13600
rect 112380 -13620 112620 -13600
rect 112880 -13620 113120 -13600
rect 113380 -13620 113620 -13600
rect 113880 -13620 114120 -13600
rect 114380 -13620 114620 -13600
rect 114880 -13620 115120 -13600
rect 115380 -13620 115620 -13600
rect 115880 -13620 116120 -13600
rect 116380 -13620 116620 -13600
rect 116880 -13620 117120 -13600
rect 117380 -13620 117620 -13600
rect 117880 -13620 118120 -13600
rect 118380 -13620 118620 -13600
rect 118880 -13620 119120 -13600
rect 119380 -13620 119620 -13600
rect 119880 -13620 120120 -13600
rect 120380 -13620 120620 -13600
rect 120880 -13620 121120 -13600
rect 121380 -13620 121620 -13600
rect 121880 -13620 122120 -13600
rect 122380 -13620 122620 -13600
rect 122880 -13620 123120 -13600
rect 123380 -13620 123620 -13600
rect 123880 -13620 124120 -13600
rect 124380 -13620 124620 -13600
rect 124880 -13620 125120 -13600
rect 125380 -13620 125620 -13600
rect 125880 -13620 126120 -13600
rect 126380 -13620 126620 -13600
rect 126880 -13620 127120 -13600
rect 127380 -13620 127620 -13600
rect 127880 -13620 128120 -13600
rect 128380 -13620 128620 -13600
rect 128880 -13620 129120 -13600
rect 129380 -13620 129620 -13600
rect 129880 -13620 130120 -13600
rect 130380 -13620 130620 -13600
rect 130880 -13620 131120 -13600
rect 131380 -13620 131620 -13600
rect 131880 -13620 132120 -13600
rect 132380 -13620 132620 -13600
rect 132880 -13620 133120 -13600
rect 133380 -13620 133620 -13600
rect 133880 -13620 134120 -13600
rect 134380 -13620 134620 -13600
rect 134880 -13620 135120 -13600
rect 135380 -13620 135620 -13600
rect 135880 -13620 136120 -13600
rect 136380 -13620 136620 -13600
rect 136880 -13620 137120 -13600
rect 137380 -13620 137620 -13600
rect 137880 -13620 138120 -13600
rect 138380 -13620 138620 -13600
rect 138880 -13620 139120 -13600
rect 139380 -13620 139620 -13600
rect 139880 -13620 140000 -13600
rect 112000 -13880 112100 -13620
rect 112400 -13880 112600 -13620
rect 112900 -13880 113100 -13620
rect 113400 -13880 113600 -13620
rect 113900 -13880 114100 -13620
rect 114400 -13880 114600 -13620
rect 114900 -13880 115100 -13620
rect 115400 -13880 115600 -13620
rect 115900 -13880 116100 -13620
rect 116400 -13880 116600 -13620
rect 116900 -13880 117100 -13620
rect 117400 -13880 117600 -13620
rect 117900 -13880 118100 -13620
rect 118400 -13880 118600 -13620
rect 118900 -13880 119100 -13620
rect 119400 -13880 119600 -13620
rect 119900 -13880 120100 -13620
rect 120400 -13880 120600 -13620
rect 120900 -13880 121100 -13620
rect 121400 -13880 121600 -13620
rect 121900 -13880 122100 -13620
rect 122400 -13880 122600 -13620
rect 122900 -13880 123100 -13620
rect 123400 -13880 123600 -13620
rect 123900 -13880 124100 -13620
rect 124400 -13880 124600 -13620
rect 124900 -13880 125100 -13620
rect 125400 -13880 125600 -13620
rect 125900 -13880 126100 -13620
rect 126400 -13880 126600 -13620
rect 126900 -13880 127100 -13620
rect 127400 -13880 127600 -13620
rect 127900 -13880 128100 -13620
rect 128400 -13880 128600 -13620
rect 128900 -13880 129100 -13620
rect 129400 -13880 129600 -13620
rect 129900 -13880 130100 -13620
rect 130400 -13880 130600 -13620
rect 130900 -13880 131100 -13620
rect 131400 -13880 131600 -13620
rect 131900 -13880 132100 -13620
rect 132400 -13880 132600 -13620
rect 132900 -13880 133100 -13620
rect 133400 -13880 133600 -13620
rect 133900 -13880 134100 -13620
rect 134400 -13880 134600 -13620
rect 134900 -13880 135100 -13620
rect 135400 -13880 135600 -13620
rect 135900 -13880 136100 -13620
rect 136400 -13880 136600 -13620
rect 136900 -13880 137100 -13620
rect 137400 -13880 137600 -13620
rect 137900 -13880 138100 -13620
rect 138400 -13880 138600 -13620
rect 138900 -13880 139100 -13620
rect 139400 -13880 139600 -13620
rect 139900 -13880 140000 -13620
rect 112000 -13900 112120 -13880
rect 112380 -13900 112620 -13880
rect 112880 -13900 113120 -13880
rect 113380 -13900 113620 -13880
rect 113880 -13900 114120 -13880
rect 114380 -13900 114620 -13880
rect 114880 -13900 115120 -13880
rect 115380 -13900 115620 -13880
rect 115880 -13900 116120 -13880
rect 116380 -13900 116620 -13880
rect 116880 -13900 117120 -13880
rect 117380 -13900 117620 -13880
rect 117880 -13900 118120 -13880
rect 118380 -13900 118620 -13880
rect 118880 -13900 119120 -13880
rect 119380 -13900 119620 -13880
rect 119880 -13900 120120 -13880
rect 120380 -13900 120620 -13880
rect 120880 -13900 121120 -13880
rect 121380 -13900 121620 -13880
rect 121880 -13900 122120 -13880
rect 122380 -13900 122620 -13880
rect 122880 -13900 123120 -13880
rect 123380 -13900 123620 -13880
rect 123880 -13900 124120 -13880
rect 124380 -13900 124620 -13880
rect 124880 -13900 125120 -13880
rect 125380 -13900 125620 -13880
rect 125880 -13900 126120 -13880
rect 126380 -13900 126620 -13880
rect 126880 -13900 127120 -13880
rect 127380 -13900 127620 -13880
rect 127880 -13900 128120 -13880
rect 128380 -13900 128620 -13880
rect 128880 -13900 129120 -13880
rect 129380 -13900 129620 -13880
rect 129880 -13900 130120 -13880
rect 130380 -13900 130620 -13880
rect 130880 -13900 131120 -13880
rect 131380 -13900 131620 -13880
rect 131880 -13900 132120 -13880
rect 132380 -13900 132620 -13880
rect 132880 -13900 133120 -13880
rect 133380 -13900 133620 -13880
rect 133880 -13900 134120 -13880
rect 134380 -13900 134620 -13880
rect 134880 -13900 135120 -13880
rect 135380 -13900 135620 -13880
rect 135880 -13900 136120 -13880
rect 136380 -13900 136620 -13880
rect 136880 -13900 137120 -13880
rect 137380 -13900 137620 -13880
rect 137880 -13900 138120 -13880
rect 138380 -13900 138620 -13880
rect 138880 -13900 139120 -13880
rect 139380 -13900 139620 -13880
rect 139880 -13900 140000 -13880
rect 112000 -14000 140000 -13900
<< via1 >>
rect -15850 97910 -15650 97980
rect -15350 97910 -15150 97980
rect -14850 97910 -14650 97980
rect -14350 97910 -14150 97980
rect -13850 97910 -13650 97980
rect -13350 97910 -13150 97980
rect -12850 97910 -12650 97980
rect -12350 97910 -12150 97980
rect -11850 97910 -11650 97980
rect -11350 97910 -11150 97980
rect -10850 97910 -10650 97980
rect -10350 97910 -10150 97980
rect -9850 97910 -9650 97980
rect -9350 97910 -9150 97980
rect -8850 97910 -8650 97980
rect -8350 97910 -8150 97980
rect -7850 97910 -7650 97980
rect -7350 97910 -7150 97980
rect -6850 97910 -6650 97980
rect -6350 97910 -6150 97980
rect -5850 97910 -5650 97980
rect -5350 97910 -5150 97980
rect -4850 97910 -4650 97980
rect -4350 97910 -4150 97980
rect -3850 97910 -3650 97980
rect -3350 97910 -3150 97980
rect -2850 97910 -2650 97980
rect -2350 97910 -2150 97980
rect -1850 97910 -1650 97980
rect -1350 97910 -1150 97980
rect -850 97910 -650 97980
rect -350 97910 -150 97980
rect 150 97910 350 97980
rect 650 97910 850 97980
rect 1150 97910 1350 97980
rect 1650 97910 1850 97980
rect 2150 97910 2350 97980
rect 2650 97910 2850 97980
rect 3150 97910 3350 97980
rect 3650 97910 3850 97980
rect 4150 97910 4350 97980
rect 4650 97910 4850 97980
rect 5150 97910 5350 97980
rect 5650 97910 5850 97980
rect 6150 97910 6350 97980
rect 6650 97910 6850 97980
rect 7150 97910 7350 97980
rect 7650 97910 7850 97980
rect 8150 97910 8350 97980
rect 8650 97910 8850 97980
rect 9150 97910 9350 97980
rect 9650 97910 9850 97980
rect 10150 97910 10350 97980
rect 10650 97910 10850 97980
rect 11150 97910 11350 97980
rect 11650 97910 11850 97980
rect 12150 97910 12350 97980
rect 12650 97910 12850 97980
rect 13150 97910 13350 97980
rect 13650 97910 13850 97980
rect 14150 97910 14350 97980
rect 14650 97910 14850 97980
rect 15150 97910 15350 97980
rect 15650 97910 15850 97980
rect 16150 97910 16350 97980
rect 16650 97910 16850 97980
rect 17150 97910 17350 97980
rect 17650 97910 17850 97980
rect 18150 97910 18350 97980
rect 18650 97910 18850 97980
rect 19150 97910 19350 97980
rect 19650 97910 19850 97980
rect -15980 97650 -15910 97850
rect -15590 97650 -15520 97850
rect -15480 97650 -15410 97850
rect -15090 97650 -15020 97850
rect -14980 97650 -14910 97850
rect -14590 97650 -14520 97850
rect -14480 97650 -14410 97850
rect -14090 97650 -14020 97850
rect -13980 97650 -13910 97850
rect -13590 97650 -13520 97850
rect -13480 97650 -13410 97850
rect -13090 97650 -13020 97850
rect -12980 97650 -12910 97850
rect -12590 97650 -12520 97850
rect -12480 97650 -12410 97850
rect -12090 97650 -12020 97850
rect -11980 97650 -11910 97850
rect -11590 97650 -11520 97850
rect -11480 97650 -11410 97850
rect -11090 97650 -11020 97850
rect -10980 97650 -10910 97850
rect -10590 97650 -10520 97850
rect -10480 97650 -10410 97850
rect -10090 97650 -10020 97850
rect -9980 97650 -9910 97850
rect -9590 97650 -9520 97850
rect -9480 97650 -9410 97850
rect -9090 97650 -9020 97850
rect -8980 97650 -8910 97850
rect -8590 97650 -8520 97850
rect -8480 97650 -8410 97850
rect -8090 97650 -8020 97850
rect -7980 97650 -7910 97850
rect -7590 97650 -7520 97850
rect -7480 97650 -7410 97850
rect -7090 97650 -7020 97850
rect -6980 97650 -6910 97850
rect -6590 97650 -6520 97850
rect -6480 97650 -6410 97850
rect -6090 97650 -6020 97850
rect -5980 97650 -5910 97850
rect -5590 97650 -5520 97850
rect -5480 97650 -5410 97850
rect -5090 97650 -5020 97850
rect -4980 97650 -4910 97850
rect -4590 97650 -4520 97850
rect -4480 97650 -4410 97850
rect -4090 97650 -4020 97850
rect -3980 97650 -3910 97850
rect -3590 97650 -3520 97850
rect -3480 97650 -3410 97850
rect -3090 97650 -3020 97850
rect -2980 97650 -2910 97850
rect -2590 97650 -2520 97850
rect -2480 97650 -2410 97850
rect -2090 97650 -2020 97850
rect -1980 97650 -1910 97850
rect -1590 97650 -1520 97850
rect -1480 97650 -1410 97850
rect -1090 97650 -1020 97850
rect -980 97650 -910 97850
rect -590 97650 -520 97850
rect -480 97650 -410 97850
rect -90 97650 -20 97850
rect 20 97650 90 97850
rect 410 97650 480 97850
rect 520 97650 590 97850
rect 910 97650 980 97850
rect 1020 97650 1090 97850
rect 1410 97650 1480 97850
rect 1520 97650 1590 97850
rect 1910 97650 1980 97850
rect 2020 97650 2090 97850
rect 2410 97650 2480 97850
rect 2520 97650 2590 97850
rect 2910 97650 2980 97850
rect 3020 97650 3090 97850
rect 3410 97650 3480 97850
rect 3520 97650 3590 97850
rect 3910 97650 3980 97850
rect 4020 97650 4090 97850
rect 4410 97650 4480 97850
rect 4520 97650 4590 97850
rect 4910 97650 4980 97850
rect 5020 97650 5090 97850
rect 5410 97650 5480 97850
rect 5520 97650 5590 97850
rect 5910 97650 5980 97850
rect 6020 97650 6090 97850
rect 6410 97650 6480 97850
rect 6520 97650 6590 97850
rect 6910 97650 6980 97850
rect 7020 97650 7090 97850
rect 7410 97650 7480 97850
rect 7520 97650 7590 97850
rect 7910 97650 7980 97850
rect 8020 97650 8090 97850
rect 8410 97650 8480 97850
rect 8520 97650 8590 97850
rect 8910 97650 8980 97850
rect 9020 97650 9090 97850
rect 9410 97650 9480 97850
rect 9520 97650 9590 97850
rect 9910 97650 9980 97850
rect 10020 97650 10090 97850
rect 10410 97650 10480 97850
rect 10520 97650 10590 97850
rect 10910 97650 10980 97850
rect 11020 97650 11090 97850
rect 11410 97650 11480 97850
rect 11520 97650 11590 97850
rect 11910 97650 11980 97850
rect 12020 97650 12090 97850
rect 12410 97650 12480 97850
rect 12520 97650 12590 97850
rect 12910 97650 12980 97850
rect 13020 97650 13090 97850
rect 13410 97650 13480 97850
rect 13520 97650 13590 97850
rect 13910 97650 13980 97850
rect 14020 97650 14090 97850
rect 14410 97650 14480 97850
rect 14520 97650 14590 97850
rect 14910 97650 14980 97850
rect 15020 97650 15090 97850
rect 15410 97650 15480 97850
rect 15520 97650 15590 97850
rect 15910 97650 15980 97850
rect 16020 97650 16090 97850
rect 16410 97650 16480 97850
rect 16520 97650 16590 97850
rect 16910 97650 16980 97850
rect 17020 97650 17090 97850
rect 17410 97650 17480 97850
rect 17520 97650 17590 97850
rect 17910 97650 17980 97850
rect 18020 97650 18090 97850
rect 18410 97650 18480 97850
rect 18520 97650 18590 97850
rect 18910 97650 18980 97850
rect 19020 97650 19090 97850
rect 19410 97650 19480 97850
rect 19520 97650 19590 97850
rect 19910 97650 19980 97850
rect -15850 97520 -15650 97590
rect -15350 97520 -15150 97590
rect -14850 97520 -14650 97590
rect -14350 97520 -14150 97590
rect -13850 97520 -13650 97590
rect -13350 97520 -13150 97590
rect -12850 97520 -12650 97590
rect -12350 97520 -12150 97590
rect -11850 97520 -11650 97590
rect -11350 97520 -11150 97590
rect -10850 97520 -10650 97590
rect -10350 97520 -10150 97590
rect -9850 97520 -9650 97590
rect -9350 97520 -9150 97590
rect -8850 97520 -8650 97590
rect -8350 97520 -8150 97590
rect -7850 97520 -7650 97590
rect -7350 97520 -7150 97590
rect -6850 97520 -6650 97590
rect -6350 97520 -6150 97590
rect -5850 97520 -5650 97590
rect -5350 97520 -5150 97590
rect -4850 97520 -4650 97590
rect -4350 97520 -4150 97590
rect -3850 97520 -3650 97590
rect -3350 97520 -3150 97590
rect -2850 97520 -2650 97590
rect -2350 97520 -2150 97590
rect -1850 97520 -1650 97590
rect -1350 97520 -1150 97590
rect -850 97520 -650 97590
rect -350 97520 -150 97590
rect 150 97520 350 97590
rect 650 97520 850 97590
rect 1150 97520 1350 97590
rect 1650 97520 1850 97590
rect 2150 97520 2350 97590
rect 2650 97520 2850 97590
rect 3150 97520 3350 97590
rect 3650 97520 3850 97590
rect 4150 97520 4350 97590
rect 4650 97520 4850 97590
rect 5150 97520 5350 97590
rect 5650 97520 5850 97590
rect 6150 97520 6350 97590
rect 6650 97520 6850 97590
rect 7150 97520 7350 97590
rect 7650 97520 7850 97590
rect 8150 97520 8350 97590
rect 8650 97520 8850 97590
rect 9150 97520 9350 97590
rect 9650 97520 9850 97590
rect 10150 97520 10350 97590
rect 10650 97520 10850 97590
rect 11150 97520 11350 97590
rect 11650 97520 11850 97590
rect 12150 97520 12350 97590
rect 12650 97520 12850 97590
rect 13150 97520 13350 97590
rect 13650 97520 13850 97590
rect 14150 97520 14350 97590
rect 14650 97520 14850 97590
rect 15150 97520 15350 97590
rect 15650 97520 15850 97590
rect 16150 97520 16350 97590
rect 16650 97520 16850 97590
rect 17150 97520 17350 97590
rect 17650 97520 17850 97590
rect 18150 97520 18350 97590
rect 18650 97520 18850 97590
rect 19150 97520 19350 97590
rect 19650 97520 19850 97590
rect -15850 97410 -15650 97480
rect -15350 97410 -15150 97480
rect -14850 97410 -14650 97480
rect -14350 97410 -14150 97480
rect -13850 97410 -13650 97480
rect -13350 97410 -13150 97480
rect -12850 97410 -12650 97480
rect -12350 97410 -12150 97480
rect -11850 97410 -11650 97480
rect -11350 97410 -11150 97480
rect -10850 97410 -10650 97480
rect -10350 97410 -10150 97480
rect -9850 97410 -9650 97480
rect -9350 97410 -9150 97480
rect -8850 97410 -8650 97480
rect -8350 97410 -8150 97480
rect -7850 97410 -7650 97480
rect -7350 97410 -7150 97480
rect -6850 97410 -6650 97480
rect -6350 97410 -6150 97480
rect -5850 97410 -5650 97480
rect -5350 97410 -5150 97480
rect -4850 97410 -4650 97480
rect -4350 97410 -4150 97480
rect -3850 97410 -3650 97480
rect -3350 97410 -3150 97480
rect -2850 97410 -2650 97480
rect -2350 97410 -2150 97480
rect -1850 97410 -1650 97480
rect -1350 97410 -1150 97480
rect -850 97410 -650 97480
rect -350 97410 -150 97480
rect 150 97410 350 97480
rect 650 97410 850 97480
rect 1150 97410 1350 97480
rect 1650 97410 1850 97480
rect 2150 97410 2350 97480
rect 2650 97410 2850 97480
rect 3150 97410 3350 97480
rect 3650 97410 3850 97480
rect 4150 97410 4350 97480
rect 4650 97410 4850 97480
rect 5150 97410 5350 97480
rect 5650 97410 5850 97480
rect 6150 97410 6350 97480
rect 6650 97410 6850 97480
rect 7150 97410 7350 97480
rect 7650 97410 7850 97480
rect 8150 97410 8350 97480
rect 8650 97410 8850 97480
rect 9150 97410 9350 97480
rect 9650 97410 9850 97480
rect 10150 97410 10350 97480
rect 10650 97410 10850 97480
rect 11150 97410 11350 97480
rect 11650 97410 11850 97480
rect 12150 97410 12350 97480
rect 12650 97410 12850 97480
rect 13150 97410 13350 97480
rect 13650 97410 13850 97480
rect 14150 97410 14350 97480
rect 14650 97410 14850 97480
rect 15150 97410 15350 97480
rect 15650 97410 15850 97480
rect 16150 97410 16350 97480
rect 16650 97410 16850 97480
rect 17150 97410 17350 97480
rect 17650 97410 17850 97480
rect 18150 97410 18350 97480
rect 18650 97410 18850 97480
rect 19150 97410 19350 97480
rect 19650 97410 19850 97480
rect -15980 97150 -15910 97350
rect -15590 97150 -15520 97350
rect -15480 97150 -15410 97350
rect -15090 97150 -15020 97350
rect -14980 97150 -14910 97350
rect -14590 97150 -14520 97350
rect -14480 97150 -14410 97350
rect -14090 97150 -14020 97350
rect -13980 97150 -13910 97350
rect -13590 97150 -13520 97350
rect -13480 97150 -13410 97350
rect -13090 97150 -13020 97350
rect -12980 97150 -12910 97350
rect -12590 97150 -12520 97350
rect -12480 97150 -12410 97350
rect -12090 97150 -12020 97350
rect -11980 97150 -11910 97350
rect -11590 97150 -11520 97350
rect -11480 97150 -11410 97350
rect -11090 97150 -11020 97350
rect -10980 97150 -10910 97350
rect -10590 97150 -10520 97350
rect -10480 97150 -10410 97350
rect -10090 97150 -10020 97350
rect -9980 97150 -9910 97350
rect -9590 97150 -9520 97350
rect -9480 97150 -9410 97350
rect -9090 97150 -9020 97350
rect -8980 97150 -8910 97350
rect -8590 97150 -8520 97350
rect -8480 97150 -8410 97350
rect -8090 97150 -8020 97350
rect -7980 97150 -7910 97350
rect -7590 97150 -7520 97350
rect -7480 97150 -7410 97350
rect -7090 97150 -7020 97350
rect -6980 97150 -6910 97350
rect -6590 97150 -6520 97350
rect -6480 97150 -6410 97350
rect -6090 97150 -6020 97350
rect -5980 97150 -5910 97350
rect -5590 97150 -5520 97350
rect -5480 97150 -5410 97350
rect -5090 97150 -5020 97350
rect -4980 97150 -4910 97350
rect -4590 97150 -4520 97350
rect -4480 97150 -4410 97350
rect -4090 97150 -4020 97350
rect -3980 97150 -3910 97350
rect -3590 97150 -3520 97350
rect -3480 97150 -3410 97350
rect -3090 97150 -3020 97350
rect -2980 97150 -2910 97350
rect -2590 97150 -2520 97350
rect -2480 97150 -2410 97350
rect -2090 97150 -2020 97350
rect -1980 97150 -1910 97350
rect -1590 97150 -1520 97350
rect -1480 97150 -1410 97350
rect -1090 97150 -1020 97350
rect -980 97150 -910 97350
rect -590 97150 -520 97350
rect -480 97150 -410 97350
rect -90 97150 -20 97350
rect 20 97150 90 97350
rect 410 97150 480 97350
rect 520 97150 590 97350
rect 910 97150 980 97350
rect 1020 97150 1090 97350
rect 1410 97150 1480 97350
rect 1520 97150 1590 97350
rect 1910 97150 1980 97350
rect 2020 97150 2090 97350
rect 2410 97150 2480 97350
rect 2520 97150 2590 97350
rect 2910 97150 2980 97350
rect 3020 97150 3090 97350
rect 3410 97150 3480 97350
rect 3520 97150 3590 97350
rect 3910 97150 3980 97350
rect 4020 97150 4090 97350
rect 4410 97150 4480 97350
rect 4520 97150 4590 97350
rect 4910 97150 4980 97350
rect 5020 97150 5090 97350
rect 5410 97150 5480 97350
rect 5520 97150 5590 97350
rect 5910 97150 5980 97350
rect 6020 97150 6090 97350
rect 6410 97150 6480 97350
rect 6520 97150 6590 97350
rect 6910 97150 6980 97350
rect 7020 97150 7090 97350
rect 7410 97150 7480 97350
rect 7520 97150 7590 97350
rect 7910 97150 7980 97350
rect 8020 97150 8090 97350
rect 8410 97150 8480 97350
rect 8520 97150 8590 97350
rect 8910 97150 8980 97350
rect 9020 97150 9090 97350
rect 9410 97150 9480 97350
rect 9520 97150 9590 97350
rect 9910 97150 9980 97350
rect 10020 97150 10090 97350
rect 10410 97150 10480 97350
rect 10520 97150 10590 97350
rect 10910 97150 10980 97350
rect 11020 97150 11090 97350
rect 11410 97150 11480 97350
rect 11520 97150 11590 97350
rect 11910 97150 11980 97350
rect 12020 97150 12090 97350
rect 12410 97150 12480 97350
rect 12520 97150 12590 97350
rect 12910 97150 12980 97350
rect 13020 97150 13090 97350
rect 13410 97150 13480 97350
rect 13520 97150 13590 97350
rect 13910 97150 13980 97350
rect 14020 97150 14090 97350
rect 14410 97150 14480 97350
rect 14520 97150 14590 97350
rect 14910 97150 14980 97350
rect 15020 97150 15090 97350
rect 15410 97150 15480 97350
rect 15520 97150 15590 97350
rect 15910 97150 15980 97350
rect 16020 97150 16090 97350
rect 16410 97150 16480 97350
rect 16520 97150 16590 97350
rect 16910 97150 16980 97350
rect 17020 97150 17090 97350
rect 17410 97150 17480 97350
rect 17520 97150 17590 97350
rect 17910 97150 17980 97350
rect 18020 97150 18090 97350
rect 18410 97150 18480 97350
rect 18520 97150 18590 97350
rect 18910 97150 18980 97350
rect 19020 97150 19090 97350
rect 19410 97150 19480 97350
rect 19520 97150 19590 97350
rect 19910 97150 19980 97350
rect -15850 97020 -15650 97090
rect -15350 97020 -15150 97090
rect -14850 97020 -14650 97090
rect -14350 97020 -14150 97090
rect -13850 97020 -13650 97090
rect -13350 97020 -13150 97090
rect -12850 97020 -12650 97090
rect -12350 97020 -12150 97090
rect -11850 97020 -11650 97090
rect -11350 97020 -11150 97090
rect -10850 97020 -10650 97090
rect -10350 97020 -10150 97090
rect -9850 97020 -9650 97090
rect -9350 97020 -9150 97090
rect -8850 97020 -8650 97090
rect -8350 97020 -8150 97090
rect -7850 97020 -7650 97090
rect -7350 97020 -7150 97090
rect -6850 97020 -6650 97090
rect -6350 97020 -6150 97090
rect -5850 97020 -5650 97090
rect -5350 97020 -5150 97090
rect -4850 97020 -4650 97090
rect -4350 97020 -4150 97090
rect -3850 97020 -3650 97090
rect -3350 97020 -3150 97090
rect -2850 97020 -2650 97090
rect -2350 97020 -2150 97090
rect -1850 97020 -1650 97090
rect -1350 97020 -1150 97090
rect -850 97020 -650 97090
rect -350 97020 -150 97090
rect 150 97020 350 97090
rect 650 97020 850 97090
rect 1150 97020 1350 97090
rect 1650 97020 1850 97090
rect 2150 97020 2350 97090
rect 2650 97020 2850 97090
rect 3150 97020 3350 97090
rect 3650 97020 3850 97090
rect 4150 97020 4350 97090
rect 4650 97020 4850 97090
rect 5150 97020 5350 97090
rect 5650 97020 5850 97090
rect 6150 97020 6350 97090
rect 6650 97020 6850 97090
rect 7150 97020 7350 97090
rect 7650 97020 7850 97090
rect 8150 97020 8350 97090
rect 8650 97020 8850 97090
rect 9150 97020 9350 97090
rect 9650 97020 9850 97090
rect 10150 97020 10350 97090
rect 10650 97020 10850 97090
rect 11150 97020 11350 97090
rect 11650 97020 11850 97090
rect 12150 97020 12350 97090
rect 12650 97020 12850 97090
rect 13150 97020 13350 97090
rect 13650 97020 13850 97090
rect 14150 97020 14350 97090
rect 14650 97020 14850 97090
rect 15150 97020 15350 97090
rect 15650 97020 15850 97090
rect 16150 97020 16350 97090
rect 16650 97020 16850 97090
rect 17150 97020 17350 97090
rect 17650 97020 17850 97090
rect 18150 97020 18350 97090
rect 18650 97020 18850 97090
rect 19150 97020 19350 97090
rect 19650 97020 19850 97090
rect -15850 96910 -15650 96980
rect -15350 96910 -15150 96980
rect -14850 96910 -14650 96980
rect -14350 96910 -14150 96980
rect -13850 96910 -13650 96980
rect -13350 96910 -13150 96980
rect -12850 96910 -12650 96980
rect -12350 96910 -12150 96980
rect -11850 96910 -11650 96980
rect -11350 96910 -11150 96980
rect -10850 96910 -10650 96980
rect -10350 96910 -10150 96980
rect -9850 96910 -9650 96980
rect -9350 96910 -9150 96980
rect -8850 96910 -8650 96980
rect -8350 96910 -8150 96980
rect -7850 96910 -7650 96980
rect -7350 96910 -7150 96980
rect -6850 96910 -6650 96980
rect -6350 96910 -6150 96980
rect -5850 96910 -5650 96980
rect -5350 96910 -5150 96980
rect -4850 96910 -4650 96980
rect -4350 96910 -4150 96980
rect -3850 96910 -3650 96980
rect -3350 96910 -3150 96980
rect -2850 96910 -2650 96980
rect -2350 96910 -2150 96980
rect -1850 96910 -1650 96980
rect -1350 96910 -1150 96980
rect -850 96910 -650 96980
rect -350 96910 -150 96980
rect 150 96910 350 96980
rect 650 96910 850 96980
rect 1150 96910 1350 96980
rect 1650 96910 1850 96980
rect 2150 96910 2350 96980
rect 2650 96910 2850 96980
rect 3150 96910 3350 96980
rect 3650 96910 3850 96980
rect 4150 96910 4350 96980
rect 4650 96910 4850 96980
rect 5150 96910 5350 96980
rect 5650 96910 5850 96980
rect 6150 96910 6350 96980
rect 6650 96910 6850 96980
rect 7150 96910 7350 96980
rect 7650 96910 7850 96980
rect 8150 96910 8350 96980
rect 8650 96910 8850 96980
rect 9150 96910 9350 96980
rect 9650 96910 9850 96980
rect 10150 96910 10350 96980
rect 10650 96910 10850 96980
rect 11150 96910 11350 96980
rect 11650 96910 11850 96980
rect 12150 96910 12350 96980
rect 12650 96910 12850 96980
rect 13150 96910 13350 96980
rect 13650 96910 13850 96980
rect 14150 96910 14350 96980
rect 14650 96910 14850 96980
rect 15150 96910 15350 96980
rect 15650 96910 15850 96980
rect 16150 96910 16350 96980
rect 16650 96910 16850 96980
rect 17150 96910 17350 96980
rect 17650 96910 17850 96980
rect 18150 96910 18350 96980
rect 18650 96910 18850 96980
rect 19150 96910 19350 96980
rect 19650 96910 19850 96980
rect -15980 96650 -15910 96850
rect -15590 96650 -15520 96850
rect -15480 96650 -15410 96850
rect -15090 96650 -15020 96850
rect -14980 96650 -14910 96850
rect -14590 96650 -14520 96850
rect -14480 96650 -14410 96850
rect -14090 96650 -14020 96850
rect -13980 96650 -13910 96850
rect -13590 96650 -13520 96850
rect -13480 96650 -13410 96850
rect -13090 96650 -13020 96850
rect -12980 96650 -12910 96850
rect -12590 96650 -12520 96850
rect -12480 96650 -12410 96850
rect -12090 96650 -12020 96850
rect -11980 96650 -11910 96850
rect -11590 96650 -11520 96850
rect -11480 96650 -11410 96850
rect -11090 96650 -11020 96850
rect -10980 96650 -10910 96850
rect -10590 96650 -10520 96850
rect -10480 96650 -10410 96850
rect -10090 96650 -10020 96850
rect -9980 96650 -9910 96850
rect -9590 96650 -9520 96850
rect -9480 96650 -9410 96850
rect -9090 96650 -9020 96850
rect -8980 96650 -8910 96850
rect -8590 96650 -8520 96850
rect -8480 96650 -8410 96850
rect -8090 96650 -8020 96850
rect -7980 96650 -7910 96850
rect -7590 96650 -7520 96850
rect -7480 96650 -7410 96850
rect -7090 96650 -7020 96850
rect -6980 96650 -6910 96850
rect -6590 96650 -6520 96850
rect -6480 96650 -6410 96850
rect -6090 96650 -6020 96850
rect -5980 96650 -5910 96850
rect -5590 96650 -5520 96850
rect -5480 96650 -5410 96850
rect -5090 96650 -5020 96850
rect -4980 96650 -4910 96850
rect -4590 96650 -4520 96850
rect -4480 96650 -4410 96850
rect -4090 96650 -4020 96850
rect -3980 96650 -3910 96850
rect -3590 96650 -3520 96850
rect -3480 96650 -3410 96850
rect -3090 96650 -3020 96850
rect -2980 96650 -2910 96850
rect -2590 96650 -2520 96850
rect -2480 96650 -2410 96850
rect -2090 96650 -2020 96850
rect -1980 96650 -1910 96850
rect -1590 96650 -1520 96850
rect -1480 96650 -1410 96850
rect -1090 96650 -1020 96850
rect -980 96650 -910 96850
rect -590 96650 -520 96850
rect -480 96650 -410 96850
rect -90 96650 -20 96850
rect 20 96650 90 96850
rect 410 96650 480 96850
rect 520 96650 590 96850
rect 910 96650 980 96850
rect 1020 96650 1090 96850
rect 1410 96650 1480 96850
rect 1520 96650 1590 96850
rect 1910 96650 1980 96850
rect 2020 96650 2090 96850
rect 2410 96650 2480 96850
rect 2520 96650 2590 96850
rect 2910 96650 2980 96850
rect 3020 96650 3090 96850
rect 3410 96650 3480 96850
rect 3520 96650 3590 96850
rect 3910 96650 3980 96850
rect 4020 96650 4090 96850
rect 4410 96650 4480 96850
rect 4520 96650 4590 96850
rect 4910 96650 4980 96850
rect 5020 96650 5090 96850
rect 5410 96650 5480 96850
rect 5520 96650 5590 96850
rect 5910 96650 5980 96850
rect 6020 96650 6090 96850
rect 6410 96650 6480 96850
rect 6520 96650 6590 96850
rect 6910 96650 6980 96850
rect 7020 96650 7090 96850
rect 7410 96650 7480 96850
rect 7520 96650 7590 96850
rect 7910 96650 7980 96850
rect 8020 96650 8090 96850
rect 8410 96650 8480 96850
rect 8520 96650 8590 96850
rect 8910 96650 8980 96850
rect 9020 96650 9090 96850
rect 9410 96650 9480 96850
rect 9520 96650 9590 96850
rect 9910 96650 9980 96850
rect 10020 96650 10090 96850
rect 10410 96650 10480 96850
rect 10520 96650 10590 96850
rect 10910 96650 10980 96850
rect 11020 96650 11090 96850
rect 11410 96650 11480 96850
rect 11520 96650 11590 96850
rect 11910 96650 11980 96850
rect 12020 96650 12090 96850
rect 12410 96650 12480 96850
rect 12520 96650 12590 96850
rect 12910 96650 12980 96850
rect 13020 96650 13090 96850
rect 13410 96650 13480 96850
rect 13520 96650 13590 96850
rect 13910 96650 13980 96850
rect 14020 96650 14090 96850
rect 14410 96650 14480 96850
rect 14520 96650 14590 96850
rect 14910 96650 14980 96850
rect 15020 96650 15090 96850
rect 15410 96650 15480 96850
rect 15520 96650 15590 96850
rect 15910 96650 15980 96850
rect 16020 96650 16090 96850
rect 16410 96650 16480 96850
rect 16520 96650 16590 96850
rect 16910 96650 16980 96850
rect 17020 96650 17090 96850
rect 17410 96650 17480 96850
rect 17520 96650 17590 96850
rect 17910 96650 17980 96850
rect 18020 96650 18090 96850
rect 18410 96650 18480 96850
rect 18520 96650 18590 96850
rect 18910 96650 18980 96850
rect 19020 96650 19090 96850
rect 19410 96650 19480 96850
rect 19520 96650 19590 96850
rect 19910 96650 19980 96850
rect -15850 96520 -15650 96590
rect -15350 96520 -15150 96590
rect -14850 96520 -14650 96590
rect -14350 96520 -14150 96590
rect -13850 96520 -13650 96590
rect -13350 96520 -13150 96590
rect -12850 96520 -12650 96590
rect -12350 96520 -12150 96590
rect -11850 96520 -11650 96590
rect -11350 96520 -11150 96590
rect -10850 96520 -10650 96590
rect -10350 96520 -10150 96590
rect -9850 96520 -9650 96590
rect -9350 96520 -9150 96590
rect -8850 96520 -8650 96590
rect -8350 96520 -8150 96590
rect -7850 96520 -7650 96590
rect -7350 96520 -7150 96590
rect -6850 96520 -6650 96590
rect -6350 96520 -6150 96590
rect -5850 96520 -5650 96590
rect -5350 96520 -5150 96590
rect -4850 96520 -4650 96590
rect -4350 96520 -4150 96590
rect -3850 96520 -3650 96590
rect -3350 96520 -3150 96590
rect -2850 96520 -2650 96590
rect -2350 96520 -2150 96590
rect -1850 96520 -1650 96590
rect -1350 96520 -1150 96590
rect -850 96520 -650 96590
rect -350 96520 -150 96590
rect 150 96520 350 96590
rect 650 96520 850 96590
rect 1150 96520 1350 96590
rect 1650 96520 1850 96590
rect 2150 96520 2350 96590
rect 2650 96520 2850 96590
rect 3150 96520 3350 96590
rect 3650 96520 3850 96590
rect 4150 96520 4350 96590
rect 4650 96520 4850 96590
rect 5150 96520 5350 96590
rect 5650 96520 5850 96590
rect 6150 96520 6350 96590
rect 6650 96520 6850 96590
rect 7150 96520 7350 96590
rect 7650 96520 7850 96590
rect 8150 96520 8350 96590
rect 8650 96520 8850 96590
rect 9150 96520 9350 96590
rect 9650 96520 9850 96590
rect 10150 96520 10350 96590
rect 10650 96520 10850 96590
rect 11150 96520 11350 96590
rect 11650 96520 11850 96590
rect 12150 96520 12350 96590
rect 12650 96520 12850 96590
rect 13150 96520 13350 96590
rect 13650 96520 13850 96590
rect 14150 96520 14350 96590
rect 14650 96520 14850 96590
rect 15150 96520 15350 96590
rect 15650 96520 15850 96590
rect 16150 96520 16350 96590
rect 16650 96520 16850 96590
rect 17150 96520 17350 96590
rect 17650 96520 17850 96590
rect 18150 96520 18350 96590
rect 18650 96520 18850 96590
rect 19150 96520 19350 96590
rect 19650 96520 19850 96590
rect -15850 96410 -15650 96480
rect -15350 96410 -15150 96480
rect -14850 96410 -14650 96480
rect -14350 96410 -14150 96480
rect -13850 96410 -13650 96480
rect -13350 96410 -13150 96480
rect -12850 96410 -12650 96480
rect -12350 96410 -12150 96480
rect -11850 96410 -11650 96480
rect -11350 96410 -11150 96480
rect -10850 96410 -10650 96480
rect -10350 96410 -10150 96480
rect -9850 96410 -9650 96480
rect -9350 96410 -9150 96480
rect -8850 96410 -8650 96480
rect -8350 96410 -8150 96480
rect -7850 96410 -7650 96480
rect -7350 96410 -7150 96480
rect -6850 96410 -6650 96480
rect -6350 96410 -6150 96480
rect -5850 96410 -5650 96480
rect -5350 96410 -5150 96480
rect -4850 96410 -4650 96480
rect -4350 96410 -4150 96480
rect -3850 96410 -3650 96480
rect -3350 96410 -3150 96480
rect -2850 96410 -2650 96480
rect -2350 96410 -2150 96480
rect -1850 96410 -1650 96480
rect -1350 96410 -1150 96480
rect -850 96410 -650 96480
rect -350 96410 -150 96480
rect 150 96410 350 96480
rect 650 96410 850 96480
rect 1150 96410 1350 96480
rect 1650 96410 1850 96480
rect 2150 96410 2350 96480
rect 2650 96410 2850 96480
rect 3150 96410 3350 96480
rect 3650 96410 3850 96480
rect 4150 96410 4350 96480
rect 4650 96410 4850 96480
rect 5150 96410 5350 96480
rect 5650 96410 5850 96480
rect 6150 96410 6350 96480
rect 6650 96410 6850 96480
rect 7150 96410 7350 96480
rect 7650 96410 7850 96480
rect 8150 96410 8350 96480
rect 8650 96410 8850 96480
rect 9150 96410 9350 96480
rect 9650 96410 9850 96480
rect 10150 96410 10350 96480
rect 10650 96410 10850 96480
rect 11150 96410 11350 96480
rect 11650 96410 11850 96480
rect 12150 96410 12350 96480
rect 12650 96410 12850 96480
rect 13150 96410 13350 96480
rect 13650 96410 13850 96480
rect 14150 96410 14350 96480
rect 14650 96410 14850 96480
rect 15150 96410 15350 96480
rect 15650 96410 15850 96480
rect 16150 96410 16350 96480
rect 16650 96410 16850 96480
rect 17150 96410 17350 96480
rect 17650 96410 17850 96480
rect 18150 96410 18350 96480
rect 18650 96410 18850 96480
rect 19150 96410 19350 96480
rect 19650 96410 19850 96480
rect -15980 96150 -15910 96350
rect -15590 96150 -15520 96350
rect -15480 96150 -15410 96350
rect -15090 96150 -15020 96350
rect -14980 96150 -14910 96350
rect -14590 96150 -14520 96350
rect -14480 96150 -14410 96350
rect -14090 96150 -14020 96350
rect -13980 96150 -13910 96350
rect -13590 96150 -13520 96350
rect -13480 96150 -13410 96350
rect -13090 96150 -13020 96350
rect -12980 96150 -12910 96350
rect -12590 96150 -12520 96350
rect -12480 96150 -12410 96350
rect -12090 96150 -12020 96350
rect -11980 96150 -11910 96350
rect -11590 96150 -11520 96350
rect -11480 96150 -11410 96350
rect -11090 96150 -11020 96350
rect -10980 96150 -10910 96350
rect -10590 96150 -10520 96350
rect -10480 96150 -10410 96350
rect -10090 96150 -10020 96350
rect -9980 96150 -9910 96350
rect -9590 96150 -9520 96350
rect -9480 96150 -9410 96350
rect -9090 96150 -9020 96350
rect -8980 96150 -8910 96350
rect -8590 96150 -8520 96350
rect -8480 96150 -8410 96350
rect -8090 96150 -8020 96350
rect -7980 96150 -7910 96350
rect -7590 96150 -7520 96350
rect -7480 96150 -7410 96350
rect -7090 96150 -7020 96350
rect -6980 96150 -6910 96350
rect -6590 96150 -6520 96350
rect -6480 96150 -6410 96350
rect -6090 96150 -6020 96350
rect -5980 96150 -5910 96350
rect -5590 96150 -5520 96350
rect -5480 96150 -5410 96350
rect -5090 96150 -5020 96350
rect -4980 96150 -4910 96350
rect -4590 96150 -4520 96350
rect -4480 96150 -4410 96350
rect -4090 96150 -4020 96350
rect -3980 96150 -3910 96350
rect -3590 96150 -3520 96350
rect -3480 96150 -3410 96350
rect -3090 96150 -3020 96350
rect -2980 96150 -2910 96350
rect -2590 96150 -2520 96350
rect -2480 96150 -2410 96350
rect -2090 96150 -2020 96350
rect -1980 96150 -1910 96350
rect -1590 96150 -1520 96350
rect -1480 96150 -1410 96350
rect -1090 96150 -1020 96350
rect -980 96150 -910 96350
rect -590 96150 -520 96350
rect -480 96150 -410 96350
rect -90 96150 -20 96350
rect 20 96150 90 96350
rect 410 96150 480 96350
rect 520 96150 590 96350
rect 910 96150 980 96350
rect 1020 96150 1090 96350
rect 1410 96150 1480 96350
rect 1520 96150 1590 96350
rect 1910 96150 1980 96350
rect 2020 96150 2090 96350
rect 2410 96150 2480 96350
rect 2520 96150 2590 96350
rect 2910 96150 2980 96350
rect 3020 96150 3090 96350
rect 3410 96150 3480 96350
rect 3520 96150 3590 96350
rect 3910 96150 3980 96350
rect 4020 96150 4090 96350
rect 4410 96150 4480 96350
rect 4520 96150 4590 96350
rect 4910 96150 4980 96350
rect 5020 96150 5090 96350
rect 5410 96150 5480 96350
rect 5520 96150 5590 96350
rect 5910 96150 5980 96350
rect 6020 96150 6090 96350
rect 6410 96150 6480 96350
rect 6520 96150 6590 96350
rect 6910 96150 6980 96350
rect 7020 96150 7090 96350
rect 7410 96150 7480 96350
rect 7520 96150 7590 96350
rect 7910 96150 7980 96350
rect 8020 96150 8090 96350
rect 8410 96150 8480 96350
rect 8520 96150 8590 96350
rect 8910 96150 8980 96350
rect 9020 96150 9090 96350
rect 9410 96150 9480 96350
rect 9520 96150 9590 96350
rect 9910 96150 9980 96350
rect 10020 96150 10090 96350
rect 10410 96150 10480 96350
rect 10520 96150 10590 96350
rect 10910 96150 10980 96350
rect 11020 96150 11090 96350
rect 11410 96150 11480 96350
rect 11520 96150 11590 96350
rect 11910 96150 11980 96350
rect 12020 96150 12090 96350
rect 12410 96150 12480 96350
rect 12520 96150 12590 96350
rect 12910 96150 12980 96350
rect 13020 96150 13090 96350
rect 13410 96150 13480 96350
rect 13520 96150 13590 96350
rect 13910 96150 13980 96350
rect 14020 96150 14090 96350
rect 14410 96150 14480 96350
rect 14520 96150 14590 96350
rect 14910 96150 14980 96350
rect 15020 96150 15090 96350
rect 15410 96150 15480 96350
rect 15520 96150 15590 96350
rect 15910 96150 15980 96350
rect 16020 96150 16090 96350
rect 16410 96150 16480 96350
rect 16520 96150 16590 96350
rect 16910 96150 16980 96350
rect 17020 96150 17090 96350
rect 17410 96150 17480 96350
rect 17520 96150 17590 96350
rect 17910 96150 17980 96350
rect 18020 96150 18090 96350
rect 18410 96150 18480 96350
rect 18520 96150 18590 96350
rect 18910 96150 18980 96350
rect 19020 96150 19090 96350
rect 19410 96150 19480 96350
rect 19520 96150 19590 96350
rect 19910 96150 19980 96350
rect -15850 96020 -15650 96090
rect -15350 96020 -15150 96090
rect -14850 96020 -14650 96090
rect -14350 96020 -14150 96090
rect -13850 96020 -13650 96090
rect -13350 96020 -13150 96090
rect -12850 96020 -12650 96090
rect -12350 96020 -12150 96090
rect -11850 96020 -11650 96090
rect -11350 96020 -11150 96090
rect -10850 96020 -10650 96090
rect -10350 96020 -10150 96090
rect -9850 96020 -9650 96090
rect -9350 96020 -9150 96090
rect -8850 96020 -8650 96090
rect -8350 96020 -8150 96090
rect -7850 96020 -7650 96090
rect -7350 96020 -7150 96090
rect -6850 96020 -6650 96090
rect -6350 96020 -6150 96090
rect -5850 96020 -5650 96090
rect -5350 96020 -5150 96090
rect -4850 96020 -4650 96090
rect -4350 96020 -4150 96090
rect -3850 96020 -3650 96090
rect -3350 96020 -3150 96090
rect -2850 96020 -2650 96090
rect -2350 96020 -2150 96090
rect -1850 96020 -1650 96090
rect -1350 96020 -1150 96090
rect -850 96020 -650 96090
rect -350 96020 -150 96090
rect 150 96020 350 96090
rect 650 96020 850 96090
rect 1150 96020 1350 96090
rect 1650 96020 1850 96090
rect 2150 96020 2350 96090
rect 2650 96020 2850 96090
rect 3150 96020 3350 96090
rect 3650 96020 3850 96090
rect 4150 96020 4350 96090
rect 4650 96020 4850 96090
rect 5150 96020 5350 96090
rect 5650 96020 5850 96090
rect 6150 96020 6350 96090
rect 6650 96020 6850 96090
rect 7150 96020 7350 96090
rect 7650 96020 7850 96090
rect 8150 96020 8350 96090
rect 8650 96020 8850 96090
rect 9150 96020 9350 96090
rect 9650 96020 9850 96090
rect 10150 96020 10350 96090
rect 10650 96020 10850 96090
rect 11150 96020 11350 96090
rect 11650 96020 11850 96090
rect 12150 96020 12350 96090
rect 12650 96020 12850 96090
rect 13150 96020 13350 96090
rect 13650 96020 13850 96090
rect 14150 96020 14350 96090
rect 14650 96020 14850 96090
rect 15150 96020 15350 96090
rect 15650 96020 15850 96090
rect 16150 96020 16350 96090
rect 16650 96020 16850 96090
rect 17150 96020 17350 96090
rect 17650 96020 17850 96090
rect 18150 96020 18350 96090
rect 18650 96020 18850 96090
rect 19150 96020 19350 96090
rect 19650 96020 19850 96090
rect -15850 95910 -15650 95980
rect -15350 95910 -15150 95980
rect -14850 95910 -14650 95980
rect -14350 95910 -14150 95980
rect -13850 95910 -13650 95980
rect -13350 95910 -13150 95980
rect -12850 95910 -12650 95980
rect -12350 95910 -12150 95980
rect -11850 95910 -11650 95980
rect -11350 95910 -11150 95980
rect -10850 95910 -10650 95980
rect -10350 95910 -10150 95980
rect -9850 95910 -9650 95980
rect -9350 95910 -9150 95980
rect -8850 95910 -8650 95980
rect -8350 95910 -8150 95980
rect -7850 95910 -7650 95980
rect -7350 95910 -7150 95980
rect -6850 95910 -6650 95980
rect -6350 95910 -6150 95980
rect -5850 95910 -5650 95980
rect -5350 95910 -5150 95980
rect -4850 95910 -4650 95980
rect -4350 95910 -4150 95980
rect -3850 95910 -3650 95980
rect -3350 95910 -3150 95980
rect -2850 95910 -2650 95980
rect -2350 95910 -2150 95980
rect -1850 95910 -1650 95980
rect -1350 95910 -1150 95980
rect -850 95910 -650 95980
rect -350 95910 -150 95980
rect 150 95910 350 95980
rect 650 95910 850 95980
rect 1150 95910 1350 95980
rect 1650 95910 1850 95980
rect 2150 95910 2350 95980
rect 2650 95910 2850 95980
rect 3150 95910 3350 95980
rect 3650 95910 3850 95980
rect 4150 95910 4350 95980
rect 4650 95910 4850 95980
rect 5150 95910 5350 95980
rect 5650 95910 5850 95980
rect 6150 95910 6350 95980
rect 6650 95910 6850 95980
rect 7150 95910 7350 95980
rect 7650 95910 7850 95980
rect 8150 95910 8350 95980
rect 8650 95910 8850 95980
rect 9150 95910 9350 95980
rect 9650 95910 9850 95980
rect 10150 95910 10350 95980
rect 10650 95910 10850 95980
rect 11150 95910 11350 95980
rect 11650 95910 11850 95980
rect 12150 95910 12350 95980
rect 12650 95910 12850 95980
rect 13150 95910 13350 95980
rect 13650 95910 13850 95980
rect 14150 95910 14350 95980
rect 14650 95910 14850 95980
rect 15150 95910 15350 95980
rect 15650 95910 15850 95980
rect 16150 95910 16350 95980
rect 16650 95910 16850 95980
rect 17150 95910 17350 95980
rect 17650 95910 17850 95980
rect 18150 95910 18350 95980
rect 18650 95910 18850 95980
rect 19150 95910 19350 95980
rect 19650 95910 19850 95980
rect -15980 95650 -15910 95850
rect -15590 95650 -15520 95850
rect -15480 95650 -15410 95850
rect -15090 95650 -15020 95850
rect -14980 95650 -14910 95850
rect -14590 95650 -14520 95850
rect -14480 95650 -14410 95850
rect -14090 95650 -14020 95850
rect -13980 95650 -13910 95850
rect -13590 95650 -13520 95850
rect -13480 95650 -13410 95850
rect -13090 95650 -13020 95850
rect -12980 95650 -12910 95850
rect -12590 95650 -12520 95850
rect -12480 95650 -12410 95850
rect -12090 95650 -12020 95850
rect -11980 95650 -11910 95850
rect -11590 95650 -11520 95850
rect -11480 95650 -11410 95850
rect -11090 95650 -11020 95850
rect -10980 95650 -10910 95850
rect -10590 95650 -10520 95850
rect -10480 95650 -10410 95850
rect -10090 95650 -10020 95850
rect -9980 95650 -9910 95850
rect -9590 95650 -9520 95850
rect -9480 95650 -9410 95850
rect -9090 95650 -9020 95850
rect -8980 95650 -8910 95850
rect -8590 95650 -8520 95850
rect -8480 95650 -8410 95850
rect -8090 95650 -8020 95850
rect -7980 95650 -7910 95850
rect -7590 95650 -7520 95850
rect -7480 95650 -7410 95850
rect -7090 95650 -7020 95850
rect -6980 95650 -6910 95850
rect -6590 95650 -6520 95850
rect -6480 95650 -6410 95850
rect -6090 95650 -6020 95850
rect -5980 95650 -5910 95850
rect -5590 95650 -5520 95850
rect -5480 95650 -5410 95850
rect -5090 95650 -5020 95850
rect -4980 95650 -4910 95850
rect -4590 95650 -4520 95850
rect -4480 95650 -4410 95850
rect -4090 95650 -4020 95850
rect -3980 95650 -3910 95850
rect -3590 95650 -3520 95850
rect -3480 95650 -3410 95850
rect -3090 95650 -3020 95850
rect -2980 95650 -2910 95850
rect -2590 95650 -2520 95850
rect -2480 95650 -2410 95850
rect -2090 95650 -2020 95850
rect -1980 95650 -1910 95850
rect -1590 95650 -1520 95850
rect -1480 95650 -1410 95850
rect -1090 95650 -1020 95850
rect -980 95650 -910 95850
rect -590 95650 -520 95850
rect -480 95650 -410 95850
rect -90 95650 -20 95850
rect 20 95650 90 95850
rect 410 95650 480 95850
rect 520 95650 590 95850
rect 910 95650 980 95850
rect 1020 95650 1090 95850
rect 1410 95650 1480 95850
rect 1520 95650 1590 95850
rect 1910 95650 1980 95850
rect 2020 95650 2090 95850
rect 2410 95650 2480 95850
rect 2520 95650 2590 95850
rect 2910 95650 2980 95850
rect 3020 95650 3090 95850
rect 3410 95650 3480 95850
rect 3520 95650 3590 95850
rect 3910 95650 3980 95850
rect 4020 95650 4090 95850
rect 4410 95650 4480 95850
rect 4520 95650 4590 95850
rect 4910 95650 4980 95850
rect 5020 95650 5090 95850
rect 5410 95650 5480 95850
rect 5520 95650 5590 95850
rect 5910 95650 5980 95850
rect 6020 95650 6090 95850
rect 6410 95650 6480 95850
rect 6520 95650 6590 95850
rect 6910 95650 6980 95850
rect 7020 95650 7090 95850
rect 7410 95650 7480 95850
rect 7520 95650 7590 95850
rect 7910 95650 7980 95850
rect 8020 95650 8090 95850
rect 8410 95650 8480 95850
rect 8520 95650 8590 95850
rect 8910 95650 8980 95850
rect 9020 95650 9090 95850
rect 9410 95650 9480 95850
rect 9520 95650 9590 95850
rect 9910 95650 9980 95850
rect 10020 95650 10090 95850
rect 10410 95650 10480 95850
rect 10520 95650 10590 95850
rect 10910 95650 10980 95850
rect 11020 95650 11090 95850
rect 11410 95650 11480 95850
rect 11520 95650 11590 95850
rect 11910 95650 11980 95850
rect 12020 95650 12090 95850
rect 12410 95650 12480 95850
rect 12520 95650 12590 95850
rect 12910 95650 12980 95850
rect 13020 95650 13090 95850
rect 13410 95650 13480 95850
rect 13520 95650 13590 95850
rect 13910 95650 13980 95850
rect 14020 95650 14090 95850
rect 14410 95650 14480 95850
rect 14520 95650 14590 95850
rect 14910 95650 14980 95850
rect 15020 95650 15090 95850
rect 15410 95650 15480 95850
rect 15520 95650 15590 95850
rect 15910 95650 15980 95850
rect 16020 95650 16090 95850
rect 16410 95650 16480 95850
rect 16520 95650 16590 95850
rect 16910 95650 16980 95850
rect 17020 95650 17090 95850
rect 17410 95650 17480 95850
rect 17520 95650 17590 95850
rect 17910 95650 17980 95850
rect 18020 95650 18090 95850
rect 18410 95650 18480 95850
rect 18520 95650 18590 95850
rect 18910 95650 18980 95850
rect 19020 95650 19090 95850
rect 19410 95650 19480 95850
rect 19520 95650 19590 95850
rect 19910 95650 19980 95850
rect -15850 95520 -15650 95590
rect -15350 95520 -15150 95590
rect -14850 95520 -14650 95590
rect -14350 95520 -14150 95590
rect -13850 95520 -13650 95590
rect -13350 95520 -13150 95590
rect -12850 95520 -12650 95590
rect -12350 95520 -12150 95590
rect -11850 95520 -11650 95590
rect -11350 95520 -11150 95590
rect -10850 95520 -10650 95590
rect -10350 95520 -10150 95590
rect -9850 95520 -9650 95590
rect -9350 95520 -9150 95590
rect -8850 95520 -8650 95590
rect -8350 95520 -8150 95590
rect -7850 95520 -7650 95590
rect -7350 95520 -7150 95590
rect -6850 95520 -6650 95590
rect -6350 95520 -6150 95590
rect -5850 95520 -5650 95590
rect -5350 95520 -5150 95590
rect -4850 95520 -4650 95590
rect -4350 95520 -4150 95590
rect -3850 95520 -3650 95590
rect -3350 95520 -3150 95590
rect -2850 95520 -2650 95590
rect -2350 95520 -2150 95590
rect -1850 95520 -1650 95590
rect -1350 95520 -1150 95590
rect -850 95520 -650 95590
rect -350 95520 -150 95590
rect 150 95520 350 95590
rect 650 95520 850 95590
rect 1150 95520 1350 95590
rect 1650 95520 1850 95590
rect 2150 95520 2350 95590
rect 2650 95520 2850 95590
rect 3150 95520 3350 95590
rect 3650 95520 3850 95590
rect 4150 95520 4350 95590
rect 4650 95520 4850 95590
rect 5150 95520 5350 95590
rect 5650 95520 5850 95590
rect 6150 95520 6350 95590
rect 6650 95520 6850 95590
rect 7150 95520 7350 95590
rect 7650 95520 7850 95590
rect 8150 95520 8350 95590
rect 8650 95520 8850 95590
rect 9150 95520 9350 95590
rect 9650 95520 9850 95590
rect 10150 95520 10350 95590
rect 10650 95520 10850 95590
rect 11150 95520 11350 95590
rect 11650 95520 11850 95590
rect 12150 95520 12350 95590
rect 12650 95520 12850 95590
rect 13150 95520 13350 95590
rect 13650 95520 13850 95590
rect 14150 95520 14350 95590
rect 14650 95520 14850 95590
rect 15150 95520 15350 95590
rect 15650 95520 15850 95590
rect 16150 95520 16350 95590
rect 16650 95520 16850 95590
rect 17150 95520 17350 95590
rect 17650 95520 17850 95590
rect 18150 95520 18350 95590
rect 18650 95520 18850 95590
rect 19150 95520 19350 95590
rect 19650 95520 19850 95590
rect -15850 95410 -15650 95480
rect -15350 95410 -15150 95480
rect -14850 95410 -14650 95480
rect -14350 95410 -14150 95480
rect -13850 95410 -13650 95480
rect -13350 95410 -13150 95480
rect -12850 95410 -12650 95480
rect -12350 95410 -12150 95480
rect -11850 95410 -11650 95480
rect -11350 95410 -11150 95480
rect -10850 95410 -10650 95480
rect -10350 95410 -10150 95480
rect -9850 95410 -9650 95480
rect -9350 95410 -9150 95480
rect -8850 95410 -8650 95480
rect -8350 95410 -8150 95480
rect -7850 95410 -7650 95480
rect -7350 95410 -7150 95480
rect -6850 95410 -6650 95480
rect -6350 95410 -6150 95480
rect -5850 95410 -5650 95480
rect -5350 95410 -5150 95480
rect -4850 95410 -4650 95480
rect -4350 95410 -4150 95480
rect -3850 95410 -3650 95480
rect -3350 95410 -3150 95480
rect -2850 95410 -2650 95480
rect -2350 95410 -2150 95480
rect -1850 95410 -1650 95480
rect -1350 95410 -1150 95480
rect -850 95410 -650 95480
rect -350 95410 -150 95480
rect 150 95410 350 95480
rect 650 95410 850 95480
rect 1150 95410 1350 95480
rect 1650 95410 1850 95480
rect 2150 95410 2350 95480
rect 2650 95410 2850 95480
rect 3150 95410 3350 95480
rect 3650 95410 3850 95480
rect 4150 95410 4350 95480
rect 4650 95410 4850 95480
rect 5150 95410 5350 95480
rect 5650 95410 5850 95480
rect 6150 95410 6350 95480
rect 6650 95410 6850 95480
rect 7150 95410 7350 95480
rect 7650 95410 7850 95480
rect 8150 95410 8350 95480
rect 8650 95410 8850 95480
rect 9150 95410 9350 95480
rect 9650 95410 9850 95480
rect 10150 95410 10350 95480
rect 10650 95410 10850 95480
rect 11150 95410 11350 95480
rect 11650 95410 11850 95480
rect 12150 95410 12350 95480
rect 12650 95410 12850 95480
rect 13150 95410 13350 95480
rect 13650 95410 13850 95480
rect 14150 95410 14350 95480
rect 14650 95410 14850 95480
rect 15150 95410 15350 95480
rect 15650 95410 15850 95480
rect 16150 95410 16350 95480
rect 16650 95410 16850 95480
rect 17150 95410 17350 95480
rect 17650 95410 17850 95480
rect 18150 95410 18350 95480
rect 18650 95410 18850 95480
rect 19150 95410 19350 95480
rect 19650 95410 19850 95480
rect -15980 95150 -15910 95350
rect -15590 95150 -15520 95350
rect -15480 95150 -15410 95350
rect -15090 95150 -15020 95350
rect -14980 95150 -14910 95350
rect -14590 95150 -14520 95350
rect -14480 95150 -14410 95350
rect -14090 95150 -14020 95350
rect -13980 95150 -13910 95350
rect -13590 95150 -13520 95350
rect -13480 95150 -13410 95350
rect -13090 95150 -13020 95350
rect -12980 95150 -12910 95350
rect -12590 95150 -12520 95350
rect -12480 95150 -12410 95350
rect -12090 95150 -12020 95350
rect -11980 95150 -11910 95350
rect -11590 95150 -11520 95350
rect -11480 95150 -11410 95350
rect -11090 95150 -11020 95350
rect -10980 95150 -10910 95350
rect -10590 95150 -10520 95350
rect -10480 95150 -10410 95350
rect -10090 95150 -10020 95350
rect -9980 95150 -9910 95350
rect -9590 95150 -9520 95350
rect -9480 95150 -9410 95350
rect -9090 95150 -9020 95350
rect -8980 95150 -8910 95350
rect -8590 95150 -8520 95350
rect -8480 95150 -8410 95350
rect -8090 95150 -8020 95350
rect -7980 95150 -7910 95350
rect -7590 95150 -7520 95350
rect -7480 95150 -7410 95350
rect -7090 95150 -7020 95350
rect -6980 95150 -6910 95350
rect -6590 95150 -6520 95350
rect -6480 95150 -6410 95350
rect -6090 95150 -6020 95350
rect -5980 95150 -5910 95350
rect -5590 95150 -5520 95350
rect -5480 95150 -5410 95350
rect -5090 95150 -5020 95350
rect -4980 95150 -4910 95350
rect -4590 95150 -4520 95350
rect -4480 95150 -4410 95350
rect -4090 95150 -4020 95350
rect -3980 95150 -3910 95350
rect -3590 95150 -3520 95350
rect -3480 95150 -3410 95350
rect -3090 95150 -3020 95350
rect -2980 95150 -2910 95350
rect -2590 95150 -2520 95350
rect -2480 95150 -2410 95350
rect -2090 95150 -2020 95350
rect -1980 95150 -1910 95350
rect -1590 95150 -1520 95350
rect -1480 95150 -1410 95350
rect -1090 95150 -1020 95350
rect -980 95150 -910 95350
rect -590 95150 -520 95350
rect -480 95150 -410 95350
rect -90 95150 -20 95350
rect 20 95150 90 95350
rect 410 95150 480 95350
rect 520 95150 590 95350
rect 910 95150 980 95350
rect 1020 95150 1090 95350
rect 1410 95150 1480 95350
rect 1520 95150 1590 95350
rect 1910 95150 1980 95350
rect 2020 95150 2090 95350
rect 2410 95150 2480 95350
rect 2520 95150 2590 95350
rect 2910 95150 2980 95350
rect 3020 95150 3090 95350
rect 3410 95150 3480 95350
rect 3520 95150 3590 95350
rect 3910 95150 3980 95350
rect 4020 95150 4090 95350
rect 4410 95150 4480 95350
rect 4520 95150 4590 95350
rect 4910 95150 4980 95350
rect 5020 95150 5090 95350
rect 5410 95150 5480 95350
rect 5520 95150 5590 95350
rect 5910 95150 5980 95350
rect 6020 95150 6090 95350
rect 6410 95150 6480 95350
rect 6520 95150 6590 95350
rect 6910 95150 6980 95350
rect 7020 95150 7090 95350
rect 7410 95150 7480 95350
rect 7520 95150 7590 95350
rect 7910 95150 7980 95350
rect 8020 95150 8090 95350
rect 8410 95150 8480 95350
rect 8520 95150 8590 95350
rect 8910 95150 8980 95350
rect 9020 95150 9090 95350
rect 9410 95150 9480 95350
rect 9520 95150 9590 95350
rect 9910 95150 9980 95350
rect 10020 95150 10090 95350
rect 10410 95150 10480 95350
rect 10520 95150 10590 95350
rect 10910 95150 10980 95350
rect 11020 95150 11090 95350
rect 11410 95150 11480 95350
rect 11520 95150 11590 95350
rect 11910 95150 11980 95350
rect 12020 95150 12090 95350
rect 12410 95150 12480 95350
rect 12520 95150 12590 95350
rect 12910 95150 12980 95350
rect 13020 95150 13090 95350
rect 13410 95150 13480 95350
rect 13520 95150 13590 95350
rect 13910 95150 13980 95350
rect 14020 95150 14090 95350
rect 14410 95150 14480 95350
rect 14520 95150 14590 95350
rect 14910 95150 14980 95350
rect 15020 95150 15090 95350
rect 15410 95150 15480 95350
rect 15520 95150 15590 95350
rect 15910 95150 15980 95350
rect 16020 95150 16090 95350
rect 16410 95150 16480 95350
rect 16520 95150 16590 95350
rect 16910 95150 16980 95350
rect 17020 95150 17090 95350
rect 17410 95150 17480 95350
rect 17520 95150 17590 95350
rect 17910 95150 17980 95350
rect 18020 95150 18090 95350
rect 18410 95150 18480 95350
rect 18520 95150 18590 95350
rect 18910 95150 18980 95350
rect 19020 95150 19090 95350
rect 19410 95150 19480 95350
rect 19520 95150 19590 95350
rect 19910 95150 19980 95350
rect -15850 95020 -15650 95090
rect -15350 95020 -15150 95090
rect -14850 95020 -14650 95090
rect -14350 95020 -14150 95090
rect -13850 95020 -13650 95090
rect -13350 95020 -13150 95090
rect -12850 95020 -12650 95090
rect -12350 95020 -12150 95090
rect -11850 95020 -11650 95090
rect -11350 95020 -11150 95090
rect -10850 95020 -10650 95090
rect -10350 95020 -10150 95090
rect -9850 95020 -9650 95090
rect -9350 95020 -9150 95090
rect -8850 95020 -8650 95090
rect -8350 95020 -8150 95090
rect -7850 95020 -7650 95090
rect -7350 95020 -7150 95090
rect -6850 95020 -6650 95090
rect -6350 95020 -6150 95090
rect -5850 95020 -5650 95090
rect -5350 95020 -5150 95090
rect -4850 95020 -4650 95090
rect -4350 95020 -4150 95090
rect -3850 95020 -3650 95090
rect -3350 95020 -3150 95090
rect -2850 95020 -2650 95090
rect -2350 95020 -2150 95090
rect -1850 95020 -1650 95090
rect -1350 95020 -1150 95090
rect -850 95020 -650 95090
rect -350 95020 -150 95090
rect 150 95020 350 95090
rect 650 95020 850 95090
rect 1150 95020 1350 95090
rect 1650 95020 1850 95090
rect 2150 95020 2350 95090
rect 2650 95020 2850 95090
rect 3150 95020 3350 95090
rect 3650 95020 3850 95090
rect 4150 95020 4350 95090
rect 4650 95020 4850 95090
rect 5150 95020 5350 95090
rect 5650 95020 5850 95090
rect 6150 95020 6350 95090
rect 6650 95020 6850 95090
rect 7150 95020 7350 95090
rect 7650 95020 7850 95090
rect 8150 95020 8350 95090
rect 8650 95020 8850 95090
rect 9150 95020 9350 95090
rect 9650 95020 9850 95090
rect 10150 95020 10350 95090
rect 10650 95020 10850 95090
rect 11150 95020 11350 95090
rect 11650 95020 11850 95090
rect 12150 95020 12350 95090
rect 12650 95020 12850 95090
rect 13150 95020 13350 95090
rect 13650 95020 13850 95090
rect 14150 95020 14350 95090
rect 14650 95020 14850 95090
rect 15150 95020 15350 95090
rect 15650 95020 15850 95090
rect 16150 95020 16350 95090
rect 16650 95020 16850 95090
rect 17150 95020 17350 95090
rect 17650 95020 17850 95090
rect 18150 95020 18350 95090
rect 18650 95020 18850 95090
rect 19150 95020 19350 95090
rect 19650 95020 19850 95090
rect -15850 94910 -15650 94980
rect -15350 94910 -15150 94980
rect -14850 94910 -14650 94980
rect -14350 94910 -14150 94980
rect -13850 94910 -13650 94980
rect -13350 94910 -13150 94980
rect -12850 94910 -12650 94980
rect -12350 94910 -12150 94980
rect -11850 94910 -11650 94980
rect -11350 94910 -11150 94980
rect -10850 94910 -10650 94980
rect -10350 94910 -10150 94980
rect -9850 94910 -9650 94980
rect -9350 94910 -9150 94980
rect -8850 94910 -8650 94980
rect -8350 94910 -8150 94980
rect -7850 94910 -7650 94980
rect -7350 94910 -7150 94980
rect -6850 94910 -6650 94980
rect -6350 94910 -6150 94980
rect -5850 94910 -5650 94980
rect -5350 94910 -5150 94980
rect -4850 94910 -4650 94980
rect -4350 94910 -4150 94980
rect -3850 94910 -3650 94980
rect -3350 94910 -3150 94980
rect -2850 94910 -2650 94980
rect -2350 94910 -2150 94980
rect -1850 94910 -1650 94980
rect -1350 94910 -1150 94980
rect -850 94910 -650 94980
rect -350 94910 -150 94980
rect 150 94910 350 94980
rect 650 94910 850 94980
rect 1150 94910 1350 94980
rect 1650 94910 1850 94980
rect 2150 94910 2350 94980
rect 2650 94910 2850 94980
rect 3150 94910 3350 94980
rect 3650 94910 3850 94980
rect 4150 94910 4350 94980
rect 4650 94910 4850 94980
rect 5150 94910 5350 94980
rect 5650 94910 5850 94980
rect 6150 94910 6350 94980
rect 6650 94910 6850 94980
rect 7150 94910 7350 94980
rect 7650 94910 7850 94980
rect 8150 94910 8350 94980
rect 8650 94910 8850 94980
rect 9150 94910 9350 94980
rect 9650 94910 9850 94980
rect 10150 94910 10350 94980
rect 10650 94910 10850 94980
rect 11150 94910 11350 94980
rect 11650 94910 11850 94980
rect 12150 94910 12350 94980
rect 12650 94910 12850 94980
rect 13150 94910 13350 94980
rect 13650 94910 13850 94980
rect 14150 94910 14350 94980
rect 14650 94910 14850 94980
rect 15150 94910 15350 94980
rect 15650 94910 15850 94980
rect 16150 94910 16350 94980
rect 16650 94910 16850 94980
rect 17150 94910 17350 94980
rect 17650 94910 17850 94980
rect 18150 94910 18350 94980
rect 18650 94910 18850 94980
rect 19150 94910 19350 94980
rect 19650 94910 19850 94980
rect -15980 94650 -15910 94850
rect -15590 94650 -15520 94850
rect -15480 94650 -15410 94850
rect -15090 94650 -15020 94850
rect -14980 94650 -14910 94850
rect -14590 94650 -14520 94850
rect -14480 94650 -14410 94850
rect -14090 94650 -14020 94850
rect -13980 94650 -13910 94850
rect -13590 94650 -13520 94850
rect -13480 94650 -13410 94850
rect -13090 94650 -13020 94850
rect -12980 94650 -12910 94850
rect -12590 94650 -12520 94850
rect -12480 94650 -12410 94850
rect -12090 94650 -12020 94850
rect -11980 94650 -11910 94850
rect -11590 94650 -11520 94850
rect -11480 94650 -11410 94850
rect -11090 94650 -11020 94850
rect -10980 94650 -10910 94850
rect -10590 94650 -10520 94850
rect -10480 94650 -10410 94850
rect -10090 94650 -10020 94850
rect -9980 94650 -9910 94850
rect -9590 94650 -9520 94850
rect -9480 94650 -9410 94850
rect -9090 94650 -9020 94850
rect -8980 94650 -8910 94850
rect -8590 94650 -8520 94850
rect -8480 94650 -8410 94850
rect -8090 94650 -8020 94850
rect -7980 94650 -7910 94850
rect -7590 94650 -7520 94850
rect -7480 94650 -7410 94850
rect -7090 94650 -7020 94850
rect -6980 94650 -6910 94850
rect -6590 94650 -6520 94850
rect -6480 94650 -6410 94850
rect -6090 94650 -6020 94850
rect -5980 94650 -5910 94850
rect -5590 94650 -5520 94850
rect -5480 94650 -5410 94850
rect -5090 94650 -5020 94850
rect -4980 94650 -4910 94850
rect -4590 94650 -4520 94850
rect -4480 94650 -4410 94850
rect -4090 94650 -4020 94850
rect -3980 94650 -3910 94850
rect -3590 94650 -3520 94850
rect -3480 94650 -3410 94850
rect -3090 94650 -3020 94850
rect -2980 94650 -2910 94850
rect -2590 94650 -2520 94850
rect -2480 94650 -2410 94850
rect -2090 94650 -2020 94850
rect -1980 94650 -1910 94850
rect -1590 94650 -1520 94850
rect -1480 94650 -1410 94850
rect -1090 94650 -1020 94850
rect -980 94650 -910 94850
rect -590 94650 -520 94850
rect -480 94650 -410 94850
rect -90 94650 -20 94850
rect 20 94650 90 94850
rect 410 94650 480 94850
rect 520 94650 590 94850
rect 910 94650 980 94850
rect 1020 94650 1090 94850
rect 1410 94650 1480 94850
rect 1520 94650 1590 94850
rect 1910 94650 1980 94850
rect 2020 94650 2090 94850
rect 2410 94650 2480 94850
rect 2520 94650 2590 94850
rect 2910 94650 2980 94850
rect 3020 94650 3090 94850
rect 3410 94650 3480 94850
rect 3520 94650 3590 94850
rect 3910 94650 3980 94850
rect 4020 94650 4090 94850
rect 4410 94650 4480 94850
rect 4520 94650 4590 94850
rect 4910 94650 4980 94850
rect 5020 94650 5090 94850
rect 5410 94650 5480 94850
rect 5520 94650 5590 94850
rect 5910 94650 5980 94850
rect 6020 94650 6090 94850
rect 6410 94650 6480 94850
rect 6520 94650 6590 94850
rect 6910 94650 6980 94850
rect 7020 94650 7090 94850
rect 7410 94650 7480 94850
rect 7520 94650 7590 94850
rect 7910 94650 7980 94850
rect 8020 94650 8090 94850
rect 8410 94650 8480 94850
rect 8520 94650 8590 94850
rect 8910 94650 8980 94850
rect 9020 94650 9090 94850
rect 9410 94650 9480 94850
rect 9520 94650 9590 94850
rect 9910 94650 9980 94850
rect 10020 94650 10090 94850
rect 10410 94650 10480 94850
rect 10520 94650 10590 94850
rect 10910 94650 10980 94850
rect 11020 94650 11090 94850
rect 11410 94650 11480 94850
rect 11520 94650 11590 94850
rect 11910 94650 11980 94850
rect 12020 94650 12090 94850
rect 12410 94650 12480 94850
rect 12520 94650 12590 94850
rect 12910 94650 12980 94850
rect 13020 94650 13090 94850
rect 13410 94650 13480 94850
rect 13520 94650 13590 94850
rect 13910 94650 13980 94850
rect 14020 94650 14090 94850
rect 14410 94650 14480 94850
rect 14520 94650 14590 94850
rect 14910 94650 14980 94850
rect 15020 94650 15090 94850
rect 15410 94650 15480 94850
rect 15520 94650 15590 94850
rect 15910 94650 15980 94850
rect 16020 94650 16090 94850
rect 16410 94650 16480 94850
rect 16520 94650 16590 94850
rect 16910 94650 16980 94850
rect 17020 94650 17090 94850
rect 17410 94650 17480 94850
rect 17520 94650 17590 94850
rect 17910 94650 17980 94850
rect 18020 94650 18090 94850
rect 18410 94650 18480 94850
rect 18520 94650 18590 94850
rect 18910 94650 18980 94850
rect 19020 94650 19090 94850
rect 19410 94650 19480 94850
rect 19520 94650 19590 94850
rect 19910 94650 19980 94850
rect -15850 94520 -15650 94590
rect -15350 94520 -15150 94590
rect -14850 94520 -14650 94590
rect -14350 94520 -14150 94590
rect -13850 94520 -13650 94590
rect -13350 94520 -13150 94590
rect -12850 94520 -12650 94590
rect -12350 94520 -12150 94590
rect -11850 94520 -11650 94590
rect -11350 94520 -11150 94590
rect -10850 94520 -10650 94590
rect -10350 94520 -10150 94590
rect -9850 94520 -9650 94590
rect -9350 94520 -9150 94590
rect -8850 94520 -8650 94590
rect -8350 94520 -8150 94590
rect -7850 94520 -7650 94590
rect -7350 94520 -7150 94590
rect -6850 94520 -6650 94590
rect -6350 94520 -6150 94590
rect -5850 94520 -5650 94590
rect -5350 94520 -5150 94590
rect -4850 94520 -4650 94590
rect -4350 94520 -4150 94590
rect -3850 94520 -3650 94590
rect -3350 94520 -3150 94590
rect -2850 94520 -2650 94590
rect -2350 94520 -2150 94590
rect -1850 94520 -1650 94590
rect -1350 94520 -1150 94590
rect -850 94520 -650 94590
rect -350 94520 -150 94590
rect 150 94520 350 94590
rect 650 94520 850 94590
rect 1150 94520 1350 94590
rect 1650 94520 1850 94590
rect 2150 94520 2350 94590
rect 2650 94520 2850 94590
rect 3150 94520 3350 94590
rect 3650 94520 3850 94590
rect 4150 94520 4350 94590
rect 4650 94520 4850 94590
rect 5150 94520 5350 94590
rect 5650 94520 5850 94590
rect 6150 94520 6350 94590
rect 6650 94520 6850 94590
rect 7150 94520 7350 94590
rect 7650 94520 7850 94590
rect 8150 94520 8350 94590
rect 8650 94520 8850 94590
rect 9150 94520 9350 94590
rect 9650 94520 9850 94590
rect 10150 94520 10350 94590
rect 10650 94520 10850 94590
rect 11150 94520 11350 94590
rect 11650 94520 11850 94590
rect 12150 94520 12350 94590
rect 12650 94520 12850 94590
rect 13150 94520 13350 94590
rect 13650 94520 13850 94590
rect 14150 94520 14350 94590
rect 14650 94520 14850 94590
rect 15150 94520 15350 94590
rect 15650 94520 15850 94590
rect 16150 94520 16350 94590
rect 16650 94520 16850 94590
rect 17150 94520 17350 94590
rect 17650 94520 17850 94590
rect 18150 94520 18350 94590
rect 18650 94520 18850 94590
rect 19150 94520 19350 94590
rect 19650 94520 19850 94590
rect -15850 94410 -15650 94480
rect -15350 94410 -15150 94480
rect -14850 94410 -14650 94480
rect -14350 94410 -14150 94480
rect -13850 94410 -13650 94480
rect -13350 94410 -13150 94480
rect -12850 94410 -12650 94480
rect -12350 94410 -12150 94480
rect -11850 94410 -11650 94480
rect -11350 94410 -11150 94480
rect -10850 94410 -10650 94480
rect -10350 94410 -10150 94480
rect -9850 94410 -9650 94480
rect -9350 94410 -9150 94480
rect -8850 94410 -8650 94480
rect -8350 94410 -8150 94480
rect -7850 94410 -7650 94480
rect -7350 94410 -7150 94480
rect -6850 94410 -6650 94480
rect -6350 94410 -6150 94480
rect -5850 94410 -5650 94480
rect -5350 94410 -5150 94480
rect -4850 94410 -4650 94480
rect -4350 94410 -4150 94480
rect -3850 94410 -3650 94480
rect -3350 94410 -3150 94480
rect -2850 94410 -2650 94480
rect -2350 94410 -2150 94480
rect -1850 94410 -1650 94480
rect -1350 94410 -1150 94480
rect -850 94410 -650 94480
rect -350 94410 -150 94480
rect 150 94410 350 94480
rect 650 94410 850 94480
rect 1150 94410 1350 94480
rect 1650 94410 1850 94480
rect 2150 94410 2350 94480
rect 2650 94410 2850 94480
rect 3150 94410 3350 94480
rect 3650 94410 3850 94480
rect 4150 94410 4350 94480
rect 4650 94410 4850 94480
rect 5150 94410 5350 94480
rect 5650 94410 5850 94480
rect 6150 94410 6350 94480
rect 6650 94410 6850 94480
rect 7150 94410 7350 94480
rect 7650 94410 7850 94480
rect 8150 94410 8350 94480
rect 8650 94410 8850 94480
rect 9150 94410 9350 94480
rect 9650 94410 9850 94480
rect 10150 94410 10350 94480
rect 10650 94410 10850 94480
rect 11150 94410 11350 94480
rect 11650 94410 11850 94480
rect 12150 94410 12350 94480
rect 12650 94410 12850 94480
rect 13150 94410 13350 94480
rect 13650 94410 13850 94480
rect 14150 94410 14350 94480
rect 14650 94410 14850 94480
rect 15150 94410 15350 94480
rect 15650 94410 15850 94480
rect 16150 94410 16350 94480
rect 16650 94410 16850 94480
rect 17150 94410 17350 94480
rect 17650 94410 17850 94480
rect 18150 94410 18350 94480
rect 18650 94410 18850 94480
rect 19150 94410 19350 94480
rect 19650 94410 19850 94480
rect -15980 94150 -15910 94350
rect -15590 94150 -15520 94350
rect -15480 94150 -15410 94350
rect -15090 94150 -15020 94350
rect -14980 94150 -14910 94350
rect -14590 94150 -14520 94350
rect -14480 94150 -14410 94350
rect -14090 94150 -14020 94350
rect -13980 94150 -13910 94350
rect -13590 94150 -13520 94350
rect -13480 94150 -13410 94350
rect -13090 94150 -13020 94350
rect -12980 94150 -12910 94350
rect -12590 94150 -12520 94350
rect -12480 94150 -12410 94350
rect -12090 94150 -12020 94350
rect -11980 94150 -11910 94350
rect -11590 94150 -11520 94350
rect -11480 94150 -11410 94350
rect -11090 94150 -11020 94350
rect -10980 94150 -10910 94350
rect -10590 94150 -10520 94350
rect -10480 94150 -10410 94350
rect -10090 94150 -10020 94350
rect -9980 94150 -9910 94350
rect -9590 94150 -9520 94350
rect -9480 94150 -9410 94350
rect -9090 94150 -9020 94350
rect -8980 94150 -8910 94350
rect -8590 94150 -8520 94350
rect -8480 94150 -8410 94350
rect -8090 94150 -8020 94350
rect -7980 94150 -7910 94350
rect -7590 94150 -7520 94350
rect -7480 94150 -7410 94350
rect -7090 94150 -7020 94350
rect -6980 94150 -6910 94350
rect -6590 94150 -6520 94350
rect -6480 94150 -6410 94350
rect -6090 94150 -6020 94350
rect -5980 94150 -5910 94350
rect -5590 94150 -5520 94350
rect -5480 94150 -5410 94350
rect -5090 94150 -5020 94350
rect -4980 94150 -4910 94350
rect -4590 94150 -4520 94350
rect -4480 94150 -4410 94350
rect -4090 94150 -4020 94350
rect -3980 94150 -3910 94350
rect -3590 94150 -3520 94350
rect -3480 94150 -3410 94350
rect -3090 94150 -3020 94350
rect -2980 94150 -2910 94350
rect -2590 94150 -2520 94350
rect -2480 94150 -2410 94350
rect -2090 94150 -2020 94350
rect -1980 94150 -1910 94350
rect -1590 94150 -1520 94350
rect -1480 94150 -1410 94350
rect -1090 94150 -1020 94350
rect -980 94150 -910 94350
rect -590 94150 -520 94350
rect -480 94150 -410 94350
rect -90 94150 -20 94350
rect 20 94150 90 94350
rect 410 94150 480 94350
rect 520 94150 590 94350
rect 910 94150 980 94350
rect 1020 94150 1090 94350
rect 1410 94150 1480 94350
rect 1520 94150 1590 94350
rect 1910 94150 1980 94350
rect 2020 94150 2090 94350
rect 2410 94150 2480 94350
rect 2520 94150 2590 94350
rect 2910 94150 2980 94350
rect 3020 94150 3090 94350
rect 3410 94150 3480 94350
rect 3520 94150 3590 94350
rect 3910 94150 3980 94350
rect 4020 94150 4090 94350
rect 4410 94150 4480 94350
rect 4520 94150 4590 94350
rect 4910 94150 4980 94350
rect 5020 94150 5090 94350
rect 5410 94150 5480 94350
rect 5520 94150 5590 94350
rect 5910 94150 5980 94350
rect 6020 94150 6090 94350
rect 6410 94150 6480 94350
rect 6520 94150 6590 94350
rect 6910 94150 6980 94350
rect 7020 94150 7090 94350
rect 7410 94150 7480 94350
rect 7520 94150 7590 94350
rect 7910 94150 7980 94350
rect 8020 94150 8090 94350
rect 8410 94150 8480 94350
rect 8520 94150 8590 94350
rect 8910 94150 8980 94350
rect 9020 94150 9090 94350
rect 9410 94150 9480 94350
rect 9520 94150 9590 94350
rect 9910 94150 9980 94350
rect 10020 94150 10090 94350
rect 10410 94150 10480 94350
rect 10520 94150 10590 94350
rect 10910 94150 10980 94350
rect 11020 94150 11090 94350
rect 11410 94150 11480 94350
rect 11520 94150 11590 94350
rect 11910 94150 11980 94350
rect 12020 94150 12090 94350
rect 12410 94150 12480 94350
rect 12520 94150 12590 94350
rect 12910 94150 12980 94350
rect 13020 94150 13090 94350
rect 13410 94150 13480 94350
rect 13520 94150 13590 94350
rect 13910 94150 13980 94350
rect 14020 94150 14090 94350
rect 14410 94150 14480 94350
rect 14520 94150 14590 94350
rect 14910 94150 14980 94350
rect 15020 94150 15090 94350
rect 15410 94150 15480 94350
rect 15520 94150 15590 94350
rect 15910 94150 15980 94350
rect 16020 94150 16090 94350
rect 16410 94150 16480 94350
rect 16520 94150 16590 94350
rect 16910 94150 16980 94350
rect 17020 94150 17090 94350
rect 17410 94150 17480 94350
rect 17520 94150 17590 94350
rect 17910 94150 17980 94350
rect 18020 94150 18090 94350
rect 18410 94150 18480 94350
rect 18520 94150 18590 94350
rect 18910 94150 18980 94350
rect 19020 94150 19090 94350
rect 19410 94150 19480 94350
rect 19520 94150 19590 94350
rect 19910 94150 19980 94350
rect -15850 94020 -15650 94090
rect -15350 94020 -15150 94090
rect -14850 94020 -14650 94090
rect -14350 94020 -14150 94090
rect -13850 94020 -13650 94090
rect -13350 94020 -13150 94090
rect -12850 94020 -12650 94090
rect -12350 94020 -12150 94090
rect -11850 94020 -11650 94090
rect -11350 94020 -11150 94090
rect -10850 94020 -10650 94090
rect -10350 94020 -10150 94090
rect -9850 94020 -9650 94090
rect -9350 94020 -9150 94090
rect -8850 94020 -8650 94090
rect -8350 94020 -8150 94090
rect -7850 94020 -7650 94090
rect -7350 94020 -7150 94090
rect -6850 94020 -6650 94090
rect -6350 94020 -6150 94090
rect -5850 94020 -5650 94090
rect -5350 94020 -5150 94090
rect -4850 94020 -4650 94090
rect -4350 94020 -4150 94090
rect -3850 94020 -3650 94090
rect -3350 94020 -3150 94090
rect -2850 94020 -2650 94090
rect -2350 94020 -2150 94090
rect -1850 94020 -1650 94090
rect -1350 94020 -1150 94090
rect -850 94020 -650 94090
rect -350 94020 -150 94090
rect 150 94020 350 94090
rect 650 94020 850 94090
rect 1150 94020 1350 94090
rect 1650 94020 1850 94090
rect 2150 94020 2350 94090
rect 2650 94020 2850 94090
rect 3150 94020 3350 94090
rect 3650 94020 3850 94090
rect 4150 94020 4350 94090
rect 4650 94020 4850 94090
rect 5150 94020 5350 94090
rect 5650 94020 5850 94090
rect 6150 94020 6350 94090
rect 6650 94020 6850 94090
rect 7150 94020 7350 94090
rect 7650 94020 7850 94090
rect 8150 94020 8350 94090
rect 8650 94020 8850 94090
rect 9150 94020 9350 94090
rect 9650 94020 9850 94090
rect 10150 94020 10350 94090
rect 10650 94020 10850 94090
rect 11150 94020 11350 94090
rect 11650 94020 11850 94090
rect 12150 94020 12350 94090
rect 12650 94020 12850 94090
rect 13150 94020 13350 94090
rect 13650 94020 13850 94090
rect 14150 94020 14350 94090
rect 14650 94020 14850 94090
rect 15150 94020 15350 94090
rect 15650 94020 15850 94090
rect 16150 94020 16350 94090
rect 16650 94020 16850 94090
rect 17150 94020 17350 94090
rect 17650 94020 17850 94090
rect 18150 94020 18350 94090
rect 18650 94020 18850 94090
rect 19150 94020 19350 94090
rect 19650 94020 19850 94090
rect -15850 93910 -15650 93980
rect -15350 93910 -15150 93980
rect -14850 93910 -14650 93980
rect -14350 93910 -14150 93980
rect -13850 93910 -13650 93980
rect -13350 93910 -13150 93980
rect -12850 93910 -12650 93980
rect -12350 93910 -12150 93980
rect -15980 93650 -15910 93850
rect -15590 93650 -15520 93850
rect -15480 93650 -15410 93850
rect -15090 93650 -15020 93850
rect -14980 93650 -14910 93850
rect -14590 93650 -14520 93850
rect -14480 93650 -14410 93850
rect -14090 93650 -14020 93850
rect -13980 93650 -13910 93850
rect -13590 93650 -13520 93850
rect -13480 93650 -13410 93850
rect -13090 93650 -13020 93850
rect -12980 93650 -12910 93850
rect -12590 93650 -12520 93850
rect -12480 93650 -12410 93850
rect -12090 93650 -12020 93850
rect -15850 93520 -15650 93590
rect -15350 93520 -15150 93590
rect -14850 93520 -14650 93590
rect -14350 93520 -14150 93590
rect -13850 93520 -13650 93590
rect -13350 93520 -13150 93590
rect -12850 93520 -12650 93590
rect -12350 93520 -12150 93590
rect -15850 93410 -15650 93480
rect -15350 93410 -15150 93480
rect -14850 93410 -14650 93480
rect -14350 93410 -14150 93480
rect -13850 93410 -13650 93480
rect -13350 93410 -13150 93480
rect -12850 93410 -12650 93480
rect -12350 93410 -12150 93480
rect -15980 93150 -15910 93350
rect -15590 93150 -15520 93350
rect -15480 93150 -15410 93350
rect -15090 93150 -15020 93350
rect -14980 93150 -14910 93350
rect -14590 93150 -14520 93350
rect -14480 93150 -14410 93350
rect -14090 93150 -14020 93350
rect -13980 93150 -13910 93350
rect -13590 93150 -13520 93350
rect -13480 93150 -13410 93350
rect -13090 93150 -13020 93350
rect -12980 93150 -12910 93350
rect -12590 93150 -12520 93350
rect -12480 93150 -12410 93350
rect -12090 93150 -12020 93350
rect -15850 93020 -15650 93090
rect -15350 93020 -15150 93090
rect -14850 93020 -14650 93090
rect -14350 93020 -14150 93090
rect -13850 93020 -13650 93090
rect -13350 93020 -13150 93090
rect -12850 93020 -12650 93090
rect -12350 93020 -12150 93090
rect -15850 92910 -15650 92980
rect -15350 92910 -15150 92980
rect -14850 92910 -14650 92980
rect -14350 92910 -14150 92980
rect -13850 92910 -13650 92980
rect -13350 92910 -13150 92980
rect -12850 92910 -12650 92980
rect -12350 92910 -12150 92980
rect -15980 92650 -15910 92850
rect -15590 92650 -15520 92850
rect -15480 92650 -15410 92850
rect -15090 92650 -15020 92850
rect -14980 92650 -14910 92850
rect -14590 92650 -14520 92850
rect -14480 92650 -14410 92850
rect -14090 92650 -14020 92850
rect -13980 92650 -13910 92850
rect -13590 92650 -13520 92850
rect -13480 92650 -13410 92850
rect -13090 92650 -13020 92850
rect -12980 92650 -12910 92850
rect -12590 92650 -12520 92850
rect -12480 92650 -12410 92850
rect -12090 92650 -12020 92850
rect -15850 92520 -15650 92590
rect -15350 92520 -15150 92590
rect -14850 92520 -14650 92590
rect -14350 92520 -14150 92590
rect -13850 92520 -13650 92590
rect -13350 92520 -13150 92590
rect -12850 92520 -12650 92590
rect -12350 92520 -12150 92590
rect -15850 92410 -15650 92480
rect -15350 92410 -15150 92480
rect -14850 92410 -14650 92480
rect -14350 92410 -14150 92480
rect -13850 92410 -13650 92480
rect -13350 92410 -13150 92480
rect -12850 92410 -12650 92480
rect -12350 92410 -12150 92480
rect -15980 92150 -15910 92350
rect -15590 92150 -15520 92350
rect -15480 92150 -15410 92350
rect -15090 92150 -15020 92350
rect -14980 92150 -14910 92350
rect -14590 92150 -14520 92350
rect -14480 92150 -14410 92350
rect -14090 92150 -14020 92350
rect -13980 92150 -13910 92350
rect -13590 92150 -13520 92350
rect -13480 92150 -13410 92350
rect -13090 92150 -13020 92350
rect -12980 92150 -12910 92350
rect -12590 92150 -12520 92350
rect -12480 92150 -12410 92350
rect -12090 92150 -12020 92350
rect -15850 92020 -15650 92090
rect -15350 92020 -15150 92090
rect -14850 92020 -14650 92090
rect -14350 92020 -14150 92090
rect -13850 92020 -13650 92090
rect -13350 92020 -13150 92090
rect -12850 92020 -12650 92090
rect -12350 92020 -12150 92090
rect -15850 91910 -15650 91980
rect -15350 91910 -15150 91980
rect -14850 91910 -14650 91980
rect -14350 91910 -14150 91980
rect -13850 91910 -13650 91980
rect -13350 91910 -13150 91980
rect -12850 91910 -12650 91980
rect -12350 91910 -12150 91980
rect -15980 91650 -15910 91850
rect -15590 91650 -15520 91850
rect -15480 91650 -15410 91850
rect -15090 91650 -15020 91850
rect -14980 91650 -14910 91850
rect -14590 91650 -14520 91850
rect -14480 91650 -14410 91850
rect -14090 91650 -14020 91850
rect -13980 91650 -13910 91850
rect -13590 91650 -13520 91850
rect -13480 91650 -13410 91850
rect -13090 91650 -13020 91850
rect -12980 91650 -12910 91850
rect -12590 91650 -12520 91850
rect -12480 91650 -12410 91850
rect -12090 91650 -12020 91850
rect -15850 91520 -15650 91590
rect -15350 91520 -15150 91590
rect -14850 91520 -14650 91590
rect -14350 91520 -14150 91590
rect -13850 91520 -13650 91590
rect -13350 91520 -13150 91590
rect -12850 91520 -12650 91590
rect -12350 91520 -12150 91590
rect -15850 91410 -15650 91480
rect -15350 91410 -15150 91480
rect -14850 91410 -14650 91480
rect -14350 91410 -14150 91480
rect -13850 91410 -13650 91480
rect -13350 91410 -13150 91480
rect -12850 91410 -12650 91480
rect -12350 91410 -12150 91480
rect -15980 91150 -15910 91350
rect -15590 91150 -15520 91350
rect -15480 91150 -15410 91350
rect -15090 91150 -15020 91350
rect -14980 91150 -14910 91350
rect -14590 91150 -14520 91350
rect -14480 91150 -14410 91350
rect -14090 91150 -14020 91350
rect -13980 91150 -13910 91350
rect -13590 91150 -13520 91350
rect -13480 91150 -13410 91350
rect -13090 91150 -13020 91350
rect -12980 91150 -12910 91350
rect -12590 91150 -12520 91350
rect -12480 91150 -12410 91350
rect -12090 91150 -12020 91350
rect -15850 91020 -15650 91090
rect -15350 91020 -15150 91090
rect -14850 91020 -14650 91090
rect -14350 91020 -14150 91090
rect -13850 91020 -13650 91090
rect -13350 91020 -13150 91090
rect -12850 91020 -12650 91090
rect -12350 91020 -12150 91090
rect -15850 90910 -15650 90980
rect -15350 90910 -15150 90980
rect -14850 90910 -14650 90980
rect -14350 90910 -14150 90980
rect -13850 90910 -13650 90980
rect -13350 90910 -13150 90980
rect -12850 90910 -12650 90980
rect -12350 90910 -12150 90980
rect -15980 90650 -15910 90850
rect -15590 90650 -15520 90850
rect -15480 90650 -15410 90850
rect -15090 90650 -15020 90850
rect -14980 90650 -14910 90850
rect -14590 90650 -14520 90850
rect -14480 90650 -14410 90850
rect -14090 90650 -14020 90850
rect -13980 90650 -13910 90850
rect -13590 90650 -13520 90850
rect -13480 90650 -13410 90850
rect -13090 90650 -13020 90850
rect -12980 90650 -12910 90850
rect -12590 90650 -12520 90850
rect -12480 90650 -12410 90850
rect -12090 90650 -12020 90850
rect -15850 90520 -15650 90590
rect -15350 90520 -15150 90590
rect -14850 90520 -14650 90590
rect -14350 90520 -14150 90590
rect -13850 90520 -13650 90590
rect -13350 90520 -13150 90590
rect -12850 90520 -12650 90590
rect -12350 90520 -12150 90590
rect -15850 90410 -15650 90480
rect -15350 90410 -15150 90480
rect -14850 90410 -14650 90480
rect -14350 90410 -14150 90480
rect -13850 90410 -13650 90480
rect -13350 90410 -13150 90480
rect -12850 90410 -12650 90480
rect -12350 90410 -12150 90480
rect -15980 90150 -15910 90350
rect -15590 90150 -15520 90350
rect -15480 90150 -15410 90350
rect -15090 90150 -15020 90350
rect -14980 90150 -14910 90350
rect -14590 90150 -14520 90350
rect -14480 90150 -14410 90350
rect -14090 90150 -14020 90350
rect -13980 90150 -13910 90350
rect -13590 90150 -13520 90350
rect -13480 90150 -13410 90350
rect -13090 90150 -13020 90350
rect -12980 90150 -12910 90350
rect -12590 90150 -12520 90350
rect -12480 90150 -12410 90350
rect -12090 90150 -12020 90350
rect -15850 90020 -15650 90090
rect -15350 90020 -15150 90090
rect -14850 90020 -14650 90090
rect -14350 90020 -14150 90090
rect -13850 90020 -13650 90090
rect -13350 90020 -13150 90090
rect -12850 90020 -12650 90090
rect -12350 90020 -12150 90090
rect -15850 89910 -15650 89980
rect -15350 89910 -15150 89980
rect -14850 89910 -14650 89980
rect -14350 89910 -14150 89980
rect -13850 89910 -13650 89980
rect -13350 89910 -13150 89980
rect -12850 89910 -12650 89980
rect -12350 89910 -12150 89980
rect -15980 89650 -15910 89850
rect -15590 89650 -15520 89850
rect -15480 89650 -15410 89850
rect -15090 89650 -15020 89850
rect -14980 89650 -14910 89850
rect -14590 89650 -14520 89850
rect -14480 89650 -14410 89850
rect -14090 89650 -14020 89850
rect -13980 89650 -13910 89850
rect -13590 89650 -13520 89850
rect -13480 89650 -13410 89850
rect -13090 89650 -13020 89850
rect -12980 89650 -12910 89850
rect -12590 89650 -12520 89850
rect -12480 89650 -12410 89850
rect -12090 89650 -12020 89850
rect -15850 89520 -15650 89590
rect -15350 89520 -15150 89590
rect -14850 89520 -14650 89590
rect -14350 89520 -14150 89590
rect -13850 89520 -13650 89590
rect -13350 89520 -13150 89590
rect -12850 89520 -12650 89590
rect -12350 89520 -12150 89590
rect -15850 89410 -15650 89480
rect -15350 89410 -15150 89480
rect -14850 89410 -14650 89480
rect -14350 89410 -14150 89480
rect -13850 89410 -13650 89480
rect -13350 89410 -13150 89480
rect -12850 89410 -12650 89480
rect -12350 89410 -12150 89480
rect -15980 89150 -15910 89350
rect -15590 89150 -15520 89350
rect -15480 89150 -15410 89350
rect -15090 89150 -15020 89350
rect -14980 89150 -14910 89350
rect -14590 89150 -14520 89350
rect -14480 89150 -14410 89350
rect -14090 89150 -14020 89350
rect -13980 89150 -13910 89350
rect -13590 89150 -13520 89350
rect -13480 89150 -13410 89350
rect -13090 89150 -13020 89350
rect -12980 89150 -12910 89350
rect -12590 89150 -12520 89350
rect -12480 89150 -12410 89350
rect -12090 89150 -12020 89350
rect -15850 89020 -15650 89090
rect -15350 89020 -15150 89090
rect -14850 89020 -14650 89090
rect -14350 89020 -14150 89090
rect -13850 89020 -13650 89090
rect -13350 89020 -13150 89090
rect -12850 89020 -12650 89090
rect -12350 89020 -12150 89090
rect -15850 88910 -15650 88980
rect -15350 88910 -15150 88980
rect -14850 88910 -14650 88980
rect -14350 88910 -14150 88980
rect -13850 88910 -13650 88980
rect -13350 88910 -13150 88980
rect -12850 88910 -12650 88980
rect -12350 88910 -12150 88980
rect -15980 88650 -15910 88850
rect -15590 88650 -15520 88850
rect -15480 88650 -15410 88850
rect -15090 88650 -15020 88850
rect -14980 88650 -14910 88850
rect -14590 88650 -14520 88850
rect -14480 88650 -14410 88850
rect -14090 88650 -14020 88850
rect -13980 88650 -13910 88850
rect -13590 88650 -13520 88850
rect -13480 88650 -13410 88850
rect -13090 88650 -13020 88850
rect -12980 88650 -12910 88850
rect -12590 88650 -12520 88850
rect -12480 88650 -12410 88850
rect -12090 88650 -12020 88850
rect -15850 88520 -15650 88590
rect -15350 88520 -15150 88590
rect -14850 88520 -14650 88590
rect -14350 88520 -14150 88590
rect -13850 88520 -13650 88590
rect -13350 88520 -13150 88590
rect -12850 88520 -12650 88590
rect -12350 88520 -12150 88590
rect -15850 88410 -15650 88480
rect -15350 88410 -15150 88480
rect -14850 88410 -14650 88480
rect -14350 88410 -14150 88480
rect -13850 88410 -13650 88480
rect -13350 88410 -13150 88480
rect -12850 88410 -12650 88480
rect -12350 88410 -12150 88480
rect -15980 88150 -15910 88350
rect -15590 88150 -15520 88350
rect -15480 88150 -15410 88350
rect -15090 88150 -15020 88350
rect -14980 88150 -14910 88350
rect -14590 88150 -14520 88350
rect -14480 88150 -14410 88350
rect -14090 88150 -14020 88350
rect -13980 88150 -13910 88350
rect -13590 88150 -13520 88350
rect -13480 88150 -13410 88350
rect -13090 88150 -13020 88350
rect -12980 88150 -12910 88350
rect -12590 88150 -12520 88350
rect -12480 88150 -12410 88350
rect -12090 88150 -12020 88350
rect -15850 88020 -15650 88090
rect -15350 88020 -15150 88090
rect -14850 88020 -14650 88090
rect -14350 88020 -14150 88090
rect -13850 88020 -13650 88090
rect -13350 88020 -13150 88090
rect -12850 88020 -12650 88090
rect -12350 88020 -12150 88090
rect -15850 87910 -15650 87980
rect -15350 87910 -15150 87980
rect -14850 87910 -14650 87980
rect -14350 87910 -14150 87980
rect -13850 87910 -13650 87980
rect -13350 87910 -13150 87980
rect -12850 87910 -12650 87980
rect -12350 87910 -12150 87980
rect -15980 87650 -15910 87850
rect -15590 87650 -15520 87850
rect -15480 87650 -15410 87850
rect -15090 87650 -15020 87850
rect -14980 87650 -14910 87850
rect -14590 87650 -14520 87850
rect -14480 87650 -14410 87850
rect -14090 87650 -14020 87850
rect -13980 87650 -13910 87850
rect -13590 87650 -13520 87850
rect -13480 87650 -13410 87850
rect -13090 87650 -13020 87850
rect -12980 87650 -12910 87850
rect -12590 87650 -12520 87850
rect -12480 87650 -12410 87850
rect -12090 87650 -12020 87850
rect -15850 87520 -15650 87590
rect -15350 87520 -15150 87590
rect -14850 87520 -14650 87590
rect -14350 87520 -14150 87590
rect -13850 87520 -13650 87590
rect -13350 87520 -13150 87590
rect -12850 87520 -12650 87590
rect -12350 87520 -12150 87590
rect -15850 87410 -15650 87480
rect -15350 87410 -15150 87480
rect -14850 87410 -14650 87480
rect -14350 87410 -14150 87480
rect -13850 87410 -13650 87480
rect -13350 87410 -13150 87480
rect -12850 87410 -12650 87480
rect -12350 87410 -12150 87480
rect -15980 87150 -15910 87350
rect -15590 87150 -15520 87350
rect -15480 87150 -15410 87350
rect -15090 87150 -15020 87350
rect -14980 87150 -14910 87350
rect -14590 87150 -14520 87350
rect -14480 87150 -14410 87350
rect -14090 87150 -14020 87350
rect -13980 87150 -13910 87350
rect -13590 87150 -13520 87350
rect -13480 87150 -13410 87350
rect -13090 87150 -13020 87350
rect -12980 87150 -12910 87350
rect -12590 87150 -12520 87350
rect -12480 87150 -12410 87350
rect -12090 87150 -12020 87350
rect -15850 87020 -15650 87090
rect -15350 87020 -15150 87090
rect -14850 87020 -14650 87090
rect -14350 87020 -14150 87090
rect -13850 87020 -13650 87090
rect -13350 87020 -13150 87090
rect -12850 87020 -12650 87090
rect -12350 87020 -12150 87090
rect -15850 86910 -15650 86980
rect -15350 86910 -15150 86980
rect -14850 86910 -14650 86980
rect -14350 86910 -14150 86980
rect -13850 86910 -13650 86980
rect -13350 86910 -13150 86980
rect -12850 86910 -12650 86980
rect -12350 86910 -12150 86980
rect -15980 86650 -15910 86850
rect -15590 86650 -15520 86850
rect -15480 86650 -15410 86850
rect -15090 86650 -15020 86850
rect -14980 86650 -14910 86850
rect -14590 86650 -14520 86850
rect -14480 86650 -14410 86850
rect -14090 86650 -14020 86850
rect -13980 86650 -13910 86850
rect -13590 86650 -13520 86850
rect -13480 86650 -13410 86850
rect -13090 86650 -13020 86850
rect -12980 86650 -12910 86850
rect -12590 86650 -12520 86850
rect -12480 86650 -12410 86850
rect -12090 86650 -12020 86850
rect -15850 86520 -15650 86590
rect -15350 86520 -15150 86590
rect -14850 86520 -14650 86590
rect -14350 86520 -14150 86590
rect -13850 86520 -13650 86590
rect -13350 86520 -13150 86590
rect -12850 86520 -12650 86590
rect -12350 86520 -12150 86590
rect -15850 86410 -15650 86480
rect -15350 86410 -15150 86480
rect -14850 86410 -14650 86480
rect -14350 86410 -14150 86480
rect -13850 86410 -13650 86480
rect -13350 86410 -13150 86480
rect -12850 86410 -12650 86480
rect -12350 86410 -12150 86480
rect -15980 86150 -15910 86350
rect -15590 86150 -15520 86350
rect -15480 86150 -15410 86350
rect -15090 86150 -15020 86350
rect -14980 86150 -14910 86350
rect -14590 86150 -14520 86350
rect -14480 86150 -14410 86350
rect -14090 86150 -14020 86350
rect -13980 86150 -13910 86350
rect -13590 86150 -13520 86350
rect -13480 86150 -13410 86350
rect -13090 86150 -13020 86350
rect -12980 86150 -12910 86350
rect -12590 86150 -12520 86350
rect -12480 86150 -12410 86350
rect -12090 86150 -12020 86350
rect -15850 86020 -15650 86090
rect -15350 86020 -15150 86090
rect -14850 86020 -14650 86090
rect -14350 86020 -14150 86090
rect -13850 86020 -13650 86090
rect -13350 86020 -13150 86090
rect -12850 86020 -12650 86090
rect -12350 86020 -12150 86090
rect -15850 85910 -15650 85980
rect -15350 85910 -15150 85980
rect -14850 85910 -14650 85980
rect -14350 85910 -14150 85980
rect -13850 85910 -13650 85980
rect -13350 85910 -13150 85980
rect -12850 85910 -12650 85980
rect -12350 85910 -12150 85980
rect -15980 85650 -15910 85850
rect -15590 85650 -15520 85850
rect -15480 85650 -15410 85850
rect -15090 85650 -15020 85850
rect -14980 85650 -14910 85850
rect -14590 85650 -14520 85850
rect -14480 85650 -14410 85850
rect -14090 85650 -14020 85850
rect -13980 85650 -13910 85850
rect -13590 85650 -13520 85850
rect -13480 85650 -13410 85850
rect -13090 85650 -13020 85850
rect -12980 85650 -12910 85850
rect -12590 85650 -12520 85850
rect -12480 85650 -12410 85850
rect -12090 85650 -12020 85850
rect -15850 85520 -15650 85590
rect -15350 85520 -15150 85590
rect -14850 85520 -14650 85590
rect -14350 85520 -14150 85590
rect -13850 85520 -13650 85590
rect -13350 85520 -13150 85590
rect -12850 85520 -12650 85590
rect -12350 85520 -12150 85590
rect -15850 85410 -15650 85480
rect -15350 85410 -15150 85480
rect -14850 85410 -14650 85480
rect -14350 85410 -14150 85480
rect -13850 85410 -13650 85480
rect -13350 85410 -13150 85480
rect -12850 85410 -12650 85480
rect -12350 85410 -12150 85480
rect -15980 85150 -15910 85350
rect -15590 85150 -15520 85350
rect -15480 85150 -15410 85350
rect -15090 85150 -15020 85350
rect -14980 85150 -14910 85350
rect -14590 85150 -14520 85350
rect -14480 85150 -14410 85350
rect -14090 85150 -14020 85350
rect -13980 85150 -13910 85350
rect -13590 85150 -13520 85350
rect -13480 85150 -13410 85350
rect -13090 85150 -13020 85350
rect -12980 85150 -12910 85350
rect -12590 85150 -12520 85350
rect -12480 85150 -12410 85350
rect -12090 85150 -12020 85350
rect -15850 85020 -15650 85090
rect -15350 85020 -15150 85090
rect -14850 85020 -14650 85090
rect -14350 85020 -14150 85090
rect -13850 85020 -13650 85090
rect -13350 85020 -13150 85090
rect -12850 85020 -12650 85090
rect -12350 85020 -12150 85090
rect -15850 84910 -15650 84980
rect -15350 84910 -15150 84980
rect -14850 84910 -14650 84980
rect -14350 84910 -14150 84980
rect -13850 84910 -13650 84980
rect -13350 84910 -13150 84980
rect -12850 84910 -12650 84980
rect -12350 84910 -12150 84980
rect -15980 84650 -15910 84850
rect -15590 84650 -15520 84850
rect -15480 84650 -15410 84850
rect -15090 84650 -15020 84850
rect -14980 84650 -14910 84850
rect -14590 84650 -14520 84850
rect -14480 84650 -14410 84850
rect -14090 84650 -14020 84850
rect -13980 84650 -13910 84850
rect -13590 84650 -13520 84850
rect -13480 84650 -13410 84850
rect -13090 84650 -13020 84850
rect -12980 84650 -12910 84850
rect -12590 84650 -12520 84850
rect -12480 84650 -12410 84850
rect -12090 84650 -12020 84850
rect -15850 84520 -15650 84590
rect -15350 84520 -15150 84590
rect -14850 84520 -14650 84590
rect -14350 84520 -14150 84590
rect -13850 84520 -13650 84590
rect -13350 84520 -13150 84590
rect -12850 84520 -12650 84590
rect -12350 84520 -12150 84590
rect -15850 84410 -15650 84480
rect -15350 84410 -15150 84480
rect -14850 84410 -14650 84480
rect -14350 84410 -14150 84480
rect -13850 84410 -13650 84480
rect -13350 84410 -13150 84480
rect -12850 84410 -12650 84480
rect -12350 84410 -12150 84480
rect -15980 84150 -15910 84350
rect -15590 84150 -15520 84350
rect -15480 84150 -15410 84350
rect -15090 84150 -15020 84350
rect -14980 84150 -14910 84350
rect -14590 84150 -14520 84350
rect -14480 84150 -14410 84350
rect -14090 84150 -14020 84350
rect -13980 84150 -13910 84350
rect -13590 84150 -13520 84350
rect -13480 84150 -13410 84350
rect -13090 84150 -13020 84350
rect -12980 84150 -12910 84350
rect -12590 84150 -12520 84350
rect -12480 84150 -12410 84350
rect -12090 84150 -12020 84350
rect -15850 84020 -15650 84090
rect -15350 84020 -15150 84090
rect -14850 84020 -14650 84090
rect -14350 84020 -14150 84090
rect -13850 84020 -13650 84090
rect -13350 84020 -13150 84090
rect -12850 84020 -12650 84090
rect -12350 84020 -12150 84090
rect -15850 83910 -15650 83980
rect -15350 83910 -15150 83980
rect -14850 83910 -14650 83980
rect -14350 83910 -14150 83980
rect -13850 83910 -13650 83980
rect -13350 83910 -13150 83980
rect -12850 83910 -12650 83980
rect -12350 83910 -12150 83980
rect -15980 83650 -15910 83850
rect -15590 83650 -15520 83850
rect -15480 83650 -15410 83850
rect -15090 83650 -15020 83850
rect -14980 83650 -14910 83850
rect -14590 83650 -14520 83850
rect -14480 83650 -14410 83850
rect -14090 83650 -14020 83850
rect -13980 83650 -13910 83850
rect -13590 83650 -13520 83850
rect -13480 83650 -13410 83850
rect -13090 83650 -13020 83850
rect -12980 83650 -12910 83850
rect -12590 83650 -12520 83850
rect -12480 83650 -12410 83850
rect -12090 83650 -12020 83850
rect -15850 83520 -15650 83590
rect -15350 83520 -15150 83590
rect -14850 83520 -14650 83590
rect -14350 83520 -14150 83590
rect -13850 83520 -13650 83590
rect -13350 83520 -13150 83590
rect -12850 83520 -12650 83590
rect -12350 83520 -12150 83590
rect -15850 83410 -15650 83480
rect -15350 83410 -15150 83480
rect -14850 83410 -14650 83480
rect -14350 83410 -14150 83480
rect -13850 83410 -13650 83480
rect -13350 83410 -13150 83480
rect -12850 83410 -12650 83480
rect -12350 83410 -12150 83480
rect -15980 83150 -15910 83350
rect -15590 83150 -15520 83350
rect -15480 83150 -15410 83350
rect -15090 83150 -15020 83350
rect -14980 83150 -14910 83350
rect -14590 83150 -14520 83350
rect -14480 83150 -14410 83350
rect -14090 83150 -14020 83350
rect -13980 83150 -13910 83350
rect -13590 83150 -13520 83350
rect -13480 83150 -13410 83350
rect -13090 83150 -13020 83350
rect -12980 83150 -12910 83350
rect -12590 83150 -12520 83350
rect -12480 83150 -12410 83350
rect -12090 83150 -12020 83350
rect -15850 83020 -15650 83090
rect -15350 83020 -15150 83090
rect -14850 83020 -14650 83090
rect -14350 83020 -14150 83090
rect -13850 83020 -13650 83090
rect -13350 83020 -13150 83090
rect -12850 83020 -12650 83090
rect -12350 83020 -12150 83090
rect -15850 82910 -15650 82980
rect -15350 82910 -15150 82980
rect -14850 82910 -14650 82980
rect -14350 82910 -14150 82980
rect -13850 82910 -13650 82980
rect -13350 82910 -13150 82980
rect -12850 82910 -12650 82980
rect -12350 82910 -12150 82980
rect -15980 82650 -15910 82850
rect -15590 82650 -15520 82850
rect -15480 82650 -15410 82850
rect -15090 82650 -15020 82850
rect -14980 82650 -14910 82850
rect -14590 82650 -14520 82850
rect -14480 82650 -14410 82850
rect -14090 82650 -14020 82850
rect -13980 82650 -13910 82850
rect -13590 82650 -13520 82850
rect -13480 82650 -13410 82850
rect -13090 82650 -13020 82850
rect -12980 82650 -12910 82850
rect -12590 82650 -12520 82850
rect -12480 82650 -12410 82850
rect -12090 82650 -12020 82850
rect -15850 82520 -15650 82590
rect -15350 82520 -15150 82590
rect -14850 82520 -14650 82590
rect -14350 82520 -14150 82590
rect -13850 82520 -13650 82590
rect -13350 82520 -13150 82590
rect -12850 82520 -12650 82590
rect -12350 82520 -12150 82590
rect -15850 82410 -15650 82480
rect -15350 82410 -15150 82480
rect -14850 82410 -14650 82480
rect -14350 82410 -14150 82480
rect -13850 82410 -13650 82480
rect -13350 82410 -13150 82480
rect -12850 82410 -12650 82480
rect -12350 82410 -12150 82480
rect -15980 82150 -15910 82350
rect -15590 82150 -15520 82350
rect -15480 82150 -15410 82350
rect -15090 82150 -15020 82350
rect -14980 82150 -14910 82350
rect -14590 82150 -14520 82350
rect -14480 82150 -14410 82350
rect -14090 82150 -14020 82350
rect -13980 82150 -13910 82350
rect -13590 82150 -13520 82350
rect -13480 82150 -13410 82350
rect -13090 82150 -13020 82350
rect -12980 82150 -12910 82350
rect -12590 82150 -12520 82350
rect -12480 82150 -12410 82350
rect -12090 82150 -12020 82350
rect -15850 82020 -15650 82090
rect -15350 82020 -15150 82090
rect -14850 82020 -14650 82090
rect -14350 82020 -14150 82090
rect -13850 82020 -13650 82090
rect -13350 82020 -13150 82090
rect -12850 82020 -12650 82090
rect -12350 82020 -12150 82090
rect -15850 81910 -15650 81980
rect -15350 81910 -15150 81980
rect -14850 81910 -14650 81980
rect -14350 81910 -14150 81980
rect -13850 81910 -13650 81980
rect -13350 81910 -13150 81980
rect -12850 81910 -12650 81980
rect -12350 81910 -12150 81980
rect -15980 81650 -15910 81850
rect -15590 81650 -15520 81850
rect -15480 81650 -15410 81850
rect -15090 81650 -15020 81850
rect -14980 81650 -14910 81850
rect -14590 81650 -14520 81850
rect -14480 81650 -14410 81850
rect -14090 81650 -14020 81850
rect -13980 81650 -13910 81850
rect -13590 81650 -13520 81850
rect -13480 81650 -13410 81850
rect -13090 81650 -13020 81850
rect -12980 81650 -12910 81850
rect -12590 81650 -12520 81850
rect -12480 81650 -12410 81850
rect -12090 81650 -12020 81850
rect -15850 81520 -15650 81590
rect -15350 81520 -15150 81590
rect -14850 81520 -14650 81590
rect -14350 81520 -14150 81590
rect -13850 81520 -13650 81590
rect -13350 81520 -13150 81590
rect -12850 81520 -12650 81590
rect -12350 81520 -12150 81590
rect -15850 81410 -15650 81480
rect -15350 81410 -15150 81480
rect -14850 81410 -14650 81480
rect -14350 81410 -14150 81480
rect -13850 81410 -13650 81480
rect -13350 81410 -13150 81480
rect -12850 81410 -12650 81480
rect -12350 81410 -12150 81480
rect -15980 81150 -15910 81350
rect -15590 81150 -15520 81350
rect -15480 81150 -15410 81350
rect -15090 81150 -15020 81350
rect -14980 81150 -14910 81350
rect -14590 81150 -14520 81350
rect -14480 81150 -14410 81350
rect -14090 81150 -14020 81350
rect -13980 81150 -13910 81350
rect -13590 81150 -13520 81350
rect -13480 81150 -13410 81350
rect -13090 81150 -13020 81350
rect -12980 81150 -12910 81350
rect -12590 81150 -12520 81350
rect -12480 81150 -12410 81350
rect -12090 81150 -12020 81350
rect -15850 81020 -15650 81090
rect -15350 81020 -15150 81090
rect -14850 81020 -14650 81090
rect -14350 81020 -14150 81090
rect -13850 81020 -13650 81090
rect -13350 81020 -13150 81090
rect -12850 81020 -12650 81090
rect -12350 81020 -12150 81090
rect -15850 80910 -15650 80980
rect -15350 80910 -15150 80980
rect -14850 80910 -14650 80980
rect -14350 80910 -14150 80980
rect -13850 80910 -13650 80980
rect -13350 80910 -13150 80980
rect -12850 80910 -12650 80980
rect -12350 80910 -12150 80980
rect -15980 80650 -15910 80850
rect -15590 80650 -15520 80850
rect -15480 80650 -15410 80850
rect -15090 80650 -15020 80850
rect -14980 80650 -14910 80850
rect -14590 80650 -14520 80850
rect -14480 80650 -14410 80850
rect -14090 80650 -14020 80850
rect -13980 80650 -13910 80850
rect -13590 80650 -13520 80850
rect -13480 80650 -13410 80850
rect -13090 80650 -13020 80850
rect -12980 80650 -12910 80850
rect -12590 80650 -12520 80850
rect -12480 80650 -12410 80850
rect -12090 80650 -12020 80850
rect -15850 80520 -15650 80590
rect -15350 80520 -15150 80590
rect -14850 80520 -14650 80590
rect -14350 80520 -14150 80590
rect -13850 80520 -13650 80590
rect -13350 80520 -13150 80590
rect -12850 80520 -12650 80590
rect -12350 80520 -12150 80590
rect -15850 80410 -15650 80480
rect -15350 80410 -15150 80480
rect -14850 80410 -14650 80480
rect -14350 80410 -14150 80480
rect -13850 80410 -13650 80480
rect -13350 80410 -13150 80480
rect -12850 80410 -12650 80480
rect -12350 80410 -12150 80480
rect -15980 80150 -15910 80350
rect -15590 80150 -15520 80350
rect -15480 80150 -15410 80350
rect -15090 80150 -15020 80350
rect -14980 80150 -14910 80350
rect -14590 80150 -14520 80350
rect -14480 80150 -14410 80350
rect -14090 80150 -14020 80350
rect -13980 80150 -13910 80350
rect -13590 80150 -13520 80350
rect -13480 80150 -13410 80350
rect -13090 80150 -13020 80350
rect -12980 80150 -12910 80350
rect -12590 80150 -12520 80350
rect -12480 80150 -12410 80350
rect -12090 80150 -12020 80350
rect -15850 80020 -15650 80090
rect -15350 80020 -15150 80090
rect -14850 80020 -14650 80090
rect -14350 80020 -14150 80090
rect -13850 80020 -13650 80090
rect -13350 80020 -13150 80090
rect -12850 80020 -12650 80090
rect -12350 80020 -12150 80090
rect -15850 79910 -15650 79980
rect -15350 79910 -15150 79980
rect -14850 79910 -14650 79980
rect -14350 79910 -14150 79980
rect -13850 79910 -13650 79980
rect -13350 79910 -13150 79980
rect -12850 79910 -12650 79980
rect -12350 79910 -12150 79980
rect -15980 79650 -15910 79850
rect -15590 79650 -15520 79850
rect -15480 79650 -15410 79850
rect -15090 79650 -15020 79850
rect -14980 79650 -14910 79850
rect -14590 79650 -14520 79850
rect -14480 79650 -14410 79850
rect -14090 79650 -14020 79850
rect -13980 79650 -13910 79850
rect -13590 79650 -13520 79850
rect -13480 79650 -13410 79850
rect -13090 79650 -13020 79850
rect -12980 79650 -12910 79850
rect -12590 79650 -12520 79850
rect -12480 79650 -12410 79850
rect -12090 79650 -12020 79850
rect -15850 79520 -15650 79590
rect -15350 79520 -15150 79590
rect -14850 79520 -14650 79590
rect -14350 79520 -14150 79590
rect -13850 79520 -13650 79590
rect -13350 79520 -13150 79590
rect -12850 79520 -12650 79590
rect -12350 79520 -12150 79590
rect -15850 79410 -15650 79480
rect -15350 79410 -15150 79480
rect -14850 79410 -14650 79480
rect -14350 79410 -14150 79480
rect -13850 79410 -13650 79480
rect -13350 79410 -13150 79480
rect -12850 79410 -12650 79480
rect -12350 79410 -12150 79480
rect -15980 79150 -15910 79350
rect -15590 79150 -15520 79350
rect -15480 79150 -15410 79350
rect -15090 79150 -15020 79350
rect -14980 79150 -14910 79350
rect -14590 79150 -14520 79350
rect -14480 79150 -14410 79350
rect -14090 79150 -14020 79350
rect -13980 79150 -13910 79350
rect -13590 79150 -13520 79350
rect -13480 79150 -13410 79350
rect -13090 79150 -13020 79350
rect -12980 79150 -12910 79350
rect -12590 79150 -12520 79350
rect -12480 79150 -12410 79350
rect -12090 79150 -12020 79350
rect -15850 79020 -15650 79090
rect -15350 79020 -15150 79090
rect -14850 79020 -14650 79090
rect -14350 79020 -14150 79090
rect -13850 79020 -13650 79090
rect -13350 79020 -13150 79090
rect -12850 79020 -12650 79090
rect -12350 79020 -12150 79090
rect -15850 78910 -15650 78980
rect -15350 78910 -15150 78980
rect -14850 78910 -14650 78980
rect -14350 78910 -14150 78980
rect -13850 78910 -13650 78980
rect -13350 78910 -13150 78980
rect -12850 78910 -12650 78980
rect -12350 78910 -12150 78980
rect -15980 78650 -15910 78850
rect -15590 78650 -15520 78850
rect -15480 78650 -15410 78850
rect -15090 78650 -15020 78850
rect -14980 78650 -14910 78850
rect -14590 78650 -14520 78850
rect -14480 78650 -14410 78850
rect -14090 78650 -14020 78850
rect -13980 78650 -13910 78850
rect -13590 78650 -13520 78850
rect -13480 78650 -13410 78850
rect -13090 78650 -13020 78850
rect -12980 78650 -12910 78850
rect -12590 78650 -12520 78850
rect -12480 78650 -12410 78850
rect -12090 78650 -12020 78850
rect -15850 78520 -15650 78590
rect -15350 78520 -15150 78590
rect -14850 78520 -14650 78590
rect -14350 78520 -14150 78590
rect -13850 78520 -13650 78590
rect -13350 78520 -13150 78590
rect -12850 78520 -12650 78590
rect -12350 78520 -12150 78590
rect -15850 78410 -15650 78480
rect -15350 78410 -15150 78480
rect -14850 78410 -14650 78480
rect -14350 78410 -14150 78480
rect -13850 78410 -13650 78480
rect -13350 78410 -13150 78480
rect -12850 78410 -12650 78480
rect -12350 78410 -12150 78480
rect -15980 78150 -15910 78350
rect -15590 78150 -15520 78350
rect -15480 78150 -15410 78350
rect -15090 78150 -15020 78350
rect -14980 78150 -14910 78350
rect -14590 78150 -14520 78350
rect -14480 78150 -14410 78350
rect -14090 78150 -14020 78350
rect -13980 78150 -13910 78350
rect -13590 78150 -13520 78350
rect -13480 78150 -13410 78350
rect -13090 78150 -13020 78350
rect -12980 78150 -12910 78350
rect -12590 78150 -12520 78350
rect -12480 78150 -12410 78350
rect -12090 78150 -12020 78350
rect -15850 78020 -15650 78090
rect -15350 78020 -15150 78090
rect -14850 78020 -14650 78090
rect -14350 78020 -14150 78090
rect -13850 78020 -13650 78090
rect -13350 78020 -13150 78090
rect -12850 78020 -12650 78090
rect -12350 78020 -12150 78090
rect -15850 77910 -15650 77980
rect -15350 77910 -15150 77980
rect -14850 77910 -14650 77980
rect -14350 77910 -14150 77980
rect -13850 77910 -13650 77980
rect -13350 77910 -13150 77980
rect -12850 77910 -12650 77980
rect -12350 77910 -12150 77980
rect -15980 77650 -15910 77850
rect -15590 77650 -15520 77850
rect -15480 77650 -15410 77850
rect -15090 77650 -15020 77850
rect -14980 77650 -14910 77850
rect -14590 77650 -14520 77850
rect -14480 77650 -14410 77850
rect -14090 77650 -14020 77850
rect -13980 77650 -13910 77850
rect -13590 77650 -13520 77850
rect -13480 77650 -13410 77850
rect -13090 77650 -13020 77850
rect -12980 77650 -12910 77850
rect -12590 77650 -12520 77850
rect -12480 77650 -12410 77850
rect -12090 77650 -12020 77850
rect -15850 77520 -15650 77590
rect -15350 77520 -15150 77590
rect -14850 77520 -14650 77590
rect -14350 77520 -14150 77590
rect -13850 77520 -13650 77590
rect -13350 77520 -13150 77590
rect -12850 77520 -12650 77590
rect -12350 77520 -12150 77590
rect -15850 77410 -15650 77480
rect -15350 77410 -15150 77480
rect -14850 77410 -14650 77480
rect -14350 77410 -14150 77480
rect -13850 77410 -13650 77480
rect -13350 77410 -13150 77480
rect -12850 77410 -12650 77480
rect -12350 77410 -12150 77480
rect -15980 77150 -15910 77350
rect -15590 77150 -15520 77350
rect -15480 77150 -15410 77350
rect -15090 77150 -15020 77350
rect -14980 77150 -14910 77350
rect -14590 77150 -14520 77350
rect -14480 77150 -14410 77350
rect -14090 77150 -14020 77350
rect -13980 77150 -13910 77350
rect -13590 77150 -13520 77350
rect -13480 77150 -13410 77350
rect -13090 77150 -13020 77350
rect -12980 77150 -12910 77350
rect -12590 77150 -12520 77350
rect -12480 77150 -12410 77350
rect -12090 77150 -12020 77350
rect -15850 77020 -15650 77090
rect -15350 77020 -15150 77090
rect -14850 77020 -14650 77090
rect -14350 77020 -14150 77090
rect -13850 77020 -13650 77090
rect -13350 77020 -13150 77090
rect -12850 77020 -12650 77090
rect -12350 77020 -12150 77090
rect -15850 76910 -15650 76980
rect -15350 76910 -15150 76980
rect -14850 76910 -14650 76980
rect -14350 76910 -14150 76980
rect -13850 76910 -13650 76980
rect -13350 76910 -13150 76980
rect -12850 76910 -12650 76980
rect -12350 76910 -12150 76980
rect -15980 76650 -15910 76850
rect -15590 76650 -15520 76850
rect -15480 76650 -15410 76850
rect -15090 76650 -15020 76850
rect -14980 76650 -14910 76850
rect -14590 76650 -14520 76850
rect -14480 76650 -14410 76850
rect -14090 76650 -14020 76850
rect -13980 76650 -13910 76850
rect -13590 76650 -13520 76850
rect -13480 76650 -13410 76850
rect -13090 76650 -13020 76850
rect -12980 76650 -12910 76850
rect -12590 76650 -12520 76850
rect -12480 76650 -12410 76850
rect -12090 76650 -12020 76850
rect -15850 76520 -15650 76590
rect -15350 76520 -15150 76590
rect -14850 76520 -14650 76590
rect -14350 76520 -14150 76590
rect -13850 76520 -13650 76590
rect -13350 76520 -13150 76590
rect -12850 76520 -12650 76590
rect -12350 76520 -12150 76590
rect -15850 76410 -15650 76480
rect -15350 76410 -15150 76480
rect -14850 76410 -14650 76480
rect -14350 76410 -14150 76480
rect -13850 76410 -13650 76480
rect -13350 76410 -13150 76480
rect -12850 76410 -12650 76480
rect -12350 76410 -12150 76480
rect -15980 76150 -15910 76350
rect -15590 76150 -15520 76350
rect -15480 76150 -15410 76350
rect -15090 76150 -15020 76350
rect -14980 76150 -14910 76350
rect -14590 76150 -14520 76350
rect -14480 76150 -14410 76350
rect -14090 76150 -14020 76350
rect -13980 76150 -13910 76350
rect -13590 76150 -13520 76350
rect -13480 76150 -13410 76350
rect -13090 76150 -13020 76350
rect -12980 76150 -12910 76350
rect -12590 76150 -12520 76350
rect -12480 76150 -12410 76350
rect -12090 76150 -12020 76350
rect -15850 76020 -15650 76090
rect -15350 76020 -15150 76090
rect -14850 76020 -14650 76090
rect -14350 76020 -14150 76090
rect -13850 76020 -13650 76090
rect -13350 76020 -13150 76090
rect -12850 76020 -12650 76090
rect -12350 76020 -12150 76090
rect -15850 75910 -15650 75980
rect -15350 75910 -15150 75980
rect -14850 75910 -14650 75980
rect -14350 75910 -14150 75980
rect -13850 75910 -13650 75980
rect -13350 75910 -13150 75980
rect -12850 75910 -12650 75980
rect -12350 75910 -12150 75980
rect -15980 75650 -15910 75850
rect -15590 75650 -15520 75850
rect -15480 75650 -15410 75850
rect -15090 75650 -15020 75850
rect -14980 75650 -14910 75850
rect -14590 75650 -14520 75850
rect -14480 75650 -14410 75850
rect -14090 75650 -14020 75850
rect -13980 75650 -13910 75850
rect -13590 75650 -13520 75850
rect -13480 75650 -13410 75850
rect -13090 75650 -13020 75850
rect -12980 75650 -12910 75850
rect -12590 75650 -12520 75850
rect -12480 75650 -12410 75850
rect -12090 75650 -12020 75850
rect -15850 75520 -15650 75590
rect -15350 75520 -15150 75590
rect -14850 75520 -14650 75590
rect -14350 75520 -14150 75590
rect -13850 75520 -13650 75590
rect -13350 75520 -13150 75590
rect -12850 75520 -12650 75590
rect -12350 75520 -12150 75590
rect -15850 75410 -15650 75480
rect -15350 75410 -15150 75480
rect -14850 75410 -14650 75480
rect -14350 75410 -14150 75480
rect -13850 75410 -13650 75480
rect -13350 75410 -13150 75480
rect -12850 75410 -12650 75480
rect -12350 75410 -12150 75480
rect -15980 75150 -15910 75350
rect -15590 75150 -15520 75350
rect -15480 75150 -15410 75350
rect -15090 75150 -15020 75350
rect -14980 75150 -14910 75350
rect -14590 75150 -14520 75350
rect -14480 75150 -14410 75350
rect -14090 75150 -14020 75350
rect -13980 75150 -13910 75350
rect -13590 75150 -13520 75350
rect -13480 75150 -13410 75350
rect -13090 75150 -13020 75350
rect -12980 75150 -12910 75350
rect -12590 75150 -12520 75350
rect -12480 75150 -12410 75350
rect -12090 75150 -12020 75350
rect -15850 75020 -15650 75090
rect -15350 75020 -15150 75090
rect -14850 75020 -14650 75090
rect -14350 75020 -14150 75090
rect -13850 75020 -13650 75090
rect -13350 75020 -13150 75090
rect -12850 75020 -12650 75090
rect -12350 75020 -12150 75090
rect -15850 74910 -15650 74980
rect -15350 74910 -15150 74980
rect -14850 74910 -14650 74980
rect -14350 74910 -14150 74980
rect -13850 74910 -13650 74980
rect -13350 74910 -13150 74980
rect -12850 74910 -12650 74980
rect -12350 74910 -12150 74980
rect -15980 74650 -15910 74850
rect -15590 74650 -15520 74850
rect -15480 74650 -15410 74850
rect -15090 74650 -15020 74850
rect -14980 74650 -14910 74850
rect -14590 74650 -14520 74850
rect -14480 74650 -14410 74850
rect -14090 74650 -14020 74850
rect -13980 74650 -13910 74850
rect -13590 74650 -13520 74850
rect -13480 74650 -13410 74850
rect -13090 74650 -13020 74850
rect -12980 74650 -12910 74850
rect -12590 74650 -12520 74850
rect -12480 74650 -12410 74850
rect -12090 74650 -12020 74850
rect -15850 74520 -15650 74590
rect -15350 74520 -15150 74590
rect -14850 74520 -14650 74590
rect -14350 74520 -14150 74590
rect -13850 74520 -13650 74590
rect -13350 74520 -13150 74590
rect -12850 74520 -12650 74590
rect -12350 74520 -12150 74590
rect -15850 74410 -15650 74480
rect -15350 74410 -15150 74480
rect -14850 74410 -14650 74480
rect -14350 74410 -14150 74480
rect -13850 74410 -13650 74480
rect -13350 74410 -13150 74480
rect -12850 74410 -12650 74480
rect -12350 74410 -12150 74480
rect -15980 74150 -15910 74350
rect -15590 74150 -15520 74350
rect -15480 74150 -15410 74350
rect -15090 74150 -15020 74350
rect -14980 74150 -14910 74350
rect -14590 74150 -14520 74350
rect -14480 74150 -14410 74350
rect -14090 74150 -14020 74350
rect -13980 74150 -13910 74350
rect -13590 74150 -13520 74350
rect -13480 74150 -13410 74350
rect -13090 74150 -13020 74350
rect -12980 74150 -12910 74350
rect -12590 74150 -12520 74350
rect -12480 74150 -12410 74350
rect -12090 74150 -12020 74350
rect -15850 74020 -15650 74090
rect -15350 74020 -15150 74090
rect -14850 74020 -14650 74090
rect -14350 74020 -14150 74090
rect -13850 74020 -13650 74090
rect -13350 74020 -13150 74090
rect -12850 74020 -12650 74090
rect -12350 74020 -12150 74090
rect -15850 73910 -15650 73980
rect -15350 73910 -15150 73980
rect -14850 73910 -14650 73980
rect -14350 73910 -14150 73980
rect -13850 73910 -13650 73980
rect -13350 73910 -13150 73980
rect -12850 73910 -12650 73980
rect -12350 73910 -12150 73980
rect -15980 73650 -15910 73850
rect -15590 73650 -15520 73850
rect -15480 73650 -15410 73850
rect -15090 73650 -15020 73850
rect -14980 73650 -14910 73850
rect -14590 73650 -14520 73850
rect -14480 73650 -14410 73850
rect -14090 73650 -14020 73850
rect -13980 73650 -13910 73850
rect -13590 73650 -13520 73850
rect -13480 73650 -13410 73850
rect -13090 73650 -13020 73850
rect -12980 73650 -12910 73850
rect -12590 73650 -12520 73850
rect -12480 73650 -12410 73850
rect -12090 73650 -12020 73850
rect -15850 73520 -15650 73590
rect -15350 73520 -15150 73590
rect -14850 73520 -14650 73590
rect -14350 73520 -14150 73590
rect -13850 73520 -13650 73590
rect -13350 73520 -13150 73590
rect -12850 73520 -12650 73590
rect -12350 73520 -12150 73590
rect -15850 73410 -15650 73480
rect -15350 73410 -15150 73480
rect -14850 73410 -14650 73480
rect -14350 73410 -14150 73480
rect -13850 73410 -13650 73480
rect -13350 73410 -13150 73480
rect -12850 73410 -12650 73480
rect -12350 73410 -12150 73480
rect -15980 73150 -15910 73350
rect -15590 73150 -15520 73350
rect -15480 73150 -15410 73350
rect -15090 73150 -15020 73350
rect -14980 73150 -14910 73350
rect -14590 73150 -14520 73350
rect -14480 73150 -14410 73350
rect -14090 73150 -14020 73350
rect -13980 73150 -13910 73350
rect -13590 73150 -13520 73350
rect -13480 73150 -13410 73350
rect -13090 73150 -13020 73350
rect -12980 73150 -12910 73350
rect -12590 73150 -12520 73350
rect -12480 73150 -12410 73350
rect -12090 73150 -12020 73350
rect -15850 73020 -15650 73090
rect -15350 73020 -15150 73090
rect -14850 73020 -14650 73090
rect -14350 73020 -14150 73090
rect -13850 73020 -13650 73090
rect -13350 73020 -13150 73090
rect -12850 73020 -12650 73090
rect -12350 73020 -12150 73090
rect -15850 72910 -15650 72980
rect -15350 72910 -15150 72980
rect -14850 72910 -14650 72980
rect -14350 72910 -14150 72980
rect -13850 72910 -13650 72980
rect -13350 72910 -13150 72980
rect -12850 72910 -12650 72980
rect -12350 72910 -12150 72980
rect -15980 72650 -15910 72850
rect -15590 72650 -15520 72850
rect -15480 72650 -15410 72850
rect -15090 72650 -15020 72850
rect -14980 72650 -14910 72850
rect -14590 72650 -14520 72850
rect -14480 72650 -14410 72850
rect -14090 72650 -14020 72850
rect -13980 72650 -13910 72850
rect -13590 72650 -13520 72850
rect -13480 72650 -13410 72850
rect -13090 72650 -13020 72850
rect -12980 72650 -12910 72850
rect -12590 72650 -12520 72850
rect -12480 72650 -12410 72850
rect -12090 72650 -12020 72850
rect -15850 72520 -15650 72590
rect -15350 72520 -15150 72590
rect -14850 72520 -14650 72590
rect -14350 72520 -14150 72590
rect -13850 72520 -13650 72590
rect -13350 72520 -13150 72590
rect -12850 72520 -12650 72590
rect -12350 72520 -12150 72590
rect -15850 72410 -15650 72480
rect -15350 72410 -15150 72480
rect -14850 72410 -14650 72480
rect -14350 72410 -14150 72480
rect -13850 72410 -13650 72480
rect -13350 72410 -13150 72480
rect -12850 72410 -12650 72480
rect -12350 72410 -12150 72480
rect -15980 72150 -15910 72350
rect -15590 72150 -15520 72350
rect -15480 72150 -15410 72350
rect -15090 72150 -15020 72350
rect -14980 72150 -14910 72350
rect -14590 72150 -14520 72350
rect -14480 72150 -14410 72350
rect -14090 72150 -14020 72350
rect -13980 72150 -13910 72350
rect -13590 72150 -13520 72350
rect -13480 72150 -13410 72350
rect -13090 72150 -13020 72350
rect -12980 72150 -12910 72350
rect -12590 72150 -12520 72350
rect -12480 72150 -12410 72350
rect -12090 72150 -12020 72350
rect -15850 72020 -15650 72090
rect -15350 72020 -15150 72090
rect -14850 72020 -14650 72090
rect -14350 72020 -14150 72090
rect -13850 72020 -13650 72090
rect -13350 72020 -13150 72090
rect -12850 72020 -12650 72090
rect -12350 72020 -12150 72090
rect -15850 71910 -15650 71980
rect -15350 71910 -15150 71980
rect -14850 71910 -14650 71980
rect -14350 71910 -14150 71980
rect -13850 71910 -13650 71980
rect -13350 71910 -13150 71980
rect -12850 71910 -12650 71980
rect -12350 71910 -12150 71980
rect -15980 71650 -15910 71850
rect -15590 71650 -15520 71850
rect -15480 71650 -15410 71850
rect -15090 71650 -15020 71850
rect -14980 71650 -14910 71850
rect -14590 71650 -14520 71850
rect -14480 71650 -14410 71850
rect -14090 71650 -14020 71850
rect -13980 71650 -13910 71850
rect -13590 71650 -13520 71850
rect -13480 71650 -13410 71850
rect -13090 71650 -13020 71850
rect -12980 71650 -12910 71850
rect -12590 71650 -12520 71850
rect -12480 71650 -12410 71850
rect -12090 71650 -12020 71850
rect -15850 71520 -15650 71590
rect -15350 71520 -15150 71590
rect -14850 71520 -14650 71590
rect -14350 71520 -14150 71590
rect -13850 71520 -13650 71590
rect -13350 71520 -13150 71590
rect -12850 71520 -12650 71590
rect -12350 71520 -12150 71590
rect -15850 71410 -15650 71480
rect -15350 71410 -15150 71480
rect -14850 71410 -14650 71480
rect -14350 71410 -14150 71480
rect -13850 71410 -13650 71480
rect -13350 71410 -13150 71480
rect -12850 71410 -12650 71480
rect -12350 71410 -12150 71480
rect -15980 71150 -15910 71350
rect -15590 71150 -15520 71350
rect -15480 71150 -15410 71350
rect -15090 71150 -15020 71350
rect -14980 71150 -14910 71350
rect -14590 71150 -14520 71350
rect -14480 71150 -14410 71350
rect -14090 71150 -14020 71350
rect -13980 71150 -13910 71350
rect -13590 71150 -13520 71350
rect -13480 71150 -13410 71350
rect -13090 71150 -13020 71350
rect -12980 71150 -12910 71350
rect -12590 71150 -12520 71350
rect -12480 71150 -12410 71350
rect -12090 71150 -12020 71350
rect -15850 71020 -15650 71090
rect -15350 71020 -15150 71090
rect -14850 71020 -14650 71090
rect -14350 71020 -14150 71090
rect -13850 71020 -13650 71090
rect -13350 71020 -13150 71090
rect -12850 71020 -12650 71090
rect -12350 71020 -12150 71090
rect -15850 70910 -15650 70980
rect -15350 70910 -15150 70980
rect -14850 70910 -14650 70980
rect -14350 70910 -14150 70980
rect -13850 70910 -13650 70980
rect -13350 70910 -13150 70980
rect -12850 70910 -12650 70980
rect -12350 70910 -12150 70980
rect -15980 70650 -15910 70850
rect -15590 70650 -15520 70850
rect -15480 70650 -15410 70850
rect -15090 70650 -15020 70850
rect -14980 70650 -14910 70850
rect -14590 70650 -14520 70850
rect -14480 70650 -14410 70850
rect -14090 70650 -14020 70850
rect -13980 70650 -13910 70850
rect -13590 70650 -13520 70850
rect -13480 70650 -13410 70850
rect -13090 70650 -13020 70850
rect -12980 70650 -12910 70850
rect -12590 70650 -12520 70850
rect -12480 70650 -12410 70850
rect -12090 70650 -12020 70850
rect -15850 70520 -15650 70590
rect -15350 70520 -15150 70590
rect -14850 70520 -14650 70590
rect -14350 70520 -14150 70590
rect -13850 70520 -13650 70590
rect -13350 70520 -13150 70590
rect -12850 70520 -12650 70590
rect -12350 70520 -12150 70590
rect -15850 70410 -15650 70480
rect -15350 70410 -15150 70480
rect -14850 70410 -14650 70480
rect -14350 70410 -14150 70480
rect -13850 70410 -13650 70480
rect -13350 70410 -13150 70480
rect -12850 70410 -12650 70480
rect -12350 70410 -12150 70480
rect -15980 70150 -15910 70350
rect -15590 70150 -15520 70350
rect -15480 70150 -15410 70350
rect -15090 70150 -15020 70350
rect -14980 70150 -14910 70350
rect -14590 70150 -14520 70350
rect -14480 70150 -14410 70350
rect -14090 70150 -14020 70350
rect -13980 70150 -13910 70350
rect -13590 70150 -13520 70350
rect -13480 70150 -13410 70350
rect -13090 70150 -13020 70350
rect -12980 70150 -12910 70350
rect -12590 70150 -12520 70350
rect -12480 70150 -12410 70350
rect -12090 70150 -12020 70350
rect -15850 70020 -15650 70090
rect -15350 70020 -15150 70090
rect -14850 70020 -14650 70090
rect -14350 70020 -14150 70090
rect -13850 70020 -13650 70090
rect -13350 70020 -13150 70090
rect -12850 70020 -12650 70090
rect -12350 70020 -12150 70090
rect -15850 69910 -15650 69980
rect -15350 69910 -15150 69980
rect -14850 69910 -14650 69980
rect -14350 69910 -14150 69980
rect -13850 69910 -13650 69980
rect -13350 69910 -13150 69980
rect -12850 69910 -12650 69980
rect -12350 69910 -12150 69980
rect -15980 69650 -15910 69850
rect -15590 69650 -15520 69850
rect -15480 69650 -15410 69850
rect -15090 69650 -15020 69850
rect -14980 69650 -14910 69850
rect -14590 69650 -14520 69850
rect -14480 69650 -14410 69850
rect -14090 69650 -14020 69850
rect -13980 69650 -13910 69850
rect -13590 69650 -13520 69850
rect -13480 69650 -13410 69850
rect -13090 69650 -13020 69850
rect -12980 69650 -12910 69850
rect -12590 69650 -12520 69850
rect -12480 69650 -12410 69850
rect -12090 69650 -12020 69850
rect -15850 69520 -15650 69590
rect -15350 69520 -15150 69590
rect -14850 69520 -14650 69590
rect -14350 69520 -14150 69590
rect -13850 69520 -13650 69590
rect -13350 69520 -13150 69590
rect -12850 69520 -12650 69590
rect -12350 69520 -12150 69590
rect -15850 69410 -15650 69480
rect -15350 69410 -15150 69480
rect -14850 69410 -14650 69480
rect -14350 69410 -14150 69480
rect -13850 69410 -13650 69480
rect -13350 69410 -13150 69480
rect -12850 69410 -12650 69480
rect -12350 69410 -12150 69480
rect -15980 69150 -15910 69350
rect -15590 69150 -15520 69350
rect -15480 69150 -15410 69350
rect -15090 69150 -15020 69350
rect -14980 69150 -14910 69350
rect -14590 69150 -14520 69350
rect -14480 69150 -14410 69350
rect -14090 69150 -14020 69350
rect -13980 69150 -13910 69350
rect -13590 69150 -13520 69350
rect -13480 69150 -13410 69350
rect -13090 69150 -13020 69350
rect -12980 69150 -12910 69350
rect -12590 69150 -12520 69350
rect -12480 69150 -12410 69350
rect -12090 69150 -12020 69350
rect -15850 69020 -15650 69090
rect -15350 69020 -15150 69090
rect -14850 69020 -14650 69090
rect -14350 69020 -14150 69090
rect -13850 69020 -13650 69090
rect -13350 69020 -13150 69090
rect -12850 69020 -12650 69090
rect -12350 69020 -12150 69090
rect -15850 68910 -15650 68980
rect -15350 68910 -15150 68980
rect -14850 68910 -14650 68980
rect -14350 68910 -14150 68980
rect -13850 68910 -13650 68980
rect -13350 68910 -13150 68980
rect -12850 68910 -12650 68980
rect -12350 68910 -12150 68980
rect -15980 68650 -15910 68850
rect -15590 68650 -15520 68850
rect -15480 68650 -15410 68850
rect -15090 68650 -15020 68850
rect -14980 68650 -14910 68850
rect -14590 68650 -14520 68850
rect -14480 68650 -14410 68850
rect -14090 68650 -14020 68850
rect -13980 68650 -13910 68850
rect -13590 68650 -13520 68850
rect -13480 68650 -13410 68850
rect -13090 68650 -13020 68850
rect -12980 68650 -12910 68850
rect -12590 68650 -12520 68850
rect -12480 68650 -12410 68850
rect -12090 68650 -12020 68850
rect -15850 68520 -15650 68590
rect -15350 68520 -15150 68590
rect -14850 68520 -14650 68590
rect -14350 68520 -14150 68590
rect -13850 68520 -13650 68590
rect -13350 68520 -13150 68590
rect -12850 68520 -12650 68590
rect -12350 68520 -12150 68590
rect -15850 68410 -15650 68480
rect -15350 68410 -15150 68480
rect -14850 68410 -14650 68480
rect -14350 68410 -14150 68480
rect -13850 68410 -13650 68480
rect -13350 68410 -13150 68480
rect -12850 68410 -12650 68480
rect -12350 68410 -12150 68480
rect -15980 68150 -15910 68350
rect -15590 68150 -15520 68350
rect -15480 68150 -15410 68350
rect -15090 68150 -15020 68350
rect -14980 68150 -14910 68350
rect -14590 68150 -14520 68350
rect -14480 68150 -14410 68350
rect -14090 68150 -14020 68350
rect -13980 68150 -13910 68350
rect -13590 68150 -13520 68350
rect -13480 68150 -13410 68350
rect -13090 68150 -13020 68350
rect -12980 68150 -12910 68350
rect -12590 68150 -12520 68350
rect -12480 68150 -12410 68350
rect -12090 68150 -12020 68350
rect -15850 68020 -15650 68090
rect -15350 68020 -15150 68090
rect -14850 68020 -14650 68090
rect -14350 68020 -14150 68090
rect -13850 68020 -13650 68090
rect -13350 68020 -13150 68090
rect -12850 68020 -12650 68090
rect -12350 68020 -12150 68090
rect -15850 67910 -15650 67980
rect -15350 67910 -15150 67980
rect -14850 67910 -14650 67980
rect -14350 67910 -14150 67980
rect -13850 67910 -13650 67980
rect -13350 67910 -13150 67980
rect -12850 67910 -12650 67980
rect -12350 67910 -12150 67980
rect -15980 67650 -15910 67850
rect -15590 67650 -15520 67850
rect -15480 67650 -15410 67850
rect -15090 67650 -15020 67850
rect -14980 67650 -14910 67850
rect -14590 67650 -14520 67850
rect -14480 67650 -14410 67850
rect -14090 67650 -14020 67850
rect -13980 67650 -13910 67850
rect -13590 67650 -13520 67850
rect -13480 67650 -13410 67850
rect -13090 67650 -13020 67850
rect -12980 67650 -12910 67850
rect -12590 67650 -12520 67850
rect -12480 67650 -12410 67850
rect -12090 67650 -12020 67850
rect -15850 67520 -15650 67590
rect -15350 67520 -15150 67590
rect -14850 67520 -14650 67590
rect -14350 67520 -14150 67590
rect -13850 67520 -13650 67590
rect -13350 67520 -13150 67590
rect -12850 67520 -12650 67590
rect -12350 67520 -12150 67590
rect -15850 67410 -15650 67480
rect -15350 67410 -15150 67480
rect -14850 67410 -14650 67480
rect -14350 67410 -14150 67480
rect -13850 67410 -13650 67480
rect -13350 67410 -13150 67480
rect -12850 67410 -12650 67480
rect -12350 67410 -12150 67480
rect -15980 67150 -15910 67350
rect -15590 67150 -15520 67350
rect -15480 67150 -15410 67350
rect -15090 67150 -15020 67350
rect -14980 67150 -14910 67350
rect -14590 67150 -14520 67350
rect -14480 67150 -14410 67350
rect -14090 67150 -14020 67350
rect -13980 67150 -13910 67350
rect -13590 67150 -13520 67350
rect -13480 67150 -13410 67350
rect -13090 67150 -13020 67350
rect -12980 67150 -12910 67350
rect -12590 67150 -12520 67350
rect -12480 67150 -12410 67350
rect -12090 67150 -12020 67350
rect -15850 67020 -15650 67090
rect -15350 67020 -15150 67090
rect -14850 67020 -14650 67090
rect -14350 67020 -14150 67090
rect -13850 67020 -13650 67090
rect -13350 67020 -13150 67090
rect -12850 67020 -12650 67090
rect -12350 67020 -12150 67090
rect -15850 66910 -15650 66980
rect -15350 66910 -15150 66980
rect -14850 66910 -14650 66980
rect -14350 66910 -14150 66980
rect -13850 66910 -13650 66980
rect -13350 66910 -13150 66980
rect -12850 66910 -12650 66980
rect -12350 66910 -12150 66980
rect -15980 66650 -15910 66850
rect -15590 66650 -15520 66850
rect -15480 66650 -15410 66850
rect -15090 66650 -15020 66850
rect -14980 66650 -14910 66850
rect -14590 66650 -14520 66850
rect -14480 66650 -14410 66850
rect -14090 66650 -14020 66850
rect -13980 66650 -13910 66850
rect -13590 66650 -13520 66850
rect -13480 66650 -13410 66850
rect -13090 66650 -13020 66850
rect -12980 66650 -12910 66850
rect -12590 66650 -12520 66850
rect -12480 66650 -12410 66850
rect -12090 66650 -12020 66850
rect -15850 66520 -15650 66590
rect -15350 66520 -15150 66590
rect -14850 66520 -14650 66590
rect -14350 66520 -14150 66590
rect -13850 66520 -13650 66590
rect -13350 66520 -13150 66590
rect -12850 66520 -12650 66590
rect -12350 66520 -12150 66590
rect -15850 66410 -15650 66480
rect -15350 66410 -15150 66480
rect -14850 66410 -14650 66480
rect -14350 66410 -14150 66480
rect -13850 66410 -13650 66480
rect -13350 66410 -13150 66480
rect -12850 66410 -12650 66480
rect -12350 66410 -12150 66480
rect -15980 66150 -15910 66350
rect -15590 66150 -15520 66350
rect -15480 66150 -15410 66350
rect -15090 66150 -15020 66350
rect -14980 66150 -14910 66350
rect -14590 66150 -14520 66350
rect -14480 66150 -14410 66350
rect -14090 66150 -14020 66350
rect -13980 66150 -13910 66350
rect -13590 66150 -13520 66350
rect -13480 66150 -13410 66350
rect -13090 66150 -13020 66350
rect -12980 66150 -12910 66350
rect -12590 66150 -12520 66350
rect -12480 66150 -12410 66350
rect -12090 66150 -12020 66350
rect -15850 66020 -15650 66090
rect -15350 66020 -15150 66090
rect -14850 66020 -14650 66090
rect -14350 66020 -14150 66090
rect -13850 66020 -13650 66090
rect -13350 66020 -13150 66090
rect -12850 66020 -12650 66090
rect -12350 66020 -12150 66090
rect -15850 65910 -15650 65980
rect -15350 65910 -15150 65980
rect -14850 65910 -14650 65980
rect -14350 65910 -14150 65980
rect -13850 65910 -13650 65980
rect -13350 65910 -13150 65980
rect -12850 65910 -12650 65980
rect -12350 65910 -12150 65980
rect -15980 65650 -15910 65850
rect -15590 65650 -15520 65850
rect -15480 65650 -15410 65850
rect -15090 65650 -15020 65850
rect -14980 65650 -14910 65850
rect -14590 65650 -14520 65850
rect -14480 65650 -14410 65850
rect -14090 65650 -14020 65850
rect -13980 65650 -13910 65850
rect -13590 65650 -13520 65850
rect -13480 65650 -13410 65850
rect -13090 65650 -13020 65850
rect -12980 65650 -12910 65850
rect -12590 65650 -12520 65850
rect -12480 65650 -12410 65850
rect -12090 65650 -12020 65850
rect -15850 65520 -15650 65590
rect -15350 65520 -15150 65590
rect -14850 65520 -14650 65590
rect -14350 65520 -14150 65590
rect -13850 65520 -13650 65590
rect -13350 65520 -13150 65590
rect -12850 65520 -12650 65590
rect -12350 65520 -12150 65590
rect -15850 65410 -15650 65480
rect -15350 65410 -15150 65480
rect -14850 65410 -14650 65480
rect -14350 65410 -14150 65480
rect -13850 65410 -13650 65480
rect -13350 65410 -13150 65480
rect -12850 65410 -12650 65480
rect -12350 65410 -12150 65480
rect -15980 65150 -15910 65350
rect -15590 65150 -15520 65350
rect -15480 65150 -15410 65350
rect -15090 65150 -15020 65350
rect -14980 65150 -14910 65350
rect -14590 65150 -14520 65350
rect -14480 65150 -14410 65350
rect -14090 65150 -14020 65350
rect -13980 65150 -13910 65350
rect -13590 65150 -13520 65350
rect -13480 65150 -13410 65350
rect -13090 65150 -13020 65350
rect -12980 65150 -12910 65350
rect -12590 65150 -12520 65350
rect -12480 65150 -12410 65350
rect -12090 65150 -12020 65350
rect -15850 65020 -15650 65090
rect -15350 65020 -15150 65090
rect -14850 65020 -14650 65090
rect -14350 65020 -14150 65090
rect -13850 65020 -13650 65090
rect -13350 65020 -13150 65090
rect -12850 65020 -12650 65090
rect -12350 65020 -12150 65090
rect -15850 64910 -15650 64980
rect -15350 64910 -15150 64980
rect -14850 64910 -14650 64980
rect -14350 64910 -14150 64980
rect -13850 64910 -13650 64980
rect -13350 64910 -13150 64980
rect -12850 64910 -12650 64980
rect -12350 64910 -12150 64980
rect -15980 64650 -15910 64850
rect -15590 64650 -15520 64850
rect -15480 64650 -15410 64850
rect -15090 64650 -15020 64850
rect -14980 64650 -14910 64850
rect -14590 64650 -14520 64850
rect -14480 64650 -14410 64850
rect -14090 64650 -14020 64850
rect -13980 64650 -13910 64850
rect -13590 64650 -13520 64850
rect -13480 64650 -13410 64850
rect -13090 64650 -13020 64850
rect -12980 64650 -12910 64850
rect -12590 64650 -12520 64850
rect -12480 64650 -12410 64850
rect -12090 64650 -12020 64850
rect -15850 64520 -15650 64590
rect -15350 64520 -15150 64590
rect -14850 64520 -14650 64590
rect -14350 64520 -14150 64590
rect -13850 64520 -13650 64590
rect -13350 64520 -13150 64590
rect -12850 64520 -12650 64590
rect -12350 64520 -12150 64590
rect -15850 64410 -15650 64480
rect -15350 64410 -15150 64480
rect -14850 64410 -14650 64480
rect -14350 64410 -14150 64480
rect -13850 64410 -13650 64480
rect -13350 64410 -13150 64480
rect -12850 64410 -12650 64480
rect -12350 64410 -12150 64480
rect -15980 64150 -15910 64350
rect -15590 64150 -15520 64350
rect -15480 64150 -15410 64350
rect -15090 64150 -15020 64350
rect -14980 64150 -14910 64350
rect -14590 64150 -14520 64350
rect -14480 64150 -14410 64350
rect -14090 64150 -14020 64350
rect -13980 64150 -13910 64350
rect -13590 64150 -13520 64350
rect -13480 64150 -13410 64350
rect -13090 64150 -13020 64350
rect -12980 64150 -12910 64350
rect -12590 64150 -12520 64350
rect -12480 64150 -12410 64350
rect -12090 64150 -12020 64350
rect -15850 64020 -15650 64090
rect -15350 64020 -15150 64090
rect -14850 64020 -14650 64090
rect -14350 64020 -14150 64090
rect -13850 64020 -13650 64090
rect -13350 64020 -13150 64090
rect -12850 64020 -12650 64090
rect -12350 64020 -12150 64090
rect -15850 63910 -15650 63980
rect -15350 63910 -15150 63980
rect -14850 63910 -14650 63980
rect -14350 63910 -14150 63980
rect -13850 63910 -13650 63980
rect -13350 63910 -13150 63980
rect -12850 63910 -12650 63980
rect -12350 63910 -12150 63980
rect -15980 63650 -15910 63850
rect -15590 63650 -15520 63850
rect -15480 63650 -15410 63850
rect -15090 63650 -15020 63850
rect -14980 63650 -14910 63850
rect -14590 63650 -14520 63850
rect -14480 63650 -14410 63850
rect -14090 63650 -14020 63850
rect -13980 63650 -13910 63850
rect -13590 63650 -13520 63850
rect -13480 63650 -13410 63850
rect -13090 63650 -13020 63850
rect -12980 63650 -12910 63850
rect -12590 63650 -12520 63850
rect -12480 63650 -12410 63850
rect -12090 63650 -12020 63850
rect -15850 63520 -15650 63590
rect -15350 63520 -15150 63590
rect -14850 63520 -14650 63590
rect -14350 63520 -14150 63590
rect -13850 63520 -13650 63590
rect -13350 63520 -13150 63590
rect -12850 63520 -12650 63590
rect -12350 63520 -12150 63590
rect -15850 63410 -15650 63480
rect -15350 63410 -15150 63480
rect -14850 63410 -14650 63480
rect -14350 63410 -14150 63480
rect -13850 63410 -13650 63480
rect -13350 63410 -13150 63480
rect -12850 63410 -12650 63480
rect -12350 63410 -12150 63480
rect -15980 63150 -15910 63350
rect -15590 63150 -15520 63350
rect -15480 63150 -15410 63350
rect -15090 63150 -15020 63350
rect -14980 63150 -14910 63350
rect -14590 63150 -14520 63350
rect -14480 63150 -14410 63350
rect -14090 63150 -14020 63350
rect -13980 63150 -13910 63350
rect -13590 63150 -13520 63350
rect -13480 63150 -13410 63350
rect -13090 63150 -13020 63350
rect -12980 63150 -12910 63350
rect -12590 63150 -12520 63350
rect -12480 63150 -12410 63350
rect -12090 63150 -12020 63350
rect -15850 63020 -15650 63090
rect -15350 63020 -15150 63090
rect -14850 63020 -14650 63090
rect -14350 63020 -14150 63090
rect -13850 63020 -13650 63090
rect -13350 63020 -13150 63090
rect -12850 63020 -12650 63090
rect -12350 63020 -12150 63090
rect -15850 62910 -15650 62980
rect -15350 62910 -15150 62980
rect -14850 62910 -14650 62980
rect -14350 62910 -14150 62980
rect -13850 62910 -13650 62980
rect -13350 62910 -13150 62980
rect -12850 62910 -12650 62980
rect -12350 62910 -12150 62980
rect -15980 62650 -15910 62850
rect -15590 62650 -15520 62850
rect -15480 62650 -15410 62850
rect -15090 62650 -15020 62850
rect -14980 62650 -14910 62850
rect -14590 62650 -14520 62850
rect -14480 62650 -14410 62850
rect -14090 62650 -14020 62850
rect -13980 62650 -13910 62850
rect -13590 62650 -13520 62850
rect -13480 62650 -13410 62850
rect -13090 62650 -13020 62850
rect -12980 62650 -12910 62850
rect -12590 62650 -12520 62850
rect -12480 62650 -12410 62850
rect -12090 62650 -12020 62850
rect -15850 62520 -15650 62590
rect -15350 62520 -15150 62590
rect -14850 62520 -14650 62590
rect -14350 62520 -14150 62590
rect -13850 62520 -13650 62590
rect -13350 62520 -13150 62590
rect -12850 62520 -12650 62590
rect -12350 62520 -12150 62590
rect -15850 62410 -15650 62480
rect -15350 62410 -15150 62480
rect -14850 62410 -14650 62480
rect -14350 62410 -14150 62480
rect -13850 62410 -13650 62480
rect -13350 62410 -13150 62480
rect -12850 62410 -12650 62480
rect -12350 62410 -12150 62480
rect -15980 62150 -15910 62350
rect -15590 62150 -15520 62350
rect -15480 62150 -15410 62350
rect -15090 62150 -15020 62350
rect -14980 62150 -14910 62350
rect -14590 62150 -14520 62350
rect -14480 62150 -14410 62350
rect -14090 62150 -14020 62350
rect -13980 62150 -13910 62350
rect -13590 62150 -13520 62350
rect -13480 62150 -13410 62350
rect -13090 62150 -13020 62350
rect -12980 62150 -12910 62350
rect -12590 62150 -12520 62350
rect -12480 62150 -12410 62350
rect -12090 62150 -12020 62350
rect -15850 62020 -15650 62090
rect -15350 62020 -15150 62090
rect -14850 62020 -14650 62090
rect -14350 62020 -14150 62090
rect -13850 62020 -13650 62090
rect -13350 62020 -13150 62090
rect -12850 62020 -12650 62090
rect -12350 62020 -12150 62090
rect -15850 61910 -15650 61980
rect -15350 61910 -15150 61980
rect -14850 61910 -14650 61980
rect -14350 61910 -14150 61980
rect -13850 61910 -13650 61980
rect -13350 61910 -13150 61980
rect -12850 61910 -12650 61980
rect -12350 61910 -12150 61980
rect -15980 61650 -15910 61850
rect -15590 61650 -15520 61850
rect -15480 61650 -15410 61850
rect -15090 61650 -15020 61850
rect -14980 61650 -14910 61850
rect -14590 61650 -14520 61850
rect -14480 61650 -14410 61850
rect -14090 61650 -14020 61850
rect -13980 61650 -13910 61850
rect -13590 61650 -13520 61850
rect -13480 61650 -13410 61850
rect -13090 61650 -13020 61850
rect -12980 61650 -12910 61850
rect -12590 61650 -12520 61850
rect -12480 61650 -12410 61850
rect -12090 61650 -12020 61850
rect -15850 61520 -15650 61590
rect -15350 61520 -15150 61590
rect -14850 61520 -14650 61590
rect -14350 61520 -14150 61590
rect -13850 61520 -13650 61590
rect -13350 61520 -13150 61590
rect -12850 61520 -12650 61590
rect -12350 61520 -12150 61590
rect -15850 61410 -15650 61480
rect -15350 61410 -15150 61480
rect -14850 61410 -14650 61480
rect -14350 61410 -14150 61480
rect -13850 61410 -13650 61480
rect -13350 61410 -13150 61480
rect -12850 61410 -12650 61480
rect -12350 61410 -12150 61480
rect -15980 61150 -15910 61350
rect -15590 61150 -15520 61350
rect -15480 61150 -15410 61350
rect -15090 61150 -15020 61350
rect -14980 61150 -14910 61350
rect -14590 61150 -14520 61350
rect -14480 61150 -14410 61350
rect -14090 61150 -14020 61350
rect -13980 61150 -13910 61350
rect -13590 61150 -13520 61350
rect -13480 61150 -13410 61350
rect -13090 61150 -13020 61350
rect -12980 61150 -12910 61350
rect -12590 61150 -12520 61350
rect -12480 61150 -12410 61350
rect -12090 61150 -12020 61350
rect -15850 61020 -15650 61090
rect -15350 61020 -15150 61090
rect -14850 61020 -14650 61090
rect -14350 61020 -14150 61090
rect -13850 61020 -13650 61090
rect -13350 61020 -13150 61090
rect -12850 61020 -12650 61090
rect -12350 61020 -12150 61090
rect -15850 60910 -15650 60980
rect -15350 60910 -15150 60980
rect -14850 60910 -14650 60980
rect -14350 60910 -14150 60980
rect -13850 60910 -13650 60980
rect -13350 60910 -13150 60980
rect -12850 60910 -12650 60980
rect -12350 60910 -12150 60980
rect -15980 60650 -15910 60850
rect -15590 60650 -15520 60850
rect -15480 60650 -15410 60850
rect -15090 60650 -15020 60850
rect -14980 60650 -14910 60850
rect -14590 60650 -14520 60850
rect -14480 60650 -14410 60850
rect -14090 60650 -14020 60850
rect -13980 60650 -13910 60850
rect -13590 60650 -13520 60850
rect -13480 60650 -13410 60850
rect -13090 60650 -13020 60850
rect -12980 60650 -12910 60850
rect -12590 60650 -12520 60850
rect -12480 60650 -12410 60850
rect -12090 60650 -12020 60850
rect -15850 60520 -15650 60590
rect -15350 60520 -15150 60590
rect -14850 60520 -14650 60590
rect -14350 60520 -14150 60590
rect -13850 60520 -13650 60590
rect -13350 60520 -13150 60590
rect -12850 60520 -12650 60590
rect -12350 60520 -12150 60590
rect -15850 60410 -15650 60480
rect -15350 60410 -15150 60480
rect -14850 60410 -14650 60480
rect -14350 60410 -14150 60480
rect -13850 60410 -13650 60480
rect -13350 60410 -13150 60480
rect -12850 60410 -12650 60480
rect -12350 60410 -12150 60480
rect -15980 60150 -15910 60350
rect -15590 60150 -15520 60350
rect -15480 60150 -15410 60350
rect -15090 60150 -15020 60350
rect -14980 60150 -14910 60350
rect -14590 60150 -14520 60350
rect -14480 60150 -14410 60350
rect -14090 60150 -14020 60350
rect -13980 60150 -13910 60350
rect -13590 60150 -13520 60350
rect -13480 60150 -13410 60350
rect -13090 60150 -13020 60350
rect -12980 60150 -12910 60350
rect -12590 60150 -12520 60350
rect -12480 60150 -12410 60350
rect -12090 60150 -12020 60350
rect -15850 60020 -15650 60090
rect -15350 60020 -15150 60090
rect -14850 60020 -14650 60090
rect -14350 60020 -14150 60090
rect -13850 60020 -13650 60090
rect -13350 60020 -13150 60090
rect -12850 60020 -12650 60090
rect -12350 60020 -12150 60090
rect -15850 59910 -15650 59980
rect -15350 59910 -15150 59980
rect -14850 59910 -14650 59980
rect -14350 59910 -14150 59980
rect -13850 59910 -13650 59980
rect -13350 59910 -13150 59980
rect -12850 59910 -12650 59980
rect -12350 59910 -12150 59980
rect -15980 59650 -15910 59850
rect -15590 59650 -15520 59850
rect -15480 59650 -15410 59850
rect -15090 59650 -15020 59850
rect -14980 59650 -14910 59850
rect -14590 59650 -14520 59850
rect -14480 59650 -14410 59850
rect -14090 59650 -14020 59850
rect -13980 59650 -13910 59850
rect -13590 59650 -13520 59850
rect -13480 59650 -13410 59850
rect -13090 59650 -13020 59850
rect -12980 59650 -12910 59850
rect -12590 59650 -12520 59850
rect -12480 59650 -12410 59850
rect -12090 59650 -12020 59850
rect -15850 59520 -15650 59590
rect -15350 59520 -15150 59590
rect -14850 59520 -14650 59590
rect -14350 59520 -14150 59590
rect -13850 59520 -13650 59590
rect -13350 59520 -13150 59590
rect -12850 59520 -12650 59590
rect -12350 59520 -12150 59590
rect -15850 59410 -15650 59480
rect -15350 59410 -15150 59480
rect -14850 59410 -14650 59480
rect -14350 59410 -14150 59480
rect -13850 59410 -13650 59480
rect -13350 59410 -13150 59480
rect -12850 59410 -12650 59480
rect -12350 59410 -12150 59480
rect -15980 59150 -15910 59350
rect -15590 59150 -15520 59350
rect -15480 59150 -15410 59350
rect -15090 59150 -15020 59350
rect -14980 59150 -14910 59350
rect -14590 59150 -14520 59350
rect -14480 59150 -14410 59350
rect -14090 59150 -14020 59350
rect -13980 59150 -13910 59350
rect -13590 59150 -13520 59350
rect -13480 59150 -13410 59350
rect -13090 59150 -13020 59350
rect -12980 59150 -12910 59350
rect -12590 59150 -12520 59350
rect -12480 59150 -12410 59350
rect -12090 59150 -12020 59350
rect -15850 59020 -15650 59090
rect -15350 59020 -15150 59090
rect -14850 59020 -14650 59090
rect -14350 59020 -14150 59090
rect -13850 59020 -13650 59090
rect -13350 59020 -13150 59090
rect -12850 59020 -12650 59090
rect -12350 59020 -12150 59090
rect -15850 58910 -15650 58980
rect -15350 58910 -15150 58980
rect -14850 58910 -14650 58980
rect -14350 58910 -14150 58980
rect -13850 58910 -13650 58980
rect -13350 58910 -13150 58980
rect -12850 58910 -12650 58980
rect -12350 58910 -12150 58980
rect -15980 58650 -15910 58850
rect -15590 58650 -15520 58850
rect -15480 58650 -15410 58850
rect -15090 58650 -15020 58850
rect -14980 58650 -14910 58850
rect -14590 58650 -14520 58850
rect -14480 58650 -14410 58850
rect -14090 58650 -14020 58850
rect -13980 58650 -13910 58850
rect -13590 58650 -13520 58850
rect -13480 58650 -13410 58850
rect -13090 58650 -13020 58850
rect -12980 58650 -12910 58850
rect -12590 58650 -12520 58850
rect -12480 58650 -12410 58850
rect -12090 58650 -12020 58850
rect -15850 58520 -15650 58590
rect -15350 58520 -15150 58590
rect -14850 58520 -14650 58590
rect -14350 58520 -14150 58590
rect -13850 58520 -13650 58590
rect -13350 58520 -13150 58590
rect -12850 58520 -12650 58590
rect -12350 58520 -12150 58590
rect -15850 58410 -15650 58480
rect -15350 58410 -15150 58480
rect -14850 58410 -14650 58480
rect -14350 58410 -14150 58480
rect -13850 58410 -13650 58480
rect -13350 58410 -13150 58480
rect -12850 58410 -12650 58480
rect -12350 58410 -12150 58480
rect -15980 58150 -15910 58350
rect -15590 58150 -15520 58350
rect -15480 58150 -15410 58350
rect -15090 58150 -15020 58350
rect -14980 58150 -14910 58350
rect -14590 58150 -14520 58350
rect -14480 58150 -14410 58350
rect -14090 58150 -14020 58350
rect -13980 58150 -13910 58350
rect -13590 58150 -13520 58350
rect -13480 58150 -13410 58350
rect -13090 58150 -13020 58350
rect -12980 58150 -12910 58350
rect -12590 58150 -12520 58350
rect -12480 58150 -12410 58350
rect -12090 58150 -12020 58350
rect -15850 58020 -15650 58090
rect -15350 58020 -15150 58090
rect -14850 58020 -14650 58090
rect -14350 58020 -14150 58090
rect -13850 58020 -13650 58090
rect -13350 58020 -13150 58090
rect -12850 58020 -12650 58090
rect -12350 58020 -12150 58090
rect -15850 57910 -15650 57980
rect -15350 57910 -15150 57980
rect -14850 57910 -14650 57980
rect -14350 57910 -14150 57980
rect -13850 57910 -13650 57980
rect -13350 57910 -13150 57980
rect -12850 57910 -12650 57980
rect -12350 57910 -12150 57980
rect -15980 57650 -15910 57850
rect -15590 57650 -15520 57850
rect -15480 57650 -15410 57850
rect -15090 57650 -15020 57850
rect -14980 57650 -14910 57850
rect -14590 57650 -14520 57850
rect -14480 57650 -14410 57850
rect -14090 57650 -14020 57850
rect -13980 57650 -13910 57850
rect -13590 57650 -13520 57850
rect -13480 57650 -13410 57850
rect -13090 57650 -13020 57850
rect -12980 57650 -12910 57850
rect -12590 57650 -12520 57850
rect -12480 57650 -12410 57850
rect -12090 57650 -12020 57850
rect -15850 57520 -15650 57590
rect -15350 57520 -15150 57590
rect -14850 57520 -14650 57590
rect -14350 57520 -14150 57590
rect -13850 57520 -13650 57590
rect -13350 57520 -13150 57590
rect -12850 57520 -12650 57590
rect -12350 57520 -12150 57590
rect -15850 57410 -15650 57480
rect -15350 57410 -15150 57480
rect -14850 57410 -14650 57480
rect -14350 57410 -14150 57480
rect -13850 57410 -13650 57480
rect -13350 57410 -13150 57480
rect -12850 57410 -12650 57480
rect -12350 57410 -12150 57480
rect -15980 57150 -15910 57350
rect -15590 57150 -15520 57350
rect -15480 57150 -15410 57350
rect -15090 57150 -15020 57350
rect -14980 57150 -14910 57350
rect -14590 57150 -14520 57350
rect -14480 57150 -14410 57350
rect -14090 57150 -14020 57350
rect -13980 57150 -13910 57350
rect -13590 57150 -13520 57350
rect -13480 57150 -13410 57350
rect -13090 57150 -13020 57350
rect -12980 57150 -12910 57350
rect -12590 57150 -12520 57350
rect -12480 57150 -12410 57350
rect -12090 57150 -12020 57350
rect -15850 57020 -15650 57090
rect -15350 57020 -15150 57090
rect -14850 57020 -14650 57090
rect -14350 57020 -14150 57090
rect -13850 57020 -13650 57090
rect -13350 57020 -13150 57090
rect -12850 57020 -12650 57090
rect -12350 57020 -12150 57090
rect -15850 56910 -15650 56980
rect -15350 56910 -15150 56980
rect -14850 56910 -14650 56980
rect -14350 56910 -14150 56980
rect -13850 56910 -13650 56980
rect -13350 56910 -13150 56980
rect -12850 56910 -12650 56980
rect -12350 56910 -12150 56980
rect -15980 56650 -15910 56850
rect -15590 56650 -15520 56850
rect -15480 56650 -15410 56850
rect -15090 56650 -15020 56850
rect -14980 56650 -14910 56850
rect -14590 56650 -14520 56850
rect -14480 56650 -14410 56850
rect -14090 56650 -14020 56850
rect -13980 56650 -13910 56850
rect -13590 56650 -13520 56850
rect -13480 56650 -13410 56850
rect -13090 56650 -13020 56850
rect -12980 56650 -12910 56850
rect -12590 56650 -12520 56850
rect -12480 56650 -12410 56850
rect -12090 56650 -12020 56850
rect -15850 56520 -15650 56590
rect -15350 56520 -15150 56590
rect -14850 56520 -14650 56590
rect -14350 56520 -14150 56590
rect -13850 56520 -13650 56590
rect -13350 56520 -13150 56590
rect -12850 56520 -12650 56590
rect -12350 56520 -12150 56590
rect -15850 56410 -15650 56480
rect -15350 56410 -15150 56480
rect -14850 56410 -14650 56480
rect -14350 56410 -14150 56480
rect -13850 56410 -13650 56480
rect -13350 56410 -13150 56480
rect -12850 56410 -12650 56480
rect -12350 56410 -12150 56480
rect -15980 56150 -15910 56350
rect -15590 56150 -15520 56350
rect -15480 56150 -15410 56350
rect -15090 56150 -15020 56350
rect -14980 56150 -14910 56350
rect -14590 56150 -14520 56350
rect -14480 56150 -14410 56350
rect -14090 56150 -14020 56350
rect -13980 56150 -13910 56350
rect -13590 56150 -13520 56350
rect -13480 56150 -13410 56350
rect -13090 56150 -13020 56350
rect -12980 56150 -12910 56350
rect -12590 56150 -12520 56350
rect -12480 56150 -12410 56350
rect -12090 56150 -12020 56350
rect -15850 56020 -15650 56090
rect -15350 56020 -15150 56090
rect -14850 56020 -14650 56090
rect -14350 56020 -14150 56090
rect -13850 56020 -13650 56090
rect -13350 56020 -13150 56090
rect -12850 56020 -12650 56090
rect -12350 56020 -12150 56090
rect -15850 55910 -15650 55980
rect -15350 55910 -15150 55980
rect -14850 55910 -14650 55980
rect -14350 55910 -14150 55980
rect -13850 55910 -13650 55980
rect -13350 55910 -13150 55980
rect -12850 55910 -12650 55980
rect -12350 55910 -12150 55980
rect -15980 55650 -15910 55850
rect -15590 55650 -15520 55850
rect -15480 55650 -15410 55850
rect -15090 55650 -15020 55850
rect -14980 55650 -14910 55850
rect -14590 55650 -14520 55850
rect -14480 55650 -14410 55850
rect -14090 55650 -14020 55850
rect -13980 55650 -13910 55850
rect -13590 55650 -13520 55850
rect -13480 55650 -13410 55850
rect -13090 55650 -13020 55850
rect -12980 55650 -12910 55850
rect -12590 55650 -12520 55850
rect -12480 55650 -12410 55850
rect -12090 55650 -12020 55850
rect -15850 55520 -15650 55590
rect -15350 55520 -15150 55590
rect -14850 55520 -14650 55590
rect -14350 55520 -14150 55590
rect -13850 55520 -13650 55590
rect -13350 55520 -13150 55590
rect -12850 55520 -12650 55590
rect -12350 55520 -12150 55590
rect -15850 55410 -15650 55480
rect -15350 55410 -15150 55480
rect -14850 55410 -14650 55480
rect -14350 55410 -14150 55480
rect -13850 55410 -13650 55480
rect -13350 55410 -13150 55480
rect -12850 55410 -12650 55480
rect -12350 55410 -12150 55480
rect -15980 55150 -15910 55350
rect -15590 55150 -15520 55350
rect -15480 55150 -15410 55350
rect -15090 55150 -15020 55350
rect -14980 55150 -14910 55350
rect -14590 55150 -14520 55350
rect -14480 55150 -14410 55350
rect -14090 55150 -14020 55350
rect -13980 55150 -13910 55350
rect -13590 55150 -13520 55350
rect -13480 55150 -13410 55350
rect -13090 55150 -13020 55350
rect -12980 55150 -12910 55350
rect -12590 55150 -12520 55350
rect -12480 55150 -12410 55350
rect -12090 55150 -12020 55350
rect -15850 55020 -15650 55090
rect -15350 55020 -15150 55090
rect -14850 55020 -14650 55090
rect -14350 55020 -14150 55090
rect -13850 55020 -13650 55090
rect -13350 55020 -13150 55090
rect -12850 55020 -12650 55090
rect -12350 55020 -12150 55090
rect -15850 54910 -15650 54980
rect -15350 54910 -15150 54980
rect -14850 54910 -14650 54980
rect -14350 54910 -14150 54980
rect -13850 54910 -13650 54980
rect -13350 54910 -13150 54980
rect -12850 54910 -12650 54980
rect -12350 54910 -12150 54980
rect -15980 54650 -15910 54850
rect -15590 54650 -15520 54850
rect -15480 54650 -15410 54850
rect -15090 54650 -15020 54850
rect -14980 54650 -14910 54850
rect -14590 54650 -14520 54850
rect -14480 54650 -14410 54850
rect -14090 54650 -14020 54850
rect -13980 54650 -13910 54850
rect -13590 54650 -13520 54850
rect -13480 54650 -13410 54850
rect -13090 54650 -13020 54850
rect -12980 54650 -12910 54850
rect -12590 54650 -12520 54850
rect -12480 54650 -12410 54850
rect -12090 54650 -12020 54850
rect -15850 54520 -15650 54590
rect -15350 54520 -15150 54590
rect -14850 54520 -14650 54590
rect -14350 54520 -14150 54590
rect -13850 54520 -13650 54590
rect -13350 54520 -13150 54590
rect -12850 54520 -12650 54590
rect -12350 54520 -12150 54590
rect -15850 54410 -15650 54480
rect -15350 54410 -15150 54480
rect -14850 54410 -14650 54480
rect -14350 54410 -14150 54480
rect -13850 54410 -13650 54480
rect -13350 54410 -13150 54480
rect -12850 54410 -12650 54480
rect -12350 54410 -12150 54480
rect -15980 54150 -15910 54350
rect -15590 54150 -15520 54350
rect -15480 54150 -15410 54350
rect -15090 54150 -15020 54350
rect -14980 54150 -14910 54350
rect -14590 54150 -14520 54350
rect -14480 54150 -14410 54350
rect -14090 54150 -14020 54350
rect -13980 54150 -13910 54350
rect -13590 54150 -13520 54350
rect -13480 54150 -13410 54350
rect -13090 54150 -13020 54350
rect -12980 54150 -12910 54350
rect -12590 54150 -12520 54350
rect -12480 54150 -12410 54350
rect -12090 54150 -12020 54350
rect -15850 54020 -15650 54090
rect -15350 54020 -15150 54090
rect -14850 54020 -14650 54090
rect -14350 54020 -14150 54090
rect -13850 54020 -13650 54090
rect -13350 54020 -13150 54090
rect -12850 54020 -12650 54090
rect -12350 54020 -12150 54090
rect -15850 53910 -15650 53980
rect -15350 53910 -15150 53980
rect -14850 53910 -14650 53980
rect -14350 53910 -14150 53980
rect -13850 53910 -13650 53980
rect -13350 53910 -13150 53980
rect -12850 53910 -12650 53980
rect -12350 53910 -12150 53980
rect -15980 53650 -15910 53850
rect -15590 53650 -15520 53850
rect -15480 53650 -15410 53850
rect -15090 53650 -15020 53850
rect -14980 53650 -14910 53850
rect -14590 53650 -14520 53850
rect -14480 53650 -14410 53850
rect -14090 53650 -14020 53850
rect -13980 53650 -13910 53850
rect -13590 53650 -13520 53850
rect -13480 53650 -13410 53850
rect -13090 53650 -13020 53850
rect -12980 53650 -12910 53850
rect -12590 53650 -12520 53850
rect -12480 53650 -12410 53850
rect -12090 53650 -12020 53850
rect -15850 53520 -15650 53590
rect -15350 53520 -15150 53590
rect -14850 53520 -14650 53590
rect -14350 53520 -14150 53590
rect -13850 53520 -13650 53590
rect -13350 53520 -13150 53590
rect -12850 53520 -12650 53590
rect -12350 53520 -12150 53590
rect -15850 53410 -15650 53480
rect -15350 53410 -15150 53480
rect -14850 53410 -14650 53480
rect -14350 53410 -14150 53480
rect -13850 53410 -13650 53480
rect -13350 53410 -13150 53480
rect -12850 53410 -12650 53480
rect -12350 53410 -12150 53480
rect -15980 53150 -15910 53350
rect -15590 53150 -15520 53350
rect -15480 53150 -15410 53350
rect -15090 53150 -15020 53350
rect -14980 53150 -14910 53350
rect -14590 53150 -14520 53350
rect -14480 53150 -14410 53350
rect -14090 53150 -14020 53350
rect -13980 53150 -13910 53350
rect -13590 53150 -13520 53350
rect -13480 53150 -13410 53350
rect -13090 53150 -13020 53350
rect -12980 53150 -12910 53350
rect -12590 53150 -12520 53350
rect -12480 53150 -12410 53350
rect -12090 53150 -12020 53350
rect -15850 53020 -15650 53090
rect -15350 53020 -15150 53090
rect -14850 53020 -14650 53090
rect -14350 53020 -14150 53090
rect -13850 53020 -13650 53090
rect -13350 53020 -13150 53090
rect -12850 53020 -12650 53090
rect -12350 53020 -12150 53090
rect -15850 52910 -15650 52980
rect -15350 52910 -15150 52980
rect -14850 52910 -14650 52980
rect -14350 52910 -14150 52980
rect -13850 52910 -13650 52980
rect -13350 52910 -13150 52980
rect -12850 52910 -12650 52980
rect -12350 52910 -12150 52980
rect -15980 52650 -15910 52850
rect -15590 52650 -15520 52850
rect -15480 52650 -15410 52850
rect -15090 52650 -15020 52850
rect -14980 52650 -14910 52850
rect -14590 52650 -14520 52850
rect -14480 52650 -14410 52850
rect -14090 52650 -14020 52850
rect -13980 52650 -13910 52850
rect -13590 52650 -13520 52850
rect -13480 52650 -13410 52850
rect -13090 52650 -13020 52850
rect -12980 52650 -12910 52850
rect -12590 52650 -12520 52850
rect -12480 52650 -12410 52850
rect -12090 52650 -12020 52850
rect -15850 52520 -15650 52590
rect -15350 52520 -15150 52590
rect -14850 52520 -14650 52590
rect -14350 52520 -14150 52590
rect -13850 52520 -13650 52590
rect -13350 52520 -13150 52590
rect -12850 52520 -12650 52590
rect -12350 52520 -12150 52590
rect -15850 52410 -15650 52480
rect -15350 52410 -15150 52480
rect -14850 52410 -14650 52480
rect -14350 52410 -14150 52480
rect -13850 52410 -13650 52480
rect -13350 52410 -13150 52480
rect -12850 52410 -12650 52480
rect -12350 52410 -12150 52480
rect -15980 52150 -15910 52350
rect -15590 52150 -15520 52350
rect -15480 52150 -15410 52350
rect -15090 52150 -15020 52350
rect -14980 52150 -14910 52350
rect -14590 52150 -14520 52350
rect -14480 52150 -14410 52350
rect -14090 52150 -14020 52350
rect -13980 52150 -13910 52350
rect -13590 52150 -13520 52350
rect -13480 52150 -13410 52350
rect -13090 52150 -13020 52350
rect -12980 52150 -12910 52350
rect -12590 52150 -12520 52350
rect -12480 52150 -12410 52350
rect -12090 52150 -12020 52350
rect -15850 52020 -15650 52090
rect -15350 52020 -15150 52090
rect -14850 52020 -14650 52090
rect -14350 52020 -14150 52090
rect -13850 52020 -13650 52090
rect -13350 52020 -13150 52090
rect -12850 52020 -12650 52090
rect -12350 52020 -12150 52090
rect -15850 51910 -15650 51980
rect -15350 51910 -15150 51980
rect -14850 51910 -14650 51980
rect -14350 51910 -14150 51980
rect -13850 51910 -13650 51980
rect -13350 51910 -13150 51980
rect -12850 51910 -12650 51980
rect -12350 51910 -12150 51980
rect -15980 51650 -15910 51850
rect -15590 51650 -15520 51850
rect -15480 51650 -15410 51850
rect -15090 51650 -15020 51850
rect -14980 51650 -14910 51850
rect -14590 51650 -14520 51850
rect -14480 51650 -14410 51850
rect -14090 51650 -14020 51850
rect -13980 51650 -13910 51850
rect -13590 51650 -13520 51850
rect -13480 51650 -13410 51850
rect -13090 51650 -13020 51850
rect -12980 51650 -12910 51850
rect -12590 51650 -12520 51850
rect -12480 51650 -12410 51850
rect -12090 51650 -12020 51850
rect -15850 51520 -15650 51590
rect -15350 51520 -15150 51590
rect -14850 51520 -14650 51590
rect -14350 51520 -14150 51590
rect -13850 51520 -13650 51590
rect -13350 51520 -13150 51590
rect -12850 51520 -12650 51590
rect -12350 51520 -12150 51590
rect -15850 51410 -15650 51480
rect -15350 51410 -15150 51480
rect -14850 51410 -14650 51480
rect -14350 51410 -14150 51480
rect -13850 51410 -13650 51480
rect -13350 51410 -13150 51480
rect -12850 51410 -12650 51480
rect -12350 51410 -12150 51480
rect -15980 51150 -15910 51350
rect -15590 51150 -15520 51350
rect -15480 51150 -15410 51350
rect -15090 51150 -15020 51350
rect -14980 51150 -14910 51350
rect -14590 51150 -14520 51350
rect -14480 51150 -14410 51350
rect -14090 51150 -14020 51350
rect -13980 51150 -13910 51350
rect -13590 51150 -13520 51350
rect -13480 51150 -13410 51350
rect -13090 51150 -13020 51350
rect -12980 51150 -12910 51350
rect -12590 51150 -12520 51350
rect -12480 51150 -12410 51350
rect -12090 51150 -12020 51350
rect -15850 51020 -15650 51090
rect -15350 51020 -15150 51090
rect -14850 51020 -14650 51090
rect -14350 51020 -14150 51090
rect -13850 51020 -13650 51090
rect -13350 51020 -13150 51090
rect -12850 51020 -12650 51090
rect -12350 51020 -12150 51090
rect -15850 50910 -15650 50980
rect -15350 50910 -15150 50980
rect -14850 50910 -14650 50980
rect -14350 50910 -14150 50980
rect -13850 50910 -13650 50980
rect -13350 50910 -13150 50980
rect -12850 50910 -12650 50980
rect -12350 50910 -12150 50980
rect -15980 50650 -15910 50850
rect -15590 50650 -15520 50850
rect -15480 50650 -15410 50850
rect -15090 50650 -15020 50850
rect -14980 50650 -14910 50850
rect -14590 50650 -14520 50850
rect -14480 50650 -14410 50850
rect -14090 50650 -14020 50850
rect -13980 50650 -13910 50850
rect -13590 50650 -13520 50850
rect -13480 50650 -13410 50850
rect -13090 50650 -13020 50850
rect -12980 50650 -12910 50850
rect -12590 50650 -12520 50850
rect -12480 50650 -12410 50850
rect -12090 50650 -12020 50850
rect -15850 50520 -15650 50590
rect -15350 50520 -15150 50590
rect -14850 50520 -14650 50590
rect -14350 50520 -14150 50590
rect -13850 50520 -13650 50590
rect -13350 50520 -13150 50590
rect -12850 50520 -12650 50590
rect -12350 50520 -12150 50590
rect -15850 50410 -15650 50480
rect -15350 50410 -15150 50480
rect -14850 50410 -14650 50480
rect -14350 50410 -14150 50480
rect -13850 50410 -13650 50480
rect -13350 50410 -13150 50480
rect -12850 50410 -12650 50480
rect -12350 50410 -12150 50480
rect -15980 50150 -15910 50350
rect -15590 50150 -15520 50350
rect -15480 50150 -15410 50350
rect -15090 50150 -15020 50350
rect -14980 50150 -14910 50350
rect -14590 50150 -14520 50350
rect -14480 50150 -14410 50350
rect -14090 50150 -14020 50350
rect -13980 50150 -13910 50350
rect -13590 50150 -13520 50350
rect -13480 50150 -13410 50350
rect -13090 50150 -13020 50350
rect -12980 50150 -12910 50350
rect -12590 50150 -12520 50350
rect -12480 50150 -12410 50350
rect -12090 50150 -12020 50350
rect -15850 50020 -15650 50090
rect -15350 50020 -15150 50090
rect -14850 50020 -14650 50090
rect -14350 50020 -14150 50090
rect -13850 50020 -13650 50090
rect -13350 50020 -13150 50090
rect -12850 50020 -12650 50090
rect -12350 50020 -12150 50090
rect 96150 85910 96350 85980
rect 96650 85910 96850 85980
rect 97150 85910 97350 85980
rect 97650 85910 97850 85980
rect 98150 85910 98350 85980
rect 98650 85910 98850 85980
rect 99150 85910 99350 85980
rect 99650 85910 99850 85980
rect 96020 85650 96090 85850
rect 96410 85650 96480 85850
rect 96520 85650 96590 85850
rect 96910 85650 96980 85850
rect 97020 85650 97090 85850
rect 97410 85650 97480 85850
rect 97520 85650 97590 85850
rect 97910 85650 97980 85850
rect 98020 85650 98090 85850
rect 98410 85650 98480 85850
rect 98520 85650 98590 85850
rect 98910 85650 98980 85850
rect 99020 85650 99090 85850
rect 99410 85650 99480 85850
rect 99520 85650 99590 85850
rect 99910 85650 99980 85850
rect 96150 85520 96350 85590
rect 96650 85520 96850 85590
rect 97150 85520 97350 85590
rect 97650 85520 97850 85590
rect 98150 85520 98350 85590
rect 98650 85520 98850 85590
rect 99150 85520 99350 85590
rect 99650 85520 99850 85590
rect 96150 85410 96350 85480
rect 96650 85410 96850 85480
rect 97150 85410 97350 85480
rect 97650 85410 97850 85480
rect 98150 85410 98350 85480
rect 98650 85410 98850 85480
rect 99150 85410 99350 85480
rect 99650 85410 99850 85480
rect 96020 85150 96090 85350
rect 96410 85150 96480 85350
rect 96520 85150 96590 85350
rect 96910 85150 96980 85350
rect 97020 85150 97090 85350
rect 97410 85150 97480 85350
rect 97520 85150 97590 85350
rect 97910 85150 97980 85350
rect 98020 85150 98090 85350
rect 98410 85150 98480 85350
rect 98520 85150 98590 85350
rect 98910 85150 98980 85350
rect 99020 85150 99090 85350
rect 99410 85150 99480 85350
rect 99520 85150 99590 85350
rect 99910 85150 99980 85350
rect 96150 85020 96350 85090
rect 96650 85020 96850 85090
rect 97150 85020 97350 85090
rect 97650 85020 97850 85090
rect 98150 85020 98350 85090
rect 98650 85020 98850 85090
rect 99150 85020 99350 85090
rect 99650 85020 99850 85090
rect 96150 84910 96350 84980
rect 96650 84910 96850 84980
rect 97150 84910 97350 84980
rect 97650 84910 97850 84980
rect 98150 84910 98350 84980
rect 98650 84910 98850 84980
rect 99150 84910 99350 84980
rect 99650 84910 99850 84980
rect 96020 84650 96090 84850
rect 96410 84650 96480 84850
rect 96520 84650 96590 84850
rect 96910 84650 96980 84850
rect 97020 84650 97090 84850
rect 97410 84650 97480 84850
rect 97520 84650 97590 84850
rect 97910 84650 97980 84850
rect 98020 84650 98090 84850
rect 98410 84650 98480 84850
rect 98520 84650 98590 84850
rect 98910 84650 98980 84850
rect 99020 84650 99090 84850
rect 99410 84650 99480 84850
rect 99520 84650 99590 84850
rect 99910 84650 99980 84850
rect 96150 84520 96350 84590
rect 96650 84520 96850 84590
rect 97150 84520 97350 84590
rect 97650 84520 97850 84590
rect 98150 84520 98350 84590
rect 98650 84520 98850 84590
rect 99150 84520 99350 84590
rect 99650 84520 99850 84590
rect 96150 84410 96350 84480
rect 96650 84410 96850 84480
rect 97150 84410 97350 84480
rect 97650 84410 97850 84480
rect 98150 84410 98350 84480
rect 98650 84410 98850 84480
rect 99150 84410 99350 84480
rect 99650 84410 99850 84480
rect 96020 84150 96090 84350
rect 96410 84150 96480 84350
rect 96520 84150 96590 84350
rect 96910 84150 96980 84350
rect 97020 84150 97090 84350
rect 97410 84150 97480 84350
rect 97520 84150 97590 84350
rect 97910 84150 97980 84350
rect 98020 84150 98090 84350
rect 98410 84150 98480 84350
rect 98520 84150 98590 84350
rect 98910 84150 98980 84350
rect 99020 84150 99090 84350
rect 99410 84150 99480 84350
rect 99520 84150 99590 84350
rect 99910 84150 99980 84350
rect 96150 84020 96350 84090
rect 96650 84020 96850 84090
rect 97150 84020 97350 84090
rect 97650 84020 97850 84090
rect 98150 84020 98350 84090
rect 98650 84020 98850 84090
rect 99150 84020 99350 84090
rect 99650 84020 99850 84090
rect 96150 83910 96350 83980
rect 96650 83910 96850 83980
rect 97150 83910 97350 83980
rect 97650 83910 97850 83980
rect 98150 83910 98350 83980
rect 98650 83910 98850 83980
rect 99150 83910 99350 83980
rect 99650 83910 99850 83980
rect 96020 83650 96090 83850
rect 96410 83650 96480 83850
rect 96520 83650 96590 83850
rect 96910 83650 96980 83850
rect 97020 83650 97090 83850
rect 97410 83650 97480 83850
rect 97520 83650 97590 83850
rect 97910 83650 97980 83850
rect 98020 83650 98090 83850
rect 98410 83650 98480 83850
rect 98520 83650 98590 83850
rect 98910 83650 98980 83850
rect 99020 83650 99090 83850
rect 99410 83650 99480 83850
rect 99520 83650 99590 83850
rect 99910 83650 99980 83850
rect 96150 83520 96350 83590
rect 96650 83520 96850 83590
rect 97150 83520 97350 83590
rect 97650 83520 97850 83590
rect 98150 83520 98350 83590
rect 98650 83520 98850 83590
rect 99150 83520 99350 83590
rect 99650 83520 99850 83590
rect 96150 83410 96350 83480
rect 96650 83410 96850 83480
rect 97150 83410 97350 83480
rect 97650 83410 97850 83480
rect 98150 83410 98350 83480
rect 98650 83410 98850 83480
rect 99150 83410 99350 83480
rect 99650 83410 99850 83480
rect 96020 83150 96090 83350
rect 96410 83150 96480 83350
rect 96520 83150 96590 83350
rect 96910 83150 96980 83350
rect 97020 83150 97090 83350
rect 97410 83150 97480 83350
rect 97520 83150 97590 83350
rect 97910 83150 97980 83350
rect 98020 83150 98090 83350
rect 98410 83150 98480 83350
rect 98520 83150 98590 83350
rect 98910 83150 98980 83350
rect 99020 83150 99090 83350
rect 99410 83150 99480 83350
rect 99520 83150 99590 83350
rect 99910 83150 99980 83350
rect 96150 83020 96350 83090
rect 96650 83020 96850 83090
rect 97150 83020 97350 83090
rect 97650 83020 97850 83090
rect 98150 83020 98350 83090
rect 98650 83020 98850 83090
rect 99150 83020 99350 83090
rect 99650 83020 99850 83090
rect 96150 82910 96350 82980
rect 96650 82910 96850 82980
rect 97150 82910 97350 82980
rect 97650 82910 97850 82980
rect 98150 82910 98350 82980
rect 98650 82910 98850 82980
rect 99150 82910 99350 82980
rect 99650 82910 99850 82980
rect 96020 82650 96090 82850
rect 96410 82650 96480 82850
rect 96520 82650 96590 82850
rect 96910 82650 96980 82850
rect 97020 82650 97090 82850
rect 97410 82650 97480 82850
rect 97520 82650 97590 82850
rect 97910 82650 97980 82850
rect 98020 82650 98090 82850
rect 98410 82650 98480 82850
rect 98520 82650 98590 82850
rect 98910 82650 98980 82850
rect 99020 82650 99090 82850
rect 99410 82650 99480 82850
rect 99520 82650 99590 82850
rect 99910 82650 99980 82850
rect 96150 82520 96350 82590
rect 96650 82520 96850 82590
rect 97150 82520 97350 82590
rect 97650 82520 97850 82590
rect 98150 82520 98350 82590
rect 98650 82520 98850 82590
rect 99150 82520 99350 82590
rect 99650 82520 99850 82590
rect 96150 82410 96350 82480
rect 96650 82410 96850 82480
rect 97150 82410 97350 82480
rect 97650 82410 97850 82480
rect 98150 82410 98350 82480
rect 98650 82410 98850 82480
rect 99150 82410 99350 82480
rect 99650 82410 99850 82480
rect 96020 82150 96090 82350
rect 96410 82150 96480 82350
rect 96520 82150 96590 82350
rect 96910 82150 96980 82350
rect 97020 82150 97090 82350
rect 97410 82150 97480 82350
rect 97520 82150 97590 82350
rect 97910 82150 97980 82350
rect 98020 82150 98090 82350
rect 98410 82150 98480 82350
rect 98520 82150 98590 82350
rect 98910 82150 98980 82350
rect 99020 82150 99090 82350
rect 99410 82150 99480 82350
rect 99520 82150 99590 82350
rect 99910 82150 99980 82350
rect 96150 82020 96350 82090
rect 96650 82020 96850 82090
rect 97150 82020 97350 82090
rect 97650 82020 97850 82090
rect 98150 82020 98350 82090
rect 98650 82020 98850 82090
rect 99150 82020 99350 82090
rect 99650 82020 99850 82090
rect 96150 81910 96350 81980
rect 96650 81910 96850 81980
rect 97150 81910 97350 81980
rect 97650 81910 97850 81980
rect 98150 81910 98350 81980
rect 98650 81910 98850 81980
rect 99150 81910 99350 81980
rect 99650 81910 99850 81980
rect 96020 81650 96090 81850
rect 96410 81650 96480 81850
rect 96520 81650 96590 81850
rect 96910 81650 96980 81850
rect 97020 81650 97090 81850
rect 97410 81650 97480 81850
rect 97520 81650 97590 81850
rect 97910 81650 97980 81850
rect 98020 81650 98090 81850
rect 98410 81650 98480 81850
rect 98520 81650 98590 81850
rect 98910 81650 98980 81850
rect 99020 81650 99090 81850
rect 99410 81650 99480 81850
rect 99520 81650 99590 81850
rect 99910 81650 99980 81850
rect 96150 81520 96350 81590
rect 96650 81520 96850 81590
rect 97150 81520 97350 81590
rect 97650 81520 97850 81590
rect 98150 81520 98350 81590
rect 98650 81520 98850 81590
rect 99150 81520 99350 81590
rect 99650 81520 99850 81590
rect 96150 81410 96350 81480
rect 96650 81410 96850 81480
rect 97150 81410 97350 81480
rect 97650 81410 97850 81480
rect 98150 81410 98350 81480
rect 98650 81410 98850 81480
rect 99150 81410 99350 81480
rect 99650 81410 99850 81480
rect 96020 81150 96090 81350
rect 96410 81150 96480 81350
rect 96520 81150 96590 81350
rect 96910 81150 96980 81350
rect 97020 81150 97090 81350
rect 97410 81150 97480 81350
rect 97520 81150 97590 81350
rect 97910 81150 97980 81350
rect 98020 81150 98090 81350
rect 98410 81150 98480 81350
rect 98520 81150 98590 81350
rect 98910 81150 98980 81350
rect 99020 81150 99090 81350
rect 99410 81150 99480 81350
rect 99520 81150 99590 81350
rect 99910 81150 99980 81350
rect 96150 81020 96350 81090
rect 96650 81020 96850 81090
rect 97150 81020 97350 81090
rect 97650 81020 97850 81090
rect 98150 81020 98350 81090
rect 98650 81020 98850 81090
rect 99150 81020 99350 81090
rect 99650 81020 99850 81090
rect 96150 80910 96350 80980
rect 96650 80910 96850 80980
rect 97150 80910 97350 80980
rect 97650 80910 97850 80980
rect 98150 80910 98350 80980
rect 98650 80910 98850 80980
rect 99150 80910 99350 80980
rect 99650 80910 99850 80980
rect 96020 80650 96090 80850
rect 96410 80650 96480 80850
rect 96520 80650 96590 80850
rect 96910 80650 96980 80850
rect 97020 80650 97090 80850
rect 97410 80650 97480 80850
rect 97520 80650 97590 80850
rect 97910 80650 97980 80850
rect 98020 80650 98090 80850
rect 98410 80650 98480 80850
rect 98520 80650 98590 80850
rect 98910 80650 98980 80850
rect 99020 80650 99090 80850
rect 99410 80650 99480 80850
rect 99520 80650 99590 80850
rect 99910 80650 99980 80850
rect 96150 80520 96350 80590
rect 96650 80520 96850 80590
rect 97150 80520 97350 80590
rect 97650 80520 97850 80590
rect 98150 80520 98350 80590
rect 98650 80520 98850 80590
rect 99150 80520 99350 80590
rect 99650 80520 99850 80590
rect 96150 80410 96350 80480
rect 96650 80410 96850 80480
rect 97150 80410 97350 80480
rect 97650 80410 97850 80480
rect 98150 80410 98350 80480
rect 98650 80410 98850 80480
rect 99150 80410 99350 80480
rect 99650 80410 99850 80480
rect 96020 80150 96090 80350
rect 96410 80150 96480 80350
rect 96520 80150 96590 80350
rect 96910 80150 96980 80350
rect 97020 80150 97090 80350
rect 97410 80150 97480 80350
rect 97520 80150 97590 80350
rect 97910 80150 97980 80350
rect 98020 80150 98090 80350
rect 98410 80150 98480 80350
rect 98520 80150 98590 80350
rect 98910 80150 98980 80350
rect 99020 80150 99090 80350
rect 99410 80150 99480 80350
rect 99520 80150 99590 80350
rect 99910 80150 99980 80350
rect 96150 80020 96350 80090
rect 96650 80020 96850 80090
rect 97150 80020 97350 80090
rect 97650 80020 97850 80090
rect 98150 80020 98350 80090
rect 98650 80020 98850 80090
rect 99150 80020 99350 80090
rect 99650 80020 99850 80090
rect 96150 79910 96350 79980
rect 96650 79910 96850 79980
rect 97150 79910 97350 79980
rect 97650 79910 97850 79980
rect 98150 79910 98350 79980
rect 98650 79910 98850 79980
rect 99150 79910 99350 79980
rect 99650 79910 99850 79980
rect 96020 79650 96090 79850
rect 96410 79650 96480 79850
rect 96520 79650 96590 79850
rect 96910 79650 96980 79850
rect 97020 79650 97090 79850
rect 97410 79650 97480 79850
rect 97520 79650 97590 79850
rect 97910 79650 97980 79850
rect 98020 79650 98090 79850
rect 98410 79650 98480 79850
rect 98520 79650 98590 79850
rect 98910 79650 98980 79850
rect 99020 79650 99090 79850
rect 99410 79650 99480 79850
rect 99520 79650 99590 79850
rect 99910 79650 99980 79850
rect 96150 79520 96350 79590
rect 96650 79520 96850 79590
rect 97150 79520 97350 79590
rect 97650 79520 97850 79590
rect 98150 79520 98350 79590
rect 98650 79520 98850 79590
rect 99150 79520 99350 79590
rect 99650 79520 99850 79590
rect 96150 79410 96350 79480
rect 96650 79410 96850 79480
rect 97150 79410 97350 79480
rect 97650 79410 97850 79480
rect 98150 79410 98350 79480
rect 98650 79410 98850 79480
rect 99150 79410 99350 79480
rect 99650 79410 99850 79480
rect 96020 79150 96090 79350
rect 96410 79150 96480 79350
rect 96520 79150 96590 79350
rect 96910 79150 96980 79350
rect 97020 79150 97090 79350
rect 97410 79150 97480 79350
rect 97520 79150 97590 79350
rect 97910 79150 97980 79350
rect 98020 79150 98090 79350
rect 98410 79150 98480 79350
rect 98520 79150 98590 79350
rect 98910 79150 98980 79350
rect 99020 79150 99090 79350
rect 99410 79150 99480 79350
rect 99520 79150 99590 79350
rect 99910 79150 99980 79350
rect 96150 79020 96350 79090
rect 96650 79020 96850 79090
rect 97150 79020 97350 79090
rect 97650 79020 97850 79090
rect 98150 79020 98350 79090
rect 98650 79020 98850 79090
rect 99150 79020 99350 79090
rect 99650 79020 99850 79090
rect 96150 78910 96350 78980
rect 96650 78910 96850 78980
rect 97150 78910 97350 78980
rect 97650 78910 97850 78980
rect 98150 78910 98350 78980
rect 98650 78910 98850 78980
rect 99150 78910 99350 78980
rect 99650 78910 99850 78980
rect 96020 78650 96090 78850
rect 96410 78650 96480 78850
rect 96520 78650 96590 78850
rect 96910 78650 96980 78850
rect 97020 78650 97090 78850
rect 97410 78650 97480 78850
rect 97520 78650 97590 78850
rect 97910 78650 97980 78850
rect 98020 78650 98090 78850
rect 98410 78650 98480 78850
rect 98520 78650 98590 78850
rect 98910 78650 98980 78850
rect 99020 78650 99090 78850
rect 99410 78650 99480 78850
rect 99520 78650 99590 78850
rect 99910 78650 99980 78850
rect 96150 78520 96350 78590
rect 96650 78520 96850 78590
rect 97150 78520 97350 78590
rect 97650 78520 97850 78590
rect 98150 78520 98350 78590
rect 98650 78520 98850 78590
rect 99150 78520 99350 78590
rect 99650 78520 99850 78590
rect 96150 78410 96350 78480
rect 96650 78410 96850 78480
rect 97150 78410 97350 78480
rect 97650 78410 97850 78480
rect 98150 78410 98350 78480
rect 98650 78410 98850 78480
rect 99150 78410 99350 78480
rect 99650 78410 99850 78480
rect 96020 78150 96090 78350
rect 96410 78150 96480 78350
rect 96520 78150 96590 78350
rect 96910 78150 96980 78350
rect 97020 78150 97090 78350
rect 97410 78150 97480 78350
rect 97520 78150 97590 78350
rect 97910 78150 97980 78350
rect 98020 78150 98090 78350
rect 98410 78150 98480 78350
rect 98520 78150 98590 78350
rect 98910 78150 98980 78350
rect 99020 78150 99090 78350
rect 99410 78150 99480 78350
rect 99520 78150 99590 78350
rect 99910 78150 99980 78350
rect 96150 78020 96350 78090
rect 96650 78020 96850 78090
rect 97150 78020 97350 78090
rect 97650 78020 97850 78090
rect 98150 78020 98350 78090
rect 98650 78020 98850 78090
rect 99150 78020 99350 78090
rect 99650 78020 99850 78090
rect 96150 77910 96350 77980
rect 96650 77910 96850 77980
rect 97150 77910 97350 77980
rect 97650 77910 97850 77980
rect 98150 77910 98350 77980
rect 98650 77910 98850 77980
rect 99150 77910 99350 77980
rect 99650 77910 99850 77980
rect 96020 77650 96090 77850
rect 96410 77650 96480 77850
rect 96520 77650 96590 77850
rect 96910 77650 96980 77850
rect 97020 77650 97090 77850
rect 97410 77650 97480 77850
rect 97520 77650 97590 77850
rect 97910 77650 97980 77850
rect 98020 77650 98090 77850
rect 98410 77650 98480 77850
rect 98520 77650 98590 77850
rect 98910 77650 98980 77850
rect 99020 77650 99090 77850
rect 99410 77650 99480 77850
rect 99520 77650 99590 77850
rect 99910 77650 99980 77850
rect 96150 77520 96350 77590
rect 96650 77520 96850 77590
rect 97150 77520 97350 77590
rect 97650 77520 97850 77590
rect 98150 77520 98350 77590
rect 98650 77520 98850 77590
rect 99150 77520 99350 77590
rect 99650 77520 99850 77590
rect 96150 77410 96350 77480
rect 96650 77410 96850 77480
rect 97150 77410 97350 77480
rect 97650 77410 97850 77480
rect 98150 77410 98350 77480
rect 98650 77410 98850 77480
rect 99150 77410 99350 77480
rect 99650 77410 99850 77480
rect 96020 77150 96090 77350
rect 96410 77150 96480 77350
rect 96520 77150 96590 77350
rect 96910 77150 96980 77350
rect 97020 77150 97090 77350
rect 97410 77150 97480 77350
rect 97520 77150 97590 77350
rect 97910 77150 97980 77350
rect 98020 77150 98090 77350
rect 98410 77150 98480 77350
rect 98520 77150 98590 77350
rect 98910 77150 98980 77350
rect 99020 77150 99090 77350
rect 99410 77150 99480 77350
rect 99520 77150 99590 77350
rect 99910 77150 99980 77350
rect 96150 77020 96350 77090
rect 96650 77020 96850 77090
rect 97150 77020 97350 77090
rect 97650 77020 97850 77090
rect 98150 77020 98350 77090
rect 98650 77020 98850 77090
rect 99150 77020 99350 77090
rect 99650 77020 99850 77090
rect 96150 76910 96350 76980
rect 96650 76910 96850 76980
rect 97150 76910 97350 76980
rect 97650 76910 97850 76980
rect 98150 76910 98350 76980
rect 98650 76910 98850 76980
rect 99150 76910 99350 76980
rect 99650 76910 99850 76980
rect 96020 76650 96090 76850
rect 96410 76650 96480 76850
rect 96520 76650 96590 76850
rect 96910 76650 96980 76850
rect 97020 76650 97090 76850
rect 97410 76650 97480 76850
rect 97520 76650 97590 76850
rect 97910 76650 97980 76850
rect 98020 76650 98090 76850
rect 98410 76650 98480 76850
rect 98520 76650 98590 76850
rect 98910 76650 98980 76850
rect 99020 76650 99090 76850
rect 99410 76650 99480 76850
rect 99520 76650 99590 76850
rect 99910 76650 99980 76850
rect 96150 76520 96350 76590
rect 96650 76520 96850 76590
rect 97150 76520 97350 76590
rect 97650 76520 97850 76590
rect 98150 76520 98350 76590
rect 98650 76520 98850 76590
rect 99150 76520 99350 76590
rect 99650 76520 99850 76590
rect 96150 76410 96350 76480
rect 96650 76410 96850 76480
rect 97150 76410 97350 76480
rect 97650 76410 97850 76480
rect 98150 76410 98350 76480
rect 98650 76410 98850 76480
rect 99150 76410 99350 76480
rect 99650 76410 99850 76480
rect 96020 76150 96090 76350
rect 96410 76150 96480 76350
rect 96520 76150 96590 76350
rect 96910 76150 96980 76350
rect 97020 76150 97090 76350
rect 97410 76150 97480 76350
rect 97520 76150 97590 76350
rect 97910 76150 97980 76350
rect 98020 76150 98090 76350
rect 98410 76150 98480 76350
rect 98520 76150 98590 76350
rect 98910 76150 98980 76350
rect 99020 76150 99090 76350
rect 99410 76150 99480 76350
rect 99520 76150 99590 76350
rect 99910 76150 99980 76350
rect 96150 76020 96350 76090
rect 96650 76020 96850 76090
rect 97150 76020 97350 76090
rect 97650 76020 97850 76090
rect 98150 76020 98350 76090
rect 98650 76020 98850 76090
rect 99150 76020 99350 76090
rect 99650 76020 99850 76090
rect 96150 75910 96350 75980
rect 96650 75910 96850 75980
rect 97150 75910 97350 75980
rect 97650 75910 97850 75980
rect 98150 75910 98350 75980
rect 98650 75910 98850 75980
rect 99150 75910 99350 75980
rect 99650 75910 99850 75980
rect 96020 75650 96090 75850
rect 96410 75650 96480 75850
rect 96520 75650 96590 75850
rect 96910 75650 96980 75850
rect 97020 75650 97090 75850
rect 97410 75650 97480 75850
rect 97520 75650 97590 75850
rect 97910 75650 97980 75850
rect 98020 75650 98090 75850
rect 98410 75650 98480 75850
rect 98520 75650 98590 75850
rect 98910 75650 98980 75850
rect 99020 75650 99090 75850
rect 99410 75650 99480 75850
rect 99520 75650 99590 75850
rect 99910 75650 99980 75850
rect 96150 75520 96350 75590
rect 96650 75520 96850 75590
rect 97150 75520 97350 75590
rect 97650 75520 97850 75590
rect 98150 75520 98350 75590
rect 98650 75520 98850 75590
rect 99150 75520 99350 75590
rect 99650 75520 99850 75590
rect 96150 75410 96350 75480
rect 96650 75410 96850 75480
rect 97150 75410 97350 75480
rect 97650 75410 97850 75480
rect 98150 75410 98350 75480
rect 98650 75410 98850 75480
rect 99150 75410 99350 75480
rect 99650 75410 99850 75480
rect 96020 75150 96090 75350
rect 96410 75150 96480 75350
rect 96520 75150 96590 75350
rect 96910 75150 96980 75350
rect 97020 75150 97090 75350
rect 97410 75150 97480 75350
rect 97520 75150 97590 75350
rect 97910 75150 97980 75350
rect 98020 75150 98090 75350
rect 98410 75150 98480 75350
rect 98520 75150 98590 75350
rect 98910 75150 98980 75350
rect 99020 75150 99090 75350
rect 99410 75150 99480 75350
rect 99520 75150 99590 75350
rect 99910 75150 99980 75350
rect 96150 75020 96350 75090
rect 96650 75020 96850 75090
rect 97150 75020 97350 75090
rect 97650 75020 97850 75090
rect 98150 75020 98350 75090
rect 98650 75020 98850 75090
rect 99150 75020 99350 75090
rect 99650 75020 99850 75090
rect 96150 74910 96350 74980
rect 96650 74910 96850 74980
rect 97150 74910 97350 74980
rect 97650 74910 97850 74980
rect 98150 74910 98350 74980
rect 98650 74910 98850 74980
rect 99150 74910 99350 74980
rect 99650 74910 99850 74980
rect 96020 74650 96090 74850
rect 96410 74650 96480 74850
rect 96520 74650 96590 74850
rect 96910 74650 96980 74850
rect 97020 74650 97090 74850
rect 97410 74650 97480 74850
rect 97520 74650 97590 74850
rect 97910 74650 97980 74850
rect 98020 74650 98090 74850
rect 98410 74650 98480 74850
rect 98520 74650 98590 74850
rect 98910 74650 98980 74850
rect 99020 74650 99090 74850
rect 99410 74650 99480 74850
rect 99520 74650 99590 74850
rect 99910 74650 99980 74850
rect 96150 74520 96350 74590
rect 96650 74520 96850 74590
rect 97150 74520 97350 74590
rect 97650 74520 97850 74590
rect 98150 74520 98350 74590
rect 98650 74520 98850 74590
rect 99150 74520 99350 74590
rect 99650 74520 99850 74590
rect 96150 74410 96350 74480
rect 96650 74410 96850 74480
rect 97150 74410 97350 74480
rect 97650 74410 97850 74480
rect 98150 74410 98350 74480
rect 98650 74410 98850 74480
rect 99150 74410 99350 74480
rect 99650 74410 99850 74480
rect 96020 74150 96090 74350
rect 96410 74150 96480 74350
rect 96520 74150 96590 74350
rect 96910 74150 96980 74350
rect 97020 74150 97090 74350
rect 97410 74150 97480 74350
rect 97520 74150 97590 74350
rect 97910 74150 97980 74350
rect 98020 74150 98090 74350
rect 98410 74150 98480 74350
rect 98520 74150 98590 74350
rect 98910 74150 98980 74350
rect 99020 74150 99090 74350
rect 99410 74150 99480 74350
rect 99520 74150 99590 74350
rect 99910 74150 99980 74350
rect 96150 74020 96350 74090
rect 96650 74020 96850 74090
rect 97150 74020 97350 74090
rect 97650 74020 97850 74090
rect 98150 74020 98350 74090
rect 98650 74020 98850 74090
rect 99150 74020 99350 74090
rect 99650 74020 99850 74090
rect 96150 73910 96350 73980
rect 96650 73910 96850 73980
rect 97150 73910 97350 73980
rect 97650 73910 97850 73980
rect 98150 73910 98350 73980
rect 98650 73910 98850 73980
rect 99150 73910 99350 73980
rect 99650 73910 99850 73980
rect 96020 73650 96090 73850
rect 96410 73650 96480 73850
rect 96520 73650 96590 73850
rect 96910 73650 96980 73850
rect 97020 73650 97090 73850
rect 97410 73650 97480 73850
rect 97520 73650 97590 73850
rect 97910 73650 97980 73850
rect 98020 73650 98090 73850
rect 98410 73650 98480 73850
rect 98520 73650 98590 73850
rect 98910 73650 98980 73850
rect 99020 73650 99090 73850
rect 99410 73650 99480 73850
rect 99520 73650 99590 73850
rect 99910 73650 99980 73850
rect 96150 73520 96350 73590
rect 96650 73520 96850 73590
rect 97150 73520 97350 73590
rect 97650 73520 97850 73590
rect 98150 73520 98350 73590
rect 98650 73520 98850 73590
rect 99150 73520 99350 73590
rect 99650 73520 99850 73590
rect 96150 73410 96350 73480
rect 96650 73410 96850 73480
rect 97150 73410 97350 73480
rect 97650 73410 97850 73480
rect 98150 73410 98350 73480
rect 98650 73410 98850 73480
rect 99150 73410 99350 73480
rect 99650 73410 99850 73480
rect 96020 73150 96090 73350
rect 96410 73150 96480 73350
rect 96520 73150 96590 73350
rect 96910 73150 96980 73350
rect 97020 73150 97090 73350
rect 97410 73150 97480 73350
rect 97520 73150 97590 73350
rect 97910 73150 97980 73350
rect 98020 73150 98090 73350
rect 98410 73150 98480 73350
rect 98520 73150 98590 73350
rect 98910 73150 98980 73350
rect 99020 73150 99090 73350
rect 99410 73150 99480 73350
rect 99520 73150 99590 73350
rect 99910 73150 99980 73350
rect 96150 73020 96350 73090
rect 96650 73020 96850 73090
rect 97150 73020 97350 73090
rect 97650 73020 97850 73090
rect 98150 73020 98350 73090
rect 98650 73020 98850 73090
rect 99150 73020 99350 73090
rect 99650 73020 99850 73090
rect 96150 72910 96350 72980
rect 96650 72910 96850 72980
rect 97150 72910 97350 72980
rect 97650 72910 97850 72980
rect 98150 72910 98350 72980
rect 98650 72910 98850 72980
rect 99150 72910 99350 72980
rect 99650 72910 99850 72980
rect 96020 72650 96090 72850
rect 96410 72650 96480 72850
rect 96520 72650 96590 72850
rect 96910 72650 96980 72850
rect 97020 72650 97090 72850
rect 97410 72650 97480 72850
rect 97520 72650 97590 72850
rect 97910 72650 97980 72850
rect 98020 72650 98090 72850
rect 98410 72650 98480 72850
rect 98520 72650 98590 72850
rect 98910 72650 98980 72850
rect 99020 72650 99090 72850
rect 99410 72650 99480 72850
rect 99520 72650 99590 72850
rect 99910 72650 99980 72850
rect 96150 72520 96350 72590
rect 96650 72520 96850 72590
rect 97150 72520 97350 72590
rect 97650 72520 97850 72590
rect 98150 72520 98350 72590
rect 98650 72520 98850 72590
rect 99150 72520 99350 72590
rect 99650 72520 99850 72590
rect 96150 72410 96350 72480
rect 96650 72410 96850 72480
rect 97150 72410 97350 72480
rect 97650 72410 97850 72480
rect 98150 72410 98350 72480
rect 98650 72410 98850 72480
rect 99150 72410 99350 72480
rect 99650 72410 99850 72480
rect 96020 72150 96090 72350
rect 96410 72150 96480 72350
rect 96520 72150 96590 72350
rect 96910 72150 96980 72350
rect 97020 72150 97090 72350
rect 97410 72150 97480 72350
rect 97520 72150 97590 72350
rect 97910 72150 97980 72350
rect 98020 72150 98090 72350
rect 98410 72150 98480 72350
rect 98520 72150 98590 72350
rect 98910 72150 98980 72350
rect 99020 72150 99090 72350
rect 99410 72150 99480 72350
rect 99520 72150 99590 72350
rect 99910 72150 99980 72350
rect 96150 72020 96350 72090
rect 96650 72020 96850 72090
rect 97150 72020 97350 72090
rect 97650 72020 97850 72090
rect 98150 72020 98350 72090
rect 98650 72020 98850 72090
rect 99150 72020 99350 72090
rect 99650 72020 99850 72090
rect 96150 71910 96350 71980
rect 96650 71910 96850 71980
rect 97150 71910 97350 71980
rect 97650 71910 97850 71980
rect 98150 71910 98350 71980
rect 98650 71910 98850 71980
rect 99150 71910 99350 71980
rect 99650 71910 99850 71980
rect 96020 71650 96090 71850
rect 96410 71650 96480 71850
rect 96520 71650 96590 71850
rect 96910 71650 96980 71850
rect 97020 71650 97090 71850
rect 97410 71650 97480 71850
rect 97520 71650 97590 71850
rect 97910 71650 97980 71850
rect 98020 71650 98090 71850
rect 98410 71650 98480 71850
rect 98520 71650 98590 71850
rect 98910 71650 98980 71850
rect 99020 71650 99090 71850
rect 99410 71650 99480 71850
rect 99520 71650 99590 71850
rect 99910 71650 99980 71850
rect 96150 71520 96350 71590
rect 96650 71520 96850 71590
rect 97150 71520 97350 71590
rect 97650 71520 97850 71590
rect 98150 71520 98350 71590
rect 98650 71520 98850 71590
rect 99150 71520 99350 71590
rect 99650 71520 99850 71590
rect 96150 71410 96350 71480
rect 96650 71410 96850 71480
rect 97150 71410 97350 71480
rect 97650 71410 97850 71480
rect 98150 71410 98350 71480
rect 98650 71410 98850 71480
rect 99150 71410 99350 71480
rect 99650 71410 99850 71480
rect 96020 71150 96090 71350
rect 96410 71150 96480 71350
rect 96520 71150 96590 71350
rect 96910 71150 96980 71350
rect 97020 71150 97090 71350
rect 97410 71150 97480 71350
rect 97520 71150 97590 71350
rect 97910 71150 97980 71350
rect 98020 71150 98090 71350
rect 98410 71150 98480 71350
rect 98520 71150 98590 71350
rect 98910 71150 98980 71350
rect 99020 71150 99090 71350
rect 99410 71150 99480 71350
rect 99520 71150 99590 71350
rect 99910 71150 99980 71350
rect 96150 71020 96350 71090
rect 96650 71020 96850 71090
rect 97150 71020 97350 71090
rect 97650 71020 97850 71090
rect 98150 71020 98350 71090
rect 98650 71020 98850 71090
rect 99150 71020 99350 71090
rect 99650 71020 99850 71090
rect 96150 70910 96350 70980
rect 96650 70910 96850 70980
rect 97150 70910 97350 70980
rect 97650 70910 97850 70980
rect 98150 70910 98350 70980
rect 98650 70910 98850 70980
rect 99150 70910 99350 70980
rect 99650 70910 99850 70980
rect 96020 70650 96090 70850
rect 96410 70650 96480 70850
rect 96520 70650 96590 70850
rect 96910 70650 96980 70850
rect 97020 70650 97090 70850
rect 97410 70650 97480 70850
rect 97520 70650 97590 70850
rect 97910 70650 97980 70850
rect 98020 70650 98090 70850
rect 98410 70650 98480 70850
rect 98520 70650 98590 70850
rect 98910 70650 98980 70850
rect 99020 70650 99090 70850
rect 99410 70650 99480 70850
rect 99520 70650 99590 70850
rect 99910 70650 99980 70850
rect 96150 70520 96350 70590
rect 96650 70520 96850 70590
rect 97150 70520 97350 70590
rect 97650 70520 97850 70590
rect 98150 70520 98350 70590
rect 98650 70520 98850 70590
rect 99150 70520 99350 70590
rect 99650 70520 99850 70590
rect 96150 70410 96350 70480
rect 96650 70410 96850 70480
rect 97150 70410 97350 70480
rect 97650 70410 97850 70480
rect 98150 70410 98350 70480
rect 98650 70410 98850 70480
rect 99150 70410 99350 70480
rect 99650 70410 99850 70480
rect 96020 70150 96090 70350
rect 96410 70150 96480 70350
rect 96520 70150 96590 70350
rect 96910 70150 96980 70350
rect 97020 70150 97090 70350
rect 97410 70150 97480 70350
rect 97520 70150 97590 70350
rect 97910 70150 97980 70350
rect 98020 70150 98090 70350
rect 98410 70150 98480 70350
rect 98520 70150 98590 70350
rect 98910 70150 98980 70350
rect 99020 70150 99090 70350
rect 99410 70150 99480 70350
rect 99520 70150 99590 70350
rect 99910 70150 99980 70350
rect 96150 70020 96350 70090
rect 96650 70020 96850 70090
rect 97150 70020 97350 70090
rect 97650 70020 97850 70090
rect 98150 70020 98350 70090
rect 98650 70020 98850 70090
rect 99150 70020 99350 70090
rect 99650 70020 99850 70090
rect 96150 69910 96350 69980
rect 96650 69910 96850 69980
rect 97150 69910 97350 69980
rect 97650 69910 97850 69980
rect 98150 69910 98350 69980
rect 98650 69910 98850 69980
rect 99150 69910 99350 69980
rect 99650 69910 99850 69980
rect 96020 69650 96090 69850
rect 96410 69650 96480 69850
rect 96520 69650 96590 69850
rect 96910 69650 96980 69850
rect 97020 69650 97090 69850
rect 97410 69650 97480 69850
rect 97520 69650 97590 69850
rect 97910 69650 97980 69850
rect 98020 69650 98090 69850
rect 98410 69650 98480 69850
rect 98520 69650 98590 69850
rect 98910 69650 98980 69850
rect 99020 69650 99090 69850
rect 99410 69650 99480 69850
rect 99520 69650 99590 69850
rect 99910 69650 99980 69850
rect 96150 69520 96350 69590
rect 96650 69520 96850 69590
rect 97150 69520 97350 69590
rect 97650 69520 97850 69590
rect 98150 69520 98350 69590
rect 98650 69520 98850 69590
rect 99150 69520 99350 69590
rect 99650 69520 99850 69590
rect 96150 69410 96350 69480
rect 96650 69410 96850 69480
rect 97150 69410 97350 69480
rect 97650 69410 97850 69480
rect 98150 69410 98350 69480
rect 98650 69410 98850 69480
rect 99150 69410 99350 69480
rect 99650 69410 99850 69480
rect 96020 69150 96090 69350
rect 96410 69150 96480 69350
rect 96520 69150 96590 69350
rect 96910 69150 96980 69350
rect 97020 69150 97090 69350
rect 97410 69150 97480 69350
rect 97520 69150 97590 69350
rect 97910 69150 97980 69350
rect 98020 69150 98090 69350
rect 98410 69150 98480 69350
rect 98520 69150 98590 69350
rect 98910 69150 98980 69350
rect 99020 69150 99090 69350
rect 99410 69150 99480 69350
rect 99520 69150 99590 69350
rect 99910 69150 99980 69350
rect 96150 69020 96350 69090
rect 96650 69020 96850 69090
rect 97150 69020 97350 69090
rect 97650 69020 97850 69090
rect 98150 69020 98350 69090
rect 98650 69020 98850 69090
rect 99150 69020 99350 69090
rect 99650 69020 99850 69090
rect 96150 68910 96350 68980
rect 96650 68910 96850 68980
rect 97150 68910 97350 68980
rect 97650 68910 97850 68980
rect 98150 68910 98350 68980
rect 98650 68910 98850 68980
rect 99150 68910 99350 68980
rect 99650 68910 99850 68980
rect 96020 68650 96090 68850
rect 96410 68650 96480 68850
rect 96520 68650 96590 68850
rect 96910 68650 96980 68850
rect 97020 68650 97090 68850
rect 97410 68650 97480 68850
rect 97520 68650 97590 68850
rect 97910 68650 97980 68850
rect 98020 68650 98090 68850
rect 98410 68650 98480 68850
rect 98520 68650 98590 68850
rect 98910 68650 98980 68850
rect 99020 68650 99090 68850
rect 99410 68650 99480 68850
rect 99520 68650 99590 68850
rect 99910 68650 99980 68850
rect 96150 68520 96350 68590
rect 96650 68520 96850 68590
rect 97150 68520 97350 68590
rect 97650 68520 97850 68590
rect 98150 68520 98350 68590
rect 98650 68520 98850 68590
rect 99150 68520 99350 68590
rect 99650 68520 99850 68590
rect 96150 68410 96350 68480
rect 96650 68410 96850 68480
rect 97150 68410 97350 68480
rect 97650 68410 97850 68480
rect 98150 68410 98350 68480
rect 98650 68410 98850 68480
rect 99150 68410 99350 68480
rect 99650 68410 99850 68480
rect 96020 68150 96090 68350
rect 96410 68150 96480 68350
rect 96520 68150 96590 68350
rect 96910 68150 96980 68350
rect 97020 68150 97090 68350
rect 97410 68150 97480 68350
rect 97520 68150 97590 68350
rect 97910 68150 97980 68350
rect 98020 68150 98090 68350
rect 98410 68150 98480 68350
rect 98520 68150 98590 68350
rect 98910 68150 98980 68350
rect 99020 68150 99090 68350
rect 99410 68150 99480 68350
rect 99520 68150 99590 68350
rect 99910 68150 99980 68350
rect 96150 68020 96350 68090
rect 96650 68020 96850 68090
rect 97150 68020 97350 68090
rect 97650 68020 97850 68090
rect 98150 68020 98350 68090
rect 98650 68020 98850 68090
rect 99150 68020 99350 68090
rect 99650 68020 99850 68090
rect 96150 67910 96350 67980
rect 96650 67910 96850 67980
rect 97150 67910 97350 67980
rect 97650 67910 97850 67980
rect 98150 67910 98350 67980
rect 98650 67910 98850 67980
rect 99150 67910 99350 67980
rect 99650 67910 99850 67980
rect 96020 67650 96090 67850
rect 96410 67650 96480 67850
rect 96520 67650 96590 67850
rect 96910 67650 96980 67850
rect 97020 67650 97090 67850
rect 97410 67650 97480 67850
rect 97520 67650 97590 67850
rect 97910 67650 97980 67850
rect 98020 67650 98090 67850
rect 98410 67650 98480 67850
rect 98520 67650 98590 67850
rect 98910 67650 98980 67850
rect 99020 67650 99090 67850
rect 99410 67650 99480 67850
rect 99520 67650 99590 67850
rect 99910 67650 99980 67850
rect 96150 67520 96350 67590
rect 96650 67520 96850 67590
rect 97150 67520 97350 67590
rect 97650 67520 97850 67590
rect 98150 67520 98350 67590
rect 98650 67520 98850 67590
rect 99150 67520 99350 67590
rect 99650 67520 99850 67590
rect 96150 67410 96350 67480
rect 96650 67410 96850 67480
rect 97150 67410 97350 67480
rect 97650 67410 97850 67480
rect 98150 67410 98350 67480
rect 98650 67410 98850 67480
rect 99150 67410 99350 67480
rect 99650 67410 99850 67480
rect 96020 67150 96090 67350
rect 96410 67150 96480 67350
rect 96520 67150 96590 67350
rect 96910 67150 96980 67350
rect 97020 67150 97090 67350
rect 97410 67150 97480 67350
rect 97520 67150 97590 67350
rect 97910 67150 97980 67350
rect 98020 67150 98090 67350
rect 98410 67150 98480 67350
rect 98520 67150 98590 67350
rect 98910 67150 98980 67350
rect 99020 67150 99090 67350
rect 99410 67150 99480 67350
rect 99520 67150 99590 67350
rect 99910 67150 99980 67350
rect 96150 67020 96350 67090
rect 96650 67020 96850 67090
rect 97150 67020 97350 67090
rect 97650 67020 97850 67090
rect 98150 67020 98350 67090
rect 98650 67020 98850 67090
rect 99150 67020 99350 67090
rect 99650 67020 99850 67090
rect 96150 66910 96350 66980
rect 96650 66910 96850 66980
rect 97150 66910 97350 66980
rect 97650 66910 97850 66980
rect 98150 66910 98350 66980
rect 98650 66910 98850 66980
rect 99150 66910 99350 66980
rect 99650 66910 99850 66980
rect 96020 66650 96090 66850
rect 96410 66650 96480 66850
rect 96520 66650 96590 66850
rect 96910 66650 96980 66850
rect 97020 66650 97090 66850
rect 97410 66650 97480 66850
rect 97520 66650 97590 66850
rect 97910 66650 97980 66850
rect 98020 66650 98090 66850
rect 98410 66650 98480 66850
rect 98520 66650 98590 66850
rect 98910 66650 98980 66850
rect 99020 66650 99090 66850
rect 99410 66650 99480 66850
rect 99520 66650 99590 66850
rect 99910 66650 99980 66850
rect 96150 66520 96350 66590
rect 96650 66520 96850 66590
rect 97150 66520 97350 66590
rect 97650 66520 97850 66590
rect 98150 66520 98350 66590
rect 98650 66520 98850 66590
rect 99150 66520 99350 66590
rect 99650 66520 99850 66590
rect 96150 66410 96350 66480
rect 96650 66410 96850 66480
rect 97150 66410 97350 66480
rect 97650 66410 97850 66480
rect 98150 66410 98350 66480
rect 98650 66410 98850 66480
rect 99150 66410 99350 66480
rect 99650 66410 99850 66480
rect 96020 66150 96090 66350
rect 96410 66150 96480 66350
rect 96520 66150 96590 66350
rect 96910 66150 96980 66350
rect 97020 66150 97090 66350
rect 97410 66150 97480 66350
rect 97520 66150 97590 66350
rect 97910 66150 97980 66350
rect 98020 66150 98090 66350
rect 98410 66150 98480 66350
rect 98520 66150 98590 66350
rect 98910 66150 98980 66350
rect 99020 66150 99090 66350
rect 99410 66150 99480 66350
rect 99520 66150 99590 66350
rect 99910 66150 99980 66350
rect 96150 66020 96350 66090
rect 96650 66020 96850 66090
rect 97150 66020 97350 66090
rect 97650 66020 97850 66090
rect 98150 66020 98350 66090
rect 98650 66020 98850 66090
rect 99150 66020 99350 66090
rect 99650 66020 99850 66090
rect 96150 65910 96350 65980
rect 96650 65910 96850 65980
rect 97150 65910 97350 65980
rect 97650 65910 97850 65980
rect 98150 65910 98350 65980
rect 98650 65910 98850 65980
rect 99150 65910 99350 65980
rect 99650 65910 99850 65980
rect 96020 65650 96090 65850
rect 96410 65650 96480 65850
rect 96520 65650 96590 65850
rect 96910 65650 96980 65850
rect 97020 65650 97090 65850
rect 97410 65650 97480 65850
rect 97520 65650 97590 65850
rect 97910 65650 97980 65850
rect 98020 65650 98090 65850
rect 98410 65650 98480 65850
rect 98520 65650 98590 65850
rect 98910 65650 98980 65850
rect 99020 65650 99090 65850
rect 99410 65650 99480 65850
rect 99520 65650 99590 65850
rect 99910 65650 99980 65850
rect 96150 65520 96350 65590
rect 96650 65520 96850 65590
rect 97150 65520 97350 65590
rect 97650 65520 97850 65590
rect 98150 65520 98350 65590
rect 98650 65520 98850 65590
rect 99150 65520 99350 65590
rect 99650 65520 99850 65590
rect 96150 65410 96350 65480
rect 96650 65410 96850 65480
rect 97150 65410 97350 65480
rect 97650 65410 97850 65480
rect 98150 65410 98350 65480
rect 98650 65410 98850 65480
rect 99150 65410 99350 65480
rect 99650 65410 99850 65480
rect 96020 65150 96090 65350
rect 96410 65150 96480 65350
rect 96520 65150 96590 65350
rect 96910 65150 96980 65350
rect 97020 65150 97090 65350
rect 97410 65150 97480 65350
rect 97520 65150 97590 65350
rect 97910 65150 97980 65350
rect 98020 65150 98090 65350
rect 98410 65150 98480 65350
rect 98520 65150 98590 65350
rect 98910 65150 98980 65350
rect 99020 65150 99090 65350
rect 99410 65150 99480 65350
rect 99520 65150 99590 65350
rect 99910 65150 99980 65350
rect 96150 65020 96350 65090
rect 96650 65020 96850 65090
rect 97150 65020 97350 65090
rect 97650 65020 97850 65090
rect 98150 65020 98350 65090
rect 98650 65020 98850 65090
rect 99150 65020 99350 65090
rect 99650 65020 99850 65090
rect 96150 64910 96350 64980
rect 96650 64910 96850 64980
rect 97150 64910 97350 64980
rect 97650 64910 97850 64980
rect 98150 64910 98350 64980
rect 98650 64910 98850 64980
rect 99150 64910 99350 64980
rect 99650 64910 99850 64980
rect 96020 64650 96090 64850
rect 96410 64650 96480 64850
rect 96520 64650 96590 64850
rect 96910 64650 96980 64850
rect 97020 64650 97090 64850
rect 97410 64650 97480 64850
rect 97520 64650 97590 64850
rect 97910 64650 97980 64850
rect 98020 64650 98090 64850
rect 98410 64650 98480 64850
rect 98520 64650 98590 64850
rect 98910 64650 98980 64850
rect 99020 64650 99090 64850
rect 99410 64650 99480 64850
rect 99520 64650 99590 64850
rect 99910 64650 99980 64850
rect 96150 64520 96350 64590
rect 96650 64520 96850 64590
rect 97150 64520 97350 64590
rect 97650 64520 97850 64590
rect 98150 64520 98350 64590
rect 98650 64520 98850 64590
rect 99150 64520 99350 64590
rect 99650 64520 99850 64590
rect 96150 64410 96350 64480
rect 96650 64410 96850 64480
rect 97150 64410 97350 64480
rect 97650 64410 97850 64480
rect 98150 64410 98350 64480
rect 98650 64410 98850 64480
rect 99150 64410 99350 64480
rect 99650 64410 99850 64480
rect 96020 64150 96090 64350
rect 96410 64150 96480 64350
rect 96520 64150 96590 64350
rect 96910 64150 96980 64350
rect 97020 64150 97090 64350
rect 97410 64150 97480 64350
rect 97520 64150 97590 64350
rect 97910 64150 97980 64350
rect 98020 64150 98090 64350
rect 98410 64150 98480 64350
rect 98520 64150 98590 64350
rect 98910 64150 98980 64350
rect 99020 64150 99090 64350
rect 99410 64150 99480 64350
rect 99520 64150 99590 64350
rect 99910 64150 99980 64350
rect 96150 64020 96350 64090
rect 96650 64020 96850 64090
rect 97150 64020 97350 64090
rect 97650 64020 97850 64090
rect 98150 64020 98350 64090
rect 98650 64020 98850 64090
rect 99150 64020 99350 64090
rect 99650 64020 99850 64090
rect 96150 63910 96350 63980
rect 96650 63910 96850 63980
rect 97150 63910 97350 63980
rect 97650 63910 97850 63980
rect 98150 63910 98350 63980
rect 98650 63910 98850 63980
rect 99150 63910 99350 63980
rect 99650 63910 99850 63980
rect 96020 63650 96090 63850
rect 96410 63650 96480 63850
rect 96520 63650 96590 63850
rect 96910 63650 96980 63850
rect 97020 63650 97090 63850
rect 97410 63650 97480 63850
rect 97520 63650 97590 63850
rect 97910 63650 97980 63850
rect 98020 63650 98090 63850
rect 98410 63650 98480 63850
rect 98520 63650 98590 63850
rect 98910 63650 98980 63850
rect 99020 63650 99090 63850
rect 99410 63650 99480 63850
rect 99520 63650 99590 63850
rect 99910 63650 99980 63850
rect 96150 63520 96350 63590
rect 96650 63520 96850 63590
rect 97150 63520 97350 63590
rect 97650 63520 97850 63590
rect 98150 63520 98350 63590
rect 98650 63520 98850 63590
rect 99150 63520 99350 63590
rect 99650 63520 99850 63590
rect 96150 63410 96350 63480
rect 96650 63410 96850 63480
rect 97150 63410 97350 63480
rect 97650 63410 97850 63480
rect 98150 63410 98350 63480
rect 98650 63410 98850 63480
rect 99150 63410 99350 63480
rect 99650 63410 99850 63480
rect 96020 63150 96090 63350
rect 96410 63150 96480 63350
rect 96520 63150 96590 63350
rect 96910 63150 96980 63350
rect 97020 63150 97090 63350
rect 97410 63150 97480 63350
rect 97520 63150 97590 63350
rect 97910 63150 97980 63350
rect 98020 63150 98090 63350
rect 98410 63150 98480 63350
rect 98520 63150 98590 63350
rect 98910 63150 98980 63350
rect 99020 63150 99090 63350
rect 99410 63150 99480 63350
rect 99520 63150 99590 63350
rect 99910 63150 99980 63350
rect 96150 63020 96350 63090
rect 96650 63020 96850 63090
rect 97150 63020 97350 63090
rect 97650 63020 97850 63090
rect 98150 63020 98350 63090
rect 98650 63020 98850 63090
rect 99150 63020 99350 63090
rect 99650 63020 99850 63090
rect 96150 62910 96350 62980
rect 96650 62910 96850 62980
rect 97150 62910 97350 62980
rect 97650 62910 97850 62980
rect 98150 62910 98350 62980
rect 98650 62910 98850 62980
rect 99150 62910 99350 62980
rect 99650 62910 99850 62980
rect 96020 62650 96090 62850
rect 96410 62650 96480 62850
rect 96520 62650 96590 62850
rect 96910 62650 96980 62850
rect 97020 62650 97090 62850
rect 97410 62650 97480 62850
rect 97520 62650 97590 62850
rect 97910 62650 97980 62850
rect 98020 62650 98090 62850
rect 98410 62650 98480 62850
rect 98520 62650 98590 62850
rect 98910 62650 98980 62850
rect 99020 62650 99090 62850
rect 99410 62650 99480 62850
rect 99520 62650 99590 62850
rect 99910 62650 99980 62850
rect 96150 62520 96350 62590
rect 96650 62520 96850 62590
rect 97150 62520 97350 62590
rect 97650 62520 97850 62590
rect 98150 62520 98350 62590
rect 98650 62520 98850 62590
rect 99150 62520 99350 62590
rect 99650 62520 99850 62590
rect 96150 62410 96350 62480
rect 96650 62410 96850 62480
rect 97150 62410 97350 62480
rect 97650 62410 97850 62480
rect 98150 62410 98350 62480
rect 98650 62410 98850 62480
rect 99150 62410 99350 62480
rect 99650 62410 99850 62480
rect 96020 62150 96090 62350
rect 96410 62150 96480 62350
rect 96520 62150 96590 62350
rect 96910 62150 96980 62350
rect 97020 62150 97090 62350
rect 97410 62150 97480 62350
rect 97520 62150 97590 62350
rect 97910 62150 97980 62350
rect 98020 62150 98090 62350
rect 98410 62150 98480 62350
rect 98520 62150 98590 62350
rect 98910 62150 98980 62350
rect 99020 62150 99090 62350
rect 99410 62150 99480 62350
rect 99520 62150 99590 62350
rect 99910 62150 99980 62350
rect 96150 62020 96350 62090
rect 96650 62020 96850 62090
rect 97150 62020 97350 62090
rect 97650 62020 97850 62090
rect 98150 62020 98350 62090
rect 98650 62020 98850 62090
rect 99150 62020 99350 62090
rect 99650 62020 99850 62090
rect 96150 61910 96350 61980
rect 96650 61910 96850 61980
rect 97150 61910 97350 61980
rect 97650 61910 97850 61980
rect 98150 61910 98350 61980
rect 98650 61910 98850 61980
rect 99150 61910 99350 61980
rect 99650 61910 99850 61980
rect 96020 61650 96090 61850
rect 96410 61650 96480 61850
rect 96520 61650 96590 61850
rect 96910 61650 96980 61850
rect 97020 61650 97090 61850
rect 97410 61650 97480 61850
rect 97520 61650 97590 61850
rect 97910 61650 97980 61850
rect 98020 61650 98090 61850
rect 98410 61650 98480 61850
rect 98520 61650 98590 61850
rect 98910 61650 98980 61850
rect 99020 61650 99090 61850
rect 99410 61650 99480 61850
rect 99520 61650 99590 61850
rect 99910 61650 99980 61850
rect 96150 61520 96350 61590
rect 96650 61520 96850 61590
rect 97150 61520 97350 61590
rect 97650 61520 97850 61590
rect 98150 61520 98350 61590
rect 98650 61520 98850 61590
rect 99150 61520 99350 61590
rect 99650 61520 99850 61590
rect 96150 61410 96350 61480
rect 96650 61410 96850 61480
rect 97150 61410 97350 61480
rect 97650 61410 97850 61480
rect 98150 61410 98350 61480
rect 98650 61410 98850 61480
rect 99150 61410 99350 61480
rect 99650 61410 99850 61480
rect 96020 61150 96090 61350
rect 96410 61150 96480 61350
rect 96520 61150 96590 61350
rect 96910 61150 96980 61350
rect 97020 61150 97090 61350
rect 97410 61150 97480 61350
rect 97520 61150 97590 61350
rect 97910 61150 97980 61350
rect 98020 61150 98090 61350
rect 98410 61150 98480 61350
rect 98520 61150 98590 61350
rect 98910 61150 98980 61350
rect 99020 61150 99090 61350
rect 99410 61150 99480 61350
rect 99520 61150 99590 61350
rect 99910 61150 99980 61350
rect 96150 61020 96350 61090
rect 96650 61020 96850 61090
rect 97150 61020 97350 61090
rect 97650 61020 97850 61090
rect 98150 61020 98350 61090
rect 98650 61020 98850 61090
rect 99150 61020 99350 61090
rect 99650 61020 99850 61090
rect 96150 60910 96350 60980
rect 96650 60910 96850 60980
rect 97150 60910 97350 60980
rect 97650 60910 97850 60980
rect 98150 60910 98350 60980
rect 98650 60910 98850 60980
rect 99150 60910 99350 60980
rect 99650 60910 99850 60980
rect 96020 60650 96090 60850
rect 96410 60650 96480 60850
rect 96520 60650 96590 60850
rect 96910 60650 96980 60850
rect 97020 60650 97090 60850
rect 97410 60650 97480 60850
rect 97520 60650 97590 60850
rect 97910 60650 97980 60850
rect 98020 60650 98090 60850
rect 98410 60650 98480 60850
rect 98520 60650 98590 60850
rect 98910 60650 98980 60850
rect 99020 60650 99090 60850
rect 99410 60650 99480 60850
rect 99520 60650 99590 60850
rect 99910 60650 99980 60850
rect 96150 60520 96350 60590
rect 96650 60520 96850 60590
rect 97150 60520 97350 60590
rect 97650 60520 97850 60590
rect 98150 60520 98350 60590
rect 98650 60520 98850 60590
rect 99150 60520 99350 60590
rect 99650 60520 99850 60590
rect 96150 60410 96350 60480
rect 96650 60410 96850 60480
rect 97150 60410 97350 60480
rect 97650 60410 97850 60480
rect 98150 60410 98350 60480
rect 98650 60410 98850 60480
rect 99150 60410 99350 60480
rect 99650 60410 99850 60480
rect 96020 60150 96090 60350
rect 96410 60150 96480 60350
rect 96520 60150 96590 60350
rect 96910 60150 96980 60350
rect 97020 60150 97090 60350
rect 97410 60150 97480 60350
rect 97520 60150 97590 60350
rect 97910 60150 97980 60350
rect 98020 60150 98090 60350
rect 98410 60150 98480 60350
rect 98520 60150 98590 60350
rect 98910 60150 98980 60350
rect 99020 60150 99090 60350
rect 99410 60150 99480 60350
rect 99520 60150 99590 60350
rect 99910 60150 99980 60350
rect 96150 60020 96350 60090
rect 96650 60020 96850 60090
rect 97150 60020 97350 60090
rect 97650 60020 97850 60090
rect 98150 60020 98350 60090
rect 98650 60020 98850 60090
rect 99150 60020 99350 60090
rect 99650 60020 99850 60090
rect 96150 59910 96350 59980
rect 96650 59910 96850 59980
rect 97150 59910 97350 59980
rect 97650 59910 97850 59980
rect 98150 59910 98350 59980
rect 98650 59910 98850 59980
rect 99150 59910 99350 59980
rect 99650 59910 99850 59980
rect 96020 59650 96090 59850
rect 96410 59650 96480 59850
rect 96520 59650 96590 59850
rect 96910 59650 96980 59850
rect 97020 59650 97090 59850
rect 97410 59650 97480 59850
rect 97520 59650 97590 59850
rect 97910 59650 97980 59850
rect 98020 59650 98090 59850
rect 98410 59650 98480 59850
rect 98520 59650 98590 59850
rect 98910 59650 98980 59850
rect 99020 59650 99090 59850
rect 99410 59650 99480 59850
rect 99520 59650 99590 59850
rect 99910 59650 99980 59850
rect 96150 59520 96350 59590
rect 96650 59520 96850 59590
rect 97150 59520 97350 59590
rect 97650 59520 97850 59590
rect 98150 59520 98350 59590
rect 98650 59520 98850 59590
rect 99150 59520 99350 59590
rect 99650 59520 99850 59590
rect 96150 59410 96350 59480
rect 96650 59410 96850 59480
rect 97150 59410 97350 59480
rect 97650 59410 97850 59480
rect 98150 59410 98350 59480
rect 98650 59410 98850 59480
rect 99150 59410 99350 59480
rect 99650 59410 99850 59480
rect 96020 59150 96090 59350
rect 96410 59150 96480 59350
rect 96520 59150 96590 59350
rect 96910 59150 96980 59350
rect 97020 59150 97090 59350
rect 97410 59150 97480 59350
rect 97520 59150 97590 59350
rect 97910 59150 97980 59350
rect 98020 59150 98090 59350
rect 98410 59150 98480 59350
rect 98520 59150 98590 59350
rect 98910 59150 98980 59350
rect 99020 59150 99090 59350
rect 99410 59150 99480 59350
rect 99520 59150 99590 59350
rect 99910 59150 99980 59350
rect 96150 59020 96350 59090
rect 96650 59020 96850 59090
rect 97150 59020 97350 59090
rect 97650 59020 97850 59090
rect 98150 59020 98350 59090
rect 98650 59020 98850 59090
rect 99150 59020 99350 59090
rect 99650 59020 99850 59090
rect 96150 58910 96350 58980
rect 96650 58910 96850 58980
rect 97150 58910 97350 58980
rect 97650 58910 97850 58980
rect 98150 58910 98350 58980
rect 98650 58910 98850 58980
rect 99150 58910 99350 58980
rect 99650 58910 99850 58980
rect 96020 58650 96090 58850
rect 96410 58650 96480 58850
rect 96520 58650 96590 58850
rect 96910 58650 96980 58850
rect 97020 58650 97090 58850
rect 97410 58650 97480 58850
rect 97520 58650 97590 58850
rect 97910 58650 97980 58850
rect 98020 58650 98090 58850
rect 98410 58650 98480 58850
rect 98520 58650 98590 58850
rect 98910 58650 98980 58850
rect 99020 58650 99090 58850
rect 99410 58650 99480 58850
rect 99520 58650 99590 58850
rect 99910 58650 99980 58850
rect 96150 58520 96350 58590
rect 96650 58520 96850 58590
rect 97150 58520 97350 58590
rect 97650 58520 97850 58590
rect 98150 58520 98350 58590
rect 98650 58520 98850 58590
rect 99150 58520 99350 58590
rect 99650 58520 99850 58590
rect 96150 58410 96350 58480
rect 96650 58410 96850 58480
rect 97150 58410 97350 58480
rect 97650 58410 97850 58480
rect 98150 58410 98350 58480
rect 98650 58410 98850 58480
rect 99150 58410 99350 58480
rect 99650 58410 99850 58480
rect 96020 58150 96090 58350
rect 96410 58150 96480 58350
rect 96520 58150 96590 58350
rect 96910 58150 96980 58350
rect 97020 58150 97090 58350
rect 97410 58150 97480 58350
rect 97520 58150 97590 58350
rect 97910 58150 97980 58350
rect 98020 58150 98090 58350
rect 98410 58150 98480 58350
rect 98520 58150 98590 58350
rect 98910 58150 98980 58350
rect 99020 58150 99090 58350
rect 99410 58150 99480 58350
rect 99520 58150 99590 58350
rect 99910 58150 99980 58350
rect 96150 58020 96350 58090
rect 96650 58020 96850 58090
rect 97150 58020 97350 58090
rect 97650 58020 97850 58090
rect 98150 58020 98350 58090
rect 98650 58020 98850 58090
rect 99150 58020 99350 58090
rect 99650 58020 99850 58090
rect 96150 57910 96350 57980
rect 96650 57910 96850 57980
rect 97150 57910 97350 57980
rect 97650 57910 97850 57980
rect 98150 57910 98350 57980
rect 98650 57910 98850 57980
rect 99150 57910 99350 57980
rect 99650 57910 99850 57980
rect 96020 57650 96090 57850
rect 96410 57650 96480 57850
rect 96520 57650 96590 57850
rect 96910 57650 96980 57850
rect 97020 57650 97090 57850
rect 97410 57650 97480 57850
rect 97520 57650 97590 57850
rect 97910 57650 97980 57850
rect 98020 57650 98090 57850
rect 98410 57650 98480 57850
rect 98520 57650 98590 57850
rect 98910 57650 98980 57850
rect 99020 57650 99090 57850
rect 99410 57650 99480 57850
rect 99520 57650 99590 57850
rect 99910 57650 99980 57850
rect 96150 57520 96350 57590
rect 96650 57520 96850 57590
rect 97150 57520 97350 57590
rect 97650 57520 97850 57590
rect 98150 57520 98350 57590
rect 98650 57520 98850 57590
rect 99150 57520 99350 57590
rect 99650 57520 99850 57590
rect 96150 57410 96350 57480
rect 96650 57410 96850 57480
rect 97150 57410 97350 57480
rect 97650 57410 97850 57480
rect 98150 57410 98350 57480
rect 98650 57410 98850 57480
rect 99150 57410 99350 57480
rect 99650 57410 99850 57480
rect 96020 57150 96090 57350
rect 96410 57150 96480 57350
rect 96520 57150 96590 57350
rect 96910 57150 96980 57350
rect 97020 57150 97090 57350
rect 97410 57150 97480 57350
rect 97520 57150 97590 57350
rect 97910 57150 97980 57350
rect 98020 57150 98090 57350
rect 98410 57150 98480 57350
rect 98520 57150 98590 57350
rect 98910 57150 98980 57350
rect 99020 57150 99090 57350
rect 99410 57150 99480 57350
rect 99520 57150 99590 57350
rect 99910 57150 99980 57350
rect 96150 57020 96350 57090
rect 96650 57020 96850 57090
rect 97150 57020 97350 57090
rect 97650 57020 97850 57090
rect 98150 57020 98350 57090
rect 98650 57020 98850 57090
rect 99150 57020 99350 57090
rect 99650 57020 99850 57090
rect 96150 56910 96350 56980
rect 96650 56910 96850 56980
rect 97150 56910 97350 56980
rect 97650 56910 97850 56980
rect 98150 56910 98350 56980
rect 98650 56910 98850 56980
rect 99150 56910 99350 56980
rect 99650 56910 99850 56980
rect 96020 56650 96090 56850
rect 96410 56650 96480 56850
rect 96520 56650 96590 56850
rect 96910 56650 96980 56850
rect 97020 56650 97090 56850
rect 97410 56650 97480 56850
rect 97520 56650 97590 56850
rect 97910 56650 97980 56850
rect 98020 56650 98090 56850
rect 98410 56650 98480 56850
rect 98520 56650 98590 56850
rect 98910 56650 98980 56850
rect 99020 56650 99090 56850
rect 99410 56650 99480 56850
rect 99520 56650 99590 56850
rect 99910 56650 99980 56850
rect 96150 56520 96350 56590
rect 96650 56520 96850 56590
rect 97150 56520 97350 56590
rect 97650 56520 97850 56590
rect 98150 56520 98350 56590
rect 98650 56520 98850 56590
rect 99150 56520 99350 56590
rect 99650 56520 99850 56590
rect 96150 56410 96350 56480
rect 96650 56410 96850 56480
rect 97150 56410 97350 56480
rect 97650 56410 97850 56480
rect 98150 56410 98350 56480
rect 98650 56410 98850 56480
rect 99150 56410 99350 56480
rect 99650 56410 99850 56480
rect 96020 56150 96090 56350
rect 96410 56150 96480 56350
rect 96520 56150 96590 56350
rect 96910 56150 96980 56350
rect 97020 56150 97090 56350
rect 97410 56150 97480 56350
rect 97520 56150 97590 56350
rect 97910 56150 97980 56350
rect 98020 56150 98090 56350
rect 98410 56150 98480 56350
rect 98520 56150 98590 56350
rect 98910 56150 98980 56350
rect 99020 56150 99090 56350
rect 99410 56150 99480 56350
rect 99520 56150 99590 56350
rect 99910 56150 99980 56350
rect 96150 56020 96350 56090
rect 96650 56020 96850 56090
rect 97150 56020 97350 56090
rect 97650 56020 97850 56090
rect 98150 56020 98350 56090
rect 98650 56020 98850 56090
rect 99150 56020 99350 56090
rect 99650 56020 99850 56090
rect 96150 55910 96350 55980
rect 96650 55910 96850 55980
rect 97150 55910 97350 55980
rect 97650 55910 97850 55980
rect 98150 55910 98350 55980
rect 98650 55910 98850 55980
rect 99150 55910 99350 55980
rect 99650 55910 99850 55980
rect 96020 55650 96090 55850
rect 96410 55650 96480 55850
rect 96520 55650 96590 55850
rect 96910 55650 96980 55850
rect 97020 55650 97090 55850
rect 97410 55650 97480 55850
rect 97520 55650 97590 55850
rect 97910 55650 97980 55850
rect 98020 55650 98090 55850
rect 98410 55650 98480 55850
rect 98520 55650 98590 55850
rect 98910 55650 98980 55850
rect 99020 55650 99090 55850
rect 99410 55650 99480 55850
rect 99520 55650 99590 55850
rect 99910 55650 99980 55850
rect 96150 55520 96350 55590
rect 96650 55520 96850 55590
rect 97150 55520 97350 55590
rect 97650 55520 97850 55590
rect 98150 55520 98350 55590
rect 98650 55520 98850 55590
rect 99150 55520 99350 55590
rect 99650 55520 99850 55590
rect 96150 55410 96350 55480
rect 96650 55410 96850 55480
rect 97150 55410 97350 55480
rect 97650 55410 97850 55480
rect 98150 55410 98350 55480
rect 98650 55410 98850 55480
rect 99150 55410 99350 55480
rect 99650 55410 99850 55480
rect 96020 55150 96090 55350
rect 96410 55150 96480 55350
rect 96520 55150 96590 55350
rect 96910 55150 96980 55350
rect 97020 55150 97090 55350
rect 97410 55150 97480 55350
rect 97520 55150 97590 55350
rect 97910 55150 97980 55350
rect 98020 55150 98090 55350
rect 98410 55150 98480 55350
rect 98520 55150 98590 55350
rect 98910 55150 98980 55350
rect 99020 55150 99090 55350
rect 99410 55150 99480 55350
rect 99520 55150 99590 55350
rect 99910 55150 99980 55350
rect 96150 55020 96350 55090
rect 96650 55020 96850 55090
rect 97150 55020 97350 55090
rect 97650 55020 97850 55090
rect 98150 55020 98350 55090
rect 98650 55020 98850 55090
rect 99150 55020 99350 55090
rect 99650 55020 99850 55090
rect 96150 54910 96350 54980
rect 96650 54910 96850 54980
rect 97150 54910 97350 54980
rect 97650 54910 97850 54980
rect 98150 54910 98350 54980
rect 98650 54910 98850 54980
rect 99150 54910 99350 54980
rect 99650 54910 99850 54980
rect 96020 54650 96090 54850
rect 96410 54650 96480 54850
rect 96520 54650 96590 54850
rect 96910 54650 96980 54850
rect 97020 54650 97090 54850
rect 97410 54650 97480 54850
rect 97520 54650 97590 54850
rect 97910 54650 97980 54850
rect 98020 54650 98090 54850
rect 98410 54650 98480 54850
rect 98520 54650 98590 54850
rect 98910 54650 98980 54850
rect 99020 54650 99090 54850
rect 99410 54650 99480 54850
rect 99520 54650 99590 54850
rect 99910 54650 99980 54850
rect 96150 54520 96350 54590
rect 96650 54520 96850 54590
rect 97150 54520 97350 54590
rect 97650 54520 97850 54590
rect 98150 54520 98350 54590
rect 98650 54520 98850 54590
rect 99150 54520 99350 54590
rect 99650 54520 99850 54590
rect 96150 54410 96350 54480
rect 96650 54410 96850 54480
rect 97150 54410 97350 54480
rect 97650 54410 97850 54480
rect 98150 54410 98350 54480
rect 98650 54410 98850 54480
rect 99150 54410 99350 54480
rect 99650 54410 99850 54480
rect 96020 54150 96090 54350
rect 96410 54150 96480 54350
rect 96520 54150 96590 54350
rect 96910 54150 96980 54350
rect 97020 54150 97090 54350
rect 97410 54150 97480 54350
rect 97520 54150 97590 54350
rect 97910 54150 97980 54350
rect 98020 54150 98090 54350
rect 98410 54150 98480 54350
rect 98520 54150 98590 54350
rect 98910 54150 98980 54350
rect 99020 54150 99090 54350
rect 99410 54150 99480 54350
rect 99520 54150 99590 54350
rect 99910 54150 99980 54350
rect 96150 54020 96350 54090
rect 96650 54020 96850 54090
rect 97150 54020 97350 54090
rect 97650 54020 97850 54090
rect 98150 54020 98350 54090
rect 98650 54020 98850 54090
rect 99150 54020 99350 54090
rect 99650 54020 99850 54090
rect 96150 53910 96350 53980
rect 96650 53910 96850 53980
rect 97150 53910 97350 53980
rect 97650 53910 97850 53980
rect 98150 53910 98350 53980
rect 98650 53910 98850 53980
rect 99150 53910 99350 53980
rect 99650 53910 99850 53980
rect 96020 53650 96090 53850
rect 96410 53650 96480 53850
rect 96520 53650 96590 53850
rect 96910 53650 96980 53850
rect 97020 53650 97090 53850
rect 97410 53650 97480 53850
rect 97520 53650 97590 53850
rect 97910 53650 97980 53850
rect 98020 53650 98090 53850
rect 98410 53650 98480 53850
rect 98520 53650 98590 53850
rect 98910 53650 98980 53850
rect 99020 53650 99090 53850
rect 99410 53650 99480 53850
rect 99520 53650 99590 53850
rect 99910 53650 99980 53850
rect 96150 53520 96350 53590
rect 96650 53520 96850 53590
rect 97150 53520 97350 53590
rect 97650 53520 97850 53590
rect 98150 53520 98350 53590
rect 98650 53520 98850 53590
rect 99150 53520 99350 53590
rect 99650 53520 99850 53590
rect 96150 53410 96350 53480
rect 96650 53410 96850 53480
rect 97150 53410 97350 53480
rect 97650 53410 97850 53480
rect 98150 53410 98350 53480
rect 98650 53410 98850 53480
rect 99150 53410 99350 53480
rect 99650 53410 99850 53480
rect 96020 53150 96090 53350
rect 96410 53150 96480 53350
rect 96520 53150 96590 53350
rect 96910 53150 96980 53350
rect 97020 53150 97090 53350
rect 97410 53150 97480 53350
rect 97520 53150 97590 53350
rect 97910 53150 97980 53350
rect 98020 53150 98090 53350
rect 98410 53150 98480 53350
rect 98520 53150 98590 53350
rect 98910 53150 98980 53350
rect 99020 53150 99090 53350
rect 99410 53150 99480 53350
rect 99520 53150 99590 53350
rect 99910 53150 99980 53350
rect 96150 53020 96350 53090
rect 96650 53020 96850 53090
rect 97150 53020 97350 53090
rect 97650 53020 97850 53090
rect 98150 53020 98350 53090
rect 98650 53020 98850 53090
rect 99150 53020 99350 53090
rect 99650 53020 99850 53090
rect 96150 52910 96350 52980
rect 96650 52910 96850 52980
rect 97150 52910 97350 52980
rect 97650 52910 97850 52980
rect 98150 52910 98350 52980
rect 98650 52910 98850 52980
rect 99150 52910 99350 52980
rect 99650 52910 99850 52980
rect 96020 52650 96090 52850
rect 96410 52650 96480 52850
rect 96520 52650 96590 52850
rect 96910 52650 96980 52850
rect 97020 52650 97090 52850
rect 97410 52650 97480 52850
rect 97520 52650 97590 52850
rect 97910 52650 97980 52850
rect 98020 52650 98090 52850
rect 98410 52650 98480 52850
rect 98520 52650 98590 52850
rect 98910 52650 98980 52850
rect 99020 52650 99090 52850
rect 99410 52650 99480 52850
rect 99520 52650 99590 52850
rect 99910 52650 99980 52850
rect 96150 52520 96350 52590
rect 96650 52520 96850 52590
rect 97150 52520 97350 52590
rect 97650 52520 97850 52590
rect 98150 52520 98350 52590
rect 98650 52520 98850 52590
rect 99150 52520 99350 52590
rect 99650 52520 99850 52590
rect 96150 52410 96350 52480
rect 96650 52410 96850 52480
rect 97150 52410 97350 52480
rect 97650 52410 97850 52480
rect 98150 52410 98350 52480
rect 98650 52410 98850 52480
rect 99150 52410 99350 52480
rect 99650 52410 99850 52480
rect 96020 52150 96090 52350
rect 96410 52150 96480 52350
rect 96520 52150 96590 52350
rect 96910 52150 96980 52350
rect 97020 52150 97090 52350
rect 97410 52150 97480 52350
rect 97520 52150 97590 52350
rect 97910 52150 97980 52350
rect 98020 52150 98090 52350
rect 98410 52150 98480 52350
rect 98520 52150 98590 52350
rect 98910 52150 98980 52350
rect 99020 52150 99090 52350
rect 99410 52150 99480 52350
rect 99520 52150 99590 52350
rect 99910 52150 99980 52350
rect 96150 52020 96350 52090
rect 96650 52020 96850 52090
rect 97150 52020 97350 52090
rect 97650 52020 97850 52090
rect 98150 52020 98350 52090
rect 98650 52020 98850 52090
rect 99150 52020 99350 52090
rect 99650 52020 99850 52090
rect 96150 51910 96350 51980
rect 96650 51910 96850 51980
rect 97150 51910 97350 51980
rect 97650 51910 97850 51980
rect 98150 51910 98350 51980
rect 98650 51910 98850 51980
rect 99150 51910 99350 51980
rect 99650 51910 99850 51980
rect 96020 51650 96090 51850
rect 96410 51650 96480 51850
rect 96520 51650 96590 51850
rect 96910 51650 96980 51850
rect 97020 51650 97090 51850
rect 97410 51650 97480 51850
rect 97520 51650 97590 51850
rect 97910 51650 97980 51850
rect 98020 51650 98090 51850
rect 98410 51650 98480 51850
rect 98520 51650 98590 51850
rect 98910 51650 98980 51850
rect 99020 51650 99090 51850
rect 99410 51650 99480 51850
rect 99520 51650 99590 51850
rect 99910 51650 99980 51850
rect 96150 51520 96350 51590
rect 96650 51520 96850 51590
rect 97150 51520 97350 51590
rect 97650 51520 97850 51590
rect 98150 51520 98350 51590
rect 98650 51520 98850 51590
rect 99150 51520 99350 51590
rect 99650 51520 99850 51590
rect 96150 51410 96350 51480
rect 96650 51410 96850 51480
rect 97150 51410 97350 51480
rect 97650 51410 97850 51480
rect 98150 51410 98350 51480
rect 98650 51410 98850 51480
rect 99150 51410 99350 51480
rect 99650 51410 99850 51480
rect 96020 51150 96090 51350
rect 96410 51150 96480 51350
rect 96520 51150 96590 51350
rect 96910 51150 96980 51350
rect 97020 51150 97090 51350
rect 97410 51150 97480 51350
rect 97520 51150 97590 51350
rect 97910 51150 97980 51350
rect 98020 51150 98090 51350
rect 98410 51150 98480 51350
rect 98520 51150 98590 51350
rect 98910 51150 98980 51350
rect 99020 51150 99090 51350
rect 99410 51150 99480 51350
rect 99520 51150 99590 51350
rect 99910 51150 99980 51350
rect 96150 51020 96350 51090
rect 96650 51020 96850 51090
rect 97150 51020 97350 51090
rect 97650 51020 97850 51090
rect 98150 51020 98350 51090
rect 98650 51020 98850 51090
rect 99150 51020 99350 51090
rect 99650 51020 99850 51090
rect 96150 50910 96350 50980
rect 96650 50910 96850 50980
rect 97150 50910 97350 50980
rect 97650 50910 97850 50980
rect 98150 50910 98350 50980
rect 98650 50910 98850 50980
rect 99150 50910 99350 50980
rect 99650 50910 99850 50980
rect 96020 50650 96090 50850
rect 96410 50650 96480 50850
rect 96520 50650 96590 50850
rect 96910 50650 96980 50850
rect 97020 50650 97090 50850
rect 97410 50650 97480 50850
rect 97520 50650 97590 50850
rect 97910 50650 97980 50850
rect 98020 50650 98090 50850
rect 98410 50650 98480 50850
rect 98520 50650 98590 50850
rect 98910 50650 98980 50850
rect 99020 50650 99090 50850
rect 99410 50650 99480 50850
rect 99520 50650 99590 50850
rect 99910 50650 99980 50850
rect 96150 50520 96350 50590
rect 96650 50520 96850 50590
rect 97150 50520 97350 50590
rect 97650 50520 97850 50590
rect 98150 50520 98350 50590
rect 98650 50520 98850 50590
rect 99150 50520 99350 50590
rect 99650 50520 99850 50590
rect 96150 50410 96350 50480
rect 96650 50410 96850 50480
rect 97150 50410 97350 50480
rect 97650 50410 97850 50480
rect 98150 50410 98350 50480
rect 98650 50410 98850 50480
rect 99150 50410 99350 50480
rect 99650 50410 99850 50480
rect 96020 50150 96090 50350
rect 96410 50150 96480 50350
rect 96520 50150 96590 50350
rect 96910 50150 96980 50350
rect 97020 50150 97090 50350
rect 97410 50150 97480 50350
rect 97520 50150 97590 50350
rect 97910 50150 97980 50350
rect 98020 50150 98090 50350
rect 98410 50150 98480 50350
rect 98520 50150 98590 50350
rect 98910 50150 98980 50350
rect 99020 50150 99090 50350
rect 99410 50150 99480 50350
rect 99520 50150 99590 50350
rect 99910 50150 99980 50350
rect 96150 50020 96350 50090
rect 96650 50020 96850 50090
rect 97150 50020 97350 50090
rect 97650 50020 97850 50090
rect 98150 50020 98350 50090
rect 98650 50020 98850 50090
rect 99150 50020 99350 50090
rect 99650 50020 99850 50090
rect -15850 49910 -15650 49980
rect -15350 49910 -15150 49980
rect -14850 49910 -14650 49980
rect -14350 49910 -14150 49980
rect -13850 49910 -13650 49980
rect -13350 49910 -13150 49980
rect -12850 49910 -12650 49980
rect -12350 49910 -12150 49980
rect -15980 49650 -15910 49850
rect -15590 49650 -15520 49850
rect -15480 49650 -15410 49850
rect -15090 49650 -15020 49850
rect -14980 49650 -14910 49850
rect -14590 49650 -14520 49850
rect -14480 49650 -14410 49850
rect -14090 49650 -14020 49850
rect -13980 49650 -13910 49850
rect -13590 49650 -13520 49850
rect -13480 49650 -13410 49850
rect -13090 49650 -13020 49850
rect -12980 49650 -12910 49850
rect -12590 49650 -12520 49850
rect -12480 49650 -12410 49850
rect -12090 49650 -12020 49850
rect -15850 49520 -15650 49590
rect -15350 49520 -15150 49590
rect -14850 49520 -14650 49590
rect -14350 49520 -14150 49590
rect -13850 49520 -13650 49590
rect -13350 49520 -13150 49590
rect -12850 49520 -12650 49590
rect -12350 49520 -12150 49590
rect -15850 49410 -15650 49480
rect -15350 49410 -15150 49480
rect -14850 49410 -14650 49480
rect -14350 49410 -14150 49480
rect -13850 49410 -13650 49480
rect -13350 49410 -13150 49480
rect -12850 49410 -12650 49480
rect -12350 49410 -12150 49480
rect -15980 49150 -15910 49350
rect -15590 49150 -15520 49350
rect -15480 49150 -15410 49350
rect -15090 49150 -15020 49350
rect -14980 49150 -14910 49350
rect -14590 49150 -14520 49350
rect -14480 49150 -14410 49350
rect -14090 49150 -14020 49350
rect -13980 49150 -13910 49350
rect -13590 49150 -13520 49350
rect -13480 49150 -13410 49350
rect -13090 49150 -13020 49350
rect -12980 49150 -12910 49350
rect -12590 49150 -12520 49350
rect -12480 49150 -12410 49350
rect -12090 49150 -12020 49350
rect -15850 49020 -15650 49090
rect -15350 49020 -15150 49090
rect -14850 49020 -14650 49090
rect -14350 49020 -14150 49090
rect -13850 49020 -13650 49090
rect -13350 49020 -13150 49090
rect -12850 49020 -12650 49090
rect -12350 49020 -12150 49090
rect -15850 48910 -15650 48980
rect -15350 48910 -15150 48980
rect -14850 48910 -14650 48980
rect -14350 48910 -14150 48980
rect -13850 48910 -13650 48980
rect -13350 48910 -13150 48980
rect -12850 48910 -12650 48980
rect -12350 48910 -12150 48980
rect -15980 48650 -15910 48850
rect -15590 48650 -15520 48850
rect -15480 48650 -15410 48850
rect -15090 48650 -15020 48850
rect -14980 48650 -14910 48850
rect -14590 48650 -14520 48850
rect -14480 48650 -14410 48850
rect -14090 48650 -14020 48850
rect -13980 48650 -13910 48850
rect -13590 48650 -13520 48850
rect -13480 48650 -13410 48850
rect -13090 48650 -13020 48850
rect -12980 48650 -12910 48850
rect -12590 48650 -12520 48850
rect -12480 48650 -12410 48850
rect -12090 48650 -12020 48850
rect -15850 48520 -15650 48590
rect -15350 48520 -15150 48590
rect -14850 48520 -14650 48590
rect -14350 48520 -14150 48590
rect -13850 48520 -13650 48590
rect -13350 48520 -13150 48590
rect -12850 48520 -12650 48590
rect -12350 48520 -12150 48590
rect -15850 48410 -15650 48480
rect -15350 48410 -15150 48480
rect -14850 48410 -14650 48480
rect -14350 48410 -14150 48480
rect -13850 48410 -13650 48480
rect -13350 48410 -13150 48480
rect -12850 48410 -12650 48480
rect -12350 48410 -12150 48480
rect -15980 48150 -15910 48350
rect -15590 48150 -15520 48350
rect -15480 48150 -15410 48350
rect -15090 48150 -15020 48350
rect -14980 48150 -14910 48350
rect -14590 48150 -14520 48350
rect -14480 48150 -14410 48350
rect -14090 48150 -14020 48350
rect -13980 48150 -13910 48350
rect -13590 48150 -13520 48350
rect -13480 48150 -13410 48350
rect -13090 48150 -13020 48350
rect -12980 48150 -12910 48350
rect -12590 48150 -12520 48350
rect -12480 48150 -12410 48350
rect -12090 48150 -12020 48350
rect -15850 48020 -15650 48090
rect -15350 48020 -15150 48090
rect -14850 48020 -14650 48090
rect -14350 48020 -14150 48090
rect -13850 48020 -13650 48090
rect -13350 48020 -13150 48090
rect -12850 48020 -12650 48090
rect -12350 48020 -12150 48090
rect -15850 47910 -15650 47980
rect -15350 47910 -15150 47980
rect -14850 47910 -14650 47980
rect -14350 47910 -14150 47980
rect -13850 47910 -13650 47980
rect -13350 47910 -13150 47980
rect -12850 47910 -12650 47980
rect -12350 47910 -12150 47980
rect -15980 47650 -15910 47850
rect -15590 47650 -15520 47850
rect -15480 47650 -15410 47850
rect -15090 47650 -15020 47850
rect -14980 47650 -14910 47850
rect -14590 47650 -14520 47850
rect -14480 47650 -14410 47850
rect -14090 47650 -14020 47850
rect -13980 47650 -13910 47850
rect -13590 47650 -13520 47850
rect -13480 47650 -13410 47850
rect -13090 47650 -13020 47850
rect -12980 47650 -12910 47850
rect -12590 47650 -12520 47850
rect -12480 47650 -12410 47850
rect -12090 47650 -12020 47850
rect -15850 47520 -15650 47590
rect -15350 47520 -15150 47590
rect -14850 47520 -14650 47590
rect -14350 47520 -14150 47590
rect -13850 47520 -13650 47590
rect -13350 47520 -13150 47590
rect -12850 47520 -12650 47590
rect -12350 47520 -12150 47590
rect -15850 47410 -15650 47480
rect -15350 47410 -15150 47480
rect -14850 47410 -14650 47480
rect -14350 47410 -14150 47480
rect -13850 47410 -13650 47480
rect -13350 47410 -13150 47480
rect -12850 47410 -12650 47480
rect -12350 47410 -12150 47480
rect -15980 47150 -15910 47350
rect -15590 47150 -15520 47350
rect -15480 47150 -15410 47350
rect -15090 47150 -15020 47350
rect -14980 47150 -14910 47350
rect -14590 47150 -14520 47350
rect -14480 47150 -14410 47350
rect -14090 47150 -14020 47350
rect -13980 47150 -13910 47350
rect -13590 47150 -13520 47350
rect -13480 47150 -13410 47350
rect -13090 47150 -13020 47350
rect -12980 47150 -12910 47350
rect -12590 47150 -12520 47350
rect -12480 47150 -12410 47350
rect -12090 47150 -12020 47350
rect -15850 47020 -15650 47090
rect -15350 47020 -15150 47090
rect -14850 47020 -14650 47090
rect -14350 47020 -14150 47090
rect -13850 47020 -13650 47090
rect -13350 47020 -13150 47090
rect -12850 47020 -12650 47090
rect -12350 47020 -12150 47090
rect -15850 46910 -15650 46980
rect -15350 46910 -15150 46980
rect -14850 46910 -14650 46980
rect -14350 46910 -14150 46980
rect -13850 46910 -13650 46980
rect -13350 46910 -13150 46980
rect -12850 46910 -12650 46980
rect -12350 46910 -12150 46980
rect -15980 46650 -15910 46850
rect -15590 46650 -15520 46850
rect -15480 46650 -15410 46850
rect -15090 46650 -15020 46850
rect -14980 46650 -14910 46850
rect -14590 46650 -14520 46850
rect -14480 46650 -14410 46850
rect -14090 46650 -14020 46850
rect -13980 46650 -13910 46850
rect -13590 46650 -13520 46850
rect -13480 46650 -13410 46850
rect -13090 46650 -13020 46850
rect -12980 46650 -12910 46850
rect -12590 46650 -12520 46850
rect -12480 46650 -12410 46850
rect -12090 46650 -12020 46850
rect -15850 46520 -15650 46590
rect -15350 46520 -15150 46590
rect -14850 46520 -14650 46590
rect -14350 46520 -14150 46590
rect -13850 46520 -13650 46590
rect -13350 46520 -13150 46590
rect -12850 46520 -12650 46590
rect -12350 46520 -12150 46590
rect -15850 46410 -15650 46480
rect -15350 46410 -15150 46480
rect -14850 46410 -14650 46480
rect -14350 46410 -14150 46480
rect -13850 46410 -13650 46480
rect -13350 46410 -13150 46480
rect -12850 46410 -12650 46480
rect -12350 46410 -12150 46480
rect -15980 46150 -15910 46350
rect -15590 46150 -15520 46350
rect -15480 46150 -15410 46350
rect -15090 46150 -15020 46350
rect -14980 46150 -14910 46350
rect -14590 46150 -14520 46350
rect -14480 46150 -14410 46350
rect -14090 46150 -14020 46350
rect -13980 46150 -13910 46350
rect -13590 46150 -13520 46350
rect -13480 46150 -13410 46350
rect -13090 46150 -13020 46350
rect -12980 46150 -12910 46350
rect -12590 46150 -12520 46350
rect -12480 46150 -12410 46350
rect -12090 46150 -12020 46350
rect -15850 46020 -15650 46090
rect -15350 46020 -15150 46090
rect -14850 46020 -14650 46090
rect -14350 46020 -14150 46090
rect -13850 46020 -13650 46090
rect -13350 46020 -13150 46090
rect -12850 46020 -12650 46090
rect -12350 46020 -12150 46090
rect -15850 45910 -15650 45980
rect -15350 45910 -15150 45980
rect -14850 45910 -14650 45980
rect -14350 45910 -14150 45980
rect -13850 45910 -13650 45980
rect -13350 45910 -13150 45980
rect -12850 45910 -12650 45980
rect -12350 45910 -12150 45980
rect -15980 45650 -15910 45850
rect -15590 45650 -15520 45850
rect -15480 45650 -15410 45850
rect -15090 45650 -15020 45850
rect -14980 45650 -14910 45850
rect -14590 45650 -14520 45850
rect -14480 45650 -14410 45850
rect -14090 45650 -14020 45850
rect -13980 45650 -13910 45850
rect -13590 45650 -13520 45850
rect -13480 45650 -13410 45850
rect -13090 45650 -13020 45850
rect -12980 45650 -12910 45850
rect -12590 45650 -12520 45850
rect -12480 45650 -12410 45850
rect -12090 45650 -12020 45850
rect -15850 45520 -15650 45590
rect -15350 45520 -15150 45590
rect -14850 45520 -14650 45590
rect -14350 45520 -14150 45590
rect -13850 45520 -13650 45590
rect -13350 45520 -13150 45590
rect -12850 45520 -12650 45590
rect -12350 45520 -12150 45590
rect -15850 45410 -15650 45480
rect -15350 45410 -15150 45480
rect -14850 45410 -14650 45480
rect -14350 45410 -14150 45480
rect -13850 45410 -13650 45480
rect -13350 45410 -13150 45480
rect -12850 45410 -12650 45480
rect -12350 45410 -12150 45480
rect -15980 45150 -15910 45350
rect -15590 45150 -15520 45350
rect -15480 45150 -15410 45350
rect -15090 45150 -15020 45350
rect -14980 45150 -14910 45350
rect -14590 45150 -14520 45350
rect -14480 45150 -14410 45350
rect -14090 45150 -14020 45350
rect -13980 45150 -13910 45350
rect -13590 45150 -13520 45350
rect -13480 45150 -13410 45350
rect -13090 45150 -13020 45350
rect -12980 45150 -12910 45350
rect -12590 45150 -12520 45350
rect -12480 45150 -12410 45350
rect -12090 45150 -12020 45350
rect -15850 45020 -15650 45090
rect -15350 45020 -15150 45090
rect -14850 45020 -14650 45090
rect -14350 45020 -14150 45090
rect -13850 45020 -13650 45090
rect -13350 45020 -13150 45090
rect -12850 45020 -12650 45090
rect -12350 45020 -12150 45090
rect -15850 44910 -15650 44980
rect -15350 44910 -15150 44980
rect -14850 44910 -14650 44980
rect -14350 44910 -14150 44980
rect -13850 44910 -13650 44980
rect -13350 44910 -13150 44980
rect -12850 44910 -12650 44980
rect -12350 44910 -12150 44980
rect -15980 44650 -15910 44850
rect -15590 44650 -15520 44850
rect -15480 44650 -15410 44850
rect -15090 44650 -15020 44850
rect -14980 44650 -14910 44850
rect -14590 44650 -14520 44850
rect -14480 44650 -14410 44850
rect -14090 44650 -14020 44850
rect -13980 44650 -13910 44850
rect -13590 44650 -13520 44850
rect -13480 44650 -13410 44850
rect -13090 44650 -13020 44850
rect -12980 44650 -12910 44850
rect -12590 44650 -12520 44850
rect -12480 44650 -12410 44850
rect -12090 44650 -12020 44850
rect -15850 44520 -15650 44590
rect -15350 44520 -15150 44590
rect -14850 44520 -14650 44590
rect -14350 44520 -14150 44590
rect -13850 44520 -13650 44590
rect -13350 44520 -13150 44590
rect -12850 44520 -12650 44590
rect -12350 44520 -12150 44590
rect -15850 44410 -15650 44480
rect -15350 44410 -15150 44480
rect -14850 44410 -14650 44480
rect -14350 44410 -14150 44480
rect -13850 44410 -13650 44480
rect -13350 44410 -13150 44480
rect -12850 44410 -12650 44480
rect -12350 44410 -12150 44480
rect -15980 44150 -15910 44350
rect -15590 44150 -15520 44350
rect -15480 44150 -15410 44350
rect -15090 44150 -15020 44350
rect -14980 44150 -14910 44350
rect -14590 44150 -14520 44350
rect -14480 44150 -14410 44350
rect -14090 44150 -14020 44350
rect -13980 44150 -13910 44350
rect -13590 44150 -13520 44350
rect -13480 44150 -13410 44350
rect -13090 44150 -13020 44350
rect -12980 44150 -12910 44350
rect -12590 44150 -12520 44350
rect -12480 44150 -12410 44350
rect -12090 44150 -12020 44350
rect -15850 44020 -15650 44090
rect -15350 44020 -15150 44090
rect -14850 44020 -14650 44090
rect -14350 44020 -14150 44090
rect -13850 44020 -13650 44090
rect -13350 44020 -13150 44090
rect -12850 44020 -12650 44090
rect -12350 44020 -12150 44090
rect -15850 43910 -15650 43980
rect -15350 43910 -15150 43980
rect -14850 43910 -14650 43980
rect -14350 43910 -14150 43980
rect -13850 43910 -13650 43980
rect -13350 43910 -13150 43980
rect -12850 43910 -12650 43980
rect -12350 43910 -12150 43980
rect -15980 43650 -15910 43850
rect -15590 43650 -15520 43850
rect -15480 43650 -15410 43850
rect -15090 43650 -15020 43850
rect -14980 43650 -14910 43850
rect -14590 43650 -14520 43850
rect -14480 43650 -14410 43850
rect -14090 43650 -14020 43850
rect -13980 43650 -13910 43850
rect -13590 43650 -13520 43850
rect -13480 43650 -13410 43850
rect -13090 43650 -13020 43850
rect -12980 43650 -12910 43850
rect -12590 43650 -12520 43850
rect -12480 43650 -12410 43850
rect -12090 43650 -12020 43850
rect -15850 43520 -15650 43590
rect -15350 43520 -15150 43590
rect -14850 43520 -14650 43590
rect -14350 43520 -14150 43590
rect -13850 43520 -13650 43590
rect -13350 43520 -13150 43590
rect -12850 43520 -12650 43590
rect -12350 43520 -12150 43590
rect -15850 43410 -15650 43480
rect -15350 43410 -15150 43480
rect -14850 43410 -14650 43480
rect -14350 43410 -14150 43480
rect -13850 43410 -13650 43480
rect -13350 43410 -13150 43480
rect -12850 43410 -12650 43480
rect -12350 43410 -12150 43480
rect -15980 43150 -15910 43350
rect -15590 43150 -15520 43350
rect -15480 43150 -15410 43350
rect -15090 43150 -15020 43350
rect -14980 43150 -14910 43350
rect -14590 43150 -14520 43350
rect -14480 43150 -14410 43350
rect -14090 43150 -14020 43350
rect -13980 43150 -13910 43350
rect -13590 43150 -13520 43350
rect -13480 43150 -13410 43350
rect -13090 43150 -13020 43350
rect -12980 43150 -12910 43350
rect -12590 43150 -12520 43350
rect -12480 43150 -12410 43350
rect -12090 43150 -12020 43350
rect -15850 43020 -15650 43090
rect -15350 43020 -15150 43090
rect -14850 43020 -14650 43090
rect -14350 43020 -14150 43090
rect -13850 43020 -13650 43090
rect -13350 43020 -13150 43090
rect -12850 43020 -12650 43090
rect -12350 43020 -12150 43090
rect -15850 42910 -15650 42980
rect -15350 42910 -15150 42980
rect -14850 42910 -14650 42980
rect -14350 42910 -14150 42980
rect -13850 42910 -13650 42980
rect -13350 42910 -13150 42980
rect -12850 42910 -12650 42980
rect -12350 42910 -12150 42980
rect -15980 42650 -15910 42850
rect -15590 42650 -15520 42850
rect -15480 42650 -15410 42850
rect -15090 42650 -15020 42850
rect -14980 42650 -14910 42850
rect -14590 42650 -14520 42850
rect -14480 42650 -14410 42850
rect -14090 42650 -14020 42850
rect -13980 42650 -13910 42850
rect -13590 42650 -13520 42850
rect -13480 42650 -13410 42850
rect -13090 42650 -13020 42850
rect -12980 42650 -12910 42850
rect -12590 42650 -12520 42850
rect -12480 42650 -12410 42850
rect -12090 42650 -12020 42850
rect -15850 42520 -15650 42590
rect -15350 42520 -15150 42590
rect -14850 42520 -14650 42590
rect -14350 42520 -14150 42590
rect -13850 42520 -13650 42590
rect -13350 42520 -13150 42590
rect -12850 42520 -12650 42590
rect -12350 42520 -12150 42590
rect -15850 42410 -15650 42480
rect -15350 42410 -15150 42480
rect -14850 42410 -14650 42480
rect -14350 42410 -14150 42480
rect -13850 42410 -13650 42480
rect -13350 42410 -13150 42480
rect -12850 42410 -12650 42480
rect -12350 42410 -12150 42480
rect -15980 42150 -15910 42350
rect -15590 42150 -15520 42350
rect -15480 42150 -15410 42350
rect -15090 42150 -15020 42350
rect -14980 42150 -14910 42350
rect -14590 42150 -14520 42350
rect -14480 42150 -14410 42350
rect -14090 42150 -14020 42350
rect -13980 42150 -13910 42350
rect -13590 42150 -13520 42350
rect -13480 42150 -13410 42350
rect -13090 42150 -13020 42350
rect -12980 42150 -12910 42350
rect -12590 42150 -12520 42350
rect -12480 42150 -12410 42350
rect -12090 42150 -12020 42350
rect -15850 42020 -15650 42090
rect -15350 42020 -15150 42090
rect -14850 42020 -14650 42090
rect -14350 42020 -14150 42090
rect -13850 42020 -13650 42090
rect -13350 42020 -13150 42090
rect -12850 42020 -12650 42090
rect -12350 42020 -12150 42090
rect -15850 41910 -15650 41980
rect -15350 41910 -15150 41980
rect -14850 41910 -14650 41980
rect -14350 41910 -14150 41980
rect -13850 41910 -13650 41980
rect -13350 41910 -13150 41980
rect -12850 41910 -12650 41980
rect -12350 41910 -12150 41980
rect -11850 41910 -11650 41980
rect -11350 41910 -11150 41980
rect -10850 41910 -10650 41980
rect -10350 41910 -10150 41980
rect -9850 41910 -9650 41980
rect -9350 41910 -9150 41980
rect -8850 41910 -8650 41980
rect -8350 41910 -8150 41980
rect -7850 41910 -7650 41980
rect -7350 41910 -7150 41980
rect -6850 41910 -6650 41980
rect -6350 41910 -6150 41980
rect -5850 41910 -5650 41980
rect -5350 41910 -5150 41980
rect -4850 41910 -4650 41980
rect -4350 41910 -4150 41980
rect -3850 41910 -3650 41980
rect -3350 41910 -3150 41980
rect -2850 41910 -2650 41980
rect -2350 41910 -2150 41980
rect -1850 41910 -1650 41980
rect -1350 41910 -1150 41980
rect -850 41910 -650 41980
rect -350 41910 -150 41980
rect 150 41910 350 41980
rect 650 41910 850 41980
rect 1150 41910 1350 41980
rect 1650 41910 1850 41980
rect 2150 41910 2350 41980
rect 2650 41910 2850 41980
rect 3150 41910 3350 41980
rect 3650 41910 3850 41980
rect -15980 41650 -15910 41850
rect -15590 41650 -15520 41850
rect -15480 41650 -15410 41850
rect -15090 41650 -15020 41850
rect -14980 41650 -14910 41850
rect -14590 41650 -14520 41850
rect -14480 41650 -14410 41850
rect -14090 41650 -14020 41850
rect -13980 41650 -13910 41850
rect -13590 41650 -13520 41850
rect -13480 41650 -13410 41850
rect -13090 41650 -13020 41850
rect -12980 41650 -12910 41850
rect -12590 41650 -12520 41850
rect -12480 41650 -12410 41850
rect -12090 41650 -12020 41850
rect -11980 41650 -11910 41850
rect -11590 41650 -11520 41850
rect -11480 41650 -11410 41850
rect -11090 41650 -11020 41850
rect -10980 41650 -10910 41850
rect -10590 41650 -10520 41850
rect -10480 41650 -10410 41850
rect -10090 41650 -10020 41850
rect -9980 41650 -9910 41850
rect -9590 41650 -9520 41850
rect -9480 41650 -9410 41850
rect -9090 41650 -9020 41850
rect -8980 41650 -8910 41850
rect -8590 41650 -8520 41850
rect -8480 41650 -8410 41850
rect -8090 41650 -8020 41850
rect -7980 41650 -7910 41850
rect -7590 41650 -7520 41850
rect -7480 41650 -7410 41850
rect -7090 41650 -7020 41850
rect -6980 41650 -6910 41850
rect -6590 41650 -6520 41850
rect -6480 41650 -6410 41850
rect -6090 41650 -6020 41850
rect -5980 41650 -5910 41850
rect -5590 41650 -5520 41850
rect -5480 41650 -5410 41850
rect -5090 41650 -5020 41850
rect -4980 41650 -4910 41850
rect -4590 41650 -4520 41850
rect -4480 41650 -4410 41850
rect -4090 41650 -4020 41850
rect -3980 41650 -3910 41850
rect -3590 41650 -3520 41850
rect -3480 41650 -3410 41850
rect -3090 41650 -3020 41850
rect -2980 41650 -2910 41850
rect -2590 41650 -2520 41850
rect -2480 41650 -2410 41850
rect -2090 41650 -2020 41850
rect -1980 41650 -1910 41850
rect -1590 41650 -1520 41850
rect -1480 41650 -1410 41850
rect -1090 41650 -1020 41850
rect -980 41650 -910 41850
rect -590 41650 -520 41850
rect -480 41650 -410 41850
rect -90 41650 -20 41850
rect 20 41650 90 41850
rect 410 41650 480 41850
rect 520 41650 590 41850
rect 910 41650 980 41850
rect 1020 41650 1090 41850
rect 1410 41650 1480 41850
rect 1520 41650 1590 41850
rect 1910 41650 1980 41850
rect 2020 41650 2090 41850
rect 2410 41650 2480 41850
rect 2520 41650 2590 41850
rect 2910 41650 2980 41850
rect 3020 41650 3090 41850
rect 3410 41650 3480 41850
rect 3520 41650 3590 41850
rect 3910 41650 3980 41850
rect -15850 41520 -15650 41590
rect -15350 41520 -15150 41590
rect -14850 41520 -14650 41590
rect -14350 41520 -14150 41590
rect -13850 41520 -13650 41590
rect -13350 41520 -13150 41590
rect -12850 41520 -12650 41590
rect -12350 41520 -12150 41590
rect -11850 41520 -11650 41590
rect -11350 41520 -11150 41590
rect -10850 41520 -10650 41590
rect -10350 41520 -10150 41590
rect -9850 41520 -9650 41590
rect -9350 41520 -9150 41590
rect -8850 41520 -8650 41590
rect -8350 41520 -8150 41590
rect -7850 41520 -7650 41590
rect -7350 41520 -7150 41590
rect -6850 41520 -6650 41590
rect -6350 41520 -6150 41590
rect -5850 41520 -5650 41590
rect -5350 41520 -5150 41590
rect -4850 41520 -4650 41590
rect -4350 41520 -4150 41590
rect -3850 41520 -3650 41590
rect -3350 41520 -3150 41590
rect -2850 41520 -2650 41590
rect -2350 41520 -2150 41590
rect -1850 41520 -1650 41590
rect -1350 41520 -1150 41590
rect -850 41520 -650 41590
rect -350 41520 -150 41590
rect 150 41520 350 41590
rect 650 41520 850 41590
rect 1150 41520 1350 41590
rect 1650 41520 1850 41590
rect 2150 41520 2350 41590
rect 2650 41520 2850 41590
rect 3150 41520 3350 41590
rect 3650 41520 3850 41590
rect -15850 41410 -15650 41480
rect -15350 41410 -15150 41480
rect -14850 41410 -14650 41480
rect -14350 41410 -14150 41480
rect -13850 41410 -13650 41480
rect -13350 41410 -13150 41480
rect -12850 41410 -12650 41480
rect -12350 41410 -12150 41480
rect -11850 41410 -11650 41480
rect -11350 41410 -11150 41480
rect -10850 41410 -10650 41480
rect -10350 41410 -10150 41480
rect -9850 41410 -9650 41480
rect -9350 41410 -9150 41480
rect -8850 41410 -8650 41480
rect -8350 41410 -8150 41480
rect -7850 41410 -7650 41480
rect -7350 41410 -7150 41480
rect -6850 41410 -6650 41480
rect -6350 41410 -6150 41480
rect -5850 41410 -5650 41480
rect -5350 41410 -5150 41480
rect -4850 41410 -4650 41480
rect -4350 41410 -4150 41480
rect -3850 41410 -3650 41480
rect -3350 41410 -3150 41480
rect -2850 41410 -2650 41480
rect -2350 41410 -2150 41480
rect -1850 41410 -1650 41480
rect -1350 41410 -1150 41480
rect -850 41410 -650 41480
rect -350 41410 -150 41480
rect 150 41410 350 41480
rect 650 41410 850 41480
rect 1150 41410 1350 41480
rect 1650 41410 1850 41480
rect 2150 41410 2350 41480
rect 2650 41410 2850 41480
rect 3150 41410 3350 41480
rect 3650 41410 3850 41480
rect -15980 41150 -15910 41350
rect -15590 41150 -15520 41350
rect -15480 41150 -15410 41350
rect -15090 41150 -15020 41350
rect -14980 41150 -14910 41350
rect -14590 41150 -14520 41350
rect -14480 41150 -14410 41350
rect -14090 41150 -14020 41350
rect -13980 41150 -13910 41350
rect -13590 41150 -13520 41350
rect -13480 41150 -13410 41350
rect -13090 41150 -13020 41350
rect -12980 41150 -12910 41350
rect -12590 41150 -12520 41350
rect -12480 41150 -12410 41350
rect -12090 41150 -12020 41350
rect -11980 41150 -11910 41350
rect -11590 41150 -11520 41350
rect -11480 41150 -11410 41350
rect -11090 41150 -11020 41350
rect -10980 41150 -10910 41350
rect -10590 41150 -10520 41350
rect -10480 41150 -10410 41350
rect -10090 41150 -10020 41350
rect -9980 41150 -9910 41350
rect -9590 41150 -9520 41350
rect -9480 41150 -9410 41350
rect -9090 41150 -9020 41350
rect -8980 41150 -8910 41350
rect -8590 41150 -8520 41350
rect -8480 41150 -8410 41350
rect -8090 41150 -8020 41350
rect -7980 41150 -7910 41350
rect -7590 41150 -7520 41350
rect -7480 41150 -7410 41350
rect -7090 41150 -7020 41350
rect -6980 41150 -6910 41350
rect -6590 41150 -6520 41350
rect -6480 41150 -6410 41350
rect -6090 41150 -6020 41350
rect -5980 41150 -5910 41350
rect -5590 41150 -5520 41350
rect -5480 41150 -5410 41350
rect -5090 41150 -5020 41350
rect -4980 41150 -4910 41350
rect -4590 41150 -4520 41350
rect -4480 41150 -4410 41350
rect -4090 41150 -4020 41350
rect -3980 41150 -3910 41350
rect -3590 41150 -3520 41350
rect -3480 41150 -3410 41350
rect -3090 41150 -3020 41350
rect -2980 41150 -2910 41350
rect -2590 41150 -2520 41350
rect -2480 41150 -2410 41350
rect -2090 41150 -2020 41350
rect -1980 41150 -1910 41350
rect -1590 41150 -1520 41350
rect -1480 41150 -1410 41350
rect -1090 41150 -1020 41350
rect -980 41150 -910 41350
rect -590 41150 -520 41350
rect -480 41150 -410 41350
rect -90 41150 -20 41350
rect 20 41150 90 41350
rect 410 41150 480 41350
rect 520 41150 590 41350
rect 910 41150 980 41350
rect 1020 41150 1090 41350
rect 1410 41150 1480 41350
rect 1520 41150 1590 41350
rect 1910 41150 1980 41350
rect 2020 41150 2090 41350
rect 2410 41150 2480 41350
rect 2520 41150 2590 41350
rect 2910 41150 2980 41350
rect 3020 41150 3090 41350
rect 3410 41150 3480 41350
rect 3520 41150 3590 41350
rect 3910 41150 3980 41350
rect -15850 41020 -15650 41090
rect -15350 41020 -15150 41090
rect -14850 41020 -14650 41090
rect -14350 41020 -14150 41090
rect -13850 41020 -13650 41090
rect -13350 41020 -13150 41090
rect -12850 41020 -12650 41090
rect -12350 41020 -12150 41090
rect -11850 41020 -11650 41090
rect -11350 41020 -11150 41090
rect -10850 41020 -10650 41090
rect -10350 41020 -10150 41090
rect -9850 41020 -9650 41090
rect -9350 41020 -9150 41090
rect -8850 41020 -8650 41090
rect -8350 41020 -8150 41090
rect -7850 41020 -7650 41090
rect -7350 41020 -7150 41090
rect -6850 41020 -6650 41090
rect -6350 41020 -6150 41090
rect -5850 41020 -5650 41090
rect -5350 41020 -5150 41090
rect -4850 41020 -4650 41090
rect -4350 41020 -4150 41090
rect -3850 41020 -3650 41090
rect -3350 41020 -3150 41090
rect -2850 41020 -2650 41090
rect -2350 41020 -2150 41090
rect -1850 41020 -1650 41090
rect -1350 41020 -1150 41090
rect -850 41020 -650 41090
rect -350 41020 -150 41090
rect 150 41020 350 41090
rect 650 41020 850 41090
rect 1150 41020 1350 41090
rect 1650 41020 1850 41090
rect 2150 41020 2350 41090
rect 2650 41020 2850 41090
rect 3150 41020 3350 41090
rect 3650 41020 3850 41090
rect -15850 40910 -15650 40980
rect -15350 40910 -15150 40980
rect -14850 40910 -14650 40980
rect -14350 40910 -14150 40980
rect -13850 40910 -13650 40980
rect -13350 40910 -13150 40980
rect -12850 40910 -12650 40980
rect -12350 40910 -12150 40980
rect -11850 40910 -11650 40980
rect -11350 40910 -11150 40980
rect -10850 40910 -10650 40980
rect -10350 40910 -10150 40980
rect -9850 40910 -9650 40980
rect -9350 40910 -9150 40980
rect -8850 40910 -8650 40980
rect -8350 40910 -8150 40980
rect -7850 40910 -7650 40980
rect -7350 40910 -7150 40980
rect -6850 40910 -6650 40980
rect -6350 40910 -6150 40980
rect -5850 40910 -5650 40980
rect -5350 40910 -5150 40980
rect -4850 40910 -4650 40980
rect -4350 40910 -4150 40980
rect -3850 40910 -3650 40980
rect -3350 40910 -3150 40980
rect -2850 40910 -2650 40980
rect -2350 40910 -2150 40980
rect -1850 40910 -1650 40980
rect -1350 40910 -1150 40980
rect -850 40910 -650 40980
rect -350 40910 -150 40980
rect 150 40910 350 40980
rect 650 40910 850 40980
rect 1150 40910 1350 40980
rect 1650 40910 1850 40980
rect 2150 40910 2350 40980
rect 2650 40910 2850 40980
rect 3150 40910 3350 40980
rect 3650 40910 3850 40980
rect -15980 40650 -15910 40850
rect -15590 40650 -15520 40850
rect -15480 40650 -15410 40850
rect -15090 40650 -15020 40850
rect -14980 40650 -14910 40850
rect -14590 40650 -14520 40850
rect -14480 40650 -14410 40850
rect -14090 40650 -14020 40850
rect -13980 40650 -13910 40850
rect -13590 40650 -13520 40850
rect -13480 40650 -13410 40850
rect -13090 40650 -13020 40850
rect -12980 40650 -12910 40850
rect -12590 40650 -12520 40850
rect -12480 40650 -12410 40850
rect -12090 40650 -12020 40850
rect -11980 40650 -11910 40850
rect -11590 40650 -11520 40850
rect -11480 40650 -11410 40850
rect -11090 40650 -11020 40850
rect -10980 40650 -10910 40850
rect -10590 40650 -10520 40850
rect -10480 40650 -10410 40850
rect -10090 40650 -10020 40850
rect -9980 40650 -9910 40850
rect -9590 40650 -9520 40850
rect -9480 40650 -9410 40850
rect -9090 40650 -9020 40850
rect -8980 40650 -8910 40850
rect -8590 40650 -8520 40850
rect -8480 40650 -8410 40850
rect -8090 40650 -8020 40850
rect -7980 40650 -7910 40850
rect -7590 40650 -7520 40850
rect -7480 40650 -7410 40850
rect -7090 40650 -7020 40850
rect -6980 40650 -6910 40850
rect -6590 40650 -6520 40850
rect -6480 40650 -6410 40850
rect -6090 40650 -6020 40850
rect -5980 40650 -5910 40850
rect -5590 40650 -5520 40850
rect -5480 40650 -5410 40850
rect -5090 40650 -5020 40850
rect -4980 40650 -4910 40850
rect -4590 40650 -4520 40850
rect -4480 40650 -4410 40850
rect -4090 40650 -4020 40850
rect -3980 40650 -3910 40850
rect -3590 40650 -3520 40850
rect -3480 40650 -3410 40850
rect -3090 40650 -3020 40850
rect -2980 40650 -2910 40850
rect -2590 40650 -2520 40850
rect -2480 40650 -2410 40850
rect -2090 40650 -2020 40850
rect -1980 40650 -1910 40850
rect -1590 40650 -1520 40850
rect -1480 40650 -1410 40850
rect -1090 40650 -1020 40850
rect -980 40650 -910 40850
rect -590 40650 -520 40850
rect -480 40650 -410 40850
rect -90 40650 -20 40850
rect 20 40650 90 40850
rect 410 40650 480 40850
rect 520 40650 590 40850
rect 910 40650 980 40850
rect 1020 40650 1090 40850
rect 1410 40650 1480 40850
rect 1520 40650 1590 40850
rect 1910 40650 1980 40850
rect 2020 40650 2090 40850
rect 2410 40650 2480 40850
rect 2520 40650 2590 40850
rect 2910 40650 2980 40850
rect 3020 40650 3090 40850
rect 3410 40650 3480 40850
rect 3520 40650 3590 40850
rect 3910 40650 3980 40850
rect -15850 40520 -15650 40590
rect -15350 40520 -15150 40590
rect -14850 40520 -14650 40590
rect -14350 40520 -14150 40590
rect -13850 40520 -13650 40590
rect -13350 40520 -13150 40590
rect -12850 40520 -12650 40590
rect -12350 40520 -12150 40590
rect -11850 40520 -11650 40590
rect -11350 40520 -11150 40590
rect -10850 40520 -10650 40590
rect -10350 40520 -10150 40590
rect -9850 40520 -9650 40590
rect -9350 40520 -9150 40590
rect -8850 40520 -8650 40590
rect -8350 40520 -8150 40590
rect -7850 40520 -7650 40590
rect -7350 40520 -7150 40590
rect -6850 40520 -6650 40590
rect -6350 40520 -6150 40590
rect -5850 40520 -5650 40590
rect -5350 40520 -5150 40590
rect -4850 40520 -4650 40590
rect -4350 40520 -4150 40590
rect -3850 40520 -3650 40590
rect -3350 40520 -3150 40590
rect -2850 40520 -2650 40590
rect -2350 40520 -2150 40590
rect -1850 40520 -1650 40590
rect -1350 40520 -1150 40590
rect -850 40520 -650 40590
rect -350 40520 -150 40590
rect 150 40520 350 40590
rect 650 40520 850 40590
rect 1150 40520 1350 40590
rect 1650 40520 1850 40590
rect 2150 40520 2350 40590
rect 2650 40520 2850 40590
rect 3150 40520 3350 40590
rect 3650 40520 3850 40590
rect -15850 40410 -15650 40480
rect -15350 40410 -15150 40480
rect -14850 40410 -14650 40480
rect -14350 40410 -14150 40480
rect -13850 40410 -13650 40480
rect -13350 40410 -13150 40480
rect -12850 40410 -12650 40480
rect -12350 40410 -12150 40480
rect -11850 40410 -11650 40480
rect -11350 40410 -11150 40480
rect -10850 40410 -10650 40480
rect -10350 40410 -10150 40480
rect -9850 40410 -9650 40480
rect -9350 40410 -9150 40480
rect -8850 40410 -8650 40480
rect -8350 40410 -8150 40480
rect -7850 40410 -7650 40480
rect -7350 40410 -7150 40480
rect -6850 40410 -6650 40480
rect -6350 40410 -6150 40480
rect -5850 40410 -5650 40480
rect -5350 40410 -5150 40480
rect -4850 40410 -4650 40480
rect -4350 40410 -4150 40480
rect -3850 40410 -3650 40480
rect -3350 40410 -3150 40480
rect -2850 40410 -2650 40480
rect -2350 40410 -2150 40480
rect -1850 40410 -1650 40480
rect -1350 40410 -1150 40480
rect -850 40410 -650 40480
rect -350 40410 -150 40480
rect 150 40410 350 40480
rect 650 40410 850 40480
rect 1150 40410 1350 40480
rect 1650 40410 1850 40480
rect 2150 40410 2350 40480
rect 2650 40410 2850 40480
rect 3150 40410 3350 40480
rect 3650 40410 3850 40480
rect -15980 40150 -15910 40350
rect -15590 40150 -15520 40350
rect -15480 40150 -15410 40350
rect -15090 40150 -15020 40350
rect -14980 40150 -14910 40350
rect -14590 40150 -14520 40350
rect -14480 40150 -14410 40350
rect -14090 40150 -14020 40350
rect -13980 40150 -13910 40350
rect -13590 40150 -13520 40350
rect -13480 40150 -13410 40350
rect -13090 40150 -13020 40350
rect -12980 40150 -12910 40350
rect -12590 40150 -12520 40350
rect -12480 40150 -12410 40350
rect -12090 40150 -12020 40350
rect -11980 40150 -11910 40350
rect -11590 40150 -11520 40350
rect -11480 40150 -11410 40350
rect -11090 40150 -11020 40350
rect -10980 40150 -10910 40350
rect -10590 40150 -10520 40350
rect -10480 40150 -10410 40350
rect -10090 40150 -10020 40350
rect -9980 40150 -9910 40350
rect -9590 40150 -9520 40350
rect -9480 40150 -9410 40350
rect -9090 40150 -9020 40350
rect -8980 40150 -8910 40350
rect -8590 40150 -8520 40350
rect -8480 40150 -8410 40350
rect -8090 40150 -8020 40350
rect -7980 40150 -7910 40350
rect -7590 40150 -7520 40350
rect -7480 40150 -7410 40350
rect -7090 40150 -7020 40350
rect -6980 40150 -6910 40350
rect -6590 40150 -6520 40350
rect -6480 40150 -6410 40350
rect -6090 40150 -6020 40350
rect -5980 40150 -5910 40350
rect -5590 40150 -5520 40350
rect -5480 40150 -5410 40350
rect -5090 40150 -5020 40350
rect -4980 40150 -4910 40350
rect -4590 40150 -4520 40350
rect -4480 40150 -4410 40350
rect -4090 40150 -4020 40350
rect -3980 40150 -3910 40350
rect -3590 40150 -3520 40350
rect -3480 40150 -3410 40350
rect -3090 40150 -3020 40350
rect -2980 40150 -2910 40350
rect -2590 40150 -2520 40350
rect -2480 40150 -2410 40350
rect -2090 40150 -2020 40350
rect -1980 40150 -1910 40350
rect -1590 40150 -1520 40350
rect -1480 40150 -1410 40350
rect -1090 40150 -1020 40350
rect -980 40150 -910 40350
rect -590 40150 -520 40350
rect -480 40150 -410 40350
rect -90 40150 -20 40350
rect 20 40150 90 40350
rect 410 40150 480 40350
rect 520 40150 590 40350
rect 910 40150 980 40350
rect 1020 40150 1090 40350
rect 1410 40150 1480 40350
rect 1520 40150 1590 40350
rect 1910 40150 1980 40350
rect 2020 40150 2090 40350
rect 2410 40150 2480 40350
rect 2520 40150 2590 40350
rect 2910 40150 2980 40350
rect 3020 40150 3090 40350
rect 3410 40150 3480 40350
rect 3520 40150 3590 40350
rect 3910 40150 3980 40350
rect -15850 40020 -15650 40090
rect -15350 40020 -15150 40090
rect -14850 40020 -14650 40090
rect -14350 40020 -14150 40090
rect -13850 40020 -13650 40090
rect -13350 40020 -13150 40090
rect -12850 40020 -12650 40090
rect -12350 40020 -12150 40090
rect -11850 40020 -11650 40090
rect -11350 40020 -11150 40090
rect -10850 40020 -10650 40090
rect -10350 40020 -10150 40090
rect -9850 40020 -9650 40090
rect -9350 40020 -9150 40090
rect -8850 40020 -8650 40090
rect -8350 40020 -8150 40090
rect -7850 40020 -7650 40090
rect -7350 40020 -7150 40090
rect -6850 40020 -6650 40090
rect -6350 40020 -6150 40090
rect -5850 40020 -5650 40090
rect -5350 40020 -5150 40090
rect -4850 40020 -4650 40090
rect -4350 40020 -4150 40090
rect -3850 40020 -3650 40090
rect -3350 40020 -3150 40090
rect -2850 40020 -2650 40090
rect -2350 40020 -2150 40090
rect -1850 40020 -1650 40090
rect -1350 40020 -1150 40090
rect -850 40020 -650 40090
rect -350 40020 -150 40090
rect 150 40020 350 40090
rect 650 40020 850 40090
rect 1150 40020 1350 40090
rect 1650 40020 1850 40090
rect 2150 40020 2350 40090
rect 2650 40020 2850 40090
rect 3150 40020 3350 40090
rect 3650 40020 3850 40090
rect -27850 39910 -27650 39980
rect -27350 39910 -27150 39980
rect -26850 39910 -26650 39980
rect -26350 39910 -26150 39980
rect -25850 39910 -25650 39980
rect -25350 39910 -25150 39980
rect -24850 39910 -24650 39980
rect -24350 39910 -24150 39980
rect -23850 39910 -23650 39980
rect -23350 39910 -23150 39980
rect -22850 39910 -22650 39980
rect -22350 39910 -22150 39980
rect -21850 39910 -21650 39980
rect -21350 39910 -21150 39980
rect -20850 39910 -20650 39980
rect -20350 39910 -20150 39980
rect -19850 39910 -19650 39980
rect -19350 39910 -19150 39980
rect -18850 39910 -18650 39980
rect -18350 39910 -18150 39980
rect -17850 39910 -17650 39980
rect -17350 39910 -17150 39980
rect -16850 39910 -16650 39980
rect -16350 39910 -16150 39980
rect -15850 39910 -15650 39980
rect -15350 39910 -15150 39980
rect -14850 39910 -14650 39980
rect -14350 39910 -14150 39980
rect -13850 39910 -13650 39980
rect -13350 39910 -13150 39980
rect -12850 39910 -12650 39980
rect -12350 39910 -12150 39980
rect -11850 39910 -11650 39980
rect -11350 39910 -11150 39980
rect -10850 39910 -10650 39980
rect -10350 39910 -10150 39980
rect -9850 39910 -9650 39980
rect -9350 39910 -9150 39980
rect -8850 39910 -8650 39980
rect -8350 39910 -8150 39980
rect -7850 39910 -7650 39980
rect -7350 39910 -7150 39980
rect -6850 39910 -6650 39980
rect -6350 39910 -6150 39980
rect -5850 39910 -5650 39980
rect -5350 39910 -5150 39980
rect -4850 39910 -4650 39980
rect -4350 39910 -4150 39980
rect -3850 39910 -3650 39980
rect -3350 39910 -3150 39980
rect -2850 39910 -2650 39980
rect -2350 39910 -2150 39980
rect -1850 39910 -1650 39980
rect -1350 39910 -1150 39980
rect -850 39910 -650 39980
rect -350 39910 -150 39980
rect 150 39910 350 39980
rect 650 39910 850 39980
rect 1150 39910 1350 39980
rect 1650 39910 1850 39980
rect 2150 39910 2350 39980
rect 2650 39910 2850 39980
rect 3150 39910 3350 39980
rect 3650 39910 3850 39980
rect -27980 39650 -27910 39850
rect -27590 39650 -27520 39850
rect -27480 39650 -27410 39850
rect -27090 39650 -27020 39850
rect -26980 39650 -26910 39850
rect -26590 39650 -26520 39850
rect -26480 39650 -26410 39850
rect -26090 39650 -26020 39850
rect -25980 39650 -25910 39850
rect -25590 39650 -25520 39850
rect -25480 39650 -25410 39850
rect -25090 39650 -25020 39850
rect -24980 39650 -24910 39850
rect -24590 39650 -24520 39850
rect -24480 39650 -24410 39850
rect -24090 39650 -24020 39850
rect -23980 39650 -23910 39850
rect -23590 39650 -23520 39850
rect -23480 39650 -23410 39850
rect -23090 39650 -23020 39850
rect -22980 39650 -22910 39850
rect -22590 39650 -22520 39850
rect -22480 39650 -22410 39850
rect -22090 39650 -22020 39850
rect -21980 39650 -21910 39850
rect -21590 39650 -21520 39850
rect -21480 39650 -21410 39850
rect -21090 39650 -21020 39850
rect -20980 39650 -20910 39850
rect -20590 39650 -20520 39850
rect -20480 39650 -20410 39850
rect -20090 39650 -20020 39850
rect -19980 39650 -19910 39850
rect -19590 39650 -19520 39850
rect -19480 39650 -19410 39850
rect -19090 39650 -19020 39850
rect -18980 39650 -18910 39850
rect -18590 39650 -18520 39850
rect -18480 39650 -18410 39850
rect -18090 39650 -18020 39850
rect -17980 39650 -17910 39850
rect -17590 39650 -17520 39850
rect -17480 39650 -17410 39850
rect -17090 39650 -17020 39850
rect -16980 39650 -16910 39850
rect -16590 39650 -16520 39850
rect -16480 39650 -16410 39850
rect -16090 39650 -16020 39850
rect -15980 39650 -15910 39850
rect -15590 39650 -15520 39850
rect -15480 39650 -15410 39850
rect -15090 39650 -15020 39850
rect -14980 39650 -14910 39850
rect -14590 39650 -14520 39850
rect -14480 39650 -14410 39850
rect -14090 39650 -14020 39850
rect -13980 39650 -13910 39850
rect -13590 39650 -13520 39850
rect -13480 39650 -13410 39850
rect -13090 39650 -13020 39850
rect -12980 39650 -12910 39850
rect -12590 39650 -12520 39850
rect -12480 39650 -12410 39850
rect -12090 39650 -12020 39850
rect -11980 39650 -11910 39850
rect -11590 39650 -11520 39850
rect -11480 39650 -11410 39850
rect -11090 39650 -11020 39850
rect -10980 39650 -10910 39850
rect -10590 39650 -10520 39850
rect -10480 39650 -10410 39850
rect -10090 39650 -10020 39850
rect -9980 39650 -9910 39850
rect -9590 39650 -9520 39850
rect -9480 39650 -9410 39850
rect -9090 39650 -9020 39850
rect -8980 39650 -8910 39850
rect -8590 39650 -8520 39850
rect -8480 39650 -8410 39850
rect -8090 39650 -8020 39850
rect -7980 39650 -7910 39850
rect -7590 39650 -7520 39850
rect -7480 39650 -7410 39850
rect -7090 39650 -7020 39850
rect -6980 39650 -6910 39850
rect -6590 39650 -6520 39850
rect -6480 39650 -6410 39850
rect -6090 39650 -6020 39850
rect -5980 39650 -5910 39850
rect -5590 39650 -5520 39850
rect -5480 39650 -5410 39850
rect -5090 39650 -5020 39850
rect -4980 39650 -4910 39850
rect -4590 39650 -4520 39850
rect -4480 39650 -4410 39850
rect -4090 39650 -4020 39850
rect -3980 39650 -3910 39850
rect -3590 39650 -3520 39850
rect -3480 39650 -3410 39850
rect -3090 39650 -3020 39850
rect -2980 39650 -2910 39850
rect -2590 39650 -2520 39850
rect -2480 39650 -2410 39850
rect -2090 39650 -2020 39850
rect -1980 39650 -1910 39850
rect -1590 39650 -1520 39850
rect -1480 39650 -1410 39850
rect -1090 39650 -1020 39850
rect -980 39650 -910 39850
rect -590 39650 -520 39850
rect -480 39650 -410 39850
rect -90 39650 -20 39850
rect 20 39650 90 39850
rect 410 39650 480 39850
rect 520 39650 590 39850
rect 910 39650 980 39850
rect 1020 39650 1090 39850
rect 1410 39650 1480 39850
rect 1520 39650 1590 39850
rect 1910 39650 1980 39850
rect 2020 39650 2090 39850
rect 2410 39650 2480 39850
rect 2520 39650 2590 39850
rect 2910 39650 2980 39850
rect 3020 39650 3090 39850
rect 3410 39650 3480 39850
rect 3520 39650 3590 39850
rect 3910 39650 3980 39850
rect -27850 39520 -27650 39590
rect -27350 39520 -27150 39590
rect -26850 39520 -26650 39590
rect -26350 39520 -26150 39590
rect -25850 39520 -25650 39590
rect -25350 39520 -25150 39590
rect -24850 39520 -24650 39590
rect -24350 39520 -24150 39590
rect -23850 39520 -23650 39590
rect -23350 39520 -23150 39590
rect -22850 39520 -22650 39590
rect -22350 39520 -22150 39590
rect -21850 39520 -21650 39590
rect -21350 39520 -21150 39590
rect -20850 39520 -20650 39590
rect -20350 39520 -20150 39590
rect -19850 39520 -19650 39590
rect -19350 39520 -19150 39590
rect -18850 39520 -18650 39590
rect -18350 39520 -18150 39590
rect -17850 39520 -17650 39590
rect -17350 39520 -17150 39590
rect -16850 39520 -16650 39590
rect -16350 39520 -16150 39590
rect -15850 39520 -15650 39590
rect -15350 39520 -15150 39590
rect -14850 39520 -14650 39590
rect -14350 39520 -14150 39590
rect -13850 39520 -13650 39590
rect -13350 39520 -13150 39590
rect -12850 39520 -12650 39590
rect -12350 39520 -12150 39590
rect -11850 39520 -11650 39590
rect -11350 39520 -11150 39590
rect -10850 39520 -10650 39590
rect -10350 39520 -10150 39590
rect -9850 39520 -9650 39590
rect -9350 39520 -9150 39590
rect -8850 39520 -8650 39590
rect -8350 39520 -8150 39590
rect -7850 39520 -7650 39590
rect -7350 39520 -7150 39590
rect -6850 39520 -6650 39590
rect -6350 39520 -6150 39590
rect -5850 39520 -5650 39590
rect -5350 39520 -5150 39590
rect -4850 39520 -4650 39590
rect -4350 39520 -4150 39590
rect -3850 39520 -3650 39590
rect -3350 39520 -3150 39590
rect -2850 39520 -2650 39590
rect -2350 39520 -2150 39590
rect -1850 39520 -1650 39590
rect -1350 39520 -1150 39590
rect -850 39520 -650 39590
rect -350 39520 -150 39590
rect 150 39520 350 39590
rect 650 39520 850 39590
rect 1150 39520 1350 39590
rect 1650 39520 1850 39590
rect 2150 39520 2350 39590
rect 2650 39520 2850 39590
rect 3150 39520 3350 39590
rect 3650 39520 3850 39590
rect -27850 39410 -27650 39480
rect -27350 39410 -27150 39480
rect -26850 39410 -26650 39480
rect -26350 39410 -26150 39480
rect -25850 39410 -25650 39480
rect -25350 39410 -25150 39480
rect -24850 39410 -24650 39480
rect -24350 39410 -24150 39480
rect -23850 39410 -23650 39480
rect -23350 39410 -23150 39480
rect -22850 39410 -22650 39480
rect -22350 39410 -22150 39480
rect -21850 39410 -21650 39480
rect -21350 39410 -21150 39480
rect -20850 39410 -20650 39480
rect -20350 39410 -20150 39480
rect -19850 39410 -19650 39480
rect -19350 39410 -19150 39480
rect -18850 39410 -18650 39480
rect -18350 39410 -18150 39480
rect -17850 39410 -17650 39480
rect -17350 39410 -17150 39480
rect -16850 39410 -16650 39480
rect -16350 39410 -16150 39480
rect -15850 39410 -15650 39480
rect -15350 39410 -15150 39480
rect -14850 39410 -14650 39480
rect -14350 39410 -14150 39480
rect -13850 39410 -13650 39480
rect -13350 39410 -13150 39480
rect -12850 39410 -12650 39480
rect -12350 39410 -12150 39480
rect -11850 39410 -11650 39480
rect -11350 39410 -11150 39480
rect -10850 39410 -10650 39480
rect -10350 39410 -10150 39480
rect -9850 39410 -9650 39480
rect -9350 39410 -9150 39480
rect -8850 39410 -8650 39480
rect -8350 39410 -8150 39480
rect -7850 39410 -7650 39480
rect -7350 39410 -7150 39480
rect -6850 39410 -6650 39480
rect -6350 39410 -6150 39480
rect -5850 39410 -5650 39480
rect -5350 39410 -5150 39480
rect -4850 39410 -4650 39480
rect -4350 39410 -4150 39480
rect -3850 39410 -3650 39480
rect -3350 39410 -3150 39480
rect -2850 39410 -2650 39480
rect -2350 39410 -2150 39480
rect -1850 39410 -1650 39480
rect -1350 39410 -1150 39480
rect -850 39410 -650 39480
rect -350 39410 -150 39480
rect 150 39410 350 39480
rect 650 39410 850 39480
rect 1150 39410 1350 39480
rect 1650 39410 1850 39480
rect 2150 39410 2350 39480
rect 2650 39410 2850 39480
rect 3150 39410 3350 39480
rect 3650 39410 3850 39480
rect -27980 39150 -27910 39350
rect -27590 39150 -27520 39350
rect -27480 39150 -27410 39350
rect -27090 39150 -27020 39350
rect -26980 39150 -26910 39350
rect -26590 39150 -26520 39350
rect -26480 39150 -26410 39350
rect -26090 39150 -26020 39350
rect -25980 39150 -25910 39350
rect -25590 39150 -25520 39350
rect -25480 39150 -25410 39350
rect -25090 39150 -25020 39350
rect -24980 39150 -24910 39350
rect -24590 39150 -24520 39350
rect -24480 39150 -24410 39350
rect -24090 39150 -24020 39350
rect -23980 39150 -23910 39350
rect -23590 39150 -23520 39350
rect -23480 39150 -23410 39350
rect -23090 39150 -23020 39350
rect -22980 39150 -22910 39350
rect -22590 39150 -22520 39350
rect -22480 39150 -22410 39350
rect -22090 39150 -22020 39350
rect -21980 39150 -21910 39350
rect -21590 39150 -21520 39350
rect -21480 39150 -21410 39350
rect -21090 39150 -21020 39350
rect -20980 39150 -20910 39350
rect -20590 39150 -20520 39350
rect -20480 39150 -20410 39350
rect -20090 39150 -20020 39350
rect -19980 39150 -19910 39350
rect -19590 39150 -19520 39350
rect -19480 39150 -19410 39350
rect -19090 39150 -19020 39350
rect -18980 39150 -18910 39350
rect -18590 39150 -18520 39350
rect -18480 39150 -18410 39350
rect -18090 39150 -18020 39350
rect -17980 39150 -17910 39350
rect -17590 39150 -17520 39350
rect -17480 39150 -17410 39350
rect -17090 39150 -17020 39350
rect -16980 39150 -16910 39350
rect -16590 39150 -16520 39350
rect -16480 39150 -16410 39350
rect -16090 39150 -16020 39350
rect -15980 39150 -15910 39350
rect -15590 39150 -15520 39350
rect -15480 39150 -15410 39350
rect -15090 39150 -15020 39350
rect -14980 39150 -14910 39350
rect -14590 39150 -14520 39350
rect -14480 39150 -14410 39350
rect -14090 39150 -14020 39350
rect -13980 39150 -13910 39350
rect -13590 39150 -13520 39350
rect -13480 39150 -13410 39350
rect -13090 39150 -13020 39350
rect -12980 39150 -12910 39350
rect -12590 39150 -12520 39350
rect -12480 39150 -12410 39350
rect -12090 39150 -12020 39350
rect -11980 39150 -11910 39350
rect -11590 39150 -11520 39350
rect -11480 39150 -11410 39350
rect -11090 39150 -11020 39350
rect -10980 39150 -10910 39350
rect -10590 39150 -10520 39350
rect -10480 39150 -10410 39350
rect -10090 39150 -10020 39350
rect -9980 39150 -9910 39350
rect -9590 39150 -9520 39350
rect -9480 39150 -9410 39350
rect -9090 39150 -9020 39350
rect -8980 39150 -8910 39350
rect -8590 39150 -8520 39350
rect -8480 39150 -8410 39350
rect -8090 39150 -8020 39350
rect -7980 39150 -7910 39350
rect -7590 39150 -7520 39350
rect -7480 39150 -7410 39350
rect -7090 39150 -7020 39350
rect -6980 39150 -6910 39350
rect -6590 39150 -6520 39350
rect -6480 39150 -6410 39350
rect -6090 39150 -6020 39350
rect -5980 39150 -5910 39350
rect -5590 39150 -5520 39350
rect -5480 39150 -5410 39350
rect -5090 39150 -5020 39350
rect -4980 39150 -4910 39350
rect -4590 39150 -4520 39350
rect -4480 39150 -4410 39350
rect -4090 39150 -4020 39350
rect -3980 39150 -3910 39350
rect -3590 39150 -3520 39350
rect -3480 39150 -3410 39350
rect -3090 39150 -3020 39350
rect -2980 39150 -2910 39350
rect -2590 39150 -2520 39350
rect -2480 39150 -2410 39350
rect -2090 39150 -2020 39350
rect -1980 39150 -1910 39350
rect -1590 39150 -1520 39350
rect -1480 39150 -1410 39350
rect -1090 39150 -1020 39350
rect -980 39150 -910 39350
rect -590 39150 -520 39350
rect -480 39150 -410 39350
rect -90 39150 -20 39350
rect 20 39150 90 39350
rect 410 39150 480 39350
rect 520 39150 590 39350
rect 910 39150 980 39350
rect 1020 39150 1090 39350
rect 1410 39150 1480 39350
rect 1520 39150 1590 39350
rect 1910 39150 1980 39350
rect 2020 39150 2090 39350
rect 2410 39150 2480 39350
rect 2520 39150 2590 39350
rect 2910 39150 2980 39350
rect 3020 39150 3090 39350
rect 3410 39150 3480 39350
rect 3520 39150 3590 39350
rect 3910 39150 3980 39350
rect -27850 39020 -27650 39090
rect -27350 39020 -27150 39090
rect -26850 39020 -26650 39090
rect -26350 39020 -26150 39090
rect -25850 39020 -25650 39090
rect -25350 39020 -25150 39090
rect -24850 39020 -24650 39090
rect -24350 39020 -24150 39090
rect -23850 39020 -23650 39090
rect -23350 39020 -23150 39090
rect -22850 39020 -22650 39090
rect -22350 39020 -22150 39090
rect -21850 39020 -21650 39090
rect -21350 39020 -21150 39090
rect -20850 39020 -20650 39090
rect -20350 39020 -20150 39090
rect -19850 39020 -19650 39090
rect -19350 39020 -19150 39090
rect -18850 39020 -18650 39090
rect -18350 39020 -18150 39090
rect -17850 39020 -17650 39090
rect -17350 39020 -17150 39090
rect -16850 39020 -16650 39090
rect -16350 39020 -16150 39090
rect -15850 39020 -15650 39090
rect -15350 39020 -15150 39090
rect -14850 39020 -14650 39090
rect -14350 39020 -14150 39090
rect -13850 39020 -13650 39090
rect -13350 39020 -13150 39090
rect -12850 39020 -12650 39090
rect -12350 39020 -12150 39090
rect -11850 39020 -11650 39090
rect -11350 39020 -11150 39090
rect -10850 39020 -10650 39090
rect -10350 39020 -10150 39090
rect -9850 39020 -9650 39090
rect -9350 39020 -9150 39090
rect -8850 39020 -8650 39090
rect -8350 39020 -8150 39090
rect -7850 39020 -7650 39090
rect -7350 39020 -7150 39090
rect -6850 39020 -6650 39090
rect -6350 39020 -6150 39090
rect -5850 39020 -5650 39090
rect -5350 39020 -5150 39090
rect -4850 39020 -4650 39090
rect -4350 39020 -4150 39090
rect -3850 39020 -3650 39090
rect -3350 39020 -3150 39090
rect -2850 39020 -2650 39090
rect -2350 39020 -2150 39090
rect -1850 39020 -1650 39090
rect -1350 39020 -1150 39090
rect -850 39020 -650 39090
rect -350 39020 -150 39090
rect 150 39020 350 39090
rect 650 39020 850 39090
rect 1150 39020 1350 39090
rect 1650 39020 1850 39090
rect 2150 39020 2350 39090
rect 2650 39020 2850 39090
rect 3150 39020 3350 39090
rect 3650 39020 3850 39090
rect -27850 38910 -27650 38980
rect -27350 38910 -27150 38980
rect -26850 38910 -26650 38980
rect -26350 38910 -26150 38980
rect -25850 38910 -25650 38980
rect -25350 38910 -25150 38980
rect -24850 38910 -24650 38980
rect -24350 38910 -24150 38980
rect -23850 38910 -23650 38980
rect -23350 38910 -23150 38980
rect -22850 38910 -22650 38980
rect -22350 38910 -22150 38980
rect -21850 38910 -21650 38980
rect -21350 38910 -21150 38980
rect -20850 38910 -20650 38980
rect -20350 38910 -20150 38980
rect -19850 38910 -19650 38980
rect -19350 38910 -19150 38980
rect -18850 38910 -18650 38980
rect -18350 38910 -18150 38980
rect -17850 38910 -17650 38980
rect -17350 38910 -17150 38980
rect -16850 38910 -16650 38980
rect -16350 38910 -16150 38980
rect -15850 38910 -15650 38980
rect -15350 38910 -15150 38980
rect -14850 38910 -14650 38980
rect -14350 38910 -14150 38980
rect -13850 38910 -13650 38980
rect -13350 38910 -13150 38980
rect -12850 38910 -12650 38980
rect -12350 38910 -12150 38980
rect -11850 38910 -11650 38980
rect -11350 38910 -11150 38980
rect -10850 38910 -10650 38980
rect -10350 38910 -10150 38980
rect -9850 38910 -9650 38980
rect -9350 38910 -9150 38980
rect -8850 38910 -8650 38980
rect -8350 38910 -8150 38980
rect -7850 38910 -7650 38980
rect -7350 38910 -7150 38980
rect -6850 38910 -6650 38980
rect -6350 38910 -6150 38980
rect -5850 38910 -5650 38980
rect -5350 38910 -5150 38980
rect -4850 38910 -4650 38980
rect -4350 38910 -4150 38980
rect -3850 38910 -3650 38980
rect -3350 38910 -3150 38980
rect -2850 38910 -2650 38980
rect -2350 38910 -2150 38980
rect -1850 38910 -1650 38980
rect -1350 38910 -1150 38980
rect -850 38910 -650 38980
rect -350 38910 -150 38980
rect 150 38910 350 38980
rect 650 38910 850 38980
rect 1150 38910 1350 38980
rect 1650 38910 1850 38980
rect 2150 38910 2350 38980
rect 2650 38910 2850 38980
rect 3150 38910 3350 38980
rect 3650 38910 3850 38980
rect -27980 38650 -27910 38850
rect -27590 38650 -27520 38850
rect -27480 38650 -27410 38850
rect -27090 38650 -27020 38850
rect -26980 38650 -26910 38850
rect -26590 38650 -26520 38850
rect -26480 38650 -26410 38850
rect -26090 38650 -26020 38850
rect -25980 38650 -25910 38850
rect -25590 38650 -25520 38850
rect -25480 38650 -25410 38850
rect -25090 38650 -25020 38850
rect -24980 38650 -24910 38850
rect -24590 38650 -24520 38850
rect -24480 38650 -24410 38850
rect -24090 38650 -24020 38850
rect -23980 38650 -23910 38850
rect -23590 38650 -23520 38850
rect -23480 38650 -23410 38850
rect -23090 38650 -23020 38850
rect -22980 38650 -22910 38850
rect -22590 38650 -22520 38850
rect -22480 38650 -22410 38850
rect -22090 38650 -22020 38850
rect -21980 38650 -21910 38850
rect -21590 38650 -21520 38850
rect -21480 38650 -21410 38850
rect -21090 38650 -21020 38850
rect -20980 38650 -20910 38850
rect -20590 38650 -20520 38850
rect -20480 38650 -20410 38850
rect -20090 38650 -20020 38850
rect -19980 38650 -19910 38850
rect -19590 38650 -19520 38850
rect -19480 38650 -19410 38850
rect -19090 38650 -19020 38850
rect -18980 38650 -18910 38850
rect -18590 38650 -18520 38850
rect -18480 38650 -18410 38850
rect -18090 38650 -18020 38850
rect -17980 38650 -17910 38850
rect -17590 38650 -17520 38850
rect -17480 38650 -17410 38850
rect -17090 38650 -17020 38850
rect -16980 38650 -16910 38850
rect -16590 38650 -16520 38850
rect -16480 38650 -16410 38850
rect -16090 38650 -16020 38850
rect -15980 38650 -15910 38850
rect -15590 38650 -15520 38850
rect -15480 38650 -15410 38850
rect -15090 38650 -15020 38850
rect -14980 38650 -14910 38850
rect -14590 38650 -14520 38850
rect -14480 38650 -14410 38850
rect -14090 38650 -14020 38850
rect -13980 38650 -13910 38850
rect -13590 38650 -13520 38850
rect -13480 38650 -13410 38850
rect -13090 38650 -13020 38850
rect -12980 38650 -12910 38850
rect -12590 38650 -12520 38850
rect -12480 38650 -12410 38850
rect -12090 38650 -12020 38850
rect -11980 38650 -11910 38850
rect -11590 38650 -11520 38850
rect -11480 38650 -11410 38850
rect -11090 38650 -11020 38850
rect -10980 38650 -10910 38850
rect -10590 38650 -10520 38850
rect -10480 38650 -10410 38850
rect -10090 38650 -10020 38850
rect -9980 38650 -9910 38850
rect -9590 38650 -9520 38850
rect -9480 38650 -9410 38850
rect -9090 38650 -9020 38850
rect -8980 38650 -8910 38850
rect -8590 38650 -8520 38850
rect -8480 38650 -8410 38850
rect -8090 38650 -8020 38850
rect -7980 38650 -7910 38850
rect -7590 38650 -7520 38850
rect -7480 38650 -7410 38850
rect -7090 38650 -7020 38850
rect -6980 38650 -6910 38850
rect -6590 38650 -6520 38850
rect -6480 38650 -6410 38850
rect -6090 38650 -6020 38850
rect -5980 38650 -5910 38850
rect -5590 38650 -5520 38850
rect -5480 38650 -5410 38850
rect -5090 38650 -5020 38850
rect -4980 38650 -4910 38850
rect -4590 38650 -4520 38850
rect -4480 38650 -4410 38850
rect -4090 38650 -4020 38850
rect -3980 38650 -3910 38850
rect -3590 38650 -3520 38850
rect -3480 38650 -3410 38850
rect -3090 38650 -3020 38850
rect -2980 38650 -2910 38850
rect -2590 38650 -2520 38850
rect -2480 38650 -2410 38850
rect -2090 38650 -2020 38850
rect -1980 38650 -1910 38850
rect -1590 38650 -1520 38850
rect -1480 38650 -1410 38850
rect -1090 38650 -1020 38850
rect -980 38650 -910 38850
rect -590 38650 -520 38850
rect -480 38650 -410 38850
rect -90 38650 -20 38850
rect 20 38650 90 38850
rect 410 38650 480 38850
rect 520 38650 590 38850
rect 910 38650 980 38850
rect 1020 38650 1090 38850
rect 1410 38650 1480 38850
rect 1520 38650 1590 38850
rect 1910 38650 1980 38850
rect 2020 38650 2090 38850
rect 2410 38650 2480 38850
rect 2520 38650 2590 38850
rect 2910 38650 2980 38850
rect 3020 38650 3090 38850
rect 3410 38650 3480 38850
rect 3520 38650 3590 38850
rect 3910 38650 3980 38850
rect -27850 38520 -27650 38590
rect -27350 38520 -27150 38590
rect -26850 38520 -26650 38590
rect -26350 38520 -26150 38590
rect -25850 38520 -25650 38590
rect -25350 38520 -25150 38590
rect -24850 38520 -24650 38590
rect -24350 38520 -24150 38590
rect -23850 38520 -23650 38590
rect -23350 38520 -23150 38590
rect -22850 38520 -22650 38590
rect -22350 38520 -22150 38590
rect -21850 38520 -21650 38590
rect -21350 38520 -21150 38590
rect -20850 38520 -20650 38590
rect -20350 38520 -20150 38590
rect -19850 38520 -19650 38590
rect -19350 38520 -19150 38590
rect -18850 38520 -18650 38590
rect -18350 38520 -18150 38590
rect -17850 38520 -17650 38590
rect -17350 38520 -17150 38590
rect -16850 38520 -16650 38590
rect -16350 38520 -16150 38590
rect -15850 38520 -15650 38590
rect -15350 38520 -15150 38590
rect -14850 38520 -14650 38590
rect -14350 38520 -14150 38590
rect -13850 38520 -13650 38590
rect -13350 38520 -13150 38590
rect -12850 38520 -12650 38590
rect -12350 38520 -12150 38590
rect -11850 38520 -11650 38590
rect -11350 38520 -11150 38590
rect -10850 38520 -10650 38590
rect -10350 38520 -10150 38590
rect -9850 38520 -9650 38590
rect -9350 38520 -9150 38590
rect -8850 38520 -8650 38590
rect -8350 38520 -8150 38590
rect -7850 38520 -7650 38590
rect -7350 38520 -7150 38590
rect -6850 38520 -6650 38590
rect -6350 38520 -6150 38590
rect -5850 38520 -5650 38590
rect -5350 38520 -5150 38590
rect -4850 38520 -4650 38590
rect -4350 38520 -4150 38590
rect -3850 38520 -3650 38590
rect -3350 38520 -3150 38590
rect -2850 38520 -2650 38590
rect -2350 38520 -2150 38590
rect -1850 38520 -1650 38590
rect -1350 38520 -1150 38590
rect -850 38520 -650 38590
rect -350 38520 -150 38590
rect 150 38520 350 38590
rect 650 38520 850 38590
rect 1150 38520 1350 38590
rect 1650 38520 1850 38590
rect 2150 38520 2350 38590
rect 2650 38520 2850 38590
rect 3150 38520 3350 38590
rect 3650 38520 3850 38590
rect -27850 38410 -27650 38480
rect -27350 38410 -27150 38480
rect -26850 38410 -26650 38480
rect -26350 38410 -26150 38480
rect -25850 38410 -25650 38480
rect -25350 38410 -25150 38480
rect -24850 38410 -24650 38480
rect -24350 38410 -24150 38480
rect -23850 38410 -23650 38480
rect -23350 38410 -23150 38480
rect -22850 38410 -22650 38480
rect -22350 38410 -22150 38480
rect -21850 38410 -21650 38480
rect -21350 38410 -21150 38480
rect -20850 38410 -20650 38480
rect -20350 38410 -20150 38480
rect -19850 38410 -19650 38480
rect -19350 38410 -19150 38480
rect -18850 38410 -18650 38480
rect -18350 38410 -18150 38480
rect -17850 38410 -17650 38480
rect -17350 38410 -17150 38480
rect -16850 38410 -16650 38480
rect -16350 38410 -16150 38480
rect -15850 38410 -15650 38480
rect -15350 38410 -15150 38480
rect -14850 38410 -14650 38480
rect -14350 38410 -14150 38480
rect -13850 38410 -13650 38480
rect -13350 38410 -13150 38480
rect -12850 38410 -12650 38480
rect -12350 38410 -12150 38480
rect -11850 38410 -11650 38480
rect -11350 38410 -11150 38480
rect -10850 38410 -10650 38480
rect -10350 38410 -10150 38480
rect -9850 38410 -9650 38480
rect -9350 38410 -9150 38480
rect -8850 38410 -8650 38480
rect -8350 38410 -8150 38480
rect -7850 38410 -7650 38480
rect -7350 38410 -7150 38480
rect -6850 38410 -6650 38480
rect -6350 38410 -6150 38480
rect -5850 38410 -5650 38480
rect -5350 38410 -5150 38480
rect -4850 38410 -4650 38480
rect -4350 38410 -4150 38480
rect -3850 38410 -3650 38480
rect -3350 38410 -3150 38480
rect -2850 38410 -2650 38480
rect -2350 38410 -2150 38480
rect -1850 38410 -1650 38480
rect -1350 38410 -1150 38480
rect -850 38410 -650 38480
rect -350 38410 -150 38480
rect 150 38410 350 38480
rect 650 38410 850 38480
rect 1150 38410 1350 38480
rect 1650 38410 1850 38480
rect 2150 38410 2350 38480
rect 2650 38410 2850 38480
rect 3150 38410 3350 38480
rect 3650 38410 3850 38480
rect -27980 38150 -27910 38350
rect -27590 38150 -27520 38350
rect -27480 38150 -27410 38350
rect -27090 38150 -27020 38350
rect -26980 38150 -26910 38350
rect -26590 38150 -26520 38350
rect -26480 38150 -26410 38350
rect -26090 38150 -26020 38350
rect -25980 38150 -25910 38350
rect -25590 38150 -25520 38350
rect -25480 38150 -25410 38350
rect -25090 38150 -25020 38350
rect -24980 38150 -24910 38350
rect -24590 38150 -24520 38350
rect -24480 38150 -24410 38350
rect -24090 38150 -24020 38350
rect -23980 38150 -23910 38350
rect -23590 38150 -23520 38350
rect -23480 38150 -23410 38350
rect -23090 38150 -23020 38350
rect -22980 38150 -22910 38350
rect -22590 38150 -22520 38350
rect -22480 38150 -22410 38350
rect -22090 38150 -22020 38350
rect -21980 38150 -21910 38350
rect -21590 38150 -21520 38350
rect -21480 38150 -21410 38350
rect -21090 38150 -21020 38350
rect -20980 38150 -20910 38350
rect -20590 38150 -20520 38350
rect -20480 38150 -20410 38350
rect -20090 38150 -20020 38350
rect -19980 38150 -19910 38350
rect -19590 38150 -19520 38350
rect -19480 38150 -19410 38350
rect -19090 38150 -19020 38350
rect -18980 38150 -18910 38350
rect -18590 38150 -18520 38350
rect -18480 38150 -18410 38350
rect -18090 38150 -18020 38350
rect -17980 38150 -17910 38350
rect -17590 38150 -17520 38350
rect -17480 38150 -17410 38350
rect -17090 38150 -17020 38350
rect -16980 38150 -16910 38350
rect -16590 38150 -16520 38350
rect -16480 38150 -16410 38350
rect -16090 38150 -16020 38350
rect -15980 38150 -15910 38350
rect -15590 38150 -15520 38350
rect -15480 38150 -15410 38350
rect -15090 38150 -15020 38350
rect -14980 38150 -14910 38350
rect -14590 38150 -14520 38350
rect -14480 38150 -14410 38350
rect -14090 38150 -14020 38350
rect -13980 38150 -13910 38350
rect -13590 38150 -13520 38350
rect -13480 38150 -13410 38350
rect -13090 38150 -13020 38350
rect -12980 38150 -12910 38350
rect -12590 38150 -12520 38350
rect -12480 38150 -12410 38350
rect -12090 38150 -12020 38350
rect -11980 38150 -11910 38350
rect -11590 38150 -11520 38350
rect -11480 38150 -11410 38350
rect -11090 38150 -11020 38350
rect -10980 38150 -10910 38350
rect -10590 38150 -10520 38350
rect -10480 38150 -10410 38350
rect -10090 38150 -10020 38350
rect -9980 38150 -9910 38350
rect -9590 38150 -9520 38350
rect -9480 38150 -9410 38350
rect -9090 38150 -9020 38350
rect -8980 38150 -8910 38350
rect -8590 38150 -8520 38350
rect -8480 38150 -8410 38350
rect -8090 38150 -8020 38350
rect -7980 38150 -7910 38350
rect -7590 38150 -7520 38350
rect -7480 38150 -7410 38350
rect -7090 38150 -7020 38350
rect -6980 38150 -6910 38350
rect -6590 38150 -6520 38350
rect -6480 38150 -6410 38350
rect -6090 38150 -6020 38350
rect -5980 38150 -5910 38350
rect -5590 38150 -5520 38350
rect -5480 38150 -5410 38350
rect -5090 38150 -5020 38350
rect -4980 38150 -4910 38350
rect -4590 38150 -4520 38350
rect -4480 38150 -4410 38350
rect -4090 38150 -4020 38350
rect -3980 38150 -3910 38350
rect -3590 38150 -3520 38350
rect -3480 38150 -3410 38350
rect -3090 38150 -3020 38350
rect -2980 38150 -2910 38350
rect -2590 38150 -2520 38350
rect -2480 38150 -2410 38350
rect -2090 38150 -2020 38350
rect -1980 38150 -1910 38350
rect -1590 38150 -1520 38350
rect -1480 38150 -1410 38350
rect -1090 38150 -1020 38350
rect -980 38150 -910 38350
rect -590 38150 -520 38350
rect -480 38150 -410 38350
rect -90 38150 -20 38350
rect 20 38150 90 38350
rect 410 38150 480 38350
rect 520 38150 590 38350
rect 910 38150 980 38350
rect 1020 38150 1090 38350
rect 1410 38150 1480 38350
rect 1520 38150 1590 38350
rect 1910 38150 1980 38350
rect 2020 38150 2090 38350
rect 2410 38150 2480 38350
rect 2520 38150 2590 38350
rect 2910 38150 2980 38350
rect 3020 38150 3090 38350
rect 3410 38150 3480 38350
rect 3520 38150 3590 38350
rect 3910 38150 3980 38350
rect -27850 38020 -27650 38090
rect -27350 38020 -27150 38090
rect -26850 38020 -26650 38090
rect -26350 38020 -26150 38090
rect -25850 38020 -25650 38090
rect -25350 38020 -25150 38090
rect -24850 38020 -24650 38090
rect -24350 38020 -24150 38090
rect -23850 38020 -23650 38090
rect -23350 38020 -23150 38090
rect -22850 38020 -22650 38090
rect -22350 38020 -22150 38090
rect -21850 38020 -21650 38090
rect -21350 38020 -21150 38090
rect -20850 38020 -20650 38090
rect -20350 38020 -20150 38090
rect -19850 38020 -19650 38090
rect -19350 38020 -19150 38090
rect -18850 38020 -18650 38090
rect -18350 38020 -18150 38090
rect -17850 38020 -17650 38090
rect -17350 38020 -17150 38090
rect -16850 38020 -16650 38090
rect -16350 38020 -16150 38090
rect -15850 38020 -15650 38090
rect -15350 38020 -15150 38090
rect -14850 38020 -14650 38090
rect -14350 38020 -14150 38090
rect -13850 38020 -13650 38090
rect -13350 38020 -13150 38090
rect -12850 38020 -12650 38090
rect -12350 38020 -12150 38090
rect -11850 38020 -11650 38090
rect -11350 38020 -11150 38090
rect -10850 38020 -10650 38090
rect -10350 38020 -10150 38090
rect -9850 38020 -9650 38090
rect -9350 38020 -9150 38090
rect -8850 38020 -8650 38090
rect -8350 38020 -8150 38090
rect -7850 38020 -7650 38090
rect -7350 38020 -7150 38090
rect -6850 38020 -6650 38090
rect -6350 38020 -6150 38090
rect -5850 38020 -5650 38090
rect -5350 38020 -5150 38090
rect -4850 38020 -4650 38090
rect -4350 38020 -4150 38090
rect -3850 38020 -3650 38090
rect -3350 38020 -3150 38090
rect -2850 38020 -2650 38090
rect -2350 38020 -2150 38090
rect -1850 38020 -1650 38090
rect -1350 38020 -1150 38090
rect -850 38020 -650 38090
rect -350 38020 -150 38090
rect 150 38020 350 38090
rect 650 38020 850 38090
rect 1150 38020 1350 38090
rect 1650 38020 1850 38090
rect 2150 38020 2350 38090
rect 2650 38020 2850 38090
rect 3150 38020 3350 38090
rect 3650 38020 3850 38090
rect 128150 10910 128350 10980
rect 128650 10910 128850 10980
rect 129150 10910 129350 10980
rect 129650 10910 129850 10980
rect 130150 10910 130350 10980
rect 130650 10910 130850 10980
rect 131150 10910 131350 10980
rect 131650 10910 131850 10980
rect 132150 10910 132350 10980
rect 132650 10910 132850 10980
rect 133150 10910 133350 10980
rect 133650 10910 133850 10980
rect 134150 10910 134350 10980
rect 134650 10910 134850 10980
rect 135150 10910 135350 10980
rect 135650 10910 135850 10980
rect 136150 10910 136350 10980
rect 136650 10910 136850 10980
rect 137150 10910 137350 10980
rect 137650 10910 137850 10980
rect 138150 10910 138350 10980
rect 138650 10910 138850 10980
rect 139150 10910 139350 10980
rect 139650 10910 139850 10980
rect 128020 10650 128090 10850
rect 128410 10650 128480 10850
rect 128520 10650 128590 10850
rect 128910 10650 128980 10850
rect 129020 10650 129090 10850
rect 129410 10650 129480 10850
rect 129520 10650 129590 10850
rect 129910 10650 129980 10850
rect 130020 10650 130090 10850
rect 130410 10650 130480 10850
rect 130520 10650 130590 10850
rect 130910 10650 130980 10850
rect 131020 10650 131090 10850
rect 131410 10650 131480 10850
rect 131520 10650 131590 10850
rect 131910 10650 131980 10850
rect 132020 10650 132090 10850
rect 132410 10650 132480 10850
rect 132520 10650 132590 10850
rect 132910 10650 132980 10850
rect 133020 10650 133090 10850
rect 133410 10650 133480 10850
rect 133520 10650 133590 10850
rect 133910 10650 133980 10850
rect 134020 10650 134090 10850
rect 134410 10650 134480 10850
rect 134520 10650 134590 10850
rect 134910 10650 134980 10850
rect 135020 10650 135090 10850
rect 135410 10650 135480 10850
rect 135520 10650 135590 10850
rect 135910 10650 135980 10850
rect 136020 10650 136090 10850
rect 136410 10650 136480 10850
rect 136520 10650 136590 10850
rect 136910 10650 136980 10850
rect 137020 10650 137090 10850
rect 137410 10650 137480 10850
rect 137520 10650 137590 10850
rect 137910 10650 137980 10850
rect 138020 10650 138090 10850
rect 138410 10650 138480 10850
rect 138520 10650 138590 10850
rect 138910 10650 138980 10850
rect 139020 10650 139090 10850
rect 139410 10650 139480 10850
rect 139520 10650 139590 10850
rect 139910 10650 139980 10850
rect 128150 10520 128350 10590
rect 128650 10520 128850 10590
rect 129150 10520 129350 10590
rect 129650 10520 129850 10590
rect 130150 10520 130350 10590
rect 130650 10520 130850 10590
rect 131150 10520 131350 10590
rect 131650 10520 131850 10590
rect 132150 10520 132350 10590
rect 132650 10520 132850 10590
rect 133150 10520 133350 10590
rect 133650 10520 133850 10590
rect 134150 10520 134350 10590
rect 134650 10520 134850 10590
rect 135150 10520 135350 10590
rect 135650 10520 135850 10590
rect 136150 10520 136350 10590
rect 136650 10520 136850 10590
rect 137150 10520 137350 10590
rect 137650 10520 137850 10590
rect 138150 10520 138350 10590
rect 138650 10520 138850 10590
rect 139150 10520 139350 10590
rect 139650 10520 139850 10590
rect 128150 10410 128350 10480
rect 128650 10410 128850 10480
rect 129150 10410 129350 10480
rect 129650 10410 129850 10480
rect 130150 10410 130350 10480
rect 130650 10410 130850 10480
rect 131150 10410 131350 10480
rect 131650 10410 131850 10480
rect 132150 10410 132350 10480
rect 132650 10410 132850 10480
rect 133150 10410 133350 10480
rect 133650 10410 133850 10480
rect 134150 10410 134350 10480
rect 134650 10410 134850 10480
rect 135150 10410 135350 10480
rect 135650 10410 135850 10480
rect 136150 10410 136350 10480
rect 136650 10410 136850 10480
rect 137150 10410 137350 10480
rect 137650 10410 137850 10480
rect 138150 10410 138350 10480
rect 138650 10410 138850 10480
rect 139150 10410 139350 10480
rect 139650 10410 139850 10480
rect 128020 10150 128090 10350
rect 128410 10150 128480 10350
rect 128520 10150 128590 10350
rect 128910 10150 128980 10350
rect 129020 10150 129090 10350
rect 129410 10150 129480 10350
rect 129520 10150 129590 10350
rect 129910 10150 129980 10350
rect 130020 10150 130090 10350
rect 130410 10150 130480 10350
rect 130520 10150 130590 10350
rect 130910 10150 130980 10350
rect 131020 10150 131090 10350
rect 131410 10150 131480 10350
rect 131520 10150 131590 10350
rect 131910 10150 131980 10350
rect 132020 10150 132090 10350
rect 132410 10150 132480 10350
rect 132520 10150 132590 10350
rect 132910 10150 132980 10350
rect 133020 10150 133090 10350
rect 133410 10150 133480 10350
rect 133520 10150 133590 10350
rect 133910 10150 133980 10350
rect 134020 10150 134090 10350
rect 134410 10150 134480 10350
rect 134520 10150 134590 10350
rect 134910 10150 134980 10350
rect 135020 10150 135090 10350
rect 135410 10150 135480 10350
rect 135520 10150 135590 10350
rect 135910 10150 135980 10350
rect 136020 10150 136090 10350
rect 136410 10150 136480 10350
rect 136520 10150 136590 10350
rect 136910 10150 136980 10350
rect 137020 10150 137090 10350
rect 137410 10150 137480 10350
rect 137520 10150 137590 10350
rect 137910 10150 137980 10350
rect 138020 10150 138090 10350
rect 138410 10150 138480 10350
rect 138520 10150 138590 10350
rect 138910 10150 138980 10350
rect 139020 10150 139090 10350
rect 139410 10150 139480 10350
rect 139520 10150 139590 10350
rect 139910 10150 139980 10350
rect 128150 10020 128350 10090
rect 128650 10020 128850 10090
rect 129150 10020 129350 10090
rect 129650 10020 129850 10090
rect 130150 10020 130350 10090
rect 130650 10020 130850 10090
rect 131150 10020 131350 10090
rect 131650 10020 131850 10090
rect 132150 10020 132350 10090
rect 132650 10020 132850 10090
rect 133150 10020 133350 10090
rect 133650 10020 133850 10090
rect 134150 10020 134350 10090
rect 134650 10020 134850 10090
rect 135150 10020 135350 10090
rect 135650 10020 135850 10090
rect 136150 10020 136350 10090
rect 136650 10020 136850 10090
rect 137150 10020 137350 10090
rect 137650 10020 137850 10090
rect 138150 10020 138350 10090
rect 138650 10020 138850 10090
rect 139150 10020 139350 10090
rect 139650 10020 139850 10090
rect 128150 9910 128350 9980
rect 128650 9910 128850 9980
rect 129150 9910 129350 9980
rect 129650 9910 129850 9980
rect 130150 9910 130350 9980
rect 130650 9910 130850 9980
rect 131150 9910 131350 9980
rect 131650 9910 131850 9980
rect 132150 9910 132350 9980
rect 132650 9910 132850 9980
rect 133150 9910 133350 9980
rect 133650 9910 133850 9980
rect 134150 9910 134350 9980
rect 134650 9910 134850 9980
rect 135150 9910 135350 9980
rect 135650 9910 135850 9980
rect 136150 9910 136350 9980
rect 136650 9910 136850 9980
rect 137150 9910 137350 9980
rect 137650 9910 137850 9980
rect 138150 9910 138350 9980
rect 138650 9910 138850 9980
rect 139150 9910 139350 9980
rect 139650 9910 139850 9980
rect 128020 9650 128090 9850
rect 128410 9650 128480 9850
rect 128520 9650 128590 9850
rect 128910 9650 128980 9850
rect 129020 9650 129090 9850
rect 129410 9650 129480 9850
rect 129520 9650 129590 9850
rect 129910 9650 129980 9850
rect 130020 9650 130090 9850
rect 130410 9650 130480 9850
rect 130520 9650 130590 9850
rect 130910 9650 130980 9850
rect 131020 9650 131090 9850
rect 131410 9650 131480 9850
rect 131520 9650 131590 9850
rect 131910 9650 131980 9850
rect 132020 9650 132090 9850
rect 132410 9650 132480 9850
rect 132520 9650 132590 9850
rect 132910 9650 132980 9850
rect 133020 9650 133090 9850
rect 133410 9650 133480 9850
rect 133520 9650 133590 9850
rect 133910 9650 133980 9850
rect 134020 9650 134090 9850
rect 134410 9650 134480 9850
rect 134520 9650 134590 9850
rect 134910 9650 134980 9850
rect 135020 9650 135090 9850
rect 135410 9650 135480 9850
rect 135520 9650 135590 9850
rect 135910 9650 135980 9850
rect 136020 9650 136090 9850
rect 136410 9650 136480 9850
rect 136520 9650 136590 9850
rect 136910 9650 136980 9850
rect 137020 9650 137090 9850
rect 137410 9650 137480 9850
rect 137520 9650 137590 9850
rect 137910 9650 137980 9850
rect 138020 9650 138090 9850
rect 138410 9650 138480 9850
rect 138520 9650 138590 9850
rect 138910 9650 138980 9850
rect 139020 9650 139090 9850
rect 139410 9650 139480 9850
rect 139520 9650 139590 9850
rect 139910 9650 139980 9850
rect 128150 9520 128350 9590
rect 128650 9520 128850 9590
rect 129150 9520 129350 9590
rect 129650 9520 129850 9590
rect 130150 9520 130350 9590
rect 130650 9520 130850 9590
rect 131150 9520 131350 9590
rect 131650 9520 131850 9590
rect 132150 9520 132350 9590
rect 132650 9520 132850 9590
rect 133150 9520 133350 9590
rect 133650 9520 133850 9590
rect 134150 9520 134350 9590
rect 134650 9520 134850 9590
rect 135150 9520 135350 9590
rect 135650 9520 135850 9590
rect 136150 9520 136350 9590
rect 136650 9520 136850 9590
rect 137150 9520 137350 9590
rect 137650 9520 137850 9590
rect 138150 9520 138350 9590
rect 138650 9520 138850 9590
rect 139150 9520 139350 9590
rect 139650 9520 139850 9590
rect 128150 9410 128350 9480
rect 128650 9410 128850 9480
rect 129150 9410 129350 9480
rect 129650 9410 129850 9480
rect 130150 9410 130350 9480
rect 130650 9410 130850 9480
rect 131150 9410 131350 9480
rect 131650 9410 131850 9480
rect 132150 9410 132350 9480
rect 132650 9410 132850 9480
rect 133150 9410 133350 9480
rect 133650 9410 133850 9480
rect 134150 9410 134350 9480
rect 134650 9410 134850 9480
rect 135150 9410 135350 9480
rect 135650 9410 135850 9480
rect 136150 9410 136350 9480
rect 136650 9410 136850 9480
rect 137150 9410 137350 9480
rect 137650 9410 137850 9480
rect 138150 9410 138350 9480
rect 138650 9410 138850 9480
rect 139150 9410 139350 9480
rect 139650 9410 139850 9480
rect 128020 9150 128090 9350
rect 128410 9150 128480 9350
rect 128520 9150 128590 9350
rect 128910 9150 128980 9350
rect 129020 9150 129090 9350
rect 129410 9150 129480 9350
rect 129520 9150 129590 9350
rect 129910 9150 129980 9350
rect 130020 9150 130090 9350
rect 130410 9150 130480 9350
rect 130520 9150 130590 9350
rect 130910 9150 130980 9350
rect 131020 9150 131090 9350
rect 131410 9150 131480 9350
rect 131520 9150 131590 9350
rect 131910 9150 131980 9350
rect 132020 9150 132090 9350
rect 132410 9150 132480 9350
rect 132520 9150 132590 9350
rect 132910 9150 132980 9350
rect 133020 9150 133090 9350
rect 133410 9150 133480 9350
rect 133520 9150 133590 9350
rect 133910 9150 133980 9350
rect 134020 9150 134090 9350
rect 134410 9150 134480 9350
rect 134520 9150 134590 9350
rect 134910 9150 134980 9350
rect 135020 9150 135090 9350
rect 135410 9150 135480 9350
rect 135520 9150 135590 9350
rect 135910 9150 135980 9350
rect 136020 9150 136090 9350
rect 136410 9150 136480 9350
rect 136520 9150 136590 9350
rect 136910 9150 136980 9350
rect 137020 9150 137090 9350
rect 137410 9150 137480 9350
rect 137520 9150 137590 9350
rect 137910 9150 137980 9350
rect 138020 9150 138090 9350
rect 138410 9150 138480 9350
rect 138520 9150 138590 9350
rect 138910 9150 138980 9350
rect 139020 9150 139090 9350
rect 139410 9150 139480 9350
rect 139520 9150 139590 9350
rect 139910 9150 139980 9350
rect 128150 9020 128350 9090
rect 128650 9020 128850 9090
rect 129150 9020 129350 9090
rect 129650 9020 129850 9090
rect 130150 9020 130350 9090
rect 130650 9020 130850 9090
rect 131150 9020 131350 9090
rect 131650 9020 131850 9090
rect 132150 9020 132350 9090
rect 132650 9020 132850 9090
rect 133150 9020 133350 9090
rect 133650 9020 133850 9090
rect 134150 9020 134350 9090
rect 134650 9020 134850 9090
rect 135150 9020 135350 9090
rect 135650 9020 135850 9090
rect 136150 9020 136350 9090
rect 136650 9020 136850 9090
rect 137150 9020 137350 9090
rect 137650 9020 137850 9090
rect 138150 9020 138350 9090
rect 138650 9020 138850 9090
rect 139150 9020 139350 9090
rect 139650 9020 139850 9090
rect 128150 8910 128350 8980
rect 128650 8910 128850 8980
rect 129150 8910 129350 8980
rect 129650 8910 129850 8980
rect 130150 8910 130350 8980
rect 130650 8910 130850 8980
rect 131150 8910 131350 8980
rect 131650 8910 131850 8980
rect 132150 8910 132350 8980
rect 132650 8910 132850 8980
rect 133150 8910 133350 8980
rect 133650 8910 133850 8980
rect 134150 8910 134350 8980
rect 134650 8910 134850 8980
rect 135150 8910 135350 8980
rect 135650 8910 135850 8980
rect 136150 8910 136350 8980
rect 136650 8910 136850 8980
rect 137150 8910 137350 8980
rect 137650 8910 137850 8980
rect 138150 8910 138350 8980
rect 138650 8910 138850 8980
rect 139150 8910 139350 8980
rect 139650 8910 139850 8980
rect 128020 8650 128090 8850
rect 128410 8650 128480 8850
rect 128520 8650 128590 8850
rect 128910 8650 128980 8850
rect 129020 8650 129090 8850
rect 129410 8650 129480 8850
rect 129520 8650 129590 8850
rect 129910 8650 129980 8850
rect 130020 8650 130090 8850
rect 130410 8650 130480 8850
rect 130520 8650 130590 8850
rect 130910 8650 130980 8850
rect 131020 8650 131090 8850
rect 131410 8650 131480 8850
rect 131520 8650 131590 8850
rect 131910 8650 131980 8850
rect 132020 8650 132090 8850
rect 132410 8650 132480 8850
rect 132520 8650 132590 8850
rect 132910 8650 132980 8850
rect 133020 8650 133090 8850
rect 133410 8650 133480 8850
rect 133520 8650 133590 8850
rect 133910 8650 133980 8850
rect 134020 8650 134090 8850
rect 134410 8650 134480 8850
rect 134520 8650 134590 8850
rect 134910 8650 134980 8850
rect 135020 8650 135090 8850
rect 135410 8650 135480 8850
rect 135520 8650 135590 8850
rect 135910 8650 135980 8850
rect 136020 8650 136090 8850
rect 136410 8650 136480 8850
rect 136520 8650 136590 8850
rect 136910 8650 136980 8850
rect 137020 8650 137090 8850
rect 137410 8650 137480 8850
rect 137520 8650 137590 8850
rect 137910 8650 137980 8850
rect 138020 8650 138090 8850
rect 138410 8650 138480 8850
rect 138520 8650 138590 8850
rect 138910 8650 138980 8850
rect 139020 8650 139090 8850
rect 139410 8650 139480 8850
rect 139520 8650 139590 8850
rect 139910 8650 139980 8850
rect 128150 8520 128350 8590
rect 128650 8520 128850 8590
rect 129150 8520 129350 8590
rect 129650 8520 129850 8590
rect 130150 8520 130350 8590
rect 130650 8520 130850 8590
rect 131150 8520 131350 8590
rect 131650 8520 131850 8590
rect 132150 8520 132350 8590
rect 132650 8520 132850 8590
rect 133150 8520 133350 8590
rect 133650 8520 133850 8590
rect 134150 8520 134350 8590
rect 134650 8520 134850 8590
rect 135150 8520 135350 8590
rect 135650 8520 135850 8590
rect 136150 8520 136350 8590
rect 136650 8520 136850 8590
rect 137150 8520 137350 8590
rect 137650 8520 137850 8590
rect 138150 8520 138350 8590
rect 138650 8520 138850 8590
rect 139150 8520 139350 8590
rect 139650 8520 139850 8590
rect 128150 8410 128350 8480
rect 128650 8410 128850 8480
rect 129150 8410 129350 8480
rect 129650 8410 129850 8480
rect 130150 8410 130350 8480
rect 130650 8410 130850 8480
rect 131150 8410 131350 8480
rect 131650 8410 131850 8480
rect 132150 8410 132350 8480
rect 132650 8410 132850 8480
rect 133150 8410 133350 8480
rect 133650 8410 133850 8480
rect 134150 8410 134350 8480
rect 134650 8410 134850 8480
rect 135150 8410 135350 8480
rect 135650 8410 135850 8480
rect 136150 8410 136350 8480
rect 136650 8410 136850 8480
rect 137150 8410 137350 8480
rect 137650 8410 137850 8480
rect 138150 8410 138350 8480
rect 138650 8410 138850 8480
rect 139150 8410 139350 8480
rect 139650 8410 139850 8480
rect 128020 8150 128090 8350
rect 128410 8150 128480 8350
rect 128520 8150 128590 8350
rect 128910 8150 128980 8350
rect 129020 8150 129090 8350
rect 129410 8150 129480 8350
rect 129520 8150 129590 8350
rect 129910 8150 129980 8350
rect 130020 8150 130090 8350
rect 130410 8150 130480 8350
rect 130520 8150 130590 8350
rect 130910 8150 130980 8350
rect 131020 8150 131090 8350
rect 131410 8150 131480 8350
rect 131520 8150 131590 8350
rect 131910 8150 131980 8350
rect 132020 8150 132090 8350
rect 132410 8150 132480 8350
rect 132520 8150 132590 8350
rect 132910 8150 132980 8350
rect 133020 8150 133090 8350
rect 133410 8150 133480 8350
rect 133520 8150 133590 8350
rect 133910 8150 133980 8350
rect 134020 8150 134090 8350
rect 134410 8150 134480 8350
rect 134520 8150 134590 8350
rect 134910 8150 134980 8350
rect 135020 8150 135090 8350
rect 135410 8150 135480 8350
rect 135520 8150 135590 8350
rect 135910 8150 135980 8350
rect 136020 8150 136090 8350
rect 136410 8150 136480 8350
rect 136520 8150 136590 8350
rect 136910 8150 136980 8350
rect 137020 8150 137090 8350
rect 137410 8150 137480 8350
rect 137520 8150 137590 8350
rect 137910 8150 137980 8350
rect 138020 8150 138090 8350
rect 138410 8150 138480 8350
rect 138520 8150 138590 8350
rect 138910 8150 138980 8350
rect 139020 8150 139090 8350
rect 139410 8150 139480 8350
rect 139520 8150 139590 8350
rect 139910 8150 139980 8350
rect 128150 8020 128350 8090
rect 128650 8020 128850 8090
rect 129150 8020 129350 8090
rect 129650 8020 129850 8090
rect 130150 8020 130350 8090
rect 130650 8020 130850 8090
rect 131150 8020 131350 8090
rect 131650 8020 131850 8090
rect 132150 8020 132350 8090
rect 132650 8020 132850 8090
rect 133150 8020 133350 8090
rect 133650 8020 133850 8090
rect 134150 8020 134350 8090
rect 134650 8020 134850 8090
rect 135150 8020 135350 8090
rect 135650 8020 135850 8090
rect 136150 8020 136350 8090
rect 136650 8020 136850 8090
rect 137150 8020 137350 8090
rect 137650 8020 137850 8090
rect 138150 8020 138350 8090
rect 138650 8020 138850 8090
rect 139150 8020 139350 8090
rect 139650 8020 139850 8090
rect 128150 7910 128350 7980
rect 128650 7910 128850 7980
rect 129150 7910 129350 7980
rect 129650 7910 129850 7980
rect 130150 7910 130350 7980
rect 130650 7910 130850 7980
rect 131150 7910 131350 7980
rect 131650 7910 131850 7980
rect 132150 7910 132350 7980
rect 132650 7910 132850 7980
rect 133150 7910 133350 7980
rect 133650 7910 133850 7980
rect 134150 7910 134350 7980
rect 134650 7910 134850 7980
rect 135150 7910 135350 7980
rect 135650 7910 135850 7980
rect 136150 7910 136350 7980
rect 136650 7910 136850 7980
rect 137150 7910 137350 7980
rect 137650 7910 137850 7980
rect 138150 7910 138350 7980
rect 138650 7910 138850 7980
rect 139150 7910 139350 7980
rect 139650 7910 139850 7980
rect 128020 7650 128090 7850
rect 128410 7650 128480 7850
rect 128520 7650 128590 7850
rect 128910 7650 128980 7850
rect 129020 7650 129090 7850
rect 129410 7650 129480 7850
rect 129520 7650 129590 7850
rect 129910 7650 129980 7850
rect 130020 7650 130090 7850
rect 130410 7650 130480 7850
rect 130520 7650 130590 7850
rect 130910 7650 130980 7850
rect 131020 7650 131090 7850
rect 131410 7650 131480 7850
rect 131520 7650 131590 7850
rect 131910 7650 131980 7850
rect 132020 7650 132090 7850
rect 132410 7650 132480 7850
rect 132520 7650 132590 7850
rect 132910 7650 132980 7850
rect 133020 7650 133090 7850
rect 133410 7650 133480 7850
rect 133520 7650 133590 7850
rect 133910 7650 133980 7850
rect 134020 7650 134090 7850
rect 134410 7650 134480 7850
rect 134520 7650 134590 7850
rect 134910 7650 134980 7850
rect 135020 7650 135090 7850
rect 135410 7650 135480 7850
rect 135520 7650 135590 7850
rect 135910 7650 135980 7850
rect 136020 7650 136090 7850
rect 136410 7650 136480 7850
rect 136520 7650 136590 7850
rect 136910 7650 136980 7850
rect 137020 7650 137090 7850
rect 137410 7650 137480 7850
rect 137520 7650 137590 7850
rect 137910 7650 137980 7850
rect 138020 7650 138090 7850
rect 138410 7650 138480 7850
rect 138520 7650 138590 7850
rect 138910 7650 138980 7850
rect 139020 7650 139090 7850
rect 139410 7650 139480 7850
rect 139520 7650 139590 7850
rect 139910 7650 139980 7850
rect 128150 7520 128350 7590
rect 128650 7520 128850 7590
rect 129150 7520 129350 7590
rect 129650 7520 129850 7590
rect 130150 7520 130350 7590
rect 130650 7520 130850 7590
rect 131150 7520 131350 7590
rect 131650 7520 131850 7590
rect 132150 7520 132350 7590
rect 132650 7520 132850 7590
rect 133150 7520 133350 7590
rect 133650 7520 133850 7590
rect 134150 7520 134350 7590
rect 134650 7520 134850 7590
rect 135150 7520 135350 7590
rect 135650 7520 135850 7590
rect 136150 7520 136350 7590
rect 136650 7520 136850 7590
rect 137150 7520 137350 7590
rect 137650 7520 137850 7590
rect 138150 7520 138350 7590
rect 138650 7520 138850 7590
rect 139150 7520 139350 7590
rect 139650 7520 139850 7590
rect 128150 7410 128350 7480
rect 128650 7410 128850 7480
rect 129150 7410 129350 7480
rect 129650 7410 129850 7480
rect 130150 7410 130350 7480
rect 130650 7410 130850 7480
rect 131150 7410 131350 7480
rect 131650 7410 131850 7480
rect 132150 7410 132350 7480
rect 132650 7410 132850 7480
rect 133150 7410 133350 7480
rect 133650 7410 133850 7480
rect 134150 7410 134350 7480
rect 134650 7410 134850 7480
rect 135150 7410 135350 7480
rect 135650 7410 135850 7480
rect 136150 7410 136350 7480
rect 136650 7410 136850 7480
rect 137150 7410 137350 7480
rect 137650 7410 137850 7480
rect 138150 7410 138350 7480
rect 138650 7410 138850 7480
rect 139150 7410 139350 7480
rect 139650 7410 139850 7480
rect 128020 7150 128090 7350
rect 128410 7150 128480 7350
rect 128520 7150 128590 7350
rect 128910 7150 128980 7350
rect 129020 7150 129090 7350
rect 129410 7150 129480 7350
rect 129520 7150 129590 7350
rect 129910 7150 129980 7350
rect 130020 7150 130090 7350
rect 130410 7150 130480 7350
rect 130520 7150 130590 7350
rect 130910 7150 130980 7350
rect 131020 7150 131090 7350
rect 131410 7150 131480 7350
rect 131520 7150 131590 7350
rect 131910 7150 131980 7350
rect 132020 7150 132090 7350
rect 132410 7150 132480 7350
rect 132520 7150 132590 7350
rect 132910 7150 132980 7350
rect 133020 7150 133090 7350
rect 133410 7150 133480 7350
rect 133520 7150 133590 7350
rect 133910 7150 133980 7350
rect 134020 7150 134090 7350
rect 134410 7150 134480 7350
rect 134520 7150 134590 7350
rect 134910 7150 134980 7350
rect 135020 7150 135090 7350
rect 135410 7150 135480 7350
rect 135520 7150 135590 7350
rect 135910 7150 135980 7350
rect 136020 7150 136090 7350
rect 136410 7150 136480 7350
rect 136520 7150 136590 7350
rect 136910 7150 136980 7350
rect 137020 7150 137090 7350
rect 137410 7150 137480 7350
rect 137520 7150 137590 7350
rect 137910 7150 137980 7350
rect 138020 7150 138090 7350
rect 138410 7150 138480 7350
rect 138520 7150 138590 7350
rect 138910 7150 138980 7350
rect 139020 7150 139090 7350
rect 139410 7150 139480 7350
rect 139520 7150 139590 7350
rect 139910 7150 139980 7350
rect 128150 7020 128350 7090
rect 128650 7020 128850 7090
rect 129150 7020 129350 7090
rect 129650 7020 129850 7090
rect 130150 7020 130350 7090
rect 130650 7020 130850 7090
rect 131150 7020 131350 7090
rect 131650 7020 131850 7090
rect 132150 7020 132350 7090
rect 132650 7020 132850 7090
rect 133150 7020 133350 7090
rect 133650 7020 133850 7090
rect 134150 7020 134350 7090
rect 134650 7020 134850 7090
rect 135150 7020 135350 7090
rect 135650 7020 135850 7090
rect 136150 7020 136350 7090
rect 136650 7020 136850 7090
rect 137150 7020 137350 7090
rect 137650 7020 137850 7090
rect 138150 7020 138350 7090
rect 138650 7020 138850 7090
rect 139150 7020 139350 7090
rect 139650 7020 139850 7090
rect 128150 6910 128350 6980
rect 128650 6910 128850 6980
rect 129150 6910 129350 6980
rect 129650 6910 129850 6980
rect 130150 6910 130350 6980
rect 130650 6910 130850 6980
rect 131150 6910 131350 6980
rect 131650 6910 131850 6980
rect 132150 6910 132350 6980
rect 132650 6910 132850 6980
rect 133150 6910 133350 6980
rect 133650 6910 133850 6980
rect 134150 6910 134350 6980
rect 134650 6910 134850 6980
rect 135150 6910 135350 6980
rect 135650 6910 135850 6980
rect 136150 6910 136350 6980
rect 136650 6910 136850 6980
rect 137150 6910 137350 6980
rect 137650 6910 137850 6980
rect 138150 6910 138350 6980
rect 138650 6910 138850 6980
rect 139150 6910 139350 6980
rect 139650 6910 139850 6980
rect 128020 6650 128090 6850
rect 128410 6650 128480 6850
rect 128520 6650 128590 6850
rect 128910 6650 128980 6850
rect 129020 6650 129090 6850
rect 129410 6650 129480 6850
rect 129520 6650 129590 6850
rect 129910 6650 129980 6850
rect 130020 6650 130090 6850
rect 130410 6650 130480 6850
rect 130520 6650 130590 6850
rect 130910 6650 130980 6850
rect 131020 6650 131090 6850
rect 131410 6650 131480 6850
rect 131520 6650 131590 6850
rect 131910 6650 131980 6850
rect 132020 6650 132090 6850
rect 132410 6650 132480 6850
rect 132520 6650 132590 6850
rect 132910 6650 132980 6850
rect 133020 6650 133090 6850
rect 133410 6650 133480 6850
rect 133520 6650 133590 6850
rect 133910 6650 133980 6850
rect 134020 6650 134090 6850
rect 134410 6650 134480 6850
rect 134520 6650 134590 6850
rect 134910 6650 134980 6850
rect 135020 6650 135090 6850
rect 135410 6650 135480 6850
rect 135520 6650 135590 6850
rect 135910 6650 135980 6850
rect 136020 6650 136090 6850
rect 136410 6650 136480 6850
rect 136520 6650 136590 6850
rect 136910 6650 136980 6850
rect 137020 6650 137090 6850
rect 137410 6650 137480 6850
rect 137520 6650 137590 6850
rect 137910 6650 137980 6850
rect 138020 6650 138090 6850
rect 138410 6650 138480 6850
rect 138520 6650 138590 6850
rect 138910 6650 138980 6850
rect 139020 6650 139090 6850
rect 139410 6650 139480 6850
rect 139520 6650 139590 6850
rect 139910 6650 139980 6850
rect 128150 6520 128350 6590
rect 128650 6520 128850 6590
rect 129150 6520 129350 6590
rect 129650 6520 129850 6590
rect 130150 6520 130350 6590
rect 130650 6520 130850 6590
rect 131150 6520 131350 6590
rect 131650 6520 131850 6590
rect 132150 6520 132350 6590
rect 132650 6520 132850 6590
rect 133150 6520 133350 6590
rect 133650 6520 133850 6590
rect 134150 6520 134350 6590
rect 134650 6520 134850 6590
rect 135150 6520 135350 6590
rect 135650 6520 135850 6590
rect 136150 6520 136350 6590
rect 136650 6520 136850 6590
rect 137150 6520 137350 6590
rect 137650 6520 137850 6590
rect 138150 6520 138350 6590
rect 138650 6520 138850 6590
rect 139150 6520 139350 6590
rect 139650 6520 139850 6590
rect 128150 6410 128350 6480
rect 128650 6410 128850 6480
rect 129150 6410 129350 6480
rect 129650 6410 129850 6480
rect 130150 6410 130350 6480
rect 130650 6410 130850 6480
rect 131150 6410 131350 6480
rect 131650 6410 131850 6480
rect 132150 6410 132350 6480
rect 132650 6410 132850 6480
rect 133150 6410 133350 6480
rect 133650 6410 133850 6480
rect 134150 6410 134350 6480
rect 134650 6410 134850 6480
rect 135150 6410 135350 6480
rect 135650 6410 135850 6480
rect 136150 6410 136350 6480
rect 136650 6410 136850 6480
rect 137150 6410 137350 6480
rect 137650 6410 137850 6480
rect 138150 6410 138350 6480
rect 138650 6410 138850 6480
rect 139150 6410 139350 6480
rect 139650 6410 139850 6480
rect 128020 6150 128090 6350
rect 128410 6150 128480 6350
rect 128520 6150 128590 6350
rect 128910 6150 128980 6350
rect 129020 6150 129090 6350
rect 129410 6150 129480 6350
rect 129520 6150 129590 6350
rect 129910 6150 129980 6350
rect 130020 6150 130090 6350
rect 130410 6150 130480 6350
rect 130520 6150 130590 6350
rect 130910 6150 130980 6350
rect 131020 6150 131090 6350
rect 131410 6150 131480 6350
rect 131520 6150 131590 6350
rect 131910 6150 131980 6350
rect 132020 6150 132090 6350
rect 132410 6150 132480 6350
rect 132520 6150 132590 6350
rect 132910 6150 132980 6350
rect 133020 6150 133090 6350
rect 133410 6150 133480 6350
rect 133520 6150 133590 6350
rect 133910 6150 133980 6350
rect 134020 6150 134090 6350
rect 134410 6150 134480 6350
rect 134520 6150 134590 6350
rect 134910 6150 134980 6350
rect 135020 6150 135090 6350
rect 135410 6150 135480 6350
rect 135520 6150 135590 6350
rect 135910 6150 135980 6350
rect 136020 6150 136090 6350
rect 136410 6150 136480 6350
rect 136520 6150 136590 6350
rect 136910 6150 136980 6350
rect 137020 6150 137090 6350
rect 137410 6150 137480 6350
rect 137520 6150 137590 6350
rect 137910 6150 137980 6350
rect 138020 6150 138090 6350
rect 138410 6150 138480 6350
rect 138520 6150 138590 6350
rect 138910 6150 138980 6350
rect 139020 6150 139090 6350
rect 139410 6150 139480 6350
rect 139520 6150 139590 6350
rect 139910 6150 139980 6350
rect 128150 6020 128350 6090
rect 128650 6020 128850 6090
rect 129150 6020 129350 6090
rect 129650 6020 129850 6090
rect 130150 6020 130350 6090
rect 130650 6020 130850 6090
rect 131150 6020 131350 6090
rect 131650 6020 131850 6090
rect 132150 6020 132350 6090
rect 132650 6020 132850 6090
rect 133150 6020 133350 6090
rect 133650 6020 133850 6090
rect 134150 6020 134350 6090
rect 134650 6020 134850 6090
rect 135150 6020 135350 6090
rect 135650 6020 135850 6090
rect 136150 6020 136350 6090
rect 136650 6020 136850 6090
rect 137150 6020 137350 6090
rect 137650 6020 137850 6090
rect 138150 6020 138350 6090
rect 138650 6020 138850 6090
rect 139150 6020 139350 6090
rect 139650 6020 139850 6090
rect 136150 5910 136350 5980
rect 136650 5910 136850 5980
rect 137150 5910 137350 5980
rect 137650 5910 137850 5980
rect 138150 5910 138350 5980
rect 138650 5910 138850 5980
rect 139150 5910 139350 5980
rect 139650 5910 139850 5980
rect 136020 5650 136090 5850
rect 136410 5650 136480 5850
rect 136520 5650 136590 5850
rect 136910 5650 136980 5850
rect 137020 5650 137090 5850
rect 137410 5650 137480 5850
rect 137520 5650 137590 5850
rect 137910 5650 137980 5850
rect 138020 5650 138090 5850
rect 138410 5650 138480 5850
rect 138520 5650 138590 5850
rect 138910 5650 138980 5850
rect 139020 5650 139090 5850
rect 139410 5650 139480 5850
rect 139520 5650 139590 5850
rect 139910 5650 139980 5850
rect 136150 5520 136350 5590
rect 136650 5520 136850 5590
rect 137150 5520 137350 5590
rect 137650 5520 137850 5590
rect 138150 5520 138350 5590
rect 138650 5520 138850 5590
rect 139150 5520 139350 5590
rect 139650 5520 139850 5590
rect 136150 5410 136350 5480
rect 136650 5410 136850 5480
rect 137150 5410 137350 5480
rect 137650 5410 137850 5480
rect 138150 5410 138350 5480
rect 138650 5410 138850 5480
rect 139150 5410 139350 5480
rect 139650 5410 139850 5480
rect 136020 5150 136090 5350
rect 136410 5150 136480 5350
rect 136520 5150 136590 5350
rect 136910 5150 136980 5350
rect 137020 5150 137090 5350
rect 137410 5150 137480 5350
rect 137520 5150 137590 5350
rect 137910 5150 137980 5350
rect 138020 5150 138090 5350
rect 138410 5150 138480 5350
rect 138520 5150 138590 5350
rect 138910 5150 138980 5350
rect 139020 5150 139090 5350
rect 139410 5150 139480 5350
rect 139520 5150 139590 5350
rect 139910 5150 139980 5350
rect 136150 5020 136350 5090
rect 136650 5020 136850 5090
rect 137150 5020 137350 5090
rect 137650 5020 137850 5090
rect 138150 5020 138350 5090
rect 138650 5020 138850 5090
rect 139150 5020 139350 5090
rect 139650 5020 139850 5090
rect 136150 4910 136350 4980
rect 136650 4910 136850 4980
rect 137150 4910 137350 4980
rect 137650 4910 137850 4980
rect 138150 4910 138350 4980
rect 138650 4910 138850 4980
rect 139150 4910 139350 4980
rect 139650 4910 139850 4980
rect 136020 4650 136090 4850
rect 136410 4650 136480 4850
rect 136520 4650 136590 4850
rect 136910 4650 136980 4850
rect 137020 4650 137090 4850
rect 137410 4650 137480 4850
rect 137520 4650 137590 4850
rect 137910 4650 137980 4850
rect 138020 4650 138090 4850
rect 138410 4650 138480 4850
rect 138520 4650 138590 4850
rect 138910 4650 138980 4850
rect 139020 4650 139090 4850
rect 139410 4650 139480 4850
rect 139520 4650 139590 4850
rect 139910 4650 139980 4850
rect 136150 4520 136350 4590
rect 136650 4520 136850 4590
rect 137150 4520 137350 4590
rect 137650 4520 137850 4590
rect 138150 4520 138350 4590
rect 138650 4520 138850 4590
rect 139150 4520 139350 4590
rect 139650 4520 139850 4590
rect 136150 4410 136350 4480
rect 136650 4410 136850 4480
rect 137150 4410 137350 4480
rect 137650 4410 137850 4480
rect 138150 4410 138350 4480
rect 138650 4410 138850 4480
rect 139150 4410 139350 4480
rect 139650 4410 139850 4480
rect 136020 4150 136090 4350
rect 136410 4150 136480 4350
rect 136520 4150 136590 4350
rect 136910 4150 136980 4350
rect 137020 4150 137090 4350
rect 137410 4150 137480 4350
rect 137520 4150 137590 4350
rect 137910 4150 137980 4350
rect 138020 4150 138090 4350
rect 138410 4150 138480 4350
rect 138520 4150 138590 4350
rect 138910 4150 138980 4350
rect 139020 4150 139090 4350
rect 139410 4150 139480 4350
rect 139520 4150 139590 4350
rect 139910 4150 139980 4350
rect 136150 4020 136350 4090
rect 136650 4020 136850 4090
rect 137150 4020 137350 4090
rect 137650 4020 137850 4090
rect 138150 4020 138350 4090
rect 138650 4020 138850 4090
rect 139150 4020 139350 4090
rect 139650 4020 139850 4090
rect 136150 3910 136350 3980
rect 136650 3910 136850 3980
rect 137150 3910 137350 3980
rect 137650 3910 137850 3980
rect 138150 3910 138350 3980
rect 138650 3910 138850 3980
rect 139150 3910 139350 3980
rect 139650 3910 139850 3980
rect 136020 3650 136090 3850
rect 136410 3650 136480 3850
rect 136520 3650 136590 3850
rect 136910 3650 136980 3850
rect 137020 3650 137090 3850
rect 137410 3650 137480 3850
rect 137520 3650 137590 3850
rect 137910 3650 137980 3850
rect 138020 3650 138090 3850
rect 138410 3650 138480 3850
rect 138520 3650 138590 3850
rect 138910 3650 138980 3850
rect 139020 3650 139090 3850
rect 139410 3650 139480 3850
rect 139520 3650 139590 3850
rect 139910 3650 139980 3850
rect 136150 3520 136350 3590
rect 136650 3520 136850 3590
rect 137150 3520 137350 3590
rect 137650 3520 137850 3590
rect 138150 3520 138350 3590
rect 138650 3520 138850 3590
rect 139150 3520 139350 3590
rect 139650 3520 139850 3590
rect 136150 3410 136350 3480
rect 136650 3410 136850 3480
rect 137150 3410 137350 3480
rect 137650 3410 137850 3480
rect 138150 3410 138350 3480
rect 138650 3410 138850 3480
rect 139150 3410 139350 3480
rect 139650 3410 139850 3480
rect 136020 3150 136090 3350
rect 136410 3150 136480 3350
rect 136520 3150 136590 3350
rect 136910 3150 136980 3350
rect 137020 3150 137090 3350
rect 137410 3150 137480 3350
rect 137520 3150 137590 3350
rect 137910 3150 137980 3350
rect 138020 3150 138090 3350
rect 138410 3150 138480 3350
rect 138520 3150 138590 3350
rect 138910 3150 138980 3350
rect 139020 3150 139090 3350
rect 139410 3150 139480 3350
rect 139520 3150 139590 3350
rect 139910 3150 139980 3350
rect 136150 3020 136350 3090
rect 136650 3020 136850 3090
rect 137150 3020 137350 3090
rect 137650 3020 137850 3090
rect 138150 3020 138350 3090
rect 138650 3020 138850 3090
rect 139150 3020 139350 3090
rect 139650 3020 139850 3090
rect 136150 2910 136350 2980
rect 136650 2910 136850 2980
rect 137150 2910 137350 2980
rect 137650 2910 137850 2980
rect 138150 2910 138350 2980
rect 138650 2910 138850 2980
rect 139150 2910 139350 2980
rect 139650 2910 139850 2980
rect 136020 2650 136090 2850
rect 136410 2650 136480 2850
rect 136520 2650 136590 2850
rect 136910 2650 136980 2850
rect 137020 2650 137090 2850
rect 137410 2650 137480 2850
rect 137520 2650 137590 2850
rect 137910 2650 137980 2850
rect 138020 2650 138090 2850
rect 138410 2650 138480 2850
rect 138520 2650 138590 2850
rect 138910 2650 138980 2850
rect 139020 2650 139090 2850
rect 139410 2650 139480 2850
rect 139520 2650 139590 2850
rect 139910 2650 139980 2850
rect 136150 2520 136350 2590
rect 136650 2520 136850 2590
rect 137150 2520 137350 2590
rect 137650 2520 137850 2590
rect 138150 2520 138350 2590
rect 138650 2520 138850 2590
rect 139150 2520 139350 2590
rect 139650 2520 139850 2590
rect 136150 2410 136350 2480
rect 136650 2410 136850 2480
rect 137150 2410 137350 2480
rect 137650 2410 137850 2480
rect 138150 2410 138350 2480
rect 138650 2410 138850 2480
rect 139150 2410 139350 2480
rect 139650 2410 139850 2480
rect 136020 2150 136090 2350
rect 136410 2150 136480 2350
rect 136520 2150 136590 2350
rect 136910 2150 136980 2350
rect 137020 2150 137090 2350
rect 137410 2150 137480 2350
rect 137520 2150 137590 2350
rect 137910 2150 137980 2350
rect 138020 2150 138090 2350
rect 138410 2150 138480 2350
rect 138520 2150 138590 2350
rect 138910 2150 138980 2350
rect 139020 2150 139090 2350
rect 139410 2150 139480 2350
rect 139520 2150 139590 2350
rect 139910 2150 139980 2350
rect 136150 2020 136350 2090
rect 136650 2020 136850 2090
rect 137150 2020 137350 2090
rect 137650 2020 137850 2090
rect 138150 2020 138350 2090
rect 138650 2020 138850 2090
rect 139150 2020 139350 2090
rect 139650 2020 139850 2090
rect 136150 1910 136350 1980
rect 136650 1910 136850 1980
rect 137150 1910 137350 1980
rect 137650 1910 137850 1980
rect 138150 1910 138350 1980
rect 138650 1910 138850 1980
rect 139150 1910 139350 1980
rect 139650 1910 139850 1980
rect 136020 1650 136090 1850
rect 136410 1650 136480 1850
rect 136520 1650 136590 1850
rect 136910 1650 136980 1850
rect 137020 1650 137090 1850
rect 137410 1650 137480 1850
rect 137520 1650 137590 1850
rect 137910 1650 137980 1850
rect 138020 1650 138090 1850
rect 138410 1650 138480 1850
rect 138520 1650 138590 1850
rect 138910 1650 138980 1850
rect 139020 1650 139090 1850
rect 139410 1650 139480 1850
rect 139520 1650 139590 1850
rect 139910 1650 139980 1850
rect 136150 1520 136350 1590
rect 136650 1520 136850 1590
rect 137150 1520 137350 1590
rect 137650 1520 137850 1590
rect 138150 1520 138350 1590
rect 138650 1520 138850 1590
rect 139150 1520 139350 1590
rect 139650 1520 139850 1590
rect 136150 1410 136350 1480
rect 136650 1410 136850 1480
rect 137150 1410 137350 1480
rect 137650 1410 137850 1480
rect 138150 1410 138350 1480
rect 138650 1410 138850 1480
rect 139150 1410 139350 1480
rect 139650 1410 139850 1480
rect 136020 1150 136090 1350
rect 136410 1150 136480 1350
rect 136520 1150 136590 1350
rect 136910 1150 136980 1350
rect 137020 1150 137090 1350
rect 137410 1150 137480 1350
rect 137520 1150 137590 1350
rect 137910 1150 137980 1350
rect 138020 1150 138090 1350
rect 138410 1150 138480 1350
rect 138520 1150 138590 1350
rect 138910 1150 138980 1350
rect 139020 1150 139090 1350
rect 139410 1150 139480 1350
rect 139520 1150 139590 1350
rect 139910 1150 139980 1350
rect 136150 1020 136350 1090
rect 136650 1020 136850 1090
rect 137150 1020 137350 1090
rect 137650 1020 137850 1090
rect 138150 1020 138350 1090
rect 138650 1020 138850 1090
rect 139150 1020 139350 1090
rect 139650 1020 139850 1090
rect 136150 910 136350 980
rect 136650 910 136850 980
rect 137150 910 137350 980
rect 137650 910 137850 980
rect 138150 910 138350 980
rect 138650 910 138850 980
rect 139150 910 139350 980
rect 139650 910 139850 980
rect 136020 650 136090 850
rect 136410 650 136480 850
rect 136520 650 136590 850
rect 136910 650 136980 850
rect 137020 650 137090 850
rect 137410 650 137480 850
rect 137520 650 137590 850
rect 137910 650 137980 850
rect 138020 650 138090 850
rect 138410 650 138480 850
rect 138520 650 138590 850
rect 138910 650 138980 850
rect 139020 650 139090 850
rect 139410 650 139480 850
rect 139520 650 139590 850
rect 139910 650 139980 850
rect 136150 520 136350 590
rect 136650 520 136850 590
rect 137150 520 137350 590
rect 137650 520 137850 590
rect 138150 520 138350 590
rect 138650 520 138850 590
rect 139150 520 139350 590
rect 139650 520 139850 590
rect 136150 410 136350 480
rect 136650 410 136850 480
rect 137150 410 137350 480
rect 137650 410 137850 480
rect 138150 410 138350 480
rect 138650 410 138850 480
rect 139150 410 139350 480
rect 139650 410 139850 480
rect 136020 150 136090 350
rect 136410 150 136480 350
rect 136520 150 136590 350
rect 136910 150 136980 350
rect 137020 150 137090 350
rect 137410 150 137480 350
rect 137520 150 137590 350
rect 137910 150 137980 350
rect 138020 150 138090 350
rect 138410 150 138480 350
rect 138520 150 138590 350
rect 138910 150 138980 350
rect 139020 150 139090 350
rect 139410 150 139480 350
rect 139520 150 139590 350
rect 139910 150 139980 350
rect 136150 20 136350 90
rect 136650 20 136850 90
rect 137150 20 137350 90
rect 137650 20 137850 90
rect 138150 20 138350 90
rect 138650 20 138850 90
rect 139150 20 139350 90
rect 139650 20 139850 90
rect 136150 -90 136350 -20
rect 136650 -90 136850 -20
rect 137150 -90 137350 -20
rect 137650 -90 137850 -20
rect 138150 -90 138350 -20
rect 138650 -90 138850 -20
rect 139150 -90 139350 -20
rect 139650 -90 139850 -20
rect 136020 -350 136090 -150
rect 136410 -350 136480 -150
rect 136520 -350 136590 -150
rect 136910 -350 136980 -150
rect 137020 -350 137090 -150
rect 137410 -350 137480 -150
rect 137520 -350 137590 -150
rect 137910 -350 137980 -150
rect 138020 -350 138090 -150
rect 138410 -350 138480 -150
rect 138520 -350 138590 -150
rect 138910 -350 138980 -150
rect 139020 -350 139090 -150
rect 139410 -350 139480 -150
rect 139520 -350 139590 -150
rect 139910 -350 139980 -150
rect 136150 -480 136350 -410
rect 136650 -480 136850 -410
rect 137150 -480 137350 -410
rect 137650 -480 137850 -410
rect 138150 -480 138350 -410
rect 138650 -480 138850 -410
rect 139150 -480 139350 -410
rect 139650 -480 139850 -410
rect 136150 -590 136350 -520
rect 136650 -590 136850 -520
rect 137150 -590 137350 -520
rect 137650 -590 137850 -520
rect 138150 -590 138350 -520
rect 138650 -590 138850 -520
rect 139150 -590 139350 -520
rect 139650 -590 139850 -520
rect 136020 -850 136090 -650
rect 136410 -850 136480 -650
rect 136520 -850 136590 -650
rect 136910 -850 136980 -650
rect 137020 -850 137090 -650
rect 137410 -850 137480 -650
rect 137520 -850 137590 -650
rect 137910 -850 137980 -650
rect 138020 -850 138090 -650
rect 138410 -850 138480 -650
rect 138520 -850 138590 -650
rect 138910 -850 138980 -650
rect 139020 -850 139090 -650
rect 139410 -850 139480 -650
rect 139520 -850 139590 -650
rect 139910 -850 139980 -650
rect 136150 -980 136350 -910
rect 136650 -980 136850 -910
rect 137150 -980 137350 -910
rect 137650 -980 137850 -910
rect 138150 -980 138350 -910
rect 138650 -980 138850 -910
rect 139150 -980 139350 -910
rect 139650 -980 139850 -910
rect 136150 -1090 136350 -1020
rect 136650 -1090 136850 -1020
rect 137150 -1090 137350 -1020
rect 137650 -1090 137850 -1020
rect 138150 -1090 138350 -1020
rect 138650 -1090 138850 -1020
rect 139150 -1090 139350 -1020
rect 139650 -1090 139850 -1020
rect 136020 -1350 136090 -1150
rect 136410 -1350 136480 -1150
rect 136520 -1350 136590 -1150
rect 136910 -1350 136980 -1150
rect 137020 -1350 137090 -1150
rect 137410 -1350 137480 -1150
rect 137520 -1350 137590 -1150
rect 137910 -1350 137980 -1150
rect 138020 -1350 138090 -1150
rect 138410 -1350 138480 -1150
rect 138520 -1350 138590 -1150
rect 138910 -1350 138980 -1150
rect 139020 -1350 139090 -1150
rect 139410 -1350 139480 -1150
rect 139520 -1350 139590 -1150
rect 139910 -1350 139980 -1150
rect 136150 -1480 136350 -1410
rect 136650 -1480 136850 -1410
rect 137150 -1480 137350 -1410
rect 137650 -1480 137850 -1410
rect 138150 -1480 138350 -1410
rect 138650 -1480 138850 -1410
rect 139150 -1480 139350 -1410
rect 139650 -1480 139850 -1410
rect 136150 -1590 136350 -1520
rect 136650 -1590 136850 -1520
rect 137150 -1590 137350 -1520
rect 137650 -1590 137850 -1520
rect 138150 -1590 138350 -1520
rect 138650 -1590 138850 -1520
rect 139150 -1590 139350 -1520
rect 139650 -1590 139850 -1520
rect 136020 -1850 136090 -1650
rect 136410 -1850 136480 -1650
rect 136520 -1850 136590 -1650
rect 136910 -1850 136980 -1650
rect 137020 -1850 137090 -1650
rect 137410 -1850 137480 -1650
rect 137520 -1850 137590 -1650
rect 137910 -1850 137980 -1650
rect 138020 -1850 138090 -1650
rect 138410 -1850 138480 -1650
rect 138520 -1850 138590 -1650
rect 138910 -1850 138980 -1650
rect 139020 -1850 139090 -1650
rect 139410 -1850 139480 -1650
rect 139520 -1850 139590 -1650
rect 139910 -1850 139980 -1650
rect 136150 -1980 136350 -1910
rect 136650 -1980 136850 -1910
rect 137150 -1980 137350 -1910
rect 137650 -1980 137850 -1910
rect 138150 -1980 138350 -1910
rect 138650 -1980 138850 -1910
rect 139150 -1980 139350 -1910
rect 139650 -1980 139850 -1910
<< metal2 >>
rect -15860 97980 -15640 98000
rect -15860 97910 -15850 97980
rect -15650 97910 -15640 97980
rect -15860 97860 -15640 97910
rect -15360 97980 -15140 98000
rect -15360 97910 -15350 97980
rect -15150 97910 -15140 97980
rect -15360 97860 -15140 97910
rect -14860 97980 -14640 98000
rect -14860 97910 -14850 97980
rect -14650 97910 -14640 97980
rect -14860 97860 -14640 97910
rect -14360 97980 -14140 98000
rect -14360 97910 -14350 97980
rect -14150 97910 -14140 97980
rect -14360 97860 -14140 97910
rect -13860 97980 -13640 98000
rect -13860 97910 -13850 97980
rect -13650 97910 -13640 97980
rect -13860 97860 -13640 97910
rect -13360 97980 -13140 98000
rect -13360 97910 -13350 97980
rect -13150 97910 -13140 97980
rect -13360 97860 -13140 97910
rect -12860 97980 -12640 98000
rect -12860 97910 -12850 97980
rect -12650 97910 -12640 97980
rect -12860 97860 -12640 97910
rect -12360 97980 -12140 98000
rect -12360 97910 -12350 97980
rect -12150 97910 -12140 97980
rect -12360 97860 -12140 97910
rect -11860 97980 -11640 98000
rect -11860 97910 -11850 97980
rect -11650 97910 -11640 97980
rect -11860 97860 -11640 97910
rect -11360 97980 -11140 98000
rect -11360 97910 -11350 97980
rect -11150 97910 -11140 97980
rect -11360 97860 -11140 97910
rect -10860 97980 -10640 98000
rect -10860 97910 -10850 97980
rect -10650 97910 -10640 97980
rect -10860 97860 -10640 97910
rect -10360 97980 -10140 98000
rect -10360 97910 -10350 97980
rect -10150 97910 -10140 97980
rect -10360 97860 -10140 97910
rect -9860 97980 -9640 98000
rect -9860 97910 -9850 97980
rect -9650 97910 -9640 97980
rect -9860 97860 -9640 97910
rect -9360 97980 -9140 98000
rect -9360 97910 -9350 97980
rect -9150 97910 -9140 97980
rect -9360 97860 -9140 97910
rect -8860 97980 -8640 98000
rect -8860 97910 -8850 97980
rect -8650 97910 -8640 97980
rect -8860 97860 -8640 97910
rect -8360 97980 -8140 98000
rect -8360 97910 -8350 97980
rect -8150 97910 -8140 97980
rect -8360 97860 -8140 97910
rect -7860 97980 -7640 98000
rect -7860 97910 -7850 97980
rect -7650 97910 -7640 97980
rect -7860 97860 -7640 97910
rect -7360 97980 -7140 98000
rect -7360 97910 -7350 97980
rect -7150 97910 -7140 97980
rect -7360 97860 -7140 97910
rect -6860 97980 -6640 98000
rect -6860 97910 -6850 97980
rect -6650 97910 -6640 97980
rect -6860 97860 -6640 97910
rect -6360 97980 -6140 98000
rect -6360 97910 -6350 97980
rect -6150 97910 -6140 97980
rect -6360 97860 -6140 97910
rect -5860 97980 -5640 98000
rect -5860 97910 -5850 97980
rect -5650 97910 -5640 97980
rect -5860 97860 -5640 97910
rect -5360 97980 -5140 98000
rect -5360 97910 -5350 97980
rect -5150 97910 -5140 97980
rect -5360 97860 -5140 97910
rect -4860 97980 -4640 98000
rect -4860 97910 -4850 97980
rect -4650 97910 -4640 97980
rect -4860 97860 -4640 97910
rect -4360 97980 -4140 98000
rect -4360 97910 -4350 97980
rect -4150 97910 -4140 97980
rect -4360 97860 -4140 97910
rect -3860 97980 -3640 98000
rect -3860 97910 -3850 97980
rect -3650 97910 -3640 97980
rect -3860 97860 -3640 97910
rect -3360 97980 -3140 98000
rect -3360 97910 -3350 97980
rect -3150 97910 -3140 97980
rect -3360 97860 -3140 97910
rect -2860 97980 -2640 98000
rect -2860 97910 -2850 97980
rect -2650 97910 -2640 97980
rect -2860 97860 -2640 97910
rect -2360 97980 -2140 98000
rect -2360 97910 -2350 97980
rect -2150 97910 -2140 97980
rect -2360 97860 -2140 97910
rect -1860 97980 -1640 98000
rect -1860 97910 -1850 97980
rect -1650 97910 -1640 97980
rect -1860 97860 -1640 97910
rect -1360 97980 -1140 98000
rect -1360 97910 -1350 97980
rect -1150 97910 -1140 97980
rect -1360 97860 -1140 97910
rect -860 97980 -640 98000
rect -860 97910 -850 97980
rect -650 97910 -640 97980
rect -860 97860 -640 97910
rect -360 97980 -140 98000
rect -360 97910 -350 97980
rect -150 97910 -140 97980
rect -360 97860 -140 97910
rect 140 97980 360 98000
rect 140 97910 150 97980
rect 350 97910 360 97980
rect 140 97860 360 97910
rect 640 97980 860 98000
rect 640 97910 650 97980
rect 850 97910 860 97980
rect 640 97860 860 97910
rect 1140 97980 1360 98000
rect 1140 97910 1150 97980
rect 1350 97910 1360 97980
rect 1140 97860 1360 97910
rect 1640 97980 1860 98000
rect 1640 97910 1650 97980
rect 1850 97910 1860 97980
rect 1640 97860 1860 97910
rect 2140 97980 2360 98000
rect 2140 97910 2150 97980
rect 2350 97910 2360 97980
rect 2140 97860 2360 97910
rect 2640 97980 2860 98000
rect 2640 97910 2650 97980
rect 2850 97910 2860 97980
rect 2640 97860 2860 97910
rect 3140 97980 3360 98000
rect 3140 97910 3150 97980
rect 3350 97910 3360 97980
rect 3140 97860 3360 97910
rect 3640 97980 3860 98000
rect 3640 97910 3650 97980
rect 3850 97910 3860 97980
rect 3640 97860 3860 97910
rect 4140 97980 4360 98000
rect 4140 97910 4150 97980
rect 4350 97910 4360 97980
rect 4140 97860 4360 97910
rect 4640 97980 4860 98000
rect 4640 97910 4650 97980
rect 4850 97910 4860 97980
rect 4640 97860 4860 97910
rect 5140 97980 5360 98000
rect 5140 97910 5150 97980
rect 5350 97910 5360 97980
rect 5140 97860 5360 97910
rect 5640 97980 5860 98000
rect 5640 97910 5650 97980
rect 5850 97910 5860 97980
rect 5640 97860 5860 97910
rect 6140 97980 6360 98000
rect 6140 97910 6150 97980
rect 6350 97910 6360 97980
rect 6140 97860 6360 97910
rect 6640 97980 6860 98000
rect 6640 97910 6650 97980
rect 6850 97910 6860 97980
rect 6640 97860 6860 97910
rect 7140 97980 7360 98000
rect 7140 97910 7150 97980
rect 7350 97910 7360 97980
rect 7140 97860 7360 97910
rect 7640 97980 7860 98000
rect 7640 97910 7650 97980
rect 7850 97910 7860 97980
rect 7640 97860 7860 97910
rect 8140 97980 8360 98000
rect 8140 97910 8150 97980
rect 8350 97910 8360 97980
rect 8140 97860 8360 97910
rect 8640 97980 8860 98000
rect 8640 97910 8650 97980
rect 8850 97910 8860 97980
rect 8640 97860 8860 97910
rect 9140 97980 9360 98000
rect 9140 97910 9150 97980
rect 9350 97910 9360 97980
rect 9140 97860 9360 97910
rect 9640 97980 9860 98000
rect 9640 97910 9650 97980
rect 9850 97910 9860 97980
rect 9640 97860 9860 97910
rect 10140 97980 10360 98000
rect 10140 97910 10150 97980
rect 10350 97910 10360 97980
rect 10140 97860 10360 97910
rect 10640 97980 10860 98000
rect 10640 97910 10650 97980
rect 10850 97910 10860 97980
rect 10640 97860 10860 97910
rect 11140 97980 11360 98000
rect 11140 97910 11150 97980
rect 11350 97910 11360 97980
rect 11140 97860 11360 97910
rect 11640 97980 11860 98000
rect 11640 97910 11650 97980
rect 11850 97910 11860 97980
rect 11640 97860 11860 97910
rect 12140 97980 12360 98000
rect 12140 97910 12150 97980
rect 12350 97910 12360 97980
rect 12140 97860 12360 97910
rect 12640 97980 12860 98000
rect 12640 97910 12650 97980
rect 12850 97910 12860 97980
rect 12640 97860 12860 97910
rect 13140 97980 13360 98000
rect 13140 97910 13150 97980
rect 13350 97910 13360 97980
rect 13140 97860 13360 97910
rect 13640 97980 13860 98000
rect 13640 97910 13650 97980
rect 13850 97910 13860 97980
rect 13640 97860 13860 97910
rect 14140 97980 14360 98000
rect 14140 97910 14150 97980
rect 14350 97910 14360 97980
rect 14140 97860 14360 97910
rect 14640 97980 14860 98000
rect 14640 97910 14650 97980
rect 14850 97910 14860 97980
rect 14640 97860 14860 97910
rect 15140 97980 15360 98000
rect 15140 97910 15150 97980
rect 15350 97910 15360 97980
rect 15140 97860 15360 97910
rect 15640 97980 15860 98000
rect 15640 97910 15650 97980
rect 15850 97910 15860 97980
rect 15640 97860 15860 97910
rect 16140 97980 16360 98000
rect 16140 97910 16150 97980
rect 16350 97910 16360 97980
rect 16140 97860 16360 97910
rect 16640 97980 16860 98000
rect 16640 97910 16650 97980
rect 16850 97910 16860 97980
rect 16640 97860 16860 97910
rect 17140 97980 17360 98000
rect 17140 97910 17150 97980
rect 17350 97910 17360 97980
rect 17140 97860 17360 97910
rect 17640 97980 17860 98000
rect 17640 97910 17650 97980
rect 17850 97910 17860 97980
rect 17640 97860 17860 97910
rect 18140 97980 18360 98000
rect 18140 97910 18150 97980
rect 18350 97910 18360 97980
rect 18140 97860 18360 97910
rect 18640 97980 18860 98000
rect 18640 97910 18650 97980
rect 18850 97910 18860 97980
rect 18640 97860 18860 97910
rect 19140 97980 19360 98000
rect 19140 97910 19150 97980
rect 19350 97910 19360 97980
rect 19140 97860 19360 97910
rect 19640 97980 19860 98000
rect 19640 97910 19650 97980
rect 19850 97910 19860 97980
rect 19640 97860 19860 97910
rect -16000 97850 20000 97860
rect -16000 97650 -15980 97850
rect -15910 97650 -15590 97850
rect -15520 97650 -15480 97850
rect -15410 97650 -15090 97850
rect -15020 97650 -14980 97850
rect -14910 97650 -14590 97850
rect -14520 97650 -14480 97850
rect -14410 97650 -14090 97850
rect -14020 97650 -13980 97850
rect -13910 97650 -13590 97850
rect -13520 97650 -13480 97850
rect -13410 97650 -13090 97850
rect -13020 97650 -12980 97850
rect -12910 97650 -12590 97850
rect -12520 97650 -12480 97850
rect -12410 97650 -12090 97850
rect -12020 97650 -11980 97850
rect -11910 97650 -11590 97850
rect -11520 97650 -11480 97850
rect -11410 97650 -11090 97850
rect -11020 97650 -10980 97850
rect -10910 97650 -10590 97850
rect -10520 97650 -10480 97850
rect -10410 97650 -10090 97850
rect -10020 97650 -9980 97850
rect -9910 97650 -9590 97850
rect -9520 97650 -9480 97850
rect -9410 97650 -9090 97850
rect -9020 97650 -8980 97850
rect -8910 97650 -8590 97850
rect -8520 97650 -8480 97850
rect -8410 97650 -8090 97850
rect -8020 97650 -7980 97850
rect -7910 97650 -7590 97850
rect -7520 97650 -7480 97850
rect -7410 97650 -7090 97850
rect -7020 97650 -6980 97850
rect -6910 97650 -6590 97850
rect -6520 97650 -6480 97850
rect -6410 97650 -6090 97850
rect -6020 97650 -5980 97850
rect -5910 97650 -5590 97850
rect -5520 97650 -5480 97850
rect -5410 97650 -5090 97850
rect -5020 97650 -4980 97850
rect -4910 97650 -4590 97850
rect -4520 97650 -4480 97850
rect -4410 97650 -4090 97850
rect -4020 97650 -3980 97850
rect -3910 97650 -3590 97850
rect -3520 97650 -3480 97850
rect -3410 97650 -3090 97850
rect -3020 97650 -2980 97850
rect -2910 97650 -2590 97850
rect -2520 97650 -2480 97850
rect -2410 97650 -2090 97850
rect -2020 97650 -1980 97850
rect -1910 97650 -1590 97850
rect -1520 97650 -1480 97850
rect -1410 97650 -1090 97850
rect -1020 97650 -980 97850
rect -910 97650 -590 97850
rect -520 97650 -480 97850
rect -410 97650 -90 97850
rect -20 97650 20 97850
rect 90 97650 410 97850
rect 480 97650 520 97850
rect 590 97650 910 97850
rect 980 97650 1020 97850
rect 1090 97650 1410 97850
rect 1480 97650 1520 97850
rect 1590 97650 1910 97850
rect 1980 97650 2020 97850
rect 2090 97650 2410 97850
rect 2480 97650 2520 97850
rect 2590 97650 2910 97850
rect 2980 97650 3020 97850
rect 3090 97650 3410 97850
rect 3480 97650 3520 97850
rect 3590 97650 3910 97850
rect 3980 97650 4020 97850
rect 4090 97650 4410 97850
rect 4480 97650 4520 97850
rect 4590 97650 4910 97850
rect 4980 97650 5020 97850
rect 5090 97650 5410 97850
rect 5480 97650 5520 97850
rect 5590 97650 5910 97850
rect 5980 97650 6020 97850
rect 6090 97650 6410 97850
rect 6480 97650 6520 97850
rect 6590 97650 6910 97850
rect 6980 97650 7020 97850
rect 7090 97650 7410 97850
rect 7480 97650 7520 97850
rect 7590 97650 7910 97850
rect 7980 97650 8020 97850
rect 8090 97650 8410 97850
rect 8480 97650 8520 97850
rect 8590 97650 8910 97850
rect 8980 97650 9020 97850
rect 9090 97650 9410 97850
rect 9480 97650 9520 97850
rect 9590 97650 9910 97850
rect 9980 97650 10020 97850
rect 10090 97650 10410 97850
rect 10480 97650 10520 97850
rect 10590 97650 10910 97850
rect 10980 97650 11020 97850
rect 11090 97650 11410 97850
rect 11480 97650 11520 97850
rect 11590 97650 11910 97850
rect 11980 97650 12020 97850
rect 12090 97650 12410 97850
rect 12480 97650 12520 97850
rect 12590 97650 12910 97850
rect 12980 97650 13020 97850
rect 13090 97650 13410 97850
rect 13480 97650 13520 97850
rect 13590 97650 13910 97850
rect 13980 97650 14020 97850
rect 14090 97650 14410 97850
rect 14480 97650 14520 97850
rect 14590 97650 14910 97850
rect 14980 97650 15020 97850
rect 15090 97650 15410 97850
rect 15480 97650 15520 97850
rect 15590 97650 15910 97850
rect 15980 97650 16020 97850
rect 16090 97650 16410 97850
rect 16480 97650 16520 97850
rect 16590 97650 16910 97850
rect 16980 97650 17020 97850
rect 17090 97650 17410 97850
rect 17480 97650 17520 97850
rect 17590 97650 17910 97850
rect 17980 97650 18020 97850
rect 18090 97650 18410 97850
rect 18480 97650 18520 97850
rect 18590 97650 18910 97850
rect 18980 97650 19020 97850
rect 19090 97650 19410 97850
rect 19480 97650 19520 97850
rect 19590 97650 19910 97850
rect 19980 97650 20000 97850
rect -16000 97640 20000 97650
rect -15860 97590 -15640 97640
rect -15860 97520 -15850 97590
rect -15650 97520 -15640 97590
rect -15860 97480 -15640 97520
rect -15860 97410 -15850 97480
rect -15650 97410 -15640 97480
rect -15860 97360 -15640 97410
rect -15360 97590 -15140 97640
rect -15360 97520 -15350 97590
rect -15150 97520 -15140 97590
rect -15360 97480 -15140 97520
rect -15360 97410 -15350 97480
rect -15150 97410 -15140 97480
rect -15360 97360 -15140 97410
rect -14860 97590 -14640 97640
rect -14860 97520 -14850 97590
rect -14650 97520 -14640 97590
rect -14860 97480 -14640 97520
rect -14860 97410 -14850 97480
rect -14650 97410 -14640 97480
rect -14860 97360 -14640 97410
rect -14360 97590 -14140 97640
rect -14360 97520 -14350 97590
rect -14150 97520 -14140 97590
rect -14360 97480 -14140 97520
rect -14360 97410 -14350 97480
rect -14150 97410 -14140 97480
rect -14360 97360 -14140 97410
rect -13860 97590 -13640 97640
rect -13860 97520 -13850 97590
rect -13650 97520 -13640 97590
rect -13860 97480 -13640 97520
rect -13860 97410 -13850 97480
rect -13650 97410 -13640 97480
rect -13860 97360 -13640 97410
rect -13360 97590 -13140 97640
rect -13360 97520 -13350 97590
rect -13150 97520 -13140 97590
rect -13360 97480 -13140 97520
rect -13360 97410 -13350 97480
rect -13150 97410 -13140 97480
rect -13360 97360 -13140 97410
rect -12860 97590 -12640 97640
rect -12860 97520 -12850 97590
rect -12650 97520 -12640 97590
rect -12860 97480 -12640 97520
rect -12860 97410 -12850 97480
rect -12650 97410 -12640 97480
rect -12860 97360 -12640 97410
rect -12360 97590 -12140 97640
rect -12360 97520 -12350 97590
rect -12150 97520 -12140 97590
rect -12360 97480 -12140 97520
rect -12360 97410 -12350 97480
rect -12150 97410 -12140 97480
rect -12360 97360 -12140 97410
rect -11860 97590 -11640 97640
rect -11860 97520 -11850 97590
rect -11650 97520 -11640 97590
rect -11860 97480 -11640 97520
rect -11860 97410 -11850 97480
rect -11650 97410 -11640 97480
rect -11860 97360 -11640 97410
rect -11360 97590 -11140 97640
rect -11360 97520 -11350 97590
rect -11150 97520 -11140 97590
rect -11360 97480 -11140 97520
rect -11360 97410 -11350 97480
rect -11150 97410 -11140 97480
rect -11360 97360 -11140 97410
rect -10860 97590 -10640 97640
rect -10860 97520 -10850 97590
rect -10650 97520 -10640 97590
rect -10860 97480 -10640 97520
rect -10860 97410 -10850 97480
rect -10650 97410 -10640 97480
rect -10860 97360 -10640 97410
rect -10360 97590 -10140 97640
rect -10360 97520 -10350 97590
rect -10150 97520 -10140 97590
rect -10360 97480 -10140 97520
rect -10360 97410 -10350 97480
rect -10150 97410 -10140 97480
rect -10360 97360 -10140 97410
rect -9860 97590 -9640 97640
rect -9860 97520 -9850 97590
rect -9650 97520 -9640 97590
rect -9860 97480 -9640 97520
rect -9860 97410 -9850 97480
rect -9650 97410 -9640 97480
rect -9860 97360 -9640 97410
rect -9360 97590 -9140 97640
rect -9360 97520 -9350 97590
rect -9150 97520 -9140 97590
rect -9360 97480 -9140 97520
rect -9360 97410 -9350 97480
rect -9150 97410 -9140 97480
rect -9360 97360 -9140 97410
rect -8860 97590 -8640 97640
rect -8860 97520 -8850 97590
rect -8650 97520 -8640 97590
rect -8860 97480 -8640 97520
rect -8860 97410 -8850 97480
rect -8650 97410 -8640 97480
rect -8860 97360 -8640 97410
rect -8360 97590 -8140 97640
rect -8360 97520 -8350 97590
rect -8150 97520 -8140 97590
rect -8360 97480 -8140 97520
rect -8360 97410 -8350 97480
rect -8150 97410 -8140 97480
rect -8360 97360 -8140 97410
rect -7860 97590 -7640 97640
rect -7860 97520 -7850 97590
rect -7650 97520 -7640 97590
rect -7860 97480 -7640 97520
rect -7860 97410 -7850 97480
rect -7650 97410 -7640 97480
rect -7860 97360 -7640 97410
rect -7360 97590 -7140 97640
rect -7360 97520 -7350 97590
rect -7150 97520 -7140 97590
rect -7360 97480 -7140 97520
rect -7360 97410 -7350 97480
rect -7150 97410 -7140 97480
rect -7360 97360 -7140 97410
rect -6860 97590 -6640 97640
rect -6860 97520 -6850 97590
rect -6650 97520 -6640 97590
rect -6860 97480 -6640 97520
rect -6860 97410 -6850 97480
rect -6650 97410 -6640 97480
rect -6860 97360 -6640 97410
rect -6360 97590 -6140 97640
rect -6360 97520 -6350 97590
rect -6150 97520 -6140 97590
rect -6360 97480 -6140 97520
rect -6360 97410 -6350 97480
rect -6150 97410 -6140 97480
rect -6360 97360 -6140 97410
rect -5860 97590 -5640 97640
rect -5860 97520 -5850 97590
rect -5650 97520 -5640 97590
rect -5860 97480 -5640 97520
rect -5860 97410 -5850 97480
rect -5650 97410 -5640 97480
rect -5860 97360 -5640 97410
rect -5360 97590 -5140 97640
rect -5360 97520 -5350 97590
rect -5150 97520 -5140 97590
rect -5360 97480 -5140 97520
rect -5360 97410 -5350 97480
rect -5150 97410 -5140 97480
rect -5360 97360 -5140 97410
rect -4860 97590 -4640 97640
rect -4860 97520 -4850 97590
rect -4650 97520 -4640 97590
rect -4860 97480 -4640 97520
rect -4860 97410 -4850 97480
rect -4650 97410 -4640 97480
rect -4860 97360 -4640 97410
rect -4360 97590 -4140 97640
rect -4360 97520 -4350 97590
rect -4150 97520 -4140 97590
rect -4360 97480 -4140 97520
rect -4360 97410 -4350 97480
rect -4150 97410 -4140 97480
rect -4360 97360 -4140 97410
rect -3860 97590 -3640 97640
rect -3860 97520 -3850 97590
rect -3650 97520 -3640 97590
rect -3860 97480 -3640 97520
rect -3860 97410 -3850 97480
rect -3650 97410 -3640 97480
rect -3860 97360 -3640 97410
rect -3360 97590 -3140 97640
rect -3360 97520 -3350 97590
rect -3150 97520 -3140 97590
rect -3360 97480 -3140 97520
rect -3360 97410 -3350 97480
rect -3150 97410 -3140 97480
rect -3360 97360 -3140 97410
rect -2860 97590 -2640 97640
rect -2860 97520 -2850 97590
rect -2650 97520 -2640 97590
rect -2860 97480 -2640 97520
rect -2860 97410 -2850 97480
rect -2650 97410 -2640 97480
rect -2860 97360 -2640 97410
rect -2360 97590 -2140 97640
rect -2360 97520 -2350 97590
rect -2150 97520 -2140 97590
rect -2360 97480 -2140 97520
rect -2360 97410 -2350 97480
rect -2150 97410 -2140 97480
rect -2360 97360 -2140 97410
rect -1860 97590 -1640 97640
rect -1860 97520 -1850 97590
rect -1650 97520 -1640 97590
rect -1860 97480 -1640 97520
rect -1860 97410 -1850 97480
rect -1650 97410 -1640 97480
rect -1860 97360 -1640 97410
rect -1360 97590 -1140 97640
rect -1360 97520 -1350 97590
rect -1150 97520 -1140 97590
rect -1360 97480 -1140 97520
rect -1360 97410 -1350 97480
rect -1150 97410 -1140 97480
rect -1360 97360 -1140 97410
rect -860 97590 -640 97640
rect -860 97520 -850 97590
rect -650 97520 -640 97590
rect -860 97480 -640 97520
rect -860 97410 -850 97480
rect -650 97410 -640 97480
rect -860 97360 -640 97410
rect -360 97590 -140 97640
rect -360 97520 -350 97590
rect -150 97520 -140 97590
rect -360 97480 -140 97520
rect -360 97410 -350 97480
rect -150 97410 -140 97480
rect -360 97360 -140 97410
rect 140 97590 360 97640
rect 140 97520 150 97590
rect 350 97520 360 97590
rect 140 97480 360 97520
rect 140 97410 150 97480
rect 350 97410 360 97480
rect 140 97360 360 97410
rect 640 97590 860 97640
rect 640 97520 650 97590
rect 850 97520 860 97590
rect 640 97480 860 97520
rect 640 97410 650 97480
rect 850 97410 860 97480
rect 640 97360 860 97410
rect 1140 97590 1360 97640
rect 1140 97520 1150 97590
rect 1350 97520 1360 97590
rect 1140 97480 1360 97520
rect 1140 97410 1150 97480
rect 1350 97410 1360 97480
rect 1140 97360 1360 97410
rect 1640 97590 1860 97640
rect 1640 97520 1650 97590
rect 1850 97520 1860 97590
rect 1640 97480 1860 97520
rect 1640 97410 1650 97480
rect 1850 97410 1860 97480
rect 1640 97360 1860 97410
rect 2140 97590 2360 97640
rect 2140 97520 2150 97590
rect 2350 97520 2360 97590
rect 2140 97480 2360 97520
rect 2140 97410 2150 97480
rect 2350 97410 2360 97480
rect 2140 97360 2360 97410
rect 2640 97590 2860 97640
rect 2640 97520 2650 97590
rect 2850 97520 2860 97590
rect 2640 97480 2860 97520
rect 2640 97410 2650 97480
rect 2850 97410 2860 97480
rect 2640 97360 2860 97410
rect 3140 97590 3360 97640
rect 3140 97520 3150 97590
rect 3350 97520 3360 97590
rect 3140 97480 3360 97520
rect 3140 97410 3150 97480
rect 3350 97410 3360 97480
rect 3140 97360 3360 97410
rect 3640 97590 3860 97640
rect 3640 97520 3650 97590
rect 3850 97520 3860 97590
rect 3640 97480 3860 97520
rect 3640 97410 3650 97480
rect 3850 97410 3860 97480
rect 3640 97360 3860 97410
rect 4140 97590 4360 97640
rect 4140 97520 4150 97590
rect 4350 97520 4360 97590
rect 4140 97480 4360 97520
rect 4140 97410 4150 97480
rect 4350 97410 4360 97480
rect 4140 97360 4360 97410
rect 4640 97590 4860 97640
rect 4640 97520 4650 97590
rect 4850 97520 4860 97590
rect 4640 97480 4860 97520
rect 4640 97410 4650 97480
rect 4850 97410 4860 97480
rect 4640 97360 4860 97410
rect 5140 97590 5360 97640
rect 5140 97520 5150 97590
rect 5350 97520 5360 97590
rect 5140 97480 5360 97520
rect 5140 97410 5150 97480
rect 5350 97410 5360 97480
rect 5140 97360 5360 97410
rect 5640 97590 5860 97640
rect 5640 97520 5650 97590
rect 5850 97520 5860 97590
rect 5640 97480 5860 97520
rect 5640 97410 5650 97480
rect 5850 97410 5860 97480
rect 5640 97360 5860 97410
rect 6140 97590 6360 97640
rect 6140 97520 6150 97590
rect 6350 97520 6360 97590
rect 6140 97480 6360 97520
rect 6140 97410 6150 97480
rect 6350 97410 6360 97480
rect 6140 97360 6360 97410
rect 6640 97590 6860 97640
rect 6640 97520 6650 97590
rect 6850 97520 6860 97590
rect 6640 97480 6860 97520
rect 6640 97410 6650 97480
rect 6850 97410 6860 97480
rect 6640 97360 6860 97410
rect 7140 97590 7360 97640
rect 7140 97520 7150 97590
rect 7350 97520 7360 97590
rect 7140 97480 7360 97520
rect 7140 97410 7150 97480
rect 7350 97410 7360 97480
rect 7140 97360 7360 97410
rect 7640 97590 7860 97640
rect 7640 97520 7650 97590
rect 7850 97520 7860 97590
rect 7640 97480 7860 97520
rect 7640 97410 7650 97480
rect 7850 97410 7860 97480
rect 7640 97360 7860 97410
rect 8140 97590 8360 97640
rect 8140 97520 8150 97590
rect 8350 97520 8360 97590
rect 8140 97480 8360 97520
rect 8140 97410 8150 97480
rect 8350 97410 8360 97480
rect 8140 97360 8360 97410
rect 8640 97590 8860 97640
rect 8640 97520 8650 97590
rect 8850 97520 8860 97590
rect 8640 97480 8860 97520
rect 8640 97410 8650 97480
rect 8850 97410 8860 97480
rect 8640 97360 8860 97410
rect 9140 97590 9360 97640
rect 9140 97520 9150 97590
rect 9350 97520 9360 97590
rect 9140 97480 9360 97520
rect 9140 97410 9150 97480
rect 9350 97410 9360 97480
rect 9140 97360 9360 97410
rect 9640 97590 9860 97640
rect 9640 97520 9650 97590
rect 9850 97520 9860 97590
rect 9640 97480 9860 97520
rect 9640 97410 9650 97480
rect 9850 97410 9860 97480
rect 9640 97360 9860 97410
rect 10140 97590 10360 97640
rect 10140 97520 10150 97590
rect 10350 97520 10360 97590
rect 10140 97480 10360 97520
rect 10140 97410 10150 97480
rect 10350 97410 10360 97480
rect 10140 97360 10360 97410
rect 10640 97590 10860 97640
rect 10640 97520 10650 97590
rect 10850 97520 10860 97590
rect 10640 97480 10860 97520
rect 10640 97410 10650 97480
rect 10850 97410 10860 97480
rect 10640 97360 10860 97410
rect 11140 97590 11360 97640
rect 11140 97520 11150 97590
rect 11350 97520 11360 97590
rect 11140 97480 11360 97520
rect 11140 97410 11150 97480
rect 11350 97410 11360 97480
rect 11140 97360 11360 97410
rect 11640 97590 11860 97640
rect 11640 97520 11650 97590
rect 11850 97520 11860 97590
rect 11640 97480 11860 97520
rect 11640 97410 11650 97480
rect 11850 97410 11860 97480
rect 11640 97360 11860 97410
rect 12140 97590 12360 97640
rect 12140 97520 12150 97590
rect 12350 97520 12360 97590
rect 12140 97480 12360 97520
rect 12140 97410 12150 97480
rect 12350 97410 12360 97480
rect 12140 97360 12360 97410
rect 12640 97590 12860 97640
rect 12640 97520 12650 97590
rect 12850 97520 12860 97590
rect 12640 97480 12860 97520
rect 12640 97410 12650 97480
rect 12850 97410 12860 97480
rect 12640 97360 12860 97410
rect 13140 97590 13360 97640
rect 13140 97520 13150 97590
rect 13350 97520 13360 97590
rect 13140 97480 13360 97520
rect 13140 97410 13150 97480
rect 13350 97410 13360 97480
rect 13140 97360 13360 97410
rect 13640 97590 13860 97640
rect 13640 97520 13650 97590
rect 13850 97520 13860 97590
rect 13640 97480 13860 97520
rect 13640 97410 13650 97480
rect 13850 97410 13860 97480
rect 13640 97360 13860 97410
rect 14140 97590 14360 97640
rect 14140 97520 14150 97590
rect 14350 97520 14360 97590
rect 14140 97480 14360 97520
rect 14140 97410 14150 97480
rect 14350 97410 14360 97480
rect 14140 97360 14360 97410
rect 14640 97590 14860 97640
rect 14640 97520 14650 97590
rect 14850 97520 14860 97590
rect 14640 97480 14860 97520
rect 14640 97410 14650 97480
rect 14850 97410 14860 97480
rect 14640 97360 14860 97410
rect 15140 97590 15360 97640
rect 15140 97520 15150 97590
rect 15350 97520 15360 97590
rect 15140 97480 15360 97520
rect 15140 97410 15150 97480
rect 15350 97410 15360 97480
rect 15140 97360 15360 97410
rect 15640 97590 15860 97640
rect 15640 97520 15650 97590
rect 15850 97520 15860 97590
rect 15640 97480 15860 97520
rect 15640 97410 15650 97480
rect 15850 97410 15860 97480
rect 15640 97360 15860 97410
rect 16140 97590 16360 97640
rect 16140 97520 16150 97590
rect 16350 97520 16360 97590
rect 16140 97480 16360 97520
rect 16140 97410 16150 97480
rect 16350 97410 16360 97480
rect 16140 97360 16360 97410
rect 16640 97590 16860 97640
rect 16640 97520 16650 97590
rect 16850 97520 16860 97590
rect 16640 97480 16860 97520
rect 16640 97410 16650 97480
rect 16850 97410 16860 97480
rect 16640 97360 16860 97410
rect 17140 97590 17360 97640
rect 17140 97520 17150 97590
rect 17350 97520 17360 97590
rect 17140 97480 17360 97520
rect 17140 97410 17150 97480
rect 17350 97410 17360 97480
rect 17140 97360 17360 97410
rect 17640 97590 17860 97640
rect 17640 97520 17650 97590
rect 17850 97520 17860 97590
rect 17640 97480 17860 97520
rect 17640 97410 17650 97480
rect 17850 97410 17860 97480
rect 17640 97360 17860 97410
rect 18140 97590 18360 97640
rect 18140 97520 18150 97590
rect 18350 97520 18360 97590
rect 18140 97480 18360 97520
rect 18140 97410 18150 97480
rect 18350 97410 18360 97480
rect 18140 97360 18360 97410
rect 18640 97590 18860 97640
rect 18640 97520 18650 97590
rect 18850 97520 18860 97590
rect 18640 97480 18860 97520
rect 18640 97410 18650 97480
rect 18850 97410 18860 97480
rect 18640 97360 18860 97410
rect 19140 97590 19360 97640
rect 19140 97520 19150 97590
rect 19350 97520 19360 97590
rect 19140 97480 19360 97520
rect 19140 97410 19150 97480
rect 19350 97410 19360 97480
rect 19140 97360 19360 97410
rect 19640 97590 19860 97640
rect 19640 97520 19650 97590
rect 19850 97520 19860 97590
rect 19640 97480 19860 97520
rect 19640 97410 19650 97480
rect 19850 97410 19860 97480
rect 19640 97360 19860 97410
rect -16000 97350 20000 97360
rect -16000 97150 -15980 97350
rect -15910 97150 -15590 97350
rect -15520 97150 -15480 97350
rect -15410 97150 -15090 97350
rect -15020 97150 -14980 97350
rect -14910 97150 -14590 97350
rect -14520 97150 -14480 97350
rect -14410 97150 -14090 97350
rect -14020 97150 -13980 97350
rect -13910 97150 -13590 97350
rect -13520 97150 -13480 97350
rect -13410 97150 -13090 97350
rect -13020 97150 -12980 97350
rect -12910 97150 -12590 97350
rect -12520 97150 -12480 97350
rect -12410 97150 -12090 97350
rect -12020 97150 -11980 97350
rect -11910 97150 -11590 97350
rect -11520 97150 -11480 97350
rect -11410 97150 -11090 97350
rect -11020 97150 -10980 97350
rect -10910 97150 -10590 97350
rect -10520 97150 -10480 97350
rect -10410 97150 -10090 97350
rect -10020 97150 -9980 97350
rect -9910 97150 -9590 97350
rect -9520 97150 -9480 97350
rect -9410 97150 -9090 97350
rect -9020 97150 -8980 97350
rect -8910 97150 -8590 97350
rect -8520 97150 -8480 97350
rect -8410 97150 -8090 97350
rect -8020 97150 -7980 97350
rect -7910 97150 -7590 97350
rect -7520 97150 -7480 97350
rect -7410 97150 -7090 97350
rect -7020 97150 -6980 97350
rect -6910 97150 -6590 97350
rect -6520 97150 -6480 97350
rect -6410 97150 -6090 97350
rect -6020 97150 -5980 97350
rect -5910 97150 -5590 97350
rect -5520 97150 -5480 97350
rect -5410 97150 -5090 97350
rect -5020 97150 -4980 97350
rect -4910 97150 -4590 97350
rect -4520 97150 -4480 97350
rect -4410 97150 -4090 97350
rect -4020 97150 -3980 97350
rect -3910 97150 -3590 97350
rect -3520 97150 -3480 97350
rect -3410 97150 -3090 97350
rect -3020 97150 -2980 97350
rect -2910 97150 -2590 97350
rect -2520 97150 -2480 97350
rect -2410 97150 -2090 97350
rect -2020 97150 -1980 97350
rect -1910 97150 -1590 97350
rect -1520 97150 -1480 97350
rect -1410 97150 -1090 97350
rect -1020 97150 -980 97350
rect -910 97150 -590 97350
rect -520 97150 -480 97350
rect -410 97150 -90 97350
rect -20 97150 20 97350
rect 90 97150 410 97350
rect 480 97150 520 97350
rect 590 97150 910 97350
rect 980 97150 1020 97350
rect 1090 97150 1410 97350
rect 1480 97150 1520 97350
rect 1590 97150 1910 97350
rect 1980 97150 2020 97350
rect 2090 97150 2410 97350
rect 2480 97150 2520 97350
rect 2590 97150 2910 97350
rect 2980 97150 3020 97350
rect 3090 97150 3410 97350
rect 3480 97150 3520 97350
rect 3590 97150 3910 97350
rect 3980 97150 4020 97350
rect 4090 97150 4410 97350
rect 4480 97150 4520 97350
rect 4590 97150 4910 97350
rect 4980 97150 5020 97350
rect 5090 97150 5410 97350
rect 5480 97150 5520 97350
rect 5590 97150 5910 97350
rect 5980 97150 6020 97350
rect 6090 97150 6410 97350
rect 6480 97150 6520 97350
rect 6590 97150 6910 97350
rect 6980 97150 7020 97350
rect 7090 97150 7410 97350
rect 7480 97150 7520 97350
rect 7590 97150 7910 97350
rect 7980 97150 8020 97350
rect 8090 97150 8410 97350
rect 8480 97150 8520 97350
rect 8590 97150 8910 97350
rect 8980 97150 9020 97350
rect 9090 97150 9410 97350
rect 9480 97150 9520 97350
rect 9590 97150 9910 97350
rect 9980 97150 10020 97350
rect 10090 97150 10410 97350
rect 10480 97150 10520 97350
rect 10590 97150 10910 97350
rect 10980 97150 11020 97350
rect 11090 97150 11410 97350
rect 11480 97150 11520 97350
rect 11590 97150 11910 97350
rect 11980 97150 12020 97350
rect 12090 97150 12410 97350
rect 12480 97150 12520 97350
rect 12590 97150 12910 97350
rect 12980 97150 13020 97350
rect 13090 97150 13410 97350
rect 13480 97150 13520 97350
rect 13590 97150 13910 97350
rect 13980 97150 14020 97350
rect 14090 97150 14410 97350
rect 14480 97150 14520 97350
rect 14590 97150 14910 97350
rect 14980 97150 15020 97350
rect 15090 97150 15410 97350
rect 15480 97150 15520 97350
rect 15590 97150 15910 97350
rect 15980 97150 16020 97350
rect 16090 97150 16410 97350
rect 16480 97150 16520 97350
rect 16590 97150 16910 97350
rect 16980 97150 17020 97350
rect 17090 97150 17410 97350
rect 17480 97150 17520 97350
rect 17590 97150 17910 97350
rect 17980 97150 18020 97350
rect 18090 97150 18410 97350
rect 18480 97150 18520 97350
rect 18590 97150 18910 97350
rect 18980 97150 19020 97350
rect 19090 97150 19410 97350
rect 19480 97150 19520 97350
rect 19590 97150 19910 97350
rect 19980 97150 20000 97350
rect -16000 97140 20000 97150
rect -15860 97090 -15640 97140
rect -15860 97020 -15850 97090
rect -15650 97020 -15640 97090
rect -15860 96980 -15640 97020
rect -15860 96910 -15850 96980
rect -15650 96910 -15640 96980
rect -15860 96860 -15640 96910
rect -15360 97090 -15140 97140
rect -15360 97020 -15350 97090
rect -15150 97020 -15140 97090
rect -15360 96980 -15140 97020
rect -15360 96910 -15350 96980
rect -15150 96910 -15140 96980
rect -15360 96860 -15140 96910
rect -14860 97090 -14640 97140
rect -14860 97020 -14850 97090
rect -14650 97020 -14640 97090
rect -14860 96980 -14640 97020
rect -14860 96910 -14850 96980
rect -14650 96910 -14640 96980
rect -14860 96860 -14640 96910
rect -14360 97090 -14140 97140
rect -14360 97020 -14350 97090
rect -14150 97020 -14140 97090
rect -14360 96980 -14140 97020
rect -14360 96910 -14350 96980
rect -14150 96910 -14140 96980
rect -14360 96860 -14140 96910
rect -13860 97090 -13640 97140
rect -13860 97020 -13850 97090
rect -13650 97020 -13640 97090
rect -13860 96980 -13640 97020
rect -13860 96910 -13850 96980
rect -13650 96910 -13640 96980
rect -13860 96860 -13640 96910
rect -13360 97090 -13140 97140
rect -13360 97020 -13350 97090
rect -13150 97020 -13140 97090
rect -13360 96980 -13140 97020
rect -13360 96910 -13350 96980
rect -13150 96910 -13140 96980
rect -13360 96860 -13140 96910
rect -12860 97090 -12640 97140
rect -12860 97020 -12850 97090
rect -12650 97020 -12640 97090
rect -12860 96980 -12640 97020
rect -12860 96910 -12850 96980
rect -12650 96910 -12640 96980
rect -12860 96860 -12640 96910
rect -12360 97090 -12140 97140
rect -12360 97020 -12350 97090
rect -12150 97020 -12140 97090
rect -12360 96980 -12140 97020
rect -12360 96910 -12350 96980
rect -12150 96910 -12140 96980
rect -12360 96860 -12140 96910
rect -11860 97090 -11640 97140
rect -11860 97020 -11850 97090
rect -11650 97020 -11640 97090
rect -11860 96980 -11640 97020
rect -11860 96910 -11850 96980
rect -11650 96910 -11640 96980
rect -11860 96860 -11640 96910
rect -11360 97090 -11140 97140
rect -11360 97020 -11350 97090
rect -11150 97020 -11140 97090
rect -11360 96980 -11140 97020
rect -11360 96910 -11350 96980
rect -11150 96910 -11140 96980
rect -11360 96860 -11140 96910
rect -10860 97090 -10640 97140
rect -10860 97020 -10850 97090
rect -10650 97020 -10640 97090
rect -10860 96980 -10640 97020
rect -10860 96910 -10850 96980
rect -10650 96910 -10640 96980
rect -10860 96860 -10640 96910
rect -10360 97090 -10140 97140
rect -10360 97020 -10350 97090
rect -10150 97020 -10140 97090
rect -10360 96980 -10140 97020
rect -10360 96910 -10350 96980
rect -10150 96910 -10140 96980
rect -10360 96860 -10140 96910
rect -9860 97090 -9640 97140
rect -9860 97020 -9850 97090
rect -9650 97020 -9640 97090
rect -9860 96980 -9640 97020
rect -9860 96910 -9850 96980
rect -9650 96910 -9640 96980
rect -9860 96860 -9640 96910
rect -9360 97090 -9140 97140
rect -9360 97020 -9350 97090
rect -9150 97020 -9140 97090
rect -9360 96980 -9140 97020
rect -9360 96910 -9350 96980
rect -9150 96910 -9140 96980
rect -9360 96860 -9140 96910
rect -8860 97090 -8640 97140
rect -8860 97020 -8850 97090
rect -8650 97020 -8640 97090
rect -8860 96980 -8640 97020
rect -8860 96910 -8850 96980
rect -8650 96910 -8640 96980
rect -8860 96860 -8640 96910
rect -8360 97090 -8140 97140
rect -8360 97020 -8350 97090
rect -8150 97020 -8140 97090
rect -8360 96980 -8140 97020
rect -8360 96910 -8350 96980
rect -8150 96910 -8140 96980
rect -8360 96860 -8140 96910
rect -7860 97090 -7640 97140
rect -7860 97020 -7850 97090
rect -7650 97020 -7640 97090
rect -7860 96980 -7640 97020
rect -7860 96910 -7850 96980
rect -7650 96910 -7640 96980
rect -7860 96860 -7640 96910
rect -7360 97090 -7140 97140
rect -7360 97020 -7350 97090
rect -7150 97020 -7140 97090
rect -7360 96980 -7140 97020
rect -7360 96910 -7350 96980
rect -7150 96910 -7140 96980
rect -7360 96860 -7140 96910
rect -6860 97090 -6640 97140
rect -6860 97020 -6850 97090
rect -6650 97020 -6640 97090
rect -6860 96980 -6640 97020
rect -6860 96910 -6850 96980
rect -6650 96910 -6640 96980
rect -6860 96860 -6640 96910
rect -6360 97090 -6140 97140
rect -6360 97020 -6350 97090
rect -6150 97020 -6140 97090
rect -6360 96980 -6140 97020
rect -6360 96910 -6350 96980
rect -6150 96910 -6140 96980
rect -6360 96860 -6140 96910
rect -5860 97090 -5640 97140
rect -5860 97020 -5850 97090
rect -5650 97020 -5640 97090
rect -5860 96980 -5640 97020
rect -5860 96910 -5850 96980
rect -5650 96910 -5640 96980
rect -5860 96860 -5640 96910
rect -5360 97090 -5140 97140
rect -5360 97020 -5350 97090
rect -5150 97020 -5140 97090
rect -5360 96980 -5140 97020
rect -5360 96910 -5350 96980
rect -5150 96910 -5140 96980
rect -5360 96860 -5140 96910
rect -4860 97090 -4640 97140
rect -4860 97020 -4850 97090
rect -4650 97020 -4640 97090
rect -4860 96980 -4640 97020
rect -4860 96910 -4850 96980
rect -4650 96910 -4640 96980
rect -4860 96860 -4640 96910
rect -4360 97090 -4140 97140
rect -4360 97020 -4350 97090
rect -4150 97020 -4140 97090
rect -4360 96980 -4140 97020
rect -4360 96910 -4350 96980
rect -4150 96910 -4140 96980
rect -4360 96860 -4140 96910
rect -3860 97090 -3640 97140
rect -3860 97020 -3850 97090
rect -3650 97020 -3640 97090
rect -3860 96980 -3640 97020
rect -3860 96910 -3850 96980
rect -3650 96910 -3640 96980
rect -3860 96860 -3640 96910
rect -3360 97090 -3140 97140
rect -3360 97020 -3350 97090
rect -3150 97020 -3140 97090
rect -3360 96980 -3140 97020
rect -3360 96910 -3350 96980
rect -3150 96910 -3140 96980
rect -3360 96860 -3140 96910
rect -2860 97090 -2640 97140
rect -2860 97020 -2850 97090
rect -2650 97020 -2640 97090
rect -2860 96980 -2640 97020
rect -2860 96910 -2850 96980
rect -2650 96910 -2640 96980
rect -2860 96860 -2640 96910
rect -2360 97090 -2140 97140
rect -2360 97020 -2350 97090
rect -2150 97020 -2140 97090
rect -2360 96980 -2140 97020
rect -2360 96910 -2350 96980
rect -2150 96910 -2140 96980
rect -2360 96860 -2140 96910
rect -1860 97090 -1640 97140
rect -1860 97020 -1850 97090
rect -1650 97020 -1640 97090
rect -1860 96980 -1640 97020
rect -1860 96910 -1850 96980
rect -1650 96910 -1640 96980
rect -1860 96860 -1640 96910
rect -1360 97090 -1140 97140
rect -1360 97020 -1350 97090
rect -1150 97020 -1140 97090
rect -1360 96980 -1140 97020
rect -1360 96910 -1350 96980
rect -1150 96910 -1140 96980
rect -1360 96860 -1140 96910
rect -860 97090 -640 97140
rect -860 97020 -850 97090
rect -650 97020 -640 97090
rect -860 96980 -640 97020
rect -860 96910 -850 96980
rect -650 96910 -640 96980
rect -860 96860 -640 96910
rect -360 97090 -140 97140
rect -360 97020 -350 97090
rect -150 97020 -140 97090
rect -360 96980 -140 97020
rect -360 96910 -350 96980
rect -150 96910 -140 96980
rect -360 96860 -140 96910
rect 140 97090 360 97140
rect 140 97020 150 97090
rect 350 97020 360 97090
rect 140 96980 360 97020
rect 140 96910 150 96980
rect 350 96910 360 96980
rect 140 96860 360 96910
rect 640 97090 860 97140
rect 640 97020 650 97090
rect 850 97020 860 97090
rect 640 96980 860 97020
rect 640 96910 650 96980
rect 850 96910 860 96980
rect 640 96860 860 96910
rect 1140 97090 1360 97140
rect 1140 97020 1150 97090
rect 1350 97020 1360 97090
rect 1140 96980 1360 97020
rect 1140 96910 1150 96980
rect 1350 96910 1360 96980
rect 1140 96860 1360 96910
rect 1640 97090 1860 97140
rect 1640 97020 1650 97090
rect 1850 97020 1860 97090
rect 1640 96980 1860 97020
rect 1640 96910 1650 96980
rect 1850 96910 1860 96980
rect 1640 96860 1860 96910
rect 2140 97090 2360 97140
rect 2140 97020 2150 97090
rect 2350 97020 2360 97090
rect 2140 96980 2360 97020
rect 2140 96910 2150 96980
rect 2350 96910 2360 96980
rect 2140 96860 2360 96910
rect 2640 97090 2860 97140
rect 2640 97020 2650 97090
rect 2850 97020 2860 97090
rect 2640 96980 2860 97020
rect 2640 96910 2650 96980
rect 2850 96910 2860 96980
rect 2640 96860 2860 96910
rect 3140 97090 3360 97140
rect 3140 97020 3150 97090
rect 3350 97020 3360 97090
rect 3140 96980 3360 97020
rect 3140 96910 3150 96980
rect 3350 96910 3360 96980
rect 3140 96860 3360 96910
rect 3640 97090 3860 97140
rect 3640 97020 3650 97090
rect 3850 97020 3860 97090
rect 3640 96980 3860 97020
rect 3640 96910 3650 96980
rect 3850 96910 3860 96980
rect 3640 96860 3860 96910
rect 4140 97090 4360 97140
rect 4140 97020 4150 97090
rect 4350 97020 4360 97090
rect 4140 96980 4360 97020
rect 4140 96910 4150 96980
rect 4350 96910 4360 96980
rect 4140 96860 4360 96910
rect 4640 97090 4860 97140
rect 4640 97020 4650 97090
rect 4850 97020 4860 97090
rect 4640 96980 4860 97020
rect 4640 96910 4650 96980
rect 4850 96910 4860 96980
rect 4640 96860 4860 96910
rect 5140 97090 5360 97140
rect 5140 97020 5150 97090
rect 5350 97020 5360 97090
rect 5140 96980 5360 97020
rect 5140 96910 5150 96980
rect 5350 96910 5360 96980
rect 5140 96860 5360 96910
rect 5640 97090 5860 97140
rect 5640 97020 5650 97090
rect 5850 97020 5860 97090
rect 5640 96980 5860 97020
rect 5640 96910 5650 96980
rect 5850 96910 5860 96980
rect 5640 96860 5860 96910
rect 6140 97090 6360 97140
rect 6140 97020 6150 97090
rect 6350 97020 6360 97090
rect 6140 96980 6360 97020
rect 6140 96910 6150 96980
rect 6350 96910 6360 96980
rect 6140 96860 6360 96910
rect 6640 97090 6860 97140
rect 6640 97020 6650 97090
rect 6850 97020 6860 97090
rect 6640 96980 6860 97020
rect 6640 96910 6650 96980
rect 6850 96910 6860 96980
rect 6640 96860 6860 96910
rect 7140 97090 7360 97140
rect 7140 97020 7150 97090
rect 7350 97020 7360 97090
rect 7140 96980 7360 97020
rect 7140 96910 7150 96980
rect 7350 96910 7360 96980
rect 7140 96860 7360 96910
rect 7640 97090 7860 97140
rect 7640 97020 7650 97090
rect 7850 97020 7860 97090
rect 7640 96980 7860 97020
rect 7640 96910 7650 96980
rect 7850 96910 7860 96980
rect 7640 96860 7860 96910
rect 8140 97090 8360 97140
rect 8140 97020 8150 97090
rect 8350 97020 8360 97090
rect 8140 96980 8360 97020
rect 8140 96910 8150 96980
rect 8350 96910 8360 96980
rect 8140 96860 8360 96910
rect 8640 97090 8860 97140
rect 8640 97020 8650 97090
rect 8850 97020 8860 97090
rect 8640 96980 8860 97020
rect 8640 96910 8650 96980
rect 8850 96910 8860 96980
rect 8640 96860 8860 96910
rect 9140 97090 9360 97140
rect 9140 97020 9150 97090
rect 9350 97020 9360 97090
rect 9140 96980 9360 97020
rect 9140 96910 9150 96980
rect 9350 96910 9360 96980
rect 9140 96860 9360 96910
rect 9640 97090 9860 97140
rect 9640 97020 9650 97090
rect 9850 97020 9860 97090
rect 9640 96980 9860 97020
rect 9640 96910 9650 96980
rect 9850 96910 9860 96980
rect 9640 96860 9860 96910
rect 10140 97090 10360 97140
rect 10140 97020 10150 97090
rect 10350 97020 10360 97090
rect 10140 96980 10360 97020
rect 10140 96910 10150 96980
rect 10350 96910 10360 96980
rect 10140 96860 10360 96910
rect 10640 97090 10860 97140
rect 10640 97020 10650 97090
rect 10850 97020 10860 97090
rect 10640 96980 10860 97020
rect 10640 96910 10650 96980
rect 10850 96910 10860 96980
rect 10640 96860 10860 96910
rect 11140 97090 11360 97140
rect 11140 97020 11150 97090
rect 11350 97020 11360 97090
rect 11140 96980 11360 97020
rect 11140 96910 11150 96980
rect 11350 96910 11360 96980
rect 11140 96860 11360 96910
rect 11640 97090 11860 97140
rect 11640 97020 11650 97090
rect 11850 97020 11860 97090
rect 11640 96980 11860 97020
rect 11640 96910 11650 96980
rect 11850 96910 11860 96980
rect 11640 96860 11860 96910
rect 12140 97090 12360 97140
rect 12140 97020 12150 97090
rect 12350 97020 12360 97090
rect 12140 96980 12360 97020
rect 12140 96910 12150 96980
rect 12350 96910 12360 96980
rect 12140 96860 12360 96910
rect 12640 97090 12860 97140
rect 12640 97020 12650 97090
rect 12850 97020 12860 97090
rect 12640 96980 12860 97020
rect 12640 96910 12650 96980
rect 12850 96910 12860 96980
rect 12640 96860 12860 96910
rect 13140 97090 13360 97140
rect 13140 97020 13150 97090
rect 13350 97020 13360 97090
rect 13140 96980 13360 97020
rect 13140 96910 13150 96980
rect 13350 96910 13360 96980
rect 13140 96860 13360 96910
rect 13640 97090 13860 97140
rect 13640 97020 13650 97090
rect 13850 97020 13860 97090
rect 13640 96980 13860 97020
rect 13640 96910 13650 96980
rect 13850 96910 13860 96980
rect 13640 96860 13860 96910
rect 14140 97090 14360 97140
rect 14140 97020 14150 97090
rect 14350 97020 14360 97090
rect 14140 96980 14360 97020
rect 14140 96910 14150 96980
rect 14350 96910 14360 96980
rect 14140 96860 14360 96910
rect 14640 97090 14860 97140
rect 14640 97020 14650 97090
rect 14850 97020 14860 97090
rect 14640 96980 14860 97020
rect 14640 96910 14650 96980
rect 14850 96910 14860 96980
rect 14640 96860 14860 96910
rect 15140 97090 15360 97140
rect 15140 97020 15150 97090
rect 15350 97020 15360 97090
rect 15140 96980 15360 97020
rect 15140 96910 15150 96980
rect 15350 96910 15360 96980
rect 15140 96860 15360 96910
rect 15640 97090 15860 97140
rect 15640 97020 15650 97090
rect 15850 97020 15860 97090
rect 15640 96980 15860 97020
rect 15640 96910 15650 96980
rect 15850 96910 15860 96980
rect 15640 96860 15860 96910
rect 16140 97090 16360 97140
rect 16140 97020 16150 97090
rect 16350 97020 16360 97090
rect 16140 96980 16360 97020
rect 16140 96910 16150 96980
rect 16350 96910 16360 96980
rect 16140 96860 16360 96910
rect 16640 97090 16860 97140
rect 16640 97020 16650 97090
rect 16850 97020 16860 97090
rect 16640 96980 16860 97020
rect 16640 96910 16650 96980
rect 16850 96910 16860 96980
rect 16640 96860 16860 96910
rect 17140 97090 17360 97140
rect 17140 97020 17150 97090
rect 17350 97020 17360 97090
rect 17140 96980 17360 97020
rect 17140 96910 17150 96980
rect 17350 96910 17360 96980
rect 17140 96860 17360 96910
rect 17640 97090 17860 97140
rect 17640 97020 17650 97090
rect 17850 97020 17860 97090
rect 17640 96980 17860 97020
rect 17640 96910 17650 96980
rect 17850 96910 17860 96980
rect 17640 96860 17860 96910
rect 18140 97090 18360 97140
rect 18140 97020 18150 97090
rect 18350 97020 18360 97090
rect 18140 96980 18360 97020
rect 18140 96910 18150 96980
rect 18350 96910 18360 96980
rect 18140 96860 18360 96910
rect 18640 97090 18860 97140
rect 18640 97020 18650 97090
rect 18850 97020 18860 97090
rect 18640 96980 18860 97020
rect 18640 96910 18650 96980
rect 18850 96910 18860 96980
rect 18640 96860 18860 96910
rect 19140 97090 19360 97140
rect 19140 97020 19150 97090
rect 19350 97020 19360 97090
rect 19140 96980 19360 97020
rect 19140 96910 19150 96980
rect 19350 96910 19360 96980
rect 19140 96860 19360 96910
rect 19640 97090 19860 97140
rect 19640 97020 19650 97090
rect 19850 97020 19860 97090
rect 19640 96980 19860 97020
rect 19640 96910 19650 96980
rect 19850 96910 19860 96980
rect 19640 96860 19860 96910
rect -16000 96850 20000 96860
rect -16000 96650 -15980 96850
rect -15910 96650 -15590 96850
rect -15520 96650 -15480 96850
rect -15410 96650 -15090 96850
rect -15020 96650 -14980 96850
rect -14910 96650 -14590 96850
rect -14520 96650 -14480 96850
rect -14410 96650 -14090 96850
rect -14020 96650 -13980 96850
rect -13910 96650 -13590 96850
rect -13520 96650 -13480 96850
rect -13410 96650 -13090 96850
rect -13020 96650 -12980 96850
rect -12910 96650 -12590 96850
rect -12520 96650 -12480 96850
rect -12410 96650 -12090 96850
rect -12020 96650 -11980 96850
rect -11910 96650 -11590 96850
rect -11520 96650 -11480 96850
rect -11410 96650 -11090 96850
rect -11020 96650 -10980 96850
rect -10910 96650 -10590 96850
rect -10520 96650 -10480 96850
rect -10410 96650 -10090 96850
rect -10020 96650 -9980 96850
rect -9910 96650 -9590 96850
rect -9520 96650 -9480 96850
rect -9410 96650 -9090 96850
rect -9020 96650 -8980 96850
rect -8910 96650 -8590 96850
rect -8520 96650 -8480 96850
rect -8410 96650 -8090 96850
rect -8020 96650 -7980 96850
rect -7910 96650 -7590 96850
rect -7520 96650 -7480 96850
rect -7410 96650 -7090 96850
rect -7020 96650 -6980 96850
rect -6910 96650 -6590 96850
rect -6520 96650 -6480 96850
rect -6410 96650 -6090 96850
rect -6020 96650 -5980 96850
rect -5910 96650 -5590 96850
rect -5520 96650 -5480 96850
rect -5410 96650 -5090 96850
rect -5020 96650 -4980 96850
rect -4910 96650 -4590 96850
rect -4520 96650 -4480 96850
rect -4410 96650 -4090 96850
rect -4020 96650 -3980 96850
rect -3910 96650 -3590 96850
rect -3520 96650 -3480 96850
rect -3410 96650 -3090 96850
rect -3020 96650 -2980 96850
rect -2910 96650 -2590 96850
rect -2520 96650 -2480 96850
rect -2410 96650 -2090 96850
rect -2020 96650 -1980 96850
rect -1910 96650 -1590 96850
rect -1520 96650 -1480 96850
rect -1410 96650 -1090 96850
rect -1020 96650 -980 96850
rect -910 96650 -590 96850
rect -520 96650 -480 96850
rect -410 96650 -90 96850
rect -20 96650 20 96850
rect 90 96650 410 96850
rect 480 96650 520 96850
rect 590 96650 910 96850
rect 980 96650 1020 96850
rect 1090 96650 1410 96850
rect 1480 96650 1520 96850
rect 1590 96650 1910 96850
rect 1980 96650 2020 96850
rect 2090 96650 2410 96850
rect 2480 96650 2520 96850
rect 2590 96650 2910 96850
rect 2980 96650 3020 96850
rect 3090 96650 3410 96850
rect 3480 96650 3520 96850
rect 3590 96650 3910 96850
rect 3980 96650 4020 96850
rect 4090 96650 4410 96850
rect 4480 96650 4520 96850
rect 4590 96650 4910 96850
rect 4980 96650 5020 96850
rect 5090 96650 5410 96850
rect 5480 96650 5520 96850
rect 5590 96650 5910 96850
rect 5980 96650 6020 96850
rect 6090 96650 6410 96850
rect 6480 96650 6520 96850
rect 6590 96650 6910 96850
rect 6980 96650 7020 96850
rect 7090 96650 7410 96850
rect 7480 96650 7520 96850
rect 7590 96650 7910 96850
rect 7980 96650 8020 96850
rect 8090 96650 8410 96850
rect 8480 96650 8520 96850
rect 8590 96650 8910 96850
rect 8980 96650 9020 96850
rect 9090 96650 9410 96850
rect 9480 96650 9520 96850
rect 9590 96650 9910 96850
rect 9980 96650 10020 96850
rect 10090 96650 10410 96850
rect 10480 96650 10520 96850
rect 10590 96650 10910 96850
rect 10980 96650 11020 96850
rect 11090 96650 11410 96850
rect 11480 96650 11520 96850
rect 11590 96650 11910 96850
rect 11980 96650 12020 96850
rect 12090 96650 12410 96850
rect 12480 96650 12520 96850
rect 12590 96650 12910 96850
rect 12980 96650 13020 96850
rect 13090 96650 13410 96850
rect 13480 96650 13520 96850
rect 13590 96650 13910 96850
rect 13980 96650 14020 96850
rect 14090 96650 14410 96850
rect 14480 96650 14520 96850
rect 14590 96650 14910 96850
rect 14980 96650 15020 96850
rect 15090 96650 15410 96850
rect 15480 96650 15520 96850
rect 15590 96650 15910 96850
rect 15980 96650 16020 96850
rect 16090 96650 16410 96850
rect 16480 96650 16520 96850
rect 16590 96650 16910 96850
rect 16980 96650 17020 96850
rect 17090 96650 17410 96850
rect 17480 96650 17520 96850
rect 17590 96650 17910 96850
rect 17980 96650 18020 96850
rect 18090 96650 18410 96850
rect 18480 96650 18520 96850
rect 18590 96650 18910 96850
rect 18980 96650 19020 96850
rect 19090 96650 19410 96850
rect 19480 96650 19520 96850
rect 19590 96650 19910 96850
rect 19980 96650 20000 96850
rect -16000 96640 20000 96650
rect -15860 96590 -15640 96640
rect -15860 96520 -15850 96590
rect -15650 96520 -15640 96590
rect -15860 96480 -15640 96520
rect -15860 96410 -15850 96480
rect -15650 96410 -15640 96480
rect -15860 96360 -15640 96410
rect -15360 96590 -15140 96640
rect -15360 96520 -15350 96590
rect -15150 96520 -15140 96590
rect -15360 96480 -15140 96520
rect -15360 96410 -15350 96480
rect -15150 96410 -15140 96480
rect -15360 96360 -15140 96410
rect -14860 96590 -14640 96640
rect -14860 96520 -14850 96590
rect -14650 96520 -14640 96590
rect -14860 96480 -14640 96520
rect -14860 96410 -14850 96480
rect -14650 96410 -14640 96480
rect -14860 96360 -14640 96410
rect -14360 96590 -14140 96640
rect -14360 96520 -14350 96590
rect -14150 96520 -14140 96590
rect -14360 96480 -14140 96520
rect -14360 96410 -14350 96480
rect -14150 96410 -14140 96480
rect -14360 96360 -14140 96410
rect -13860 96590 -13640 96640
rect -13860 96520 -13850 96590
rect -13650 96520 -13640 96590
rect -13860 96480 -13640 96520
rect -13860 96410 -13850 96480
rect -13650 96410 -13640 96480
rect -13860 96360 -13640 96410
rect -13360 96590 -13140 96640
rect -13360 96520 -13350 96590
rect -13150 96520 -13140 96590
rect -13360 96480 -13140 96520
rect -13360 96410 -13350 96480
rect -13150 96410 -13140 96480
rect -13360 96360 -13140 96410
rect -12860 96590 -12640 96640
rect -12860 96520 -12850 96590
rect -12650 96520 -12640 96590
rect -12860 96480 -12640 96520
rect -12860 96410 -12850 96480
rect -12650 96410 -12640 96480
rect -12860 96360 -12640 96410
rect -12360 96590 -12140 96640
rect -12360 96520 -12350 96590
rect -12150 96520 -12140 96590
rect -12360 96480 -12140 96520
rect -12360 96410 -12350 96480
rect -12150 96410 -12140 96480
rect -12360 96360 -12140 96410
rect -11860 96590 -11640 96640
rect -11860 96520 -11850 96590
rect -11650 96520 -11640 96590
rect -11860 96480 -11640 96520
rect -11860 96410 -11850 96480
rect -11650 96410 -11640 96480
rect -11860 96360 -11640 96410
rect -11360 96590 -11140 96640
rect -11360 96520 -11350 96590
rect -11150 96520 -11140 96590
rect -11360 96480 -11140 96520
rect -11360 96410 -11350 96480
rect -11150 96410 -11140 96480
rect -11360 96360 -11140 96410
rect -10860 96590 -10640 96640
rect -10860 96520 -10850 96590
rect -10650 96520 -10640 96590
rect -10860 96480 -10640 96520
rect -10860 96410 -10850 96480
rect -10650 96410 -10640 96480
rect -10860 96360 -10640 96410
rect -10360 96590 -10140 96640
rect -10360 96520 -10350 96590
rect -10150 96520 -10140 96590
rect -10360 96480 -10140 96520
rect -10360 96410 -10350 96480
rect -10150 96410 -10140 96480
rect -10360 96360 -10140 96410
rect -9860 96590 -9640 96640
rect -9860 96520 -9850 96590
rect -9650 96520 -9640 96590
rect -9860 96480 -9640 96520
rect -9860 96410 -9850 96480
rect -9650 96410 -9640 96480
rect -9860 96360 -9640 96410
rect -9360 96590 -9140 96640
rect -9360 96520 -9350 96590
rect -9150 96520 -9140 96590
rect -9360 96480 -9140 96520
rect -9360 96410 -9350 96480
rect -9150 96410 -9140 96480
rect -9360 96360 -9140 96410
rect -8860 96590 -8640 96640
rect -8860 96520 -8850 96590
rect -8650 96520 -8640 96590
rect -8860 96480 -8640 96520
rect -8860 96410 -8850 96480
rect -8650 96410 -8640 96480
rect -8860 96360 -8640 96410
rect -8360 96590 -8140 96640
rect -8360 96520 -8350 96590
rect -8150 96520 -8140 96590
rect -8360 96480 -8140 96520
rect -8360 96410 -8350 96480
rect -8150 96410 -8140 96480
rect -8360 96360 -8140 96410
rect -7860 96590 -7640 96640
rect -7860 96520 -7850 96590
rect -7650 96520 -7640 96590
rect -7860 96480 -7640 96520
rect -7860 96410 -7850 96480
rect -7650 96410 -7640 96480
rect -7860 96360 -7640 96410
rect -7360 96590 -7140 96640
rect -7360 96520 -7350 96590
rect -7150 96520 -7140 96590
rect -7360 96480 -7140 96520
rect -7360 96410 -7350 96480
rect -7150 96410 -7140 96480
rect -7360 96360 -7140 96410
rect -6860 96590 -6640 96640
rect -6860 96520 -6850 96590
rect -6650 96520 -6640 96590
rect -6860 96480 -6640 96520
rect -6860 96410 -6850 96480
rect -6650 96410 -6640 96480
rect -6860 96360 -6640 96410
rect -6360 96590 -6140 96640
rect -6360 96520 -6350 96590
rect -6150 96520 -6140 96590
rect -6360 96480 -6140 96520
rect -6360 96410 -6350 96480
rect -6150 96410 -6140 96480
rect -6360 96360 -6140 96410
rect -5860 96590 -5640 96640
rect -5860 96520 -5850 96590
rect -5650 96520 -5640 96590
rect -5860 96480 -5640 96520
rect -5860 96410 -5850 96480
rect -5650 96410 -5640 96480
rect -5860 96360 -5640 96410
rect -5360 96590 -5140 96640
rect -5360 96520 -5350 96590
rect -5150 96520 -5140 96590
rect -5360 96480 -5140 96520
rect -5360 96410 -5350 96480
rect -5150 96410 -5140 96480
rect -5360 96360 -5140 96410
rect -4860 96590 -4640 96640
rect -4860 96520 -4850 96590
rect -4650 96520 -4640 96590
rect -4860 96480 -4640 96520
rect -4860 96410 -4850 96480
rect -4650 96410 -4640 96480
rect -4860 96360 -4640 96410
rect -4360 96590 -4140 96640
rect -4360 96520 -4350 96590
rect -4150 96520 -4140 96590
rect -4360 96480 -4140 96520
rect -4360 96410 -4350 96480
rect -4150 96410 -4140 96480
rect -4360 96360 -4140 96410
rect -3860 96590 -3640 96640
rect -3860 96520 -3850 96590
rect -3650 96520 -3640 96590
rect -3860 96480 -3640 96520
rect -3860 96410 -3850 96480
rect -3650 96410 -3640 96480
rect -3860 96360 -3640 96410
rect -3360 96590 -3140 96640
rect -3360 96520 -3350 96590
rect -3150 96520 -3140 96590
rect -3360 96480 -3140 96520
rect -3360 96410 -3350 96480
rect -3150 96410 -3140 96480
rect -3360 96360 -3140 96410
rect -2860 96590 -2640 96640
rect -2860 96520 -2850 96590
rect -2650 96520 -2640 96590
rect -2860 96480 -2640 96520
rect -2860 96410 -2850 96480
rect -2650 96410 -2640 96480
rect -2860 96360 -2640 96410
rect -2360 96590 -2140 96640
rect -2360 96520 -2350 96590
rect -2150 96520 -2140 96590
rect -2360 96480 -2140 96520
rect -2360 96410 -2350 96480
rect -2150 96410 -2140 96480
rect -2360 96360 -2140 96410
rect -1860 96590 -1640 96640
rect -1860 96520 -1850 96590
rect -1650 96520 -1640 96590
rect -1860 96480 -1640 96520
rect -1860 96410 -1850 96480
rect -1650 96410 -1640 96480
rect -1860 96360 -1640 96410
rect -1360 96590 -1140 96640
rect -1360 96520 -1350 96590
rect -1150 96520 -1140 96590
rect -1360 96480 -1140 96520
rect -1360 96410 -1350 96480
rect -1150 96410 -1140 96480
rect -1360 96360 -1140 96410
rect -860 96590 -640 96640
rect -860 96520 -850 96590
rect -650 96520 -640 96590
rect -860 96480 -640 96520
rect -860 96410 -850 96480
rect -650 96410 -640 96480
rect -860 96360 -640 96410
rect -360 96590 -140 96640
rect -360 96520 -350 96590
rect -150 96520 -140 96590
rect -360 96480 -140 96520
rect -360 96410 -350 96480
rect -150 96410 -140 96480
rect -360 96360 -140 96410
rect 140 96590 360 96640
rect 140 96520 150 96590
rect 350 96520 360 96590
rect 140 96480 360 96520
rect 140 96410 150 96480
rect 350 96410 360 96480
rect 140 96360 360 96410
rect 640 96590 860 96640
rect 640 96520 650 96590
rect 850 96520 860 96590
rect 640 96480 860 96520
rect 640 96410 650 96480
rect 850 96410 860 96480
rect 640 96360 860 96410
rect 1140 96590 1360 96640
rect 1140 96520 1150 96590
rect 1350 96520 1360 96590
rect 1140 96480 1360 96520
rect 1140 96410 1150 96480
rect 1350 96410 1360 96480
rect 1140 96360 1360 96410
rect 1640 96590 1860 96640
rect 1640 96520 1650 96590
rect 1850 96520 1860 96590
rect 1640 96480 1860 96520
rect 1640 96410 1650 96480
rect 1850 96410 1860 96480
rect 1640 96360 1860 96410
rect 2140 96590 2360 96640
rect 2140 96520 2150 96590
rect 2350 96520 2360 96590
rect 2140 96480 2360 96520
rect 2140 96410 2150 96480
rect 2350 96410 2360 96480
rect 2140 96360 2360 96410
rect 2640 96590 2860 96640
rect 2640 96520 2650 96590
rect 2850 96520 2860 96590
rect 2640 96480 2860 96520
rect 2640 96410 2650 96480
rect 2850 96410 2860 96480
rect 2640 96360 2860 96410
rect 3140 96590 3360 96640
rect 3140 96520 3150 96590
rect 3350 96520 3360 96590
rect 3140 96480 3360 96520
rect 3140 96410 3150 96480
rect 3350 96410 3360 96480
rect 3140 96360 3360 96410
rect 3640 96590 3860 96640
rect 3640 96520 3650 96590
rect 3850 96520 3860 96590
rect 3640 96480 3860 96520
rect 3640 96410 3650 96480
rect 3850 96410 3860 96480
rect 3640 96360 3860 96410
rect 4140 96590 4360 96640
rect 4140 96520 4150 96590
rect 4350 96520 4360 96590
rect 4140 96480 4360 96520
rect 4140 96410 4150 96480
rect 4350 96410 4360 96480
rect 4140 96360 4360 96410
rect 4640 96590 4860 96640
rect 4640 96520 4650 96590
rect 4850 96520 4860 96590
rect 4640 96480 4860 96520
rect 4640 96410 4650 96480
rect 4850 96410 4860 96480
rect 4640 96360 4860 96410
rect 5140 96590 5360 96640
rect 5140 96520 5150 96590
rect 5350 96520 5360 96590
rect 5140 96480 5360 96520
rect 5140 96410 5150 96480
rect 5350 96410 5360 96480
rect 5140 96360 5360 96410
rect 5640 96590 5860 96640
rect 5640 96520 5650 96590
rect 5850 96520 5860 96590
rect 5640 96480 5860 96520
rect 5640 96410 5650 96480
rect 5850 96410 5860 96480
rect 5640 96360 5860 96410
rect 6140 96590 6360 96640
rect 6140 96520 6150 96590
rect 6350 96520 6360 96590
rect 6140 96480 6360 96520
rect 6140 96410 6150 96480
rect 6350 96410 6360 96480
rect 6140 96360 6360 96410
rect 6640 96590 6860 96640
rect 6640 96520 6650 96590
rect 6850 96520 6860 96590
rect 6640 96480 6860 96520
rect 6640 96410 6650 96480
rect 6850 96410 6860 96480
rect 6640 96360 6860 96410
rect 7140 96590 7360 96640
rect 7140 96520 7150 96590
rect 7350 96520 7360 96590
rect 7140 96480 7360 96520
rect 7140 96410 7150 96480
rect 7350 96410 7360 96480
rect 7140 96360 7360 96410
rect 7640 96590 7860 96640
rect 7640 96520 7650 96590
rect 7850 96520 7860 96590
rect 7640 96480 7860 96520
rect 7640 96410 7650 96480
rect 7850 96410 7860 96480
rect 7640 96360 7860 96410
rect 8140 96590 8360 96640
rect 8140 96520 8150 96590
rect 8350 96520 8360 96590
rect 8140 96480 8360 96520
rect 8140 96410 8150 96480
rect 8350 96410 8360 96480
rect 8140 96360 8360 96410
rect 8640 96590 8860 96640
rect 8640 96520 8650 96590
rect 8850 96520 8860 96590
rect 8640 96480 8860 96520
rect 8640 96410 8650 96480
rect 8850 96410 8860 96480
rect 8640 96360 8860 96410
rect 9140 96590 9360 96640
rect 9140 96520 9150 96590
rect 9350 96520 9360 96590
rect 9140 96480 9360 96520
rect 9140 96410 9150 96480
rect 9350 96410 9360 96480
rect 9140 96360 9360 96410
rect 9640 96590 9860 96640
rect 9640 96520 9650 96590
rect 9850 96520 9860 96590
rect 9640 96480 9860 96520
rect 9640 96410 9650 96480
rect 9850 96410 9860 96480
rect 9640 96360 9860 96410
rect 10140 96590 10360 96640
rect 10140 96520 10150 96590
rect 10350 96520 10360 96590
rect 10140 96480 10360 96520
rect 10140 96410 10150 96480
rect 10350 96410 10360 96480
rect 10140 96360 10360 96410
rect 10640 96590 10860 96640
rect 10640 96520 10650 96590
rect 10850 96520 10860 96590
rect 10640 96480 10860 96520
rect 10640 96410 10650 96480
rect 10850 96410 10860 96480
rect 10640 96360 10860 96410
rect 11140 96590 11360 96640
rect 11140 96520 11150 96590
rect 11350 96520 11360 96590
rect 11140 96480 11360 96520
rect 11140 96410 11150 96480
rect 11350 96410 11360 96480
rect 11140 96360 11360 96410
rect 11640 96590 11860 96640
rect 11640 96520 11650 96590
rect 11850 96520 11860 96590
rect 11640 96480 11860 96520
rect 11640 96410 11650 96480
rect 11850 96410 11860 96480
rect 11640 96360 11860 96410
rect 12140 96590 12360 96640
rect 12140 96520 12150 96590
rect 12350 96520 12360 96590
rect 12140 96480 12360 96520
rect 12140 96410 12150 96480
rect 12350 96410 12360 96480
rect 12140 96360 12360 96410
rect 12640 96590 12860 96640
rect 12640 96520 12650 96590
rect 12850 96520 12860 96590
rect 12640 96480 12860 96520
rect 12640 96410 12650 96480
rect 12850 96410 12860 96480
rect 12640 96360 12860 96410
rect 13140 96590 13360 96640
rect 13140 96520 13150 96590
rect 13350 96520 13360 96590
rect 13140 96480 13360 96520
rect 13140 96410 13150 96480
rect 13350 96410 13360 96480
rect 13140 96360 13360 96410
rect 13640 96590 13860 96640
rect 13640 96520 13650 96590
rect 13850 96520 13860 96590
rect 13640 96480 13860 96520
rect 13640 96410 13650 96480
rect 13850 96410 13860 96480
rect 13640 96360 13860 96410
rect 14140 96590 14360 96640
rect 14140 96520 14150 96590
rect 14350 96520 14360 96590
rect 14140 96480 14360 96520
rect 14140 96410 14150 96480
rect 14350 96410 14360 96480
rect 14140 96360 14360 96410
rect 14640 96590 14860 96640
rect 14640 96520 14650 96590
rect 14850 96520 14860 96590
rect 14640 96480 14860 96520
rect 14640 96410 14650 96480
rect 14850 96410 14860 96480
rect 14640 96360 14860 96410
rect 15140 96590 15360 96640
rect 15140 96520 15150 96590
rect 15350 96520 15360 96590
rect 15140 96480 15360 96520
rect 15140 96410 15150 96480
rect 15350 96410 15360 96480
rect 15140 96360 15360 96410
rect 15640 96590 15860 96640
rect 15640 96520 15650 96590
rect 15850 96520 15860 96590
rect 15640 96480 15860 96520
rect 15640 96410 15650 96480
rect 15850 96410 15860 96480
rect 15640 96360 15860 96410
rect 16140 96590 16360 96640
rect 16140 96520 16150 96590
rect 16350 96520 16360 96590
rect 16140 96480 16360 96520
rect 16140 96410 16150 96480
rect 16350 96410 16360 96480
rect 16140 96360 16360 96410
rect 16640 96590 16860 96640
rect 16640 96520 16650 96590
rect 16850 96520 16860 96590
rect 16640 96480 16860 96520
rect 16640 96410 16650 96480
rect 16850 96410 16860 96480
rect 16640 96360 16860 96410
rect 17140 96590 17360 96640
rect 17140 96520 17150 96590
rect 17350 96520 17360 96590
rect 17140 96480 17360 96520
rect 17140 96410 17150 96480
rect 17350 96410 17360 96480
rect 17140 96360 17360 96410
rect 17640 96590 17860 96640
rect 17640 96520 17650 96590
rect 17850 96520 17860 96590
rect 17640 96480 17860 96520
rect 17640 96410 17650 96480
rect 17850 96410 17860 96480
rect 17640 96360 17860 96410
rect 18140 96590 18360 96640
rect 18140 96520 18150 96590
rect 18350 96520 18360 96590
rect 18140 96480 18360 96520
rect 18140 96410 18150 96480
rect 18350 96410 18360 96480
rect 18140 96360 18360 96410
rect 18640 96590 18860 96640
rect 18640 96520 18650 96590
rect 18850 96520 18860 96590
rect 18640 96480 18860 96520
rect 18640 96410 18650 96480
rect 18850 96410 18860 96480
rect 18640 96360 18860 96410
rect 19140 96590 19360 96640
rect 19140 96520 19150 96590
rect 19350 96520 19360 96590
rect 19140 96480 19360 96520
rect 19140 96410 19150 96480
rect 19350 96410 19360 96480
rect 19140 96360 19360 96410
rect 19640 96590 19860 96640
rect 19640 96520 19650 96590
rect 19850 96520 19860 96590
rect 19640 96480 19860 96520
rect 19640 96410 19650 96480
rect 19850 96410 19860 96480
rect 19640 96360 19860 96410
rect -16000 96350 20000 96360
rect -16000 96150 -15980 96350
rect -15910 96150 -15590 96350
rect -15520 96150 -15480 96350
rect -15410 96150 -15090 96350
rect -15020 96150 -14980 96350
rect -14910 96150 -14590 96350
rect -14520 96150 -14480 96350
rect -14410 96150 -14090 96350
rect -14020 96150 -13980 96350
rect -13910 96150 -13590 96350
rect -13520 96150 -13480 96350
rect -13410 96150 -13090 96350
rect -13020 96150 -12980 96350
rect -12910 96150 -12590 96350
rect -12520 96150 -12480 96350
rect -12410 96150 -12090 96350
rect -12020 96150 -11980 96350
rect -11910 96150 -11590 96350
rect -11520 96150 -11480 96350
rect -11410 96150 -11090 96350
rect -11020 96150 -10980 96350
rect -10910 96150 -10590 96350
rect -10520 96150 -10480 96350
rect -10410 96150 -10090 96350
rect -10020 96150 -9980 96350
rect -9910 96150 -9590 96350
rect -9520 96150 -9480 96350
rect -9410 96150 -9090 96350
rect -9020 96150 -8980 96350
rect -8910 96150 -8590 96350
rect -8520 96150 -8480 96350
rect -8410 96150 -8090 96350
rect -8020 96150 -7980 96350
rect -7910 96150 -7590 96350
rect -7520 96150 -7480 96350
rect -7410 96150 -7090 96350
rect -7020 96150 -6980 96350
rect -6910 96150 -6590 96350
rect -6520 96150 -6480 96350
rect -6410 96150 -6090 96350
rect -6020 96150 -5980 96350
rect -5910 96150 -5590 96350
rect -5520 96150 -5480 96350
rect -5410 96150 -5090 96350
rect -5020 96150 -4980 96350
rect -4910 96150 -4590 96350
rect -4520 96150 -4480 96350
rect -4410 96150 -4090 96350
rect -4020 96150 -3980 96350
rect -3910 96150 -3590 96350
rect -3520 96150 -3480 96350
rect -3410 96150 -3090 96350
rect -3020 96150 -2980 96350
rect -2910 96150 -2590 96350
rect -2520 96150 -2480 96350
rect -2410 96150 -2090 96350
rect -2020 96150 -1980 96350
rect -1910 96150 -1590 96350
rect -1520 96150 -1480 96350
rect -1410 96150 -1090 96350
rect -1020 96150 -980 96350
rect -910 96150 -590 96350
rect -520 96150 -480 96350
rect -410 96150 -90 96350
rect -20 96150 20 96350
rect 90 96150 410 96350
rect 480 96150 520 96350
rect 590 96150 910 96350
rect 980 96150 1020 96350
rect 1090 96150 1410 96350
rect 1480 96150 1520 96350
rect 1590 96150 1910 96350
rect 1980 96150 2020 96350
rect 2090 96150 2410 96350
rect 2480 96150 2520 96350
rect 2590 96150 2910 96350
rect 2980 96150 3020 96350
rect 3090 96150 3410 96350
rect 3480 96150 3520 96350
rect 3590 96150 3910 96350
rect 3980 96150 4020 96350
rect 4090 96150 4410 96350
rect 4480 96150 4520 96350
rect 4590 96150 4910 96350
rect 4980 96150 5020 96350
rect 5090 96150 5410 96350
rect 5480 96150 5520 96350
rect 5590 96150 5910 96350
rect 5980 96150 6020 96350
rect 6090 96150 6410 96350
rect 6480 96150 6520 96350
rect 6590 96150 6910 96350
rect 6980 96150 7020 96350
rect 7090 96150 7410 96350
rect 7480 96150 7520 96350
rect 7590 96150 7910 96350
rect 7980 96150 8020 96350
rect 8090 96150 8410 96350
rect 8480 96150 8520 96350
rect 8590 96150 8910 96350
rect 8980 96150 9020 96350
rect 9090 96150 9410 96350
rect 9480 96150 9520 96350
rect 9590 96150 9910 96350
rect 9980 96150 10020 96350
rect 10090 96150 10410 96350
rect 10480 96150 10520 96350
rect 10590 96150 10910 96350
rect 10980 96150 11020 96350
rect 11090 96150 11410 96350
rect 11480 96150 11520 96350
rect 11590 96150 11910 96350
rect 11980 96150 12020 96350
rect 12090 96150 12410 96350
rect 12480 96150 12520 96350
rect 12590 96150 12910 96350
rect 12980 96150 13020 96350
rect 13090 96150 13410 96350
rect 13480 96150 13520 96350
rect 13590 96150 13910 96350
rect 13980 96150 14020 96350
rect 14090 96150 14410 96350
rect 14480 96150 14520 96350
rect 14590 96150 14910 96350
rect 14980 96150 15020 96350
rect 15090 96150 15410 96350
rect 15480 96150 15520 96350
rect 15590 96150 15910 96350
rect 15980 96150 16020 96350
rect 16090 96150 16410 96350
rect 16480 96150 16520 96350
rect 16590 96150 16910 96350
rect 16980 96150 17020 96350
rect 17090 96150 17410 96350
rect 17480 96150 17520 96350
rect 17590 96150 17910 96350
rect 17980 96150 18020 96350
rect 18090 96150 18410 96350
rect 18480 96150 18520 96350
rect 18590 96150 18910 96350
rect 18980 96150 19020 96350
rect 19090 96150 19410 96350
rect 19480 96150 19520 96350
rect 19590 96150 19910 96350
rect 19980 96150 20000 96350
rect -16000 96140 20000 96150
rect -15860 96090 -15640 96140
rect -15860 96020 -15850 96090
rect -15650 96020 -15640 96090
rect -15860 95980 -15640 96020
rect -15860 95910 -15850 95980
rect -15650 95910 -15640 95980
rect -15860 95860 -15640 95910
rect -15360 96090 -15140 96140
rect -15360 96020 -15350 96090
rect -15150 96020 -15140 96090
rect -15360 95980 -15140 96020
rect -15360 95910 -15350 95980
rect -15150 95910 -15140 95980
rect -15360 95860 -15140 95910
rect -14860 96090 -14640 96140
rect -14860 96020 -14850 96090
rect -14650 96020 -14640 96090
rect -14860 95980 -14640 96020
rect -14860 95910 -14850 95980
rect -14650 95910 -14640 95980
rect -14860 95860 -14640 95910
rect -14360 96090 -14140 96140
rect -14360 96020 -14350 96090
rect -14150 96020 -14140 96090
rect -14360 95980 -14140 96020
rect -14360 95910 -14350 95980
rect -14150 95910 -14140 95980
rect -14360 95860 -14140 95910
rect -13860 96090 -13640 96140
rect -13860 96020 -13850 96090
rect -13650 96020 -13640 96090
rect -13860 95980 -13640 96020
rect -13860 95910 -13850 95980
rect -13650 95910 -13640 95980
rect -13860 95860 -13640 95910
rect -13360 96090 -13140 96140
rect -13360 96020 -13350 96090
rect -13150 96020 -13140 96090
rect -13360 95980 -13140 96020
rect -13360 95910 -13350 95980
rect -13150 95910 -13140 95980
rect -13360 95860 -13140 95910
rect -12860 96090 -12640 96140
rect -12860 96020 -12850 96090
rect -12650 96020 -12640 96090
rect -12860 95980 -12640 96020
rect -12860 95910 -12850 95980
rect -12650 95910 -12640 95980
rect -12860 95860 -12640 95910
rect -12360 96090 -12140 96140
rect -12360 96020 -12350 96090
rect -12150 96020 -12140 96090
rect -12360 95980 -12140 96020
rect -12360 95910 -12350 95980
rect -12150 95910 -12140 95980
rect -12360 95860 -12140 95910
rect -11860 96090 -11640 96140
rect -11860 96020 -11850 96090
rect -11650 96020 -11640 96090
rect -11860 95980 -11640 96020
rect -11860 95910 -11850 95980
rect -11650 95910 -11640 95980
rect -11860 95860 -11640 95910
rect -11360 96090 -11140 96140
rect -11360 96020 -11350 96090
rect -11150 96020 -11140 96090
rect -11360 95980 -11140 96020
rect -11360 95910 -11350 95980
rect -11150 95910 -11140 95980
rect -11360 95860 -11140 95910
rect -10860 96090 -10640 96140
rect -10860 96020 -10850 96090
rect -10650 96020 -10640 96090
rect -10860 95980 -10640 96020
rect -10860 95910 -10850 95980
rect -10650 95910 -10640 95980
rect -10860 95860 -10640 95910
rect -10360 96090 -10140 96140
rect -10360 96020 -10350 96090
rect -10150 96020 -10140 96090
rect -10360 95980 -10140 96020
rect -10360 95910 -10350 95980
rect -10150 95910 -10140 95980
rect -10360 95860 -10140 95910
rect -9860 96090 -9640 96140
rect -9860 96020 -9850 96090
rect -9650 96020 -9640 96090
rect -9860 95980 -9640 96020
rect -9860 95910 -9850 95980
rect -9650 95910 -9640 95980
rect -9860 95860 -9640 95910
rect -9360 96090 -9140 96140
rect -9360 96020 -9350 96090
rect -9150 96020 -9140 96090
rect -9360 95980 -9140 96020
rect -9360 95910 -9350 95980
rect -9150 95910 -9140 95980
rect -9360 95860 -9140 95910
rect -8860 96090 -8640 96140
rect -8860 96020 -8850 96090
rect -8650 96020 -8640 96090
rect -8860 95980 -8640 96020
rect -8860 95910 -8850 95980
rect -8650 95910 -8640 95980
rect -8860 95860 -8640 95910
rect -8360 96090 -8140 96140
rect -8360 96020 -8350 96090
rect -8150 96020 -8140 96090
rect -8360 95980 -8140 96020
rect -8360 95910 -8350 95980
rect -8150 95910 -8140 95980
rect -8360 95860 -8140 95910
rect -7860 96090 -7640 96140
rect -7860 96020 -7850 96090
rect -7650 96020 -7640 96090
rect -7860 95980 -7640 96020
rect -7860 95910 -7850 95980
rect -7650 95910 -7640 95980
rect -7860 95860 -7640 95910
rect -7360 96090 -7140 96140
rect -7360 96020 -7350 96090
rect -7150 96020 -7140 96090
rect -7360 95980 -7140 96020
rect -7360 95910 -7350 95980
rect -7150 95910 -7140 95980
rect -7360 95860 -7140 95910
rect -6860 96090 -6640 96140
rect -6860 96020 -6850 96090
rect -6650 96020 -6640 96090
rect -6860 95980 -6640 96020
rect -6860 95910 -6850 95980
rect -6650 95910 -6640 95980
rect -6860 95860 -6640 95910
rect -6360 96090 -6140 96140
rect -6360 96020 -6350 96090
rect -6150 96020 -6140 96090
rect -6360 95980 -6140 96020
rect -6360 95910 -6350 95980
rect -6150 95910 -6140 95980
rect -6360 95860 -6140 95910
rect -5860 96090 -5640 96140
rect -5860 96020 -5850 96090
rect -5650 96020 -5640 96090
rect -5860 95980 -5640 96020
rect -5860 95910 -5850 95980
rect -5650 95910 -5640 95980
rect -5860 95860 -5640 95910
rect -5360 96090 -5140 96140
rect -5360 96020 -5350 96090
rect -5150 96020 -5140 96090
rect -5360 95980 -5140 96020
rect -5360 95910 -5350 95980
rect -5150 95910 -5140 95980
rect -5360 95860 -5140 95910
rect -4860 96090 -4640 96140
rect -4860 96020 -4850 96090
rect -4650 96020 -4640 96090
rect -4860 95980 -4640 96020
rect -4860 95910 -4850 95980
rect -4650 95910 -4640 95980
rect -4860 95860 -4640 95910
rect -4360 96090 -4140 96140
rect -4360 96020 -4350 96090
rect -4150 96020 -4140 96090
rect -4360 95980 -4140 96020
rect -4360 95910 -4350 95980
rect -4150 95910 -4140 95980
rect -4360 95860 -4140 95910
rect -3860 96090 -3640 96140
rect -3860 96020 -3850 96090
rect -3650 96020 -3640 96090
rect -3860 95980 -3640 96020
rect -3860 95910 -3850 95980
rect -3650 95910 -3640 95980
rect -3860 95860 -3640 95910
rect -3360 96090 -3140 96140
rect -3360 96020 -3350 96090
rect -3150 96020 -3140 96090
rect -3360 95980 -3140 96020
rect -3360 95910 -3350 95980
rect -3150 95910 -3140 95980
rect -3360 95860 -3140 95910
rect -2860 96090 -2640 96140
rect -2860 96020 -2850 96090
rect -2650 96020 -2640 96090
rect -2860 95980 -2640 96020
rect -2860 95910 -2850 95980
rect -2650 95910 -2640 95980
rect -2860 95860 -2640 95910
rect -2360 96090 -2140 96140
rect -2360 96020 -2350 96090
rect -2150 96020 -2140 96090
rect -2360 95980 -2140 96020
rect -2360 95910 -2350 95980
rect -2150 95910 -2140 95980
rect -2360 95860 -2140 95910
rect -1860 96090 -1640 96140
rect -1860 96020 -1850 96090
rect -1650 96020 -1640 96090
rect -1860 95980 -1640 96020
rect -1860 95910 -1850 95980
rect -1650 95910 -1640 95980
rect -1860 95860 -1640 95910
rect -1360 96090 -1140 96140
rect -1360 96020 -1350 96090
rect -1150 96020 -1140 96090
rect -1360 95980 -1140 96020
rect -1360 95910 -1350 95980
rect -1150 95910 -1140 95980
rect -1360 95860 -1140 95910
rect -860 96090 -640 96140
rect -860 96020 -850 96090
rect -650 96020 -640 96090
rect -860 95980 -640 96020
rect -860 95910 -850 95980
rect -650 95910 -640 95980
rect -860 95860 -640 95910
rect -360 96090 -140 96140
rect -360 96020 -350 96090
rect -150 96020 -140 96090
rect -360 95980 -140 96020
rect -360 95910 -350 95980
rect -150 95910 -140 95980
rect -360 95860 -140 95910
rect 140 96090 360 96140
rect 140 96020 150 96090
rect 350 96020 360 96090
rect 140 95980 360 96020
rect 140 95910 150 95980
rect 350 95910 360 95980
rect 140 95860 360 95910
rect 640 96090 860 96140
rect 640 96020 650 96090
rect 850 96020 860 96090
rect 640 95980 860 96020
rect 640 95910 650 95980
rect 850 95910 860 95980
rect 640 95860 860 95910
rect 1140 96090 1360 96140
rect 1140 96020 1150 96090
rect 1350 96020 1360 96090
rect 1140 95980 1360 96020
rect 1140 95910 1150 95980
rect 1350 95910 1360 95980
rect 1140 95860 1360 95910
rect 1640 96090 1860 96140
rect 1640 96020 1650 96090
rect 1850 96020 1860 96090
rect 1640 95980 1860 96020
rect 1640 95910 1650 95980
rect 1850 95910 1860 95980
rect 1640 95860 1860 95910
rect 2140 96090 2360 96140
rect 2140 96020 2150 96090
rect 2350 96020 2360 96090
rect 2140 95980 2360 96020
rect 2140 95910 2150 95980
rect 2350 95910 2360 95980
rect 2140 95860 2360 95910
rect 2640 96090 2860 96140
rect 2640 96020 2650 96090
rect 2850 96020 2860 96090
rect 2640 95980 2860 96020
rect 2640 95910 2650 95980
rect 2850 95910 2860 95980
rect 2640 95860 2860 95910
rect 3140 96090 3360 96140
rect 3140 96020 3150 96090
rect 3350 96020 3360 96090
rect 3140 95980 3360 96020
rect 3140 95910 3150 95980
rect 3350 95910 3360 95980
rect 3140 95860 3360 95910
rect 3640 96090 3860 96140
rect 3640 96020 3650 96090
rect 3850 96020 3860 96090
rect 3640 95980 3860 96020
rect 3640 95910 3650 95980
rect 3850 95910 3860 95980
rect 3640 95860 3860 95910
rect 4140 96090 4360 96140
rect 4140 96020 4150 96090
rect 4350 96020 4360 96090
rect 4140 95980 4360 96020
rect 4140 95910 4150 95980
rect 4350 95910 4360 95980
rect 4140 95860 4360 95910
rect 4640 96090 4860 96140
rect 4640 96020 4650 96090
rect 4850 96020 4860 96090
rect 4640 95980 4860 96020
rect 4640 95910 4650 95980
rect 4850 95910 4860 95980
rect 4640 95860 4860 95910
rect 5140 96090 5360 96140
rect 5140 96020 5150 96090
rect 5350 96020 5360 96090
rect 5140 95980 5360 96020
rect 5140 95910 5150 95980
rect 5350 95910 5360 95980
rect 5140 95860 5360 95910
rect 5640 96090 5860 96140
rect 5640 96020 5650 96090
rect 5850 96020 5860 96090
rect 5640 95980 5860 96020
rect 5640 95910 5650 95980
rect 5850 95910 5860 95980
rect 5640 95860 5860 95910
rect 6140 96090 6360 96140
rect 6140 96020 6150 96090
rect 6350 96020 6360 96090
rect 6140 95980 6360 96020
rect 6140 95910 6150 95980
rect 6350 95910 6360 95980
rect 6140 95860 6360 95910
rect 6640 96090 6860 96140
rect 6640 96020 6650 96090
rect 6850 96020 6860 96090
rect 6640 95980 6860 96020
rect 6640 95910 6650 95980
rect 6850 95910 6860 95980
rect 6640 95860 6860 95910
rect 7140 96090 7360 96140
rect 7140 96020 7150 96090
rect 7350 96020 7360 96090
rect 7140 95980 7360 96020
rect 7140 95910 7150 95980
rect 7350 95910 7360 95980
rect 7140 95860 7360 95910
rect 7640 96090 7860 96140
rect 7640 96020 7650 96090
rect 7850 96020 7860 96090
rect 7640 95980 7860 96020
rect 7640 95910 7650 95980
rect 7850 95910 7860 95980
rect 7640 95860 7860 95910
rect 8140 96090 8360 96140
rect 8140 96020 8150 96090
rect 8350 96020 8360 96090
rect 8140 95980 8360 96020
rect 8140 95910 8150 95980
rect 8350 95910 8360 95980
rect 8140 95860 8360 95910
rect 8640 96090 8860 96140
rect 8640 96020 8650 96090
rect 8850 96020 8860 96090
rect 8640 95980 8860 96020
rect 8640 95910 8650 95980
rect 8850 95910 8860 95980
rect 8640 95860 8860 95910
rect 9140 96090 9360 96140
rect 9140 96020 9150 96090
rect 9350 96020 9360 96090
rect 9140 95980 9360 96020
rect 9140 95910 9150 95980
rect 9350 95910 9360 95980
rect 9140 95860 9360 95910
rect 9640 96090 9860 96140
rect 9640 96020 9650 96090
rect 9850 96020 9860 96090
rect 9640 95980 9860 96020
rect 9640 95910 9650 95980
rect 9850 95910 9860 95980
rect 9640 95860 9860 95910
rect 10140 96090 10360 96140
rect 10140 96020 10150 96090
rect 10350 96020 10360 96090
rect 10140 95980 10360 96020
rect 10140 95910 10150 95980
rect 10350 95910 10360 95980
rect 10140 95860 10360 95910
rect 10640 96090 10860 96140
rect 10640 96020 10650 96090
rect 10850 96020 10860 96090
rect 10640 95980 10860 96020
rect 10640 95910 10650 95980
rect 10850 95910 10860 95980
rect 10640 95860 10860 95910
rect 11140 96090 11360 96140
rect 11140 96020 11150 96090
rect 11350 96020 11360 96090
rect 11140 95980 11360 96020
rect 11140 95910 11150 95980
rect 11350 95910 11360 95980
rect 11140 95860 11360 95910
rect 11640 96090 11860 96140
rect 11640 96020 11650 96090
rect 11850 96020 11860 96090
rect 11640 95980 11860 96020
rect 11640 95910 11650 95980
rect 11850 95910 11860 95980
rect 11640 95860 11860 95910
rect 12140 96090 12360 96140
rect 12140 96020 12150 96090
rect 12350 96020 12360 96090
rect 12140 95980 12360 96020
rect 12140 95910 12150 95980
rect 12350 95910 12360 95980
rect 12140 95860 12360 95910
rect 12640 96090 12860 96140
rect 12640 96020 12650 96090
rect 12850 96020 12860 96090
rect 12640 95980 12860 96020
rect 12640 95910 12650 95980
rect 12850 95910 12860 95980
rect 12640 95860 12860 95910
rect 13140 96090 13360 96140
rect 13140 96020 13150 96090
rect 13350 96020 13360 96090
rect 13140 95980 13360 96020
rect 13140 95910 13150 95980
rect 13350 95910 13360 95980
rect 13140 95860 13360 95910
rect 13640 96090 13860 96140
rect 13640 96020 13650 96090
rect 13850 96020 13860 96090
rect 13640 95980 13860 96020
rect 13640 95910 13650 95980
rect 13850 95910 13860 95980
rect 13640 95860 13860 95910
rect 14140 96090 14360 96140
rect 14140 96020 14150 96090
rect 14350 96020 14360 96090
rect 14140 95980 14360 96020
rect 14140 95910 14150 95980
rect 14350 95910 14360 95980
rect 14140 95860 14360 95910
rect 14640 96090 14860 96140
rect 14640 96020 14650 96090
rect 14850 96020 14860 96090
rect 14640 95980 14860 96020
rect 14640 95910 14650 95980
rect 14850 95910 14860 95980
rect 14640 95860 14860 95910
rect 15140 96090 15360 96140
rect 15140 96020 15150 96090
rect 15350 96020 15360 96090
rect 15140 95980 15360 96020
rect 15140 95910 15150 95980
rect 15350 95910 15360 95980
rect 15140 95860 15360 95910
rect 15640 96090 15860 96140
rect 15640 96020 15650 96090
rect 15850 96020 15860 96090
rect 15640 95980 15860 96020
rect 15640 95910 15650 95980
rect 15850 95910 15860 95980
rect 15640 95860 15860 95910
rect 16140 96090 16360 96140
rect 16140 96020 16150 96090
rect 16350 96020 16360 96090
rect 16140 95980 16360 96020
rect 16140 95910 16150 95980
rect 16350 95910 16360 95980
rect 16140 95860 16360 95910
rect 16640 96090 16860 96140
rect 16640 96020 16650 96090
rect 16850 96020 16860 96090
rect 16640 95980 16860 96020
rect 16640 95910 16650 95980
rect 16850 95910 16860 95980
rect 16640 95860 16860 95910
rect 17140 96090 17360 96140
rect 17140 96020 17150 96090
rect 17350 96020 17360 96090
rect 17140 95980 17360 96020
rect 17140 95910 17150 95980
rect 17350 95910 17360 95980
rect 17140 95860 17360 95910
rect 17640 96090 17860 96140
rect 17640 96020 17650 96090
rect 17850 96020 17860 96090
rect 17640 95980 17860 96020
rect 17640 95910 17650 95980
rect 17850 95910 17860 95980
rect 17640 95860 17860 95910
rect 18140 96090 18360 96140
rect 18140 96020 18150 96090
rect 18350 96020 18360 96090
rect 18140 95980 18360 96020
rect 18140 95910 18150 95980
rect 18350 95910 18360 95980
rect 18140 95860 18360 95910
rect 18640 96090 18860 96140
rect 18640 96020 18650 96090
rect 18850 96020 18860 96090
rect 18640 95980 18860 96020
rect 18640 95910 18650 95980
rect 18850 95910 18860 95980
rect 18640 95860 18860 95910
rect 19140 96090 19360 96140
rect 19140 96020 19150 96090
rect 19350 96020 19360 96090
rect 19140 95980 19360 96020
rect 19140 95910 19150 95980
rect 19350 95910 19360 95980
rect 19140 95860 19360 95910
rect 19640 96090 19860 96140
rect 19640 96020 19650 96090
rect 19850 96020 19860 96090
rect 19640 95980 19860 96020
rect 19640 95910 19650 95980
rect 19850 95910 19860 95980
rect 19640 95860 19860 95910
rect -16000 95850 20000 95860
rect -16000 95650 -15980 95850
rect -15910 95650 -15590 95850
rect -15520 95650 -15480 95850
rect -15410 95650 -15090 95850
rect -15020 95650 -14980 95850
rect -14910 95650 -14590 95850
rect -14520 95650 -14480 95850
rect -14410 95650 -14090 95850
rect -14020 95650 -13980 95850
rect -13910 95650 -13590 95850
rect -13520 95650 -13480 95850
rect -13410 95650 -13090 95850
rect -13020 95650 -12980 95850
rect -12910 95650 -12590 95850
rect -12520 95650 -12480 95850
rect -12410 95650 -12090 95850
rect -12020 95650 -11980 95850
rect -11910 95650 -11590 95850
rect -11520 95650 -11480 95850
rect -11410 95650 -11090 95850
rect -11020 95650 -10980 95850
rect -10910 95650 -10590 95850
rect -10520 95650 -10480 95850
rect -10410 95650 -10090 95850
rect -10020 95650 -9980 95850
rect -9910 95650 -9590 95850
rect -9520 95650 -9480 95850
rect -9410 95650 -9090 95850
rect -9020 95650 -8980 95850
rect -8910 95650 -8590 95850
rect -8520 95650 -8480 95850
rect -8410 95650 -8090 95850
rect -8020 95650 -7980 95850
rect -7910 95650 -7590 95850
rect -7520 95650 -7480 95850
rect -7410 95650 -7090 95850
rect -7020 95650 -6980 95850
rect -6910 95650 -6590 95850
rect -6520 95650 -6480 95850
rect -6410 95650 -6090 95850
rect -6020 95650 -5980 95850
rect -5910 95650 -5590 95850
rect -5520 95650 -5480 95850
rect -5410 95650 -5090 95850
rect -5020 95650 -4980 95850
rect -4910 95650 -4590 95850
rect -4520 95650 -4480 95850
rect -4410 95650 -4090 95850
rect -4020 95650 -3980 95850
rect -3910 95650 -3590 95850
rect -3520 95650 -3480 95850
rect -3410 95650 -3090 95850
rect -3020 95650 -2980 95850
rect -2910 95650 -2590 95850
rect -2520 95650 -2480 95850
rect -2410 95650 -2090 95850
rect -2020 95650 -1980 95850
rect -1910 95650 -1590 95850
rect -1520 95650 -1480 95850
rect -1410 95650 -1090 95850
rect -1020 95650 -980 95850
rect -910 95650 -590 95850
rect -520 95650 -480 95850
rect -410 95650 -90 95850
rect -20 95650 20 95850
rect 90 95650 410 95850
rect 480 95650 520 95850
rect 590 95650 910 95850
rect 980 95650 1020 95850
rect 1090 95650 1410 95850
rect 1480 95650 1520 95850
rect 1590 95650 1910 95850
rect 1980 95650 2020 95850
rect 2090 95650 2410 95850
rect 2480 95650 2520 95850
rect 2590 95650 2910 95850
rect 2980 95650 3020 95850
rect 3090 95650 3410 95850
rect 3480 95650 3520 95850
rect 3590 95650 3910 95850
rect 3980 95650 4020 95850
rect 4090 95650 4410 95850
rect 4480 95650 4520 95850
rect 4590 95650 4910 95850
rect 4980 95650 5020 95850
rect 5090 95650 5410 95850
rect 5480 95650 5520 95850
rect 5590 95650 5910 95850
rect 5980 95650 6020 95850
rect 6090 95650 6410 95850
rect 6480 95650 6520 95850
rect 6590 95650 6910 95850
rect 6980 95650 7020 95850
rect 7090 95650 7410 95850
rect 7480 95650 7520 95850
rect 7590 95650 7910 95850
rect 7980 95650 8020 95850
rect 8090 95650 8410 95850
rect 8480 95650 8520 95850
rect 8590 95650 8910 95850
rect 8980 95650 9020 95850
rect 9090 95650 9410 95850
rect 9480 95650 9520 95850
rect 9590 95650 9910 95850
rect 9980 95650 10020 95850
rect 10090 95650 10410 95850
rect 10480 95650 10520 95850
rect 10590 95650 10910 95850
rect 10980 95650 11020 95850
rect 11090 95650 11410 95850
rect 11480 95650 11520 95850
rect 11590 95650 11910 95850
rect 11980 95650 12020 95850
rect 12090 95650 12410 95850
rect 12480 95650 12520 95850
rect 12590 95650 12910 95850
rect 12980 95650 13020 95850
rect 13090 95650 13410 95850
rect 13480 95650 13520 95850
rect 13590 95650 13910 95850
rect 13980 95650 14020 95850
rect 14090 95650 14410 95850
rect 14480 95650 14520 95850
rect 14590 95650 14910 95850
rect 14980 95650 15020 95850
rect 15090 95650 15410 95850
rect 15480 95650 15520 95850
rect 15590 95650 15910 95850
rect 15980 95650 16020 95850
rect 16090 95650 16410 95850
rect 16480 95650 16520 95850
rect 16590 95650 16910 95850
rect 16980 95650 17020 95850
rect 17090 95650 17410 95850
rect 17480 95650 17520 95850
rect 17590 95650 17910 95850
rect 17980 95650 18020 95850
rect 18090 95650 18410 95850
rect 18480 95650 18520 95850
rect 18590 95650 18910 95850
rect 18980 95650 19020 95850
rect 19090 95650 19410 95850
rect 19480 95650 19520 95850
rect 19590 95650 19910 95850
rect 19980 95650 20000 95850
rect -16000 95640 20000 95650
rect -15860 95590 -15640 95640
rect -15860 95520 -15850 95590
rect -15650 95520 -15640 95590
rect -15860 95480 -15640 95520
rect -15860 95410 -15850 95480
rect -15650 95410 -15640 95480
rect -15860 95360 -15640 95410
rect -15360 95590 -15140 95640
rect -15360 95520 -15350 95590
rect -15150 95520 -15140 95590
rect -15360 95480 -15140 95520
rect -15360 95410 -15350 95480
rect -15150 95410 -15140 95480
rect -15360 95360 -15140 95410
rect -14860 95590 -14640 95640
rect -14860 95520 -14850 95590
rect -14650 95520 -14640 95590
rect -14860 95480 -14640 95520
rect -14860 95410 -14850 95480
rect -14650 95410 -14640 95480
rect -14860 95360 -14640 95410
rect -14360 95590 -14140 95640
rect -14360 95520 -14350 95590
rect -14150 95520 -14140 95590
rect -14360 95480 -14140 95520
rect -14360 95410 -14350 95480
rect -14150 95410 -14140 95480
rect -14360 95360 -14140 95410
rect -13860 95590 -13640 95640
rect -13860 95520 -13850 95590
rect -13650 95520 -13640 95590
rect -13860 95480 -13640 95520
rect -13860 95410 -13850 95480
rect -13650 95410 -13640 95480
rect -13860 95360 -13640 95410
rect -13360 95590 -13140 95640
rect -13360 95520 -13350 95590
rect -13150 95520 -13140 95590
rect -13360 95480 -13140 95520
rect -13360 95410 -13350 95480
rect -13150 95410 -13140 95480
rect -13360 95360 -13140 95410
rect -12860 95590 -12640 95640
rect -12860 95520 -12850 95590
rect -12650 95520 -12640 95590
rect -12860 95480 -12640 95520
rect -12860 95410 -12850 95480
rect -12650 95410 -12640 95480
rect -12860 95360 -12640 95410
rect -12360 95590 -12140 95640
rect -12360 95520 -12350 95590
rect -12150 95520 -12140 95590
rect -12360 95480 -12140 95520
rect -12360 95410 -12350 95480
rect -12150 95410 -12140 95480
rect -12360 95360 -12140 95410
rect -11860 95590 -11640 95640
rect -11860 95520 -11850 95590
rect -11650 95520 -11640 95590
rect -11860 95480 -11640 95520
rect -11860 95410 -11850 95480
rect -11650 95410 -11640 95480
rect -11860 95360 -11640 95410
rect -11360 95590 -11140 95640
rect -11360 95520 -11350 95590
rect -11150 95520 -11140 95590
rect -11360 95480 -11140 95520
rect -11360 95410 -11350 95480
rect -11150 95410 -11140 95480
rect -11360 95360 -11140 95410
rect -10860 95590 -10640 95640
rect -10860 95520 -10850 95590
rect -10650 95520 -10640 95590
rect -10860 95480 -10640 95520
rect -10860 95410 -10850 95480
rect -10650 95410 -10640 95480
rect -10860 95360 -10640 95410
rect -10360 95590 -10140 95640
rect -10360 95520 -10350 95590
rect -10150 95520 -10140 95590
rect -10360 95480 -10140 95520
rect -10360 95410 -10350 95480
rect -10150 95410 -10140 95480
rect -10360 95360 -10140 95410
rect -9860 95590 -9640 95640
rect -9860 95520 -9850 95590
rect -9650 95520 -9640 95590
rect -9860 95480 -9640 95520
rect -9860 95410 -9850 95480
rect -9650 95410 -9640 95480
rect -9860 95360 -9640 95410
rect -9360 95590 -9140 95640
rect -9360 95520 -9350 95590
rect -9150 95520 -9140 95590
rect -9360 95480 -9140 95520
rect -9360 95410 -9350 95480
rect -9150 95410 -9140 95480
rect -9360 95360 -9140 95410
rect -8860 95590 -8640 95640
rect -8860 95520 -8850 95590
rect -8650 95520 -8640 95590
rect -8860 95480 -8640 95520
rect -8860 95410 -8850 95480
rect -8650 95410 -8640 95480
rect -8860 95360 -8640 95410
rect -8360 95590 -8140 95640
rect -8360 95520 -8350 95590
rect -8150 95520 -8140 95590
rect -8360 95480 -8140 95520
rect -8360 95410 -8350 95480
rect -8150 95410 -8140 95480
rect -8360 95360 -8140 95410
rect -7860 95590 -7640 95640
rect -7860 95520 -7850 95590
rect -7650 95520 -7640 95590
rect -7860 95480 -7640 95520
rect -7860 95410 -7850 95480
rect -7650 95410 -7640 95480
rect -7860 95360 -7640 95410
rect -7360 95590 -7140 95640
rect -7360 95520 -7350 95590
rect -7150 95520 -7140 95590
rect -7360 95480 -7140 95520
rect -7360 95410 -7350 95480
rect -7150 95410 -7140 95480
rect -7360 95360 -7140 95410
rect -6860 95590 -6640 95640
rect -6860 95520 -6850 95590
rect -6650 95520 -6640 95590
rect -6860 95480 -6640 95520
rect -6860 95410 -6850 95480
rect -6650 95410 -6640 95480
rect -6860 95360 -6640 95410
rect -6360 95590 -6140 95640
rect -6360 95520 -6350 95590
rect -6150 95520 -6140 95590
rect -6360 95480 -6140 95520
rect -6360 95410 -6350 95480
rect -6150 95410 -6140 95480
rect -6360 95360 -6140 95410
rect -5860 95590 -5640 95640
rect -5860 95520 -5850 95590
rect -5650 95520 -5640 95590
rect -5860 95480 -5640 95520
rect -5860 95410 -5850 95480
rect -5650 95410 -5640 95480
rect -5860 95360 -5640 95410
rect -5360 95590 -5140 95640
rect -5360 95520 -5350 95590
rect -5150 95520 -5140 95590
rect -5360 95480 -5140 95520
rect -5360 95410 -5350 95480
rect -5150 95410 -5140 95480
rect -5360 95360 -5140 95410
rect -4860 95590 -4640 95640
rect -4860 95520 -4850 95590
rect -4650 95520 -4640 95590
rect -4860 95480 -4640 95520
rect -4860 95410 -4850 95480
rect -4650 95410 -4640 95480
rect -4860 95360 -4640 95410
rect -4360 95590 -4140 95640
rect -4360 95520 -4350 95590
rect -4150 95520 -4140 95590
rect -4360 95480 -4140 95520
rect -4360 95410 -4350 95480
rect -4150 95410 -4140 95480
rect -4360 95360 -4140 95410
rect -3860 95590 -3640 95640
rect -3860 95520 -3850 95590
rect -3650 95520 -3640 95590
rect -3860 95480 -3640 95520
rect -3860 95410 -3850 95480
rect -3650 95410 -3640 95480
rect -3860 95360 -3640 95410
rect -3360 95590 -3140 95640
rect -3360 95520 -3350 95590
rect -3150 95520 -3140 95590
rect -3360 95480 -3140 95520
rect -3360 95410 -3350 95480
rect -3150 95410 -3140 95480
rect -3360 95360 -3140 95410
rect -2860 95590 -2640 95640
rect -2860 95520 -2850 95590
rect -2650 95520 -2640 95590
rect -2860 95480 -2640 95520
rect -2860 95410 -2850 95480
rect -2650 95410 -2640 95480
rect -2860 95360 -2640 95410
rect -2360 95590 -2140 95640
rect -2360 95520 -2350 95590
rect -2150 95520 -2140 95590
rect -2360 95480 -2140 95520
rect -2360 95410 -2350 95480
rect -2150 95410 -2140 95480
rect -2360 95360 -2140 95410
rect -1860 95590 -1640 95640
rect -1860 95520 -1850 95590
rect -1650 95520 -1640 95590
rect -1860 95480 -1640 95520
rect -1860 95410 -1850 95480
rect -1650 95410 -1640 95480
rect -1860 95360 -1640 95410
rect -1360 95590 -1140 95640
rect -1360 95520 -1350 95590
rect -1150 95520 -1140 95590
rect -1360 95480 -1140 95520
rect -1360 95410 -1350 95480
rect -1150 95410 -1140 95480
rect -1360 95360 -1140 95410
rect -860 95590 -640 95640
rect -860 95520 -850 95590
rect -650 95520 -640 95590
rect -860 95480 -640 95520
rect -860 95410 -850 95480
rect -650 95410 -640 95480
rect -860 95360 -640 95410
rect -360 95590 -140 95640
rect -360 95520 -350 95590
rect -150 95520 -140 95590
rect -360 95480 -140 95520
rect -360 95410 -350 95480
rect -150 95410 -140 95480
rect -360 95360 -140 95410
rect 140 95590 360 95640
rect 140 95520 150 95590
rect 350 95520 360 95590
rect 140 95480 360 95520
rect 140 95410 150 95480
rect 350 95410 360 95480
rect 140 95360 360 95410
rect 640 95590 860 95640
rect 640 95520 650 95590
rect 850 95520 860 95590
rect 640 95480 860 95520
rect 640 95410 650 95480
rect 850 95410 860 95480
rect 640 95360 860 95410
rect 1140 95590 1360 95640
rect 1140 95520 1150 95590
rect 1350 95520 1360 95590
rect 1140 95480 1360 95520
rect 1140 95410 1150 95480
rect 1350 95410 1360 95480
rect 1140 95360 1360 95410
rect 1640 95590 1860 95640
rect 1640 95520 1650 95590
rect 1850 95520 1860 95590
rect 1640 95480 1860 95520
rect 1640 95410 1650 95480
rect 1850 95410 1860 95480
rect 1640 95360 1860 95410
rect 2140 95590 2360 95640
rect 2140 95520 2150 95590
rect 2350 95520 2360 95590
rect 2140 95480 2360 95520
rect 2140 95410 2150 95480
rect 2350 95410 2360 95480
rect 2140 95360 2360 95410
rect 2640 95590 2860 95640
rect 2640 95520 2650 95590
rect 2850 95520 2860 95590
rect 2640 95480 2860 95520
rect 2640 95410 2650 95480
rect 2850 95410 2860 95480
rect 2640 95360 2860 95410
rect 3140 95590 3360 95640
rect 3140 95520 3150 95590
rect 3350 95520 3360 95590
rect 3140 95480 3360 95520
rect 3140 95410 3150 95480
rect 3350 95410 3360 95480
rect 3140 95360 3360 95410
rect 3640 95590 3860 95640
rect 3640 95520 3650 95590
rect 3850 95520 3860 95590
rect 3640 95480 3860 95520
rect 3640 95410 3650 95480
rect 3850 95410 3860 95480
rect 3640 95360 3860 95410
rect 4140 95590 4360 95640
rect 4140 95520 4150 95590
rect 4350 95520 4360 95590
rect 4140 95480 4360 95520
rect 4140 95410 4150 95480
rect 4350 95410 4360 95480
rect 4140 95360 4360 95410
rect 4640 95590 4860 95640
rect 4640 95520 4650 95590
rect 4850 95520 4860 95590
rect 4640 95480 4860 95520
rect 4640 95410 4650 95480
rect 4850 95410 4860 95480
rect 4640 95360 4860 95410
rect 5140 95590 5360 95640
rect 5140 95520 5150 95590
rect 5350 95520 5360 95590
rect 5140 95480 5360 95520
rect 5140 95410 5150 95480
rect 5350 95410 5360 95480
rect 5140 95360 5360 95410
rect 5640 95590 5860 95640
rect 5640 95520 5650 95590
rect 5850 95520 5860 95590
rect 5640 95480 5860 95520
rect 5640 95410 5650 95480
rect 5850 95410 5860 95480
rect 5640 95360 5860 95410
rect 6140 95590 6360 95640
rect 6140 95520 6150 95590
rect 6350 95520 6360 95590
rect 6140 95480 6360 95520
rect 6140 95410 6150 95480
rect 6350 95410 6360 95480
rect 6140 95360 6360 95410
rect 6640 95590 6860 95640
rect 6640 95520 6650 95590
rect 6850 95520 6860 95590
rect 6640 95480 6860 95520
rect 6640 95410 6650 95480
rect 6850 95410 6860 95480
rect 6640 95360 6860 95410
rect 7140 95590 7360 95640
rect 7140 95520 7150 95590
rect 7350 95520 7360 95590
rect 7140 95480 7360 95520
rect 7140 95410 7150 95480
rect 7350 95410 7360 95480
rect 7140 95360 7360 95410
rect 7640 95590 7860 95640
rect 7640 95520 7650 95590
rect 7850 95520 7860 95590
rect 7640 95480 7860 95520
rect 7640 95410 7650 95480
rect 7850 95410 7860 95480
rect 7640 95360 7860 95410
rect 8140 95590 8360 95640
rect 8140 95520 8150 95590
rect 8350 95520 8360 95590
rect 8140 95480 8360 95520
rect 8140 95410 8150 95480
rect 8350 95410 8360 95480
rect 8140 95360 8360 95410
rect 8640 95590 8860 95640
rect 8640 95520 8650 95590
rect 8850 95520 8860 95590
rect 8640 95480 8860 95520
rect 8640 95410 8650 95480
rect 8850 95410 8860 95480
rect 8640 95360 8860 95410
rect 9140 95590 9360 95640
rect 9140 95520 9150 95590
rect 9350 95520 9360 95590
rect 9140 95480 9360 95520
rect 9140 95410 9150 95480
rect 9350 95410 9360 95480
rect 9140 95360 9360 95410
rect 9640 95590 9860 95640
rect 9640 95520 9650 95590
rect 9850 95520 9860 95590
rect 9640 95480 9860 95520
rect 9640 95410 9650 95480
rect 9850 95410 9860 95480
rect 9640 95360 9860 95410
rect 10140 95590 10360 95640
rect 10140 95520 10150 95590
rect 10350 95520 10360 95590
rect 10140 95480 10360 95520
rect 10140 95410 10150 95480
rect 10350 95410 10360 95480
rect 10140 95360 10360 95410
rect 10640 95590 10860 95640
rect 10640 95520 10650 95590
rect 10850 95520 10860 95590
rect 10640 95480 10860 95520
rect 10640 95410 10650 95480
rect 10850 95410 10860 95480
rect 10640 95360 10860 95410
rect 11140 95590 11360 95640
rect 11140 95520 11150 95590
rect 11350 95520 11360 95590
rect 11140 95480 11360 95520
rect 11140 95410 11150 95480
rect 11350 95410 11360 95480
rect 11140 95360 11360 95410
rect 11640 95590 11860 95640
rect 11640 95520 11650 95590
rect 11850 95520 11860 95590
rect 11640 95480 11860 95520
rect 11640 95410 11650 95480
rect 11850 95410 11860 95480
rect 11640 95360 11860 95410
rect 12140 95590 12360 95640
rect 12140 95520 12150 95590
rect 12350 95520 12360 95590
rect 12140 95480 12360 95520
rect 12140 95410 12150 95480
rect 12350 95410 12360 95480
rect 12140 95360 12360 95410
rect 12640 95590 12860 95640
rect 12640 95520 12650 95590
rect 12850 95520 12860 95590
rect 12640 95480 12860 95520
rect 12640 95410 12650 95480
rect 12850 95410 12860 95480
rect 12640 95360 12860 95410
rect 13140 95590 13360 95640
rect 13140 95520 13150 95590
rect 13350 95520 13360 95590
rect 13140 95480 13360 95520
rect 13140 95410 13150 95480
rect 13350 95410 13360 95480
rect 13140 95360 13360 95410
rect 13640 95590 13860 95640
rect 13640 95520 13650 95590
rect 13850 95520 13860 95590
rect 13640 95480 13860 95520
rect 13640 95410 13650 95480
rect 13850 95410 13860 95480
rect 13640 95360 13860 95410
rect 14140 95590 14360 95640
rect 14140 95520 14150 95590
rect 14350 95520 14360 95590
rect 14140 95480 14360 95520
rect 14140 95410 14150 95480
rect 14350 95410 14360 95480
rect 14140 95360 14360 95410
rect 14640 95590 14860 95640
rect 14640 95520 14650 95590
rect 14850 95520 14860 95590
rect 14640 95480 14860 95520
rect 14640 95410 14650 95480
rect 14850 95410 14860 95480
rect 14640 95360 14860 95410
rect 15140 95590 15360 95640
rect 15140 95520 15150 95590
rect 15350 95520 15360 95590
rect 15140 95480 15360 95520
rect 15140 95410 15150 95480
rect 15350 95410 15360 95480
rect 15140 95360 15360 95410
rect 15640 95590 15860 95640
rect 15640 95520 15650 95590
rect 15850 95520 15860 95590
rect 15640 95480 15860 95520
rect 15640 95410 15650 95480
rect 15850 95410 15860 95480
rect 15640 95360 15860 95410
rect 16140 95590 16360 95640
rect 16140 95520 16150 95590
rect 16350 95520 16360 95590
rect 16140 95480 16360 95520
rect 16140 95410 16150 95480
rect 16350 95410 16360 95480
rect 16140 95360 16360 95410
rect 16640 95590 16860 95640
rect 16640 95520 16650 95590
rect 16850 95520 16860 95590
rect 16640 95480 16860 95520
rect 16640 95410 16650 95480
rect 16850 95410 16860 95480
rect 16640 95360 16860 95410
rect 17140 95590 17360 95640
rect 17140 95520 17150 95590
rect 17350 95520 17360 95590
rect 17140 95480 17360 95520
rect 17140 95410 17150 95480
rect 17350 95410 17360 95480
rect 17140 95360 17360 95410
rect 17640 95590 17860 95640
rect 17640 95520 17650 95590
rect 17850 95520 17860 95590
rect 17640 95480 17860 95520
rect 17640 95410 17650 95480
rect 17850 95410 17860 95480
rect 17640 95360 17860 95410
rect 18140 95590 18360 95640
rect 18140 95520 18150 95590
rect 18350 95520 18360 95590
rect 18140 95480 18360 95520
rect 18140 95410 18150 95480
rect 18350 95410 18360 95480
rect 18140 95360 18360 95410
rect 18640 95590 18860 95640
rect 18640 95520 18650 95590
rect 18850 95520 18860 95590
rect 18640 95480 18860 95520
rect 18640 95410 18650 95480
rect 18850 95410 18860 95480
rect 18640 95360 18860 95410
rect 19140 95590 19360 95640
rect 19140 95520 19150 95590
rect 19350 95520 19360 95590
rect 19140 95480 19360 95520
rect 19140 95410 19150 95480
rect 19350 95410 19360 95480
rect 19140 95360 19360 95410
rect 19640 95590 19860 95640
rect 19640 95520 19650 95590
rect 19850 95520 19860 95590
rect 19640 95480 19860 95520
rect 19640 95410 19650 95480
rect 19850 95410 19860 95480
rect 19640 95360 19860 95410
rect -16000 95350 20000 95360
rect -16000 95150 -15980 95350
rect -15910 95150 -15590 95350
rect -15520 95150 -15480 95350
rect -15410 95150 -15090 95350
rect -15020 95150 -14980 95350
rect -14910 95150 -14590 95350
rect -14520 95150 -14480 95350
rect -14410 95150 -14090 95350
rect -14020 95150 -13980 95350
rect -13910 95150 -13590 95350
rect -13520 95150 -13480 95350
rect -13410 95150 -13090 95350
rect -13020 95150 -12980 95350
rect -12910 95150 -12590 95350
rect -12520 95150 -12480 95350
rect -12410 95150 -12090 95350
rect -12020 95150 -11980 95350
rect -11910 95150 -11590 95350
rect -11520 95150 -11480 95350
rect -11410 95150 -11090 95350
rect -11020 95150 -10980 95350
rect -10910 95150 -10590 95350
rect -10520 95150 -10480 95350
rect -10410 95150 -10090 95350
rect -10020 95150 -9980 95350
rect -9910 95150 -9590 95350
rect -9520 95150 -9480 95350
rect -9410 95150 -9090 95350
rect -9020 95150 -8980 95350
rect -8910 95150 -8590 95350
rect -8520 95150 -8480 95350
rect -8410 95150 -8090 95350
rect -8020 95150 -7980 95350
rect -7910 95150 -7590 95350
rect -7520 95150 -7480 95350
rect -7410 95150 -7090 95350
rect -7020 95150 -6980 95350
rect -6910 95150 -6590 95350
rect -6520 95150 -6480 95350
rect -6410 95150 -6090 95350
rect -6020 95150 -5980 95350
rect -5910 95150 -5590 95350
rect -5520 95150 -5480 95350
rect -5410 95150 -5090 95350
rect -5020 95150 -4980 95350
rect -4910 95150 -4590 95350
rect -4520 95150 -4480 95350
rect -4410 95150 -4090 95350
rect -4020 95150 -3980 95350
rect -3910 95150 -3590 95350
rect -3520 95150 -3480 95350
rect -3410 95150 -3090 95350
rect -3020 95150 -2980 95350
rect -2910 95150 -2590 95350
rect -2520 95150 -2480 95350
rect -2410 95150 -2090 95350
rect -2020 95150 -1980 95350
rect -1910 95150 -1590 95350
rect -1520 95150 -1480 95350
rect -1410 95150 -1090 95350
rect -1020 95150 -980 95350
rect -910 95150 -590 95350
rect -520 95150 -480 95350
rect -410 95150 -90 95350
rect -20 95150 20 95350
rect 90 95150 410 95350
rect 480 95150 520 95350
rect 590 95150 910 95350
rect 980 95150 1020 95350
rect 1090 95150 1410 95350
rect 1480 95150 1520 95350
rect 1590 95150 1910 95350
rect 1980 95150 2020 95350
rect 2090 95150 2410 95350
rect 2480 95150 2520 95350
rect 2590 95150 2910 95350
rect 2980 95150 3020 95350
rect 3090 95150 3410 95350
rect 3480 95150 3520 95350
rect 3590 95150 3910 95350
rect 3980 95150 4020 95350
rect 4090 95150 4410 95350
rect 4480 95150 4520 95350
rect 4590 95150 4910 95350
rect 4980 95150 5020 95350
rect 5090 95150 5410 95350
rect 5480 95150 5520 95350
rect 5590 95150 5910 95350
rect 5980 95150 6020 95350
rect 6090 95150 6410 95350
rect 6480 95150 6520 95350
rect 6590 95150 6910 95350
rect 6980 95150 7020 95350
rect 7090 95150 7410 95350
rect 7480 95150 7520 95350
rect 7590 95150 7910 95350
rect 7980 95150 8020 95350
rect 8090 95150 8410 95350
rect 8480 95150 8520 95350
rect 8590 95150 8910 95350
rect 8980 95150 9020 95350
rect 9090 95150 9410 95350
rect 9480 95150 9520 95350
rect 9590 95150 9910 95350
rect 9980 95150 10020 95350
rect 10090 95150 10410 95350
rect 10480 95150 10520 95350
rect 10590 95150 10910 95350
rect 10980 95150 11020 95350
rect 11090 95150 11410 95350
rect 11480 95150 11520 95350
rect 11590 95150 11910 95350
rect 11980 95150 12020 95350
rect 12090 95150 12410 95350
rect 12480 95150 12520 95350
rect 12590 95150 12910 95350
rect 12980 95150 13020 95350
rect 13090 95150 13410 95350
rect 13480 95150 13520 95350
rect 13590 95150 13910 95350
rect 13980 95150 14020 95350
rect 14090 95150 14410 95350
rect 14480 95150 14520 95350
rect 14590 95150 14910 95350
rect 14980 95150 15020 95350
rect 15090 95150 15410 95350
rect 15480 95150 15520 95350
rect 15590 95150 15910 95350
rect 15980 95150 16020 95350
rect 16090 95150 16410 95350
rect 16480 95150 16520 95350
rect 16590 95150 16910 95350
rect 16980 95150 17020 95350
rect 17090 95150 17410 95350
rect 17480 95150 17520 95350
rect 17590 95150 17910 95350
rect 17980 95150 18020 95350
rect 18090 95150 18410 95350
rect 18480 95150 18520 95350
rect 18590 95150 18910 95350
rect 18980 95150 19020 95350
rect 19090 95150 19410 95350
rect 19480 95150 19520 95350
rect 19590 95150 19910 95350
rect 19980 95150 20000 95350
rect -16000 95140 20000 95150
rect -15860 95090 -15640 95140
rect -15860 95020 -15850 95090
rect -15650 95020 -15640 95090
rect -15860 94980 -15640 95020
rect -15860 94910 -15850 94980
rect -15650 94910 -15640 94980
rect -15860 94860 -15640 94910
rect -15360 95090 -15140 95140
rect -15360 95020 -15350 95090
rect -15150 95020 -15140 95090
rect -15360 94980 -15140 95020
rect -15360 94910 -15350 94980
rect -15150 94910 -15140 94980
rect -15360 94860 -15140 94910
rect -14860 95090 -14640 95140
rect -14860 95020 -14850 95090
rect -14650 95020 -14640 95090
rect -14860 94980 -14640 95020
rect -14860 94910 -14850 94980
rect -14650 94910 -14640 94980
rect -14860 94860 -14640 94910
rect -14360 95090 -14140 95140
rect -14360 95020 -14350 95090
rect -14150 95020 -14140 95090
rect -14360 94980 -14140 95020
rect -14360 94910 -14350 94980
rect -14150 94910 -14140 94980
rect -14360 94860 -14140 94910
rect -13860 95090 -13640 95140
rect -13860 95020 -13850 95090
rect -13650 95020 -13640 95090
rect -13860 94980 -13640 95020
rect -13860 94910 -13850 94980
rect -13650 94910 -13640 94980
rect -13860 94860 -13640 94910
rect -13360 95090 -13140 95140
rect -13360 95020 -13350 95090
rect -13150 95020 -13140 95090
rect -13360 94980 -13140 95020
rect -13360 94910 -13350 94980
rect -13150 94910 -13140 94980
rect -13360 94860 -13140 94910
rect -12860 95090 -12640 95140
rect -12860 95020 -12850 95090
rect -12650 95020 -12640 95090
rect -12860 94980 -12640 95020
rect -12860 94910 -12850 94980
rect -12650 94910 -12640 94980
rect -12860 94860 -12640 94910
rect -12360 95090 -12140 95140
rect -12360 95020 -12350 95090
rect -12150 95020 -12140 95090
rect -12360 94980 -12140 95020
rect -12360 94910 -12350 94980
rect -12150 94910 -12140 94980
rect -12360 94860 -12140 94910
rect -11860 95090 -11640 95140
rect -11860 95020 -11850 95090
rect -11650 95020 -11640 95090
rect -11860 94980 -11640 95020
rect -11860 94910 -11850 94980
rect -11650 94910 -11640 94980
rect -11860 94860 -11640 94910
rect -11360 95090 -11140 95140
rect -11360 95020 -11350 95090
rect -11150 95020 -11140 95090
rect -11360 94980 -11140 95020
rect -11360 94910 -11350 94980
rect -11150 94910 -11140 94980
rect -11360 94860 -11140 94910
rect -10860 95090 -10640 95140
rect -10860 95020 -10850 95090
rect -10650 95020 -10640 95090
rect -10860 94980 -10640 95020
rect -10860 94910 -10850 94980
rect -10650 94910 -10640 94980
rect -10860 94860 -10640 94910
rect -10360 95090 -10140 95140
rect -10360 95020 -10350 95090
rect -10150 95020 -10140 95090
rect -10360 94980 -10140 95020
rect -10360 94910 -10350 94980
rect -10150 94910 -10140 94980
rect -10360 94860 -10140 94910
rect -9860 95090 -9640 95140
rect -9860 95020 -9850 95090
rect -9650 95020 -9640 95090
rect -9860 94980 -9640 95020
rect -9860 94910 -9850 94980
rect -9650 94910 -9640 94980
rect -9860 94860 -9640 94910
rect -9360 95090 -9140 95140
rect -9360 95020 -9350 95090
rect -9150 95020 -9140 95090
rect -9360 94980 -9140 95020
rect -9360 94910 -9350 94980
rect -9150 94910 -9140 94980
rect -9360 94860 -9140 94910
rect -8860 95090 -8640 95140
rect -8860 95020 -8850 95090
rect -8650 95020 -8640 95090
rect -8860 94980 -8640 95020
rect -8860 94910 -8850 94980
rect -8650 94910 -8640 94980
rect -8860 94860 -8640 94910
rect -8360 95090 -8140 95140
rect -8360 95020 -8350 95090
rect -8150 95020 -8140 95090
rect -8360 94980 -8140 95020
rect -8360 94910 -8350 94980
rect -8150 94910 -8140 94980
rect -8360 94860 -8140 94910
rect -7860 95090 -7640 95140
rect -7860 95020 -7850 95090
rect -7650 95020 -7640 95090
rect -7860 94980 -7640 95020
rect -7860 94910 -7850 94980
rect -7650 94910 -7640 94980
rect -7860 94860 -7640 94910
rect -7360 95090 -7140 95140
rect -7360 95020 -7350 95090
rect -7150 95020 -7140 95090
rect -7360 94980 -7140 95020
rect -7360 94910 -7350 94980
rect -7150 94910 -7140 94980
rect -7360 94860 -7140 94910
rect -6860 95090 -6640 95140
rect -6860 95020 -6850 95090
rect -6650 95020 -6640 95090
rect -6860 94980 -6640 95020
rect -6860 94910 -6850 94980
rect -6650 94910 -6640 94980
rect -6860 94860 -6640 94910
rect -6360 95090 -6140 95140
rect -6360 95020 -6350 95090
rect -6150 95020 -6140 95090
rect -6360 94980 -6140 95020
rect -6360 94910 -6350 94980
rect -6150 94910 -6140 94980
rect -6360 94860 -6140 94910
rect -5860 95090 -5640 95140
rect -5860 95020 -5850 95090
rect -5650 95020 -5640 95090
rect -5860 94980 -5640 95020
rect -5860 94910 -5850 94980
rect -5650 94910 -5640 94980
rect -5860 94860 -5640 94910
rect -5360 95090 -5140 95140
rect -5360 95020 -5350 95090
rect -5150 95020 -5140 95090
rect -5360 94980 -5140 95020
rect -5360 94910 -5350 94980
rect -5150 94910 -5140 94980
rect -5360 94860 -5140 94910
rect -4860 95090 -4640 95140
rect -4860 95020 -4850 95090
rect -4650 95020 -4640 95090
rect -4860 94980 -4640 95020
rect -4860 94910 -4850 94980
rect -4650 94910 -4640 94980
rect -4860 94860 -4640 94910
rect -4360 95090 -4140 95140
rect -4360 95020 -4350 95090
rect -4150 95020 -4140 95090
rect -4360 94980 -4140 95020
rect -4360 94910 -4350 94980
rect -4150 94910 -4140 94980
rect -4360 94860 -4140 94910
rect -3860 95090 -3640 95140
rect -3860 95020 -3850 95090
rect -3650 95020 -3640 95090
rect -3860 94980 -3640 95020
rect -3860 94910 -3850 94980
rect -3650 94910 -3640 94980
rect -3860 94860 -3640 94910
rect -3360 95090 -3140 95140
rect -3360 95020 -3350 95090
rect -3150 95020 -3140 95090
rect -3360 94980 -3140 95020
rect -3360 94910 -3350 94980
rect -3150 94910 -3140 94980
rect -3360 94860 -3140 94910
rect -2860 95090 -2640 95140
rect -2860 95020 -2850 95090
rect -2650 95020 -2640 95090
rect -2860 94980 -2640 95020
rect -2860 94910 -2850 94980
rect -2650 94910 -2640 94980
rect -2860 94860 -2640 94910
rect -2360 95090 -2140 95140
rect -2360 95020 -2350 95090
rect -2150 95020 -2140 95090
rect -2360 94980 -2140 95020
rect -2360 94910 -2350 94980
rect -2150 94910 -2140 94980
rect -2360 94860 -2140 94910
rect -1860 95090 -1640 95140
rect -1860 95020 -1850 95090
rect -1650 95020 -1640 95090
rect -1860 94980 -1640 95020
rect -1860 94910 -1850 94980
rect -1650 94910 -1640 94980
rect -1860 94860 -1640 94910
rect -1360 95090 -1140 95140
rect -1360 95020 -1350 95090
rect -1150 95020 -1140 95090
rect -1360 94980 -1140 95020
rect -1360 94910 -1350 94980
rect -1150 94910 -1140 94980
rect -1360 94860 -1140 94910
rect -860 95090 -640 95140
rect -860 95020 -850 95090
rect -650 95020 -640 95090
rect -860 94980 -640 95020
rect -860 94910 -850 94980
rect -650 94910 -640 94980
rect -860 94860 -640 94910
rect -360 95090 -140 95140
rect -360 95020 -350 95090
rect -150 95020 -140 95090
rect -360 94980 -140 95020
rect -360 94910 -350 94980
rect -150 94910 -140 94980
rect -360 94860 -140 94910
rect 140 95090 360 95140
rect 140 95020 150 95090
rect 350 95020 360 95090
rect 140 94980 360 95020
rect 140 94910 150 94980
rect 350 94910 360 94980
rect 140 94860 360 94910
rect 640 95090 860 95140
rect 640 95020 650 95090
rect 850 95020 860 95090
rect 640 94980 860 95020
rect 640 94910 650 94980
rect 850 94910 860 94980
rect 640 94860 860 94910
rect 1140 95090 1360 95140
rect 1140 95020 1150 95090
rect 1350 95020 1360 95090
rect 1140 94980 1360 95020
rect 1140 94910 1150 94980
rect 1350 94910 1360 94980
rect 1140 94860 1360 94910
rect 1640 95090 1860 95140
rect 1640 95020 1650 95090
rect 1850 95020 1860 95090
rect 1640 94980 1860 95020
rect 1640 94910 1650 94980
rect 1850 94910 1860 94980
rect 1640 94860 1860 94910
rect 2140 95090 2360 95140
rect 2140 95020 2150 95090
rect 2350 95020 2360 95090
rect 2140 94980 2360 95020
rect 2140 94910 2150 94980
rect 2350 94910 2360 94980
rect 2140 94860 2360 94910
rect 2640 95090 2860 95140
rect 2640 95020 2650 95090
rect 2850 95020 2860 95090
rect 2640 94980 2860 95020
rect 2640 94910 2650 94980
rect 2850 94910 2860 94980
rect 2640 94860 2860 94910
rect 3140 95090 3360 95140
rect 3140 95020 3150 95090
rect 3350 95020 3360 95090
rect 3140 94980 3360 95020
rect 3140 94910 3150 94980
rect 3350 94910 3360 94980
rect 3140 94860 3360 94910
rect 3640 95090 3860 95140
rect 3640 95020 3650 95090
rect 3850 95020 3860 95090
rect 3640 94980 3860 95020
rect 3640 94910 3650 94980
rect 3850 94910 3860 94980
rect 3640 94860 3860 94910
rect 4140 95090 4360 95140
rect 4140 95020 4150 95090
rect 4350 95020 4360 95090
rect 4140 94980 4360 95020
rect 4140 94910 4150 94980
rect 4350 94910 4360 94980
rect 4140 94860 4360 94910
rect 4640 95090 4860 95140
rect 4640 95020 4650 95090
rect 4850 95020 4860 95090
rect 4640 94980 4860 95020
rect 4640 94910 4650 94980
rect 4850 94910 4860 94980
rect 4640 94860 4860 94910
rect 5140 95090 5360 95140
rect 5140 95020 5150 95090
rect 5350 95020 5360 95090
rect 5140 94980 5360 95020
rect 5140 94910 5150 94980
rect 5350 94910 5360 94980
rect 5140 94860 5360 94910
rect 5640 95090 5860 95140
rect 5640 95020 5650 95090
rect 5850 95020 5860 95090
rect 5640 94980 5860 95020
rect 5640 94910 5650 94980
rect 5850 94910 5860 94980
rect 5640 94860 5860 94910
rect 6140 95090 6360 95140
rect 6140 95020 6150 95090
rect 6350 95020 6360 95090
rect 6140 94980 6360 95020
rect 6140 94910 6150 94980
rect 6350 94910 6360 94980
rect 6140 94860 6360 94910
rect 6640 95090 6860 95140
rect 6640 95020 6650 95090
rect 6850 95020 6860 95090
rect 6640 94980 6860 95020
rect 6640 94910 6650 94980
rect 6850 94910 6860 94980
rect 6640 94860 6860 94910
rect 7140 95090 7360 95140
rect 7140 95020 7150 95090
rect 7350 95020 7360 95090
rect 7140 94980 7360 95020
rect 7140 94910 7150 94980
rect 7350 94910 7360 94980
rect 7140 94860 7360 94910
rect 7640 95090 7860 95140
rect 7640 95020 7650 95090
rect 7850 95020 7860 95090
rect 7640 94980 7860 95020
rect 7640 94910 7650 94980
rect 7850 94910 7860 94980
rect 7640 94860 7860 94910
rect 8140 95090 8360 95140
rect 8140 95020 8150 95090
rect 8350 95020 8360 95090
rect 8140 94980 8360 95020
rect 8140 94910 8150 94980
rect 8350 94910 8360 94980
rect 8140 94860 8360 94910
rect 8640 95090 8860 95140
rect 8640 95020 8650 95090
rect 8850 95020 8860 95090
rect 8640 94980 8860 95020
rect 8640 94910 8650 94980
rect 8850 94910 8860 94980
rect 8640 94860 8860 94910
rect 9140 95090 9360 95140
rect 9140 95020 9150 95090
rect 9350 95020 9360 95090
rect 9140 94980 9360 95020
rect 9140 94910 9150 94980
rect 9350 94910 9360 94980
rect 9140 94860 9360 94910
rect 9640 95090 9860 95140
rect 9640 95020 9650 95090
rect 9850 95020 9860 95090
rect 9640 94980 9860 95020
rect 9640 94910 9650 94980
rect 9850 94910 9860 94980
rect 9640 94860 9860 94910
rect 10140 95090 10360 95140
rect 10140 95020 10150 95090
rect 10350 95020 10360 95090
rect 10140 94980 10360 95020
rect 10140 94910 10150 94980
rect 10350 94910 10360 94980
rect 10140 94860 10360 94910
rect 10640 95090 10860 95140
rect 10640 95020 10650 95090
rect 10850 95020 10860 95090
rect 10640 94980 10860 95020
rect 10640 94910 10650 94980
rect 10850 94910 10860 94980
rect 10640 94860 10860 94910
rect 11140 95090 11360 95140
rect 11140 95020 11150 95090
rect 11350 95020 11360 95090
rect 11140 94980 11360 95020
rect 11140 94910 11150 94980
rect 11350 94910 11360 94980
rect 11140 94860 11360 94910
rect 11640 95090 11860 95140
rect 11640 95020 11650 95090
rect 11850 95020 11860 95090
rect 11640 94980 11860 95020
rect 11640 94910 11650 94980
rect 11850 94910 11860 94980
rect 11640 94860 11860 94910
rect 12140 95090 12360 95140
rect 12140 95020 12150 95090
rect 12350 95020 12360 95090
rect 12140 94980 12360 95020
rect 12140 94910 12150 94980
rect 12350 94910 12360 94980
rect 12140 94860 12360 94910
rect 12640 95090 12860 95140
rect 12640 95020 12650 95090
rect 12850 95020 12860 95090
rect 12640 94980 12860 95020
rect 12640 94910 12650 94980
rect 12850 94910 12860 94980
rect 12640 94860 12860 94910
rect 13140 95090 13360 95140
rect 13140 95020 13150 95090
rect 13350 95020 13360 95090
rect 13140 94980 13360 95020
rect 13140 94910 13150 94980
rect 13350 94910 13360 94980
rect 13140 94860 13360 94910
rect 13640 95090 13860 95140
rect 13640 95020 13650 95090
rect 13850 95020 13860 95090
rect 13640 94980 13860 95020
rect 13640 94910 13650 94980
rect 13850 94910 13860 94980
rect 13640 94860 13860 94910
rect 14140 95090 14360 95140
rect 14140 95020 14150 95090
rect 14350 95020 14360 95090
rect 14140 94980 14360 95020
rect 14140 94910 14150 94980
rect 14350 94910 14360 94980
rect 14140 94860 14360 94910
rect 14640 95090 14860 95140
rect 14640 95020 14650 95090
rect 14850 95020 14860 95090
rect 14640 94980 14860 95020
rect 14640 94910 14650 94980
rect 14850 94910 14860 94980
rect 14640 94860 14860 94910
rect 15140 95090 15360 95140
rect 15140 95020 15150 95090
rect 15350 95020 15360 95090
rect 15140 94980 15360 95020
rect 15140 94910 15150 94980
rect 15350 94910 15360 94980
rect 15140 94860 15360 94910
rect 15640 95090 15860 95140
rect 15640 95020 15650 95090
rect 15850 95020 15860 95090
rect 15640 94980 15860 95020
rect 15640 94910 15650 94980
rect 15850 94910 15860 94980
rect 15640 94860 15860 94910
rect 16140 95090 16360 95140
rect 16140 95020 16150 95090
rect 16350 95020 16360 95090
rect 16140 94980 16360 95020
rect 16140 94910 16150 94980
rect 16350 94910 16360 94980
rect 16140 94860 16360 94910
rect 16640 95090 16860 95140
rect 16640 95020 16650 95090
rect 16850 95020 16860 95090
rect 16640 94980 16860 95020
rect 16640 94910 16650 94980
rect 16850 94910 16860 94980
rect 16640 94860 16860 94910
rect 17140 95090 17360 95140
rect 17140 95020 17150 95090
rect 17350 95020 17360 95090
rect 17140 94980 17360 95020
rect 17140 94910 17150 94980
rect 17350 94910 17360 94980
rect 17140 94860 17360 94910
rect 17640 95090 17860 95140
rect 17640 95020 17650 95090
rect 17850 95020 17860 95090
rect 17640 94980 17860 95020
rect 17640 94910 17650 94980
rect 17850 94910 17860 94980
rect 17640 94860 17860 94910
rect 18140 95090 18360 95140
rect 18140 95020 18150 95090
rect 18350 95020 18360 95090
rect 18140 94980 18360 95020
rect 18140 94910 18150 94980
rect 18350 94910 18360 94980
rect 18140 94860 18360 94910
rect 18640 95090 18860 95140
rect 18640 95020 18650 95090
rect 18850 95020 18860 95090
rect 18640 94980 18860 95020
rect 18640 94910 18650 94980
rect 18850 94910 18860 94980
rect 18640 94860 18860 94910
rect 19140 95090 19360 95140
rect 19140 95020 19150 95090
rect 19350 95020 19360 95090
rect 19140 94980 19360 95020
rect 19140 94910 19150 94980
rect 19350 94910 19360 94980
rect 19140 94860 19360 94910
rect 19640 95090 19860 95140
rect 19640 95020 19650 95090
rect 19850 95020 19860 95090
rect 19640 94980 19860 95020
rect 19640 94910 19650 94980
rect 19850 94910 19860 94980
rect 19640 94860 19860 94910
rect -16000 94850 20000 94860
rect -16000 94650 -15980 94850
rect -15910 94650 -15590 94850
rect -15520 94650 -15480 94850
rect -15410 94650 -15090 94850
rect -15020 94650 -14980 94850
rect -14910 94650 -14590 94850
rect -14520 94650 -14480 94850
rect -14410 94650 -14090 94850
rect -14020 94650 -13980 94850
rect -13910 94650 -13590 94850
rect -13520 94650 -13480 94850
rect -13410 94650 -13090 94850
rect -13020 94650 -12980 94850
rect -12910 94650 -12590 94850
rect -12520 94650 -12480 94850
rect -12410 94650 -12090 94850
rect -12020 94650 -11980 94850
rect -11910 94650 -11590 94850
rect -11520 94650 -11480 94850
rect -11410 94650 -11090 94850
rect -11020 94650 -10980 94850
rect -10910 94650 -10590 94850
rect -10520 94650 -10480 94850
rect -10410 94650 -10090 94850
rect -10020 94650 -9980 94850
rect -9910 94650 -9590 94850
rect -9520 94650 -9480 94850
rect -9410 94650 -9090 94850
rect -9020 94650 -8980 94850
rect -8910 94650 -8590 94850
rect -8520 94650 -8480 94850
rect -8410 94650 -8090 94850
rect -8020 94650 -7980 94850
rect -7910 94650 -7590 94850
rect -7520 94650 -7480 94850
rect -7410 94650 -7090 94850
rect -7020 94650 -6980 94850
rect -6910 94650 -6590 94850
rect -6520 94650 -6480 94850
rect -6410 94650 -6090 94850
rect -6020 94650 -5980 94850
rect -5910 94650 -5590 94850
rect -5520 94650 -5480 94850
rect -5410 94650 -5090 94850
rect -5020 94650 -4980 94850
rect -4910 94650 -4590 94850
rect -4520 94650 -4480 94850
rect -4410 94650 -4090 94850
rect -4020 94650 -3980 94850
rect -3910 94650 -3590 94850
rect -3520 94650 -3480 94850
rect -3410 94650 -3090 94850
rect -3020 94650 -2980 94850
rect -2910 94650 -2590 94850
rect -2520 94650 -2480 94850
rect -2410 94650 -2090 94850
rect -2020 94650 -1980 94850
rect -1910 94650 -1590 94850
rect -1520 94650 -1480 94850
rect -1410 94650 -1090 94850
rect -1020 94650 -980 94850
rect -910 94650 -590 94850
rect -520 94650 -480 94850
rect -410 94650 -90 94850
rect -20 94650 20 94850
rect 90 94650 410 94850
rect 480 94650 520 94850
rect 590 94650 910 94850
rect 980 94650 1020 94850
rect 1090 94650 1410 94850
rect 1480 94650 1520 94850
rect 1590 94650 1910 94850
rect 1980 94650 2020 94850
rect 2090 94650 2410 94850
rect 2480 94650 2520 94850
rect 2590 94650 2910 94850
rect 2980 94650 3020 94850
rect 3090 94650 3410 94850
rect 3480 94650 3520 94850
rect 3590 94650 3910 94850
rect 3980 94650 4020 94850
rect 4090 94650 4410 94850
rect 4480 94650 4520 94850
rect 4590 94650 4910 94850
rect 4980 94650 5020 94850
rect 5090 94650 5410 94850
rect 5480 94650 5520 94850
rect 5590 94650 5910 94850
rect 5980 94650 6020 94850
rect 6090 94650 6410 94850
rect 6480 94650 6520 94850
rect 6590 94650 6910 94850
rect 6980 94650 7020 94850
rect 7090 94650 7410 94850
rect 7480 94650 7520 94850
rect 7590 94650 7910 94850
rect 7980 94650 8020 94850
rect 8090 94650 8410 94850
rect 8480 94650 8520 94850
rect 8590 94650 8910 94850
rect 8980 94650 9020 94850
rect 9090 94650 9410 94850
rect 9480 94650 9520 94850
rect 9590 94650 9910 94850
rect 9980 94650 10020 94850
rect 10090 94650 10410 94850
rect 10480 94650 10520 94850
rect 10590 94650 10910 94850
rect 10980 94650 11020 94850
rect 11090 94650 11410 94850
rect 11480 94650 11520 94850
rect 11590 94650 11910 94850
rect 11980 94650 12020 94850
rect 12090 94650 12410 94850
rect 12480 94650 12520 94850
rect 12590 94650 12910 94850
rect 12980 94650 13020 94850
rect 13090 94650 13410 94850
rect 13480 94650 13520 94850
rect 13590 94650 13910 94850
rect 13980 94650 14020 94850
rect 14090 94650 14410 94850
rect 14480 94650 14520 94850
rect 14590 94650 14910 94850
rect 14980 94650 15020 94850
rect 15090 94650 15410 94850
rect 15480 94650 15520 94850
rect 15590 94650 15910 94850
rect 15980 94650 16020 94850
rect 16090 94650 16410 94850
rect 16480 94650 16520 94850
rect 16590 94650 16910 94850
rect 16980 94650 17020 94850
rect 17090 94650 17410 94850
rect 17480 94650 17520 94850
rect 17590 94650 17910 94850
rect 17980 94650 18020 94850
rect 18090 94650 18410 94850
rect 18480 94650 18520 94850
rect 18590 94650 18910 94850
rect 18980 94650 19020 94850
rect 19090 94650 19410 94850
rect 19480 94650 19520 94850
rect 19590 94650 19910 94850
rect 19980 94650 20000 94850
rect -16000 94640 20000 94650
rect -15860 94590 -15640 94640
rect -15860 94520 -15850 94590
rect -15650 94520 -15640 94590
rect -15860 94480 -15640 94520
rect -15860 94410 -15850 94480
rect -15650 94410 -15640 94480
rect -15860 94360 -15640 94410
rect -15360 94590 -15140 94640
rect -15360 94520 -15350 94590
rect -15150 94520 -15140 94590
rect -15360 94480 -15140 94520
rect -15360 94410 -15350 94480
rect -15150 94410 -15140 94480
rect -15360 94360 -15140 94410
rect -14860 94590 -14640 94640
rect -14860 94520 -14850 94590
rect -14650 94520 -14640 94590
rect -14860 94480 -14640 94520
rect -14860 94410 -14850 94480
rect -14650 94410 -14640 94480
rect -14860 94360 -14640 94410
rect -14360 94590 -14140 94640
rect -14360 94520 -14350 94590
rect -14150 94520 -14140 94590
rect -14360 94480 -14140 94520
rect -14360 94410 -14350 94480
rect -14150 94410 -14140 94480
rect -14360 94360 -14140 94410
rect -13860 94590 -13640 94640
rect -13860 94520 -13850 94590
rect -13650 94520 -13640 94590
rect -13860 94480 -13640 94520
rect -13860 94410 -13850 94480
rect -13650 94410 -13640 94480
rect -13860 94360 -13640 94410
rect -13360 94590 -13140 94640
rect -13360 94520 -13350 94590
rect -13150 94520 -13140 94590
rect -13360 94480 -13140 94520
rect -13360 94410 -13350 94480
rect -13150 94410 -13140 94480
rect -13360 94360 -13140 94410
rect -12860 94590 -12640 94640
rect -12860 94520 -12850 94590
rect -12650 94520 -12640 94590
rect -12860 94480 -12640 94520
rect -12860 94410 -12850 94480
rect -12650 94410 -12640 94480
rect -12860 94360 -12640 94410
rect -12360 94590 -12140 94640
rect -12360 94520 -12350 94590
rect -12150 94520 -12140 94590
rect -12360 94480 -12140 94520
rect -12360 94410 -12350 94480
rect -12150 94410 -12140 94480
rect -12360 94360 -12140 94410
rect -11860 94590 -11640 94640
rect -11860 94520 -11850 94590
rect -11650 94520 -11640 94590
rect -11860 94480 -11640 94520
rect -11860 94410 -11850 94480
rect -11650 94410 -11640 94480
rect -11860 94360 -11640 94410
rect -11360 94590 -11140 94640
rect -11360 94520 -11350 94590
rect -11150 94520 -11140 94590
rect -11360 94480 -11140 94520
rect -11360 94410 -11350 94480
rect -11150 94410 -11140 94480
rect -11360 94360 -11140 94410
rect -10860 94590 -10640 94640
rect -10860 94520 -10850 94590
rect -10650 94520 -10640 94590
rect -10860 94480 -10640 94520
rect -10860 94410 -10850 94480
rect -10650 94410 -10640 94480
rect -10860 94360 -10640 94410
rect -10360 94590 -10140 94640
rect -10360 94520 -10350 94590
rect -10150 94520 -10140 94590
rect -10360 94480 -10140 94520
rect -10360 94410 -10350 94480
rect -10150 94410 -10140 94480
rect -10360 94360 -10140 94410
rect -9860 94590 -9640 94640
rect -9860 94520 -9850 94590
rect -9650 94520 -9640 94590
rect -9860 94480 -9640 94520
rect -9860 94410 -9850 94480
rect -9650 94410 -9640 94480
rect -9860 94360 -9640 94410
rect -9360 94590 -9140 94640
rect -9360 94520 -9350 94590
rect -9150 94520 -9140 94590
rect -9360 94480 -9140 94520
rect -9360 94410 -9350 94480
rect -9150 94410 -9140 94480
rect -9360 94360 -9140 94410
rect -8860 94590 -8640 94640
rect -8860 94520 -8850 94590
rect -8650 94520 -8640 94590
rect -8860 94480 -8640 94520
rect -8860 94410 -8850 94480
rect -8650 94410 -8640 94480
rect -8860 94360 -8640 94410
rect -8360 94590 -8140 94640
rect -8360 94520 -8350 94590
rect -8150 94520 -8140 94590
rect -8360 94480 -8140 94520
rect -8360 94410 -8350 94480
rect -8150 94410 -8140 94480
rect -8360 94360 -8140 94410
rect -7860 94590 -7640 94640
rect -7860 94520 -7850 94590
rect -7650 94520 -7640 94590
rect -7860 94480 -7640 94520
rect -7860 94410 -7850 94480
rect -7650 94410 -7640 94480
rect -7860 94360 -7640 94410
rect -7360 94590 -7140 94640
rect -7360 94520 -7350 94590
rect -7150 94520 -7140 94590
rect -7360 94480 -7140 94520
rect -7360 94410 -7350 94480
rect -7150 94410 -7140 94480
rect -7360 94360 -7140 94410
rect -6860 94590 -6640 94640
rect -6860 94520 -6850 94590
rect -6650 94520 -6640 94590
rect -6860 94480 -6640 94520
rect -6860 94410 -6850 94480
rect -6650 94410 -6640 94480
rect -6860 94360 -6640 94410
rect -6360 94590 -6140 94640
rect -6360 94520 -6350 94590
rect -6150 94520 -6140 94590
rect -6360 94480 -6140 94520
rect -6360 94410 -6350 94480
rect -6150 94410 -6140 94480
rect -6360 94360 -6140 94410
rect -5860 94590 -5640 94640
rect -5860 94520 -5850 94590
rect -5650 94520 -5640 94590
rect -5860 94480 -5640 94520
rect -5860 94410 -5850 94480
rect -5650 94410 -5640 94480
rect -5860 94360 -5640 94410
rect -5360 94590 -5140 94640
rect -5360 94520 -5350 94590
rect -5150 94520 -5140 94590
rect -5360 94480 -5140 94520
rect -5360 94410 -5350 94480
rect -5150 94410 -5140 94480
rect -5360 94360 -5140 94410
rect -4860 94590 -4640 94640
rect -4860 94520 -4850 94590
rect -4650 94520 -4640 94590
rect -4860 94480 -4640 94520
rect -4860 94410 -4850 94480
rect -4650 94410 -4640 94480
rect -4860 94360 -4640 94410
rect -4360 94590 -4140 94640
rect -4360 94520 -4350 94590
rect -4150 94520 -4140 94590
rect -4360 94480 -4140 94520
rect -4360 94410 -4350 94480
rect -4150 94410 -4140 94480
rect -4360 94360 -4140 94410
rect -3860 94590 -3640 94640
rect -3860 94520 -3850 94590
rect -3650 94520 -3640 94590
rect -3860 94480 -3640 94520
rect -3860 94410 -3850 94480
rect -3650 94410 -3640 94480
rect -3860 94360 -3640 94410
rect -3360 94590 -3140 94640
rect -3360 94520 -3350 94590
rect -3150 94520 -3140 94590
rect -3360 94480 -3140 94520
rect -3360 94410 -3350 94480
rect -3150 94410 -3140 94480
rect -3360 94360 -3140 94410
rect -2860 94590 -2640 94640
rect -2860 94520 -2850 94590
rect -2650 94520 -2640 94590
rect -2860 94480 -2640 94520
rect -2860 94410 -2850 94480
rect -2650 94410 -2640 94480
rect -2860 94360 -2640 94410
rect -2360 94590 -2140 94640
rect -2360 94520 -2350 94590
rect -2150 94520 -2140 94590
rect -2360 94480 -2140 94520
rect -2360 94410 -2350 94480
rect -2150 94410 -2140 94480
rect -2360 94360 -2140 94410
rect -1860 94590 -1640 94640
rect -1860 94520 -1850 94590
rect -1650 94520 -1640 94590
rect -1860 94480 -1640 94520
rect -1860 94410 -1850 94480
rect -1650 94410 -1640 94480
rect -1860 94360 -1640 94410
rect -1360 94590 -1140 94640
rect -1360 94520 -1350 94590
rect -1150 94520 -1140 94590
rect -1360 94480 -1140 94520
rect -1360 94410 -1350 94480
rect -1150 94410 -1140 94480
rect -1360 94360 -1140 94410
rect -860 94590 -640 94640
rect -860 94520 -850 94590
rect -650 94520 -640 94590
rect -860 94480 -640 94520
rect -860 94410 -850 94480
rect -650 94410 -640 94480
rect -860 94360 -640 94410
rect -360 94590 -140 94640
rect -360 94520 -350 94590
rect -150 94520 -140 94590
rect -360 94480 -140 94520
rect -360 94410 -350 94480
rect -150 94410 -140 94480
rect -360 94360 -140 94410
rect 140 94590 360 94640
rect 140 94520 150 94590
rect 350 94520 360 94590
rect 140 94480 360 94520
rect 140 94410 150 94480
rect 350 94410 360 94480
rect 140 94360 360 94410
rect 640 94590 860 94640
rect 640 94520 650 94590
rect 850 94520 860 94590
rect 640 94480 860 94520
rect 640 94410 650 94480
rect 850 94410 860 94480
rect 640 94360 860 94410
rect 1140 94590 1360 94640
rect 1140 94520 1150 94590
rect 1350 94520 1360 94590
rect 1140 94480 1360 94520
rect 1140 94410 1150 94480
rect 1350 94410 1360 94480
rect 1140 94360 1360 94410
rect 1640 94590 1860 94640
rect 1640 94520 1650 94590
rect 1850 94520 1860 94590
rect 1640 94480 1860 94520
rect 1640 94410 1650 94480
rect 1850 94410 1860 94480
rect 1640 94360 1860 94410
rect 2140 94590 2360 94640
rect 2140 94520 2150 94590
rect 2350 94520 2360 94590
rect 2140 94480 2360 94520
rect 2140 94410 2150 94480
rect 2350 94410 2360 94480
rect 2140 94360 2360 94410
rect 2640 94590 2860 94640
rect 2640 94520 2650 94590
rect 2850 94520 2860 94590
rect 2640 94480 2860 94520
rect 2640 94410 2650 94480
rect 2850 94410 2860 94480
rect 2640 94360 2860 94410
rect 3140 94590 3360 94640
rect 3140 94520 3150 94590
rect 3350 94520 3360 94590
rect 3140 94480 3360 94520
rect 3140 94410 3150 94480
rect 3350 94410 3360 94480
rect 3140 94360 3360 94410
rect 3640 94590 3860 94640
rect 3640 94520 3650 94590
rect 3850 94520 3860 94590
rect 3640 94480 3860 94520
rect 3640 94410 3650 94480
rect 3850 94410 3860 94480
rect 3640 94360 3860 94410
rect 4140 94590 4360 94640
rect 4140 94520 4150 94590
rect 4350 94520 4360 94590
rect 4140 94480 4360 94520
rect 4140 94410 4150 94480
rect 4350 94410 4360 94480
rect 4140 94360 4360 94410
rect 4640 94590 4860 94640
rect 4640 94520 4650 94590
rect 4850 94520 4860 94590
rect 4640 94480 4860 94520
rect 4640 94410 4650 94480
rect 4850 94410 4860 94480
rect 4640 94360 4860 94410
rect 5140 94590 5360 94640
rect 5140 94520 5150 94590
rect 5350 94520 5360 94590
rect 5140 94480 5360 94520
rect 5140 94410 5150 94480
rect 5350 94410 5360 94480
rect 5140 94360 5360 94410
rect 5640 94590 5860 94640
rect 5640 94520 5650 94590
rect 5850 94520 5860 94590
rect 5640 94480 5860 94520
rect 5640 94410 5650 94480
rect 5850 94410 5860 94480
rect 5640 94360 5860 94410
rect 6140 94590 6360 94640
rect 6140 94520 6150 94590
rect 6350 94520 6360 94590
rect 6140 94480 6360 94520
rect 6140 94410 6150 94480
rect 6350 94410 6360 94480
rect 6140 94360 6360 94410
rect 6640 94590 6860 94640
rect 6640 94520 6650 94590
rect 6850 94520 6860 94590
rect 6640 94480 6860 94520
rect 6640 94410 6650 94480
rect 6850 94410 6860 94480
rect 6640 94360 6860 94410
rect 7140 94590 7360 94640
rect 7140 94520 7150 94590
rect 7350 94520 7360 94590
rect 7140 94480 7360 94520
rect 7140 94410 7150 94480
rect 7350 94410 7360 94480
rect 7140 94360 7360 94410
rect 7640 94590 7860 94640
rect 7640 94520 7650 94590
rect 7850 94520 7860 94590
rect 7640 94480 7860 94520
rect 7640 94410 7650 94480
rect 7850 94410 7860 94480
rect 7640 94360 7860 94410
rect 8140 94590 8360 94640
rect 8140 94520 8150 94590
rect 8350 94520 8360 94590
rect 8140 94480 8360 94520
rect 8140 94410 8150 94480
rect 8350 94410 8360 94480
rect 8140 94360 8360 94410
rect 8640 94590 8860 94640
rect 8640 94520 8650 94590
rect 8850 94520 8860 94590
rect 8640 94480 8860 94520
rect 8640 94410 8650 94480
rect 8850 94410 8860 94480
rect 8640 94360 8860 94410
rect 9140 94590 9360 94640
rect 9140 94520 9150 94590
rect 9350 94520 9360 94590
rect 9140 94480 9360 94520
rect 9140 94410 9150 94480
rect 9350 94410 9360 94480
rect 9140 94360 9360 94410
rect 9640 94590 9860 94640
rect 9640 94520 9650 94590
rect 9850 94520 9860 94590
rect 9640 94480 9860 94520
rect 9640 94410 9650 94480
rect 9850 94410 9860 94480
rect 9640 94360 9860 94410
rect 10140 94590 10360 94640
rect 10140 94520 10150 94590
rect 10350 94520 10360 94590
rect 10140 94480 10360 94520
rect 10140 94410 10150 94480
rect 10350 94410 10360 94480
rect 10140 94360 10360 94410
rect 10640 94590 10860 94640
rect 10640 94520 10650 94590
rect 10850 94520 10860 94590
rect 10640 94480 10860 94520
rect 10640 94410 10650 94480
rect 10850 94410 10860 94480
rect 10640 94360 10860 94410
rect 11140 94590 11360 94640
rect 11140 94520 11150 94590
rect 11350 94520 11360 94590
rect 11140 94480 11360 94520
rect 11140 94410 11150 94480
rect 11350 94410 11360 94480
rect 11140 94360 11360 94410
rect 11640 94590 11860 94640
rect 11640 94520 11650 94590
rect 11850 94520 11860 94590
rect 11640 94480 11860 94520
rect 11640 94410 11650 94480
rect 11850 94410 11860 94480
rect 11640 94360 11860 94410
rect 12140 94590 12360 94640
rect 12140 94520 12150 94590
rect 12350 94520 12360 94590
rect 12140 94480 12360 94520
rect 12140 94410 12150 94480
rect 12350 94410 12360 94480
rect 12140 94360 12360 94410
rect 12640 94590 12860 94640
rect 12640 94520 12650 94590
rect 12850 94520 12860 94590
rect 12640 94480 12860 94520
rect 12640 94410 12650 94480
rect 12850 94410 12860 94480
rect 12640 94360 12860 94410
rect 13140 94590 13360 94640
rect 13140 94520 13150 94590
rect 13350 94520 13360 94590
rect 13140 94480 13360 94520
rect 13140 94410 13150 94480
rect 13350 94410 13360 94480
rect 13140 94360 13360 94410
rect 13640 94590 13860 94640
rect 13640 94520 13650 94590
rect 13850 94520 13860 94590
rect 13640 94480 13860 94520
rect 13640 94410 13650 94480
rect 13850 94410 13860 94480
rect 13640 94360 13860 94410
rect 14140 94590 14360 94640
rect 14140 94520 14150 94590
rect 14350 94520 14360 94590
rect 14140 94480 14360 94520
rect 14140 94410 14150 94480
rect 14350 94410 14360 94480
rect 14140 94360 14360 94410
rect 14640 94590 14860 94640
rect 14640 94520 14650 94590
rect 14850 94520 14860 94590
rect 14640 94480 14860 94520
rect 14640 94410 14650 94480
rect 14850 94410 14860 94480
rect 14640 94360 14860 94410
rect 15140 94590 15360 94640
rect 15140 94520 15150 94590
rect 15350 94520 15360 94590
rect 15140 94480 15360 94520
rect 15140 94410 15150 94480
rect 15350 94410 15360 94480
rect 15140 94360 15360 94410
rect 15640 94590 15860 94640
rect 15640 94520 15650 94590
rect 15850 94520 15860 94590
rect 15640 94480 15860 94520
rect 15640 94410 15650 94480
rect 15850 94410 15860 94480
rect 15640 94360 15860 94410
rect 16140 94590 16360 94640
rect 16140 94520 16150 94590
rect 16350 94520 16360 94590
rect 16140 94480 16360 94520
rect 16140 94410 16150 94480
rect 16350 94410 16360 94480
rect 16140 94360 16360 94410
rect 16640 94590 16860 94640
rect 16640 94520 16650 94590
rect 16850 94520 16860 94590
rect 16640 94480 16860 94520
rect 16640 94410 16650 94480
rect 16850 94410 16860 94480
rect 16640 94360 16860 94410
rect 17140 94590 17360 94640
rect 17140 94520 17150 94590
rect 17350 94520 17360 94590
rect 17140 94480 17360 94520
rect 17140 94410 17150 94480
rect 17350 94410 17360 94480
rect 17140 94360 17360 94410
rect 17640 94590 17860 94640
rect 17640 94520 17650 94590
rect 17850 94520 17860 94590
rect 17640 94480 17860 94520
rect 17640 94410 17650 94480
rect 17850 94410 17860 94480
rect 17640 94360 17860 94410
rect 18140 94590 18360 94640
rect 18140 94520 18150 94590
rect 18350 94520 18360 94590
rect 18140 94480 18360 94520
rect 18140 94410 18150 94480
rect 18350 94410 18360 94480
rect 18140 94360 18360 94410
rect 18640 94590 18860 94640
rect 18640 94520 18650 94590
rect 18850 94520 18860 94590
rect 18640 94480 18860 94520
rect 18640 94410 18650 94480
rect 18850 94410 18860 94480
rect 18640 94360 18860 94410
rect 19140 94590 19360 94640
rect 19140 94520 19150 94590
rect 19350 94520 19360 94590
rect 19140 94480 19360 94520
rect 19140 94410 19150 94480
rect 19350 94410 19360 94480
rect 19140 94360 19360 94410
rect 19640 94590 19860 94640
rect 19640 94520 19650 94590
rect 19850 94520 19860 94590
rect 19640 94480 19860 94520
rect 19640 94410 19650 94480
rect 19850 94410 19860 94480
rect 19640 94360 19860 94410
rect -16000 94350 20000 94360
rect -16000 94150 -15980 94350
rect -15910 94150 -15590 94350
rect -15520 94150 -15480 94350
rect -15410 94150 -15090 94350
rect -15020 94150 -14980 94350
rect -14910 94150 -14590 94350
rect -14520 94150 -14480 94350
rect -14410 94150 -14090 94350
rect -14020 94150 -13980 94350
rect -13910 94150 -13590 94350
rect -13520 94150 -13480 94350
rect -13410 94150 -13090 94350
rect -13020 94150 -12980 94350
rect -12910 94150 -12590 94350
rect -12520 94150 -12480 94350
rect -12410 94150 -12090 94350
rect -12020 94150 -11980 94350
rect -11910 94150 -11590 94350
rect -11520 94150 -11480 94350
rect -11410 94150 -11090 94350
rect -11020 94150 -10980 94350
rect -10910 94150 -10590 94350
rect -10520 94150 -10480 94350
rect -10410 94150 -10090 94350
rect -10020 94150 -9980 94350
rect -9910 94150 -9590 94350
rect -9520 94150 -9480 94350
rect -9410 94150 -9090 94350
rect -9020 94150 -8980 94350
rect -8910 94150 -8590 94350
rect -8520 94150 -8480 94350
rect -8410 94150 -8090 94350
rect -8020 94150 -7980 94350
rect -7910 94150 -7590 94350
rect -7520 94150 -7480 94350
rect -7410 94150 -7090 94350
rect -7020 94150 -6980 94350
rect -6910 94150 -6590 94350
rect -6520 94150 -6480 94350
rect -6410 94150 -6090 94350
rect -6020 94150 -5980 94350
rect -5910 94150 -5590 94350
rect -5520 94150 -5480 94350
rect -5410 94150 -5090 94350
rect -5020 94150 -4980 94350
rect -4910 94150 -4590 94350
rect -4520 94150 -4480 94350
rect -4410 94150 -4090 94350
rect -4020 94150 -3980 94350
rect -3910 94150 -3590 94350
rect -3520 94150 -3480 94350
rect -3410 94150 -3090 94350
rect -3020 94150 -2980 94350
rect -2910 94150 -2590 94350
rect -2520 94150 -2480 94350
rect -2410 94150 -2090 94350
rect -2020 94150 -1980 94350
rect -1910 94150 -1590 94350
rect -1520 94150 -1480 94350
rect -1410 94150 -1090 94350
rect -1020 94150 -980 94350
rect -910 94150 -590 94350
rect -520 94150 -480 94350
rect -410 94150 -90 94350
rect -20 94150 20 94350
rect 90 94150 410 94350
rect 480 94150 520 94350
rect 590 94150 910 94350
rect 980 94150 1020 94350
rect 1090 94150 1410 94350
rect 1480 94150 1520 94350
rect 1590 94150 1910 94350
rect 1980 94150 2020 94350
rect 2090 94150 2410 94350
rect 2480 94150 2520 94350
rect 2590 94150 2910 94350
rect 2980 94150 3020 94350
rect 3090 94150 3410 94350
rect 3480 94150 3520 94350
rect 3590 94150 3910 94350
rect 3980 94150 4020 94350
rect 4090 94150 4410 94350
rect 4480 94150 4520 94350
rect 4590 94150 4910 94350
rect 4980 94150 5020 94350
rect 5090 94150 5410 94350
rect 5480 94150 5520 94350
rect 5590 94150 5910 94350
rect 5980 94150 6020 94350
rect 6090 94150 6410 94350
rect 6480 94150 6520 94350
rect 6590 94150 6910 94350
rect 6980 94150 7020 94350
rect 7090 94150 7410 94350
rect 7480 94150 7520 94350
rect 7590 94150 7910 94350
rect 7980 94150 8020 94350
rect 8090 94150 8410 94350
rect 8480 94150 8520 94350
rect 8590 94150 8910 94350
rect 8980 94150 9020 94350
rect 9090 94150 9410 94350
rect 9480 94150 9520 94350
rect 9590 94150 9910 94350
rect 9980 94150 10020 94350
rect 10090 94150 10410 94350
rect 10480 94150 10520 94350
rect 10590 94150 10910 94350
rect 10980 94150 11020 94350
rect 11090 94150 11410 94350
rect 11480 94150 11520 94350
rect 11590 94150 11910 94350
rect 11980 94150 12020 94350
rect 12090 94150 12410 94350
rect 12480 94150 12520 94350
rect 12590 94150 12910 94350
rect 12980 94150 13020 94350
rect 13090 94150 13410 94350
rect 13480 94150 13520 94350
rect 13590 94150 13910 94350
rect 13980 94150 14020 94350
rect 14090 94150 14410 94350
rect 14480 94150 14520 94350
rect 14590 94150 14910 94350
rect 14980 94150 15020 94350
rect 15090 94150 15410 94350
rect 15480 94150 15520 94350
rect 15590 94150 15910 94350
rect 15980 94150 16020 94350
rect 16090 94150 16410 94350
rect 16480 94150 16520 94350
rect 16590 94150 16910 94350
rect 16980 94150 17020 94350
rect 17090 94150 17410 94350
rect 17480 94150 17520 94350
rect 17590 94150 17910 94350
rect 17980 94150 18020 94350
rect 18090 94150 18410 94350
rect 18480 94150 18520 94350
rect 18590 94150 18910 94350
rect 18980 94150 19020 94350
rect 19090 94150 19410 94350
rect 19480 94150 19520 94350
rect 19590 94150 19910 94350
rect 19980 94150 20000 94350
rect -16000 94140 20000 94150
rect -15860 94090 -15640 94140
rect -15860 94020 -15850 94090
rect -15650 94020 -15640 94090
rect -15860 93980 -15640 94020
rect -15860 93910 -15850 93980
rect -15650 93910 -15640 93980
rect -15860 93860 -15640 93910
rect -15360 94090 -15140 94140
rect -15360 94020 -15350 94090
rect -15150 94020 -15140 94090
rect -15360 93980 -15140 94020
rect -15360 93910 -15350 93980
rect -15150 93910 -15140 93980
rect -15360 93860 -15140 93910
rect -14860 94090 -14640 94140
rect -14860 94020 -14850 94090
rect -14650 94020 -14640 94090
rect -14860 93980 -14640 94020
rect -14860 93910 -14850 93980
rect -14650 93910 -14640 93980
rect -14860 93860 -14640 93910
rect -14360 94090 -14140 94140
rect -14360 94020 -14350 94090
rect -14150 94020 -14140 94090
rect -14360 93980 -14140 94020
rect -14360 93910 -14350 93980
rect -14150 93910 -14140 93980
rect -14360 93860 -14140 93910
rect -13860 94090 -13640 94140
rect -13860 94020 -13850 94090
rect -13650 94020 -13640 94090
rect -13860 93980 -13640 94020
rect -13860 93910 -13850 93980
rect -13650 93910 -13640 93980
rect -13860 93860 -13640 93910
rect -13360 94090 -13140 94140
rect -13360 94020 -13350 94090
rect -13150 94020 -13140 94090
rect -13360 93980 -13140 94020
rect -13360 93910 -13350 93980
rect -13150 93910 -13140 93980
rect -13360 93860 -13140 93910
rect -12860 94090 -12640 94140
rect -12860 94020 -12850 94090
rect -12650 94020 -12640 94090
rect -12860 93980 -12640 94020
rect -12860 93910 -12850 93980
rect -12650 93910 -12640 93980
rect -12860 93860 -12640 93910
rect -12360 94090 -12140 94140
rect -12360 94020 -12350 94090
rect -12150 94020 -12140 94090
rect -12360 93980 -12140 94020
rect -11860 94090 -11640 94140
rect -11860 94020 -11850 94090
rect -11650 94020 -11640 94090
rect -11860 94000 -11640 94020
rect -11360 94090 -11140 94140
rect -11360 94020 -11350 94090
rect -11150 94020 -11140 94090
rect -11360 94000 -11140 94020
rect -10860 94090 -10640 94140
rect -10860 94020 -10850 94090
rect -10650 94020 -10640 94090
rect -10860 94000 -10640 94020
rect -10360 94090 -10140 94140
rect -10360 94020 -10350 94090
rect -10150 94020 -10140 94090
rect -10360 94000 -10140 94020
rect -9860 94090 -9640 94140
rect -9860 94020 -9850 94090
rect -9650 94020 -9640 94090
rect -9860 94000 -9640 94020
rect -9360 94090 -9140 94140
rect -9360 94020 -9350 94090
rect -9150 94020 -9140 94090
rect -9360 94000 -9140 94020
rect -8860 94090 -8640 94140
rect -8860 94020 -8850 94090
rect -8650 94020 -8640 94090
rect -8860 94000 -8640 94020
rect -8360 94090 -8140 94140
rect -8360 94020 -8350 94090
rect -8150 94020 -8140 94090
rect -8360 94000 -8140 94020
rect -7860 94090 -7640 94140
rect -7860 94020 -7850 94090
rect -7650 94020 -7640 94090
rect -7860 94000 -7640 94020
rect -7360 94090 -7140 94140
rect -7360 94020 -7350 94090
rect -7150 94020 -7140 94090
rect -7360 94000 -7140 94020
rect -6860 94090 -6640 94140
rect -6860 94020 -6850 94090
rect -6650 94020 -6640 94090
rect -6860 94000 -6640 94020
rect -6360 94090 -6140 94140
rect -6360 94020 -6350 94090
rect -6150 94020 -6140 94090
rect -6360 94000 -6140 94020
rect -5860 94090 -5640 94140
rect -5860 94020 -5850 94090
rect -5650 94020 -5640 94090
rect -5860 94000 -5640 94020
rect -5360 94090 -5140 94140
rect -5360 94020 -5350 94090
rect -5150 94020 -5140 94090
rect -5360 94000 -5140 94020
rect -4860 94090 -4640 94140
rect -4860 94020 -4850 94090
rect -4650 94020 -4640 94090
rect -4860 94000 -4640 94020
rect -4360 94090 -4140 94140
rect -4360 94020 -4350 94090
rect -4150 94020 -4140 94090
rect -4360 94000 -4140 94020
rect -3860 94090 -3640 94140
rect -3860 94020 -3850 94090
rect -3650 94020 -3640 94090
rect -3860 94000 -3640 94020
rect -3360 94090 -3140 94140
rect -3360 94020 -3350 94090
rect -3150 94020 -3140 94090
rect -3360 94000 -3140 94020
rect -2860 94090 -2640 94140
rect -2860 94020 -2850 94090
rect -2650 94020 -2640 94090
rect -2860 94000 -2640 94020
rect -2360 94090 -2140 94140
rect -2360 94020 -2350 94090
rect -2150 94020 -2140 94090
rect -2360 94000 -2140 94020
rect -1860 94090 -1640 94140
rect -1860 94020 -1850 94090
rect -1650 94020 -1640 94090
rect -1860 94000 -1640 94020
rect -1360 94090 -1140 94140
rect -1360 94020 -1350 94090
rect -1150 94020 -1140 94090
rect -1360 94000 -1140 94020
rect -860 94090 -640 94140
rect -860 94020 -850 94090
rect -650 94020 -640 94090
rect -860 94000 -640 94020
rect -360 94090 -140 94140
rect -360 94020 -350 94090
rect -150 94020 -140 94090
rect -360 94000 -140 94020
rect 140 94090 360 94140
rect 140 94020 150 94090
rect 350 94020 360 94090
rect 140 94000 360 94020
rect 640 94090 860 94140
rect 640 94020 650 94090
rect 850 94020 860 94090
rect 640 94000 860 94020
rect 1140 94090 1360 94140
rect 1140 94020 1150 94090
rect 1350 94020 1360 94090
rect 1140 94000 1360 94020
rect 1640 94090 1860 94140
rect 1640 94020 1650 94090
rect 1850 94020 1860 94090
rect 1640 94000 1860 94020
rect 2140 94090 2360 94140
rect 2140 94020 2150 94090
rect 2350 94020 2360 94090
rect 2140 94000 2360 94020
rect 2640 94090 2860 94140
rect 2640 94020 2650 94090
rect 2850 94020 2860 94090
rect 2640 94000 2860 94020
rect 3140 94090 3360 94140
rect 3140 94020 3150 94090
rect 3350 94020 3360 94090
rect 3140 94000 3360 94020
rect 3640 94090 3860 94140
rect 3640 94020 3650 94090
rect 3850 94020 3860 94090
rect 3640 94000 3860 94020
rect 4140 94090 4360 94140
rect 4140 94020 4150 94090
rect 4350 94020 4360 94090
rect 4140 94000 4360 94020
rect 4640 94090 4860 94140
rect 4640 94020 4650 94090
rect 4850 94020 4860 94090
rect 4640 94000 4860 94020
rect 5140 94090 5360 94140
rect 5140 94020 5150 94090
rect 5350 94020 5360 94090
rect 5140 94000 5360 94020
rect 5640 94090 5860 94140
rect 5640 94020 5650 94090
rect 5850 94020 5860 94090
rect 5640 94000 5860 94020
rect 6140 94090 6360 94140
rect 6140 94020 6150 94090
rect 6350 94020 6360 94090
rect 6140 94000 6360 94020
rect 6640 94090 6860 94140
rect 6640 94020 6650 94090
rect 6850 94020 6860 94090
rect 6640 94000 6860 94020
rect 7140 94090 7360 94140
rect 7140 94020 7150 94090
rect 7350 94020 7360 94090
rect 7140 94000 7360 94020
rect 7640 94090 7860 94140
rect 7640 94020 7650 94090
rect 7850 94020 7860 94090
rect 7640 94000 7860 94020
rect 8140 94090 8360 94140
rect 8140 94020 8150 94090
rect 8350 94020 8360 94090
rect 8140 94000 8360 94020
rect 8640 94090 8860 94140
rect 8640 94020 8650 94090
rect 8850 94020 8860 94090
rect 8640 94000 8860 94020
rect 9140 94090 9360 94140
rect 9140 94020 9150 94090
rect 9350 94020 9360 94090
rect 9140 94000 9360 94020
rect 9640 94090 9860 94140
rect 9640 94020 9650 94090
rect 9850 94020 9860 94090
rect 9640 94000 9860 94020
rect 10140 94090 10360 94140
rect 10140 94020 10150 94090
rect 10350 94020 10360 94090
rect 10140 94000 10360 94020
rect 10640 94090 10860 94140
rect 10640 94020 10650 94090
rect 10850 94020 10860 94090
rect 10640 94000 10860 94020
rect 11140 94090 11360 94140
rect 11140 94020 11150 94090
rect 11350 94020 11360 94090
rect 11140 94000 11360 94020
rect 11640 94090 11860 94140
rect 11640 94020 11650 94090
rect 11850 94020 11860 94090
rect 11640 94000 11860 94020
rect 12140 94090 12360 94140
rect 12140 94020 12150 94090
rect 12350 94020 12360 94090
rect 12140 94000 12360 94020
rect 12640 94090 12860 94140
rect 12640 94020 12650 94090
rect 12850 94020 12860 94090
rect 12640 94000 12860 94020
rect 13140 94090 13360 94140
rect 13140 94020 13150 94090
rect 13350 94020 13360 94090
rect 13140 94000 13360 94020
rect 13640 94090 13860 94140
rect 13640 94020 13650 94090
rect 13850 94020 13860 94090
rect 13640 94000 13860 94020
rect 14140 94090 14360 94140
rect 14140 94020 14150 94090
rect 14350 94020 14360 94090
rect 14140 94000 14360 94020
rect 14640 94090 14860 94140
rect 14640 94020 14650 94090
rect 14850 94020 14860 94090
rect 14640 94000 14860 94020
rect 15140 94090 15360 94140
rect 15140 94020 15150 94090
rect 15350 94020 15360 94090
rect 15140 94000 15360 94020
rect 15640 94090 15860 94140
rect 15640 94020 15650 94090
rect 15850 94020 15860 94090
rect 15640 94000 15860 94020
rect 16140 94090 16360 94140
rect 16140 94020 16150 94090
rect 16350 94020 16360 94090
rect 16140 94000 16360 94020
rect 16640 94090 16860 94140
rect 16640 94020 16650 94090
rect 16850 94020 16860 94090
rect 16640 94000 16860 94020
rect 17140 94090 17360 94140
rect 17140 94020 17150 94090
rect 17350 94020 17360 94090
rect 17140 94000 17360 94020
rect 17640 94090 17860 94140
rect 17640 94020 17650 94090
rect 17850 94020 17860 94090
rect 17640 94000 17860 94020
rect 18140 94090 18360 94140
rect 18140 94020 18150 94090
rect 18350 94020 18360 94090
rect 18140 94000 18360 94020
rect 18640 94090 18860 94140
rect 18640 94020 18650 94090
rect 18850 94020 18860 94090
rect 18640 94000 18860 94020
rect 19140 94090 19360 94140
rect 19140 94020 19150 94090
rect 19350 94020 19360 94090
rect 19140 94000 19360 94020
rect 19640 94090 19860 94140
rect 19640 94020 19650 94090
rect 19850 94020 19860 94090
rect 19640 94000 19860 94020
rect -12360 93910 -12350 93980
rect -12150 93910 -12140 93980
rect -12360 93860 -12140 93910
rect -16000 93850 -12000 93860
rect -16000 93650 -15980 93850
rect -15910 93650 -15590 93850
rect -15520 93650 -15480 93850
rect -15410 93650 -15090 93850
rect -15020 93650 -14980 93850
rect -14910 93650 -14590 93850
rect -14520 93650 -14480 93850
rect -14410 93650 -14090 93850
rect -14020 93650 -13980 93850
rect -13910 93650 -13590 93850
rect -13520 93650 -13480 93850
rect -13410 93650 -13090 93850
rect -13020 93650 -12980 93850
rect -12910 93650 -12590 93850
rect -12520 93650 -12480 93850
rect -12410 93650 -12090 93850
rect -12020 93650 -12000 93850
rect -16000 93640 -12000 93650
rect -15860 93590 -15640 93640
rect -15860 93520 -15850 93590
rect -15650 93520 -15640 93590
rect -15860 93480 -15640 93520
rect -15860 93410 -15850 93480
rect -15650 93410 -15640 93480
rect -15860 93360 -15640 93410
rect -15360 93590 -15140 93640
rect -15360 93520 -15350 93590
rect -15150 93520 -15140 93590
rect -15360 93480 -15140 93520
rect -15360 93410 -15350 93480
rect -15150 93410 -15140 93480
rect -15360 93360 -15140 93410
rect -14860 93590 -14640 93640
rect -14860 93520 -14850 93590
rect -14650 93520 -14640 93590
rect -14860 93480 -14640 93520
rect -14860 93410 -14850 93480
rect -14650 93410 -14640 93480
rect -14860 93360 -14640 93410
rect -14360 93590 -14140 93640
rect -14360 93520 -14350 93590
rect -14150 93520 -14140 93590
rect -14360 93480 -14140 93520
rect -14360 93410 -14350 93480
rect -14150 93410 -14140 93480
rect -14360 93360 -14140 93410
rect -13860 93590 -13640 93640
rect -13860 93520 -13850 93590
rect -13650 93520 -13640 93590
rect -13860 93480 -13640 93520
rect -13860 93410 -13850 93480
rect -13650 93410 -13640 93480
rect -13860 93360 -13640 93410
rect -13360 93590 -13140 93640
rect -13360 93520 -13350 93590
rect -13150 93520 -13140 93590
rect -13360 93480 -13140 93520
rect -13360 93410 -13350 93480
rect -13150 93410 -13140 93480
rect -13360 93360 -13140 93410
rect -12860 93590 -12640 93640
rect -12860 93520 -12850 93590
rect -12650 93520 -12640 93590
rect -12860 93480 -12640 93520
rect -12860 93410 -12850 93480
rect -12650 93410 -12640 93480
rect -12860 93360 -12640 93410
rect -12360 93590 -12140 93640
rect -12360 93520 -12350 93590
rect -12150 93520 -12140 93590
rect -12360 93480 -12140 93520
rect -12360 93410 -12350 93480
rect -12150 93410 -12140 93480
rect -12360 93360 -12140 93410
rect -16000 93350 -12000 93360
rect -16000 93150 -15980 93350
rect -15910 93150 -15590 93350
rect -15520 93150 -15480 93350
rect -15410 93150 -15090 93350
rect -15020 93150 -14980 93350
rect -14910 93150 -14590 93350
rect -14520 93150 -14480 93350
rect -14410 93150 -14090 93350
rect -14020 93150 -13980 93350
rect -13910 93150 -13590 93350
rect -13520 93150 -13480 93350
rect -13410 93150 -13090 93350
rect -13020 93150 -12980 93350
rect -12910 93150 -12590 93350
rect -12520 93150 -12480 93350
rect -12410 93150 -12090 93350
rect -12020 93150 -12000 93350
rect -16000 93140 -12000 93150
rect -15860 93090 -15640 93140
rect -15860 93020 -15850 93090
rect -15650 93020 -15640 93090
rect -15860 92980 -15640 93020
rect -15860 92910 -15850 92980
rect -15650 92910 -15640 92980
rect -15860 92860 -15640 92910
rect -15360 93090 -15140 93140
rect -15360 93020 -15350 93090
rect -15150 93020 -15140 93090
rect -15360 92980 -15140 93020
rect -15360 92910 -15350 92980
rect -15150 92910 -15140 92980
rect -15360 92860 -15140 92910
rect -14860 93090 -14640 93140
rect -14860 93020 -14850 93090
rect -14650 93020 -14640 93090
rect -14860 92980 -14640 93020
rect -14860 92910 -14850 92980
rect -14650 92910 -14640 92980
rect -14860 92860 -14640 92910
rect -14360 93090 -14140 93140
rect -14360 93020 -14350 93090
rect -14150 93020 -14140 93090
rect -14360 92980 -14140 93020
rect -14360 92910 -14350 92980
rect -14150 92910 -14140 92980
rect -14360 92860 -14140 92910
rect -13860 93090 -13640 93140
rect -13860 93020 -13850 93090
rect -13650 93020 -13640 93090
rect -13860 92980 -13640 93020
rect -13860 92910 -13850 92980
rect -13650 92910 -13640 92980
rect -13860 92860 -13640 92910
rect -13360 93090 -13140 93140
rect -13360 93020 -13350 93090
rect -13150 93020 -13140 93090
rect -13360 92980 -13140 93020
rect -13360 92910 -13350 92980
rect -13150 92910 -13140 92980
rect -13360 92860 -13140 92910
rect -12860 93090 -12640 93140
rect -12860 93020 -12850 93090
rect -12650 93020 -12640 93090
rect -12860 92980 -12640 93020
rect -12860 92910 -12850 92980
rect -12650 92910 -12640 92980
rect -12860 92860 -12640 92910
rect -12360 93090 -12140 93140
rect -12360 93020 -12350 93090
rect -12150 93020 -12140 93090
rect -12360 92980 -12140 93020
rect -12360 92910 -12350 92980
rect -12150 92910 -12140 92980
rect -12360 92860 -12140 92910
rect -16000 92850 -12000 92860
rect -16000 92650 -15980 92850
rect -15910 92650 -15590 92850
rect -15520 92650 -15480 92850
rect -15410 92650 -15090 92850
rect -15020 92650 -14980 92850
rect -14910 92650 -14590 92850
rect -14520 92650 -14480 92850
rect -14410 92650 -14090 92850
rect -14020 92650 -13980 92850
rect -13910 92650 -13590 92850
rect -13520 92650 -13480 92850
rect -13410 92650 -13090 92850
rect -13020 92650 -12980 92850
rect -12910 92650 -12590 92850
rect -12520 92650 -12480 92850
rect -12410 92650 -12090 92850
rect -12020 92650 -12000 92850
rect -16000 92640 -12000 92650
rect -15860 92590 -15640 92640
rect -15860 92520 -15850 92590
rect -15650 92520 -15640 92590
rect -15860 92480 -15640 92520
rect -15860 92410 -15850 92480
rect -15650 92410 -15640 92480
rect -15860 92360 -15640 92410
rect -15360 92590 -15140 92640
rect -15360 92520 -15350 92590
rect -15150 92520 -15140 92590
rect -15360 92480 -15140 92520
rect -15360 92410 -15350 92480
rect -15150 92410 -15140 92480
rect -15360 92360 -15140 92410
rect -14860 92590 -14640 92640
rect -14860 92520 -14850 92590
rect -14650 92520 -14640 92590
rect -14860 92480 -14640 92520
rect -14860 92410 -14850 92480
rect -14650 92410 -14640 92480
rect -14860 92360 -14640 92410
rect -14360 92590 -14140 92640
rect -14360 92520 -14350 92590
rect -14150 92520 -14140 92590
rect -14360 92480 -14140 92520
rect -14360 92410 -14350 92480
rect -14150 92410 -14140 92480
rect -14360 92360 -14140 92410
rect -13860 92590 -13640 92640
rect -13860 92520 -13850 92590
rect -13650 92520 -13640 92590
rect -13860 92480 -13640 92520
rect -13860 92410 -13850 92480
rect -13650 92410 -13640 92480
rect -13860 92360 -13640 92410
rect -13360 92590 -13140 92640
rect -13360 92520 -13350 92590
rect -13150 92520 -13140 92590
rect -13360 92480 -13140 92520
rect -13360 92410 -13350 92480
rect -13150 92410 -13140 92480
rect -13360 92360 -13140 92410
rect -12860 92590 -12640 92640
rect -12860 92520 -12850 92590
rect -12650 92520 -12640 92590
rect -12860 92480 -12640 92520
rect -12860 92410 -12850 92480
rect -12650 92410 -12640 92480
rect -12860 92360 -12640 92410
rect -12360 92590 -12140 92640
rect -12360 92520 -12350 92590
rect -12150 92520 -12140 92590
rect -12360 92480 -12140 92520
rect -12360 92410 -12350 92480
rect -12150 92410 -12140 92480
rect -12360 92360 -12140 92410
rect -16000 92350 -12000 92360
rect -16000 92150 -15980 92350
rect -15910 92150 -15590 92350
rect -15520 92150 -15480 92350
rect -15410 92150 -15090 92350
rect -15020 92150 -14980 92350
rect -14910 92150 -14590 92350
rect -14520 92150 -14480 92350
rect -14410 92150 -14090 92350
rect -14020 92150 -13980 92350
rect -13910 92150 -13590 92350
rect -13520 92150 -13480 92350
rect -13410 92150 -13090 92350
rect -13020 92150 -12980 92350
rect -12910 92150 -12590 92350
rect -12520 92150 -12480 92350
rect -12410 92150 -12090 92350
rect -12020 92150 -12000 92350
rect -16000 92140 -12000 92150
rect -15860 92090 -15640 92140
rect -15860 92020 -15850 92090
rect -15650 92020 -15640 92090
rect -15860 91980 -15640 92020
rect -15860 91910 -15850 91980
rect -15650 91910 -15640 91980
rect -15860 91860 -15640 91910
rect -15360 92090 -15140 92140
rect -15360 92020 -15350 92090
rect -15150 92020 -15140 92090
rect -15360 91980 -15140 92020
rect -15360 91910 -15350 91980
rect -15150 91910 -15140 91980
rect -15360 91860 -15140 91910
rect -14860 92090 -14640 92140
rect -14860 92020 -14850 92090
rect -14650 92020 -14640 92090
rect -14860 91980 -14640 92020
rect -14860 91910 -14850 91980
rect -14650 91910 -14640 91980
rect -14860 91860 -14640 91910
rect -14360 92090 -14140 92140
rect -14360 92020 -14350 92090
rect -14150 92020 -14140 92090
rect -14360 91980 -14140 92020
rect -14360 91910 -14350 91980
rect -14150 91910 -14140 91980
rect -14360 91860 -14140 91910
rect -13860 92090 -13640 92140
rect -13860 92020 -13850 92090
rect -13650 92020 -13640 92090
rect -13860 91980 -13640 92020
rect -13860 91910 -13850 91980
rect -13650 91910 -13640 91980
rect -13860 91860 -13640 91910
rect -13360 92090 -13140 92140
rect -13360 92020 -13350 92090
rect -13150 92020 -13140 92090
rect -13360 91980 -13140 92020
rect -13360 91910 -13350 91980
rect -13150 91910 -13140 91980
rect -13360 91860 -13140 91910
rect -12860 92090 -12640 92140
rect -12860 92020 -12850 92090
rect -12650 92020 -12640 92090
rect -12860 91980 -12640 92020
rect -12860 91910 -12850 91980
rect -12650 91910 -12640 91980
rect -12860 91860 -12640 91910
rect -12360 92090 -12140 92140
rect -12360 92020 -12350 92090
rect -12150 92020 -12140 92090
rect -12360 91980 -12140 92020
rect -12360 91910 -12350 91980
rect -12150 91910 -12140 91980
rect -12360 91860 -12140 91910
rect -16000 91850 -12000 91860
rect -16000 91650 -15980 91850
rect -15910 91650 -15590 91850
rect -15520 91650 -15480 91850
rect -15410 91650 -15090 91850
rect -15020 91650 -14980 91850
rect -14910 91650 -14590 91850
rect -14520 91650 -14480 91850
rect -14410 91650 -14090 91850
rect -14020 91650 -13980 91850
rect -13910 91650 -13590 91850
rect -13520 91650 -13480 91850
rect -13410 91650 -13090 91850
rect -13020 91650 -12980 91850
rect -12910 91650 -12590 91850
rect -12520 91650 -12480 91850
rect -12410 91650 -12090 91850
rect -12020 91650 -12000 91850
rect -16000 91640 -12000 91650
rect -15860 91590 -15640 91640
rect -15860 91520 -15850 91590
rect -15650 91520 -15640 91590
rect -15860 91480 -15640 91520
rect -15860 91410 -15850 91480
rect -15650 91410 -15640 91480
rect -15860 91360 -15640 91410
rect -15360 91590 -15140 91640
rect -15360 91520 -15350 91590
rect -15150 91520 -15140 91590
rect -15360 91480 -15140 91520
rect -15360 91410 -15350 91480
rect -15150 91410 -15140 91480
rect -15360 91360 -15140 91410
rect -14860 91590 -14640 91640
rect -14860 91520 -14850 91590
rect -14650 91520 -14640 91590
rect -14860 91480 -14640 91520
rect -14860 91410 -14850 91480
rect -14650 91410 -14640 91480
rect -14860 91360 -14640 91410
rect -14360 91590 -14140 91640
rect -14360 91520 -14350 91590
rect -14150 91520 -14140 91590
rect -14360 91480 -14140 91520
rect -14360 91410 -14350 91480
rect -14150 91410 -14140 91480
rect -14360 91360 -14140 91410
rect -13860 91590 -13640 91640
rect -13860 91520 -13850 91590
rect -13650 91520 -13640 91590
rect -13860 91480 -13640 91520
rect -13860 91410 -13850 91480
rect -13650 91410 -13640 91480
rect -13860 91360 -13640 91410
rect -13360 91590 -13140 91640
rect -13360 91520 -13350 91590
rect -13150 91520 -13140 91590
rect -13360 91480 -13140 91520
rect -13360 91410 -13350 91480
rect -13150 91410 -13140 91480
rect -13360 91360 -13140 91410
rect -12860 91590 -12640 91640
rect -12860 91520 -12850 91590
rect -12650 91520 -12640 91590
rect -12860 91480 -12640 91520
rect -12860 91410 -12850 91480
rect -12650 91410 -12640 91480
rect -12860 91360 -12640 91410
rect -12360 91590 -12140 91640
rect -12360 91520 -12350 91590
rect -12150 91520 -12140 91590
rect -12360 91480 -12140 91520
rect -12360 91410 -12350 91480
rect -12150 91410 -12140 91480
rect -12360 91360 -12140 91410
rect -16000 91350 -12000 91360
rect -16000 91150 -15980 91350
rect -15910 91150 -15590 91350
rect -15520 91150 -15480 91350
rect -15410 91150 -15090 91350
rect -15020 91150 -14980 91350
rect -14910 91150 -14590 91350
rect -14520 91150 -14480 91350
rect -14410 91150 -14090 91350
rect -14020 91150 -13980 91350
rect -13910 91150 -13590 91350
rect -13520 91150 -13480 91350
rect -13410 91150 -13090 91350
rect -13020 91150 -12980 91350
rect -12910 91150 -12590 91350
rect -12520 91150 -12480 91350
rect -12410 91150 -12090 91350
rect -12020 91150 -12000 91350
rect -16000 91140 -12000 91150
rect -15860 91090 -15640 91140
rect -15860 91020 -15850 91090
rect -15650 91020 -15640 91090
rect -15860 90980 -15640 91020
rect -15860 90910 -15850 90980
rect -15650 90910 -15640 90980
rect -15860 90860 -15640 90910
rect -15360 91090 -15140 91140
rect -15360 91020 -15350 91090
rect -15150 91020 -15140 91090
rect -15360 90980 -15140 91020
rect -15360 90910 -15350 90980
rect -15150 90910 -15140 90980
rect -15360 90860 -15140 90910
rect -14860 91090 -14640 91140
rect -14860 91020 -14850 91090
rect -14650 91020 -14640 91090
rect -14860 90980 -14640 91020
rect -14860 90910 -14850 90980
rect -14650 90910 -14640 90980
rect -14860 90860 -14640 90910
rect -14360 91090 -14140 91140
rect -14360 91020 -14350 91090
rect -14150 91020 -14140 91090
rect -14360 90980 -14140 91020
rect -14360 90910 -14350 90980
rect -14150 90910 -14140 90980
rect -14360 90860 -14140 90910
rect -13860 91090 -13640 91140
rect -13860 91020 -13850 91090
rect -13650 91020 -13640 91090
rect -13860 90980 -13640 91020
rect -13860 90910 -13850 90980
rect -13650 90910 -13640 90980
rect -13860 90860 -13640 90910
rect -13360 91090 -13140 91140
rect -13360 91020 -13350 91090
rect -13150 91020 -13140 91090
rect -13360 90980 -13140 91020
rect -13360 90910 -13350 90980
rect -13150 90910 -13140 90980
rect -13360 90860 -13140 90910
rect -12860 91090 -12640 91140
rect -12860 91020 -12850 91090
rect -12650 91020 -12640 91090
rect -12860 90980 -12640 91020
rect -12860 90910 -12850 90980
rect -12650 90910 -12640 90980
rect -12860 90860 -12640 90910
rect -12360 91090 -12140 91140
rect -12360 91020 -12350 91090
rect -12150 91020 -12140 91090
rect -12360 90980 -12140 91020
rect -12360 90910 -12350 90980
rect -12150 90910 -12140 90980
rect -12360 90860 -12140 90910
rect -16000 90850 -12000 90860
rect -16000 90650 -15980 90850
rect -15910 90650 -15590 90850
rect -15520 90650 -15480 90850
rect -15410 90650 -15090 90850
rect -15020 90650 -14980 90850
rect -14910 90650 -14590 90850
rect -14520 90650 -14480 90850
rect -14410 90650 -14090 90850
rect -14020 90650 -13980 90850
rect -13910 90650 -13590 90850
rect -13520 90650 -13480 90850
rect -13410 90650 -13090 90850
rect -13020 90650 -12980 90850
rect -12910 90650 -12590 90850
rect -12520 90650 -12480 90850
rect -12410 90650 -12090 90850
rect -12020 90650 -12000 90850
rect -16000 90640 -12000 90650
rect -15860 90590 -15640 90640
rect -15860 90520 -15850 90590
rect -15650 90520 -15640 90590
rect -15860 90480 -15640 90520
rect -15860 90410 -15850 90480
rect -15650 90410 -15640 90480
rect -15860 90360 -15640 90410
rect -15360 90590 -15140 90640
rect -15360 90520 -15350 90590
rect -15150 90520 -15140 90590
rect -15360 90480 -15140 90520
rect -15360 90410 -15350 90480
rect -15150 90410 -15140 90480
rect -15360 90360 -15140 90410
rect -14860 90590 -14640 90640
rect -14860 90520 -14850 90590
rect -14650 90520 -14640 90590
rect -14860 90480 -14640 90520
rect -14860 90410 -14850 90480
rect -14650 90410 -14640 90480
rect -14860 90360 -14640 90410
rect -14360 90590 -14140 90640
rect -14360 90520 -14350 90590
rect -14150 90520 -14140 90590
rect -14360 90480 -14140 90520
rect -14360 90410 -14350 90480
rect -14150 90410 -14140 90480
rect -14360 90360 -14140 90410
rect -13860 90590 -13640 90640
rect -13860 90520 -13850 90590
rect -13650 90520 -13640 90590
rect -13860 90480 -13640 90520
rect -13860 90410 -13850 90480
rect -13650 90410 -13640 90480
rect -13860 90360 -13640 90410
rect -13360 90590 -13140 90640
rect -13360 90520 -13350 90590
rect -13150 90520 -13140 90590
rect -13360 90480 -13140 90520
rect -13360 90410 -13350 90480
rect -13150 90410 -13140 90480
rect -13360 90360 -13140 90410
rect -12860 90590 -12640 90640
rect -12860 90520 -12850 90590
rect -12650 90520 -12640 90590
rect -12860 90480 -12640 90520
rect -12860 90410 -12850 90480
rect -12650 90410 -12640 90480
rect -12860 90360 -12640 90410
rect -12360 90590 -12140 90640
rect -12360 90520 -12350 90590
rect -12150 90520 -12140 90590
rect -12360 90480 -12140 90520
rect -12360 90410 -12350 90480
rect -12150 90410 -12140 90480
rect -12360 90360 -12140 90410
rect -16000 90350 -12000 90360
rect -16000 90150 -15980 90350
rect -15910 90150 -15590 90350
rect -15520 90150 -15480 90350
rect -15410 90150 -15090 90350
rect -15020 90150 -14980 90350
rect -14910 90150 -14590 90350
rect -14520 90150 -14480 90350
rect -14410 90150 -14090 90350
rect -14020 90150 -13980 90350
rect -13910 90150 -13590 90350
rect -13520 90150 -13480 90350
rect -13410 90150 -13090 90350
rect -13020 90150 -12980 90350
rect -12910 90150 -12590 90350
rect -12520 90150 -12480 90350
rect -12410 90150 -12090 90350
rect -12020 90150 -12000 90350
rect -16000 90140 -12000 90150
rect -15860 90090 -15640 90140
rect -15860 90020 -15850 90090
rect -15650 90020 -15640 90090
rect -15860 89980 -15640 90020
rect -15860 89910 -15850 89980
rect -15650 89910 -15640 89980
rect -15860 89860 -15640 89910
rect -15360 90090 -15140 90140
rect -15360 90020 -15350 90090
rect -15150 90020 -15140 90090
rect -15360 89980 -15140 90020
rect -15360 89910 -15350 89980
rect -15150 89910 -15140 89980
rect -15360 89860 -15140 89910
rect -14860 90090 -14640 90140
rect -14860 90020 -14850 90090
rect -14650 90020 -14640 90090
rect -14860 89980 -14640 90020
rect -14860 89910 -14850 89980
rect -14650 89910 -14640 89980
rect -14860 89860 -14640 89910
rect -14360 90090 -14140 90140
rect -14360 90020 -14350 90090
rect -14150 90020 -14140 90090
rect -14360 89980 -14140 90020
rect -14360 89910 -14350 89980
rect -14150 89910 -14140 89980
rect -14360 89860 -14140 89910
rect -13860 90090 -13640 90140
rect -13860 90020 -13850 90090
rect -13650 90020 -13640 90090
rect -13860 89980 -13640 90020
rect -13860 89910 -13850 89980
rect -13650 89910 -13640 89980
rect -13860 89860 -13640 89910
rect -13360 90090 -13140 90140
rect -13360 90020 -13350 90090
rect -13150 90020 -13140 90090
rect -13360 89980 -13140 90020
rect -13360 89910 -13350 89980
rect -13150 89910 -13140 89980
rect -13360 89860 -13140 89910
rect -12860 90090 -12640 90140
rect -12860 90020 -12850 90090
rect -12650 90020 -12640 90090
rect -12860 89980 -12640 90020
rect -12860 89910 -12850 89980
rect -12650 89910 -12640 89980
rect -12860 89860 -12640 89910
rect -12360 90090 -12140 90140
rect -12360 90020 -12350 90090
rect -12150 90020 -12140 90090
rect -12360 89980 -12140 90020
rect -12360 89910 -12350 89980
rect -12150 89910 -12140 89980
rect -12360 89860 -12140 89910
rect -16000 89850 -12000 89860
rect -16000 89650 -15980 89850
rect -15910 89650 -15590 89850
rect -15520 89650 -15480 89850
rect -15410 89650 -15090 89850
rect -15020 89650 -14980 89850
rect -14910 89650 -14590 89850
rect -14520 89650 -14480 89850
rect -14410 89650 -14090 89850
rect -14020 89650 -13980 89850
rect -13910 89650 -13590 89850
rect -13520 89650 -13480 89850
rect -13410 89650 -13090 89850
rect -13020 89650 -12980 89850
rect -12910 89650 -12590 89850
rect -12520 89650 -12480 89850
rect -12410 89650 -12090 89850
rect -12020 89650 -12000 89850
rect -16000 89640 -12000 89650
rect -15860 89590 -15640 89640
rect -15860 89520 -15850 89590
rect -15650 89520 -15640 89590
rect -15860 89480 -15640 89520
rect -15860 89410 -15850 89480
rect -15650 89410 -15640 89480
rect -15860 89360 -15640 89410
rect -15360 89590 -15140 89640
rect -15360 89520 -15350 89590
rect -15150 89520 -15140 89590
rect -15360 89480 -15140 89520
rect -15360 89410 -15350 89480
rect -15150 89410 -15140 89480
rect -15360 89360 -15140 89410
rect -14860 89590 -14640 89640
rect -14860 89520 -14850 89590
rect -14650 89520 -14640 89590
rect -14860 89480 -14640 89520
rect -14860 89410 -14850 89480
rect -14650 89410 -14640 89480
rect -14860 89360 -14640 89410
rect -14360 89590 -14140 89640
rect -14360 89520 -14350 89590
rect -14150 89520 -14140 89590
rect -14360 89480 -14140 89520
rect -14360 89410 -14350 89480
rect -14150 89410 -14140 89480
rect -14360 89360 -14140 89410
rect -13860 89590 -13640 89640
rect -13860 89520 -13850 89590
rect -13650 89520 -13640 89590
rect -13860 89480 -13640 89520
rect -13860 89410 -13850 89480
rect -13650 89410 -13640 89480
rect -13860 89360 -13640 89410
rect -13360 89590 -13140 89640
rect -13360 89520 -13350 89590
rect -13150 89520 -13140 89590
rect -13360 89480 -13140 89520
rect -13360 89410 -13350 89480
rect -13150 89410 -13140 89480
rect -13360 89360 -13140 89410
rect -12860 89590 -12640 89640
rect -12860 89520 -12850 89590
rect -12650 89520 -12640 89590
rect -12860 89480 -12640 89520
rect -12860 89410 -12850 89480
rect -12650 89410 -12640 89480
rect -12860 89360 -12640 89410
rect -12360 89590 -12140 89640
rect -12360 89520 -12350 89590
rect -12150 89520 -12140 89590
rect -12360 89480 -12140 89520
rect -12360 89410 -12350 89480
rect -12150 89410 -12140 89480
rect -12360 89360 -12140 89410
rect -16000 89350 -12000 89360
rect -16000 89150 -15980 89350
rect -15910 89150 -15590 89350
rect -15520 89150 -15480 89350
rect -15410 89150 -15090 89350
rect -15020 89150 -14980 89350
rect -14910 89150 -14590 89350
rect -14520 89150 -14480 89350
rect -14410 89150 -14090 89350
rect -14020 89150 -13980 89350
rect -13910 89150 -13590 89350
rect -13520 89150 -13480 89350
rect -13410 89150 -13090 89350
rect -13020 89150 -12980 89350
rect -12910 89150 -12590 89350
rect -12520 89150 -12480 89350
rect -12410 89150 -12090 89350
rect -12020 89150 -12000 89350
rect -16000 89140 -12000 89150
rect -15860 89090 -15640 89140
rect -15860 89020 -15850 89090
rect -15650 89020 -15640 89090
rect -15860 88980 -15640 89020
rect -15860 88910 -15850 88980
rect -15650 88910 -15640 88980
rect -15860 88860 -15640 88910
rect -15360 89090 -15140 89140
rect -15360 89020 -15350 89090
rect -15150 89020 -15140 89090
rect -15360 88980 -15140 89020
rect -15360 88910 -15350 88980
rect -15150 88910 -15140 88980
rect -15360 88860 -15140 88910
rect -14860 89090 -14640 89140
rect -14860 89020 -14850 89090
rect -14650 89020 -14640 89090
rect -14860 88980 -14640 89020
rect -14860 88910 -14850 88980
rect -14650 88910 -14640 88980
rect -14860 88860 -14640 88910
rect -14360 89090 -14140 89140
rect -14360 89020 -14350 89090
rect -14150 89020 -14140 89090
rect -14360 88980 -14140 89020
rect -14360 88910 -14350 88980
rect -14150 88910 -14140 88980
rect -14360 88860 -14140 88910
rect -13860 89090 -13640 89140
rect -13860 89020 -13850 89090
rect -13650 89020 -13640 89090
rect -13860 88980 -13640 89020
rect -13860 88910 -13850 88980
rect -13650 88910 -13640 88980
rect -13860 88860 -13640 88910
rect -13360 89090 -13140 89140
rect -13360 89020 -13350 89090
rect -13150 89020 -13140 89090
rect -13360 88980 -13140 89020
rect -13360 88910 -13350 88980
rect -13150 88910 -13140 88980
rect -13360 88860 -13140 88910
rect -12860 89090 -12640 89140
rect -12860 89020 -12850 89090
rect -12650 89020 -12640 89090
rect -12860 88980 -12640 89020
rect -12860 88910 -12850 88980
rect -12650 88910 -12640 88980
rect -12860 88860 -12640 88910
rect -12360 89090 -12140 89140
rect -12360 89020 -12350 89090
rect -12150 89020 -12140 89090
rect -12360 88980 -12140 89020
rect -12360 88910 -12350 88980
rect -12150 88910 -12140 88980
rect -12360 88860 -12140 88910
rect -16000 88850 -12000 88860
rect -16000 88650 -15980 88850
rect -15910 88650 -15590 88850
rect -15520 88650 -15480 88850
rect -15410 88650 -15090 88850
rect -15020 88650 -14980 88850
rect -14910 88650 -14590 88850
rect -14520 88650 -14480 88850
rect -14410 88650 -14090 88850
rect -14020 88650 -13980 88850
rect -13910 88650 -13590 88850
rect -13520 88650 -13480 88850
rect -13410 88650 -13090 88850
rect -13020 88650 -12980 88850
rect -12910 88650 -12590 88850
rect -12520 88650 -12480 88850
rect -12410 88650 -12090 88850
rect -12020 88650 -12000 88850
rect -16000 88640 -12000 88650
rect -15860 88590 -15640 88640
rect -15860 88520 -15850 88590
rect -15650 88520 -15640 88590
rect -15860 88480 -15640 88520
rect -15860 88410 -15850 88480
rect -15650 88410 -15640 88480
rect -15860 88360 -15640 88410
rect -15360 88590 -15140 88640
rect -15360 88520 -15350 88590
rect -15150 88520 -15140 88590
rect -15360 88480 -15140 88520
rect -15360 88410 -15350 88480
rect -15150 88410 -15140 88480
rect -15360 88360 -15140 88410
rect -14860 88590 -14640 88640
rect -14860 88520 -14850 88590
rect -14650 88520 -14640 88590
rect -14860 88480 -14640 88520
rect -14860 88410 -14850 88480
rect -14650 88410 -14640 88480
rect -14860 88360 -14640 88410
rect -14360 88590 -14140 88640
rect -14360 88520 -14350 88590
rect -14150 88520 -14140 88590
rect -14360 88480 -14140 88520
rect -14360 88410 -14350 88480
rect -14150 88410 -14140 88480
rect -14360 88360 -14140 88410
rect -13860 88590 -13640 88640
rect -13860 88520 -13850 88590
rect -13650 88520 -13640 88590
rect -13860 88480 -13640 88520
rect -13860 88410 -13850 88480
rect -13650 88410 -13640 88480
rect -13860 88360 -13640 88410
rect -13360 88590 -13140 88640
rect -13360 88520 -13350 88590
rect -13150 88520 -13140 88590
rect -13360 88480 -13140 88520
rect -13360 88410 -13350 88480
rect -13150 88410 -13140 88480
rect -13360 88360 -13140 88410
rect -12860 88590 -12640 88640
rect -12860 88520 -12850 88590
rect -12650 88520 -12640 88590
rect -12860 88480 -12640 88520
rect -12860 88410 -12850 88480
rect -12650 88410 -12640 88480
rect -12860 88360 -12640 88410
rect -12360 88590 -12140 88640
rect -12360 88520 -12350 88590
rect -12150 88520 -12140 88590
rect -12360 88480 -12140 88520
rect -12360 88410 -12350 88480
rect -12150 88410 -12140 88480
rect -12360 88360 -12140 88410
rect -16000 88350 -12000 88360
rect -16000 88150 -15980 88350
rect -15910 88150 -15590 88350
rect -15520 88150 -15480 88350
rect -15410 88150 -15090 88350
rect -15020 88150 -14980 88350
rect -14910 88150 -14590 88350
rect -14520 88150 -14480 88350
rect -14410 88150 -14090 88350
rect -14020 88150 -13980 88350
rect -13910 88150 -13590 88350
rect -13520 88150 -13480 88350
rect -13410 88150 -13090 88350
rect -13020 88150 -12980 88350
rect -12910 88150 -12590 88350
rect -12520 88150 -12480 88350
rect -12410 88150 -12090 88350
rect -12020 88150 -12000 88350
rect -16000 88140 -12000 88150
rect -15860 88090 -15640 88140
rect -15860 88020 -15850 88090
rect -15650 88020 -15640 88090
rect -15860 87980 -15640 88020
rect -15860 87910 -15850 87980
rect -15650 87910 -15640 87980
rect -15860 87860 -15640 87910
rect -15360 88090 -15140 88140
rect -15360 88020 -15350 88090
rect -15150 88020 -15140 88090
rect -15360 87980 -15140 88020
rect -15360 87910 -15350 87980
rect -15150 87910 -15140 87980
rect -15360 87860 -15140 87910
rect -14860 88090 -14640 88140
rect -14860 88020 -14850 88090
rect -14650 88020 -14640 88090
rect -14860 87980 -14640 88020
rect -14860 87910 -14850 87980
rect -14650 87910 -14640 87980
rect -14860 87860 -14640 87910
rect -14360 88090 -14140 88140
rect -14360 88020 -14350 88090
rect -14150 88020 -14140 88090
rect -14360 87980 -14140 88020
rect -14360 87910 -14350 87980
rect -14150 87910 -14140 87980
rect -14360 87860 -14140 87910
rect -13860 88090 -13640 88140
rect -13860 88020 -13850 88090
rect -13650 88020 -13640 88090
rect -13860 87980 -13640 88020
rect -13860 87910 -13850 87980
rect -13650 87910 -13640 87980
rect -13860 87860 -13640 87910
rect -13360 88090 -13140 88140
rect -13360 88020 -13350 88090
rect -13150 88020 -13140 88090
rect -13360 87980 -13140 88020
rect -13360 87910 -13350 87980
rect -13150 87910 -13140 87980
rect -13360 87860 -13140 87910
rect -12860 88090 -12640 88140
rect -12860 88020 -12850 88090
rect -12650 88020 -12640 88090
rect -12860 87980 -12640 88020
rect -12860 87910 -12850 87980
rect -12650 87910 -12640 87980
rect -12860 87860 -12640 87910
rect -12360 88090 -12140 88140
rect -12360 88020 -12350 88090
rect -12150 88020 -12140 88090
rect -12360 87980 -12140 88020
rect -12360 87910 -12350 87980
rect -12150 87910 -12140 87980
rect -12360 87860 -12140 87910
rect -16000 87850 -12000 87860
rect -16000 87650 -15980 87850
rect -15910 87650 -15590 87850
rect -15520 87650 -15480 87850
rect -15410 87650 -15090 87850
rect -15020 87650 -14980 87850
rect -14910 87650 -14590 87850
rect -14520 87650 -14480 87850
rect -14410 87650 -14090 87850
rect -14020 87650 -13980 87850
rect -13910 87650 -13590 87850
rect -13520 87650 -13480 87850
rect -13410 87650 -13090 87850
rect -13020 87650 -12980 87850
rect -12910 87650 -12590 87850
rect -12520 87650 -12480 87850
rect -12410 87650 -12090 87850
rect -12020 87650 -12000 87850
rect -16000 87640 -12000 87650
rect -15860 87590 -15640 87640
rect -15860 87520 -15850 87590
rect -15650 87520 -15640 87590
rect -15860 87480 -15640 87520
rect -15860 87410 -15850 87480
rect -15650 87410 -15640 87480
rect -15860 87360 -15640 87410
rect -15360 87590 -15140 87640
rect -15360 87520 -15350 87590
rect -15150 87520 -15140 87590
rect -15360 87480 -15140 87520
rect -15360 87410 -15350 87480
rect -15150 87410 -15140 87480
rect -15360 87360 -15140 87410
rect -14860 87590 -14640 87640
rect -14860 87520 -14850 87590
rect -14650 87520 -14640 87590
rect -14860 87480 -14640 87520
rect -14860 87410 -14850 87480
rect -14650 87410 -14640 87480
rect -14860 87360 -14640 87410
rect -14360 87590 -14140 87640
rect -14360 87520 -14350 87590
rect -14150 87520 -14140 87590
rect -14360 87480 -14140 87520
rect -14360 87410 -14350 87480
rect -14150 87410 -14140 87480
rect -14360 87360 -14140 87410
rect -13860 87590 -13640 87640
rect -13860 87520 -13850 87590
rect -13650 87520 -13640 87590
rect -13860 87480 -13640 87520
rect -13860 87410 -13850 87480
rect -13650 87410 -13640 87480
rect -13860 87360 -13640 87410
rect -13360 87590 -13140 87640
rect -13360 87520 -13350 87590
rect -13150 87520 -13140 87590
rect -13360 87480 -13140 87520
rect -13360 87410 -13350 87480
rect -13150 87410 -13140 87480
rect -13360 87360 -13140 87410
rect -12860 87590 -12640 87640
rect -12860 87520 -12850 87590
rect -12650 87520 -12640 87590
rect -12860 87480 -12640 87520
rect -12860 87410 -12850 87480
rect -12650 87410 -12640 87480
rect -12860 87360 -12640 87410
rect -12360 87590 -12140 87640
rect -12360 87520 -12350 87590
rect -12150 87520 -12140 87590
rect -12360 87480 -12140 87520
rect -12360 87410 -12350 87480
rect -12150 87410 -12140 87480
rect -12360 87360 -12140 87410
rect -16000 87350 -12000 87360
rect -16000 87150 -15980 87350
rect -15910 87150 -15590 87350
rect -15520 87150 -15480 87350
rect -15410 87150 -15090 87350
rect -15020 87150 -14980 87350
rect -14910 87150 -14590 87350
rect -14520 87150 -14480 87350
rect -14410 87150 -14090 87350
rect -14020 87150 -13980 87350
rect -13910 87150 -13590 87350
rect -13520 87150 -13480 87350
rect -13410 87150 -13090 87350
rect -13020 87150 -12980 87350
rect -12910 87150 -12590 87350
rect -12520 87150 -12480 87350
rect -12410 87150 -12090 87350
rect -12020 87150 -12000 87350
rect -16000 87140 -12000 87150
rect -15860 87090 -15640 87140
rect -15860 87020 -15850 87090
rect -15650 87020 -15640 87090
rect -15860 86980 -15640 87020
rect -15860 86910 -15850 86980
rect -15650 86910 -15640 86980
rect -15860 86860 -15640 86910
rect -15360 87090 -15140 87140
rect -15360 87020 -15350 87090
rect -15150 87020 -15140 87090
rect -15360 86980 -15140 87020
rect -15360 86910 -15350 86980
rect -15150 86910 -15140 86980
rect -15360 86860 -15140 86910
rect -14860 87090 -14640 87140
rect -14860 87020 -14850 87090
rect -14650 87020 -14640 87090
rect -14860 86980 -14640 87020
rect -14860 86910 -14850 86980
rect -14650 86910 -14640 86980
rect -14860 86860 -14640 86910
rect -14360 87090 -14140 87140
rect -14360 87020 -14350 87090
rect -14150 87020 -14140 87090
rect -14360 86980 -14140 87020
rect -14360 86910 -14350 86980
rect -14150 86910 -14140 86980
rect -14360 86860 -14140 86910
rect -13860 87090 -13640 87140
rect -13860 87020 -13850 87090
rect -13650 87020 -13640 87090
rect -13860 86980 -13640 87020
rect -13860 86910 -13850 86980
rect -13650 86910 -13640 86980
rect -13860 86860 -13640 86910
rect -13360 87090 -13140 87140
rect -13360 87020 -13350 87090
rect -13150 87020 -13140 87090
rect -13360 86980 -13140 87020
rect -13360 86910 -13350 86980
rect -13150 86910 -13140 86980
rect -13360 86860 -13140 86910
rect -12860 87090 -12640 87140
rect -12860 87020 -12850 87090
rect -12650 87020 -12640 87090
rect -12860 86980 -12640 87020
rect -12860 86910 -12850 86980
rect -12650 86910 -12640 86980
rect -12860 86860 -12640 86910
rect -12360 87090 -12140 87140
rect -12360 87020 -12350 87090
rect -12150 87020 -12140 87090
rect -12360 86980 -12140 87020
rect -12360 86910 -12350 86980
rect -12150 86910 -12140 86980
rect -12360 86860 -12140 86910
rect -16000 86850 -12000 86860
rect -16000 86650 -15980 86850
rect -15910 86650 -15590 86850
rect -15520 86650 -15480 86850
rect -15410 86650 -15090 86850
rect -15020 86650 -14980 86850
rect -14910 86650 -14590 86850
rect -14520 86650 -14480 86850
rect -14410 86650 -14090 86850
rect -14020 86650 -13980 86850
rect -13910 86650 -13590 86850
rect -13520 86650 -13480 86850
rect -13410 86650 -13090 86850
rect -13020 86650 -12980 86850
rect -12910 86650 -12590 86850
rect -12520 86650 -12480 86850
rect -12410 86650 -12090 86850
rect -12020 86650 -12000 86850
rect -16000 86640 -12000 86650
rect -15860 86590 -15640 86640
rect -15860 86520 -15850 86590
rect -15650 86520 -15640 86590
rect -15860 86480 -15640 86520
rect -15860 86410 -15850 86480
rect -15650 86410 -15640 86480
rect -15860 86360 -15640 86410
rect -15360 86590 -15140 86640
rect -15360 86520 -15350 86590
rect -15150 86520 -15140 86590
rect -15360 86480 -15140 86520
rect -15360 86410 -15350 86480
rect -15150 86410 -15140 86480
rect -15360 86360 -15140 86410
rect -14860 86590 -14640 86640
rect -14860 86520 -14850 86590
rect -14650 86520 -14640 86590
rect -14860 86480 -14640 86520
rect -14860 86410 -14850 86480
rect -14650 86410 -14640 86480
rect -14860 86360 -14640 86410
rect -14360 86590 -14140 86640
rect -14360 86520 -14350 86590
rect -14150 86520 -14140 86590
rect -14360 86480 -14140 86520
rect -14360 86410 -14350 86480
rect -14150 86410 -14140 86480
rect -14360 86360 -14140 86410
rect -13860 86590 -13640 86640
rect -13860 86520 -13850 86590
rect -13650 86520 -13640 86590
rect -13860 86480 -13640 86520
rect -13860 86410 -13850 86480
rect -13650 86410 -13640 86480
rect -13860 86360 -13640 86410
rect -13360 86590 -13140 86640
rect -13360 86520 -13350 86590
rect -13150 86520 -13140 86590
rect -13360 86480 -13140 86520
rect -13360 86410 -13350 86480
rect -13150 86410 -13140 86480
rect -13360 86360 -13140 86410
rect -12860 86590 -12640 86640
rect -12860 86520 -12850 86590
rect -12650 86520 -12640 86590
rect -12860 86480 -12640 86520
rect -12860 86410 -12850 86480
rect -12650 86410 -12640 86480
rect -12860 86360 -12640 86410
rect -12360 86590 -12140 86640
rect -12360 86520 -12350 86590
rect -12150 86520 -12140 86590
rect -12360 86480 -12140 86520
rect -12360 86410 -12350 86480
rect -12150 86410 -12140 86480
rect -12360 86360 -12140 86410
rect -16000 86350 -12000 86360
rect -16000 86150 -15980 86350
rect -15910 86150 -15590 86350
rect -15520 86150 -15480 86350
rect -15410 86150 -15090 86350
rect -15020 86150 -14980 86350
rect -14910 86150 -14590 86350
rect -14520 86150 -14480 86350
rect -14410 86150 -14090 86350
rect -14020 86150 -13980 86350
rect -13910 86150 -13590 86350
rect -13520 86150 -13480 86350
rect -13410 86150 -13090 86350
rect -13020 86150 -12980 86350
rect -12910 86150 -12590 86350
rect -12520 86150 -12480 86350
rect -12410 86150 -12090 86350
rect -12020 86150 -12000 86350
rect -16000 86140 -12000 86150
rect -15860 86090 -15640 86140
rect -15860 86020 -15850 86090
rect -15650 86020 -15640 86090
rect -15860 85980 -15640 86020
rect -15860 85910 -15850 85980
rect -15650 85910 -15640 85980
rect -15860 85860 -15640 85910
rect -15360 86090 -15140 86140
rect -15360 86020 -15350 86090
rect -15150 86020 -15140 86090
rect -15360 85980 -15140 86020
rect -15360 85910 -15350 85980
rect -15150 85910 -15140 85980
rect -15360 85860 -15140 85910
rect -14860 86090 -14640 86140
rect -14860 86020 -14850 86090
rect -14650 86020 -14640 86090
rect -14860 85980 -14640 86020
rect -14860 85910 -14850 85980
rect -14650 85910 -14640 85980
rect -14860 85860 -14640 85910
rect -14360 86090 -14140 86140
rect -14360 86020 -14350 86090
rect -14150 86020 -14140 86090
rect -14360 85980 -14140 86020
rect -14360 85910 -14350 85980
rect -14150 85910 -14140 85980
rect -14360 85860 -14140 85910
rect -13860 86090 -13640 86140
rect -13860 86020 -13850 86090
rect -13650 86020 -13640 86090
rect -13860 85980 -13640 86020
rect -13860 85910 -13850 85980
rect -13650 85910 -13640 85980
rect -13860 85860 -13640 85910
rect -13360 86090 -13140 86140
rect -13360 86020 -13350 86090
rect -13150 86020 -13140 86090
rect -13360 85980 -13140 86020
rect -13360 85910 -13350 85980
rect -13150 85910 -13140 85980
rect -13360 85860 -13140 85910
rect -12860 86090 -12640 86140
rect -12860 86020 -12850 86090
rect -12650 86020 -12640 86090
rect -12860 85980 -12640 86020
rect -12860 85910 -12850 85980
rect -12650 85910 -12640 85980
rect -12860 85860 -12640 85910
rect -12360 86090 -12140 86140
rect -12360 86020 -12350 86090
rect -12150 86020 -12140 86090
rect -12360 85980 -12140 86020
rect -12360 85910 -12350 85980
rect -12150 85910 -12140 85980
rect -12360 85860 -12140 85910
rect 96140 85980 96360 86000
rect 96140 85910 96150 85980
rect 96350 85910 96360 85980
rect 96140 85860 96360 85910
rect 96640 85980 96860 86000
rect 96640 85910 96650 85980
rect 96850 85910 96860 85980
rect 96640 85860 96860 85910
rect 97140 85980 97360 86000
rect 97140 85910 97150 85980
rect 97350 85910 97360 85980
rect 97140 85860 97360 85910
rect 97640 85980 97860 86000
rect 97640 85910 97650 85980
rect 97850 85910 97860 85980
rect 97640 85860 97860 85910
rect 98140 85980 98360 86000
rect 98140 85910 98150 85980
rect 98350 85910 98360 85980
rect 98140 85860 98360 85910
rect 98640 85980 98860 86000
rect 98640 85910 98650 85980
rect 98850 85910 98860 85980
rect 98640 85860 98860 85910
rect 99140 85980 99360 86000
rect 99140 85910 99150 85980
rect 99350 85910 99360 85980
rect 99140 85860 99360 85910
rect 99640 85980 99860 86000
rect 99640 85910 99650 85980
rect 99850 85910 99860 85980
rect 99640 85860 99860 85910
rect -16000 85850 -12000 85860
rect -16000 85650 -15980 85850
rect -15910 85650 -15590 85850
rect -15520 85650 -15480 85850
rect -15410 85650 -15090 85850
rect -15020 85650 -14980 85850
rect -14910 85650 -14590 85850
rect -14520 85650 -14480 85850
rect -14410 85650 -14090 85850
rect -14020 85650 -13980 85850
rect -13910 85650 -13590 85850
rect -13520 85650 -13480 85850
rect -13410 85650 -13090 85850
rect -13020 85650 -12980 85850
rect -12910 85650 -12590 85850
rect -12520 85650 -12480 85850
rect -12410 85650 -12090 85850
rect -12020 85650 -12000 85850
rect -16000 85640 -12000 85650
rect 96000 85850 100000 85860
rect 96000 85650 96020 85850
rect 96090 85650 96410 85850
rect 96480 85650 96520 85850
rect 96590 85650 96910 85850
rect 96980 85650 97020 85850
rect 97090 85650 97410 85850
rect 97480 85650 97520 85850
rect 97590 85650 97910 85850
rect 97980 85650 98020 85850
rect 98090 85650 98410 85850
rect 98480 85650 98520 85850
rect 98590 85650 98910 85850
rect 98980 85650 99020 85850
rect 99090 85650 99410 85850
rect 99480 85650 99520 85850
rect 99590 85650 99910 85850
rect 99980 85650 100000 85850
rect 96000 85640 100000 85650
rect -15860 85590 -15640 85640
rect -15860 85520 -15850 85590
rect -15650 85520 -15640 85590
rect -15860 85480 -15640 85520
rect -15860 85410 -15850 85480
rect -15650 85410 -15640 85480
rect -15860 85360 -15640 85410
rect -15360 85590 -15140 85640
rect -15360 85520 -15350 85590
rect -15150 85520 -15140 85590
rect -15360 85480 -15140 85520
rect -15360 85410 -15350 85480
rect -15150 85410 -15140 85480
rect -15360 85360 -15140 85410
rect -14860 85590 -14640 85640
rect -14860 85520 -14850 85590
rect -14650 85520 -14640 85590
rect -14860 85480 -14640 85520
rect -14860 85410 -14850 85480
rect -14650 85410 -14640 85480
rect -14860 85360 -14640 85410
rect -14360 85590 -14140 85640
rect -14360 85520 -14350 85590
rect -14150 85520 -14140 85590
rect -14360 85480 -14140 85520
rect -14360 85410 -14350 85480
rect -14150 85410 -14140 85480
rect -14360 85360 -14140 85410
rect -13860 85590 -13640 85640
rect -13860 85520 -13850 85590
rect -13650 85520 -13640 85590
rect -13860 85480 -13640 85520
rect -13860 85410 -13850 85480
rect -13650 85410 -13640 85480
rect -13860 85360 -13640 85410
rect -13360 85590 -13140 85640
rect -13360 85520 -13350 85590
rect -13150 85520 -13140 85590
rect -13360 85480 -13140 85520
rect -13360 85410 -13350 85480
rect -13150 85410 -13140 85480
rect -13360 85360 -13140 85410
rect -12860 85590 -12640 85640
rect -12860 85520 -12850 85590
rect -12650 85520 -12640 85590
rect -12860 85480 -12640 85520
rect -12860 85410 -12850 85480
rect -12650 85410 -12640 85480
rect -12860 85360 -12640 85410
rect -12360 85590 -12140 85640
rect -12360 85520 -12350 85590
rect -12150 85520 -12140 85590
rect -12360 85480 -12140 85520
rect -12360 85410 -12350 85480
rect -12150 85410 -12140 85480
rect -12360 85360 -12140 85410
rect 96140 85590 96360 85640
rect 96140 85520 96150 85590
rect 96350 85520 96360 85590
rect 96140 85480 96360 85520
rect 96140 85410 96150 85480
rect 96350 85410 96360 85480
rect 96140 85360 96360 85410
rect 96640 85590 96860 85640
rect 96640 85520 96650 85590
rect 96850 85520 96860 85590
rect 96640 85480 96860 85520
rect 96640 85410 96650 85480
rect 96850 85410 96860 85480
rect 96640 85360 96860 85410
rect 97140 85590 97360 85640
rect 97140 85520 97150 85590
rect 97350 85520 97360 85590
rect 97140 85480 97360 85520
rect 97140 85410 97150 85480
rect 97350 85410 97360 85480
rect 97140 85360 97360 85410
rect 97640 85590 97860 85640
rect 97640 85520 97650 85590
rect 97850 85520 97860 85590
rect 97640 85480 97860 85520
rect 97640 85410 97650 85480
rect 97850 85410 97860 85480
rect 97640 85360 97860 85410
rect 98140 85590 98360 85640
rect 98140 85520 98150 85590
rect 98350 85520 98360 85590
rect 98140 85480 98360 85520
rect 98140 85410 98150 85480
rect 98350 85410 98360 85480
rect 98140 85360 98360 85410
rect 98640 85590 98860 85640
rect 98640 85520 98650 85590
rect 98850 85520 98860 85590
rect 98640 85480 98860 85520
rect 98640 85410 98650 85480
rect 98850 85410 98860 85480
rect 98640 85360 98860 85410
rect 99140 85590 99360 85640
rect 99140 85520 99150 85590
rect 99350 85520 99360 85590
rect 99140 85480 99360 85520
rect 99140 85410 99150 85480
rect 99350 85410 99360 85480
rect 99140 85360 99360 85410
rect 99640 85590 99860 85640
rect 99640 85520 99650 85590
rect 99850 85520 99860 85590
rect 99640 85480 99860 85520
rect 99640 85410 99650 85480
rect 99850 85410 99860 85480
rect 99640 85360 99860 85410
rect -16000 85350 -12000 85360
rect -16000 85150 -15980 85350
rect -15910 85150 -15590 85350
rect -15520 85150 -15480 85350
rect -15410 85150 -15090 85350
rect -15020 85150 -14980 85350
rect -14910 85150 -14590 85350
rect -14520 85150 -14480 85350
rect -14410 85150 -14090 85350
rect -14020 85150 -13980 85350
rect -13910 85150 -13590 85350
rect -13520 85150 -13480 85350
rect -13410 85150 -13090 85350
rect -13020 85150 -12980 85350
rect -12910 85150 -12590 85350
rect -12520 85150 -12480 85350
rect -12410 85150 -12090 85350
rect -12020 85150 -12000 85350
rect -16000 85140 -12000 85150
rect 96000 85350 100000 85360
rect 96000 85150 96020 85350
rect 96090 85150 96410 85350
rect 96480 85150 96520 85350
rect 96590 85150 96910 85350
rect 96980 85150 97020 85350
rect 97090 85150 97410 85350
rect 97480 85150 97520 85350
rect 97590 85150 97910 85350
rect 97980 85150 98020 85350
rect 98090 85150 98410 85350
rect 98480 85150 98520 85350
rect 98590 85150 98910 85350
rect 98980 85150 99020 85350
rect 99090 85150 99410 85350
rect 99480 85150 99520 85350
rect 99590 85150 99910 85350
rect 99980 85150 100000 85350
rect 96000 85140 100000 85150
rect -15860 85090 -15640 85140
rect -15860 85020 -15850 85090
rect -15650 85020 -15640 85090
rect -15860 84980 -15640 85020
rect -15860 84910 -15850 84980
rect -15650 84910 -15640 84980
rect -15860 84860 -15640 84910
rect -15360 85090 -15140 85140
rect -15360 85020 -15350 85090
rect -15150 85020 -15140 85090
rect -15360 84980 -15140 85020
rect -15360 84910 -15350 84980
rect -15150 84910 -15140 84980
rect -15360 84860 -15140 84910
rect -14860 85090 -14640 85140
rect -14860 85020 -14850 85090
rect -14650 85020 -14640 85090
rect -14860 84980 -14640 85020
rect -14860 84910 -14850 84980
rect -14650 84910 -14640 84980
rect -14860 84860 -14640 84910
rect -14360 85090 -14140 85140
rect -14360 85020 -14350 85090
rect -14150 85020 -14140 85090
rect -14360 84980 -14140 85020
rect -14360 84910 -14350 84980
rect -14150 84910 -14140 84980
rect -14360 84860 -14140 84910
rect -13860 85090 -13640 85140
rect -13860 85020 -13850 85090
rect -13650 85020 -13640 85090
rect -13860 84980 -13640 85020
rect -13860 84910 -13850 84980
rect -13650 84910 -13640 84980
rect -13860 84860 -13640 84910
rect -13360 85090 -13140 85140
rect -13360 85020 -13350 85090
rect -13150 85020 -13140 85090
rect -13360 84980 -13140 85020
rect -13360 84910 -13350 84980
rect -13150 84910 -13140 84980
rect -13360 84860 -13140 84910
rect -12860 85090 -12640 85140
rect -12860 85020 -12850 85090
rect -12650 85020 -12640 85090
rect -12860 84980 -12640 85020
rect -12860 84910 -12850 84980
rect -12650 84910 -12640 84980
rect -12860 84860 -12640 84910
rect -12360 85090 -12140 85140
rect -12360 85020 -12350 85090
rect -12150 85020 -12140 85090
rect -12360 84980 -12140 85020
rect -12360 84910 -12350 84980
rect -12150 84910 -12140 84980
rect -12360 84860 -12140 84910
rect 96140 85090 96360 85140
rect 96140 85020 96150 85090
rect 96350 85020 96360 85090
rect 96140 84980 96360 85020
rect 96140 84910 96150 84980
rect 96350 84910 96360 84980
rect 96140 84860 96360 84910
rect 96640 85090 96860 85140
rect 96640 85020 96650 85090
rect 96850 85020 96860 85090
rect 96640 84980 96860 85020
rect 96640 84910 96650 84980
rect 96850 84910 96860 84980
rect 96640 84860 96860 84910
rect 97140 85090 97360 85140
rect 97140 85020 97150 85090
rect 97350 85020 97360 85090
rect 97140 84980 97360 85020
rect 97140 84910 97150 84980
rect 97350 84910 97360 84980
rect 97140 84860 97360 84910
rect 97640 85090 97860 85140
rect 97640 85020 97650 85090
rect 97850 85020 97860 85090
rect 97640 84980 97860 85020
rect 97640 84910 97650 84980
rect 97850 84910 97860 84980
rect 97640 84860 97860 84910
rect 98140 85090 98360 85140
rect 98140 85020 98150 85090
rect 98350 85020 98360 85090
rect 98140 84980 98360 85020
rect 98140 84910 98150 84980
rect 98350 84910 98360 84980
rect 98140 84860 98360 84910
rect 98640 85090 98860 85140
rect 98640 85020 98650 85090
rect 98850 85020 98860 85090
rect 98640 84980 98860 85020
rect 98640 84910 98650 84980
rect 98850 84910 98860 84980
rect 98640 84860 98860 84910
rect 99140 85090 99360 85140
rect 99140 85020 99150 85090
rect 99350 85020 99360 85090
rect 99140 84980 99360 85020
rect 99140 84910 99150 84980
rect 99350 84910 99360 84980
rect 99140 84860 99360 84910
rect 99640 85090 99860 85140
rect 99640 85020 99650 85090
rect 99850 85020 99860 85090
rect 99640 84980 99860 85020
rect 99640 84910 99650 84980
rect 99850 84910 99860 84980
rect 99640 84860 99860 84910
rect -16000 84850 -12000 84860
rect -16000 84650 -15980 84850
rect -15910 84650 -15590 84850
rect -15520 84650 -15480 84850
rect -15410 84650 -15090 84850
rect -15020 84650 -14980 84850
rect -14910 84650 -14590 84850
rect -14520 84650 -14480 84850
rect -14410 84650 -14090 84850
rect -14020 84650 -13980 84850
rect -13910 84650 -13590 84850
rect -13520 84650 -13480 84850
rect -13410 84650 -13090 84850
rect -13020 84650 -12980 84850
rect -12910 84650 -12590 84850
rect -12520 84650 -12480 84850
rect -12410 84650 -12090 84850
rect -12020 84650 -12000 84850
rect -16000 84640 -12000 84650
rect 96000 84850 100000 84860
rect 96000 84650 96020 84850
rect 96090 84650 96410 84850
rect 96480 84650 96520 84850
rect 96590 84650 96910 84850
rect 96980 84650 97020 84850
rect 97090 84650 97410 84850
rect 97480 84650 97520 84850
rect 97590 84650 97910 84850
rect 97980 84650 98020 84850
rect 98090 84650 98410 84850
rect 98480 84650 98520 84850
rect 98590 84650 98910 84850
rect 98980 84650 99020 84850
rect 99090 84650 99410 84850
rect 99480 84650 99520 84850
rect 99590 84650 99910 84850
rect 99980 84650 100000 84850
rect 96000 84640 100000 84650
rect -15860 84590 -15640 84640
rect -15860 84520 -15850 84590
rect -15650 84520 -15640 84590
rect -15860 84480 -15640 84520
rect -15860 84410 -15850 84480
rect -15650 84410 -15640 84480
rect -15860 84360 -15640 84410
rect -15360 84590 -15140 84640
rect -15360 84520 -15350 84590
rect -15150 84520 -15140 84590
rect -15360 84480 -15140 84520
rect -15360 84410 -15350 84480
rect -15150 84410 -15140 84480
rect -15360 84360 -15140 84410
rect -14860 84590 -14640 84640
rect -14860 84520 -14850 84590
rect -14650 84520 -14640 84590
rect -14860 84480 -14640 84520
rect -14860 84410 -14850 84480
rect -14650 84410 -14640 84480
rect -14860 84360 -14640 84410
rect -14360 84590 -14140 84640
rect -14360 84520 -14350 84590
rect -14150 84520 -14140 84590
rect -14360 84480 -14140 84520
rect -14360 84410 -14350 84480
rect -14150 84410 -14140 84480
rect -14360 84360 -14140 84410
rect -13860 84590 -13640 84640
rect -13860 84520 -13850 84590
rect -13650 84520 -13640 84590
rect -13860 84480 -13640 84520
rect -13860 84410 -13850 84480
rect -13650 84410 -13640 84480
rect -13860 84360 -13640 84410
rect -13360 84590 -13140 84640
rect -13360 84520 -13350 84590
rect -13150 84520 -13140 84590
rect -13360 84480 -13140 84520
rect -13360 84410 -13350 84480
rect -13150 84410 -13140 84480
rect -13360 84360 -13140 84410
rect -12860 84590 -12640 84640
rect -12860 84520 -12850 84590
rect -12650 84520 -12640 84590
rect -12860 84480 -12640 84520
rect -12860 84410 -12850 84480
rect -12650 84410 -12640 84480
rect -12860 84360 -12640 84410
rect -12360 84590 -12140 84640
rect -12360 84520 -12350 84590
rect -12150 84520 -12140 84590
rect -12360 84480 -12140 84520
rect -12360 84410 -12350 84480
rect -12150 84410 -12140 84480
rect -12360 84360 -12140 84410
rect 96140 84590 96360 84640
rect 96140 84520 96150 84590
rect 96350 84520 96360 84590
rect 96140 84480 96360 84520
rect 96140 84410 96150 84480
rect 96350 84410 96360 84480
rect 96140 84360 96360 84410
rect 96640 84590 96860 84640
rect 96640 84520 96650 84590
rect 96850 84520 96860 84590
rect 96640 84480 96860 84520
rect 96640 84410 96650 84480
rect 96850 84410 96860 84480
rect 96640 84360 96860 84410
rect 97140 84590 97360 84640
rect 97140 84520 97150 84590
rect 97350 84520 97360 84590
rect 97140 84480 97360 84520
rect 97140 84410 97150 84480
rect 97350 84410 97360 84480
rect 97140 84360 97360 84410
rect 97640 84590 97860 84640
rect 97640 84520 97650 84590
rect 97850 84520 97860 84590
rect 97640 84480 97860 84520
rect 97640 84410 97650 84480
rect 97850 84410 97860 84480
rect 97640 84360 97860 84410
rect 98140 84590 98360 84640
rect 98140 84520 98150 84590
rect 98350 84520 98360 84590
rect 98140 84480 98360 84520
rect 98140 84410 98150 84480
rect 98350 84410 98360 84480
rect 98140 84360 98360 84410
rect 98640 84590 98860 84640
rect 98640 84520 98650 84590
rect 98850 84520 98860 84590
rect 98640 84480 98860 84520
rect 98640 84410 98650 84480
rect 98850 84410 98860 84480
rect 98640 84360 98860 84410
rect 99140 84590 99360 84640
rect 99140 84520 99150 84590
rect 99350 84520 99360 84590
rect 99140 84480 99360 84520
rect 99140 84410 99150 84480
rect 99350 84410 99360 84480
rect 99140 84360 99360 84410
rect 99640 84590 99860 84640
rect 99640 84520 99650 84590
rect 99850 84520 99860 84590
rect 99640 84480 99860 84520
rect 99640 84410 99650 84480
rect 99850 84410 99860 84480
rect 99640 84360 99860 84410
rect -16000 84350 -12000 84360
rect -16000 84150 -15980 84350
rect -15910 84150 -15590 84350
rect -15520 84150 -15480 84350
rect -15410 84150 -15090 84350
rect -15020 84150 -14980 84350
rect -14910 84150 -14590 84350
rect -14520 84150 -14480 84350
rect -14410 84150 -14090 84350
rect -14020 84150 -13980 84350
rect -13910 84150 -13590 84350
rect -13520 84150 -13480 84350
rect -13410 84150 -13090 84350
rect -13020 84150 -12980 84350
rect -12910 84150 -12590 84350
rect -12520 84150 -12480 84350
rect -12410 84150 -12090 84350
rect -12020 84150 -12000 84350
rect -16000 84140 -12000 84150
rect 96000 84350 100000 84360
rect 96000 84150 96020 84350
rect 96090 84150 96410 84350
rect 96480 84150 96520 84350
rect 96590 84150 96910 84350
rect 96980 84150 97020 84350
rect 97090 84150 97410 84350
rect 97480 84150 97520 84350
rect 97590 84150 97910 84350
rect 97980 84150 98020 84350
rect 98090 84150 98410 84350
rect 98480 84150 98520 84350
rect 98590 84150 98910 84350
rect 98980 84150 99020 84350
rect 99090 84150 99410 84350
rect 99480 84150 99520 84350
rect 99590 84150 99910 84350
rect 99980 84150 100000 84350
rect 96000 84140 100000 84150
rect -15860 84090 -15640 84140
rect -15860 84020 -15850 84090
rect -15650 84020 -15640 84090
rect -15860 83980 -15640 84020
rect -15860 83910 -15850 83980
rect -15650 83910 -15640 83980
rect -15860 83860 -15640 83910
rect -15360 84090 -15140 84140
rect -15360 84020 -15350 84090
rect -15150 84020 -15140 84090
rect -15360 83980 -15140 84020
rect -15360 83910 -15350 83980
rect -15150 83910 -15140 83980
rect -15360 83860 -15140 83910
rect -14860 84090 -14640 84140
rect -14860 84020 -14850 84090
rect -14650 84020 -14640 84090
rect -14860 83980 -14640 84020
rect -14860 83910 -14850 83980
rect -14650 83910 -14640 83980
rect -14860 83860 -14640 83910
rect -14360 84090 -14140 84140
rect -14360 84020 -14350 84090
rect -14150 84020 -14140 84090
rect -14360 83980 -14140 84020
rect -14360 83910 -14350 83980
rect -14150 83910 -14140 83980
rect -14360 83860 -14140 83910
rect -13860 84090 -13640 84140
rect -13860 84020 -13850 84090
rect -13650 84020 -13640 84090
rect -13860 83980 -13640 84020
rect -13860 83910 -13850 83980
rect -13650 83910 -13640 83980
rect -13860 83860 -13640 83910
rect -13360 84090 -13140 84140
rect -13360 84020 -13350 84090
rect -13150 84020 -13140 84090
rect -13360 83980 -13140 84020
rect -13360 83910 -13350 83980
rect -13150 83910 -13140 83980
rect -13360 83860 -13140 83910
rect -12860 84090 -12640 84140
rect -12860 84020 -12850 84090
rect -12650 84020 -12640 84090
rect -12860 83980 -12640 84020
rect -12860 83910 -12850 83980
rect -12650 83910 -12640 83980
rect -12860 83860 -12640 83910
rect -12360 84090 -12140 84140
rect -12360 84020 -12350 84090
rect -12150 84020 -12140 84090
rect -12360 83980 -12140 84020
rect -12360 83910 -12350 83980
rect -12150 83910 -12140 83980
rect -12360 83860 -12140 83910
rect 96140 84090 96360 84140
rect 96140 84020 96150 84090
rect 96350 84020 96360 84090
rect 96140 83980 96360 84020
rect 96140 83910 96150 83980
rect 96350 83910 96360 83980
rect 96140 83860 96360 83910
rect 96640 84090 96860 84140
rect 96640 84020 96650 84090
rect 96850 84020 96860 84090
rect 96640 83980 96860 84020
rect 96640 83910 96650 83980
rect 96850 83910 96860 83980
rect 96640 83860 96860 83910
rect 97140 84090 97360 84140
rect 97140 84020 97150 84090
rect 97350 84020 97360 84090
rect 97140 83980 97360 84020
rect 97140 83910 97150 83980
rect 97350 83910 97360 83980
rect 97140 83860 97360 83910
rect 97640 84090 97860 84140
rect 97640 84020 97650 84090
rect 97850 84020 97860 84090
rect 97640 83980 97860 84020
rect 97640 83910 97650 83980
rect 97850 83910 97860 83980
rect 97640 83860 97860 83910
rect 98140 84090 98360 84140
rect 98140 84020 98150 84090
rect 98350 84020 98360 84090
rect 98140 83980 98360 84020
rect 98140 83910 98150 83980
rect 98350 83910 98360 83980
rect 98140 83860 98360 83910
rect 98640 84090 98860 84140
rect 98640 84020 98650 84090
rect 98850 84020 98860 84090
rect 98640 83980 98860 84020
rect 98640 83910 98650 83980
rect 98850 83910 98860 83980
rect 98640 83860 98860 83910
rect 99140 84090 99360 84140
rect 99140 84020 99150 84090
rect 99350 84020 99360 84090
rect 99140 83980 99360 84020
rect 99140 83910 99150 83980
rect 99350 83910 99360 83980
rect 99140 83860 99360 83910
rect 99640 84090 99860 84140
rect 99640 84020 99650 84090
rect 99850 84020 99860 84090
rect 99640 83980 99860 84020
rect 99640 83910 99650 83980
rect 99850 83910 99860 83980
rect 99640 83860 99860 83910
rect -16000 83850 -12000 83860
rect -16000 83650 -15980 83850
rect -15910 83650 -15590 83850
rect -15520 83650 -15480 83850
rect -15410 83650 -15090 83850
rect -15020 83650 -14980 83850
rect -14910 83650 -14590 83850
rect -14520 83650 -14480 83850
rect -14410 83650 -14090 83850
rect -14020 83650 -13980 83850
rect -13910 83650 -13590 83850
rect -13520 83650 -13480 83850
rect -13410 83650 -13090 83850
rect -13020 83650 -12980 83850
rect -12910 83650 -12590 83850
rect -12520 83650 -12480 83850
rect -12410 83650 -12090 83850
rect -12020 83650 -12000 83850
rect -16000 83640 -12000 83650
rect 96000 83850 100000 83860
rect 96000 83650 96020 83850
rect 96090 83650 96410 83850
rect 96480 83650 96520 83850
rect 96590 83650 96910 83850
rect 96980 83650 97020 83850
rect 97090 83650 97410 83850
rect 97480 83650 97520 83850
rect 97590 83650 97910 83850
rect 97980 83650 98020 83850
rect 98090 83650 98410 83850
rect 98480 83650 98520 83850
rect 98590 83650 98910 83850
rect 98980 83650 99020 83850
rect 99090 83650 99410 83850
rect 99480 83650 99520 83850
rect 99590 83650 99910 83850
rect 99980 83650 100000 83850
rect 96000 83640 100000 83650
rect -15860 83590 -15640 83640
rect -15860 83520 -15850 83590
rect -15650 83520 -15640 83590
rect -15860 83480 -15640 83520
rect -15860 83410 -15850 83480
rect -15650 83410 -15640 83480
rect -15860 83360 -15640 83410
rect -15360 83590 -15140 83640
rect -15360 83520 -15350 83590
rect -15150 83520 -15140 83590
rect -15360 83480 -15140 83520
rect -15360 83410 -15350 83480
rect -15150 83410 -15140 83480
rect -15360 83360 -15140 83410
rect -14860 83590 -14640 83640
rect -14860 83520 -14850 83590
rect -14650 83520 -14640 83590
rect -14860 83480 -14640 83520
rect -14860 83410 -14850 83480
rect -14650 83410 -14640 83480
rect -14860 83360 -14640 83410
rect -14360 83590 -14140 83640
rect -14360 83520 -14350 83590
rect -14150 83520 -14140 83590
rect -14360 83480 -14140 83520
rect -14360 83410 -14350 83480
rect -14150 83410 -14140 83480
rect -14360 83360 -14140 83410
rect -13860 83590 -13640 83640
rect -13860 83520 -13850 83590
rect -13650 83520 -13640 83590
rect -13860 83480 -13640 83520
rect -13860 83410 -13850 83480
rect -13650 83410 -13640 83480
rect -13860 83360 -13640 83410
rect -13360 83590 -13140 83640
rect -13360 83520 -13350 83590
rect -13150 83520 -13140 83590
rect -13360 83480 -13140 83520
rect -13360 83410 -13350 83480
rect -13150 83410 -13140 83480
rect -13360 83360 -13140 83410
rect -12860 83590 -12640 83640
rect -12860 83520 -12850 83590
rect -12650 83520 -12640 83590
rect -12860 83480 -12640 83520
rect -12860 83410 -12850 83480
rect -12650 83410 -12640 83480
rect -12860 83360 -12640 83410
rect -12360 83590 -12140 83640
rect -12360 83520 -12350 83590
rect -12150 83520 -12140 83590
rect -12360 83480 -12140 83520
rect -12360 83410 -12350 83480
rect -12150 83410 -12140 83480
rect -12360 83360 -12140 83410
rect 96140 83590 96360 83640
rect 96140 83520 96150 83590
rect 96350 83520 96360 83590
rect 96140 83480 96360 83520
rect 96140 83410 96150 83480
rect 96350 83410 96360 83480
rect 96140 83360 96360 83410
rect 96640 83590 96860 83640
rect 96640 83520 96650 83590
rect 96850 83520 96860 83590
rect 96640 83480 96860 83520
rect 96640 83410 96650 83480
rect 96850 83410 96860 83480
rect 96640 83360 96860 83410
rect 97140 83590 97360 83640
rect 97140 83520 97150 83590
rect 97350 83520 97360 83590
rect 97140 83480 97360 83520
rect 97140 83410 97150 83480
rect 97350 83410 97360 83480
rect 97140 83360 97360 83410
rect 97640 83590 97860 83640
rect 97640 83520 97650 83590
rect 97850 83520 97860 83590
rect 97640 83480 97860 83520
rect 97640 83410 97650 83480
rect 97850 83410 97860 83480
rect 97640 83360 97860 83410
rect 98140 83590 98360 83640
rect 98140 83520 98150 83590
rect 98350 83520 98360 83590
rect 98140 83480 98360 83520
rect 98140 83410 98150 83480
rect 98350 83410 98360 83480
rect 98140 83360 98360 83410
rect 98640 83590 98860 83640
rect 98640 83520 98650 83590
rect 98850 83520 98860 83590
rect 98640 83480 98860 83520
rect 98640 83410 98650 83480
rect 98850 83410 98860 83480
rect 98640 83360 98860 83410
rect 99140 83590 99360 83640
rect 99140 83520 99150 83590
rect 99350 83520 99360 83590
rect 99140 83480 99360 83520
rect 99140 83410 99150 83480
rect 99350 83410 99360 83480
rect 99140 83360 99360 83410
rect 99640 83590 99860 83640
rect 99640 83520 99650 83590
rect 99850 83520 99860 83590
rect 99640 83480 99860 83520
rect 99640 83410 99650 83480
rect 99850 83410 99860 83480
rect 99640 83360 99860 83410
rect -16000 83350 -12000 83360
rect -16000 83150 -15980 83350
rect -15910 83150 -15590 83350
rect -15520 83150 -15480 83350
rect -15410 83150 -15090 83350
rect -15020 83150 -14980 83350
rect -14910 83150 -14590 83350
rect -14520 83150 -14480 83350
rect -14410 83150 -14090 83350
rect -14020 83150 -13980 83350
rect -13910 83150 -13590 83350
rect -13520 83150 -13480 83350
rect -13410 83150 -13090 83350
rect -13020 83150 -12980 83350
rect -12910 83150 -12590 83350
rect -12520 83150 -12480 83350
rect -12410 83150 -12090 83350
rect -12020 83150 -12000 83350
rect -16000 83140 -12000 83150
rect 96000 83350 100000 83360
rect 96000 83150 96020 83350
rect 96090 83150 96410 83350
rect 96480 83150 96520 83350
rect 96590 83150 96910 83350
rect 96980 83150 97020 83350
rect 97090 83150 97410 83350
rect 97480 83150 97520 83350
rect 97590 83150 97910 83350
rect 97980 83150 98020 83350
rect 98090 83150 98410 83350
rect 98480 83150 98520 83350
rect 98590 83150 98910 83350
rect 98980 83150 99020 83350
rect 99090 83150 99410 83350
rect 99480 83150 99520 83350
rect 99590 83150 99910 83350
rect 99980 83150 100000 83350
rect 96000 83140 100000 83150
rect -15860 83090 -15640 83140
rect -15860 83020 -15850 83090
rect -15650 83020 -15640 83090
rect -15860 82980 -15640 83020
rect -15860 82910 -15850 82980
rect -15650 82910 -15640 82980
rect -15860 82860 -15640 82910
rect -15360 83090 -15140 83140
rect -15360 83020 -15350 83090
rect -15150 83020 -15140 83090
rect -15360 82980 -15140 83020
rect -15360 82910 -15350 82980
rect -15150 82910 -15140 82980
rect -15360 82860 -15140 82910
rect -14860 83090 -14640 83140
rect -14860 83020 -14850 83090
rect -14650 83020 -14640 83090
rect -14860 82980 -14640 83020
rect -14860 82910 -14850 82980
rect -14650 82910 -14640 82980
rect -14860 82860 -14640 82910
rect -14360 83090 -14140 83140
rect -14360 83020 -14350 83090
rect -14150 83020 -14140 83090
rect -14360 82980 -14140 83020
rect -14360 82910 -14350 82980
rect -14150 82910 -14140 82980
rect -14360 82860 -14140 82910
rect -13860 83090 -13640 83140
rect -13860 83020 -13850 83090
rect -13650 83020 -13640 83090
rect -13860 82980 -13640 83020
rect -13860 82910 -13850 82980
rect -13650 82910 -13640 82980
rect -13860 82860 -13640 82910
rect -13360 83090 -13140 83140
rect -13360 83020 -13350 83090
rect -13150 83020 -13140 83090
rect -13360 82980 -13140 83020
rect -13360 82910 -13350 82980
rect -13150 82910 -13140 82980
rect -13360 82860 -13140 82910
rect -12860 83090 -12640 83140
rect -12860 83020 -12850 83090
rect -12650 83020 -12640 83090
rect -12860 82980 -12640 83020
rect -12860 82910 -12850 82980
rect -12650 82910 -12640 82980
rect -12860 82860 -12640 82910
rect -12360 83090 -12140 83140
rect -12360 83020 -12350 83090
rect -12150 83020 -12140 83090
rect -12360 82980 -12140 83020
rect -12360 82910 -12350 82980
rect -12150 82910 -12140 82980
rect -12360 82860 -12140 82910
rect 96140 83090 96360 83140
rect 96140 83020 96150 83090
rect 96350 83020 96360 83090
rect 96140 82980 96360 83020
rect 96140 82910 96150 82980
rect 96350 82910 96360 82980
rect 96140 82860 96360 82910
rect 96640 83090 96860 83140
rect 96640 83020 96650 83090
rect 96850 83020 96860 83090
rect 96640 82980 96860 83020
rect 96640 82910 96650 82980
rect 96850 82910 96860 82980
rect 96640 82860 96860 82910
rect 97140 83090 97360 83140
rect 97140 83020 97150 83090
rect 97350 83020 97360 83090
rect 97140 82980 97360 83020
rect 97140 82910 97150 82980
rect 97350 82910 97360 82980
rect 97140 82860 97360 82910
rect 97640 83090 97860 83140
rect 97640 83020 97650 83090
rect 97850 83020 97860 83090
rect 97640 82980 97860 83020
rect 97640 82910 97650 82980
rect 97850 82910 97860 82980
rect 97640 82860 97860 82910
rect 98140 83090 98360 83140
rect 98140 83020 98150 83090
rect 98350 83020 98360 83090
rect 98140 82980 98360 83020
rect 98140 82910 98150 82980
rect 98350 82910 98360 82980
rect 98140 82860 98360 82910
rect 98640 83090 98860 83140
rect 98640 83020 98650 83090
rect 98850 83020 98860 83090
rect 98640 82980 98860 83020
rect 98640 82910 98650 82980
rect 98850 82910 98860 82980
rect 98640 82860 98860 82910
rect 99140 83090 99360 83140
rect 99140 83020 99150 83090
rect 99350 83020 99360 83090
rect 99140 82980 99360 83020
rect 99140 82910 99150 82980
rect 99350 82910 99360 82980
rect 99140 82860 99360 82910
rect 99640 83090 99860 83140
rect 99640 83020 99650 83090
rect 99850 83020 99860 83090
rect 99640 82980 99860 83020
rect 99640 82910 99650 82980
rect 99850 82910 99860 82980
rect 99640 82860 99860 82910
rect -16000 82850 -12000 82860
rect -16000 82650 -15980 82850
rect -15910 82650 -15590 82850
rect -15520 82650 -15480 82850
rect -15410 82650 -15090 82850
rect -15020 82650 -14980 82850
rect -14910 82650 -14590 82850
rect -14520 82650 -14480 82850
rect -14410 82650 -14090 82850
rect -14020 82650 -13980 82850
rect -13910 82650 -13590 82850
rect -13520 82650 -13480 82850
rect -13410 82650 -13090 82850
rect -13020 82650 -12980 82850
rect -12910 82650 -12590 82850
rect -12520 82650 -12480 82850
rect -12410 82650 -12090 82850
rect -12020 82650 -12000 82850
rect -16000 82640 -12000 82650
rect 96000 82850 100000 82860
rect 96000 82650 96020 82850
rect 96090 82650 96410 82850
rect 96480 82650 96520 82850
rect 96590 82650 96910 82850
rect 96980 82650 97020 82850
rect 97090 82650 97410 82850
rect 97480 82650 97520 82850
rect 97590 82650 97910 82850
rect 97980 82650 98020 82850
rect 98090 82650 98410 82850
rect 98480 82650 98520 82850
rect 98590 82650 98910 82850
rect 98980 82650 99020 82850
rect 99090 82650 99410 82850
rect 99480 82650 99520 82850
rect 99590 82650 99910 82850
rect 99980 82650 100000 82850
rect 96000 82640 100000 82650
rect -15860 82590 -15640 82640
rect -15860 82520 -15850 82590
rect -15650 82520 -15640 82590
rect -15860 82480 -15640 82520
rect -15860 82410 -15850 82480
rect -15650 82410 -15640 82480
rect -15860 82360 -15640 82410
rect -15360 82590 -15140 82640
rect -15360 82520 -15350 82590
rect -15150 82520 -15140 82590
rect -15360 82480 -15140 82520
rect -15360 82410 -15350 82480
rect -15150 82410 -15140 82480
rect -15360 82360 -15140 82410
rect -14860 82590 -14640 82640
rect -14860 82520 -14850 82590
rect -14650 82520 -14640 82590
rect -14860 82480 -14640 82520
rect -14860 82410 -14850 82480
rect -14650 82410 -14640 82480
rect -14860 82360 -14640 82410
rect -14360 82590 -14140 82640
rect -14360 82520 -14350 82590
rect -14150 82520 -14140 82590
rect -14360 82480 -14140 82520
rect -14360 82410 -14350 82480
rect -14150 82410 -14140 82480
rect -14360 82360 -14140 82410
rect -13860 82590 -13640 82640
rect -13860 82520 -13850 82590
rect -13650 82520 -13640 82590
rect -13860 82480 -13640 82520
rect -13860 82410 -13850 82480
rect -13650 82410 -13640 82480
rect -13860 82360 -13640 82410
rect -13360 82590 -13140 82640
rect -13360 82520 -13350 82590
rect -13150 82520 -13140 82590
rect -13360 82480 -13140 82520
rect -13360 82410 -13350 82480
rect -13150 82410 -13140 82480
rect -13360 82360 -13140 82410
rect -12860 82590 -12640 82640
rect -12860 82520 -12850 82590
rect -12650 82520 -12640 82590
rect -12860 82480 -12640 82520
rect -12860 82410 -12850 82480
rect -12650 82410 -12640 82480
rect -12860 82360 -12640 82410
rect -12360 82590 -12140 82640
rect -12360 82520 -12350 82590
rect -12150 82520 -12140 82590
rect -12360 82480 -12140 82520
rect -12360 82410 -12350 82480
rect -12150 82410 -12140 82480
rect -12360 82360 -12140 82410
rect 96140 82590 96360 82640
rect 96140 82520 96150 82590
rect 96350 82520 96360 82590
rect 96140 82480 96360 82520
rect 96140 82410 96150 82480
rect 96350 82410 96360 82480
rect 96140 82360 96360 82410
rect 96640 82590 96860 82640
rect 96640 82520 96650 82590
rect 96850 82520 96860 82590
rect 96640 82480 96860 82520
rect 96640 82410 96650 82480
rect 96850 82410 96860 82480
rect 96640 82360 96860 82410
rect 97140 82590 97360 82640
rect 97140 82520 97150 82590
rect 97350 82520 97360 82590
rect 97140 82480 97360 82520
rect 97140 82410 97150 82480
rect 97350 82410 97360 82480
rect 97140 82360 97360 82410
rect 97640 82590 97860 82640
rect 97640 82520 97650 82590
rect 97850 82520 97860 82590
rect 97640 82480 97860 82520
rect 97640 82410 97650 82480
rect 97850 82410 97860 82480
rect 97640 82360 97860 82410
rect 98140 82590 98360 82640
rect 98140 82520 98150 82590
rect 98350 82520 98360 82590
rect 98140 82480 98360 82520
rect 98140 82410 98150 82480
rect 98350 82410 98360 82480
rect 98140 82360 98360 82410
rect 98640 82590 98860 82640
rect 98640 82520 98650 82590
rect 98850 82520 98860 82590
rect 98640 82480 98860 82520
rect 98640 82410 98650 82480
rect 98850 82410 98860 82480
rect 98640 82360 98860 82410
rect 99140 82590 99360 82640
rect 99140 82520 99150 82590
rect 99350 82520 99360 82590
rect 99140 82480 99360 82520
rect 99140 82410 99150 82480
rect 99350 82410 99360 82480
rect 99140 82360 99360 82410
rect 99640 82590 99860 82640
rect 99640 82520 99650 82590
rect 99850 82520 99860 82590
rect 99640 82480 99860 82520
rect 99640 82410 99650 82480
rect 99850 82410 99860 82480
rect 99640 82360 99860 82410
rect -16000 82350 -12000 82360
rect -16000 82150 -15980 82350
rect -15910 82150 -15590 82350
rect -15520 82150 -15480 82350
rect -15410 82150 -15090 82350
rect -15020 82150 -14980 82350
rect -14910 82150 -14590 82350
rect -14520 82150 -14480 82350
rect -14410 82150 -14090 82350
rect -14020 82150 -13980 82350
rect -13910 82150 -13590 82350
rect -13520 82150 -13480 82350
rect -13410 82150 -13090 82350
rect -13020 82150 -12980 82350
rect -12910 82150 -12590 82350
rect -12520 82150 -12480 82350
rect -12410 82150 -12090 82350
rect -12020 82150 -12000 82350
rect -16000 82140 -12000 82150
rect 96000 82350 100000 82360
rect 96000 82150 96020 82350
rect 96090 82150 96410 82350
rect 96480 82150 96520 82350
rect 96590 82150 96910 82350
rect 96980 82150 97020 82350
rect 97090 82150 97410 82350
rect 97480 82150 97520 82350
rect 97590 82150 97910 82350
rect 97980 82150 98020 82350
rect 98090 82150 98410 82350
rect 98480 82150 98520 82350
rect 98590 82150 98910 82350
rect 98980 82150 99020 82350
rect 99090 82150 99410 82350
rect 99480 82150 99520 82350
rect 99590 82150 99910 82350
rect 99980 82150 100000 82350
rect 96000 82140 100000 82150
rect -15860 82090 -15640 82140
rect -15860 82020 -15850 82090
rect -15650 82020 -15640 82090
rect -15860 81980 -15640 82020
rect -15860 81910 -15850 81980
rect -15650 81910 -15640 81980
rect -15860 81860 -15640 81910
rect -15360 82090 -15140 82140
rect -15360 82020 -15350 82090
rect -15150 82020 -15140 82090
rect -15360 81980 -15140 82020
rect -15360 81910 -15350 81980
rect -15150 81910 -15140 81980
rect -15360 81860 -15140 81910
rect -14860 82090 -14640 82140
rect -14860 82020 -14850 82090
rect -14650 82020 -14640 82090
rect -14860 81980 -14640 82020
rect -14860 81910 -14850 81980
rect -14650 81910 -14640 81980
rect -14860 81860 -14640 81910
rect -14360 82090 -14140 82140
rect -14360 82020 -14350 82090
rect -14150 82020 -14140 82090
rect -14360 81980 -14140 82020
rect -14360 81910 -14350 81980
rect -14150 81910 -14140 81980
rect -14360 81860 -14140 81910
rect -13860 82090 -13640 82140
rect -13860 82020 -13850 82090
rect -13650 82020 -13640 82090
rect -13860 81980 -13640 82020
rect -13860 81910 -13850 81980
rect -13650 81910 -13640 81980
rect -13860 81860 -13640 81910
rect -13360 82090 -13140 82140
rect -13360 82020 -13350 82090
rect -13150 82020 -13140 82090
rect -13360 81980 -13140 82020
rect -13360 81910 -13350 81980
rect -13150 81910 -13140 81980
rect -13360 81860 -13140 81910
rect -12860 82090 -12640 82140
rect -12860 82020 -12850 82090
rect -12650 82020 -12640 82090
rect -12860 81980 -12640 82020
rect -12860 81910 -12850 81980
rect -12650 81910 -12640 81980
rect -12860 81860 -12640 81910
rect -12360 82090 -12140 82140
rect -12360 82020 -12350 82090
rect -12150 82020 -12140 82090
rect -12360 81980 -12140 82020
rect -12360 81910 -12350 81980
rect -12150 81910 -12140 81980
rect -12360 81860 -12140 81910
rect 96140 82090 96360 82140
rect 96140 82020 96150 82090
rect 96350 82020 96360 82090
rect 96140 81980 96360 82020
rect 96140 81910 96150 81980
rect 96350 81910 96360 81980
rect 96140 81860 96360 81910
rect 96640 82090 96860 82140
rect 96640 82020 96650 82090
rect 96850 82020 96860 82090
rect 96640 81980 96860 82020
rect 96640 81910 96650 81980
rect 96850 81910 96860 81980
rect 96640 81860 96860 81910
rect 97140 82090 97360 82140
rect 97140 82020 97150 82090
rect 97350 82020 97360 82090
rect 97140 81980 97360 82020
rect 97140 81910 97150 81980
rect 97350 81910 97360 81980
rect 97140 81860 97360 81910
rect 97640 82090 97860 82140
rect 97640 82020 97650 82090
rect 97850 82020 97860 82090
rect 97640 81980 97860 82020
rect 97640 81910 97650 81980
rect 97850 81910 97860 81980
rect 97640 81860 97860 81910
rect 98140 82090 98360 82140
rect 98140 82020 98150 82090
rect 98350 82020 98360 82090
rect 98140 81980 98360 82020
rect 98140 81910 98150 81980
rect 98350 81910 98360 81980
rect 98140 81860 98360 81910
rect 98640 82090 98860 82140
rect 98640 82020 98650 82090
rect 98850 82020 98860 82090
rect 98640 81980 98860 82020
rect 98640 81910 98650 81980
rect 98850 81910 98860 81980
rect 98640 81860 98860 81910
rect 99140 82090 99360 82140
rect 99140 82020 99150 82090
rect 99350 82020 99360 82090
rect 99140 81980 99360 82020
rect 99140 81910 99150 81980
rect 99350 81910 99360 81980
rect 99140 81860 99360 81910
rect 99640 82090 99860 82140
rect 99640 82020 99650 82090
rect 99850 82020 99860 82090
rect 99640 81980 99860 82020
rect 99640 81910 99650 81980
rect 99850 81910 99860 81980
rect 99640 81860 99860 81910
rect -16000 81850 -12000 81860
rect -16000 81650 -15980 81850
rect -15910 81650 -15590 81850
rect -15520 81650 -15480 81850
rect -15410 81650 -15090 81850
rect -15020 81650 -14980 81850
rect -14910 81650 -14590 81850
rect -14520 81650 -14480 81850
rect -14410 81650 -14090 81850
rect -14020 81650 -13980 81850
rect -13910 81650 -13590 81850
rect -13520 81650 -13480 81850
rect -13410 81650 -13090 81850
rect -13020 81650 -12980 81850
rect -12910 81650 -12590 81850
rect -12520 81650 -12480 81850
rect -12410 81650 -12090 81850
rect -12020 81650 -12000 81850
rect -16000 81640 -12000 81650
rect 96000 81850 100000 81860
rect 96000 81650 96020 81850
rect 96090 81650 96410 81850
rect 96480 81650 96520 81850
rect 96590 81650 96910 81850
rect 96980 81650 97020 81850
rect 97090 81650 97410 81850
rect 97480 81650 97520 81850
rect 97590 81650 97910 81850
rect 97980 81650 98020 81850
rect 98090 81650 98410 81850
rect 98480 81650 98520 81850
rect 98590 81650 98910 81850
rect 98980 81650 99020 81850
rect 99090 81650 99410 81850
rect 99480 81650 99520 81850
rect 99590 81650 99910 81850
rect 99980 81650 100000 81850
rect 96000 81640 100000 81650
rect -15860 81590 -15640 81640
rect -15860 81520 -15850 81590
rect -15650 81520 -15640 81590
rect -15860 81480 -15640 81520
rect -15860 81410 -15850 81480
rect -15650 81410 -15640 81480
rect -15860 81360 -15640 81410
rect -15360 81590 -15140 81640
rect -15360 81520 -15350 81590
rect -15150 81520 -15140 81590
rect -15360 81480 -15140 81520
rect -15360 81410 -15350 81480
rect -15150 81410 -15140 81480
rect -15360 81360 -15140 81410
rect -14860 81590 -14640 81640
rect -14860 81520 -14850 81590
rect -14650 81520 -14640 81590
rect -14860 81480 -14640 81520
rect -14860 81410 -14850 81480
rect -14650 81410 -14640 81480
rect -14860 81360 -14640 81410
rect -14360 81590 -14140 81640
rect -14360 81520 -14350 81590
rect -14150 81520 -14140 81590
rect -14360 81480 -14140 81520
rect -14360 81410 -14350 81480
rect -14150 81410 -14140 81480
rect -14360 81360 -14140 81410
rect -13860 81590 -13640 81640
rect -13860 81520 -13850 81590
rect -13650 81520 -13640 81590
rect -13860 81480 -13640 81520
rect -13860 81410 -13850 81480
rect -13650 81410 -13640 81480
rect -13860 81360 -13640 81410
rect -13360 81590 -13140 81640
rect -13360 81520 -13350 81590
rect -13150 81520 -13140 81590
rect -13360 81480 -13140 81520
rect -13360 81410 -13350 81480
rect -13150 81410 -13140 81480
rect -13360 81360 -13140 81410
rect -12860 81590 -12640 81640
rect -12860 81520 -12850 81590
rect -12650 81520 -12640 81590
rect -12860 81480 -12640 81520
rect -12860 81410 -12850 81480
rect -12650 81410 -12640 81480
rect -12860 81360 -12640 81410
rect -12360 81590 -12140 81640
rect -12360 81520 -12350 81590
rect -12150 81520 -12140 81590
rect -12360 81480 -12140 81520
rect -12360 81410 -12350 81480
rect -12150 81410 -12140 81480
rect -12360 81360 -12140 81410
rect 96140 81590 96360 81640
rect 96140 81520 96150 81590
rect 96350 81520 96360 81590
rect 96140 81480 96360 81520
rect 96140 81410 96150 81480
rect 96350 81410 96360 81480
rect 96140 81360 96360 81410
rect 96640 81590 96860 81640
rect 96640 81520 96650 81590
rect 96850 81520 96860 81590
rect 96640 81480 96860 81520
rect 96640 81410 96650 81480
rect 96850 81410 96860 81480
rect 96640 81360 96860 81410
rect 97140 81590 97360 81640
rect 97140 81520 97150 81590
rect 97350 81520 97360 81590
rect 97140 81480 97360 81520
rect 97140 81410 97150 81480
rect 97350 81410 97360 81480
rect 97140 81360 97360 81410
rect 97640 81590 97860 81640
rect 97640 81520 97650 81590
rect 97850 81520 97860 81590
rect 97640 81480 97860 81520
rect 97640 81410 97650 81480
rect 97850 81410 97860 81480
rect 97640 81360 97860 81410
rect 98140 81590 98360 81640
rect 98140 81520 98150 81590
rect 98350 81520 98360 81590
rect 98140 81480 98360 81520
rect 98140 81410 98150 81480
rect 98350 81410 98360 81480
rect 98140 81360 98360 81410
rect 98640 81590 98860 81640
rect 98640 81520 98650 81590
rect 98850 81520 98860 81590
rect 98640 81480 98860 81520
rect 98640 81410 98650 81480
rect 98850 81410 98860 81480
rect 98640 81360 98860 81410
rect 99140 81590 99360 81640
rect 99140 81520 99150 81590
rect 99350 81520 99360 81590
rect 99140 81480 99360 81520
rect 99140 81410 99150 81480
rect 99350 81410 99360 81480
rect 99140 81360 99360 81410
rect 99640 81590 99860 81640
rect 99640 81520 99650 81590
rect 99850 81520 99860 81590
rect 99640 81480 99860 81520
rect 99640 81410 99650 81480
rect 99850 81410 99860 81480
rect 99640 81360 99860 81410
rect -16000 81350 -12000 81360
rect -16000 81150 -15980 81350
rect -15910 81150 -15590 81350
rect -15520 81150 -15480 81350
rect -15410 81150 -15090 81350
rect -15020 81150 -14980 81350
rect -14910 81150 -14590 81350
rect -14520 81150 -14480 81350
rect -14410 81150 -14090 81350
rect -14020 81150 -13980 81350
rect -13910 81150 -13590 81350
rect -13520 81150 -13480 81350
rect -13410 81150 -13090 81350
rect -13020 81150 -12980 81350
rect -12910 81150 -12590 81350
rect -12520 81150 -12480 81350
rect -12410 81150 -12090 81350
rect -12020 81150 -12000 81350
rect -16000 81140 -12000 81150
rect 96000 81350 100000 81360
rect 96000 81150 96020 81350
rect 96090 81150 96410 81350
rect 96480 81150 96520 81350
rect 96590 81150 96910 81350
rect 96980 81150 97020 81350
rect 97090 81150 97410 81350
rect 97480 81150 97520 81350
rect 97590 81150 97910 81350
rect 97980 81150 98020 81350
rect 98090 81150 98410 81350
rect 98480 81150 98520 81350
rect 98590 81150 98910 81350
rect 98980 81150 99020 81350
rect 99090 81150 99410 81350
rect 99480 81150 99520 81350
rect 99590 81150 99910 81350
rect 99980 81150 100000 81350
rect 96000 81140 100000 81150
rect -15860 81090 -15640 81140
rect -15860 81020 -15850 81090
rect -15650 81020 -15640 81090
rect -15860 80980 -15640 81020
rect -15860 80910 -15850 80980
rect -15650 80910 -15640 80980
rect -15860 80860 -15640 80910
rect -15360 81090 -15140 81140
rect -15360 81020 -15350 81090
rect -15150 81020 -15140 81090
rect -15360 80980 -15140 81020
rect -15360 80910 -15350 80980
rect -15150 80910 -15140 80980
rect -15360 80860 -15140 80910
rect -14860 81090 -14640 81140
rect -14860 81020 -14850 81090
rect -14650 81020 -14640 81090
rect -14860 80980 -14640 81020
rect -14860 80910 -14850 80980
rect -14650 80910 -14640 80980
rect -14860 80860 -14640 80910
rect -14360 81090 -14140 81140
rect -14360 81020 -14350 81090
rect -14150 81020 -14140 81090
rect -14360 80980 -14140 81020
rect -14360 80910 -14350 80980
rect -14150 80910 -14140 80980
rect -14360 80860 -14140 80910
rect -13860 81090 -13640 81140
rect -13860 81020 -13850 81090
rect -13650 81020 -13640 81090
rect -13860 80980 -13640 81020
rect -13860 80910 -13850 80980
rect -13650 80910 -13640 80980
rect -13860 80860 -13640 80910
rect -13360 81090 -13140 81140
rect -13360 81020 -13350 81090
rect -13150 81020 -13140 81090
rect -13360 80980 -13140 81020
rect -13360 80910 -13350 80980
rect -13150 80910 -13140 80980
rect -13360 80860 -13140 80910
rect -12860 81090 -12640 81140
rect -12860 81020 -12850 81090
rect -12650 81020 -12640 81090
rect -12860 80980 -12640 81020
rect -12860 80910 -12850 80980
rect -12650 80910 -12640 80980
rect -12860 80860 -12640 80910
rect -12360 81090 -12140 81140
rect -12360 81020 -12350 81090
rect -12150 81020 -12140 81090
rect -12360 80980 -12140 81020
rect -12360 80910 -12350 80980
rect -12150 80910 -12140 80980
rect -12360 80860 -12140 80910
rect 96140 81090 96360 81140
rect 96140 81020 96150 81090
rect 96350 81020 96360 81090
rect 96140 80980 96360 81020
rect 96140 80910 96150 80980
rect 96350 80910 96360 80980
rect 96140 80860 96360 80910
rect 96640 81090 96860 81140
rect 96640 81020 96650 81090
rect 96850 81020 96860 81090
rect 96640 80980 96860 81020
rect 96640 80910 96650 80980
rect 96850 80910 96860 80980
rect 96640 80860 96860 80910
rect 97140 81090 97360 81140
rect 97140 81020 97150 81090
rect 97350 81020 97360 81090
rect 97140 80980 97360 81020
rect 97140 80910 97150 80980
rect 97350 80910 97360 80980
rect 97140 80860 97360 80910
rect 97640 81090 97860 81140
rect 97640 81020 97650 81090
rect 97850 81020 97860 81090
rect 97640 80980 97860 81020
rect 97640 80910 97650 80980
rect 97850 80910 97860 80980
rect 97640 80860 97860 80910
rect 98140 81090 98360 81140
rect 98140 81020 98150 81090
rect 98350 81020 98360 81090
rect 98140 80980 98360 81020
rect 98140 80910 98150 80980
rect 98350 80910 98360 80980
rect 98140 80860 98360 80910
rect 98640 81090 98860 81140
rect 98640 81020 98650 81090
rect 98850 81020 98860 81090
rect 98640 80980 98860 81020
rect 98640 80910 98650 80980
rect 98850 80910 98860 80980
rect 98640 80860 98860 80910
rect 99140 81090 99360 81140
rect 99140 81020 99150 81090
rect 99350 81020 99360 81090
rect 99140 80980 99360 81020
rect 99140 80910 99150 80980
rect 99350 80910 99360 80980
rect 99140 80860 99360 80910
rect 99640 81090 99860 81140
rect 99640 81020 99650 81090
rect 99850 81020 99860 81090
rect 99640 80980 99860 81020
rect 99640 80910 99650 80980
rect 99850 80910 99860 80980
rect 99640 80860 99860 80910
rect -16000 80850 -12000 80860
rect -16000 80650 -15980 80850
rect -15910 80650 -15590 80850
rect -15520 80650 -15480 80850
rect -15410 80650 -15090 80850
rect -15020 80650 -14980 80850
rect -14910 80650 -14590 80850
rect -14520 80650 -14480 80850
rect -14410 80650 -14090 80850
rect -14020 80650 -13980 80850
rect -13910 80650 -13590 80850
rect -13520 80650 -13480 80850
rect -13410 80650 -13090 80850
rect -13020 80650 -12980 80850
rect -12910 80650 -12590 80850
rect -12520 80650 -12480 80850
rect -12410 80650 -12090 80850
rect -12020 80650 -12000 80850
rect -16000 80640 -12000 80650
rect 96000 80850 100000 80860
rect 96000 80650 96020 80850
rect 96090 80650 96410 80850
rect 96480 80650 96520 80850
rect 96590 80650 96910 80850
rect 96980 80650 97020 80850
rect 97090 80650 97410 80850
rect 97480 80650 97520 80850
rect 97590 80650 97910 80850
rect 97980 80650 98020 80850
rect 98090 80650 98410 80850
rect 98480 80650 98520 80850
rect 98590 80650 98910 80850
rect 98980 80650 99020 80850
rect 99090 80650 99410 80850
rect 99480 80650 99520 80850
rect 99590 80650 99910 80850
rect 99980 80650 100000 80850
rect 96000 80640 100000 80650
rect -15860 80590 -15640 80640
rect -15860 80520 -15850 80590
rect -15650 80520 -15640 80590
rect -15860 80480 -15640 80520
rect -15860 80410 -15850 80480
rect -15650 80410 -15640 80480
rect -15860 80360 -15640 80410
rect -15360 80590 -15140 80640
rect -15360 80520 -15350 80590
rect -15150 80520 -15140 80590
rect -15360 80480 -15140 80520
rect -15360 80410 -15350 80480
rect -15150 80410 -15140 80480
rect -15360 80360 -15140 80410
rect -14860 80590 -14640 80640
rect -14860 80520 -14850 80590
rect -14650 80520 -14640 80590
rect -14860 80480 -14640 80520
rect -14860 80410 -14850 80480
rect -14650 80410 -14640 80480
rect -14860 80360 -14640 80410
rect -14360 80590 -14140 80640
rect -14360 80520 -14350 80590
rect -14150 80520 -14140 80590
rect -14360 80480 -14140 80520
rect -14360 80410 -14350 80480
rect -14150 80410 -14140 80480
rect -14360 80360 -14140 80410
rect -13860 80590 -13640 80640
rect -13860 80520 -13850 80590
rect -13650 80520 -13640 80590
rect -13860 80480 -13640 80520
rect -13860 80410 -13850 80480
rect -13650 80410 -13640 80480
rect -13860 80360 -13640 80410
rect -13360 80590 -13140 80640
rect -13360 80520 -13350 80590
rect -13150 80520 -13140 80590
rect -13360 80480 -13140 80520
rect -13360 80410 -13350 80480
rect -13150 80410 -13140 80480
rect -13360 80360 -13140 80410
rect -12860 80590 -12640 80640
rect -12860 80520 -12850 80590
rect -12650 80520 -12640 80590
rect -12860 80480 -12640 80520
rect -12860 80410 -12850 80480
rect -12650 80410 -12640 80480
rect -12860 80360 -12640 80410
rect -12360 80590 -12140 80640
rect -12360 80520 -12350 80590
rect -12150 80520 -12140 80590
rect -12360 80480 -12140 80520
rect -12360 80410 -12350 80480
rect -12150 80410 -12140 80480
rect -12360 80360 -12140 80410
rect 96140 80590 96360 80640
rect 96140 80520 96150 80590
rect 96350 80520 96360 80590
rect 96140 80480 96360 80520
rect 96140 80410 96150 80480
rect 96350 80410 96360 80480
rect 96140 80360 96360 80410
rect 96640 80590 96860 80640
rect 96640 80520 96650 80590
rect 96850 80520 96860 80590
rect 96640 80480 96860 80520
rect 96640 80410 96650 80480
rect 96850 80410 96860 80480
rect 96640 80360 96860 80410
rect 97140 80590 97360 80640
rect 97140 80520 97150 80590
rect 97350 80520 97360 80590
rect 97140 80480 97360 80520
rect 97140 80410 97150 80480
rect 97350 80410 97360 80480
rect 97140 80360 97360 80410
rect 97640 80590 97860 80640
rect 97640 80520 97650 80590
rect 97850 80520 97860 80590
rect 97640 80480 97860 80520
rect 97640 80410 97650 80480
rect 97850 80410 97860 80480
rect 97640 80360 97860 80410
rect 98140 80590 98360 80640
rect 98140 80520 98150 80590
rect 98350 80520 98360 80590
rect 98140 80480 98360 80520
rect 98140 80410 98150 80480
rect 98350 80410 98360 80480
rect 98140 80360 98360 80410
rect 98640 80590 98860 80640
rect 98640 80520 98650 80590
rect 98850 80520 98860 80590
rect 98640 80480 98860 80520
rect 98640 80410 98650 80480
rect 98850 80410 98860 80480
rect 98640 80360 98860 80410
rect 99140 80590 99360 80640
rect 99140 80520 99150 80590
rect 99350 80520 99360 80590
rect 99140 80480 99360 80520
rect 99140 80410 99150 80480
rect 99350 80410 99360 80480
rect 99140 80360 99360 80410
rect 99640 80590 99860 80640
rect 99640 80520 99650 80590
rect 99850 80520 99860 80590
rect 99640 80480 99860 80520
rect 99640 80410 99650 80480
rect 99850 80410 99860 80480
rect 99640 80360 99860 80410
rect -16000 80350 -12000 80360
rect -16000 80150 -15980 80350
rect -15910 80150 -15590 80350
rect -15520 80150 -15480 80350
rect -15410 80150 -15090 80350
rect -15020 80150 -14980 80350
rect -14910 80150 -14590 80350
rect -14520 80150 -14480 80350
rect -14410 80150 -14090 80350
rect -14020 80150 -13980 80350
rect -13910 80150 -13590 80350
rect -13520 80150 -13480 80350
rect -13410 80150 -13090 80350
rect -13020 80150 -12980 80350
rect -12910 80150 -12590 80350
rect -12520 80150 -12480 80350
rect -12410 80150 -12090 80350
rect -12020 80150 -12000 80350
rect -16000 80140 -12000 80150
rect 96000 80350 100000 80360
rect 96000 80150 96020 80350
rect 96090 80150 96410 80350
rect 96480 80150 96520 80350
rect 96590 80150 96910 80350
rect 96980 80150 97020 80350
rect 97090 80150 97410 80350
rect 97480 80150 97520 80350
rect 97590 80150 97910 80350
rect 97980 80150 98020 80350
rect 98090 80150 98410 80350
rect 98480 80150 98520 80350
rect 98590 80150 98910 80350
rect 98980 80150 99020 80350
rect 99090 80150 99410 80350
rect 99480 80150 99520 80350
rect 99590 80150 99910 80350
rect 99980 80150 100000 80350
rect 96000 80140 100000 80150
rect -15860 80090 -15640 80140
rect -15860 80020 -15850 80090
rect -15650 80020 -15640 80090
rect -15860 79980 -15640 80020
rect -15860 79910 -15850 79980
rect -15650 79910 -15640 79980
rect -15860 79860 -15640 79910
rect -15360 80090 -15140 80140
rect -15360 80020 -15350 80090
rect -15150 80020 -15140 80090
rect -15360 79980 -15140 80020
rect -15360 79910 -15350 79980
rect -15150 79910 -15140 79980
rect -15360 79860 -15140 79910
rect -14860 80090 -14640 80140
rect -14860 80020 -14850 80090
rect -14650 80020 -14640 80090
rect -14860 79980 -14640 80020
rect -14860 79910 -14850 79980
rect -14650 79910 -14640 79980
rect -14860 79860 -14640 79910
rect -14360 80090 -14140 80140
rect -14360 80020 -14350 80090
rect -14150 80020 -14140 80090
rect -14360 79980 -14140 80020
rect -14360 79910 -14350 79980
rect -14150 79910 -14140 79980
rect -14360 79860 -14140 79910
rect -13860 80090 -13640 80140
rect -13860 80020 -13850 80090
rect -13650 80020 -13640 80090
rect -13860 79980 -13640 80020
rect -13860 79910 -13850 79980
rect -13650 79910 -13640 79980
rect -13860 79860 -13640 79910
rect -13360 80090 -13140 80140
rect -13360 80020 -13350 80090
rect -13150 80020 -13140 80090
rect -13360 79980 -13140 80020
rect -13360 79910 -13350 79980
rect -13150 79910 -13140 79980
rect -13360 79860 -13140 79910
rect -12860 80090 -12640 80140
rect -12860 80020 -12850 80090
rect -12650 80020 -12640 80090
rect -12860 79980 -12640 80020
rect -12860 79910 -12850 79980
rect -12650 79910 -12640 79980
rect -12860 79860 -12640 79910
rect -12360 80090 -12140 80140
rect -12360 80020 -12350 80090
rect -12150 80020 -12140 80090
rect -12360 79980 -12140 80020
rect -12360 79910 -12350 79980
rect -12150 79910 -12140 79980
rect -12360 79860 -12140 79910
rect 96140 80090 96360 80140
rect 96140 80020 96150 80090
rect 96350 80020 96360 80090
rect 96140 79980 96360 80020
rect 96140 79910 96150 79980
rect 96350 79910 96360 79980
rect 96140 79860 96360 79910
rect 96640 80090 96860 80140
rect 96640 80020 96650 80090
rect 96850 80020 96860 80090
rect 96640 79980 96860 80020
rect 96640 79910 96650 79980
rect 96850 79910 96860 79980
rect 96640 79860 96860 79910
rect 97140 80090 97360 80140
rect 97140 80020 97150 80090
rect 97350 80020 97360 80090
rect 97140 79980 97360 80020
rect 97140 79910 97150 79980
rect 97350 79910 97360 79980
rect 97140 79860 97360 79910
rect 97640 80090 97860 80140
rect 97640 80020 97650 80090
rect 97850 80020 97860 80090
rect 97640 79980 97860 80020
rect 97640 79910 97650 79980
rect 97850 79910 97860 79980
rect 97640 79860 97860 79910
rect 98140 80090 98360 80140
rect 98140 80020 98150 80090
rect 98350 80020 98360 80090
rect 98140 79980 98360 80020
rect 98140 79910 98150 79980
rect 98350 79910 98360 79980
rect 98140 79860 98360 79910
rect 98640 80090 98860 80140
rect 98640 80020 98650 80090
rect 98850 80020 98860 80090
rect 98640 79980 98860 80020
rect 98640 79910 98650 79980
rect 98850 79910 98860 79980
rect 98640 79860 98860 79910
rect 99140 80090 99360 80140
rect 99140 80020 99150 80090
rect 99350 80020 99360 80090
rect 99140 79980 99360 80020
rect 99140 79910 99150 79980
rect 99350 79910 99360 79980
rect 99140 79860 99360 79910
rect 99640 80090 99860 80140
rect 99640 80020 99650 80090
rect 99850 80020 99860 80090
rect 99640 79980 99860 80020
rect 99640 79910 99650 79980
rect 99850 79910 99860 79980
rect 99640 79860 99860 79910
rect -16000 79850 -12000 79860
rect -16000 79650 -15980 79850
rect -15910 79650 -15590 79850
rect -15520 79650 -15480 79850
rect -15410 79650 -15090 79850
rect -15020 79650 -14980 79850
rect -14910 79650 -14590 79850
rect -14520 79650 -14480 79850
rect -14410 79650 -14090 79850
rect -14020 79650 -13980 79850
rect -13910 79650 -13590 79850
rect -13520 79650 -13480 79850
rect -13410 79650 -13090 79850
rect -13020 79650 -12980 79850
rect -12910 79650 -12590 79850
rect -12520 79650 -12480 79850
rect -12410 79650 -12090 79850
rect -12020 79650 -12000 79850
rect -16000 79640 -12000 79650
rect 96000 79850 100000 79860
rect 96000 79650 96020 79850
rect 96090 79650 96410 79850
rect 96480 79650 96520 79850
rect 96590 79650 96910 79850
rect 96980 79650 97020 79850
rect 97090 79650 97410 79850
rect 97480 79650 97520 79850
rect 97590 79650 97910 79850
rect 97980 79650 98020 79850
rect 98090 79650 98410 79850
rect 98480 79650 98520 79850
rect 98590 79650 98910 79850
rect 98980 79650 99020 79850
rect 99090 79650 99410 79850
rect 99480 79650 99520 79850
rect 99590 79650 99910 79850
rect 99980 79650 100000 79850
rect 96000 79640 100000 79650
rect -15860 79590 -15640 79640
rect -15860 79520 -15850 79590
rect -15650 79520 -15640 79590
rect -15860 79480 -15640 79520
rect -15860 79410 -15850 79480
rect -15650 79410 -15640 79480
rect -15860 79360 -15640 79410
rect -15360 79590 -15140 79640
rect -15360 79520 -15350 79590
rect -15150 79520 -15140 79590
rect -15360 79480 -15140 79520
rect -15360 79410 -15350 79480
rect -15150 79410 -15140 79480
rect -15360 79360 -15140 79410
rect -14860 79590 -14640 79640
rect -14860 79520 -14850 79590
rect -14650 79520 -14640 79590
rect -14860 79480 -14640 79520
rect -14860 79410 -14850 79480
rect -14650 79410 -14640 79480
rect -14860 79360 -14640 79410
rect -14360 79590 -14140 79640
rect -14360 79520 -14350 79590
rect -14150 79520 -14140 79590
rect -14360 79480 -14140 79520
rect -14360 79410 -14350 79480
rect -14150 79410 -14140 79480
rect -14360 79360 -14140 79410
rect -13860 79590 -13640 79640
rect -13860 79520 -13850 79590
rect -13650 79520 -13640 79590
rect -13860 79480 -13640 79520
rect -13860 79410 -13850 79480
rect -13650 79410 -13640 79480
rect -13860 79360 -13640 79410
rect -13360 79590 -13140 79640
rect -13360 79520 -13350 79590
rect -13150 79520 -13140 79590
rect -13360 79480 -13140 79520
rect -13360 79410 -13350 79480
rect -13150 79410 -13140 79480
rect -13360 79360 -13140 79410
rect -12860 79590 -12640 79640
rect -12860 79520 -12850 79590
rect -12650 79520 -12640 79590
rect -12860 79480 -12640 79520
rect -12860 79410 -12850 79480
rect -12650 79410 -12640 79480
rect -12860 79360 -12640 79410
rect -12360 79590 -12140 79640
rect -12360 79520 -12350 79590
rect -12150 79520 -12140 79590
rect -12360 79480 -12140 79520
rect -12360 79410 -12350 79480
rect -12150 79410 -12140 79480
rect -12360 79360 -12140 79410
rect 96140 79590 96360 79640
rect 96140 79520 96150 79590
rect 96350 79520 96360 79590
rect 96140 79480 96360 79520
rect 96140 79410 96150 79480
rect 96350 79410 96360 79480
rect 96140 79360 96360 79410
rect 96640 79590 96860 79640
rect 96640 79520 96650 79590
rect 96850 79520 96860 79590
rect 96640 79480 96860 79520
rect 96640 79410 96650 79480
rect 96850 79410 96860 79480
rect 96640 79360 96860 79410
rect 97140 79590 97360 79640
rect 97140 79520 97150 79590
rect 97350 79520 97360 79590
rect 97140 79480 97360 79520
rect 97140 79410 97150 79480
rect 97350 79410 97360 79480
rect 97140 79360 97360 79410
rect 97640 79590 97860 79640
rect 97640 79520 97650 79590
rect 97850 79520 97860 79590
rect 97640 79480 97860 79520
rect 97640 79410 97650 79480
rect 97850 79410 97860 79480
rect 97640 79360 97860 79410
rect 98140 79590 98360 79640
rect 98140 79520 98150 79590
rect 98350 79520 98360 79590
rect 98140 79480 98360 79520
rect 98140 79410 98150 79480
rect 98350 79410 98360 79480
rect 98140 79360 98360 79410
rect 98640 79590 98860 79640
rect 98640 79520 98650 79590
rect 98850 79520 98860 79590
rect 98640 79480 98860 79520
rect 98640 79410 98650 79480
rect 98850 79410 98860 79480
rect 98640 79360 98860 79410
rect 99140 79590 99360 79640
rect 99140 79520 99150 79590
rect 99350 79520 99360 79590
rect 99140 79480 99360 79520
rect 99140 79410 99150 79480
rect 99350 79410 99360 79480
rect 99140 79360 99360 79410
rect 99640 79590 99860 79640
rect 99640 79520 99650 79590
rect 99850 79520 99860 79590
rect 99640 79480 99860 79520
rect 99640 79410 99650 79480
rect 99850 79410 99860 79480
rect 99640 79360 99860 79410
rect -16000 79350 -12000 79360
rect -16000 79150 -15980 79350
rect -15910 79150 -15590 79350
rect -15520 79150 -15480 79350
rect -15410 79150 -15090 79350
rect -15020 79150 -14980 79350
rect -14910 79150 -14590 79350
rect -14520 79150 -14480 79350
rect -14410 79150 -14090 79350
rect -14020 79150 -13980 79350
rect -13910 79150 -13590 79350
rect -13520 79150 -13480 79350
rect -13410 79150 -13090 79350
rect -13020 79150 -12980 79350
rect -12910 79150 -12590 79350
rect -12520 79150 -12480 79350
rect -12410 79150 -12090 79350
rect -12020 79150 -12000 79350
rect -16000 79140 -12000 79150
rect 96000 79350 100000 79360
rect 96000 79150 96020 79350
rect 96090 79150 96410 79350
rect 96480 79150 96520 79350
rect 96590 79150 96910 79350
rect 96980 79150 97020 79350
rect 97090 79150 97410 79350
rect 97480 79150 97520 79350
rect 97590 79150 97910 79350
rect 97980 79150 98020 79350
rect 98090 79150 98410 79350
rect 98480 79150 98520 79350
rect 98590 79150 98910 79350
rect 98980 79150 99020 79350
rect 99090 79150 99410 79350
rect 99480 79150 99520 79350
rect 99590 79150 99910 79350
rect 99980 79150 100000 79350
rect 96000 79140 100000 79150
rect -15860 79090 -15640 79140
rect -15860 79020 -15850 79090
rect -15650 79020 -15640 79090
rect -15860 78980 -15640 79020
rect -15860 78910 -15850 78980
rect -15650 78910 -15640 78980
rect -15860 78860 -15640 78910
rect -15360 79090 -15140 79140
rect -15360 79020 -15350 79090
rect -15150 79020 -15140 79090
rect -15360 78980 -15140 79020
rect -15360 78910 -15350 78980
rect -15150 78910 -15140 78980
rect -15360 78860 -15140 78910
rect -14860 79090 -14640 79140
rect -14860 79020 -14850 79090
rect -14650 79020 -14640 79090
rect -14860 78980 -14640 79020
rect -14860 78910 -14850 78980
rect -14650 78910 -14640 78980
rect -14860 78860 -14640 78910
rect -14360 79090 -14140 79140
rect -14360 79020 -14350 79090
rect -14150 79020 -14140 79090
rect -14360 78980 -14140 79020
rect -14360 78910 -14350 78980
rect -14150 78910 -14140 78980
rect -14360 78860 -14140 78910
rect -13860 79090 -13640 79140
rect -13860 79020 -13850 79090
rect -13650 79020 -13640 79090
rect -13860 78980 -13640 79020
rect -13860 78910 -13850 78980
rect -13650 78910 -13640 78980
rect -13860 78860 -13640 78910
rect -13360 79090 -13140 79140
rect -13360 79020 -13350 79090
rect -13150 79020 -13140 79090
rect -13360 78980 -13140 79020
rect -13360 78910 -13350 78980
rect -13150 78910 -13140 78980
rect -13360 78860 -13140 78910
rect -12860 79090 -12640 79140
rect -12860 79020 -12850 79090
rect -12650 79020 -12640 79090
rect -12860 78980 -12640 79020
rect -12860 78910 -12850 78980
rect -12650 78910 -12640 78980
rect -12860 78860 -12640 78910
rect -12360 79090 -12140 79140
rect -12360 79020 -12350 79090
rect -12150 79020 -12140 79090
rect -12360 78980 -12140 79020
rect -12360 78910 -12350 78980
rect -12150 78910 -12140 78980
rect -12360 78860 -12140 78910
rect 96140 79090 96360 79140
rect 96140 79020 96150 79090
rect 96350 79020 96360 79090
rect 96140 78980 96360 79020
rect 96140 78910 96150 78980
rect 96350 78910 96360 78980
rect 96140 78860 96360 78910
rect 96640 79090 96860 79140
rect 96640 79020 96650 79090
rect 96850 79020 96860 79090
rect 96640 78980 96860 79020
rect 96640 78910 96650 78980
rect 96850 78910 96860 78980
rect 96640 78860 96860 78910
rect 97140 79090 97360 79140
rect 97140 79020 97150 79090
rect 97350 79020 97360 79090
rect 97140 78980 97360 79020
rect 97140 78910 97150 78980
rect 97350 78910 97360 78980
rect 97140 78860 97360 78910
rect 97640 79090 97860 79140
rect 97640 79020 97650 79090
rect 97850 79020 97860 79090
rect 97640 78980 97860 79020
rect 97640 78910 97650 78980
rect 97850 78910 97860 78980
rect 97640 78860 97860 78910
rect 98140 79090 98360 79140
rect 98140 79020 98150 79090
rect 98350 79020 98360 79090
rect 98140 78980 98360 79020
rect 98140 78910 98150 78980
rect 98350 78910 98360 78980
rect 98140 78860 98360 78910
rect 98640 79090 98860 79140
rect 98640 79020 98650 79090
rect 98850 79020 98860 79090
rect 98640 78980 98860 79020
rect 98640 78910 98650 78980
rect 98850 78910 98860 78980
rect 98640 78860 98860 78910
rect 99140 79090 99360 79140
rect 99140 79020 99150 79090
rect 99350 79020 99360 79090
rect 99140 78980 99360 79020
rect 99140 78910 99150 78980
rect 99350 78910 99360 78980
rect 99140 78860 99360 78910
rect 99640 79090 99860 79140
rect 99640 79020 99650 79090
rect 99850 79020 99860 79090
rect 99640 78980 99860 79020
rect 99640 78910 99650 78980
rect 99850 78910 99860 78980
rect 99640 78860 99860 78910
rect -16000 78850 -12000 78860
rect -16000 78650 -15980 78850
rect -15910 78650 -15590 78850
rect -15520 78650 -15480 78850
rect -15410 78650 -15090 78850
rect -15020 78650 -14980 78850
rect -14910 78650 -14590 78850
rect -14520 78650 -14480 78850
rect -14410 78650 -14090 78850
rect -14020 78650 -13980 78850
rect -13910 78650 -13590 78850
rect -13520 78650 -13480 78850
rect -13410 78650 -13090 78850
rect -13020 78650 -12980 78850
rect -12910 78650 -12590 78850
rect -12520 78650 -12480 78850
rect -12410 78650 -12090 78850
rect -12020 78650 -12000 78850
rect -16000 78640 -12000 78650
rect 96000 78850 100000 78860
rect 96000 78650 96020 78850
rect 96090 78650 96410 78850
rect 96480 78650 96520 78850
rect 96590 78650 96910 78850
rect 96980 78650 97020 78850
rect 97090 78650 97410 78850
rect 97480 78650 97520 78850
rect 97590 78650 97910 78850
rect 97980 78650 98020 78850
rect 98090 78650 98410 78850
rect 98480 78650 98520 78850
rect 98590 78650 98910 78850
rect 98980 78650 99020 78850
rect 99090 78650 99410 78850
rect 99480 78650 99520 78850
rect 99590 78650 99910 78850
rect 99980 78650 100000 78850
rect 96000 78640 100000 78650
rect -15860 78590 -15640 78640
rect -15860 78520 -15850 78590
rect -15650 78520 -15640 78590
rect -15860 78480 -15640 78520
rect -15860 78410 -15850 78480
rect -15650 78410 -15640 78480
rect -15860 78360 -15640 78410
rect -15360 78590 -15140 78640
rect -15360 78520 -15350 78590
rect -15150 78520 -15140 78590
rect -15360 78480 -15140 78520
rect -15360 78410 -15350 78480
rect -15150 78410 -15140 78480
rect -15360 78360 -15140 78410
rect -14860 78590 -14640 78640
rect -14860 78520 -14850 78590
rect -14650 78520 -14640 78590
rect -14860 78480 -14640 78520
rect -14860 78410 -14850 78480
rect -14650 78410 -14640 78480
rect -14860 78360 -14640 78410
rect -14360 78590 -14140 78640
rect -14360 78520 -14350 78590
rect -14150 78520 -14140 78590
rect -14360 78480 -14140 78520
rect -14360 78410 -14350 78480
rect -14150 78410 -14140 78480
rect -14360 78360 -14140 78410
rect -13860 78590 -13640 78640
rect -13860 78520 -13850 78590
rect -13650 78520 -13640 78590
rect -13860 78480 -13640 78520
rect -13860 78410 -13850 78480
rect -13650 78410 -13640 78480
rect -13860 78360 -13640 78410
rect -13360 78590 -13140 78640
rect -13360 78520 -13350 78590
rect -13150 78520 -13140 78590
rect -13360 78480 -13140 78520
rect -13360 78410 -13350 78480
rect -13150 78410 -13140 78480
rect -13360 78360 -13140 78410
rect -12860 78590 -12640 78640
rect -12860 78520 -12850 78590
rect -12650 78520 -12640 78590
rect -12860 78480 -12640 78520
rect -12860 78410 -12850 78480
rect -12650 78410 -12640 78480
rect -12860 78360 -12640 78410
rect -12360 78590 -12140 78640
rect -12360 78520 -12350 78590
rect -12150 78520 -12140 78590
rect -12360 78480 -12140 78520
rect -12360 78410 -12350 78480
rect -12150 78410 -12140 78480
rect -12360 78360 -12140 78410
rect 96140 78590 96360 78640
rect 96140 78520 96150 78590
rect 96350 78520 96360 78590
rect 96140 78480 96360 78520
rect 96140 78410 96150 78480
rect 96350 78410 96360 78480
rect 96140 78360 96360 78410
rect 96640 78590 96860 78640
rect 96640 78520 96650 78590
rect 96850 78520 96860 78590
rect 96640 78480 96860 78520
rect 96640 78410 96650 78480
rect 96850 78410 96860 78480
rect 96640 78360 96860 78410
rect 97140 78590 97360 78640
rect 97140 78520 97150 78590
rect 97350 78520 97360 78590
rect 97140 78480 97360 78520
rect 97140 78410 97150 78480
rect 97350 78410 97360 78480
rect 97140 78360 97360 78410
rect 97640 78590 97860 78640
rect 97640 78520 97650 78590
rect 97850 78520 97860 78590
rect 97640 78480 97860 78520
rect 97640 78410 97650 78480
rect 97850 78410 97860 78480
rect 97640 78360 97860 78410
rect 98140 78590 98360 78640
rect 98140 78520 98150 78590
rect 98350 78520 98360 78590
rect 98140 78480 98360 78520
rect 98140 78410 98150 78480
rect 98350 78410 98360 78480
rect 98140 78360 98360 78410
rect 98640 78590 98860 78640
rect 98640 78520 98650 78590
rect 98850 78520 98860 78590
rect 98640 78480 98860 78520
rect 98640 78410 98650 78480
rect 98850 78410 98860 78480
rect 98640 78360 98860 78410
rect 99140 78590 99360 78640
rect 99140 78520 99150 78590
rect 99350 78520 99360 78590
rect 99140 78480 99360 78520
rect 99140 78410 99150 78480
rect 99350 78410 99360 78480
rect 99140 78360 99360 78410
rect 99640 78590 99860 78640
rect 99640 78520 99650 78590
rect 99850 78520 99860 78590
rect 99640 78480 99860 78520
rect 99640 78410 99650 78480
rect 99850 78410 99860 78480
rect 99640 78360 99860 78410
rect -16000 78350 -12000 78360
rect -16000 78150 -15980 78350
rect -15910 78150 -15590 78350
rect -15520 78150 -15480 78350
rect -15410 78150 -15090 78350
rect -15020 78150 -14980 78350
rect -14910 78150 -14590 78350
rect -14520 78150 -14480 78350
rect -14410 78150 -14090 78350
rect -14020 78150 -13980 78350
rect -13910 78150 -13590 78350
rect -13520 78150 -13480 78350
rect -13410 78150 -13090 78350
rect -13020 78150 -12980 78350
rect -12910 78150 -12590 78350
rect -12520 78150 -12480 78350
rect -12410 78150 -12090 78350
rect -12020 78150 -12000 78350
rect -16000 78140 -12000 78150
rect 96000 78350 100000 78360
rect 96000 78150 96020 78350
rect 96090 78150 96410 78350
rect 96480 78150 96520 78350
rect 96590 78150 96910 78350
rect 96980 78150 97020 78350
rect 97090 78150 97410 78350
rect 97480 78150 97520 78350
rect 97590 78150 97910 78350
rect 97980 78150 98020 78350
rect 98090 78150 98410 78350
rect 98480 78150 98520 78350
rect 98590 78150 98910 78350
rect 98980 78150 99020 78350
rect 99090 78150 99410 78350
rect 99480 78150 99520 78350
rect 99590 78150 99910 78350
rect 99980 78150 100000 78350
rect 96000 78140 100000 78150
rect -15860 78090 -15640 78140
rect -15860 78020 -15850 78090
rect -15650 78020 -15640 78090
rect -15860 77980 -15640 78020
rect -15860 77910 -15850 77980
rect -15650 77910 -15640 77980
rect -15860 77860 -15640 77910
rect -15360 78090 -15140 78140
rect -15360 78020 -15350 78090
rect -15150 78020 -15140 78090
rect -15360 77980 -15140 78020
rect -15360 77910 -15350 77980
rect -15150 77910 -15140 77980
rect -15360 77860 -15140 77910
rect -14860 78090 -14640 78140
rect -14860 78020 -14850 78090
rect -14650 78020 -14640 78090
rect -14860 77980 -14640 78020
rect -14860 77910 -14850 77980
rect -14650 77910 -14640 77980
rect -14860 77860 -14640 77910
rect -14360 78090 -14140 78140
rect -14360 78020 -14350 78090
rect -14150 78020 -14140 78090
rect -14360 77980 -14140 78020
rect -14360 77910 -14350 77980
rect -14150 77910 -14140 77980
rect -14360 77860 -14140 77910
rect -13860 78090 -13640 78140
rect -13860 78020 -13850 78090
rect -13650 78020 -13640 78090
rect -13860 77980 -13640 78020
rect -13860 77910 -13850 77980
rect -13650 77910 -13640 77980
rect -13860 77860 -13640 77910
rect -13360 78090 -13140 78140
rect -13360 78020 -13350 78090
rect -13150 78020 -13140 78090
rect -13360 77980 -13140 78020
rect -13360 77910 -13350 77980
rect -13150 77910 -13140 77980
rect -13360 77860 -13140 77910
rect -12860 78090 -12640 78140
rect -12860 78020 -12850 78090
rect -12650 78020 -12640 78090
rect -12860 77980 -12640 78020
rect -12860 77910 -12850 77980
rect -12650 77910 -12640 77980
rect -12860 77860 -12640 77910
rect -12360 78090 -12140 78140
rect -12360 78020 -12350 78090
rect -12150 78020 -12140 78090
rect -12360 77980 -12140 78020
rect -12360 77910 -12350 77980
rect -12150 77910 -12140 77980
rect -12360 77860 -12140 77910
rect 96140 78090 96360 78140
rect 96140 78020 96150 78090
rect 96350 78020 96360 78090
rect 96140 77980 96360 78020
rect 96140 77910 96150 77980
rect 96350 77910 96360 77980
rect 96140 77860 96360 77910
rect 96640 78090 96860 78140
rect 96640 78020 96650 78090
rect 96850 78020 96860 78090
rect 96640 77980 96860 78020
rect 96640 77910 96650 77980
rect 96850 77910 96860 77980
rect 96640 77860 96860 77910
rect 97140 78090 97360 78140
rect 97140 78020 97150 78090
rect 97350 78020 97360 78090
rect 97140 77980 97360 78020
rect 97140 77910 97150 77980
rect 97350 77910 97360 77980
rect 97140 77860 97360 77910
rect 97640 78090 97860 78140
rect 97640 78020 97650 78090
rect 97850 78020 97860 78090
rect 97640 77980 97860 78020
rect 97640 77910 97650 77980
rect 97850 77910 97860 77980
rect 97640 77860 97860 77910
rect 98140 78090 98360 78140
rect 98140 78020 98150 78090
rect 98350 78020 98360 78090
rect 98140 77980 98360 78020
rect 98140 77910 98150 77980
rect 98350 77910 98360 77980
rect 98140 77860 98360 77910
rect 98640 78090 98860 78140
rect 98640 78020 98650 78090
rect 98850 78020 98860 78090
rect 98640 77980 98860 78020
rect 98640 77910 98650 77980
rect 98850 77910 98860 77980
rect 98640 77860 98860 77910
rect 99140 78090 99360 78140
rect 99140 78020 99150 78090
rect 99350 78020 99360 78090
rect 99140 77980 99360 78020
rect 99140 77910 99150 77980
rect 99350 77910 99360 77980
rect 99140 77860 99360 77910
rect 99640 78090 99860 78140
rect 99640 78020 99650 78090
rect 99850 78020 99860 78090
rect 99640 77980 99860 78020
rect 99640 77910 99650 77980
rect 99850 77910 99860 77980
rect 99640 77860 99860 77910
rect -16000 77850 -12000 77860
rect -16000 77650 -15980 77850
rect -15910 77650 -15590 77850
rect -15520 77650 -15480 77850
rect -15410 77650 -15090 77850
rect -15020 77650 -14980 77850
rect -14910 77650 -14590 77850
rect -14520 77650 -14480 77850
rect -14410 77650 -14090 77850
rect -14020 77650 -13980 77850
rect -13910 77650 -13590 77850
rect -13520 77650 -13480 77850
rect -13410 77650 -13090 77850
rect -13020 77650 -12980 77850
rect -12910 77650 -12590 77850
rect -12520 77650 -12480 77850
rect -12410 77650 -12090 77850
rect -12020 77650 -12000 77850
rect -16000 77640 -12000 77650
rect 96000 77850 100000 77860
rect 96000 77650 96020 77850
rect 96090 77650 96410 77850
rect 96480 77650 96520 77850
rect 96590 77650 96910 77850
rect 96980 77650 97020 77850
rect 97090 77650 97410 77850
rect 97480 77650 97520 77850
rect 97590 77650 97910 77850
rect 97980 77650 98020 77850
rect 98090 77650 98410 77850
rect 98480 77650 98520 77850
rect 98590 77650 98910 77850
rect 98980 77650 99020 77850
rect 99090 77650 99410 77850
rect 99480 77650 99520 77850
rect 99590 77650 99910 77850
rect 99980 77650 100000 77850
rect 96000 77640 100000 77650
rect -15860 77590 -15640 77640
rect -15860 77520 -15850 77590
rect -15650 77520 -15640 77590
rect -15860 77480 -15640 77520
rect -15860 77410 -15850 77480
rect -15650 77410 -15640 77480
rect -15860 77360 -15640 77410
rect -15360 77590 -15140 77640
rect -15360 77520 -15350 77590
rect -15150 77520 -15140 77590
rect -15360 77480 -15140 77520
rect -15360 77410 -15350 77480
rect -15150 77410 -15140 77480
rect -15360 77360 -15140 77410
rect -14860 77590 -14640 77640
rect -14860 77520 -14850 77590
rect -14650 77520 -14640 77590
rect -14860 77480 -14640 77520
rect -14860 77410 -14850 77480
rect -14650 77410 -14640 77480
rect -14860 77360 -14640 77410
rect -14360 77590 -14140 77640
rect -14360 77520 -14350 77590
rect -14150 77520 -14140 77590
rect -14360 77480 -14140 77520
rect -14360 77410 -14350 77480
rect -14150 77410 -14140 77480
rect -14360 77360 -14140 77410
rect -13860 77590 -13640 77640
rect -13860 77520 -13850 77590
rect -13650 77520 -13640 77590
rect -13860 77480 -13640 77520
rect -13860 77410 -13850 77480
rect -13650 77410 -13640 77480
rect -13860 77360 -13640 77410
rect -13360 77590 -13140 77640
rect -13360 77520 -13350 77590
rect -13150 77520 -13140 77590
rect -13360 77480 -13140 77520
rect -13360 77410 -13350 77480
rect -13150 77410 -13140 77480
rect -13360 77360 -13140 77410
rect -12860 77590 -12640 77640
rect -12860 77520 -12850 77590
rect -12650 77520 -12640 77590
rect -12860 77480 -12640 77520
rect -12860 77410 -12850 77480
rect -12650 77410 -12640 77480
rect -12860 77360 -12640 77410
rect -12360 77590 -12140 77640
rect -12360 77520 -12350 77590
rect -12150 77520 -12140 77590
rect -12360 77480 -12140 77520
rect -12360 77410 -12350 77480
rect -12150 77410 -12140 77480
rect -12360 77360 -12140 77410
rect 96140 77590 96360 77640
rect 96140 77520 96150 77590
rect 96350 77520 96360 77590
rect 96140 77480 96360 77520
rect 96140 77410 96150 77480
rect 96350 77410 96360 77480
rect 96140 77360 96360 77410
rect 96640 77590 96860 77640
rect 96640 77520 96650 77590
rect 96850 77520 96860 77590
rect 96640 77480 96860 77520
rect 96640 77410 96650 77480
rect 96850 77410 96860 77480
rect 96640 77360 96860 77410
rect 97140 77590 97360 77640
rect 97140 77520 97150 77590
rect 97350 77520 97360 77590
rect 97140 77480 97360 77520
rect 97140 77410 97150 77480
rect 97350 77410 97360 77480
rect 97140 77360 97360 77410
rect 97640 77590 97860 77640
rect 97640 77520 97650 77590
rect 97850 77520 97860 77590
rect 97640 77480 97860 77520
rect 97640 77410 97650 77480
rect 97850 77410 97860 77480
rect 97640 77360 97860 77410
rect 98140 77590 98360 77640
rect 98140 77520 98150 77590
rect 98350 77520 98360 77590
rect 98140 77480 98360 77520
rect 98140 77410 98150 77480
rect 98350 77410 98360 77480
rect 98140 77360 98360 77410
rect 98640 77590 98860 77640
rect 98640 77520 98650 77590
rect 98850 77520 98860 77590
rect 98640 77480 98860 77520
rect 98640 77410 98650 77480
rect 98850 77410 98860 77480
rect 98640 77360 98860 77410
rect 99140 77590 99360 77640
rect 99140 77520 99150 77590
rect 99350 77520 99360 77590
rect 99140 77480 99360 77520
rect 99140 77410 99150 77480
rect 99350 77410 99360 77480
rect 99140 77360 99360 77410
rect 99640 77590 99860 77640
rect 99640 77520 99650 77590
rect 99850 77520 99860 77590
rect 99640 77480 99860 77520
rect 99640 77410 99650 77480
rect 99850 77410 99860 77480
rect 99640 77360 99860 77410
rect -16000 77350 -12000 77360
rect -16000 77150 -15980 77350
rect -15910 77150 -15590 77350
rect -15520 77150 -15480 77350
rect -15410 77150 -15090 77350
rect -15020 77150 -14980 77350
rect -14910 77150 -14590 77350
rect -14520 77150 -14480 77350
rect -14410 77150 -14090 77350
rect -14020 77150 -13980 77350
rect -13910 77150 -13590 77350
rect -13520 77150 -13480 77350
rect -13410 77150 -13090 77350
rect -13020 77150 -12980 77350
rect -12910 77150 -12590 77350
rect -12520 77150 -12480 77350
rect -12410 77150 -12090 77350
rect -12020 77150 -12000 77350
rect -16000 77140 -12000 77150
rect 96000 77350 100000 77360
rect 96000 77150 96020 77350
rect 96090 77150 96410 77350
rect 96480 77150 96520 77350
rect 96590 77150 96910 77350
rect 96980 77150 97020 77350
rect 97090 77150 97410 77350
rect 97480 77150 97520 77350
rect 97590 77150 97910 77350
rect 97980 77150 98020 77350
rect 98090 77150 98410 77350
rect 98480 77150 98520 77350
rect 98590 77150 98910 77350
rect 98980 77150 99020 77350
rect 99090 77150 99410 77350
rect 99480 77150 99520 77350
rect 99590 77150 99910 77350
rect 99980 77150 100000 77350
rect 96000 77140 100000 77150
rect -15860 77090 -15640 77140
rect -15860 77020 -15850 77090
rect -15650 77020 -15640 77090
rect -15860 76980 -15640 77020
rect -15860 76910 -15850 76980
rect -15650 76910 -15640 76980
rect -15860 76860 -15640 76910
rect -15360 77090 -15140 77140
rect -15360 77020 -15350 77090
rect -15150 77020 -15140 77090
rect -15360 76980 -15140 77020
rect -15360 76910 -15350 76980
rect -15150 76910 -15140 76980
rect -15360 76860 -15140 76910
rect -14860 77090 -14640 77140
rect -14860 77020 -14850 77090
rect -14650 77020 -14640 77090
rect -14860 76980 -14640 77020
rect -14860 76910 -14850 76980
rect -14650 76910 -14640 76980
rect -14860 76860 -14640 76910
rect -14360 77090 -14140 77140
rect -14360 77020 -14350 77090
rect -14150 77020 -14140 77090
rect -14360 76980 -14140 77020
rect -14360 76910 -14350 76980
rect -14150 76910 -14140 76980
rect -14360 76860 -14140 76910
rect -13860 77090 -13640 77140
rect -13860 77020 -13850 77090
rect -13650 77020 -13640 77090
rect -13860 76980 -13640 77020
rect -13860 76910 -13850 76980
rect -13650 76910 -13640 76980
rect -13860 76860 -13640 76910
rect -13360 77090 -13140 77140
rect -13360 77020 -13350 77090
rect -13150 77020 -13140 77090
rect -13360 76980 -13140 77020
rect -13360 76910 -13350 76980
rect -13150 76910 -13140 76980
rect -13360 76860 -13140 76910
rect -12860 77090 -12640 77140
rect -12860 77020 -12850 77090
rect -12650 77020 -12640 77090
rect -12860 76980 -12640 77020
rect -12860 76910 -12850 76980
rect -12650 76910 -12640 76980
rect -12860 76860 -12640 76910
rect -12360 77090 -12140 77140
rect -12360 77020 -12350 77090
rect -12150 77020 -12140 77090
rect -12360 76980 -12140 77020
rect -12360 76910 -12350 76980
rect -12150 76910 -12140 76980
rect -12360 76860 -12140 76910
rect 96140 77090 96360 77140
rect 96140 77020 96150 77090
rect 96350 77020 96360 77090
rect 96140 76980 96360 77020
rect 96140 76910 96150 76980
rect 96350 76910 96360 76980
rect 96140 76860 96360 76910
rect 96640 77090 96860 77140
rect 96640 77020 96650 77090
rect 96850 77020 96860 77090
rect 96640 76980 96860 77020
rect 96640 76910 96650 76980
rect 96850 76910 96860 76980
rect 96640 76860 96860 76910
rect 97140 77090 97360 77140
rect 97140 77020 97150 77090
rect 97350 77020 97360 77090
rect 97140 76980 97360 77020
rect 97140 76910 97150 76980
rect 97350 76910 97360 76980
rect 97140 76860 97360 76910
rect 97640 77090 97860 77140
rect 97640 77020 97650 77090
rect 97850 77020 97860 77090
rect 97640 76980 97860 77020
rect 97640 76910 97650 76980
rect 97850 76910 97860 76980
rect 97640 76860 97860 76910
rect 98140 77090 98360 77140
rect 98140 77020 98150 77090
rect 98350 77020 98360 77090
rect 98140 76980 98360 77020
rect 98140 76910 98150 76980
rect 98350 76910 98360 76980
rect 98140 76860 98360 76910
rect 98640 77090 98860 77140
rect 98640 77020 98650 77090
rect 98850 77020 98860 77090
rect 98640 76980 98860 77020
rect 98640 76910 98650 76980
rect 98850 76910 98860 76980
rect 98640 76860 98860 76910
rect 99140 77090 99360 77140
rect 99140 77020 99150 77090
rect 99350 77020 99360 77090
rect 99140 76980 99360 77020
rect 99140 76910 99150 76980
rect 99350 76910 99360 76980
rect 99140 76860 99360 76910
rect 99640 77090 99860 77140
rect 99640 77020 99650 77090
rect 99850 77020 99860 77090
rect 99640 76980 99860 77020
rect 99640 76910 99650 76980
rect 99850 76910 99860 76980
rect 99640 76860 99860 76910
rect -16000 76850 -12000 76860
rect -16000 76650 -15980 76850
rect -15910 76650 -15590 76850
rect -15520 76650 -15480 76850
rect -15410 76650 -15090 76850
rect -15020 76650 -14980 76850
rect -14910 76650 -14590 76850
rect -14520 76650 -14480 76850
rect -14410 76650 -14090 76850
rect -14020 76650 -13980 76850
rect -13910 76650 -13590 76850
rect -13520 76650 -13480 76850
rect -13410 76650 -13090 76850
rect -13020 76650 -12980 76850
rect -12910 76650 -12590 76850
rect -12520 76650 -12480 76850
rect -12410 76650 -12090 76850
rect -12020 76650 -12000 76850
rect -16000 76640 -12000 76650
rect 96000 76850 100000 76860
rect 96000 76650 96020 76850
rect 96090 76650 96410 76850
rect 96480 76650 96520 76850
rect 96590 76650 96910 76850
rect 96980 76650 97020 76850
rect 97090 76650 97410 76850
rect 97480 76650 97520 76850
rect 97590 76650 97910 76850
rect 97980 76650 98020 76850
rect 98090 76650 98410 76850
rect 98480 76650 98520 76850
rect 98590 76650 98910 76850
rect 98980 76650 99020 76850
rect 99090 76650 99410 76850
rect 99480 76650 99520 76850
rect 99590 76650 99910 76850
rect 99980 76650 100000 76850
rect 96000 76640 100000 76650
rect -15860 76590 -15640 76640
rect -15860 76520 -15850 76590
rect -15650 76520 -15640 76590
rect -15860 76480 -15640 76520
rect -15860 76410 -15850 76480
rect -15650 76410 -15640 76480
rect -15860 76360 -15640 76410
rect -15360 76590 -15140 76640
rect -15360 76520 -15350 76590
rect -15150 76520 -15140 76590
rect -15360 76480 -15140 76520
rect -15360 76410 -15350 76480
rect -15150 76410 -15140 76480
rect -15360 76360 -15140 76410
rect -14860 76590 -14640 76640
rect -14860 76520 -14850 76590
rect -14650 76520 -14640 76590
rect -14860 76480 -14640 76520
rect -14860 76410 -14850 76480
rect -14650 76410 -14640 76480
rect -14860 76360 -14640 76410
rect -14360 76590 -14140 76640
rect -14360 76520 -14350 76590
rect -14150 76520 -14140 76590
rect -14360 76480 -14140 76520
rect -14360 76410 -14350 76480
rect -14150 76410 -14140 76480
rect -14360 76360 -14140 76410
rect -13860 76590 -13640 76640
rect -13860 76520 -13850 76590
rect -13650 76520 -13640 76590
rect -13860 76480 -13640 76520
rect -13860 76410 -13850 76480
rect -13650 76410 -13640 76480
rect -13860 76360 -13640 76410
rect -13360 76590 -13140 76640
rect -13360 76520 -13350 76590
rect -13150 76520 -13140 76590
rect -13360 76480 -13140 76520
rect -13360 76410 -13350 76480
rect -13150 76410 -13140 76480
rect -13360 76360 -13140 76410
rect -12860 76590 -12640 76640
rect -12860 76520 -12850 76590
rect -12650 76520 -12640 76590
rect -12860 76480 -12640 76520
rect -12860 76410 -12850 76480
rect -12650 76410 -12640 76480
rect -12860 76360 -12640 76410
rect -12360 76590 -12140 76640
rect -12360 76520 -12350 76590
rect -12150 76520 -12140 76590
rect -12360 76480 -12140 76520
rect -12360 76410 -12350 76480
rect -12150 76410 -12140 76480
rect -12360 76360 -12140 76410
rect 96140 76590 96360 76640
rect 96140 76520 96150 76590
rect 96350 76520 96360 76590
rect 96140 76480 96360 76520
rect 96140 76410 96150 76480
rect 96350 76410 96360 76480
rect 96140 76360 96360 76410
rect 96640 76590 96860 76640
rect 96640 76520 96650 76590
rect 96850 76520 96860 76590
rect 96640 76480 96860 76520
rect 96640 76410 96650 76480
rect 96850 76410 96860 76480
rect 96640 76360 96860 76410
rect 97140 76590 97360 76640
rect 97140 76520 97150 76590
rect 97350 76520 97360 76590
rect 97140 76480 97360 76520
rect 97140 76410 97150 76480
rect 97350 76410 97360 76480
rect 97140 76360 97360 76410
rect 97640 76590 97860 76640
rect 97640 76520 97650 76590
rect 97850 76520 97860 76590
rect 97640 76480 97860 76520
rect 97640 76410 97650 76480
rect 97850 76410 97860 76480
rect 97640 76360 97860 76410
rect 98140 76590 98360 76640
rect 98140 76520 98150 76590
rect 98350 76520 98360 76590
rect 98140 76480 98360 76520
rect 98140 76410 98150 76480
rect 98350 76410 98360 76480
rect 98140 76360 98360 76410
rect 98640 76590 98860 76640
rect 98640 76520 98650 76590
rect 98850 76520 98860 76590
rect 98640 76480 98860 76520
rect 98640 76410 98650 76480
rect 98850 76410 98860 76480
rect 98640 76360 98860 76410
rect 99140 76590 99360 76640
rect 99140 76520 99150 76590
rect 99350 76520 99360 76590
rect 99140 76480 99360 76520
rect 99140 76410 99150 76480
rect 99350 76410 99360 76480
rect 99140 76360 99360 76410
rect 99640 76590 99860 76640
rect 99640 76520 99650 76590
rect 99850 76520 99860 76590
rect 99640 76480 99860 76520
rect 99640 76410 99650 76480
rect 99850 76410 99860 76480
rect 99640 76360 99860 76410
rect -16000 76350 -12000 76360
rect -16000 76150 -15980 76350
rect -15910 76150 -15590 76350
rect -15520 76150 -15480 76350
rect -15410 76150 -15090 76350
rect -15020 76150 -14980 76350
rect -14910 76150 -14590 76350
rect -14520 76150 -14480 76350
rect -14410 76150 -14090 76350
rect -14020 76150 -13980 76350
rect -13910 76150 -13590 76350
rect -13520 76150 -13480 76350
rect -13410 76150 -13090 76350
rect -13020 76150 -12980 76350
rect -12910 76150 -12590 76350
rect -12520 76150 -12480 76350
rect -12410 76150 -12090 76350
rect -12020 76150 -12000 76350
rect -16000 76140 -12000 76150
rect 96000 76350 100000 76360
rect 96000 76150 96020 76350
rect 96090 76150 96410 76350
rect 96480 76150 96520 76350
rect 96590 76150 96910 76350
rect 96980 76150 97020 76350
rect 97090 76150 97410 76350
rect 97480 76150 97520 76350
rect 97590 76150 97910 76350
rect 97980 76150 98020 76350
rect 98090 76150 98410 76350
rect 98480 76150 98520 76350
rect 98590 76150 98910 76350
rect 98980 76150 99020 76350
rect 99090 76150 99410 76350
rect 99480 76150 99520 76350
rect 99590 76150 99910 76350
rect 99980 76150 100000 76350
rect 96000 76140 100000 76150
rect -15860 76090 -15640 76140
rect -15860 76020 -15850 76090
rect -15650 76020 -15640 76090
rect -15860 75980 -15640 76020
rect -15860 75910 -15850 75980
rect -15650 75910 -15640 75980
rect -15860 75860 -15640 75910
rect -15360 76090 -15140 76140
rect -15360 76020 -15350 76090
rect -15150 76020 -15140 76090
rect -15360 75980 -15140 76020
rect -15360 75910 -15350 75980
rect -15150 75910 -15140 75980
rect -15360 75860 -15140 75910
rect -14860 76090 -14640 76140
rect -14860 76020 -14850 76090
rect -14650 76020 -14640 76090
rect -14860 75980 -14640 76020
rect -14860 75910 -14850 75980
rect -14650 75910 -14640 75980
rect -14860 75860 -14640 75910
rect -14360 76090 -14140 76140
rect -14360 76020 -14350 76090
rect -14150 76020 -14140 76090
rect -14360 75980 -14140 76020
rect -14360 75910 -14350 75980
rect -14150 75910 -14140 75980
rect -14360 75860 -14140 75910
rect -13860 76090 -13640 76140
rect -13860 76020 -13850 76090
rect -13650 76020 -13640 76090
rect -13860 75980 -13640 76020
rect -13860 75910 -13850 75980
rect -13650 75910 -13640 75980
rect -13860 75860 -13640 75910
rect -13360 76090 -13140 76140
rect -13360 76020 -13350 76090
rect -13150 76020 -13140 76090
rect -13360 75980 -13140 76020
rect -13360 75910 -13350 75980
rect -13150 75910 -13140 75980
rect -13360 75860 -13140 75910
rect -12860 76090 -12640 76140
rect -12860 76020 -12850 76090
rect -12650 76020 -12640 76090
rect -12860 75980 -12640 76020
rect -12860 75910 -12850 75980
rect -12650 75910 -12640 75980
rect -12860 75860 -12640 75910
rect -12360 76090 -12140 76140
rect -12360 76020 -12350 76090
rect -12150 76020 -12140 76090
rect -12360 75980 -12140 76020
rect -12360 75910 -12350 75980
rect -12150 75910 -12140 75980
rect -12360 75860 -12140 75910
rect 96140 76090 96360 76140
rect 96140 76020 96150 76090
rect 96350 76020 96360 76090
rect 96140 75980 96360 76020
rect 96140 75910 96150 75980
rect 96350 75910 96360 75980
rect 96140 75860 96360 75910
rect 96640 76090 96860 76140
rect 96640 76020 96650 76090
rect 96850 76020 96860 76090
rect 96640 75980 96860 76020
rect 96640 75910 96650 75980
rect 96850 75910 96860 75980
rect 96640 75860 96860 75910
rect 97140 76090 97360 76140
rect 97140 76020 97150 76090
rect 97350 76020 97360 76090
rect 97140 75980 97360 76020
rect 97140 75910 97150 75980
rect 97350 75910 97360 75980
rect 97140 75860 97360 75910
rect 97640 76090 97860 76140
rect 97640 76020 97650 76090
rect 97850 76020 97860 76090
rect 97640 75980 97860 76020
rect 97640 75910 97650 75980
rect 97850 75910 97860 75980
rect 97640 75860 97860 75910
rect 98140 76090 98360 76140
rect 98140 76020 98150 76090
rect 98350 76020 98360 76090
rect 98140 75980 98360 76020
rect 98140 75910 98150 75980
rect 98350 75910 98360 75980
rect 98140 75860 98360 75910
rect 98640 76090 98860 76140
rect 98640 76020 98650 76090
rect 98850 76020 98860 76090
rect 98640 75980 98860 76020
rect 98640 75910 98650 75980
rect 98850 75910 98860 75980
rect 98640 75860 98860 75910
rect 99140 76090 99360 76140
rect 99140 76020 99150 76090
rect 99350 76020 99360 76090
rect 99140 75980 99360 76020
rect 99140 75910 99150 75980
rect 99350 75910 99360 75980
rect 99140 75860 99360 75910
rect 99640 76090 99860 76140
rect 99640 76020 99650 76090
rect 99850 76020 99860 76090
rect 99640 75980 99860 76020
rect 99640 75910 99650 75980
rect 99850 75910 99860 75980
rect 99640 75860 99860 75910
rect -16000 75850 -12000 75860
rect -16000 75650 -15980 75850
rect -15910 75650 -15590 75850
rect -15520 75650 -15480 75850
rect -15410 75650 -15090 75850
rect -15020 75650 -14980 75850
rect -14910 75650 -14590 75850
rect -14520 75650 -14480 75850
rect -14410 75650 -14090 75850
rect -14020 75650 -13980 75850
rect -13910 75650 -13590 75850
rect -13520 75650 -13480 75850
rect -13410 75650 -13090 75850
rect -13020 75650 -12980 75850
rect -12910 75650 -12590 75850
rect -12520 75650 -12480 75850
rect -12410 75650 -12090 75850
rect -12020 75650 -12000 75850
rect -16000 75640 -12000 75650
rect 96000 75850 100000 75860
rect 96000 75650 96020 75850
rect 96090 75650 96410 75850
rect 96480 75650 96520 75850
rect 96590 75650 96910 75850
rect 96980 75650 97020 75850
rect 97090 75650 97410 75850
rect 97480 75650 97520 75850
rect 97590 75650 97910 75850
rect 97980 75650 98020 75850
rect 98090 75650 98410 75850
rect 98480 75650 98520 75850
rect 98590 75650 98910 75850
rect 98980 75650 99020 75850
rect 99090 75650 99410 75850
rect 99480 75650 99520 75850
rect 99590 75650 99910 75850
rect 99980 75650 100000 75850
rect 96000 75640 100000 75650
rect -15860 75590 -15640 75640
rect -15860 75520 -15850 75590
rect -15650 75520 -15640 75590
rect -15860 75480 -15640 75520
rect -15860 75410 -15850 75480
rect -15650 75410 -15640 75480
rect -15860 75360 -15640 75410
rect -15360 75590 -15140 75640
rect -15360 75520 -15350 75590
rect -15150 75520 -15140 75590
rect -15360 75480 -15140 75520
rect -15360 75410 -15350 75480
rect -15150 75410 -15140 75480
rect -15360 75360 -15140 75410
rect -14860 75590 -14640 75640
rect -14860 75520 -14850 75590
rect -14650 75520 -14640 75590
rect -14860 75480 -14640 75520
rect -14860 75410 -14850 75480
rect -14650 75410 -14640 75480
rect -14860 75360 -14640 75410
rect -14360 75590 -14140 75640
rect -14360 75520 -14350 75590
rect -14150 75520 -14140 75590
rect -14360 75480 -14140 75520
rect -14360 75410 -14350 75480
rect -14150 75410 -14140 75480
rect -14360 75360 -14140 75410
rect -13860 75590 -13640 75640
rect -13860 75520 -13850 75590
rect -13650 75520 -13640 75590
rect -13860 75480 -13640 75520
rect -13860 75410 -13850 75480
rect -13650 75410 -13640 75480
rect -13860 75360 -13640 75410
rect -13360 75590 -13140 75640
rect -13360 75520 -13350 75590
rect -13150 75520 -13140 75590
rect -13360 75480 -13140 75520
rect -13360 75410 -13350 75480
rect -13150 75410 -13140 75480
rect -13360 75360 -13140 75410
rect -12860 75590 -12640 75640
rect -12860 75520 -12850 75590
rect -12650 75520 -12640 75590
rect -12860 75480 -12640 75520
rect -12860 75410 -12850 75480
rect -12650 75410 -12640 75480
rect -12860 75360 -12640 75410
rect -12360 75590 -12140 75640
rect -12360 75520 -12350 75590
rect -12150 75520 -12140 75590
rect -12360 75480 -12140 75520
rect -12360 75410 -12350 75480
rect -12150 75410 -12140 75480
rect -12360 75360 -12140 75410
rect 96140 75590 96360 75640
rect 96140 75520 96150 75590
rect 96350 75520 96360 75590
rect 96140 75480 96360 75520
rect 96140 75410 96150 75480
rect 96350 75410 96360 75480
rect 96140 75360 96360 75410
rect 96640 75590 96860 75640
rect 96640 75520 96650 75590
rect 96850 75520 96860 75590
rect 96640 75480 96860 75520
rect 96640 75410 96650 75480
rect 96850 75410 96860 75480
rect 96640 75360 96860 75410
rect 97140 75590 97360 75640
rect 97140 75520 97150 75590
rect 97350 75520 97360 75590
rect 97140 75480 97360 75520
rect 97140 75410 97150 75480
rect 97350 75410 97360 75480
rect 97140 75360 97360 75410
rect 97640 75590 97860 75640
rect 97640 75520 97650 75590
rect 97850 75520 97860 75590
rect 97640 75480 97860 75520
rect 97640 75410 97650 75480
rect 97850 75410 97860 75480
rect 97640 75360 97860 75410
rect 98140 75590 98360 75640
rect 98140 75520 98150 75590
rect 98350 75520 98360 75590
rect 98140 75480 98360 75520
rect 98140 75410 98150 75480
rect 98350 75410 98360 75480
rect 98140 75360 98360 75410
rect 98640 75590 98860 75640
rect 98640 75520 98650 75590
rect 98850 75520 98860 75590
rect 98640 75480 98860 75520
rect 98640 75410 98650 75480
rect 98850 75410 98860 75480
rect 98640 75360 98860 75410
rect 99140 75590 99360 75640
rect 99140 75520 99150 75590
rect 99350 75520 99360 75590
rect 99140 75480 99360 75520
rect 99140 75410 99150 75480
rect 99350 75410 99360 75480
rect 99140 75360 99360 75410
rect 99640 75590 99860 75640
rect 99640 75520 99650 75590
rect 99850 75520 99860 75590
rect 99640 75480 99860 75520
rect 99640 75410 99650 75480
rect 99850 75410 99860 75480
rect 99640 75360 99860 75410
rect -16000 75350 -12000 75360
rect -16000 75150 -15980 75350
rect -15910 75150 -15590 75350
rect -15520 75150 -15480 75350
rect -15410 75150 -15090 75350
rect -15020 75150 -14980 75350
rect -14910 75150 -14590 75350
rect -14520 75150 -14480 75350
rect -14410 75150 -14090 75350
rect -14020 75150 -13980 75350
rect -13910 75150 -13590 75350
rect -13520 75150 -13480 75350
rect -13410 75150 -13090 75350
rect -13020 75150 -12980 75350
rect -12910 75150 -12590 75350
rect -12520 75150 -12480 75350
rect -12410 75150 -12090 75350
rect -12020 75150 -12000 75350
rect -16000 75140 -12000 75150
rect 96000 75350 100000 75360
rect 96000 75150 96020 75350
rect 96090 75150 96410 75350
rect 96480 75150 96520 75350
rect 96590 75150 96910 75350
rect 96980 75150 97020 75350
rect 97090 75150 97410 75350
rect 97480 75150 97520 75350
rect 97590 75150 97910 75350
rect 97980 75150 98020 75350
rect 98090 75150 98410 75350
rect 98480 75150 98520 75350
rect 98590 75150 98910 75350
rect 98980 75150 99020 75350
rect 99090 75150 99410 75350
rect 99480 75150 99520 75350
rect 99590 75150 99910 75350
rect 99980 75150 100000 75350
rect 96000 75140 100000 75150
rect -15860 75090 -15640 75140
rect -15860 75020 -15850 75090
rect -15650 75020 -15640 75090
rect -15860 74980 -15640 75020
rect -15860 74910 -15850 74980
rect -15650 74910 -15640 74980
rect -15860 74860 -15640 74910
rect -15360 75090 -15140 75140
rect -15360 75020 -15350 75090
rect -15150 75020 -15140 75090
rect -15360 74980 -15140 75020
rect -15360 74910 -15350 74980
rect -15150 74910 -15140 74980
rect -15360 74860 -15140 74910
rect -14860 75090 -14640 75140
rect -14860 75020 -14850 75090
rect -14650 75020 -14640 75090
rect -14860 74980 -14640 75020
rect -14860 74910 -14850 74980
rect -14650 74910 -14640 74980
rect -14860 74860 -14640 74910
rect -14360 75090 -14140 75140
rect -14360 75020 -14350 75090
rect -14150 75020 -14140 75090
rect -14360 74980 -14140 75020
rect -14360 74910 -14350 74980
rect -14150 74910 -14140 74980
rect -14360 74860 -14140 74910
rect -13860 75090 -13640 75140
rect -13860 75020 -13850 75090
rect -13650 75020 -13640 75090
rect -13860 74980 -13640 75020
rect -13860 74910 -13850 74980
rect -13650 74910 -13640 74980
rect -13860 74860 -13640 74910
rect -13360 75090 -13140 75140
rect -13360 75020 -13350 75090
rect -13150 75020 -13140 75090
rect -13360 74980 -13140 75020
rect -13360 74910 -13350 74980
rect -13150 74910 -13140 74980
rect -13360 74860 -13140 74910
rect -12860 75090 -12640 75140
rect -12860 75020 -12850 75090
rect -12650 75020 -12640 75090
rect -12860 74980 -12640 75020
rect -12860 74910 -12850 74980
rect -12650 74910 -12640 74980
rect -12860 74860 -12640 74910
rect -12360 75090 -12140 75140
rect -12360 75020 -12350 75090
rect -12150 75020 -12140 75090
rect -12360 74980 -12140 75020
rect -12360 74910 -12350 74980
rect -12150 74910 -12140 74980
rect -12360 74860 -12140 74910
rect 96140 75090 96360 75140
rect 96140 75020 96150 75090
rect 96350 75020 96360 75090
rect 96140 74980 96360 75020
rect 96140 74910 96150 74980
rect 96350 74910 96360 74980
rect 96140 74860 96360 74910
rect 96640 75090 96860 75140
rect 96640 75020 96650 75090
rect 96850 75020 96860 75090
rect 96640 74980 96860 75020
rect 96640 74910 96650 74980
rect 96850 74910 96860 74980
rect 96640 74860 96860 74910
rect 97140 75090 97360 75140
rect 97140 75020 97150 75090
rect 97350 75020 97360 75090
rect 97140 74980 97360 75020
rect 97140 74910 97150 74980
rect 97350 74910 97360 74980
rect 97140 74860 97360 74910
rect 97640 75090 97860 75140
rect 97640 75020 97650 75090
rect 97850 75020 97860 75090
rect 97640 74980 97860 75020
rect 97640 74910 97650 74980
rect 97850 74910 97860 74980
rect 97640 74860 97860 74910
rect 98140 75090 98360 75140
rect 98140 75020 98150 75090
rect 98350 75020 98360 75090
rect 98140 74980 98360 75020
rect 98140 74910 98150 74980
rect 98350 74910 98360 74980
rect 98140 74860 98360 74910
rect 98640 75090 98860 75140
rect 98640 75020 98650 75090
rect 98850 75020 98860 75090
rect 98640 74980 98860 75020
rect 98640 74910 98650 74980
rect 98850 74910 98860 74980
rect 98640 74860 98860 74910
rect 99140 75090 99360 75140
rect 99140 75020 99150 75090
rect 99350 75020 99360 75090
rect 99140 74980 99360 75020
rect 99140 74910 99150 74980
rect 99350 74910 99360 74980
rect 99140 74860 99360 74910
rect 99640 75090 99860 75140
rect 99640 75020 99650 75090
rect 99850 75020 99860 75090
rect 99640 74980 99860 75020
rect 99640 74910 99650 74980
rect 99850 74910 99860 74980
rect 99640 74860 99860 74910
rect -16000 74850 -12000 74860
rect -16000 74650 -15980 74850
rect -15910 74650 -15590 74850
rect -15520 74650 -15480 74850
rect -15410 74650 -15090 74850
rect -15020 74650 -14980 74850
rect -14910 74650 -14590 74850
rect -14520 74650 -14480 74850
rect -14410 74650 -14090 74850
rect -14020 74650 -13980 74850
rect -13910 74650 -13590 74850
rect -13520 74650 -13480 74850
rect -13410 74650 -13090 74850
rect -13020 74650 -12980 74850
rect -12910 74650 -12590 74850
rect -12520 74650 -12480 74850
rect -12410 74650 -12090 74850
rect -12020 74650 -12000 74850
rect -16000 74640 -12000 74650
rect 96000 74850 100000 74860
rect 96000 74650 96020 74850
rect 96090 74650 96410 74850
rect 96480 74650 96520 74850
rect 96590 74650 96910 74850
rect 96980 74650 97020 74850
rect 97090 74650 97410 74850
rect 97480 74650 97520 74850
rect 97590 74650 97910 74850
rect 97980 74650 98020 74850
rect 98090 74650 98410 74850
rect 98480 74650 98520 74850
rect 98590 74650 98910 74850
rect 98980 74650 99020 74850
rect 99090 74650 99410 74850
rect 99480 74650 99520 74850
rect 99590 74650 99910 74850
rect 99980 74650 100000 74850
rect 96000 74640 100000 74650
rect -15860 74590 -15640 74640
rect -15860 74520 -15850 74590
rect -15650 74520 -15640 74590
rect -15860 74480 -15640 74520
rect -15860 74410 -15850 74480
rect -15650 74410 -15640 74480
rect -15860 74360 -15640 74410
rect -15360 74590 -15140 74640
rect -15360 74520 -15350 74590
rect -15150 74520 -15140 74590
rect -15360 74480 -15140 74520
rect -15360 74410 -15350 74480
rect -15150 74410 -15140 74480
rect -15360 74360 -15140 74410
rect -14860 74590 -14640 74640
rect -14860 74520 -14850 74590
rect -14650 74520 -14640 74590
rect -14860 74480 -14640 74520
rect -14860 74410 -14850 74480
rect -14650 74410 -14640 74480
rect -14860 74360 -14640 74410
rect -14360 74590 -14140 74640
rect -14360 74520 -14350 74590
rect -14150 74520 -14140 74590
rect -14360 74480 -14140 74520
rect -14360 74410 -14350 74480
rect -14150 74410 -14140 74480
rect -14360 74360 -14140 74410
rect -13860 74590 -13640 74640
rect -13860 74520 -13850 74590
rect -13650 74520 -13640 74590
rect -13860 74480 -13640 74520
rect -13860 74410 -13850 74480
rect -13650 74410 -13640 74480
rect -13860 74360 -13640 74410
rect -13360 74590 -13140 74640
rect -13360 74520 -13350 74590
rect -13150 74520 -13140 74590
rect -13360 74480 -13140 74520
rect -13360 74410 -13350 74480
rect -13150 74410 -13140 74480
rect -13360 74360 -13140 74410
rect -12860 74590 -12640 74640
rect -12860 74520 -12850 74590
rect -12650 74520 -12640 74590
rect -12860 74480 -12640 74520
rect -12860 74410 -12850 74480
rect -12650 74410 -12640 74480
rect -12860 74360 -12640 74410
rect -12360 74590 -12140 74640
rect -12360 74520 -12350 74590
rect -12150 74520 -12140 74590
rect -12360 74480 -12140 74520
rect -12360 74410 -12350 74480
rect -12150 74410 -12140 74480
rect -12360 74360 -12140 74410
rect 96140 74590 96360 74640
rect 96140 74520 96150 74590
rect 96350 74520 96360 74590
rect 96140 74480 96360 74520
rect 96140 74410 96150 74480
rect 96350 74410 96360 74480
rect 96140 74360 96360 74410
rect 96640 74590 96860 74640
rect 96640 74520 96650 74590
rect 96850 74520 96860 74590
rect 96640 74480 96860 74520
rect 96640 74410 96650 74480
rect 96850 74410 96860 74480
rect 96640 74360 96860 74410
rect 97140 74590 97360 74640
rect 97140 74520 97150 74590
rect 97350 74520 97360 74590
rect 97140 74480 97360 74520
rect 97140 74410 97150 74480
rect 97350 74410 97360 74480
rect 97140 74360 97360 74410
rect 97640 74590 97860 74640
rect 97640 74520 97650 74590
rect 97850 74520 97860 74590
rect 97640 74480 97860 74520
rect 97640 74410 97650 74480
rect 97850 74410 97860 74480
rect 97640 74360 97860 74410
rect 98140 74590 98360 74640
rect 98140 74520 98150 74590
rect 98350 74520 98360 74590
rect 98140 74480 98360 74520
rect 98140 74410 98150 74480
rect 98350 74410 98360 74480
rect 98140 74360 98360 74410
rect 98640 74590 98860 74640
rect 98640 74520 98650 74590
rect 98850 74520 98860 74590
rect 98640 74480 98860 74520
rect 98640 74410 98650 74480
rect 98850 74410 98860 74480
rect 98640 74360 98860 74410
rect 99140 74590 99360 74640
rect 99140 74520 99150 74590
rect 99350 74520 99360 74590
rect 99140 74480 99360 74520
rect 99140 74410 99150 74480
rect 99350 74410 99360 74480
rect 99140 74360 99360 74410
rect 99640 74590 99860 74640
rect 99640 74520 99650 74590
rect 99850 74520 99860 74590
rect 99640 74480 99860 74520
rect 99640 74410 99650 74480
rect 99850 74410 99860 74480
rect 99640 74360 99860 74410
rect -16000 74350 -12000 74360
rect -16000 74150 -15980 74350
rect -15910 74150 -15590 74350
rect -15520 74150 -15480 74350
rect -15410 74150 -15090 74350
rect -15020 74150 -14980 74350
rect -14910 74150 -14590 74350
rect -14520 74150 -14480 74350
rect -14410 74150 -14090 74350
rect -14020 74150 -13980 74350
rect -13910 74150 -13590 74350
rect -13520 74150 -13480 74350
rect -13410 74150 -13090 74350
rect -13020 74150 -12980 74350
rect -12910 74150 -12590 74350
rect -12520 74150 -12480 74350
rect -12410 74150 -12090 74350
rect -12020 74150 -12000 74350
rect -16000 74140 -12000 74150
rect 96000 74350 100000 74360
rect 96000 74150 96020 74350
rect 96090 74150 96410 74350
rect 96480 74150 96520 74350
rect 96590 74150 96910 74350
rect 96980 74150 97020 74350
rect 97090 74150 97410 74350
rect 97480 74150 97520 74350
rect 97590 74150 97910 74350
rect 97980 74150 98020 74350
rect 98090 74150 98410 74350
rect 98480 74150 98520 74350
rect 98590 74150 98910 74350
rect 98980 74150 99020 74350
rect 99090 74150 99410 74350
rect 99480 74150 99520 74350
rect 99590 74150 99910 74350
rect 99980 74150 100000 74350
rect 96000 74140 100000 74150
rect -15860 74090 -15640 74140
rect -15860 74020 -15850 74090
rect -15650 74020 -15640 74090
rect -15860 73980 -15640 74020
rect -15860 73910 -15850 73980
rect -15650 73910 -15640 73980
rect -15860 73860 -15640 73910
rect -15360 74090 -15140 74140
rect -15360 74020 -15350 74090
rect -15150 74020 -15140 74090
rect -15360 73980 -15140 74020
rect -15360 73910 -15350 73980
rect -15150 73910 -15140 73980
rect -15360 73860 -15140 73910
rect -14860 74090 -14640 74140
rect -14860 74020 -14850 74090
rect -14650 74020 -14640 74090
rect -14860 73980 -14640 74020
rect -14860 73910 -14850 73980
rect -14650 73910 -14640 73980
rect -14860 73860 -14640 73910
rect -14360 74090 -14140 74140
rect -14360 74020 -14350 74090
rect -14150 74020 -14140 74090
rect -14360 73980 -14140 74020
rect -14360 73910 -14350 73980
rect -14150 73910 -14140 73980
rect -14360 73860 -14140 73910
rect -13860 74090 -13640 74140
rect -13860 74020 -13850 74090
rect -13650 74020 -13640 74090
rect -13860 73980 -13640 74020
rect -13860 73910 -13850 73980
rect -13650 73910 -13640 73980
rect -13860 73860 -13640 73910
rect -13360 74090 -13140 74140
rect -13360 74020 -13350 74090
rect -13150 74020 -13140 74090
rect -13360 73980 -13140 74020
rect -13360 73910 -13350 73980
rect -13150 73910 -13140 73980
rect -13360 73860 -13140 73910
rect -12860 74090 -12640 74140
rect -12860 74020 -12850 74090
rect -12650 74020 -12640 74090
rect -12860 73980 -12640 74020
rect -12860 73910 -12850 73980
rect -12650 73910 -12640 73980
rect -12860 73860 -12640 73910
rect -12360 74090 -12140 74140
rect -12360 74020 -12350 74090
rect -12150 74020 -12140 74090
rect -12360 73980 -12140 74020
rect -12360 73910 -12350 73980
rect -12150 73910 -12140 73980
rect -12360 73860 -12140 73910
rect 96140 74090 96360 74140
rect 96140 74020 96150 74090
rect 96350 74020 96360 74090
rect 96140 73980 96360 74020
rect 96140 73910 96150 73980
rect 96350 73910 96360 73980
rect 96140 73860 96360 73910
rect 96640 74090 96860 74140
rect 96640 74020 96650 74090
rect 96850 74020 96860 74090
rect 96640 73980 96860 74020
rect 96640 73910 96650 73980
rect 96850 73910 96860 73980
rect 96640 73860 96860 73910
rect 97140 74090 97360 74140
rect 97140 74020 97150 74090
rect 97350 74020 97360 74090
rect 97140 73980 97360 74020
rect 97140 73910 97150 73980
rect 97350 73910 97360 73980
rect 97140 73860 97360 73910
rect 97640 74090 97860 74140
rect 97640 74020 97650 74090
rect 97850 74020 97860 74090
rect 97640 73980 97860 74020
rect 97640 73910 97650 73980
rect 97850 73910 97860 73980
rect 97640 73860 97860 73910
rect 98140 74090 98360 74140
rect 98140 74020 98150 74090
rect 98350 74020 98360 74090
rect 98140 73980 98360 74020
rect 98140 73910 98150 73980
rect 98350 73910 98360 73980
rect 98140 73860 98360 73910
rect 98640 74090 98860 74140
rect 98640 74020 98650 74090
rect 98850 74020 98860 74090
rect 98640 73980 98860 74020
rect 98640 73910 98650 73980
rect 98850 73910 98860 73980
rect 98640 73860 98860 73910
rect 99140 74090 99360 74140
rect 99140 74020 99150 74090
rect 99350 74020 99360 74090
rect 99140 73980 99360 74020
rect 99140 73910 99150 73980
rect 99350 73910 99360 73980
rect 99140 73860 99360 73910
rect 99640 74090 99860 74140
rect 99640 74020 99650 74090
rect 99850 74020 99860 74090
rect 99640 73980 99860 74020
rect 99640 73910 99650 73980
rect 99850 73910 99860 73980
rect 99640 73860 99860 73910
rect -16000 73850 -12000 73860
rect -16000 73650 -15980 73850
rect -15910 73650 -15590 73850
rect -15520 73650 -15480 73850
rect -15410 73650 -15090 73850
rect -15020 73650 -14980 73850
rect -14910 73650 -14590 73850
rect -14520 73650 -14480 73850
rect -14410 73650 -14090 73850
rect -14020 73650 -13980 73850
rect -13910 73650 -13590 73850
rect -13520 73650 -13480 73850
rect -13410 73650 -13090 73850
rect -13020 73650 -12980 73850
rect -12910 73650 -12590 73850
rect -12520 73650 -12480 73850
rect -12410 73650 -12090 73850
rect -12020 73650 -12000 73850
rect -16000 73640 -12000 73650
rect 96000 73850 100000 73860
rect 96000 73650 96020 73850
rect 96090 73650 96410 73850
rect 96480 73650 96520 73850
rect 96590 73650 96910 73850
rect 96980 73650 97020 73850
rect 97090 73650 97410 73850
rect 97480 73650 97520 73850
rect 97590 73650 97910 73850
rect 97980 73650 98020 73850
rect 98090 73650 98410 73850
rect 98480 73650 98520 73850
rect 98590 73650 98910 73850
rect 98980 73650 99020 73850
rect 99090 73650 99410 73850
rect 99480 73650 99520 73850
rect 99590 73650 99910 73850
rect 99980 73650 100000 73850
rect 96000 73640 100000 73650
rect -15860 73590 -15640 73640
rect -15860 73520 -15850 73590
rect -15650 73520 -15640 73590
rect -15860 73480 -15640 73520
rect -15860 73410 -15850 73480
rect -15650 73410 -15640 73480
rect -15860 73360 -15640 73410
rect -15360 73590 -15140 73640
rect -15360 73520 -15350 73590
rect -15150 73520 -15140 73590
rect -15360 73480 -15140 73520
rect -15360 73410 -15350 73480
rect -15150 73410 -15140 73480
rect -15360 73360 -15140 73410
rect -14860 73590 -14640 73640
rect -14860 73520 -14850 73590
rect -14650 73520 -14640 73590
rect -14860 73480 -14640 73520
rect -14860 73410 -14850 73480
rect -14650 73410 -14640 73480
rect -14860 73360 -14640 73410
rect -14360 73590 -14140 73640
rect -14360 73520 -14350 73590
rect -14150 73520 -14140 73590
rect -14360 73480 -14140 73520
rect -14360 73410 -14350 73480
rect -14150 73410 -14140 73480
rect -14360 73360 -14140 73410
rect -13860 73590 -13640 73640
rect -13860 73520 -13850 73590
rect -13650 73520 -13640 73590
rect -13860 73480 -13640 73520
rect -13860 73410 -13850 73480
rect -13650 73410 -13640 73480
rect -13860 73360 -13640 73410
rect -13360 73590 -13140 73640
rect -13360 73520 -13350 73590
rect -13150 73520 -13140 73590
rect -13360 73480 -13140 73520
rect -13360 73410 -13350 73480
rect -13150 73410 -13140 73480
rect -13360 73360 -13140 73410
rect -12860 73590 -12640 73640
rect -12860 73520 -12850 73590
rect -12650 73520 -12640 73590
rect -12860 73480 -12640 73520
rect -12860 73410 -12850 73480
rect -12650 73410 -12640 73480
rect -12860 73360 -12640 73410
rect -12360 73590 -12140 73640
rect -12360 73520 -12350 73590
rect -12150 73520 -12140 73590
rect -12360 73480 -12140 73520
rect -12360 73410 -12350 73480
rect -12150 73410 -12140 73480
rect -12360 73360 -12140 73410
rect 96140 73590 96360 73640
rect 96140 73520 96150 73590
rect 96350 73520 96360 73590
rect 96140 73480 96360 73520
rect 96140 73410 96150 73480
rect 96350 73410 96360 73480
rect 96140 73360 96360 73410
rect 96640 73590 96860 73640
rect 96640 73520 96650 73590
rect 96850 73520 96860 73590
rect 96640 73480 96860 73520
rect 96640 73410 96650 73480
rect 96850 73410 96860 73480
rect 96640 73360 96860 73410
rect 97140 73590 97360 73640
rect 97140 73520 97150 73590
rect 97350 73520 97360 73590
rect 97140 73480 97360 73520
rect 97140 73410 97150 73480
rect 97350 73410 97360 73480
rect 97140 73360 97360 73410
rect 97640 73590 97860 73640
rect 97640 73520 97650 73590
rect 97850 73520 97860 73590
rect 97640 73480 97860 73520
rect 97640 73410 97650 73480
rect 97850 73410 97860 73480
rect 97640 73360 97860 73410
rect 98140 73590 98360 73640
rect 98140 73520 98150 73590
rect 98350 73520 98360 73590
rect 98140 73480 98360 73520
rect 98140 73410 98150 73480
rect 98350 73410 98360 73480
rect 98140 73360 98360 73410
rect 98640 73590 98860 73640
rect 98640 73520 98650 73590
rect 98850 73520 98860 73590
rect 98640 73480 98860 73520
rect 98640 73410 98650 73480
rect 98850 73410 98860 73480
rect 98640 73360 98860 73410
rect 99140 73590 99360 73640
rect 99140 73520 99150 73590
rect 99350 73520 99360 73590
rect 99140 73480 99360 73520
rect 99140 73410 99150 73480
rect 99350 73410 99360 73480
rect 99140 73360 99360 73410
rect 99640 73590 99860 73640
rect 99640 73520 99650 73590
rect 99850 73520 99860 73590
rect 99640 73480 99860 73520
rect 99640 73410 99650 73480
rect 99850 73410 99860 73480
rect 99640 73360 99860 73410
rect -16000 73350 -12000 73360
rect -16000 73150 -15980 73350
rect -15910 73150 -15590 73350
rect -15520 73150 -15480 73350
rect -15410 73150 -15090 73350
rect -15020 73150 -14980 73350
rect -14910 73150 -14590 73350
rect -14520 73150 -14480 73350
rect -14410 73150 -14090 73350
rect -14020 73150 -13980 73350
rect -13910 73150 -13590 73350
rect -13520 73150 -13480 73350
rect -13410 73150 -13090 73350
rect -13020 73150 -12980 73350
rect -12910 73150 -12590 73350
rect -12520 73150 -12480 73350
rect -12410 73150 -12090 73350
rect -12020 73150 -12000 73350
rect -16000 73140 -12000 73150
rect 96000 73350 100000 73360
rect 96000 73150 96020 73350
rect 96090 73150 96410 73350
rect 96480 73150 96520 73350
rect 96590 73150 96910 73350
rect 96980 73150 97020 73350
rect 97090 73150 97410 73350
rect 97480 73150 97520 73350
rect 97590 73150 97910 73350
rect 97980 73150 98020 73350
rect 98090 73150 98410 73350
rect 98480 73150 98520 73350
rect 98590 73150 98910 73350
rect 98980 73150 99020 73350
rect 99090 73150 99410 73350
rect 99480 73150 99520 73350
rect 99590 73150 99910 73350
rect 99980 73150 100000 73350
rect 96000 73140 100000 73150
rect -15860 73090 -15640 73140
rect -15860 73020 -15850 73090
rect -15650 73020 -15640 73090
rect -15860 72980 -15640 73020
rect -15860 72910 -15850 72980
rect -15650 72910 -15640 72980
rect -15860 72860 -15640 72910
rect -15360 73090 -15140 73140
rect -15360 73020 -15350 73090
rect -15150 73020 -15140 73090
rect -15360 72980 -15140 73020
rect -15360 72910 -15350 72980
rect -15150 72910 -15140 72980
rect -15360 72860 -15140 72910
rect -14860 73090 -14640 73140
rect -14860 73020 -14850 73090
rect -14650 73020 -14640 73090
rect -14860 72980 -14640 73020
rect -14860 72910 -14850 72980
rect -14650 72910 -14640 72980
rect -14860 72860 -14640 72910
rect -14360 73090 -14140 73140
rect -14360 73020 -14350 73090
rect -14150 73020 -14140 73090
rect -14360 72980 -14140 73020
rect -14360 72910 -14350 72980
rect -14150 72910 -14140 72980
rect -14360 72860 -14140 72910
rect -13860 73090 -13640 73140
rect -13860 73020 -13850 73090
rect -13650 73020 -13640 73090
rect -13860 72980 -13640 73020
rect -13860 72910 -13850 72980
rect -13650 72910 -13640 72980
rect -13860 72860 -13640 72910
rect -13360 73090 -13140 73140
rect -13360 73020 -13350 73090
rect -13150 73020 -13140 73090
rect -13360 72980 -13140 73020
rect -13360 72910 -13350 72980
rect -13150 72910 -13140 72980
rect -13360 72860 -13140 72910
rect -12860 73090 -12640 73140
rect -12860 73020 -12850 73090
rect -12650 73020 -12640 73090
rect -12860 72980 -12640 73020
rect -12860 72910 -12850 72980
rect -12650 72910 -12640 72980
rect -12860 72860 -12640 72910
rect -12360 73090 -12140 73140
rect -12360 73020 -12350 73090
rect -12150 73020 -12140 73090
rect -12360 72980 -12140 73020
rect -12360 72910 -12350 72980
rect -12150 72910 -12140 72980
rect -12360 72860 -12140 72910
rect 96140 73090 96360 73140
rect 96140 73020 96150 73090
rect 96350 73020 96360 73090
rect 96140 72980 96360 73020
rect 96140 72910 96150 72980
rect 96350 72910 96360 72980
rect 96140 72860 96360 72910
rect 96640 73090 96860 73140
rect 96640 73020 96650 73090
rect 96850 73020 96860 73090
rect 96640 72980 96860 73020
rect 96640 72910 96650 72980
rect 96850 72910 96860 72980
rect 96640 72860 96860 72910
rect 97140 73090 97360 73140
rect 97140 73020 97150 73090
rect 97350 73020 97360 73090
rect 97140 72980 97360 73020
rect 97140 72910 97150 72980
rect 97350 72910 97360 72980
rect 97140 72860 97360 72910
rect 97640 73090 97860 73140
rect 97640 73020 97650 73090
rect 97850 73020 97860 73090
rect 97640 72980 97860 73020
rect 97640 72910 97650 72980
rect 97850 72910 97860 72980
rect 97640 72860 97860 72910
rect 98140 73090 98360 73140
rect 98140 73020 98150 73090
rect 98350 73020 98360 73090
rect 98140 72980 98360 73020
rect 98140 72910 98150 72980
rect 98350 72910 98360 72980
rect 98140 72860 98360 72910
rect 98640 73090 98860 73140
rect 98640 73020 98650 73090
rect 98850 73020 98860 73090
rect 98640 72980 98860 73020
rect 98640 72910 98650 72980
rect 98850 72910 98860 72980
rect 98640 72860 98860 72910
rect 99140 73090 99360 73140
rect 99140 73020 99150 73090
rect 99350 73020 99360 73090
rect 99140 72980 99360 73020
rect 99140 72910 99150 72980
rect 99350 72910 99360 72980
rect 99140 72860 99360 72910
rect 99640 73090 99860 73140
rect 99640 73020 99650 73090
rect 99850 73020 99860 73090
rect 99640 72980 99860 73020
rect 99640 72910 99650 72980
rect 99850 72910 99860 72980
rect 99640 72860 99860 72910
rect -16000 72850 -12000 72860
rect -16000 72650 -15980 72850
rect -15910 72650 -15590 72850
rect -15520 72650 -15480 72850
rect -15410 72650 -15090 72850
rect -15020 72650 -14980 72850
rect -14910 72650 -14590 72850
rect -14520 72650 -14480 72850
rect -14410 72650 -14090 72850
rect -14020 72650 -13980 72850
rect -13910 72650 -13590 72850
rect -13520 72650 -13480 72850
rect -13410 72650 -13090 72850
rect -13020 72650 -12980 72850
rect -12910 72650 -12590 72850
rect -12520 72650 -12480 72850
rect -12410 72650 -12090 72850
rect -12020 72650 -12000 72850
rect -16000 72640 -12000 72650
rect 96000 72850 100000 72860
rect 96000 72650 96020 72850
rect 96090 72650 96410 72850
rect 96480 72650 96520 72850
rect 96590 72650 96910 72850
rect 96980 72650 97020 72850
rect 97090 72650 97410 72850
rect 97480 72650 97520 72850
rect 97590 72650 97910 72850
rect 97980 72650 98020 72850
rect 98090 72650 98410 72850
rect 98480 72650 98520 72850
rect 98590 72650 98910 72850
rect 98980 72650 99020 72850
rect 99090 72650 99410 72850
rect 99480 72650 99520 72850
rect 99590 72650 99910 72850
rect 99980 72650 100000 72850
rect 96000 72640 100000 72650
rect -15860 72590 -15640 72640
rect -15860 72520 -15850 72590
rect -15650 72520 -15640 72590
rect -15860 72480 -15640 72520
rect -15860 72410 -15850 72480
rect -15650 72410 -15640 72480
rect -15860 72360 -15640 72410
rect -15360 72590 -15140 72640
rect -15360 72520 -15350 72590
rect -15150 72520 -15140 72590
rect -15360 72480 -15140 72520
rect -15360 72410 -15350 72480
rect -15150 72410 -15140 72480
rect -15360 72360 -15140 72410
rect -14860 72590 -14640 72640
rect -14860 72520 -14850 72590
rect -14650 72520 -14640 72590
rect -14860 72480 -14640 72520
rect -14860 72410 -14850 72480
rect -14650 72410 -14640 72480
rect -14860 72360 -14640 72410
rect -14360 72590 -14140 72640
rect -14360 72520 -14350 72590
rect -14150 72520 -14140 72590
rect -14360 72480 -14140 72520
rect -14360 72410 -14350 72480
rect -14150 72410 -14140 72480
rect -14360 72360 -14140 72410
rect -13860 72590 -13640 72640
rect -13860 72520 -13850 72590
rect -13650 72520 -13640 72590
rect -13860 72480 -13640 72520
rect -13860 72410 -13850 72480
rect -13650 72410 -13640 72480
rect -13860 72360 -13640 72410
rect -13360 72590 -13140 72640
rect -13360 72520 -13350 72590
rect -13150 72520 -13140 72590
rect -13360 72480 -13140 72520
rect -13360 72410 -13350 72480
rect -13150 72410 -13140 72480
rect -13360 72360 -13140 72410
rect -12860 72590 -12640 72640
rect -12860 72520 -12850 72590
rect -12650 72520 -12640 72590
rect -12860 72480 -12640 72520
rect -12860 72410 -12850 72480
rect -12650 72410 -12640 72480
rect -12860 72360 -12640 72410
rect -12360 72590 -12140 72640
rect -12360 72520 -12350 72590
rect -12150 72520 -12140 72590
rect -12360 72480 -12140 72520
rect -12360 72410 -12350 72480
rect -12150 72410 -12140 72480
rect -12360 72360 -12140 72410
rect 96140 72590 96360 72640
rect 96140 72520 96150 72590
rect 96350 72520 96360 72590
rect 96140 72480 96360 72520
rect 96140 72410 96150 72480
rect 96350 72410 96360 72480
rect 96140 72360 96360 72410
rect 96640 72590 96860 72640
rect 96640 72520 96650 72590
rect 96850 72520 96860 72590
rect 96640 72480 96860 72520
rect 96640 72410 96650 72480
rect 96850 72410 96860 72480
rect 96640 72360 96860 72410
rect 97140 72590 97360 72640
rect 97140 72520 97150 72590
rect 97350 72520 97360 72590
rect 97140 72480 97360 72520
rect 97140 72410 97150 72480
rect 97350 72410 97360 72480
rect 97140 72360 97360 72410
rect 97640 72590 97860 72640
rect 97640 72520 97650 72590
rect 97850 72520 97860 72590
rect 97640 72480 97860 72520
rect 97640 72410 97650 72480
rect 97850 72410 97860 72480
rect 97640 72360 97860 72410
rect 98140 72590 98360 72640
rect 98140 72520 98150 72590
rect 98350 72520 98360 72590
rect 98140 72480 98360 72520
rect 98140 72410 98150 72480
rect 98350 72410 98360 72480
rect 98140 72360 98360 72410
rect 98640 72590 98860 72640
rect 98640 72520 98650 72590
rect 98850 72520 98860 72590
rect 98640 72480 98860 72520
rect 98640 72410 98650 72480
rect 98850 72410 98860 72480
rect 98640 72360 98860 72410
rect 99140 72590 99360 72640
rect 99140 72520 99150 72590
rect 99350 72520 99360 72590
rect 99140 72480 99360 72520
rect 99140 72410 99150 72480
rect 99350 72410 99360 72480
rect 99140 72360 99360 72410
rect 99640 72590 99860 72640
rect 99640 72520 99650 72590
rect 99850 72520 99860 72590
rect 99640 72480 99860 72520
rect 99640 72410 99650 72480
rect 99850 72410 99860 72480
rect 99640 72360 99860 72410
rect -16000 72350 -12000 72360
rect -16000 72150 -15980 72350
rect -15910 72150 -15590 72350
rect -15520 72150 -15480 72350
rect -15410 72150 -15090 72350
rect -15020 72150 -14980 72350
rect -14910 72150 -14590 72350
rect -14520 72150 -14480 72350
rect -14410 72150 -14090 72350
rect -14020 72150 -13980 72350
rect -13910 72150 -13590 72350
rect -13520 72150 -13480 72350
rect -13410 72150 -13090 72350
rect -13020 72150 -12980 72350
rect -12910 72150 -12590 72350
rect -12520 72150 -12480 72350
rect -12410 72150 -12090 72350
rect -12020 72150 -12000 72350
rect -16000 72140 -12000 72150
rect 96000 72350 100000 72360
rect 96000 72150 96020 72350
rect 96090 72150 96410 72350
rect 96480 72150 96520 72350
rect 96590 72150 96910 72350
rect 96980 72150 97020 72350
rect 97090 72150 97410 72350
rect 97480 72150 97520 72350
rect 97590 72150 97910 72350
rect 97980 72150 98020 72350
rect 98090 72150 98410 72350
rect 98480 72150 98520 72350
rect 98590 72150 98910 72350
rect 98980 72150 99020 72350
rect 99090 72150 99410 72350
rect 99480 72150 99520 72350
rect 99590 72150 99910 72350
rect 99980 72150 100000 72350
rect 96000 72140 100000 72150
rect -15860 72090 -15640 72140
rect -15860 72020 -15850 72090
rect -15650 72020 -15640 72090
rect -15860 71980 -15640 72020
rect -15860 71910 -15850 71980
rect -15650 71910 -15640 71980
rect -15860 71860 -15640 71910
rect -15360 72090 -15140 72140
rect -15360 72020 -15350 72090
rect -15150 72020 -15140 72090
rect -15360 71980 -15140 72020
rect -15360 71910 -15350 71980
rect -15150 71910 -15140 71980
rect -15360 71860 -15140 71910
rect -14860 72090 -14640 72140
rect -14860 72020 -14850 72090
rect -14650 72020 -14640 72090
rect -14860 71980 -14640 72020
rect -14860 71910 -14850 71980
rect -14650 71910 -14640 71980
rect -14860 71860 -14640 71910
rect -14360 72090 -14140 72140
rect -14360 72020 -14350 72090
rect -14150 72020 -14140 72090
rect -14360 71980 -14140 72020
rect -14360 71910 -14350 71980
rect -14150 71910 -14140 71980
rect -14360 71860 -14140 71910
rect -13860 72090 -13640 72140
rect -13860 72020 -13850 72090
rect -13650 72020 -13640 72090
rect -13860 71980 -13640 72020
rect -13860 71910 -13850 71980
rect -13650 71910 -13640 71980
rect -13860 71860 -13640 71910
rect -13360 72090 -13140 72140
rect -13360 72020 -13350 72090
rect -13150 72020 -13140 72090
rect -13360 71980 -13140 72020
rect -13360 71910 -13350 71980
rect -13150 71910 -13140 71980
rect -13360 71860 -13140 71910
rect -12860 72090 -12640 72140
rect -12860 72020 -12850 72090
rect -12650 72020 -12640 72090
rect -12860 71980 -12640 72020
rect -12860 71910 -12850 71980
rect -12650 71910 -12640 71980
rect -12860 71860 -12640 71910
rect -12360 72090 -12140 72140
rect -12360 72020 -12350 72090
rect -12150 72020 -12140 72090
rect -12360 71980 -12140 72020
rect -12360 71910 -12350 71980
rect -12150 71910 -12140 71980
rect -12360 71860 -12140 71910
rect 96140 72090 96360 72140
rect 96140 72020 96150 72090
rect 96350 72020 96360 72090
rect 96140 71980 96360 72020
rect 96140 71910 96150 71980
rect 96350 71910 96360 71980
rect 96140 71860 96360 71910
rect 96640 72090 96860 72140
rect 96640 72020 96650 72090
rect 96850 72020 96860 72090
rect 96640 71980 96860 72020
rect 96640 71910 96650 71980
rect 96850 71910 96860 71980
rect 96640 71860 96860 71910
rect 97140 72090 97360 72140
rect 97140 72020 97150 72090
rect 97350 72020 97360 72090
rect 97140 71980 97360 72020
rect 97140 71910 97150 71980
rect 97350 71910 97360 71980
rect 97140 71860 97360 71910
rect 97640 72090 97860 72140
rect 97640 72020 97650 72090
rect 97850 72020 97860 72090
rect 97640 71980 97860 72020
rect 97640 71910 97650 71980
rect 97850 71910 97860 71980
rect 97640 71860 97860 71910
rect 98140 72090 98360 72140
rect 98140 72020 98150 72090
rect 98350 72020 98360 72090
rect 98140 71980 98360 72020
rect 98140 71910 98150 71980
rect 98350 71910 98360 71980
rect 98140 71860 98360 71910
rect 98640 72090 98860 72140
rect 98640 72020 98650 72090
rect 98850 72020 98860 72090
rect 98640 71980 98860 72020
rect 98640 71910 98650 71980
rect 98850 71910 98860 71980
rect 98640 71860 98860 71910
rect 99140 72090 99360 72140
rect 99140 72020 99150 72090
rect 99350 72020 99360 72090
rect 99140 71980 99360 72020
rect 99140 71910 99150 71980
rect 99350 71910 99360 71980
rect 99140 71860 99360 71910
rect 99640 72090 99860 72140
rect 99640 72020 99650 72090
rect 99850 72020 99860 72090
rect 99640 71980 99860 72020
rect 99640 71910 99650 71980
rect 99850 71910 99860 71980
rect 99640 71860 99860 71910
rect -16000 71850 -12000 71860
rect -16000 71650 -15980 71850
rect -15910 71650 -15590 71850
rect -15520 71650 -15480 71850
rect -15410 71650 -15090 71850
rect -15020 71650 -14980 71850
rect -14910 71650 -14590 71850
rect -14520 71650 -14480 71850
rect -14410 71650 -14090 71850
rect -14020 71650 -13980 71850
rect -13910 71650 -13590 71850
rect -13520 71650 -13480 71850
rect -13410 71650 -13090 71850
rect -13020 71650 -12980 71850
rect -12910 71650 -12590 71850
rect -12520 71650 -12480 71850
rect -12410 71650 -12090 71850
rect -12020 71650 -12000 71850
rect -16000 71640 -12000 71650
rect 96000 71850 100000 71860
rect 96000 71650 96020 71850
rect 96090 71650 96410 71850
rect 96480 71650 96520 71850
rect 96590 71650 96910 71850
rect 96980 71650 97020 71850
rect 97090 71650 97410 71850
rect 97480 71650 97520 71850
rect 97590 71650 97910 71850
rect 97980 71650 98020 71850
rect 98090 71650 98410 71850
rect 98480 71650 98520 71850
rect 98590 71650 98910 71850
rect 98980 71650 99020 71850
rect 99090 71650 99410 71850
rect 99480 71650 99520 71850
rect 99590 71650 99910 71850
rect 99980 71650 100000 71850
rect 96000 71640 100000 71650
rect -15860 71590 -15640 71640
rect -15860 71520 -15850 71590
rect -15650 71520 -15640 71590
rect -15860 71480 -15640 71520
rect -15860 71410 -15850 71480
rect -15650 71410 -15640 71480
rect -15860 71360 -15640 71410
rect -15360 71590 -15140 71640
rect -15360 71520 -15350 71590
rect -15150 71520 -15140 71590
rect -15360 71480 -15140 71520
rect -15360 71410 -15350 71480
rect -15150 71410 -15140 71480
rect -15360 71360 -15140 71410
rect -14860 71590 -14640 71640
rect -14860 71520 -14850 71590
rect -14650 71520 -14640 71590
rect -14860 71480 -14640 71520
rect -14860 71410 -14850 71480
rect -14650 71410 -14640 71480
rect -14860 71360 -14640 71410
rect -14360 71590 -14140 71640
rect -14360 71520 -14350 71590
rect -14150 71520 -14140 71590
rect -14360 71480 -14140 71520
rect -14360 71410 -14350 71480
rect -14150 71410 -14140 71480
rect -14360 71360 -14140 71410
rect -13860 71590 -13640 71640
rect -13860 71520 -13850 71590
rect -13650 71520 -13640 71590
rect -13860 71480 -13640 71520
rect -13860 71410 -13850 71480
rect -13650 71410 -13640 71480
rect -13860 71360 -13640 71410
rect -13360 71590 -13140 71640
rect -13360 71520 -13350 71590
rect -13150 71520 -13140 71590
rect -13360 71480 -13140 71520
rect -13360 71410 -13350 71480
rect -13150 71410 -13140 71480
rect -13360 71360 -13140 71410
rect -12860 71590 -12640 71640
rect -12860 71520 -12850 71590
rect -12650 71520 -12640 71590
rect -12860 71480 -12640 71520
rect -12860 71410 -12850 71480
rect -12650 71410 -12640 71480
rect -12860 71360 -12640 71410
rect -12360 71590 -12140 71640
rect -12360 71520 -12350 71590
rect -12150 71520 -12140 71590
rect -12360 71480 -12140 71520
rect -12360 71410 -12350 71480
rect -12150 71410 -12140 71480
rect -12360 71360 -12140 71410
rect 96140 71590 96360 71640
rect 96140 71520 96150 71590
rect 96350 71520 96360 71590
rect 96140 71480 96360 71520
rect 96140 71410 96150 71480
rect 96350 71410 96360 71480
rect 96140 71360 96360 71410
rect 96640 71590 96860 71640
rect 96640 71520 96650 71590
rect 96850 71520 96860 71590
rect 96640 71480 96860 71520
rect 96640 71410 96650 71480
rect 96850 71410 96860 71480
rect 96640 71360 96860 71410
rect 97140 71590 97360 71640
rect 97140 71520 97150 71590
rect 97350 71520 97360 71590
rect 97140 71480 97360 71520
rect 97140 71410 97150 71480
rect 97350 71410 97360 71480
rect 97140 71360 97360 71410
rect 97640 71590 97860 71640
rect 97640 71520 97650 71590
rect 97850 71520 97860 71590
rect 97640 71480 97860 71520
rect 97640 71410 97650 71480
rect 97850 71410 97860 71480
rect 97640 71360 97860 71410
rect 98140 71590 98360 71640
rect 98140 71520 98150 71590
rect 98350 71520 98360 71590
rect 98140 71480 98360 71520
rect 98140 71410 98150 71480
rect 98350 71410 98360 71480
rect 98140 71360 98360 71410
rect 98640 71590 98860 71640
rect 98640 71520 98650 71590
rect 98850 71520 98860 71590
rect 98640 71480 98860 71520
rect 98640 71410 98650 71480
rect 98850 71410 98860 71480
rect 98640 71360 98860 71410
rect 99140 71590 99360 71640
rect 99140 71520 99150 71590
rect 99350 71520 99360 71590
rect 99140 71480 99360 71520
rect 99140 71410 99150 71480
rect 99350 71410 99360 71480
rect 99140 71360 99360 71410
rect 99640 71590 99860 71640
rect 99640 71520 99650 71590
rect 99850 71520 99860 71590
rect 99640 71480 99860 71520
rect 99640 71410 99650 71480
rect 99850 71410 99860 71480
rect 99640 71360 99860 71410
rect -16000 71350 -12000 71360
rect -16000 71150 -15980 71350
rect -15910 71150 -15590 71350
rect -15520 71150 -15480 71350
rect -15410 71150 -15090 71350
rect -15020 71150 -14980 71350
rect -14910 71150 -14590 71350
rect -14520 71150 -14480 71350
rect -14410 71150 -14090 71350
rect -14020 71150 -13980 71350
rect -13910 71150 -13590 71350
rect -13520 71150 -13480 71350
rect -13410 71150 -13090 71350
rect -13020 71150 -12980 71350
rect -12910 71150 -12590 71350
rect -12520 71150 -12480 71350
rect -12410 71150 -12090 71350
rect -12020 71150 -12000 71350
rect -16000 71140 -12000 71150
rect 96000 71350 100000 71360
rect 96000 71150 96020 71350
rect 96090 71150 96410 71350
rect 96480 71150 96520 71350
rect 96590 71150 96910 71350
rect 96980 71150 97020 71350
rect 97090 71150 97410 71350
rect 97480 71150 97520 71350
rect 97590 71150 97910 71350
rect 97980 71150 98020 71350
rect 98090 71150 98410 71350
rect 98480 71150 98520 71350
rect 98590 71150 98910 71350
rect 98980 71150 99020 71350
rect 99090 71150 99410 71350
rect 99480 71150 99520 71350
rect 99590 71150 99910 71350
rect 99980 71150 100000 71350
rect 96000 71140 100000 71150
rect -15860 71090 -15640 71140
rect -15860 71020 -15850 71090
rect -15650 71020 -15640 71090
rect -15860 70980 -15640 71020
rect -15860 70910 -15850 70980
rect -15650 70910 -15640 70980
rect -15860 70860 -15640 70910
rect -15360 71090 -15140 71140
rect -15360 71020 -15350 71090
rect -15150 71020 -15140 71090
rect -15360 70980 -15140 71020
rect -15360 70910 -15350 70980
rect -15150 70910 -15140 70980
rect -15360 70860 -15140 70910
rect -14860 71090 -14640 71140
rect -14860 71020 -14850 71090
rect -14650 71020 -14640 71090
rect -14860 70980 -14640 71020
rect -14860 70910 -14850 70980
rect -14650 70910 -14640 70980
rect -14860 70860 -14640 70910
rect -14360 71090 -14140 71140
rect -14360 71020 -14350 71090
rect -14150 71020 -14140 71090
rect -14360 70980 -14140 71020
rect -14360 70910 -14350 70980
rect -14150 70910 -14140 70980
rect -14360 70860 -14140 70910
rect -13860 71090 -13640 71140
rect -13860 71020 -13850 71090
rect -13650 71020 -13640 71090
rect -13860 70980 -13640 71020
rect -13860 70910 -13850 70980
rect -13650 70910 -13640 70980
rect -13860 70860 -13640 70910
rect -13360 71090 -13140 71140
rect -13360 71020 -13350 71090
rect -13150 71020 -13140 71090
rect -13360 70980 -13140 71020
rect -13360 70910 -13350 70980
rect -13150 70910 -13140 70980
rect -13360 70860 -13140 70910
rect -12860 71090 -12640 71140
rect -12860 71020 -12850 71090
rect -12650 71020 -12640 71090
rect -12860 70980 -12640 71020
rect -12860 70910 -12850 70980
rect -12650 70910 -12640 70980
rect -12860 70860 -12640 70910
rect -12360 71090 -12140 71140
rect -12360 71020 -12350 71090
rect -12150 71020 -12140 71090
rect -12360 70980 -12140 71020
rect -12360 70910 -12350 70980
rect -12150 70910 -12140 70980
rect -12360 70860 -12140 70910
rect 96140 71090 96360 71140
rect 96140 71020 96150 71090
rect 96350 71020 96360 71090
rect 96140 70980 96360 71020
rect 96140 70910 96150 70980
rect 96350 70910 96360 70980
rect 96140 70860 96360 70910
rect 96640 71090 96860 71140
rect 96640 71020 96650 71090
rect 96850 71020 96860 71090
rect 96640 70980 96860 71020
rect 96640 70910 96650 70980
rect 96850 70910 96860 70980
rect 96640 70860 96860 70910
rect 97140 71090 97360 71140
rect 97140 71020 97150 71090
rect 97350 71020 97360 71090
rect 97140 70980 97360 71020
rect 97140 70910 97150 70980
rect 97350 70910 97360 70980
rect 97140 70860 97360 70910
rect 97640 71090 97860 71140
rect 97640 71020 97650 71090
rect 97850 71020 97860 71090
rect 97640 70980 97860 71020
rect 97640 70910 97650 70980
rect 97850 70910 97860 70980
rect 97640 70860 97860 70910
rect 98140 71090 98360 71140
rect 98140 71020 98150 71090
rect 98350 71020 98360 71090
rect 98140 70980 98360 71020
rect 98140 70910 98150 70980
rect 98350 70910 98360 70980
rect 98140 70860 98360 70910
rect 98640 71090 98860 71140
rect 98640 71020 98650 71090
rect 98850 71020 98860 71090
rect 98640 70980 98860 71020
rect 98640 70910 98650 70980
rect 98850 70910 98860 70980
rect 98640 70860 98860 70910
rect 99140 71090 99360 71140
rect 99140 71020 99150 71090
rect 99350 71020 99360 71090
rect 99140 70980 99360 71020
rect 99140 70910 99150 70980
rect 99350 70910 99360 70980
rect 99140 70860 99360 70910
rect 99640 71090 99860 71140
rect 99640 71020 99650 71090
rect 99850 71020 99860 71090
rect 99640 70980 99860 71020
rect 99640 70910 99650 70980
rect 99850 70910 99860 70980
rect 99640 70860 99860 70910
rect -16000 70850 -12000 70860
rect -16000 70650 -15980 70850
rect -15910 70650 -15590 70850
rect -15520 70650 -15480 70850
rect -15410 70650 -15090 70850
rect -15020 70650 -14980 70850
rect -14910 70650 -14590 70850
rect -14520 70650 -14480 70850
rect -14410 70650 -14090 70850
rect -14020 70650 -13980 70850
rect -13910 70650 -13590 70850
rect -13520 70650 -13480 70850
rect -13410 70650 -13090 70850
rect -13020 70650 -12980 70850
rect -12910 70650 -12590 70850
rect -12520 70650 -12480 70850
rect -12410 70650 -12090 70850
rect -12020 70650 -12000 70850
rect -16000 70640 -12000 70650
rect 96000 70850 100000 70860
rect 96000 70650 96020 70850
rect 96090 70650 96410 70850
rect 96480 70650 96520 70850
rect 96590 70650 96910 70850
rect 96980 70650 97020 70850
rect 97090 70650 97410 70850
rect 97480 70650 97520 70850
rect 97590 70650 97910 70850
rect 97980 70650 98020 70850
rect 98090 70650 98410 70850
rect 98480 70650 98520 70850
rect 98590 70650 98910 70850
rect 98980 70650 99020 70850
rect 99090 70650 99410 70850
rect 99480 70650 99520 70850
rect 99590 70650 99910 70850
rect 99980 70650 100000 70850
rect 96000 70640 100000 70650
rect -15860 70590 -15640 70640
rect -15860 70520 -15850 70590
rect -15650 70520 -15640 70590
rect -15860 70480 -15640 70520
rect -15860 70410 -15850 70480
rect -15650 70410 -15640 70480
rect -15860 70360 -15640 70410
rect -15360 70590 -15140 70640
rect -15360 70520 -15350 70590
rect -15150 70520 -15140 70590
rect -15360 70480 -15140 70520
rect -15360 70410 -15350 70480
rect -15150 70410 -15140 70480
rect -15360 70360 -15140 70410
rect -14860 70590 -14640 70640
rect -14860 70520 -14850 70590
rect -14650 70520 -14640 70590
rect -14860 70480 -14640 70520
rect -14860 70410 -14850 70480
rect -14650 70410 -14640 70480
rect -14860 70360 -14640 70410
rect -14360 70590 -14140 70640
rect -14360 70520 -14350 70590
rect -14150 70520 -14140 70590
rect -14360 70480 -14140 70520
rect -14360 70410 -14350 70480
rect -14150 70410 -14140 70480
rect -14360 70360 -14140 70410
rect -13860 70590 -13640 70640
rect -13860 70520 -13850 70590
rect -13650 70520 -13640 70590
rect -13860 70480 -13640 70520
rect -13860 70410 -13850 70480
rect -13650 70410 -13640 70480
rect -13860 70360 -13640 70410
rect -13360 70590 -13140 70640
rect -13360 70520 -13350 70590
rect -13150 70520 -13140 70590
rect -13360 70480 -13140 70520
rect -13360 70410 -13350 70480
rect -13150 70410 -13140 70480
rect -13360 70360 -13140 70410
rect -12860 70590 -12640 70640
rect -12860 70520 -12850 70590
rect -12650 70520 -12640 70590
rect -12860 70480 -12640 70520
rect -12860 70410 -12850 70480
rect -12650 70410 -12640 70480
rect -12860 70360 -12640 70410
rect -12360 70590 -12140 70640
rect -12360 70520 -12350 70590
rect -12150 70520 -12140 70590
rect -12360 70480 -12140 70520
rect -12360 70410 -12350 70480
rect -12150 70410 -12140 70480
rect -12360 70360 -12140 70410
rect 96140 70590 96360 70640
rect 96140 70520 96150 70590
rect 96350 70520 96360 70590
rect 96140 70480 96360 70520
rect 96140 70410 96150 70480
rect 96350 70410 96360 70480
rect 96140 70360 96360 70410
rect 96640 70590 96860 70640
rect 96640 70520 96650 70590
rect 96850 70520 96860 70590
rect 96640 70480 96860 70520
rect 96640 70410 96650 70480
rect 96850 70410 96860 70480
rect 96640 70360 96860 70410
rect 97140 70590 97360 70640
rect 97140 70520 97150 70590
rect 97350 70520 97360 70590
rect 97140 70480 97360 70520
rect 97140 70410 97150 70480
rect 97350 70410 97360 70480
rect 97140 70360 97360 70410
rect 97640 70590 97860 70640
rect 97640 70520 97650 70590
rect 97850 70520 97860 70590
rect 97640 70480 97860 70520
rect 97640 70410 97650 70480
rect 97850 70410 97860 70480
rect 97640 70360 97860 70410
rect 98140 70590 98360 70640
rect 98140 70520 98150 70590
rect 98350 70520 98360 70590
rect 98140 70480 98360 70520
rect 98140 70410 98150 70480
rect 98350 70410 98360 70480
rect 98140 70360 98360 70410
rect 98640 70590 98860 70640
rect 98640 70520 98650 70590
rect 98850 70520 98860 70590
rect 98640 70480 98860 70520
rect 98640 70410 98650 70480
rect 98850 70410 98860 70480
rect 98640 70360 98860 70410
rect 99140 70590 99360 70640
rect 99140 70520 99150 70590
rect 99350 70520 99360 70590
rect 99140 70480 99360 70520
rect 99140 70410 99150 70480
rect 99350 70410 99360 70480
rect 99140 70360 99360 70410
rect 99640 70590 99860 70640
rect 99640 70520 99650 70590
rect 99850 70520 99860 70590
rect 99640 70480 99860 70520
rect 99640 70410 99650 70480
rect 99850 70410 99860 70480
rect 99640 70360 99860 70410
rect -16000 70350 -12000 70360
rect -16000 70150 -15980 70350
rect -15910 70150 -15590 70350
rect -15520 70150 -15480 70350
rect -15410 70150 -15090 70350
rect -15020 70150 -14980 70350
rect -14910 70150 -14590 70350
rect -14520 70150 -14480 70350
rect -14410 70150 -14090 70350
rect -14020 70150 -13980 70350
rect -13910 70150 -13590 70350
rect -13520 70150 -13480 70350
rect -13410 70150 -13090 70350
rect -13020 70150 -12980 70350
rect -12910 70150 -12590 70350
rect -12520 70150 -12480 70350
rect -12410 70150 -12090 70350
rect -12020 70150 -12000 70350
rect -16000 70140 -12000 70150
rect 96000 70350 100000 70360
rect 96000 70150 96020 70350
rect 96090 70150 96410 70350
rect 96480 70150 96520 70350
rect 96590 70150 96910 70350
rect 96980 70150 97020 70350
rect 97090 70150 97410 70350
rect 97480 70150 97520 70350
rect 97590 70150 97910 70350
rect 97980 70150 98020 70350
rect 98090 70150 98410 70350
rect 98480 70150 98520 70350
rect 98590 70150 98910 70350
rect 98980 70150 99020 70350
rect 99090 70150 99410 70350
rect 99480 70150 99520 70350
rect 99590 70150 99910 70350
rect 99980 70150 100000 70350
rect 96000 70140 100000 70150
rect -15860 70090 -15640 70140
rect -15860 70020 -15850 70090
rect -15650 70020 -15640 70090
rect -15860 69980 -15640 70020
rect -15860 69910 -15850 69980
rect -15650 69910 -15640 69980
rect -15860 69860 -15640 69910
rect -15360 70090 -15140 70140
rect -15360 70020 -15350 70090
rect -15150 70020 -15140 70090
rect -15360 69980 -15140 70020
rect -15360 69910 -15350 69980
rect -15150 69910 -15140 69980
rect -15360 69860 -15140 69910
rect -14860 70090 -14640 70140
rect -14860 70020 -14850 70090
rect -14650 70020 -14640 70090
rect -14860 69980 -14640 70020
rect -14860 69910 -14850 69980
rect -14650 69910 -14640 69980
rect -14860 69860 -14640 69910
rect -14360 70090 -14140 70140
rect -14360 70020 -14350 70090
rect -14150 70020 -14140 70090
rect -14360 69980 -14140 70020
rect -14360 69910 -14350 69980
rect -14150 69910 -14140 69980
rect -14360 69860 -14140 69910
rect -13860 70090 -13640 70140
rect -13860 70020 -13850 70090
rect -13650 70020 -13640 70090
rect -13860 69980 -13640 70020
rect -13860 69910 -13850 69980
rect -13650 69910 -13640 69980
rect -13860 69860 -13640 69910
rect -13360 70090 -13140 70140
rect -13360 70020 -13350 70090
rect -13150 70020 -13140 70090
rect -13360 69980 -13140 70020
rect -13360 69910 -13350 69980
rect -13150 69910 -13140 69980
rect -13360 69860 -13140 69910
rect -12860 70090 -12640 70140
rect -12860 70020 -12850 70090
rect -12650 70020 -12640 70090
rect -12860 69980 -12640 70020
rect -12860 69910 -12850 69980
rect -12650 69910 -12640 69980
rect -12860 69860 -12640 69910
rect -12360 70090 -12140 70140
rect -12360 70020 -12350 70090
rect -12150 70020 -12140 70090
rect -12360 69980 -12140 70020
rect -12360 69910 -12350 69980
rect -12150 69910 -12140 69980
rect -12360 69860 -12140 69910
rect 96140 70090 96360 70140
rect 96140 70020 96150 70090
rect 96350 70020 96360 70090
rect 96140 69980 96360 70020
rect 96140 69910 96150 69980
rect 96350 69910 96360 69980
rect 96140 69860 96360 69910
rect 96640 70090 96860 70140
rect 96640 70020 96650 70090
rect 96850 70020 96860 70090
rect 96640 69980 96860 70020
rect 96640 69910 96650 69980
rect 96850 69910 96860 69980
rect 96640 69860 96860 69910
rect 97140 70090 97360 70140
rect 97140 70020 97150 70090
rect 97350 70020 97360 70090
rect 97140 69980 97360 70020
rect 97140 69910 97150 69980
rect 97350 69910 97360 69980
rect 97140 69860 97360 69910
rect 97640 70090 97860 70140
rect 97640 70020 97650 70090
rect 97850 70020 97860 70090
rect 97640 69980 97860 70020
rect 97640 69910 97650 69980
rect 97850 69910 97860 69980
rect 97640 69860 97860 69910
rect 98140 70090 98360 70140
rect 98140 70020 98150 70090
rect 98350 70020 98360 70090
rect 98140 69980 98360 70020
rect 98140 69910 98150 69980
rect 98350 69910 98360 69980
rect 98140 69860 98360 69910
rect 98640 70090 98860 70140
rect 98640 70020 98650 70090
rect 98850 70020 98860 70090
rect 98640 69980 98860 70020
rect 98640 69910 98650 69980
rect 98850 69910 98860 69980
rect 98640 69860 98860 69910
rect 99140 70090 99360 70140
rect 99140 70020 99150 70090
rect 99350 70020 99360 70090
rect 99140 69980 99360 70020
rect 99140 69910 99150 69980
rect 99350 69910 99360 69980
rect 99140 69860 99360 69910
rect 99640 70090 99860 70140
rect 99640 70020 99650 70090
rect 99850 70020 99860 70090
rect 99640 69980 99860 70020
rect 99640 69910 99650 69980
rect 99850 69910 99860 69980
rect 99640 69860 99860 69910
rect -16000 69850 -12000 69860
rect -16000 69650 -15980 69850
rect -15910 69650 -15590 69850
rect -15520 69650 -15480 69850
rect -15410 69650 -15090 69850
rect -15020 69650 -14980 69850
rect -14910 69650 -14590 69850
rect -14520 69650 -14480 69850
rect -14410 69650 -14090 69850
rect -14020 69650 -13980 69850
rect -13910 69650 -13590 69850
rect -13520 69650 -13480 69850
rect -13410 69650 -13090 69850
rect -13020 69650 -12980 69850
rect -12910 69650 -12590 69850
rect -12520 69650 -12480 69850
rect -12410 69650 -12090 69850
rect -12020 69650 -12000 69850
rect -16000 69640 -12000 69650
rect 96000 69850 100000 69860
rect 96000 69650 96020 69850
rect 96090 69650 96410 69850
rect 96480 69650 96520 69850
rect 96590 69650 96910 69850
rect 96980 69650 97020 69850
rect 97090 69650 97410 69850
rect 97480 69650 97520 69850
rect 97590 69650 97910 69850
rect 97980 69650 98020 69850
rect 98090 69650 98410 69850
rect 98480 69650 98520 69850
rect 98590 69650 98910 69850
rect 98980 69650 99020 69850
rect 99090 69650 99410 69850
rect 99480 69650 99520 69850
rect 99590 69650 99910 69850
rect 99980 69650 100000 69850
rect 96000 69640 100000 69650
rect -15860 69590 -15640 69640
rect -15860 69520 -15850 69590
rect -15650 69520 -15640 69590
rect -15860 69480 -15640 69520
rect -15860 69410 -15850 69480
rect -15650 69410 -15640 69480
rect -15860 69360 -15640 69410
rect -15360 69590 -15140 69640
rect -15360 69520 -15350 69590
rect -15150 69520 -15140 69590
rect -15360 69480 -15140 69520
rect -15360 69410 -15350 69480
rect -15150 69410 -15140 69480
rect -15360 69360 -15140 69410
rect -14860 69590 -14640 69640
rect -14860 69520 -14850 69590
rect -14650 69520 -14640 69590
rect -14860 69480 -14640 69520
rect -14860 69410 -14850 69480
rect -14650 69410 -14640 69480
rect -14860 69360 -14640 69410
rect -14360 69590 -14140 69640
rect -14360 69520 -14350 69590
rect -14150 69520 -14140 69590
rect -14360 69480 -14140 69520
rect -14360 69410 -14350 69480
rect -14150 69410 -14140 69480
rect -14360 69360 -14140 69410
rect -13860 69590 -13640 69640
rect -13860 69520 -13850 69590
rect -13650 69520 -13640 69590
rect -13860 69480 -13640 69520
rect -13860 69410 -13850 69480
rect -13650 69410 -13640 69480
rect -13860 69360 -13640 69410
rect -13360 69590 -13140 69640
rect -13360 69520 -13350 69590
rect -13150 69520 -13140 69590
rect -13360 69480 -13140 69520
rect -13360 69410 -13350 69480
rect -13150 69410 -13140 69480
rect -13360 69360 -13140 69410
rect -12860 69590 -12640 69640
rect -12860 69520 -12850 69590
rect -12650 69520 -12640 69590
rect -12860 69480 -12640 69520
rect -12860 69410 -12850 69480
rect -12650 69410 -12640 69480
rect -12860 69360 -12640 69410
rect -12360 69590 -12140 69640
rect -12360 69520 -12350 69590
rect -12150 69520 -12140 69590
rect -12360 69480 -12140 69520
rect -12360 69410 -12350 69480
rect -12150 69410 -12140 69480
rect -12360 69360 -12140 69410
rect 96140 69590 96360 69640
rect 96140 69520 96150 69590
rect 96350 69520 96360 69590
rect 96140 69480 96360 69520
rect 96140 69410 96150 69480
rect 96350 69410 96360 69480
rect 96140 69360 96360 69410
rect 96640 69590 96860 69640
rect 96640 69520 96650 69590
rect 96850 69520 96860 69590
rect 96640 69480 96860 69520
rect 96640 69410 96650 69480
rect 96850 69410 96860 69480
rect 96640 69360 96860 69410
rect 97140 69590 97360 69640
rect 97140 69520 97150 69590
rect 97350 69520 97360 69590
rect 97140 69480 97360 69520
rect 97140 69410 97150 69480
rect 97350 69410 97360 69480
rect 97140 69360 97360 69410
rect 97640 69590 97860 69640
rect 97640 69520 97650 69590
rect 97850 69520 97860 69590
rect 97640 69480 97860 69520
rect 97640 69410 97650 69480
rect 97850 69410 97860 69480
rect 97640 69360 97860 69410
rect 98140 69590 98360 69640
rect 98140 69520 98150 69590
rect 98350 69520 98360 69590
rect 98140 69480 98360 69520
rect 98140 69410 98150 69480
rect 98350 69410 98360 69480
rect 98140 69360 98360 69410
rect 98640 69590 98860 69640
rect 98640 69520 98650 69590
rect 98850 69520 98860 69590
rect 98640 69480 98860 69520
rect 98640 69410 98650 69480
rect 98850 69410 98860 69480
rect 98640 69360 98860 69410
rect 99140 69590 99360 69640
rect 99140 69520 99150 69590
rect 99350 69520 99360 69590
rect 99140 69480 99360 69520
rect 99140 69410 99150 69480
rect 99350 69410 99360 69480
rect 99140 69360 99360 69410
rect 99640 69590 99860 69640
rect 99640 69520 99650 69590
rect 99850 69520 99860 69590
rect 99640 69480 99860 69520
rect 99640 69410 99650 69480
rect 99850 69410 99860 69480
rect 99640 69360 99860 69410
rect -16000 69350 -12000 69360
rect -16000 69150 -15980 69350
rect -15910 69150 -15590 69350
rect -15520 69150 -15480 69350
rect -15410 69150 -15090 69350
rect -15020 69150 -14980 69350
rect -14910 69150 -14590 69350
rect -14520 69150 -14480 69350
rect -14410 69150 -14090 69350
rect -14020 69150 -13980 69350
rect -13910 69150 -13590 69350
rect -13520 69150 -13480 69350
rect -13410 69150 -13090 69350
rect -13020 69150 -12980 69350
rect -12910 69150 -12590 69350
rect -12520 69150 -12480 69350
rect -12410 69150 -12090 69350
rect -12020 69150 -12000 69350
rect -16000 69140 -12000 69150
rect 96000 69350 100000 69360
rect 96000 69150 96020 69350
rect 96090 69150 96410 69350
rect 96480 69150 96520 69350
rect 96590 69150 96910 69350
rect 96980 69150 97020 69350
rect 97090 69150 97410 69350
rect 97480 69150 97520 69350
rect 97590 69150 97910 69350
rect 97980 69150 98020 69350
rect 98090 69150 98410 69350
rect 98480 69150 98520 69350
rect 98590 69150 98910 69350
rect 98980 69150 99020 69350
rect 99090 69150 99410 69350
rect 99480 69150 99520 69350
rect 99590 69150 99910 69350
rect 99980 69150 100000 69350
rect 96000 69140 100000 69150
rect -15860 69090 -15640 69140
rect -15860 69020 -15850 69090
rect -15650 69020 -15640 69090
rect -15860 68980 -15640 69020
rect -15860 68910 -15850 68980
rect -15650 68910 -15640 68980
rect -15860 68860 -15640 68910
rect -15360 69090 -15140 69140
rect -15360 69020 -15350 69090
rect -15150 69020 -15140 69090
rect -15360 68980 -15140 69020
rect -15360 68910 -15350 68980
rect -15150 68910 -15140 68980
rect -15360 68860 -15140 68910
rect -14860 69090 -14640 69140
rect -14860 69020 -14850 69090
rect -14650 69020 -14640 69090
rect -14860 68980 -14640 69020
rect -14860 68910 -14850 68980
rect -14650 68910 -14640 68980
rect -14860 68860 -14640 68910
rect -14360 69090 -14140 69140
rect -14360 69020 -14350 69090
rect -14150 69020 -14140 69090
rect -14360 68980 -14140 69020
rect -14360 68910 -14350 68980
rect -14150 68910 -14140 68980
rect -14360 68860 -14140 68910
rect -13860 69090 -13640 69140
rect -13860 69020 -13850 69090
rect -13650 69020 -13640 69090
rect -13860 68980 -13640 69020
rect -13860 68910 -13850 68980
rect -13650 68910 -13640 68980
rect -13860 68860 -13640 68910
rect -13360 69090 -13140 69140
rect -13360 69020 -13350 69090
rect -13150 69020 -13140 69090
rect -13360 68980 -13140 69020
rect -13360 68910 -13350 68980
rect -13150 68910 -13140 68980
rect -13360 68860 -13140 68910
rect -12860 69090 -12640 69140
rect -12860 69020 -12850 69090
rect -12650 69020 -12640 69090
rect -12860 68980 -12640 69020
rect -12860 68910 -12850 68980
rect -12650 68910 -12640 68980
rect -12860 68860 -12640 68910
rect -12360 69090 -12140 69140
rect -12360 69020 -12350 69090
rect -12150 69020 -12140 69090
rect -12360 68980 -12140 69020
rect -12360 68910 -12350 68980
rect -12150 68910 -12140 68980
rect -12360 68860 -12140 68910
rect 96140 69090 96360 69140
rect 96140 69020 96150 69090
rect 96350 69020 96360 69090
rect 96140 68980 96360 69020
rect 96140 68910 96150 68980
rect 96350 68910 96360 68980
rect 96140 68860 96360 68910
rect 96640 69090 96860 69140
rect 96640 69020 96650 69090
rect 96850 69020 96860 69090
rect 96640 68980 96860 69020
rect 96640 68910 96650 68980
rect 96850 68910 96860 68980
rect 96640 68860 96860 68910
rect 97140 69090 97360 69140
rect 97140 69020 97150 69090
rect 97350 69020 97360 69090
rect 97140 68980 97360 69020
rect 97140 68910 97150 68980
rect 97350 68910 97360 68980
rect 97140 68860 97360 68910
rect 97640 69090 97860 69140
rect 97640 69020 97650 69090
rect 97850 69020 97860 69090
rect 97640 68980 97860 69020
rect 97640 68910 97650 68980
rect 97850 68910 97860 68980
rect 97640 68860 97860 68910
rect 98140 69090 98360 69140
rect 98140 69020 98150 69090
rect 98350 69020 98360 69090
rect 98140 68980 98360 69020
rect 98140 68910 98150 68980
rect 98350 68910 98360 68980
rect 98140 68860 98360 68910
rect 98640 69090 98860 69140
rect 98640 69020 98650 69090
rect 98850 69020 98860 69090
rect 98640 68980 98860 69020
rect 98640 68910 98650 68980
rect 98850 68910 98860 68980
rect 98640 68860 98860 68910
rect 99140 69090 99360 69140
rect 99140 69020 99150 69090
rect 99350 69020 99360 69090
rect 99140 68980 99360 69020
rect 99140 68910 99150 68980
rect 99350 68910 99360 68980
rect 99140 68860 99360 68910
rect 99640 69090 99860 69140
rect 99640 69020 99650 69090
rect 99850 69020 99860 69090
rect 99640 68980 99860 69020
rect 99640 68910 99650 68980
rect 99850 68910 99860 68980
rect 99640 68860 99860 68910
rect -16000 68850 -12000 68860
rect -16000 68650 -15980 68850
rect -15910 68650 -15590 68850
rect -15520 68650 -15480 68850
rect -15410 68650 -15090 68850
rect -15020 68650 -14980 68850
rect -14910 68650 -14590 68850
rect -14520 68650 -14480 68850
rect -14410 68650 -14090 68850
rect -14020 68650 -13980 68850
rect -13910 68650 -13590 68850
rect -13520 68650 -13480 68850
rect -13410 68650 -13090 68850
rect -13020 68650 -12980 68850
rect -12910 68650 -12590 68850
rect -12520 68650 -12480 68850
rect -12410 68650 -12090 68850
rect -12020 68650 -12000 68850
rect -16000 68640 -12000 68650
rect 96000 68850 100000 68860
rect 96000 68650 96020 68850
rect 96090 68650 96410 68850
rect 96480 68650 96520 68850
rect 96590 68650 96910 68850
rect 96980 68650 97020 68850
rect 97090 68650 97410 68850
rect 97480 68650 97520 68850
rect 97590 68650 97910 68850
rect 97980 68650 98020 68850
rect 98090 68650 98410 68850
rect 98480 68650 98520 68850
rect 98590 68650 98910 68850
rect 98980 68650 99020 68850
rect 99090 68650 99410 68850
rect 99480 68650 99520 68850
rect 99590 68650 99910 68850
rect 99980 68650 100000 68850
rect 96000 68640 100000 68650
rect -15860 68590 -15640 68640
rect -15860 68520 -15850 68590
rect -15650 68520 -15640 68590
rect -15860 68480 -15640 68520
rect -15860 68410 -15850 68480
rect -15650 68410 -15640 68480
rect -15860 68360 -15640 68410
rect -15360 68590 -15140 68640
rect -15360 68520 -15350 68590
rect -15150 68520 -15140 68590
rect -15360 68480 -15140 68520
rect -15360 68410 -15350 68480
rect -15150 68410 -15140 68480
rect -15360 68360 -15140 68410
rect -14860 68590 -14640 68640
rect -14860 68520 -14850 68590
rect -14650 68520 -14640 68590
rect -14860 68480 -14640 68520
rect -14860 68410 -14850 68480
rect -14650 68410 -14640 68480
rect -14860 68360 -14640 68410
rect -14360 68590 -14140 68640
rect -14360 68520 -14350 68590
rect -14150 68520 -14140 68590
rect -14360 68480 -14140 68520
rect -14360 68410 -14350 68480
rect -14150 68410 -14140 68480
rect -14360 68360 -14140 68410
rect -13860 68590 -13640 68640
rect -13860 68520 -13850 68590
rect -13650 68520 -13640 68590
rect -13860 68480 -13640 68520
rect -13860 68410 -13850 68480
rect -13650 68410 -13640 68480
rect -13860 68360 -13640 68410
rect -13360 68590 -13140 68640
rect -13360 68520 -13350 68590
rect -13150 68520 -13140 68590
rect -13360 68480 -13140 68520
rect -13360 68410 -13350 68480
rect -13150 68410 -13140 68480
rect -13360 68360 -13140 68410
rect -12860 68590 -12640 68640
rect -12860 68520 -12850 68590
rect -12650 68520 -12640 68590
rect -12860 68480 -12640 68520
rect -12860 68410 -12850 68480
rect -12650 68410 -12640 68480
rect -12860 68360 -12640 68410
rect -12360 68590 -12140 68640
rect -12360 68520 -12350 68590
rect -12150 68520 -12140 68590
rect -12360 68480 -12140 68520
rect -12360 68410 -12350 68480
rect -12150 68410 -12140 68480
rect -12360 68360 -12140 68410
rect 96140 68590 96360 68640
rect 96140 68520 96150 68590
rect 96350 68520 96360 68590
rect 96140 68480 96360 68520
rect 96140 68410 96150 68480
rect 96350 68410 96360 68480
rect 96140 68360 96360 68410
rect 96640 68590 96860 68640
rect 96640 68520 96650 68590
rect 96850 68520 96860 68590
rect 96640 68480 96860 68520
rect 96640 68410 96650 68480
rect 96850 68410 96860 68480
rect 96640 68360 96860 68410
rect 97140 68590 97360 68640
rect 97140 68520 97150 68590
rect 97350 68520 97360 68590
rect 97140 68480 97360 68520
rect 97140 68410 97150 68480
rect 97350 68410 97360 68480
rect 97140 68360 97360 68410
rect 97640 68590 97860 68640
rect 97640 68520 97650 68590
rect 97850 68520 97860 68590
rect 97640 68480 97860 68520
rect 97640 68410 97650 68480
rect 97850 68410 97860 68480
rect 97640 68360 97860 68410
rect 98140 68590 98360 68640
rect 98140 68520 98150 68590
rect 98350 68520 98360 68590
rect 98140 68480 98360 68520
rect 98140 68410 98150 68480
rect 98350 68410 98360 68480
rect 98140 68360 98360 68410
rect 98640 68590 98860 68640
rect 98640 68520 98650 68590
rect 98850 68520 98860 68590
rect 98640 68480 98860 68520
rect 98640 68410 98650 68480
rect 98850 68410 98860 68480
rect 98640 68360 98860 68410
rect 99140 68590 99360 68640
rect 99140 68520 99150 68590
rect 99350 68520 99360 68590
rect 99140 68480 99360 68520
rect 99140 68410 99150 68480
rect 99350 68410 99360 68480
rect 99140 68360 99360 68410
rect 99640 68590 99860 68640
rect 99640 68520 99650 68590
rect 99850 68520 99860 68590
rect 99640 68480 99860 68520
rect 99640 68410 99650 68480
rect 99850 68410 99860 68480
rect 99640 68360 99860 68410
rect -16000 68350 -12000 68360
rect -16000 68150 -15980 68350
rect -15910 68150 -15590 68350
rect -15520 68150 -15480 68350
rect -15410 68150 -15090 68350
rect -15020 68150 -14980 68350
rect -14910 68150 -14590 68350
rect -14520 68150 -14480 68350
rect -14410 68150 -14090 68350
rect -14020 68150 -13980 68350
rect -13910 68150 -13590 68350
rect -13520 68150 -13480 68350
rect -13410 68150 -13090 68350
rect -13020 68150 -12980 68350
rect -12910 68150 -12590 68350
rect -12520 68150 -12480 68350
rect -12410 68150 -12090 68350
rect -12020 68150 -12000 68350
rect -16000 68140 -12000 68150
rect 96000 68350 100000 68360
rect 96000 68150 96020 68350
rect 96090 68150 96410 68350
rect 96480 68150 96520 68350
rect 96590 68150 96910 68350
rect 96980 68150 97020 68350
rect 97090 68150 97410 68350
rect 97480 68150 97520 68350
rect 97590 68150 97910 68350
rect 97980 68150 98020 68350
rect 98090 68150 98410 68350
rect 98480 68150 98520 68350
rect 98590 68150 98910 68350
rect 98980 68150 99020 68350
rect 99090 68150 99410 68350
rect 99480 68150 99520 68350
rect 99590 68150 99910 68350
rect 99980 68150 100000 68350
rect 96000 68140 100000 68150
rect -15860 68090 -15640 68140
rect -15860 68020 -15850 68090
rect -15650 68020 -15640 68090
rect -15860 67980 -15640 68020
rect -15860 67910 -15850 67980
rect -15650 67910 -15640 67980
rect -15860 67860 -15640 67910
rect -15360 68090 -15140 68140
rect -15360 68020 -15350 68090
rect -15150 68020 -15140 68090
rect -15360 67980 -15140 68020
rect -15360 67910 -15350 67980
rect -15150 67910 -15140 67980
rect -15360 67860 -15140 67910
rect -14860 68090 -14640 68140
rect -14860 68020 -14850 68090
rect -14650 68020 -14640 68090
rect -14860 67980 -14640 68020
rect -14860 67910 -14850 67980
rect -14650 67910 -14640 67980
rect -14860 67860 -14640 67910
rect -14360 68090 -14140 68140
rect -14360 68020 -14350 68090
rect -14150 68020 -14140 68090
rect -14360 67980 -14140 68020
rect -14360 67910 -14350 67980
rect -14150 67910 -14140 67980
rect -14360 67860 -14140 67910
rect -13860 68090 -13640 68140
rect -13860 68020 -13850 68090
rect -13650 68020 -13640 68090
rect -13860 67980 -13640 68020
rect -13860 67910 -13850 67980
rect -13650 67910 -13640 67980
rect -13860 67860 -13640 67910
rect -13360 68090 -13140 68140
rect -13360 68020 -13350 68090
rect -13150 68020 -13140 68090
rect -13360 67980 -13140 68020
rect -13360 67910 -13350 67980
rect -13150 67910 -13140 67980
rect -13360 67860 -13140 67910
rect -12860 68090 -12640 68140
rect -12860 68020 -12850 68090
rect -12650 68020 -12640 68090
rect -12860 67980 -12640 68020
rect -12860 67910 -12850 67980
rect -12650 67910 -12640 67980
rect -12860 67860 -12640 67910
rect -12360 68090 -12140 68140
rect -12360 68020 -12350 68090
rect -12150 68020 -12140 68090
rect -12360 67980 -12140 68020
rect -12360 67910 -12350 67980
rect -12150 67910 -12140 67980
rect -12360 67860 -12140 67910
rect 96140 68090 96360 68140
rect 96140 68020 96150 68090
rect 96350 68020 96360 68090
rect 96140 67980 96360 68020
rect 96140 67910 96150 67980
rect 96350 67910 96360 67980
rect 96140 67860 96360 67910
rect 96640 68090 96860 68140
rect 96640 68020 96650 68090
rect 96850 68020 96860 68090
rect 96640 67980 96860 68020
rect 96640 67910 96650 67980
rect 96850 67910 96860 67980
rect 96640 67860 96860 67910
rect 97140 68090 97360 68140
rect 97140 68020 97150 68090
rect 97350 68020 97360 68090
rect 97140 67980 97360 68020
rect 97140 67910 97150 67980
rect 97350 67910 97360 67980
rect 97140 67860 97360 67910
rect 97640 68090 97860 68140
rect 97640 68020 97650 68090
rect 97850 68020 97860 68090
rect 97640 67980 97860 68020
rect 97640 67910 97650 67980
rect 97850 67910 97860 67980
rect 97640 67860 97860 67910
rect 98140 68090 98360 68140
rect 98140 68020 98150 68090
rect 98350 68020 98360 68090
rect 98140 67980 98360 68020
rect 98140 67910 98150 67980
rect 98350 67910 98360 67980
rect 98140 67860 98360 67910
rect 98640 68090 98860 68140
rect 98640 68020 98650 68090
rect 98850 68020 98860 68090
rect 98640 67980 98860 68020
rect 98640 67910 98650 67980
rect 98850 67910 98860 67980
rect 98640 67860 98860 67910
rect 99140 68090 99360 68140
rect 99140 68020 99150 68090
rect 99350 68020 99360 68090
rect 99140 67980 99360 68020
rect 99140 67910 99150 67980
rect 99350 67910 99360 67980
rect 99140 67860 99360 67910
rect 99640 68090 99860 68140
rect 99640 68020 99650 68090
rect 99850 68020 99860 68090
rect 99640 67980 99860 68020
rect 99640 67910 99650 67980
rect 99850 67910 99860 67980
rect 99640 67860 99860 67910
rect -16000 67850 -12000 67860
rect -16000 67650 -15980 67850
rect -15910 67650 -15590 67850
rect -15520 67650 -15480 67850
rect -15410 67650 -15090 67850
rect -15020 67650 -14980 67850
rect -14910 67650 -14590 67850
rect -14520 67650 -14480 67850
rect -14410 67650 -14090 67850
rect -14020 67650 -13980 67850
rect -13910 67650 -13590 67850
rect -13520 67650 -13480 67850
rect -13410 67650 -13090 67850
rect -13020 67650 -12980 67850
rect -12910 67650 -12590 67850
rect -12520 67650 -12480 67850
rect -12410 67650 -12090 67850
rect -12020 67650 -12000 67850
rect -16000 67640 -12000 67650
rect 96000 67850 100000 67860
rect 96000 67650 96020 67850
rect 96090 67650 96410 67850
rect 96480 67650 96520 67850
rect 96590 67650 96910 67850
rect 96980 67650 97020 67850
rect 97090 67650 97410 67850
rect 97480 67650 97520 67850
rect 97590 67650 97910 67850
rect 97980 67650 98020 67850
rect 98090 67650 98410 67850
rect 98480 67650 98520 67850
rect 98590 67650 98910 67850
rect 98980 67650 99020 67850
rect 99090 67650 99410 67850
rect 99480 67650 99520 67850
rect 99590 67650 99910 67850
rect 99980 67650 100000 67850
rect 96000 67640 100000 67650
rect -15860 67590 -15640 67640
rect -15860 67520 -15850 67590
rect -15650 67520 -15640 67590
rect -15860 67480 -15640 67520
rect -15860 67410 -15850 67480
rect -15650 67410 -15640 67480
rect -15860 67360 -15640 67410
rect -15360 67590 -15140 67640
rect -15360 67520 -15350 67590
rect -15150 67520 -15140 67590
rect -15360 67480 -15140 67520
rect -15360 67410 -15350 67480
rect -15150 67410 -15140 67480
rect -15360 67360 -15140 67410
rect -14860 67590 -14640 67640
rect -14860 67520 -14850 67590
rect -14650 67520 -14640 67590
rect -14860 67480 -14640 67520
rect -14860 67410 -14850 67480
rect -14650 67410 -14640 67480
rect -14860 67360 -14640 67410
rect -14360 67590 -14140 67640
rect -14360 67520 -14350 67590
rect -14150 67520 -14140 67590
rect -14360 67480 -14140 67520
rect -14360 67410 -14350 67480
rect -14150 67410 -14140 67480
rect -14360 67360 -14140 67410
rect -13860 67590 -13640 67640
rect -13860 67520 -13850 67590
rect -13650 67520 -13640 67590
rect -13860 67480 -13640 67520
rect -13860 67410 -13850 67480
rect -13650 67410 -13640 67480
rect -13860 67360 -13640 67410
rect -13360 67590 -13140 67640
rect -13360 67520 -13350 67590
rect -13150 67520 -13140 67590
rect -13360 67480 -13140 67520
rect -13360 67410 -13350 67480
rect -13150 67410 -13140 67480
rect -13360 67360 -13140 67410
rect -12860 67590 -12640 67640
rect -12860 67520 -12850 67590
rect -12650 67520 -12640 67590
rect -12860 67480 -12640 67520
rect -12860 67410 -12850 67480
rect -12650 67410 -12640 67480
rect -12860 67360 -12640 67410
rect -12360 67590 -12140 67640
rect -12360 67520 -12350 67590
rect -12150 67520 -12140 67590
rect -12360 67480 -12140 67520
rect -12360 67410 -12350 67480
rect -12150 67410 -12140 67480
rect -12360 67360 -12140 67410
rect 96140 67590 96360 67640
rect 96140 67520 96150 67590
rect 96350 67520 96360 67590
rect 96140 67480 96360 67520
rect 96140 67410 96150 67480
rect 96350 67410 96360 67480
rect 96140 67360 96360 67410
rect 96640 67590 96860 67640
rect 96640 67520 96650 67590
rect 96850 67520 96860 67590
rect 96640 67480 96860 67520
rect 96640 67410 96650 67480
rect 96850 67410 96860 67480
rect 96640 67360 96860 67410
rect 97140 67590 97360 67640
rect 97140 67520 97150 67590
rect 97350 67520 97360 67590
rect 97140 67480 97360 67520
rect 97140 67410 97150 67480
rect 97350 67410 97360 67480
rect 97140 67360 97360 67410
rect 97640 67590 97860 67640
rect 97640 67520 97650 67590
rect 97850 67520 97860 67590
rect 97640 67480 97860 67520
rect 97640 67410 97650 67480
rect 97850 67410 97860 67480
rect 97640 67360 97860 67410
rect 98140 67590 98360 67640
rect 98140 67520 98150 67590
rect 98350 67520 98360 67590
rect 98140 67480 98360 67520
rect 98140 67410 98150 67480
rect 98350 67410 98360 67480
rect 98140 67360 98360 67410
rect 98640 67590 98860 67640
rect 98640 67520 98650 67590
rect 98850 67520 98860 67590
rect 98640 67480 98860 67520
rect 98640 67410 98650 67480
rect 98850 67410 98860 67480
rect 98640 67360 98860 67410
rect 99140 67590 99360 67640
rect 99140 67520 99150 67590
rect 99350 67520 99360 67590
rect 99140 67480 99360 67520
rect 99140 67410 99150 67480
rect 99350 67410 99360 67480
rect 99140 67360 99360 67410
rect 99640 67590 99860 67640
rect 99640 67520 99650 67590
rect 99850 67520 99860 67590
rect 99640 67480 99860 67520
rect 99640 67410 99650 67480
rect 99850 67410 99860 67480
rect 99640 67360 99860 67410
rect -16000 67350 -12000 67360
rect -16000 67150 -15980 67350
rect -15910 67150 -15590 67350
rect -15520 67150 -15480 67350
rect -15410 67150 -15090 67350
rect -15020 67150 -14980 67350
rect -14910 67150 -14590 67350
rect -14520 67150 -14480 67350
rect -14410 67150 -14090 67350
rect -14020 67150 -13980 67350
rect -13910 67150 -13590 67350
rect -13520 67150 -13480 67350
rect -13410 67150 -13090 67350
rect -13020 67150 -12980 67350
rect -12910 67150 -12590 67350
rect -12520 67150 -12480 67350
rect -12410 67150 -12090 67350
rect -12020 67150 -12000 67350
rect -16000 67140 -12000 67150
rect 96000 67350 100000 67360
rect 96000 67150 96020 67350
rect 96090 67150 96410 67350
rect 96480 67150 96520 67350
rect 96590 67150 96910 67350
rect 96980 67150 97020 67350
rect 97090 67150 97410 67350
rect 97480 67150 97520 67350
rect 97590 67150 97910 67350
rect 97980 67150 98020 67350
rect 98090 67150 98410 67350
rect 98480 67150 98520 67350
rect 98590 67150 98910 67350
rect 98980 67150 99020 67350
rect 99090 67150 99410 67350
rect 99480 67150 99520 67350
rect 99590 67150 99910 67350
rect 99980 67150 100000 67350
rect 96000 67140 100000 67150
rect -15860 67090 -15640 67140
rect -15860 67020 -15850 67090
rect -15650 67020 -15640 67090
rect -15860 66980 -15640 67020
rect -15860 66910 -15850 66980
rect -15650 66910 -15640 66980
rect -15860 66860 -15640 66910
rect -15360 67090 -15140 67140
rect -15360 67020 -15350 67090
rect -15150 67020 -15140 67090
rect -15360 66980 -15140 67020
rect -15360 66910 -15350 66980
rect -15150 66910 -15140 66980
rect -15360 66860 -15140 66910
rect -14860 67090 -14640 67140
rect -14860 67020 -14850 67090
rect -14650 67020 -14640 67090
rect -14860 66980 -14640 67020
rect -14860 66910 -14850 66980
rect -14650 66910 -14640 66980
rect -14860 66860 -14640 66910
rect -14360 67090 -14140 67140
rect -14360 67020 -14350 67090
rect -14150 67020 -14140 67090
rect -14360 66980 -14140 67020
rect -14360 66910 -14350 66980
rect -14150 66910 -14140 66980
rect -14360 66860 -14140 66910
rect -13860 67090 -13640 67140
rect -13860 67020 -13850 67090
rect -13650 67020 -13640 67090
rect -13860 66980 -13640 67020
rect -13860 66910 -13850 66980
rect -13650 66910 -13640 66980
rect -13860 66860 -13640 66910
rect -13360 67090 -13140 67140
rect -13360 67020 -13350 67090
rect -13150 67020 -13140 67090
rect -13360 66980 -13140 67020
rect -13360 66910 -13350 66980
rect -13150 66910 -13140 66980
rect -13360 66860 -13140 66910
rect -12860 67090 -12640 67140
rect -12860 67020 -12850 67090
rect -12650 67020 -12640 67090
rect -12860 66980 -12640 67020
rect -12860 66910 -12850 66980
rect -12650 66910 -12640 66980
rect -12860 66860 -12640 66910
rect -12360 67090 -12140 67140
rect -12360 67020 -12350 67090
rect -12150 67020 -12140 67090
rect -12360 66980 -12140 67020
rect -12360 66910 -12350 66980
rect -12150 66910 -12140 66980
rect -12360 66860 -12140 66910
rect 96140 67090 96360 67140
rect 96140 67020 96150 67090
rect 96350 67020 96360 67090
rect 96140 66980 96360 67020
rect 96140 66910 96150 66980
rect 96350 66910 96360 66980
rect 96140 66860 96360 66910
rect 96640 67090 96860 67140
rect 96640 67020 96650 67090
rect 96850 67020 96860 67090
rect 96640 66980 96860 67020
rect 96640 66910 96650 66980
rect 96850 66910 96860 66980
rect 96640 66860 96860 66910
rect 97140 67090 97360 67140
rect 97140 67020 97150 67090
rect 97350 67020 97360 67090
rect 97140 66980 97360 67020
rect 97140 66910 97150 66980
rect 97350 66910 97360 66980
rect 97140 66860 97360 66910
rect 97640 67090 97860 67140
rect 97640 67020 97650 67090
rect 97850 67020 97860 67090
rect 97640 66980 97860 67020
rect 97640 66910 97650 66980
rect 97850 66910 97860 66980
rect 97640 66860 97860 66910
rect 98140 67090 98360 67140
rect 98140 67020 98150 67090
rect 98350 67020 98360 67090
rect 98140 66980 98360 67020
rect 98140 66910 98150 66980
rect 98350 66910 98360 66980
rect 98140 66860 98360 66910
rect 98640 67090 98860 67140
rect 98640 67020 98650 67090
rect 98850 67020 98860 67090
rect 98640 66980 98860 67020
rect 98640 66910 98650 66980
rect 98850 66910 98860 66980
rect 98640 66860 98860 66910
rect 99140 67090 99360 67140
rect 99140 67020 99150 67090
rect 99350 67020 99360 67090
rect 99140 66980 99360 67020
rect 99140 66910 99150 66980
rect 99350 66910 99360 66980
rect 99140 66860 99360 66910
rect 99640 67090 99860 67140
rect 99640 67020 99650 67090
rect 99850 67020 99860 67090
rect 99640 66980 99860 67020
rect 99640 66910 99650 66980
rect 99850 66910 99860 66980
rect 99640 66860 99860 66910
rect -16000 66850 -12000 66860
rect -16000 66650 -15980 66850
rect -15910 66650 -15590 66850
rect -15520 66650 -15480 66850
rect -15410 66650 -15090 66850
rect -15020 66650 -14980 66850
rect -14910 66650 -14590 66850
rect -14520 66650 -14480 66850
rect -14410 66650 -14090 66850
rect -14020 66650 -13980 66850
rect -13910 66650 -13590 66850
rect -13520 66650 -13480 66850
rect -13410 66650 -13090 66850
rect -13020 66650 -12980 66850
rect -12910 66650 -12590 66850
rect -12520 66650 -12480 66850
rect -12410 66650 -12090 66850
rect -12020 66650 -12000 66850
rect -16000 66640 -12000 66650
rect 96000 66850 100000 66860
rect 96000 66650 96020 66850
rect 96090 66650 96410 66850
rect 96480 66650 96520 66850
rect 96590 66650 96910 66850
rect 96980 66650 97020 66850
rect 97090 66650 97410 66850
rect 97480 66650 97520 66850
rect 97590 66650 97910 66850
rect 97980 66650 98020 66850
rect 98090 66650 98410 66850
rect 98480 66650 98520 66850
rect 98590 66650 98910 66850
rect 98980 66650 99020 66850
rect 99090 66650 99410 66850
rect 99480 66650 99520 66850
rect 99590 66650 99910 66850
rect 99980 66650 100000 66850
rect 96000 66640 100000 66650
rect -15860 66590 -15640 66640
rect -15860 66520 -15850 66590
rect -15650 66520 -15640 66590
rect -15860 66480 -15640 66520
rect -15860 66410 -15850 66480
rect -15650 66410 -15640 66480
rect -15860 66360 -15640 66410
rect -15360 66590 -15140 66640
rect -15360 66520 -15350 66590
rect -15150 66520 -15140 66590
rect -15360 66480 -15140 66520
rect -15360 66410 -15350 66480
rect -15150 66410 -15140 66480
rect -15360 66360 -15140 66410
rect -14860 66590 -14640 66640
rect -14860 66520 -14850 66590
rect -14650 66520 -14640 66590
rect -14860 66480 -14640 66520
rect -14860 66410 -14850 66480
rect -14650 66410 -14640 66480
rect -14860 66360 -14640 66410
rect -14360 66590 -14140 66640
rect -14360 66520 -14350 66590
rect -14150 66520 -14140 66590
rect -14360 66480 -14140 66520
rect -14360 66410 -14350 66480
rect -14150 66410 -14140 66480
rect -14360 66360 -14140 66410
rect -13860 66590 -13640 66640
rect -13860 66520 -13850 66590
rect -13650 66520 -13640 66590
rect -13860 66480 -13640 66520
rect -13860 66410 -13850 66480
rect -13650 66410 -13640 66480
rect -13860 66360 -13640 66410
rect -13360 66590 -13140 66640
rect -13360 66520 -13350 66590
rect -13150 66520 -13140 66590
rect -13360 66480 -13140 66520
rect -13360 66410 -13350 66480
rect -13150 66410 -13140 66480
rect -13360 66360 -13140 66410
rect -12860 66590 -12640 66640
rect -12860 66520 -12850 66590
rect -12650 66520 -12640 66590
rect -12860 66480 -12640 66520
rect -12860 66410 -12850 66480
rect -12650 66410 -12640 66480
rect -12860 66360 -12640 66410
rect -12360 66590 -12140 66640
rect -12360 66520 -12350 66590
rect -12150 66520 -12140 66590
rect -12360 66480 -12140 66520
rect -12360 66410 -12350 66480
rect -12150 66410 -12140 66480
rect -12360 66360 -12140 66410
rect 96140 66590 96360 66640
rect 96140 66520 96150 66590
rect 96350 66520 96360 66590
rect 96140 66480 96360 66520
rect 96140 66410 96150 66480
rect 96350 66410 96360 66480
rect 96140 66360 96360 66410
rect 96640 66590 96860 66640
rect 96640 66520 96650 66590
rect 96850 66520 96860 66590
rect 96640 66480 96860 66520
rect 96640 66410 96650 66480
rect 96850 66410 96860 66480
rect 96640 66360 96860 66410
rect 97140 66590 97360 66640
rect 97140 66520 97150 66590
rect 97350 66520 97360 66590
rect 97140 66480 97360 66520
rect 97140 66410 97150 66480
rect 97350 66410 97360 66480
rect 97140 66360 97360 66410
rect 97640 66590 97860 66640
rect 97640 66520 97650 66590
rect 97850 66520 97860 66590
rect 97640 66480 97860 66520
rect 97640 66410 97650 66480
rect 97850 66410 97860 66480
rect 97640 66360 97860 66410
rect 98140 66590 98360 66640
rect 98140 66520 98150 66590
rect 98350 66520 98360 66590
rect 98140 66480 98360 66520
rect 98140 66410 98150 66480
rect 98350 66410 98360 66480
rect 98140 66360 98360 66410
rect 98640 66590 98860 66640
rect 98640 66520 98650 66590
rect 98850 66520 98860 66590
rect 98640 66480 98860 66520
rect 98640 66410 98650 66480
rect 98850 66410 98860 66480
rect 98640 66360 98860 66410
rect 99140 66590 99360 66640
rect 99140 66520 99150 66590
rect 99350 66520 99360 66590
rect 99140 66480 99360 66520
rect 99140 66410 99150 66480
rect 99350 66410 99360 66480
rect 99140 66360 99360 66410
rect 99640 66590 99860 66640
rect 99640 66520 99650 66590
rect 99850 66520 99860 66590
rect 99640 66480 99860 66520
rect 99640 66410 99650 66480
rect 99850 66410 99860 66480
rect 99640 66360 99860 66410
rect -16000 66350 -12000 66360
rect -16000 66150 -15980 66350
rect -15910 66150 -15590 66350
rect -15520 66150 -15480 66350
rect -15410 66150 -15090 66350
rect -15020 66150 -14980 66350
rect -14910 66150 -14590 66350
rect -14520 66150 -14480 66350
rect -14410 66150 -14090 66350
rect -14020 66150 -13980 66350
rect -13910 66150 -13590 66350
rect -13520 66150 -13480 66350
rect -13410 66150 -13090 66350
rect -13020 66150 -12980 66350
rect -12910 66150 -12590 66350
rect -12520 66150 -12480 66350
rect -12410 66150 -12090 66350
rect -12020 66150 -12000 66350
rect -16000 66140 -12000 66150
rect 96000 66350 100000 66360
rect 96000 66150 96020 66350
rect 96090 66150 96410 66350
rect 96480 66150 96520 66350
rect 96590 66150 96910 66350
rect 96980 66150 97020 66350
rect 97090 66150 97410 66350
rect 97480 66150 97520 66350
rect 97590 66150 97910 66350
rect 97980 66150 98020 66350
rect 98090 66150 98410 66350
rect 98480 66150 98520 66350
rect 98590 66150 98910 66350
rect 98980 66150 99020 66350
rect 99090 66150 99410 66350
rect 99480 66150 99520 66350
rect 99590 66150 99910 66350
rect 99980 66150 100000 66350
rect 96000 66140 100000 66150
rect -15860 66090 -15640 66140
rect -15860 66020 -15850 66090
rect -15650 66020 -15640 66090
rect -15860 65980 -15640 66020
rect -15860 65910 -15850 65980
rect -15650 65910 -15640 65980
rect -15860 65860 -15640 65910
rect -15360 66090 -15140 66140
rect -15360 66020 -15350 66090
rect -15150 66020 -15140 66090
rect -15360 65980 -15140 66020
rect -15360 65910 -15350 65980
rect -15150 65910 -15140 65980
rect -15360 65860 -15140 65910
rect -14860 66090 -14640 66140
rect -14860 66020 -14850 66090
rect -14650 66020 -14640 66090
rect -14860 65980 -14640 66020
rect -14860 65910 -14850 65980
rect -14650 65910 -14640 65980
rect -14860 65860 -14640 65910
rect -14360 66090 -14140 66140
rect -14360 66020 -14350 66090
rect -14150 66020 -14140 66090
rect -14360 65980 -14140 66020
rect -14360 65910 -14350 65980
rect -14150 65910 -14140 65980
rect -14360 65860 -14140 65910
rect -13860 66090 -13640 66140
rect -13860 66020 -13850 66090
rect -13650 66020 -13640 66090
rect -13860 65980 -13640 66020
rect -13860 65910 -13850 65980
rect -13650 65910 -13640 65980
rect -13860 65860 -13640 65910
rect -13360 66090 -13140 66140
rect -13360 66020 -13350 66090
rect -13150 66020 -13140 66090
rect -13360 65980 -13140 66020
rect -13360 65910 -13350 65980
rect -13150 65910 -13140 65980
rect -13360 65860 -13140 65910
rect -12860 66090 -12640 66140
rect -12860 66020 -12850 66090
rect -12650 66020 -12640 66090
rect -12860 65980 -12640 66020
rect -12860 65910 -12850 65980
rect -12650 65910 -12640 65980
rect -12860 65860 -12640 65910
rect -12360 66090 -12140 66140
rect -12360 66020 -12350 66090
rect -12150 66020 -12140 66090
rect -12360 65980 -12140 66020
rect -12360 65910 -12350 65980
rect -12150 65910 -12140 65980
rect -12360 65860 -12140 65910
rect 96140 66090 96360 66140
rect 96140 66020 96150 66090
rect 96350 66020 96360 66090
rect 96140 65980 96360 66020
rect 96140 65910 96150 65980
rect 96350 65910 96360 65980
rect 96140 65860 96360 65910
rect 96640 66090 96860 66140
rect 96640 66020 96650 66090
rect 96850 66020 96860 66090
rect 96640 65980 96860 66020
rect 96640 65910 96650 65980
rect 96850 65910 96860 65980
rect 96640 65860 96860 65910
rect 97140 66090 97360 66140
rect 97140 66020 97150 66090
rect 97350 66020 97360 66090
rect 97140 65980 97360 66020
rect 97140 65910 97150 65980
rect 97350 65910 97360 65980
rect 97140 65860 97360 65910
rect 97640 66090 97860 66140
rect 97640 66020 97650 66090
rect 97850 66020 97860 66090
rect 97640 65980 97860 66020
rect 97640 65910 97650 65980
rect 97850 65910 97860 65980
rect 97640 65860 97860 65910
rect 98140 66090 98360 66140
rect 98140 66020 98150 66090
rect 98350 66020 98360 66090
rect 98140 65980 98360 66020
rect 98140 65910 98150 65980
rect 98350 65910 98360 65980
rect 98140 65860 98360 65910
rect 98640 66090 98860 66140
rect 98640 66020 98650 66090
rect 98850 66020 98860 66090
rect 98640 65980 98860 66020
rect 98640 65910 98650 65980
rect 98850 65910 98860 65980
rect 98640 65860 98860 65910
rect 99140 66090 99360 66140
rect 99140 66020 99150 66090
rect 99350 66020 99360 66090
rect 99140 65980 99360 66020
rect 99140 65910 99150 65980
rect 99350 65910 99360 65980
rect 99140 65860 99360 65910
rect 99640 66090 99860 66140
rect 99640 66020 99650 66090
rect 99850 66020 99860 66090
rect 99640 65980 99860 66020
rect 99640 65910 99650 65980
rect 99850 65910 99860 65980
rect 99640 65860 99860 65910
rect -16000 65850 -12000 65860
rect -16000 65650 -15980 65850
rect -15910 65650 -15590 65850
rect -15520 65650 -15480 65850
rect -15410 65650 -15090 65850
rect -15020 65650 -14980 65850
rect -14910 65650 -14590 65850
rect -14520 65650 -14480 65850
rect -14410 65650 -14090 65850
rect -14020 65650 -13980 65850
rect -13910 65650 -13590 65850
rect -13520 65650 -13480 65850
rect -13410 65650 -13090 65850
rect -13020 65650 -12980 65850
rect -12910 65650 -12590 65850
rect -12520 65650 -12480 65850
rect -12410 65650 -12090 65850
rect -12020 65650 -12000 65850
rect -16000 65640 -12000 65650
rect 96000 65850 100000 65860
rect 96000 65650 96020 65850
rect 96090 65650 96410 65850
rect 96480 65650 96520 65850
rect 96590 65650 96910 65850
rect 96980 65650 97020 65850
rect 97090 65650 97410 65850
rect 97480 65650 97520 65850
rect 97590 65650 97910 65850
rect 97980 65650 98020 65850
rect 98090 65650 98410 65850
rect 98480 65650 98520 65850
rect 98590 65650 98910 65850
rect 98980 65650 99020 65850
rect 99090 65650 99410 65850
rect 99480 65650 99520 65850
rect 99590 65650 99910 65850
rect 99980 65650 100000 65850
rect 96000 65640 100000 65650
rect -15860 65590 -15640 65640
rect -15860 65520 -15850 65590
rect -15650 65520 -15640 65590
rect -15860 65480 -15640 65520
rect -15860 65410 -15850 65480
rect -15650 65410 -15640 65480
rect -15860 65360 -15640 65410
rect -15360 65590 -15140 65640
rect -15360 65520 -15350 65590
rect -15150 65520 -15140 65590
rect -15360 65480 -15140 65520
rect -15360 65410 -15350 65480
rect -15150 65410 -15140 65480
rect -15360 65360 -15140 65410
rect -14860 65590 -14640 65640
rect -14860 65520 -14850 65590
rect -14650 65520 -14640 65590
rect -14860 65480 -14640 65520
rect -14860 65410 -14850 65480
rect -14650 65410 -14640 65480
rect -14860 65360 -14640 65410
rect -14360 65590 -14140 65640
rect -14360 65520 -14350 65590
rect -14150 65520 -14140 65590
rect -14360 65480 -14140 65520
rect -14360 65410 -14350 65480
rect -14150 65410 -14140 65480
rect -14360 65360 -14140 65410
rect -13860 65590 -13640 65640
rect -13860 65520 -13850 65590
rect -13650 65520 -13640 65590
rect -13860 65480 -13640 65520
rect -13860 65410 -13850 65480
rect -13650 65410 -13640 65480
rect -13860 65360 -13640 65410
rect -13360 65590 -13140 65640
rect -13360 65520 -13350 65590
rect -13150 65520 -13140 65590
rect -13360 65480 -13140 65520
rect -13360 65410 -13350 65480
rect -13150 65410 -13140 65480
rect -13360 65360 -13140 65410
rect -12860 65590 -12640 65640
rect -12860 65520 -12850 65590
rect -12650 65520 -12640 65590
rect -12860 65480 -12640 65520
rect -12860 65410 -12850 65480
rect -12650 65410 -12640 65480
rect -12860 65360 -12640 65410
rect -12360 65590 -12140 65640
rect -12360 65520 -12350 65590
rect -12150 65520 -12140 65590
rect -12360 65480 -12140 65520
rect -12360 65410 -12350 65480
rect -12150 65410 -12140 65480
rect -12360 65360 -12140 65410
rect 96140 65590 96360 65640
rect 96140 65520 96150 65590
rect 96350 65520 96360 65590
rect 96140 65480 96360 65520
rect 96140 65410 96150 65480
rect 96350 65410 96360 65480
rect 96140 65360 96360 65410
rect 96640 65590 96860 65640
rect 96640 65520 96650 65590
rect 96850 65520 96860 65590
rect 96640 65480 96860 65520
rect 96640 65410 96650 65480
rect 96850 65410 96860 65480
rect 96640 65360 96860 65410
rect 97140 65590 97360 65640
rect 97140 65520 97150 65590
rect 97350 65520 97360 65590
rect 97140 65480 97360 65520
rect 97140 65410 97150 65480
rect 97350 65410 97360 65480
rect 97140 65360 97360 65410
rect 97640 65590 97860 65640
rect 97640 65520 97650 65590
rect 97850 65520 97860 65590
rect 97640 65480 97860 65520
rect 97640 65410 97650 65480
rect 97850 65410 97860 65480
rect 97640 65360 97860 65410
rect 98140 65590 98360 65640
rect 98140 65520 98150 65590
rect 98350 65520 98360 65590
rect 98140 65480 98360 65520
rect 98140 65410 98150 65480
rect 98350 65410 98360 65480
rect 98140 65360 98360 65410
rect 98640 65590 98860 65640
rect 98640 65520 98650 65590
rect 98850 65520 98860 65590
rect 98640 65480 98860 65520
rect 98640 65410 98650 65480
rect 98850 65410 98860 65480
rect 98640 65360 98860 65410
rect 99140 65590 99360 65640
rect 99140 65520 99150 65590
rect 99350 65520 99360 65590
rect 99140 65480 99360 65520
rect 99140 65410 99150 65480
rect 99350 65410 99360 65480
rect 99140 65360 99360 65410
rect 99640 65590 99860 65640
rect 99640 65520 99650 65590
rect 99850 65520 99860 65590
rect 99640 65480 99860 65520
rect 99640 65410 99650 65480
rect 99850 65410 99860 65480
rect 99640 65360 99860 65410
rect -16000 65350 -12000 65360
rect -16000 65150 -15980 65350
rect -15910 65150 -15590 65350
rect -15520 65150 -15480 65350
rect -15410 65150 -15090 65350
rect -15020 65150 -14980 65350
rect -14910 65150 -14590 65350
rect -14520 65150 -14480 65350
rect -14410 65150 -14090 65350
rect -14020 65150 -13980 65350
rect -13910 65150 -13590 65350
rect -13520 65150 -13480 65350
rect -13410 65150 -13090 65350
rect -13020 65150 -12980 65350
rect -12910 65150 -12590 65350
rect -12520 65150 -12480 65350
rect -12410 65150 -12090 65350
rect -12020 65150 -12000 65350
rect -16000 65140 -12000 65150
rect 96000 65350 100000 65360
rect 96000 65150 96020 65350
rect 96090 65150 96410 65350
rect 96480 65150 96520 65350
rect 96590 65150 96910 65350
rect 96980 65150 97020 65350
rect 97090 65150 97410 65350
rect 97480 65150 97520 65350
rect 97590 65150 97910 65350
rect 97980 65150 98020 65350
rect 98090 65150 98410 65350
rect 98480 65150 98520 65350
rect 98590 65150 98910 65350
rect 98980 65150 99020 65350
rect 99090 65150 99410 65350
rect 99480 65150 99520 65350
rect 99590 65150 99910 65350
rect 99980 65150 100000 65350
rect 96000 65140 100000 65150
rect -15860 65090 -15640 65140
rect -15860 65020 -15850 65090
rect -15650 65020 -15640 65090
rect -15860 64980 -15640 65020
rect -15860 64910 -15850 64980
rect -15650 64910 -15640 64980
rect -15860 64860 -15640 64910
rect -15360 65090 -15140 65140
rect -15360 65020 -15350 65090
rect -15150 65020 -15140 65090
rect -15360 64980 -15140 65020
rect -15360 64910 -15350 64980
rect -15150 64910 -15140 64980
rect -15360 64860 -15140 64910
rect -14860 65090 -14640 65140
rect -14860 65020 -14850 65090
rect -14650 65020 -14640 65090
rect -14860 64980 -14640 65020
rect -14860 64910 -14850 64980
rect -14650 64910 -14640 64980
rect -14860 64860 -14640 64910
rect -14360 65090 -14140 65140
rect -14360 65020 -14350 65090
rect -14150 65020 -14140 65090
rect -14360 64980 -14140 65020
rect -14360 64910 -14350 64980
rect -14150 64910 -14140 64980
rect -14360 64860 -14140 64910
rect -13860 65090 -13640 65140
rect -13860 65020 -13850 65090
rect -13650 65020 -13640 65090
rect -13860 64980 -13640 65020
rect -13860 64910 -13850 64980
rect -13650 64910 -13640 64980
rect -13860 64860 -13640 64910
rect -13360 65090 -13140 65140
rect -13360 65020 -13350 65090
rect -13150 65020 -13140 65090
rect -13360 64980 -13140 65020
rect -13360 64910 -13350 64980
rect -13150 64910 -13140 64980
rect -13360 64860 -13140 64910
rect -12860 65090 -12640 65140
rect -12860 65020 -12850 65090
rect -12650 65020 -12640 65090
rect -12860 64980 -12640 65020
rect -12860 64910 -12850 64980
rect -12650 64910 -12640 64980
rect -12860 64860 -12640 64910
rect -12360 65090 -12140 65140
rect -12360 65020 -12350 65090
rect -12150 65020 -12140 65090
rect -12360 64980 -12140 65020
rect -12360 64910 -12350 64980
rect -12150 64910 -12140 64980
rect -12360 64860 -12140 64910
rect 96140 65090 96360 65140
rect 96140 65020 96150 65090
rect 96350 65020 96360 65090
rect 96140 64980 96360 65020
rect 96140 64910 96150 64980
rect 96350 64910 96360 64980
rect 96140 64860 96360 64910
rect 96640 65090 96860 65140
rect 96640 65020 96650 65090
rect 96850 65020 96860 65090
rect 96640 64980 96860 65020
rect 96640 64910 96650 64980
rect 96850 64910 96860 64980
rect 96640 64860 96860 64910
rect 97140 65090 97360 65140
rect 97140 65020 97150 65090
rect 97350 65020 97360 65090
rect 97140 64980 97360 65020
rect 97140 64910 97150 64980
rect 97350 64910 97360 64980
rect 97140 64860 97360 64910
rect 97640 65090 97860 65140
rect 97640 65020 97650 65090
rect 97850 65020 97860 65090
rect 97640 64980 97860 65020
rect 97640 64910 97650 64980
rect 97850 64910 97860 64980
rect 97640 64860 97860 64910
rect 98140 65090 98360 65140
rect 98140 65020 98150 65090
rect 98350 65020 98360 65090
rect 98140 64980 98360 65020
rect 98140 64910 98150 64980
rect 98350 64910 98360 64980
rect 98140 64860 98360 64910
rect 98640 65090 98860 65140
rect 98640 65020 98650 65090
rect 98850 65020 98860 65090
rect 98640 64980 98860 65020
rect 98640 64910 98650 64980
rect 98850 64910 98860 64980
rect 98640 64860 98860 64910
rect 99140 65090 99360 65140
rect 99140 65020 99150 65090
rect 99350 65020 99360 65090
rect 99140 64980 99360 65020
rect 99140 64910 99150 64980
rect 99350 64910 99360 64980
rect 99140 64860 99360 64910
rect 99640 65090 99860 65140
rect 99640 65020 99650 65090
rect 99850 65020 99860 65090
rect 99640 64980 99860 65020
rect 99640 64910 99650 64980
rect 99850 64910 99860 64980
rect 99640 64860 99860 64910
rect -16000 64850 -12000 64860
rect -16000 64650 -15980 64850
rect -15910 64650 -15590 64850
rect -15520 64650 -15480 64850
rect -15410 64650 -15090 64850
rect -15020 64650 -14980 64850
rect -14910 64650 -14590 64850
rect -14520 64650 -14480 64850
rect -14410 64650 -14090 64850
rect -14020 64650 -13980 64850
rect -13910 64650 -13590 64850
rect -13520 64650 -13480 64850
rect -13410 64650 -13090 64850
rect -13020 64650 -12980 64850
rect -12910 64650 -12590 64850
rect -12520 64650 -12480 64850
rect -12410 64650 -12090 64850
rect -12020 64650 -12000 64850
rect -16000 64640 -12000 64650
rect 96000 64850 100000 64860
rect 96000 64650 96020 64850
rect 96090 64650 96410 64850
rect 96480 64650 96520 64850
rect 96590 64650 96910 64850
rect 96980 64650 97020 64850
rect 97090 64650 97410 64850
rect 97480 64650 97520 64850
rect 97590 64650 97910 64850
rect 97980 64650 98020 64850
rect 98090 64650 98410 64850
rect 98480 64650 98520 64850
rect 98590 64650 98910 64850
rect 98980 64650 99020 64850
rect 99090 64650 99410 64850
rect 99480 64650 99520 64850
rect 99590 64650 99910 64850
rect 99980 64650 100000 64850
rect 96000 64640 100000 64650
rect -15860 64590 -15640 64640
rect -15860 64520 -15850 64590
rect -15650 64520 -15640 64590
rect -15860 64480 -15640 64520
rect -15860 64410 -15850 64480
rect -15650 64410 -15640 64480
rect -15860 64360 -15640 64410
rect -15360 64590 -15140 64640
rect -15360 64520 -15350 64590
rect -15150 64520 -15140 64590
rect -15360 64480 -15140 64520
rect -15360 64410 -15350 64480
rect -15150 64410 -15140 64480
rect -15360 64360 -15140 64410
rect -14860 64590 -14640 64640
rect -14860 64520 -14850 64590
rect -14650 64520 -14640 64590
rect -14860 64480 -14640 64520
rect -14860 64410 -14850 64480
rect -14650 64410 -14640 64480
rect -14860 64360 -14640 64410
rect -14360 64590 -14140 64640
rect -14360 64520 -14350 64590
rect -14150 64520 -14140 64590
rect -14360 64480 -14140 64520
rect -14360 64410 -14350 64480
rect -14150 64410 -14140 64480
rect -14360 64360 -14140 64410
rect -13860 64590 -13640 64640
rect -13860 64520 -13850 64590
rect -13650 64520 -13640 64590
rect -13860 64480 -13640 64520
rect -13860 64410 -13850 64480
rect -13650 64410 -13640 64480
rect -13860 64360 -13640 64410
rect -13360 64590 -13140 64640
rect -13360 64520 -13350 64590
rect -13150 64520 -13140 64590
rect -13360 64480 -13140 64520
rect -13360 64410 -13350 64480
rect -13150 64410 -13140 64480
rect -13360 64360 -13140 64410
rect -12860 64590 -12640 64640
rect -12860 64520 -12850 64590
rect -12650 64520 -12640 64590
rect -12860 64480 -12640 64520
rect -12860 64410 -12850 64480
rect -12650 64410 -12640 64480
rect -12860 64360 -12640 64410
rect -12360 64590 -12140 64640
rect -12360 64520 -12350 64590
rect -12150 64520 -12140 64590
rect -12360 64480 -12140 64520
rect -12360 64410 -12350 64480
rect -12150 64410 -12140 64480
rect -12360 64360 -12140 64410
rect 96140 64590 96360 64640
rect 96140 64520 96150 64590
rect 96350 64520 96360 64590
rect 96140 64480 96360 64520
rect 96140 64410 96150 64480
rect 96350 64410 96360 64480
rect 96140 64360 96360 64410
rect 96640 64590 96860 64640
rect 96640 64520 96650 64590
rect 96850 64520 96860 64590
rect 96640 64480 96860 64520
rect 96640 64410 96650 64480
rect 96850 64410 96860 64480
rect 96640 64360 96860 64410
rect 97140 64590 97360 64640
rect 97140 64520 97150 64590
rect 97350 64520 97360 64590
rect 97140 64480 97360 64520
rect 97140 64410 97150 64480
rect 97350 64410 97360 64480
rect 97140 64360 97360 64410
rect 97640 64590 97860 64640
rect 97640 64520 97650 64590
rect 97850 64520 97860 64590
rect 97640 64480 97860 64520
rect 97640 64410 97650 64480
rect 97850 64410 97860 64480
rect 97640 64360 97860 64410
rect 98140 64590 98360 64640
rect 98140 64520 98150 64590
rect 98350 64520 98360 64590
rect 98140 64480 98360 64520
rect 98140 64410 98150 64480
rect 98350 64410 98360 64480
rect 98140 64360 98360 64410
rect 98640 64590 98860 64640
rect 98640 64520 98650 64590
rect 98850 64520 98860 64590
rect 98640 64480 98860 64520
rect 98640 64410 98650 64480
rect 98850 64410 98860 64480
rect 98640 64360 98860 64410
rect 99140 64590 99360 64640
rect 99140 64520 99150 64590
rect 99350 64520 99360 64590
rect 99140 64480 99360 64520
rect 99140 64410 99150 64480
rect 99350 64410 99360 64480
rect 99140 64360 99360 64410
rect 99640 64590 99860 64640
rect 99640 64520 99650 64590
rect 99850 64520 99860 64590
rect 99640 64480 99860 64520
rect 99640 64410 99650 64480
rect 99850 64410 99860 64480
rect 99640 64360 99860 64410
rect -16000 64350 -12000 64360
rect -16000 64150 -15980 64350
rect -15910 64150 -15590 64350
rect -15520 64150 -15480 64350
rect -15410 64150 -15090 64350
rect -15020 64150 -14980 64350
rect -14910 64150 -14590 64350
rect -14520 64150 -14480 64350
rect -14410 64150 -14090 64350
rect -14020 64150 -13980 64350
rect -13910 64150 -13590 64350
rect -13520 64150 -13480 64350
rect -13410 64150 -13090 64350
rect -13020 64150 -12980 64350
rect -12910 64150 -12590 64350
rect -12520 64150 -12480 64350
rect -12410 64150 -12090 64350
rect -12020 64150 -12000 64350
rect -16000 64140 -12000 64150
rect 96000 64350 100000 64360
rect 96000 64150 96020 64350
rect 96090 64150 96410 64350
rect 96480 64150 96520 64350
rect 96590 64150 96910 64350
rect 96980 64150 97020 64350
rect 97090 64150 97410 64350
rect 97480 64150 97520 64350
rect 97590 64150 97910 64350
rect 97980 64150 98020 64350
rect 98090 64150 98410 64350
rect 98480 64150 98520 64350
rect 98590 64150 98910 64350
rect 98980 64150 99020 64350
rect 99090 64150 99410 64350
rect 99480 64150 99520 64350
rect 99590 64150 99910 64350
rect 99980 64150 100000 64350
rect 96000 64140 100000 64150
rect -15860 64090 -15640 64140
rect -15860 64020 -15850 64090
rect -15650 64020 -15640 64090
rect -15860 63980 -15640 64020
rect -15860 63910 -15850 63980
rect -15650 63910 -15640 63980
rect -15860 63860 -15640 63910
rect -15360 64090 -15140 64140
rect -15360 64020 -15350 64090
rect -15150 64020 -15140 64090
rect -15360 63980 -15140 64020
rect -15360 63910 -15350 63980
rect -15150 63910 -15140 63980
rect -15360 63860 -15140 63910
rect -14860 64090 -14640 64140
rect -14860 64020 -14850 64090
rect -14650 64020 -14640 64090
rect -14860 63980 -14640 64020
rect -14860 63910 -14850 63980
rect -14650 63910 -14640 63980
rect -14860 63860 -14640 63910
rect -14360 64090 -14140 64140
rect -14360 64020 -14350 64090
rect -14150 64020 -14140 64090
rect -14360 63980 -14140 64020
rect -14360 63910 -14350 63980
rect -14150 63910 -14140 63980
rect -14360 63860 -14140 63910
rect -13860 64090 -13640 64140
rect -13860 64020 -13850 64090
rect -13650 64020 -13640 64090
rect -13860 63980 -13640 64020
rect -13860 63910 -13850 63980
rect -13650 63910 -13640 63980
rect -13860 63860 -13640 63910
rect -13360 64090 -13140 64140
rect -13360 64020 -13350 64090
rect -13150 64020 -13140 64090
rect -13360 63980 -13140 64020
rect -13360 63910 -13350 63980
rect -13150 63910 -13140 63980
rect -13360 63860 -13140 63910
rect -12860 64090 -12640 64140
rect -12860 64020 -12850 64090
rect -12650 64020 -12640 64090
rect -12860 63980 -12640 64020
rect -12860 63910 -12850 63980
rect -12650 63910 -12640 63980
rect -12860 63860 -12640 63910
rect -12360 64090 -12140 64140
rect -12360 64020 -12350 64090
rect -12150 64020 -12140 64090
rect -12360 63980 -12140 64020
rect -12360 63910 -12350 63980
rect -12150 63910 -12140 63980
rect -12360 63860 -12140 63910
rect 96140 64090 96360 64140
rect 96140 64020 96150 64090
rect 96350 64020 96360 64090
rect 96140 63980 96360 64020
rect 96140 63910 96150 63980
rect 96350 63910 96360 63980
rect 96140 63860 96360 63910
rect 96640 64090 96860 64140
rect 96640 64020 96650 64090
rect 96850 64020 96860 64090
rect 96640 63980 96860 64020
rect 96640 63910 96650 63980
rect 96850 63910 96860 63980
rect 96640 63860 96860 63910
rect 97140 64090 97360 64140
rect 97140 64020 97150 64090
rect 97350 64020 97360 64090
rect 97140 63980 97360 64020
rect 97140 63910 97150 63980
rect 97350 63910 97360 63980
rect 97140 63860 97360 63910
rect 97640 64090 97860 64140
rect 97640 64020 97650 64090
rect 97850 64020 97860 64090
rect 97640 63980 97860 64020
rect 97640 63910 97650 63980
rect 97850 63910 97860 63980
rect 97640 63860 97860 63910
rect 98140 64090 98360 64140
rect 98140 64020 98150 64090
rect 98350 64020 98360 64090
rect 98140 63980 98360 64020
rect 98140 63910 98150 63980
rect 98350 63910 98360 63980
rect 98140 63860 98360 63910
rect 98640 64090 98860 64140
rect 98640 64020 98650 64090
rect 98850 64020 98860 64090
rect 98640 63980 98860 64020
rect 98640 63910 98650 63980
rect 98850 63910 98860 63980
rect 98640 63860 98860 63910
rect 99140 64090 99360 64140
rect 99140 64020 99150 64090
rect 99350 64020 99360 64090
rect 99140 63980 99360 64020
rect 99140 63910 99150 63980
rect 99350 63910 99360 63980
rect 99140 63860 99360 63910
rect 99640 64090 99860 64140
rect 99640 64020 99650 64090
rect 99850 64020 99860 64090
rect 99640 63980 99860 64020
rect 99640 63910 99650 63980
rect 99850 63910 99860 63980
rect 99640 63860 99860 63910
rect -16000 63850 -12000 63860
rect -16000 63650 -15980 63850
rect -15910 63650 -15590 63850
rect -15520 63650 -15480 63850
rect -15410 63650 -15090 63850
rect -15020 63650 -14980 63850
rect -14910 63650 -14590 63850
rect -14520 63650 -14480 63850
rect -14410 63650 -14090 63850
rect -14020 63650 -13980 63850
rect -13910 63650 -13590 63850
rect -13520 63650 -13480 63850
rect -13410 63650 -13090 63850
rect -13020 63650 -12980 63850
rect -12910 63650 -12590 63850
rect -12520 63650 -12480 63850
rect -12410 63650 -12090 63850
rect -12020 63650 -12000 63850
rect -16000 63640 -12000 63650
rect 96000 63850 100000 63860
rect 96000 63650 96020 63850
rect 96090 63650 96410 63850
rect 96480 63650 96520 63850
rect 96590 63650 96910 63850
rect 96980 63650 97020 63850
rect 97090 63650 97410 63850
rect 97480 63650 97520 63850
rect 97590 63650 97910 63850
rect 97980 63650 98020 63850
rect 98090 63650 98410 63850
rect 98480 63650 98520 63850
rect 98590 63650 98910 63850
rect 98980 63650 99020 63850
rect 99090 63650 99410 63850
rect 99480 63650 99520 63850
rect 99590 63650 99910 63850
rect 99980 63650 100000 63850
rect 96000 63640 100000 63650
rect -15860 63590 -15640 63640
rect -15860 63520 -15850 63590
rect -15650 63520 -15640 63590
rect -15860 63480 -15640 63520
rect -15860 63410 -15850 63480
rect -15650 63410 -15640 63480
rect -15860 63360 -15640 63410
rect -15360 63590 -15140 63640
rect -15360 63520 -15350 63590
rect -15150 63520 -15140 63590
rect -15360 63480 -15140 63520
rect -15360 63410 -15350 63480
rect -15150 63410 -15140 63480
rect -15360 63360 -15140 63410
rect -14860 63590 -14640 63640
rect -14860 63520 -14850 63590
rect -14650 63520 -14640 63590
rect -14860 63480 -14640 63520
rect -14860 63410 -14850 63480
rect -14650 63410 -14640 63480
rect -14860 63360 -14640 63410
rect -14360 63590 -14140 63640
rect -14360 63520 -14350 63590
rect -14150 63520 -14140 63590
rect -14360 63480 -14140 63520
rect -14360 63410 -14350 63480
rect -14150 63410 -14140 63480
rect -14360 63360 -14140 63410
rect -13860 63590 -13640 63640
rect -13860 63520 -13850 63590
rect -13650 63520 -13640 63590
rect -13860 63480 -13640 63520
rect -13860 63410 -13850 63480
rect -13650 63410 -13640 63480
rect -13860 63360 -13640 63410
rect -13360 63590 -13140 63640
rect -13360 63520 -13350 63590
rect -13150 63520 -13140 63590
rect -13360 63480 -13140 63520
rect -13360 63410 -13350 63480
rect -13150 63410 -13140 63480
rect -13360 63360 -13140 63410
rect -12860 63590 -12640 63640
rect -12860 63520 -12850 63590
rect -12650 63520 -12640 63590
rect -12860 63480 -12640 63520
rect -12860 63410 -12850 63480
rect -12650 63410 -12640 63480
rect -12860 63360 -12640 63410
rect -12360 63590 -12140 63640
rect -12360 63520 -12350 63590
rect -12150 63520 -12140 63590
rect -12360 63480 -12140 63520
rect -12360 63410 -12350 63480
rect -12150 63410 -12140 63480
rect -12360 63360 -12140 63410
rect 96140 63590 96360 63640
rect 96140 63520 96150 63590
rect 96350 63520 96360 63590
rect 96140 63480 96360 63520
rect 96140 63410 96150 63480
rect 96350 63410 96360 63480
rect 96140 63360 96360 63410
rect 96640 63590 96860 63640
rect 96640 63520 96650 63590
rect 96850 63520 96860 63590
rect 96640 63480 96860 63520
rect 96640 63410 96650 63480
rect 96850 63410 96860 63480
rect 96640 63360 96860 63410
rect 97140 63590 97360 63640
rect 97140 63520 97150 63590
rect 97350 63520 97360 63590
rect 97140 63480 97360 63520
rect 97140 63410 97150 63480
rect 97350 63410 97360 63480
rect 97140 63360 97360 63410
rect 97640 63590 97860 63640
rect 97640 63520 97650 63590
rect 97850 63520 97860 63590
rect 97640 63480 97860 63520
rect 97640 63410 97650 63480
rect 97850 63410 97860 63480
rect 97640 63360 97860 63410
rect 98140 63590 98360 63640
rect 98140 63520 98150 63590
rect 98350 63520 98360 63590
rect 98140 63480 98360 63520
rect 98140 63410 98150 63480
rect 98350 63410 98360 63480
rect 98140 63360 98360 63410
rect 98640 63590 98860 63640
rect 98640 63520 98650 63590
rect 98850 63520 98860 63590
rect 98640 63480 98860 63520
rect 98640 63410 98650 63480
rect 98850 63410 98860 63480
rect 98640 63360 98860 63410
rect 99140 63590 99360 63640
rect 99140 63520 99150 63590
rect 99350 63520 99360 63590
rect 99140 63480 99360 63520
rect 99140 63410 99150 63480
rect 99350 63410 99360 63480
rect 99140 63360 99360 63410
rect 99640 63590 99860 63640
rect 99640 63520 99650 63590
rect 99850 63520 99860 63590
rect 99640 63480 99860 63520
rect 99640 63410 99650 63480
rect 99850 63410 99860 63480
rect 99640 63360 99860 63410
rect -16000 63350 -12000 63360
rect -16000 63150 -15980 63350
rect -15910 63150 -15590 63350
rect -15520 63150 -15480 63350
rect -15410 63150 -15090 63350
rect -15020 63150 -14980 63350
rect -14910 63150 -14590 63350
rect -14520 63150 -14480 63350
rect -14410 63150 -14090 63350
rect -14020 63150 -13980 63350
rect -13910 63150 -13590 63350
rect -13520 63150 -13480 63350
rect -13410 63150 -13090 63350
rect -13020 63150 -12980 63350
rect -12910 63150 -12590 63350
rect -12520 63150 -12480 63350
rect -12410 63150 -12090 63350
rect -12020 63150 -12000 63350
rect -16000 63140 -12000 63150
rect 96000 63350 100000 63360
rect 96000 63150 96020 63350
rect 96090 63150 96410 63350
rect 96480 63150 96520 63350
rect 96590 63150 96910 63350
rect 96980 63150 97020 63350
rect 97090 63150 97410 63350
rect 97480 63150 97520 63350
rect 97590 63150 97910 63350
rect 97980 63150 98020 63350
rect 98090 63150 98410 63350
rect 98480 63150 98520 63350
rect 98590 63150 98910 63350
rect 98980 63150 99020 63350
rect 99090 63150 99410 63350
rect 99480 63150 99520 63350
rect 99590 63150 99910 63350
rect 99980 63150 100000 63350
rect 96000 63140 100000 63150
rect -15860 63090 -15640 63140
rect -15860 63020 -15850 63090
rect -15650 63020 -15640 63090
rect -15860 62980 -15640 63020
rect -15860 62910 -15850 62980
rect -15650 62910 -15640 62980
rect -15860 62860 -15640 62910
rect -15360 63090 -15140 63140
rect -15360 63020 -15350 63090
rect -15150 63020 -15140 63090
rect -15360 62980 -15140 63020
rect -15360 62910 -15350 62980
rect -15150 62910 -15140 62980
rect -15360 62860 -15140 62910
rect -14860 63090 -14640 63140
rect -14860 63020 -14850 63090
rect -14650 63020 -14640 63090
rect -14860 62980 -14640 63020
rect -14860 62910 -14850 62980
rect -14650 62910 -14640 62980
rect -14860 62860 -14640 62910
rect -14360 63090 -14140 63140
rect -14360 63020 -14350 63090
rect -14150 63020 -14140 63090
rect -14360 62980 -14140 63020
rect -14360 62910 -14350 62980
rect -14150 62910 -14140 62980
rect -14360 62860 -14140 62910
rect -13860 63090 -13640 63140
rect -13860 63020 -13850 63090
rect -13650 63020 -13640 63090
rect -13860 62980 -13640 63020
rect -13860 62910 -13850 62980
rect -13650 62910 -13640 62980
rect -13860 62860 -13640 62910
rect -13360 63090 -13140 63140
rect -13360 63020 -13350 63090
rect -13150 63020 -13140 63090
rect -13360 62980 -13140 63020
rect -13360 62910 -13350 62980
rect -13150 62910 -13140 62980
rect -13360 62860 -13140 62910
rect -12860 63090 -12640 63140
rect -12860 63020 -12850 63090
rect -12650 63020 -12640 63090
rect -12860 62980 -12640 63020
rect -12860 62910 -12850 62980
rect -12650 62910 -12640 62980
rect -12860 62860 -12640 62910
rect -12360 63090 -12140 63140
rect -12360 63020 -12350 63090
rect -12150 63020 -12140 63090
rect -12360 62980 -12140 63020
rect -12360 62910 -12350 62980
rect -12150 62910 -12140 62980
rect -12360 62860 -12140 62910
rect 96140 63090 96360 63140
rect 96140 63020 96150 63090
rect 96350 63020 96360 63090
rect 96140 62980 96360 63020
rect 96140 62910 96150 62980
rect 96350 62910 96360 62980
rect 96140 62860 96360 62910
rect 96640 63090 96860 63140
rect 96640 63020 96650 63090
rect 96850 63020 96860 63090
rect 96640 62980 96860 63020
rect 96640 62910 96650 62980
rect 96850 62910 96860 62980
rect 96640 62860 96860 62910
rect 97140 63090 97360 63140
rect 97140 63020 97150 63090
rect 97350 63020 97360 63090
rect 97140 62980 97360 63020
rect 97140 62910 97150 62980
rect 97350 62910 97360 62980
rect 97140 62860 97360 62910
rect 97640 63090 97860 63140
rect 97640 63020 97650 63090
rect 97850 63020 97860 63090
rect 97640 62980 97860 63020
rect 97640 62910 97650 62980
rect 97850 62910 97860 62980
rect 97640 62860 97860 62910
rect 98140 63090 98360 63140
rect 98140 63020 98150 63090
rect 98350 63020 98360 63090
rect 98140 62980 98360 63020
rect 98140 62910 98150 62980
rect 98350 62910 98360 62980
rect 98140 62860 98360 62910
rect 98640 63090 98860 63140
rect 98640 63020 98650 63090
rect 98850 63020 98860 63090
rect 98640 62980 98860 63020
rect 98640 62910 98650 62980
rect 98850 62910 98860 62980
rect 98640 62860 98860 62910
rect 99140 63090 99360 63140
rect 99140 63020 99150 63090
rect 99350 63020 99360 63090
rect 99140 62980 99360 63020
rect 99140 62910 99150 62980
rect 99350 62910 99360 62980
rect 99140 62860 99360 62910
rect 99640 63090 99860 63140
rect 99640 63020 99650 63090
rect 99850 63020 99860 63090
rect 99640 62980 99860 63020
rect 99640 62910 99650 62980
rect 99850 62910 99860 62980
rect 99640 62860 99860 62910
rect -16000 62850 -12000 62860
rect -16000 62650 -15980 62850
rect -15910 62650 -15590 62850
rect -15520 62650 -15480 62850
rect -15410 62650 -15090 62850
rect -15020 62650 -14980 62850
rect -14910 62650 -14590 62850
rect -14520 62650 -14480 62850
rect -14410 62650 -14090 62850
rect -14020 62650 -13980 62850
rect -13910 62650 -13590 62850
rect -13520 62650 -13480 62850
rect -13410 62650 -13090 62850
rect -13020 62650 -12980 62850
rect -12910 62650 -12590 62850
rect -12520 62650 -12480 62850
rect -12410 62650 -12090 62850
rect -12020 62650 -12000 62850
rect -16000 62640 -12000 62650
rect 96000 62850 100000 62860
rect 96000 62650 96020 62850
rect 96090 62650 96410 62850
rect 96480 62650 96520 62850
rect 96590 62650 96910 62850
rect 96980 62650 97020 62850
rect 97090 62650 97410 62850
rect 97480 62650 97520 62850
rect 97590 62650 97910 62850
rect 97980 62650 98020 62850
rect 98090 62650 98410 62850
rect 98480 62650 98520 62850
rect 98590 62650 98910 62850
rect 98980 62650 99020 62850
rect 99090 62650 99410 62850
rect 99480 62650 99520 62850
rect 99590 62650 99910 62850
rect 99980 62650 100000 62850
rect 96000 62640 100000 62650
rect -15860 62590 -15640 62640
rect -15860 62520 -15850 62590
rect -15650 62520 -15640 62590
rect -15860 62480 -15640 62520
rect -15860 62410 -15850 62480
rect -15650 62410 -15640 62480
rect -15860 62360 -15640 62410
rect -15360 62590 -15140 62640
rect -15360 62520 -15350 62590
rect -15150 62520 -15140 62590
rect -15360 62480 -15140 62520
rect -15360 62410 -15350 62480
rect -15150 62410 -15140 62480
rect -15360 62360 -15140 62410
rect -14860 62590 -14640 62640
rect -14860 62520 -14850 62590
rect -14650 62520 -14640 62590
rect -14860 62480 -14640 62520
rect -14860 62410 -14850 62480
rect -14650 62410 -14640 62480
rect -14860 62360 -14640 62410
rect -14360 62590 -14140 62640
rect -14360 62520 -14350 62590
rect -14150 62520 -14140 62590
rect -14360 62480 -14140 62520
rect -14360 62410 -14350 62480
rect -14150 62410 -14140 62480
rect -14360 62360 -14140 62410
rect -13860 62590 -13640 62640
rect -13860 62520 -13850 62590
rect -13650 62520 -13640 62590
rect -13860 62480 -13640 62520
rect -13860 62410 -13850 62480
rect -13650 62410 -13640 62480
rect -13860 62360 -13640 62410
rect -13360 62590 -13140 62640
rect -13360 62520 -13350 62590
rect -13150 62520 -13140 62590
rect -13360 62480 -13140 62520
rect -13360 62410 -13350 62480
rect -13150 62410 -13140 62480
rect -13360 62360 -13140 62410
rect -12860 62590 -12640 62640
rect -12860 62520 -12850 62590
rect -12650 62520 -12640 62590
rect -12860 62480 -12640 62520
rect -12860 62410 -12850 62480
rect -12650 62410 -12640 62480
rect -12860 62360 -12640 62410
rect -12360 62590 -12140 62640
rect -12360 62520 -12350 62590
rect -12150 62520 -12140 62590
rect -12360 62480 -12140 62520
rect -12360 62410 -12350 62480
rect -12150 62410 -12140 62480
rect -12360 62360 -12140 62410
rect 96140 62590 96360 62640
rect 96140 62520 96150 62590
rect 96350 62520 96360 62590
rect 96140 62480 96360 62520
rect 96140 62410 96150 62480
rect 96350 62410 96360 62480
rect 96140 62360 96360 62410
rect 96640 62590 96860 62640
rect 96640 62520 96650 62590
rect 96850 62520 96860 62590
rect 96640 62480 96860 62520
rect 96640 62410 96650 62480
rect 96850 62410 96860 62480
rect 96640 62360 96860 62410
rect 97140 62590 97360 62640
rect 97140 62520 97150 62590
rect 97350 62520 97360 62590
rect 97140 62480 97360 62520
rect 97140 62410 97150 62480
rect 97350 62410 97360 62480
rect 97140 62360 97360 62410
rect 97640 62590 97860 62640
rect 97640 62520 97650 62590
rect 97850 62520 97860 62590
rect 97640 62480 97860 62520
rect 97640 62410 97650 62480
rect 97850 62410 97860 62480
rect 97640 62360 97860 62410
rect 98140 62590 98360 62640
rect 98140 62520 98150 62590
rect 98350 62520 98360 62590
rect 98140 62480 98360 62520
rect 98140 62410 98150 62480
rect 98350 62410 98360 62480
rect 98140 62360 98360 62410
rect 98640 62590 98860 62640
rect 98640 62520 98650 62590
rect 98850 62520 98860 62590
rect 98640 62480 98860 62520
rect 98640 62410 98650 62480
rect 98850 62410 98860 62480
rect 98640 62360 98860 62410
rect 99140 62590 99360 62640
rect 99140 62520 99150 62590
rect 99350 62520 99360 62590
rect 99140 62480 99360 62520
rect 99140 62410 99150 62480
rect 99350 62410 99360 62480
rect 99140 62360 99360 62410
rect 99640 62590 99860 62640
rect 99640 62520 99650 62590
rect 99850 62520 99860 62590
rect 99640 62480 99860 62520
rect 99640 62410 99650 62480
rect 99850 62410 99860 62480
rect 99640 62360 99860 62410
rect -16000 62350 -12000 62360
rect -16000 62150 -15980 62350
rect -15910 62150 -15590 62350
rect -15520 62150 -15480 62350
rect -15410 62150 -15090 62350
rect -15020 62150 -14980 62350
rect -14910 62150 -14590 62350
rect -14520 62150 -14480 62350
rect -14410 62150 -14090 62350
rect -14020 62150 -13980 62350
rect -13910 62150 -13590 62350
rect -13520 62150 -13480 62350
rect -13410 62150 -13090 62350
rect -13020 62150 -12980 62350
rect -12910 62150 -12590 62350
rect -12520 62150 -12480 62350
rect -12410 62150 -12090 62350
rect -12020 62150 -12000 62350
rect -16000 62140 -12000 62150
rect 96000 62350 100000 62360
rect 96000 62150 96020 62350
rect 96090 62150 96410 62350
rect 96480 62150 96520 62350
rect 96590 62150 96910 62350
rect 96980 62150 97020 62350
rect 97090 62150 97410 62350
rect 97480 62150 97520 62350
rect 97590 62150 97910 62350
rect 97980 62150 98020 62350
rect 98090 62150 98410 62350
rect 98480 62150 98520 62350
rect 98590 62150 98910 62350
rect 98980 62150 99020 62350
rect 99090 62150 99410 62350
rect 99480 62150 99520 62350
rect 99590 62150 99910 62350
rect 99980 62150 100000 62350
rect 96000 62140 100000 62150
rect -15860 62090 -15640 62140
rect -15860 62020 -15850 62090
rect -15650 62020 -15640 62090
rect -15860 61980 -15640 62020
rect -15860 61910 -15850 61980
rect -15650 61910 -15640 61980
rect -15860 61860 -15640 61910
rect -15360 62090 -15140 62140
rect -15360 62020 -15350 62090
rect -15150 62020 -15140 62090
rect -15360 61980 -15140 62020
rect -15360 61910 -15350 61980
rect -15150 61910 -15140 61980
rect -15360 61860 -15140 61910
rect -14860 62090 -14640 62140
rect -14860 62020 -14850 62090
rect -14650 62020 -14640 62090
rect -14860 61980 -14640 62020
rect -14860 61910 -14850 61980
rect -14650 61910 -14640 61980
rect -14860 61860 -14640 61910
rect -14360 62090 -14140 62140
rect -14360 62020 -14350 62090
rect -14150 62020 -14140 62090
rect -14360 61980 -14140 62020
rect -14360 61910 -14350 61980
rect -14150 61910 -14140 61980
rect -14360 61860 -14140 61910
rect -13860 62090 -13640 62140
rect -13860 62020 -13850 62090
rect -13650 62020 -13640 62090
rect -13860 61980 -13640 62020
rect -13860 61910 -13850 61980
rect -13650 61910 -13640 61980
rect -13860 61860 -13640 61910
rect -13360 62090 -13140 62140
rect -13360 62020 -13350 62090
rect -13150 62020 -13140 62090
rect -13360 61980 -13140 62020
rect -13360 61910 -13350 61980
rect -13150 61910 -13140 61980
rect -13360 61860 -13140 61910
rect -12860 62090 -12640 62140
rect -12860 62020 -12850 62090
rect -12650 62020 -12640 62090
rect -12860 61980 -12640 62020
rect -12860 61910 -12850 61980
rect -12650 61910 -12640 61980
rect -12860 61860 -12640 61910
rect -12360 62090 -12140 62140
rect -12360 62020 -12350 62090
rect -12150 62020 -12140 62090
rect -12360 61980 -12140 62020
rect -12360 61910 -12350 61980
rect -12150 61910 -12140 61980
rect -12360 61860 -12140 61910
rect 96140 62090 96360 62140
rect 96140 62020 96150 62090
rect 96350 62020 96360 62090
rect 96140 61980 96360 62020
rect 96140 61910 96150 61980
rect 96350 61910 96360 61980
rect 96140 61860 96360 61910
rect 96640 62090 96860 62140
rect 96640 62020 96650 62090
rect 96850 62020 96860 62090
rect 96640 61980 96860 62020
rect 96640 61910 96650 61980
rect 96850 61910 96860 61980
rect 96640 61860 96860 61910
rect 97140 62090 97360 62140
rect 97140 62020 97150 62090
rect 97350 62020 97360 62090
rect 97140 61980 97360 62020
rect 97140 61910 97150 61980
rect 97350 61910 97360 61980
rect 97140 61860 97360 61910
rect 97640 62090 97860 62140
rect 97640 62020 97650 62090
rect 97850 62020 97860 62090
rect 97640 61980 97860 62020
rect 97640 61910 97650 61980
rect 97850 61910 97860 61980
rect 97640 61860 97860 61910
rect 98140 62090 98360 62140
rect 98140 62020 98150 62090
rect 98350 62020 98360 62090
rect 98140 61980 98360 62020
rect 98140 61910 98150 61980
rect 98350 61910 98360 61980
rect 98140 61860 98360 61910
rect 98640 62090 98860 62140
rect 98640 62020 98650 62090
rect 98850 62020 98860 62090
rect 98640 61980 98860 62020
rect 98640 61910 98650 61980
rect 98850 61910 98860 61980
rect 98640 61860 98860 61910
rect 99140 62090 99360 62140
rect 99140 62020 99150 62090
rect 99350 62020 99360 62090
rect 99140 61980 99360 62020
rect 99140 61910 99150 61980
rect 99350 61910 99360 61980
rect 99140 61860 99360 61910
rect 99640 62090 99860 62140
rect 99640 62020 99650 62090
rect 99850 62020 99860 62090
rect 99640 61980 99860 62020
rect 99640 61910 99650 61980
rect 99850 61910 99860 61980
rect 99640 61860 99860 61910
rect -16000 61850 -12000 61860
rect -16000 61650 -15980 61850
rect -15910 61650 -15590 61850
rect -15520 61650 -15480 61850
rect -15410 61650 -15090 61850
rect -15020 61650 -14980 61850
rect -14910 61650 -14590 61850
rect -14520 61650 -14480 61850
rect -14410 61650 -14090 61850
rect -14020 61650 -13980 61850
rect -13910 61650 -13590 61850
rect -13520 61650 -13480 61850
rect -13410 61650 -13090 61850
rect -13020 61650 -12980 61850
rect -12910 61650 -12590 61850
rect -12520 61650 -12480 61850
rect -12410 61650 -12090 61850
rect -12020 61650 -12000 61850
rect -16000 61640 -12000 61650
rect 96000 61850 100000 61860
rect 96000 61650 96020 61850
rect 96090 61650 96410 61850
rect 96480 61650 96520 61850
rect 96590 61650 96910 61850
rect 96980 61650 97020 61850
rect 97090 61650 97410 61850
rect 97480 61650 97520 61850
rect 97590 61650 97910 61850
rect 97980 61650 98020 61850
rect 98090 61650 98410 61850
rect 98480 61650 98520 61850
rect 98590 61650 98910 61850
rect 98980 61650 99020 61850
rect 99090 61650 99410 61850
rect 99480 61650 99520 61850
rect 99590 61650 99910 61850
rect 99980 61650 100000 61850
rect 96000 61640 100000 61650
rect -15860 61590 -15640 61640
rect -15860 61520 -15850 61590
rect -15650 61520 -15640 61590
rect -15860 61480 -15640 61520
rect -15860 61410 -15850 61480
rect -15650 61410 -15640 61480
rect -15860 61360 -15640 61410
rect -15360 61590 -15140 61640
rect -15360 61520 -15350 61590
rect -15150 61520 -15140 61590
rect -15360 61480 -15140 61520
rect -15360 61410 -15350 61480
rect -15150 61410 -15140 61480
rect -15360 61360 -15140 61410
rect -14860 61590 -14640 61640
rect -14860 61520 -14850 61590
rect -14650 61520 -14640 61590
rect -14860 61480 -14640 61520
rect -14860 61410 -14850 61480
rect -14650 61410 -14640 61480
rect -14860 61360 -14640 61410
rect -14360 61590 -14140 61640
rect -14360 61520 -14350 61590
rect -14150 61520 -14140 61590
rect -14360 61480 -14140 61520
rect -14360 61410 -14350 61480
rect -14150 61410 -14140 61480
rect -14360 61360 -14140 61410
rect -13860 61590 -13640 61640
rect -13860 61520 -13850 61590
rect -13650 61520 -13640 61590
rect -13860 61480 -13640 61520
rect -13860 61410 -13850 61480
rect -13650 61410 -13640 61480
rect -13860 61360 -13640 61410
rect -13360 61590 -13140 61640
rect -13360 61520 -13350 61590
rect -13150 61520 -13140 61590
rect -13360 61480 -13140 61520
rect -13360 61410 -13350 61480
rect -13150 61410 -13140 61480
rect -13360 61360 -13140 61410
rect -12860 61590 -12640 61640
rect -12860 61520 -12850 61590
rect -12650 61520 -12640 61590
rect -12860 61480 -12640 61520
rect -12860 61410 -12850 61480
rect -12650 61410 -12640 61480
rect -12860 61360 -12640 61410
rect -12360 61590 -12140 61640
rect -12360 61520 -12350 61590
rect -12150 61520 -12140 61590
rect -12360 61480 -12140 61520
rect -12360 61410 -12350 61480
rect -12150 61410 -12140 61480
rect -12360 61360 -12140 61410
rect 96140 61590 96360 61640
rect 96140 61520 96150 61590
rect 96350 61520 96360 61590
rect 96140 61480 96360 61520
rect 96140 61410 96150 61480
rect 96350 61410 96360 61480
rect 96140 61360 96360 61410
rect 96640 61590 96860 61640
rect 96640 61520 96650 61590
rect 96850 61520 96860 61590
rect 96640 61480 96860 61520
rect 96640 61410 96650 61480
rect 96850 61410 96860 61480
rect 96640 61360 96860 61410
rect 97140 61590 97360 61640
rect 97140 61520 97150 61590
rect 97350 61520 97360 61590
rect 97140 61480 97360 61520
rect 97140 61410 97150 61480
rect 97350 61410 97360 61480
rect 97140 61360 97360 61410
rect 97640 61590 97860 61640
rect 97640 61520 97650 61590
rect 97850 61520 97860 61590
rect 97640 61480 97860 61520
rect 97640 61410 97650 61480
rect 97850 61410 97860 61480
rect 97640 61360 97860 61410
rect 98140 61590 98360 61640
rect 98140 61520 98150 61590
rect 98350 61520 98360 61590
rect 98140 61480 98360 61520
rect 98140 61410 98150 61480
rect 98350 61410 98360 61480
rect 98140 61360 98360 61410
rect 98640 61590 98860 61640
rect 98640 61520 98650 61590
rect 98850 61520 98860 61590
rect 98640 61480 98860 61520
rect 98640 61410 98650 61480
rect 98850 61410 98860 61480
rect 98640 61360 98860 61410
rect 99140 61590 99360 61640
rect 99140 61520 99150 61590
rect 99350 61520 99360 61590
rect 99140 61480 99360 61520
rect 99140 61410 99150 61480
rect 99350 61410 99360 61480
rect 99140 61360 99360 61410
rect 99640 61590 99860 61640
rect 99640 61520 99650 61590
rect 99850 61520 99860 61590
rect 99640 61480 99860 61520
rect 99640 61410 99650 61480
rect 99850 61410 99860 61480
rect 99640 61360 99860 61410
rect -16000 61350 -12000 61360
rect -16000 61150 -15980 61350
rect -15910 61150 -15590 61350
rect -15520 61150 -15480 61350
rect -15410 61150 -15090 61350
rect -15020 61150 -14980 61350
rect -14910 61150 -14590 61350
rect -14520 61150 -14480 61350
rect -14410 61150 -14090 61350
rect -14020 61150 -13980 61350
rect -13910 61150 -13590 61350
rect -13520 61150 -13480 61350
rect -13410 61150 -13090 61350
rect -13020 61150 -12980 61350
rect -12910 61150 -12590 61350
rect -12520 61150 -12480 61350
rect -12410 61150 -12090 61350
rect -12020 61150 -12000 61350
rect -16000 61140 -12000 61150
rect 96000 61350 100000 61360
rect 96000 61150 96020 61350
rect 96090 61150 96410 61350
rect 96480 61150 96520 61350
rect 96590 61150 96910 61350
rect 96980 61150 97020 61350
rect 97090 61150 97410 61350
rect 97480 61150 97520 61350
rect 97590 61150 97910 61350
rect 97980 61150 98020 61350
rect 98090 61150 98410 61350
rect 98480 61150 98520 61350
rect 98590 61150 98910 61350
rect 98980 61150 99020 61350
rect 99090 61150 99410 61350
rect 99480 61150 99520 61350
rect 99590 61150 99910 61350
rect 99980 61150 100000 61350
rect 96000 61140 100000 61150
rect -15860 61090 -15640 61140
rect -15860 61020 -15850 61090
rect -15650 61020 -15640 61090
rect -15860 60980 -15640 61020
rect -15860 60910 -15850 60980
rect -15650 60910 -15640 60980
rect -15860 60860 -15640 60910
rect -15360 61090 -15140 61140
rect -15360 61020 -15350 61090
rect -15150 61020 -15140 61090
rect -15360 60980 -15140 61020
rect -15360 60910 -15350 60980
rect -15150 60910 -15140 60980
rect -15360 60860 -15140 60910
rect -14860 61090 -14640 61140
rect -14860 61020 -14850 61090
rect -14650 61020 -14640 61090
rect -14860 60980 -14640 61020
rect -14860 60910 -14850 60980
rect -14650 60910 -14640 60980
rect -14860 60860 -14640 60910
rect -14360 61090 -14140 61140
rect -14360 61020 -14350 61090
rect -14150 61020 -14140 61090
rect -14360 60980 -14140 61020
rect -14360 60910 -14350 60980
rect -14150 60910 -14140 60980
rect -14360 60860 -14140 60910
rect -13860 61090 -13640 61140
rect -13860 61020 -13850 61090
rect -13650 61020 -13640 61090
rect -13860 60980 -13640 61020
rect -13860 60910 -13850 60980
rect -13650 60910 -13640 60980
rect -13860 60860 -13640 60910
rect -13360 61090 -13140 61140
rect -13360 61020 -13350 61090
rect -13150 61020 -13140 61090
rect -13360 60980 -13140 61020
rect -13360 60910 -13350 60980
rect -13150 60910 -13140 60980
rect -13360 60860 -13140 60910
rect -12860 61090 -12640 61140
rect -12860 61020 -12850 61090
rect -12650 61020 -12640 61090
rect -12860 60980 -12640 61020
rect -12860 60910 -12850 60980
rect -12650 60910 -12640 60980
rect -12860 60860 -12640 60910
rect -12360 61090 -12140 61140
rect -12360 61020 -12350 61090
rect -12150 61020 -12140 61090
rect -12360 60980 -12140 61020
rect -12360 60910 -12350 60980
rect -12150 60910 -12140 60980
rect -12360 60860 -12140 60910
rect 96140 61090 96360 61140
rect 96140 61020 96150 61090
rect 96350 61020 96360 61090
rect 96140 60980 96360 61020
rect 96140 60910 96150 60980
rect 96350 60910 96360 60980
rect 96140 60860 96360 60910
rect 96640 61090 96860 61140
rect 96640 61020 96650 61090
rect 96850 61020 96860 61090
rect 96640 60980 96860 61020
rect 96640 60910 96650 60980
rect 96850 60910 96860 60980
rect 96640 60860 96860 60910
rect 97140 61090 97360 61140
rect 97140 61020 97150 61090
rect 97350 61020 97360 61090
rect 97140 60980 97360 61020
rect 97140 60910 97150 60980
rect 97350 60910 97360 60980
rect 97140 60860 97360 60910
rect 97640 61090 97860 61140
rect 97640 61020 97650 61090
rect 97850 61020 97860 61090
rect 97640 60980 97860 61020
rect 97640 60910 97650 60980
rect 97850 60910 97860 60980
rect 97640 60860 97860 60910
rect 98140 61090 98360 61140
rect 98140 61020 98150 61090
rect 98350 61020 98360 61090
rect 98140 60980 98360 61020
rect 98140 60910 98150 60980
rect 98350 60910 98360 60980
rect 98140 60860 98360 60910
rect 98640 61090 98860 61140
rect 98640 61020 98650 61090
rect 98850 61020 98860 61090
rect 98640 60980 98860 61020
rect 98640 60910 98650 60980
rect 98850 60910 98860 60980
rect 98640 60860 98860 60910
rect 99140 61090 99360 61140
rect 99140 61020 99150 61090
rect 99350 61020 99360 61090
rect 99140 60980 99360 61020
rect 99140 60910 99150 60980
rect 99350 60910 99360 60980
rect 99140 60860 99360 60910
rect 99640 61090 99860 61140
rect 99640 61020 99650 61090
rect 99850 61020 99860 61090
rect 99640 60980 99860 61020
rect 99640 60910 99650 60980
rect 99850 60910 99860 60980
rect 99640 60860 99860 60910
rect -16000 60850 -12000 60860
rect -16000 60650 -15980 60850
rect -15910 60650 -15590 60850
rect -15520 60650 -15480 60850
rect -15410 60650 -15090 60850
rect -15020 60650 -14980 60850
rect -14910 60650 -14590 60850
rect -14520 60650 -14480 60850
rect -14410 60650 -14090 60850
rect -14020 60650 -13980 60850
rect -13910 60650 -13590 60850
rect -13520 60650 -13480 60850
rect -13410 60650 -13090 60850
rect -13020 60650 -12980 60850
rect -12910 60650 -12590 60850
rect -12520 60650 -12480 60850
rect -12410 60650 -12090 60850
rect -12020 60650 -12000 60850
rect -16000 60640 -12000 60650
rect 96000 60850 100000 60860
rect 96000 60650 96020 60850
rect 96090 60650 96410 60850
rect 96480 60650 96520 60850
rect 96590 60650 96910 60850
rect 96980 60650 97020 60850
rect 97090 60650 97410 60850
rect 97480 60650 97520 60850
rect 97590 60650 97910 60850
rect 97980 60650 98020 60850
rect 98090 60650 98410 60850
rect 98480 60650 98520 60850
rect 98590 60650 98910 60850
rect 98980 60650 99020 60850
rect 99090 60650 99410 60850
rect 99480 60650 99520 60850
rect 99590 60650 99910 60850
rect 99980 60650 100000 60850
rect 96000 60640 100000 60650
rect -15860 60590 -15640 60640
rect -15860 60520 -15850 60590
rect -15650 60520 -15640 60590
rect -15860 60480 -15640 60520
rect -15860 60410 -15850 60480
rect -15650 60410 -15640 60480
rect -15860 60360 -15640 60410
rect -15360 60590 -15140 60640
rect -15360 60520 -15350 60590
rect -15150 60520 -15140 60590
rect -15360 60480 -15140 60520
rect -15360 60410 -15350 60480
rect -15150 60410 -15140 60480
rect -15360 60360 -15140 60410
rect -14860 60590 -14640 60640
rect -14860 60520 -14850 60590
rect -14650 60520 -14640 60590
rect -14860 60480 -14640 60520
rect -14860 60410 -14850 60480
rect -14650 60410 -14640 60480
rect -14860 60360 -14640 60410
rect -14360 60590 -14140 60640
rect -14360 60520 -14350 60590
rect -14150 60520 -14140 60590
rect -14360 60480 -14140 60520
rect -14360 60410 -14350 60480
rect -14150 60410 -14140 60480
rect -14360 60360 -14140 60410
rect -13860 60590 -13640 60640
rect -13860 60520 -13850 60590
rect -13650 60520 -13640 60590
rect -13860 60480 -13640 60520
rect -13860 60410 -13850 60480
rect -13650 60410 -13640 60480
rect -13860 60360 -13640 60410
rect -13360 60590 -13140 60640
rect -13360 60520 -13350 60590
rect -13150 60520 -13140 60590
rect -13360 60480 -13140 60520
rect -13360 60410 -13350 60480
rect -13150 60410 -13140 60480
rect -13360 60360 -13140 60410
rect -12860 60590 -12640 60640
rect -12860 60520 -12850 60590
rect -12650 60520 -12640 60590
rect -12860 60480 -12640 60520
rect -12860 60410 -12850 60480
rect -12650 60410 -12640 60480
rect -12860 60360 -12640 60410
rect -12360 60590 -12140 60640
rect -12360 60520 -12350 60590
rect -12150 60520 -12140 60590
rect -12360 60480 -12140 60520
rect -12360 60410 -12350 60480
rect -12150 60410 -12140 60480
rect -12360 60360 -12140 60410
rect 96140 60590 96360 60640
rect 96140 60520 96150 60590
rect 96350 60520 96360 60590
rect 96140 60480 96360 60520
rect 96140 60410 96150 60480
rect 96350 60410 96360 60480
rect 96140 60360 96360 60410
rect 96640 60590 96860 60640
rect 96640 60520 96650 60590
rect 96850 60520 96860 60590
rect 96640 60480 96860 60520
rect 96640 60410 96650 60480
rect 96850 60410 96860 60480
rect 96640 60360 96860 60410
rect 97140 60590 97360 60640
rect 97140 60520 97150 60590
rect 97350 60520 97360 60590
rect 97140 60480 97360 60520
rect 97140 60410 97150 60480
rect 97350 60410 97360 60480
rect 97140 60360 97360 60410
rect 97640 60590 97860 60640
rect 97640 60520 97650 60590
rect 97850 60520 97860 60590
rect 97640 60480 97860 60520
rect 97640 60410 97650 60480
rect 97850 60410 97860 60480
rect 97640 60360 97860 60410
rect 98140 60590 98360 60640
rect 98140 60520 98150 60590
rect 98350 60520 98360 60590
rect 98140 60480 98360 60520
rect 98140 60410 98150 60480
rect 98350 60410 98360 60480
rect 98140 60360 98360 60410
rect 98640 60590 98860 60640
rect 98640 60520 98650 60590
rect 98850 60520 98860 60590
rect 98640 60480 98860 60520
rect 98640 60410 98650 60480
rect 98850 60410 98860 60480
rect 98640 60360 98860 60410
rect 99140 60590 99360 60640
rect 99140 60520 99150 60590
rect 99350 60520 99360 60590
rect 99140 60480 99360 60520
rect 99140 60410 99150 60480
rect 99350 60410 99360 60480
rect 99140 60360 99360 60410
rect 99640 60590 99860 60640
rect 99640 60520 99650 60590
rect 99850 60520 99860 60590
rect 99640 60480 99860 60520
rect 99640 60410 99650 60480
rect 99850 60410 99860 60480
rect 99640 60360 99860 60410
rect -16000 60350 -12000 60360
rect -16000 60150 -15980 60350
rect -15910 60150 -15590 60350
rect -15520 60150 -15480 60350
rect -15410 60150 -15090 60350
rect -15020 60150 -14980 60350
rect -14910 60150 -14590 60350
rect -14520 60150 -14480 60350
rect -14410 60150 -14090 60350
rect -14020 60150 -13980 60350
rect -13910 60150 -13590 60350
rect -13520 60150 -13480 60350
rect -13410 60150 -13090 60350
rect -13020 60150 -12980 60350
rect -12910 60150 -12590 60350
rect -12520 60150 -12480 60350
rect -12410 60150 -12090 60350
rect -12020 60150 -12000 60350
rect -16000 60140 -12000 60150
rect 96000 60350 100000 60360
rect 96000 60150 96020 60350
rect 96090 60150 96410 60350
rect 96480 60150 96520 60350
rect 96590 60150 96910 60350
rect 96980 60150 97020 60350
rect 97090 60150 97410 60350
rect 97480 60150 97520 60350
rect 97590 60150 97910 60350
rect 97980 60150 98020 60350
rect 98090 60150 98410 60350
rect 98480 60150 98520 60350
rect 98590 60150 98910 60350
rect 98980 60150 99020 60350
rect 99090 60150 99410 60350
rect 99480 60150 99520 60350
rect 99590 60150 99910 60350
rect 99980 60150 100000 60350
rect 96000 60140 100000 60150
rect -15860 60090 -15640 60140
rect -15860 60020 -15850 60090
rect -15650 60020 -15640 60090
rect -15860 59980 -15640 60020
rect -15860 59910 -15850 59980
rect -15650 59910 -15640 59980
rect -15860 59860 -15640 59910
rect -15360 60090 -15140 60140
rect -15360 60020 -15350 60090
rect -15150 60020 -15140 60090
rect -15360 59980 -15140 60020
rect -15360 59910 -15350 59980
rect -15150 59910 -15140 59980
rect -15360 59860 -15140 59910
rect -14860 60090 -14640 60140
rect -14860 60020 -14850 60090
rect -14650 60020 -14640 60090
rect -14860 59980 -14640 60020
rect -14860 59910 -14850 59980
rect -14650 59910 -14640 59980
rect -14860 59860 -14640 59910
rect -14360 60090 -14140 60140
rect -14360 60020 -14350 60090
rect -14150 60020 -14140 60090
rect -14360 59980 -14140 60020
rect -14360 59910 -14350 59980
rect -14150 59910 -14140 59980
rect -14360 59860 -14140 59910
rect -13860 60090 -13640 60140
rect -13860 60020 -13850 60090
rect -13650 60020 -13640 60090
rect -13860 59980 -13640 60020
rect -13860 59910 -13850 59980
rect -13650 59910 -13640 59980
rect -13860 59860 -13640 59910
rect -13360 60090 -13140 60140
rect -13360 60020 -13350 60090
rect -13150 60020 -13140 60090
rect -13360 59980 -13140 60020
rect -13360 59910 -13350 59980
rect -13150 59910 -13140 59980
rect -13360 59860 -13140 59910
rect -12860 60090 -12640 60140
rect -12860 60020 -12850 60090
rect -12650 60020 -12640 60090
rect -12860 59980 -12640 60020
rect -12860 59910 -12850 59980
rect -12650 59910 -12640 59980
rect -12860 59860 -12640 59910
rect -12360 60090 -12140 60140
rect -12360 60020 -12350 60090
rect -12150 60020 -12140 60090
rect -12360 59980 -12140 60020
rect -12360 59910 -12350 59980
rect -12150 59910 -12140 59980
rect -12360 59860 -12140 59910
rect 96140 60090 96360 60140
rect 96140 60020 96150 60090
rect 96350 60020 96360 60090
rect 96140 59980 96360 60020
rect 96140 59910 96150 59980
rect 96350 59910 96360 59980
rect 96140 59860 96360 59910
rect 96640 60090 96860 60140
rect 96640 60020 96650 60090
rect 96850 60020 96860 60090
rect 96640 59980 96860 60020
rect 96640 59910 96650 59980
rect 96850 59910 96860 59980
rect 96640 59860 96860 59910
rect 97140 60090 97360 60140
rect 97140 60020 97150 60090
rect 97350 60020 97360 60090
rect 97140 59980 97360 60020
rect 97140 59910 97150 59980
rect 97350 59910 97360 59980
rect 97140 59860 97360 59910
rect 97640 60090 97860 60140
rect 97640 60020 97650 60090
rect 97850 60020 97860 60090
rect 97640 59980 97860 60020
rect 97640 59910 97650 59980
rect 97850 59910 97860 59980
rect 97640 59860 97860 59910
rect 98140 60090 98360 60140
rect 98140 60020 98150 60090
rect 98350 60020 98360 60090
rect 98140 59980 98360 60020
rect 98140 59910 98150 59980
rect 98350 59910 98360 59980
rect 98140 59860 98360 59910
rect 98640 60090 98860 60140
rect 98640 60020 98650 60090
rect 98850 60020 98860 60090
rect 98640 59980 98860 60020
rect 98640 59910 98650 59980
rect 98850 59910 98860 59980
rect 98640 59860 98860 59910
rect 99140 60090 99360 60140
rect 99140 60020 99150 60090
rect 99350 60020 99360 60090
rect 99140 59980 99360 60020
rect 99140 59910 99150 59980
rect 99350 59910 99360 59980
rect 99140 59860 99360 59910
rect 99640 60090 99860 60140
rect 99640 60020 99650 60090
rect 99850 60020 99860 60090
rect 99640 59980 99860 60020
rect 99640 59910 99650 59980
rect 99850 59910 99860 59980
rect 99640 59860 99860 59910
rect -16000 59850 -12000 59860
rect -16000 59650 -15980 59850
rect -15910 59650 -15590 59850
rect -15520 59650 -15480 59850
rect -15410 59650 -15090 59850
rect -15020 59650 -14980 59850
rect -14910 59650 -14590 59850
rect -14520 59650 -14480 59850
rect -14410 59650 -14090 59850
rect -14020 59650 -13980 59850
rect -13910 59650 -13590 59850
rect -13520 59650 -13480 59850
rect -13410 59650 -13090 59850
rect -13020 59650 -12980 59850
rect -12910 59650 -12590 59850
rect -12520 59650 -12480 59850
rect -12410 59650 -12090 59850
rect -12020 59650 -12000 59850
rect -16000 59640 -12000 59650
rect 96000 59850 100000 59860
rect 96000 59650 96020 59850
rect 96090 59650 96410 59850
rect 96480 59650 96520 59850
rect 96590 59650 96910 59850
rect 96980 59650 97020 59850
rect 97090 59650 97410 59850
rect 97480 59650 97520 59850
rect 97590 59650 97910 59850
rect 97980 59650 98020 59850
rect 98090 59650 98410 59850
rect 98480 59650 98520 59850
rect 98590 59650 98910 59850
rect 98980 59650 99020 59850
rect 99090 59650 99410 59850
rect 99480 59650 99520 59850
rect 99590 59650 99910 59850
rect 99980 59650 100000 59850
rect 96000 59640 100000 59650
rect -15860 59590 -15640 59640
rect -15860 59520 -15850 59590
rect -15650 59520 -15640 59590
rect -15860 59480 -15640 59520
rect -15860 59410 -15850 59480
rect -15650 59410 -15640 59480
rect -15860 59360 -15640 59410
rect -15360 59590 -15140 59640
rect -15360 59520 -15350 59590
rect -15150 59520 -15140 59590
rect -15360 59480 -15140 59520
rect -15360 59410 -15350 59480
rect -15150 59410 -15140 59480
rect -15360 59360 -15140 59410
rect -14860 59590 -14640 59640
rect -14860 59520 -14850 59590
rect -14650 59520 -14640 59590
rect -14860 59480 -14640 59520
rect -14860 59410 -14850 59480
rect -14650 59410 -14640 59480
rect -14860 59360 -14640 59410
rect -14360 59590 -14140 59640
rect -14360 59520 -14350 59590
rect -14150 59520 -14140 59590
rect -14360 59480 -14140 59520
rect -14360 59410 -14350 59480
rect -14150 59410 -14140 59480
rect -14360 59360 -14140 59410
rect -13860 59590 -13640 59640
rect -13860 59520 -13850 59590
rect -13650 59520 -13640 59590
rect -13860 59480 -13640 59520
rect -13860 59410 -13850 59480
rect -13650 59410 -13640 59480
rect -13860 59360 -13640 59410
rect -13360 59590 -13140 59640
rect -13360 59520 -13350 59590
rect -13150 59520 -13140 59590
rect -13360 59480 -13140 59520
rect -13360 59410 -13350 59480
rect -13150 59410 -13140 59480
rect -13360 59360 -13140 59410
rect -12860 59590 -12640 59640
rect -12860 59520 -12850 59590
rect -12650 59520 -12640 59590
rect -12860 59480 -12640 59520
rect -12860 59410 -12850 59480
rect -12650 59410 -12640 59480
rect -12860 59360 -12640 59410
rect -12360 59590 -12140 59640
rect -12360 59520 -12350 59590
rect -12150 59520 -12140 59590
rect -12360 59480 -12140 59520
rect -12360 59410 -12350 59480
rect -12150 59410 -12140 59480
rect -12360 59360 -12140 59410
rect 96140 59590 96360 59640
rect 96140 59520 96150 59590
rect 96350 59520 96360 59590
rect 96140 59480 96360 59520
rect 96140 59410 96150 59480
rect 96350 59410 96360 59480
rect 96140 59360 96360 59410
rect 96640 59590 96860 59640
rect 96640 59520 96650 59590
rect 96850 59520 96860 59590
rect 96640 59480 96860 59520
rect 96640 59410 96650 59480
rect 96850 59410 96860 59480
rect 96640 59360 96860 59410
rect 97140 59590 97360 59640
rect 97140 59520 97150 59590
rect 97350 59520 97360 59590
rect 97140 59480 97360 59520
rect 97140 59410 97150 59480
rect 97350 59410 97360 59480
rect 97140 59360 97360 59410
rect 97640 59590 97860 59640
rect 97640 59520 97650 59590
rect 97850 59520 97860 59590
rect 97640 59480 97860 59520
rect 97640 59410 97650 59480
rect 97850 59410 97860 59480
rect 97640 59360 97860 59410
rect 98140 59590 98360 59640
rect 98140 59520 98150 59590
rect 98350 59520 98360 59590
rect 98140 59480 98360 59520
rect 98140 59410 98150 59480
rect 98350 59410 98360 59480
rect 98140 59360 98360 59410
rect 98640 59590 98860 59640
rect 98640 59520 98650 59590
rect 98850 59520 98860 59590
rect 98640 59480 98860 59520
rect 98640 59410 98650 59480
rect 98850 59410 98860 59480
rect 98640 59360 98860 59410
rect 99140 59590 99360 59640
rect 99140 59520 99150 59590
rect 99350 59520 99360 59590
rect 99140 59480 99360 59520
rect 99140 59410 99150 59480
rect 99350 59410 99360 59480
rect 99140 59360 99360 59410
rect 99640 59590 99860 59640
rect 99640 59520 99650 59590
rect 99850 59520 99860 59590
rect 99640 59480 99860 59520
rect 99640 59410 99650 59480
rect 99850 59410 99860 59480
rect 99640 59360 99860 59410
rect -16000 59350 -12000 59360
rect -16000 59150 -15980 59350
rect -15910 59150 -15590 59350
rect -15520 59150 -15480 59350
rect -15410 59150 -15090 59350
rect -15020 59150 -14980 59350
rect -14910 59150 -14590 59350
rect -14520 59150 -14480 59350
rect -14410 59150 -14090 59350
rect -14020 59150 -13980 59350
rect -13910 59150 -13590 59350
rect -13520 59150 -13480 59350
rect -13410 59150 -13090 59350
rect -13020 59150 -12980 59350
rect -12910 59150 -12590 59350
rect -12520 59150 -12480 59350
rect -12410 59150 -12090 59350
rect -12020 59150 -12000 59350
rect -16000 59140 -12000 59150
rect 96000 59350 100000 59360
rect 96000 59150 96020 59350
rect 96090 59150 96410 59350
rect 96480 59150 96520 59350
rect 96590 59150 96910 59350
rect 96980 59150 97020 59350
rect 97090 59150 97410 59350
rect 97480 59150 97520 59350
rect 97590 59150 97910 59350
rect 97980 59150 98020 59350
rect 98090 59150 98410 59350
rect 98480 59150 98520 59350
rect 98590 59150 98910 59350
rect 98980 59150 99020 59350
rect 99090 59150 99410 59350
rect 99480 59150 99520 59350
rect 99590 59150 99910 59350
rect 99980 59150 100000 59350
rect 96000 59140 100000 59150
rect -15860 59090 -15640 59140
rect -15860 59020 -15850 59090
rect -15650 59020 -15640 59090
rect -15860 58980 -15640 59020
rect -15860 58910 -15850 58980
rect -15650 58910 -15640 58980
rect -15860 58860 -15640 58910
rect -15360 59090 -15140 59140
rect -15360 59020 -15350 59090
rect -15150 59020 -15140 59090
rect -15360 58980 -15140 59020
rect -15360 58910 -15350 58980
rect -15150 58910 -15140 58980
rect -15360 58860 -15140 58910
rect -14860 59090 -14640 59140
rect -14860 59020 -14850 59090
rect -14650 59020 -14640 59090
rect -14860 58980 -14640 59020
rect -14860 58910 -14850 58980
rect -14650 58910 -14640 58980
rect -14860 58860 -14640 58910
rect -14360 59090 -14140 59140
rect -14360 59020 -14350 59090
rect -14150 59020 -14140 59090
rect -14360 58980 -14140 59020
rect -14360 58910 -14350 58980
rect -14150 58910 -14140 58980
rect -14360 58860 -14140 58910
rect -13860 59090 -13640 59140
rect -13860 59020 -13850 59090
rect -13650 59020 -13640 59090
rect -13860 58980 -13640 59020
rect -13860 58910 -13850 58980
rect -13650 58910 -13640 58980
rect -13860 58860 -13640 58910
rect -13360 59090 -13140 59140
rect -13360 59020 -13350 59090
rect -13150 59020 -13140 59090
rect -13360 58980 -13140 59020
rect -13360 58910 -13350 58980
rect -13150 58910 -13140 58980
rect -13360 58860 -13140 58910
rect -12860 59090 -12640 59140
rect -12860 59020 -12850 59090
rect -12650 59020 -12640 59090
rect -12860 58980 -12640 59020
rect -12860 58910 -12850 58980
rect -12650 58910 -12640 58980
rect -12860 58860 -12640 58910
rect -12360 59090 -12140 59140
rect -12360 59020 -12350 59090
rect -12150 59020 -12140 59090
rect -12360 58980 -12140 59020
rect -12360 58910 -12350 58980
rect -12150 58910 -12140 58980
rect -12360 58860 -12140 58910
rect 96140 59090 96360 59140
rect 96140 59020 96150 59090
rect 96350 59020 96360 59090
rect 96140 58980 96360 59020
rect 96140 58910 96150 58980
rect 96350 58910 96360 58980
rect 96140 58860 96360 58910
rect 96640 59090 96860 59140
rect 96640 59020 96650 59090
rect 96850 59020 96860 59090
rect 96640 58980 96860 59020
rect 96640 58910 96650 58980
rect 96850 58910 96860 58980
rect 96640 58860 96860 58910
rect 97140 59090 97360 59140
rect 97140 59020 97150 59090
rect 97350 59020 97360 59090
rect 97140 58980 97360 59020
rect 97140 58910 97150 58980
rect 97350 58910 97360 58980
rect 97140 58860 97360 58910
rect 97640 59090 97860 59140
rect 97640 59020 97650 59090
rect 97850 59020 97860 59090
rect 97640 58980 97860 59020
rect 97640 58910 97650 58980
rect 97850 58910 97860 58980
rect 97640 58860 97860 58910
rect 98140 59090 98360 59140
rect 98140 59020 98150 59090
rect 98350 59020 98360 59090
rect 98140 58980 98360 59020
rect 98140 58910 98150 58980
rect 98350 58910 98360 58980
rect 98140 58860 98360 58910
rect 98640 59090 98860 59140
rect 98640 59020 98650 59090
rect 98850 59020 98860 59090
rect 98640 58980 98860 59020
rect 98640 58910 98650 58980
rect 98850 58910 98860 58980
rect 98640 58860 98860 58910
rect 99140 59090 99360 59140
rect 99140 59020 99150 59090
rect 99350 59020 99360 59090
rect 99140 58980 99360 59020
rect 99140 58910 99150 58980
rect 99350 58910 99360 58980
rect 99140 58860 99360 58910
rect 99640 59090 99860 59140
rect 99640 59020 99650 59090
rect 99850 59020 99860 59090
rect 99640 58980 99860 59020
rect 99640 58910 99650 58980
rect 99850 58910 99860 58980
rect 99640 58860 99860 58910
rect -16000 58850 -12000 58860
rect -16000 58650 -15980 58850
rect -15910 58650 -15590 58850
rect -15520 58650 -15480 58850
rect -15410 58650 -15090 58850
rect -15020 58650 -14980 58850
rect -14910 58650 -14590 58850
rect -14520 58650 -14480 58850
rect -14410 58650 -14090 58850
rect -14020 58650 -13980 58850
rect -13910 58650 -13590 58850
rect -13520 58650 -13480 58850
rect -13410 58650 -13090 58850
rect -13020 58650 -12980 58850
rect -12910 58650 -12590 58850
rect -12520 58650 -12480 58850
rect -12410 58650 -12090 58850
rect -12020 58650 -12000 58850
rect -16000 58640 -12000 58650
rect 96000 58850 100000 58860
rect 96000 58650 96020 58850
rect 96090 58650 96410 58850
rect 96480 58650 96520 58850
rect 96590 58650 96910 58850
rect 96980 58650 97020 58850
rect 97090 58650 97410 58850
rect 97480 58650 97520 58850
rect 97590 58650 97910 58850
rect 97980 58650 98020 58850
rect 98090 58650 98410 58850
rect 98480 58650 98520 58850
rect 98590 58650 98910 58850
rect 98980 58650 99020 58850
rect 99090 58650 99410 58850
rect 99480 58650 99520 58850
rect 99590 58650 99910 58850
rect 99980 58650 100000 58850
rect 96000 58640 100000 58650
rect -15860 58590 -15640 58640
rect -15860 58520 -15850 58590
rect -15650 58520 -15640 58590
rect -15860 58480 -15640 58520
rect -15860 58410 -15850 58480
rect -15650 58410 -15640 58480
rect -15860 58360 -15640 58410
rect -15360 58590 -15140 58640
rect -15360 58520 -15350 58590
rect -15150 58520 -15140 58590
rect -15360 58480 -15140 58520
rect -15360 58410 -15350 58480
rect -15150 58410 -15140 58480
rect -15360 58360 -15140 58410
rect -14860 58590 -14640 58640
rect -14860 58520 -14850 58590
rect -14650 58520 -14640 58590
rect -14860 58480 -14640 58520
rect -14860 58410 -14850 58480
rect -14650 58410 -14640 58480
rect -14860 58360 -14640 58410
rect -14360 58590 -14140 58640
rect -14360 58520 -14350 58590
rect -14150 58520 -14140 58590
rect -14360 58480 -14140 58520
rect -14360 58410 -14350 58480
rect -14150 58410 -14140 58480
rect -14360 58360 -14140 58410
rect -13860 58590 -13640 58640
rect -13860 58520 -13850 58590
rect -13650 58520 -13640 58590
rect -13860 58480 -13640 58520
rect -13860 58410 -13850 58480
rect -13650 58410 -13640 58480
rect -13860 58360 -13640 58410
rect -13360 58590 -13140 58640
rect -13360 58520 -13350 58590
rect -13150 58520 -13140 58590
rect -13360 58480 -13140 58520
rect -13360 58410 -13350 58480
rect -13150 58410 -13140 58480
rect -13360 58360 -13140 58410
rect -12860 58590 -12640 58640
rect -12860 58520 -12850 58590
rect -12650 58520 -12640 58590
rect -12860 58480 -12640 58520
rect -12860 58410 -12850 58480
rect -12650 58410 -12640 58480
rect -12860 58360 -12640 58410
rect -12360 58590 -12140 58640
rect -12360 58520 -12350 58590
rect -12150 58520 -12140 58590
rect -12360 58480 -12140 58520
rect -12360 58410 -12350 58480
rect -12150 58410 -12140 58480
rect -12360 58360 -12140 58410
rect 96140 58590 96360 58640
rect 96140 58520 96150 58590
rect 96350 58520 96360 58590
rect 96140 58480 96360 58520
rect 96140 58410 96150 58480
rect 96350 58410 96360 58480
rect 96140 58360 96360 58410
rect 96640 58590 96860 58640
rect 96640 58520 96650 58590
rect 96850 58520 96860 58590
rect 96640 58480 96860 58520
rect 96640 58410 96650 58480
rect 96850 58410 96860 58480
rect 96640 58360 96860 58410
rect 97140 58590 97360 58640
rect 97140 58520 97150 58590
rect 97350 58520 97360 58590
rect 97140 58480 97360 58520
rect 97140 58410 97150 58480
rect 97350 58410 97360 58480
rect 97140 58360 97360 58410
rect 97640 58590 97860 58640
rect 97640 58520 97650 58590
rect 97850 58520 97860 58590
rect 97640 58480 97860 58520
rect 97640 58410 97650 58480
rect 97850 58410 97860 58480
rect 97640 58360 97860 58410
rect 98140 58590 98360 58640
rect 98140 58520 98150 58590
rect 98350 58520 98360 58590
rect 98140 58480 98360 58520
rect 98140 58410 98150 58480
rect 98350 58410 98360 58480
rect 98140 58360 98360 58410
rect 98640 58590 98860 58640
rect 98640 58520 98650 58590
rect 98850 58520 98860 58590
rect 98640 58480 98860 58520
rect 98640 58410 98650 58480
rect 98850 58410 98860 58480
rect 98640 58360 98860 58410
rect 99140 58590 99360 58640
rect 99140 58520 99150 58590
rect 99350 58520 99360 58590
rect 99140 58480 99360 58520
rect 99140 58410 99150 58480
rect 99350 58410 99360 58480
rect 99140 58360 99360 58410
rect 99640 58590 99860 58640
rect 99640 58520 99650 58590
rect 99850 58520 99860 58590
rect 99640 58480 99860 58520
rect 99640 58410 99650 58480
rect 99850 58410 99860 58480
rect 99640 58360 99860 58410
rect -16000 58350 -12000 58360
rect -16000 58150 -15980 58350
rect -15910 58150 -15590 58350
rect -15520 58150 -15480 58350
rect -15410 58150 -15090 58350
rect -15020 58150 -14980 58350
rect -14910 58150 -14590 58350
rect -14520 58150 -14480 58350
rect -14410 58150 -14090 58350
rect -14020 58150 -13980 58350
rect -13910 58150 -13590 58350
rect -13520 58150 -13480 58350
rect -13410 58150 -13090 58350
rect -13020 58150 -12980 58350
rect -12910 58150 -12590 58350
rect -12520 58150 -12480 58350
rect -12410 58150 -12090 58350
rect -12020 58150 -12000 58350
rect -16000 58140 -12000 58150
rect 96000 58350 100000 58360
rect 96000 58150 96020 58350
rect 96090 58150 96410 58350
rect 96480 58150 96520 58350
rect 96590 58150 96910 58350
rect 96980 58150 97020 58350
rect 97090 58150 97410 58350
rect 97480 58150 97520 58350
rect 97590 58150 97910 58350
rect 97980 58150 98020 58350
rect 98090 58150 98410 58350
rect 98480 58150 98520 58350
rect 98590 58150 98910 58350
rect 98980 58150 99020 58350
rect 99090 58150 99410 58350
rect 99480 58150 99520 58350
rect 99590 58150 99910 58350
rect 99980 58150 100000 58350
rect 96000 58140 100000 58150
rect -15860 58090 -15640 58140
rect -15860 58020 -15850 58090
rect -15650 58020 -15640 58090
rect -15860 57980 -15640 58020
rect -15860 57910 -15850 57980
rect -15650 57910 -15640 57980
rect -15860 57860 -15640 57910
rect -15360 58090 -15140 58140
rect -15360 58020 -15350 58090
rect -15150 58020 -15140 58090
rect -15360 57980 -15140 58020
rect -15360 57910 -15350 57980
rect -15150 57910 -15140 57980
rect -15360 57860 -15140 57910
rect -14860 58090 -14640 58140
rect -14860 58020 -14850 58090
rect -14650 58020 -14640 58090
rect -14860 57980 -14640 58020
rect -14860 57910 -14850 57980
rect -14650 57910 -14640 57980
rect -14860 57860 -14640 57910
rect -14360 58090 -14140 58140
rect -14360 58020 -14350 58090
rect -14150 58020 -14140 58090
rect -14360 57980 -14140 58020
rect -14360 57910 -14350 57980
rect -14150 57910 -14140 57980
rect -14360 57860 -14140 57910
rect -13860 58090 -13640 58140
rect -13860 58020 -13850 58090
rect -13650 58020 -13640 58090
rect -13860 57980 -13640 58020
rect -13860 57910 -13850 57980
rect -13650 57910 -13640 57980
rect -13860 57860 -13640 57910
rect -13360 58090 -13140 58140
rect -13360 58020 -13350 58090
rect -13150 58020 -13140 58090
rect -13360 57980 -13140 58020
rect -13360 57910 -13350 57980
rect -13150 57910 -13140 57980
rect -13360 57860 -13140 57910
rect -12860 58090 -12640 58140
rect -12860 58020 -12850 58090
rect -12650 58020 -12640 58090
rect -12860 57980 -12640 58020
rect -12860 57910 -12850 57980
rect -12650 57910 -12640 57980
rect -12860 57860 -12640 57910
rect -12360 58090 -12140 58140
rect -12360 58020 -12350 58090
rect -12150 58020 -12140 58090
rect -12360 57980 -12140 58020
rect -12360 57910 -12350 57980
rect -12150 57910 -12140 57980
rect -12360 57860 -12140 57910
rect 96140 58090 96360 58140
rect 96140 58020 96150 58090
rect 96350 58020 96360 58090
rect 96140 57980 96360 58020
rect 96140 57910 96150 57980
rect 96350 57910 96360 57980
rect 96140 57860 96360 57910
rect 96640 58090 96860 58140
rect 96640 58020 96650 58090
rect 96850 58020 96860 58090
rect 96640 57980 96860 58020
rect 96640 57910 96650 57980
rect 96850 57910 96860 57980
rect 96640 57860 96860 57910
rect 97140 58090 97360 58140
rect 97140 58020 97150 58090
rect 97350 58020 97360 58090
rect 97140 57980 97360 58020
rect 97140 57910 97150 57980
rect 97350 57910 97360 57980
rect 97140 57860 97360 57910
rect 97640 58090 97860 58140
rect 97640 58020 97650 58090
rect 97850 58020 97860 58090
rect 97640 57980 97860 58020
rect 97640 57910 97650 57980
rect 97850 57910 97860 57980
rect 97640 57860 97860 57910
rect 98140 58090 98360 58140
rect 98140 58020 98150 58090
rect 98350 58020 98360 58090
rect 98140 57980 98360 58020
rect 98140 57910 98150 57980
rect 98350 57910 98360 57980
rect 98140 57860 98360 57910
rect 98640 58090 98860 58140
rect 98640 58020 98650 58090
rect 98850 58020 98860 58090
rect 98640 57980 98860 58020
rect 98640 57910 98650 57980
rect 98850 57910 98860 57980
rect 98640 57860 98860 57910
rect 99140 58090 99360 58140
rect 99140 58020 99150 58090
rect 99350 58020 99360 58090
rect 99140 57980 99360 58020
rect 99140 57910 99150 57980
rect 99350 57910 99360 57980
rect 99140 57860 99360 57910
rect 99640 58090 99860 58140
rect 99640 58020 99650 58090
rect 99850 58020 99860 58090
rect 99640 57980 99860 58020
rect 99640 57910 99650 57980
rect 99850 57910 99860 57980
rect 99640 57860 99860 57910
rect -16000 57850 -12000 57860
rect -16000 57650 -15980 57850
rect -15910 57650 -15590 57850
rect -15520 57650 -15480 57850
rect -15410 57650 -15090 57850
rect -15020 57650 -14980 57850
rect -14910 57650 -14590 57850
rect -14520 57650 -14480 57850
rect -14410 57650 -14090 57850
rect -14020 57650 -13980 57850
rect -13910 57650 -13590 57850
rect -13520 57650 -13480 57850
rect -13410 57650 -13090 57850
rect -13020 57650 -12980 57850
rect -12910 57650 -12590 57850
rect -12520 57650 -12480 57850
rect -12410 57650 -12090 57850
rect -12020 57650 -12000 57850
rect -16000 57640 -12000 57650
rect 96000 57850 100000 57860
rect 96000 57650 96020 57850
rect 96090 57650 96410 57850
rect 96480 57650 96520 57850
rect 96590 57650 96910 57850
rect 96980 57650 97020 57850
rect 97090 57650 97410 57850
rect 97480 57650 97520 57850
rect 97590 57650 97910 57850
rect 97980 57650 98020 57850
rect 98090 57650 98410 57850
rect 98480 57650 98520 57850
rect 98590 57650 98910 57850
rect 98980 57650 99020 57850
rect 99090 57650 99410 57850
rect 99480 57650 99520 57850
rect 99590 57650 99910 57850
rect 99980 57650 100000 57850
rect 96000 57640 100000 57650
rect -15860 57590 -15640 57640
rect -15860 57520 -15850 57590
rect -15650 57520 -15640 57590
rect -15860 57480 -15640 57520
rect -15860 57410 -15850 57480
rect -15650 57410 -15640 57480
rect -15860 57360 -15640 57410
rect -15360 57590 -15140 57640
rect -15360 57520 -15350 57590
rect -15150 57520 -15140 57590
rect -15360 57480 -15140 57520
rect -15360 57410 -15350 57480
rect -15150 57410 -15140 57480
rect -15360 57360 -15140 57410
rect -14860 57590 -14640 57640
rect -14860 57520 -14850 57590
rect -14650 57520 -14640 57590
rect -14860 57480 -14640 57520
rect -14860 57410 -14850 57480
rect -14650 57410 -14640 57480
rect -14860 57360 -14640 57410
rect -14360 57590 -14140 57640
rect -14360 57520 -14350 57590
rect -14150 57520 -14140 57590
rect -14360 57480 -14140 57520
rect -14360 57410 -14350 57480
rect -14150 57410 -14140 57480
rect -14360 57360 -14140 57410
rect -13860 57590 -13640 57640
rect -13860 57520 -13850 57590
rect -13650 57520 -13640 57590
rect -13860 57480 -13640 57520
rect -13860 57410 -13850 57480
rect -13650 57410 -13640 57480
rect -13860 57360 -13640 57410
rect -13360 57590 -13140 57640
rect -13360 57520 -13350 57590
rect -13150 57520 -13140 57590
rect -13360 57480 -13140 57520
rect -13360 57410 -13350 57480
rect -13150 57410 -13140 57480
rect -13360 57360 -13140 57410
rect -12860 57590 -12640 57640
rect -12860 57520 -12850 57590
rect -12650 57520 -12640 57590
rect -12860 57480 -12640 57520
rect -12860 57410 -12850 57480
rect -12650 57410 -12640 57480
rect -12860 57360 -12640 57410
rect -12360 57590 -12140 57640
rect -12360 57520 -12350 57590
rect -12150 57520 -12140 57590
rect -12360 57480 -12140 57520
rect -12360 57410 -12350 57480
rect -12150 57410 -12140 57480
rect -12360 57360 -12140 57410
rect 96140 57590 96360 57640
rect 96140 57520 96150 57590
rect 96350 57520 96360 57590
rect 96140 57480 96360 57520
rect 96140 57410 96150 57480
rect 96350 57410 96360 57480
rect 96140 57360 96360 57410
rect 96640 57590 96860 57640
rect 96640 57520 96650 57590
rect 96850 57520 96860 57590
rect 96640 57480 96860 57520
rect 96640 57410 96650 57480
rect 96850 57410 96860 57480
rect 96640 57360 96860 57410
rect 97140 57590 97360 57640
rect 97140 57520 97150 57590
rect 97350 57520 97360 57590
rect 97140 57480 97360 57520
rect 97140 57410 97150 57480
rect 97350 57410 97360 57480
rect 97140 57360 97360 57410
rect 97640 57590 97860 57640
rect 97640 57520 97650 57590
rect 97850 57520 97860 57590
rect 97640 57480 97860 57520
rect 97640 57410 97650 57480
rect 97850 57410 97860 57480
rect 97640 57360 97860 57410
rect 98140 57590 98360 57640
rect 98140 57520 98150 57590
rect 98350 57520 98360 57590
rect 98140 57480 98360 57520
rect 98140 57410 98150 57480
rect 98350 57410 98360 57480
rect 98140 57360 98360 57410
rect 98640 57590 98860 57640
rect 98640 57520 98650 57590
rect 98850 57520 98860 57590
rect 98640 57480 98860 57520
rect 98640 57410 98650 57480
rect 98850 57410 98860 57480
rect 98640 57360 98860 57410
rect 99140 57590 99360 57640
rect 99140 57520 99150 57590
rect 99350 57520 99360 57590
rect 99140 57480 99360 57520
rect 99140 57410 99150 57480
rect 99350 57410 99360 57480
rect 99140 57360 99360 57410
rect 99640 57590 99860 57640
rect 99640 57520 99650 57590
rect 99850 57520 99860 57590
rect 99640 57480 99860 57520
rect 99640 57410 99650 57480
rect 99850 57410 99860 57480
rect 99640 57360 99860 57410
rect -16000 57350 -12000 57360
rect -16000 57150 -15980 57350
rect -15910 57150 -15590 57350
rect -15520 57150 -15480 57350
rect -15410 57150 -15090 57350
rect -15020 57150 -14980 57350
rect -14910 57150 -14590 57350
rect -14520 57150 -14480 57350
rect -14410 57150 -14090 57350
rect -14020 57150 -13980 57350
rect -13910 57150 -13590 57350
rect -13520 57150 -13480 57350
rect -13410 57150 -13090 57350
rect -13020 57150 -12980 57350
rect -12910 57150 -12590 57350
rect -12520 57150 -12480 57350
rect -12410 57150 -12090 57350
rect -12020 57150 -12000 57350
rect -16000 57140 -12000 57150
rect 96000 57350 100000 57360
rect 96000 57150 96020 57350
rect 96090 57150 96410 57350
rect 96480 57150 96520 57350
rect 96590 57150 96910 57350
rect 96980 57150 97020 57350
rect 97090 57150 97410 57350
rect 97480 57150 97520 57350
rect 97590 57150 97910 57350
rect 97980 57150 98020 57350
rect 98090 57150 98410 57350
rect 98480 57150 98520 57350
rect 98590 57150 98910 57350
rect 98980 57150 99020 57350
rect 99090 57150 99410 57350
rect 99480 57150 99520 57350
rect 99590 57150 99910 57350
rect 99980 57150 100000 57350
rect 96000 57140 100000 57150
rect -15860 57090 -15640 57140
rect -15860 57020 -15850 57090
rect -15650 57020 -15640 57090
rect -15860 56980 -15640 57020
rect -15860 56910 -15850 56980
rect -15650 56910 -15640 56980
rect -15860 56860 -15640 56910
rect -15360 57090 -15140 57140
rect -15360 57020 -15350 57090
rect -15150 57020 -15140 57090
rect -15360 56980 -15140 57020
rect -15360 56910 -15350 56980
rect -15150 56910 -15140 56980
rect -15360 56860 -15140 56910
rect -14860 57090 -14640 57140
rect -14860 57020 -14850 57090
rect -14650 57020 -14640 57090
rect -14860 56980 -14640 57020
rect -14860 56910 -14850 56980
rect -14650 56910 -14640 56980
rect -14860 56860 -14640 56910
rect -14360 57090 -14140 57140
rect -14360 57020 -14350 57090
rect -14150 57020 -14140 57090
rect -14360 56980 -14140 57020
rect -14360 56910 -14350 56980
rect -14150 56910 -14140 56980
rect -14360 56860 -14140 56910
rect -13860 57090 -13640 57140
rect -13860 57020 -13850 57090
rect -13650 57020 -13640 57090
rect -13860 56980 -13640 57020
rect -13860 56910 -13850 56980
rect -13650 56910 -13640 56980
rect -13860 56860 -13640 56910
rect -13360 57090 -13140 57140
rect -13360 57020 -13350 57090
rect -13150 57020 -13140 57090
rect -13360 56980 -13140 57020
rect -13360 56910 -13350 56980
rect -13150 56910 -13140 56980
rect -13360 56860 -13140 56910
rect -12860 57090 -12640 57140
rect -12860 57020 -12850 57090
rect -12650 57020 -12640 57090
rect -12860 56980 -12640 57020
rect -12860 56910 -12850 56980
rect -12650 56910 -12640 56980
rect -12860 56860 -12640 56910
rect -12360 57090 -12140 57140
rect -12360 57020 -12350 57090
rect -12150 57020 -12140 57090
rect -12360 56980 -12140 57020
rect -12360 56910 -12350 56980
rect -12150 56910 -12140 56980
rect -12360 56860 -12140 56910
rect 96140 57090 96360 57140
rect 96140 57020 96150 57090
rect 96350 57020 96360 57090
rect 96140 56980 96360 57020
rect 96140 56910 96150 56980
rect 96350 56910 96360 56980
rect 96140 56860 96360 56910
rect 96640 57090 96860 57140
rect 96640 57020 96650 57090
rect 96850 57020 96860 57090
rect 96640 56980 96860 57020
rect 96640 56910 96650 56980
rect 96850 56910 96860 56980
rect 96640 56860 96860 56910
rect 97140 57090 97360 57140
rect 97140 57020 97150 57090
rect 97350 57020 97360 57090
rect 97140 56980 97360 57020
rect 97140 56910 97150 56980
rect 97350 56910 97360 56980
rect 97140 56860 97360 56910
rect 97640 57090 97860 57140
rect 97640 57020 97650 57090
rect 97850 57020 97860 57090
rect 97640 56980 97860 57020
rect 97640 56910 97650 56980
rect 97850 56910 97860 56980
rect 97640 56860 97860 56910
rect 98140 57090 98360 57140
rect 98140 57020 98150 57090
rect 98350 57020 98360 57090
rect 98140 56980 98360 57020
rect 98140 56910 98150 56980
rect 98350 56910 98360 56980
rect 98140 56860 98360 56910
rect 98640 57090 98860 57140
rect 98640 57020 98650 57090
rect 98850 57020 98860 57090
rect 98640 56980 98860 57020
rect 98640 56910 98650 56980
rect 98850 56910 98860 56980
rect 98640 56860 98860 56910
rect 99140 57090 99360 57140
rect 99140 57020 99150 57090
rect 99350 57020 99360 57090
rect 99140 56980 99360 57020
rect 99140 56910 99150 56980
rect 99350 56910 99360 56980
rect 99140 56860 99360 56910
rect 99640 57090 99860 57140
rect 99640 57020 99650 57090
rect 99850 57020 99860 57090
rect 99640 56980 99860 57020
rect 99640 56910 99650 56980
rect 99850 56910 99860 56980
rect 99640 56860 99860 56910
rect -16000 56850 -12000 56860
rect -16000 56650 -15980 56850
rect -15910 56650 -15590 56850
rect -15520 56650 -15480 56850
rect -15410 56650 -15090 56850
rect -15020 56650 -14980 56850
rect -14910 56650 -14590 56850
rect -14520 56650 -14480 56850
rect -14410 56650 -14090 56850
rect -14020 56650 -13980 56850
rect -13910 56650 -13590 56850
rect -13520 56650 -13480 56850
rect -13410 56650 -13090 56850
rect -13020 56650 -12980 56850
rect -12910 56650 -12590 56850
rect -12520 56650 -12480 56850
rect -12410 56650 -12090 56850
rect -12020 56650 -12000 56850
rect -16000 56640 -12000 56650
rect 96000 56850 100000 56860
rect 96000 56650 96020 56850
rect 96090 56650 96410 56850
rect 96480 56650 96520 56850
rect 96590 56650 96910 56850
rect 96980 56650 97020 56850
rect 97090 56650 97410 56850
rect 97480 56650 97520 56850
rect 97590 56650 97910 56850
rect 97980 56650 98020 56850
rect 98090 56650 98410 56850
rect 98480 56650 98520 56850
rect 98590 56650 98910 56850
rect 98980 56650 99020 56850
rect 99090 56650 99410 56850
rect 99480 56650 99520 56850
rect 99590 56650 99910 56850
rect 99980 56650 100000 56850
rect 96000 56640 100000 56650
rect -15860 56590 -15640 56640
rect -15860 56520 -15850 56590
rect -15650 56520 -15640 56590
rect -15860 56480 -15640 56520
rect -15860 56410 -15850 56480
rect -15650 56410 -15640 56480
rect -15860 56360 -15640 56410
rect -15360 56590 -15140 56640
rect -15360 56520 -15350 56590
rect -15150 56520 -15140 56590
rect -15360 56480 -15140 56520
rect -15360 56410 -15350 56480
rect -15150 56410 -15140 56480
rect -15360 56360 -15140 56410
rect -14860 56590 -14640 56640
rect -14860 56520 -14850 56590
rect -14650 56520 -14640 56590
rect -14860 56480 -14640 56520
rect -14860 56410 -14850 56480
rect -14650 56410 -14640 56480
rect -14860 56360 -14640 56410
rect -14360 56590 -14140 56640
rect -14360 56520 -14350 56590
rect -14150 56520 -14140 56590
rect -14360 56480 -14140 56520
rect -14360 56410 -14350 56480
rect -14150 56410 -14140 56480
rect -14360 56360 -14140 56410
rect -13860 56590 -13640 56640
rect -13860 56520 -13850 56590
rect -13650 56520 -13640 56590
rect -13860 56480 -13640 56520
rect -13860 56410 -13850 56480
rect -13650 56410 -13640 56480
rect -13860 56360 -13640 56410
rect -13360 56590 -13140 56640
rect -13360 56520 -13350 56590
rect -13150 56520 -13140 56590
rect -13360 56480 -13140 56520
rect -13360 56410 -13350 56480
rect -13150 56410 -13140 56480
rect -13360 56360 -13140 56410
rect -12860 56590 -12640 56640
rect -12860 56520 -12850 56590
rect -12650 56520 -12640 56590
rect -12860 56480 -12640 56520
rect -12860 56410 -12850 56480
rect -12650 56410 -12640 56480
rect -12860 56360 -12640 56410
rect -12360 56590 -12140 56640
rect -12360 56520 -12350 56590
rect -12150 56520 -12140 56590
rect -12360 56480 -12140 56520
rect -12360 56410 -12350 56480
rect -12150 56410 -12140 56480
rect -12360 56360 -12140 56410
rect 96140 56590 96360 56640
rect 96140 56520 96150 56590
rect 96350 56520 96360 56590
rect 96140 56480 96360 56520
rect 96140 56410 96150 56480
rect 96350 56410 96360 56480
rect 96140 56360 96360 56410
rect 96640 56590 96860 56640
rect 96640 56520 96650 56590
rect 96850 56520 96860 56590
rect 96640 56480 96860 56520
rect 96640 56410 96650 56480
rect 96850 56410 96860 56480
rect 96640 56360 96860 56410
rect 97140 56590 97360 56640
rect 97140 56520 97150 56590
rect 97350 56520 97360 56590
rect 97140 56480 97360 56520
rect 97140 56410 97150 56480
rect 97350 56410 97360 56480
rect 97140 56360 97360 56410
rect 97640 56590 97860 56640
rect 97640 56520 97650 56590
rect 97850 56520 97860 56590
rect 97640 56480 97860 56520
rect 97640 56410 97650 56480
rect 97850 56410 97860 56480
rect 97640 56360 97860 56410
rect 98140 56590 98360 56640
rect 98140 56520 98150 56590
rect 98350 56520 98360 56590
rect 98140 56480 98360 56520
rect 98140 56410 98150 56480
rect 98350 56410 98360 56480
rect 98140 56360 98360 56410
rect 98640 56590 98860 56640
rect 98640 56520 98650 56590
rect 98850 56520 98860 56590
rect 98640 56480 98860 56520
rect 98640 56410 98650 56480
rect 98850 56410 98860 56480
rect 98640 56360 98860 56410
rect 99140 56590 99360 56640
rect 99140 56520 99150 56590
rect 99350 56520 99360 56590
rect 99140 56480 99360 56520
rect 99140 56410 99150 56480
rect 99350 56410 99360 56480
rect 99140 56360 99360 56410
rect 99640 56590 99860 56640
rect 99640 56520 99650 56590
rect 99850 56520 99860 56590
rect 99640 56480 99860 56520
rect 99640 56410 99650 56480
rect 99850 56410 99860 56480
rect 99640 56360 99860 56410
rect -16000 56350 -12000 56360
rect -16000 56150 -15980 56350
rect -15910 56150 -15590 56350
rect -15520 56150 -15480 56350
rect -15410 56150 -15090 56350
rect -15020 56150 -14980 56350
rect -14910 56150 -14590 56350
rect -14520 56150 -14480 56350
rect -14410 56150 -14090 56350
rect -14020 56150 -13980 56350
rect -13910 56150 -13590 56350
rect -13520 56150 -13480 56350
rect -13410 56150 -13090 56350
rect -13020 56150 -12980 56350
rect -12910 56150 -12590 56350
rect -12520 56150 -12480 56350
rect -12410 56150 -12090 56350
rect -12020 56150 -12000 56350
rect -16000 56140 -12000 56150
rect 96000 56350 100000 56360
rect 96000 56150 96020 56350
rect 96090 56150 96410 56350
rect 96480 56150 96520 56350
rect 96590 56150 96910 56350
rect 96980 56150 97020 56350
rect 97090 56150 97410 56350
rect 97480 56150 97520 56350
rect 97590 56150 97910 56350
rect 97980 56150 98020 56350
rect 98090 56150 98410 56350
rect 98480 56150 98520 56350
rect 98590 56150 98910 56350
rect 98980 56150 99020 56350
rect 99090 56150 99410 56350
rect 99480 56150 99520 56350
rect 99590 56150 99910 56350
rect 99980 56150 100000 56350
rect 96000 56140 100000 56150
rect -15860 56090 -15640 56140
rect -15860 56020 -15850 56090
rect -15650 56020 -15640 56090
rect -15860 55980 -15640 56020
rect -15860 55910 -15850 55980
rect -15650 55910 -15640 55980
rect -15860 55860 -15640 55910
rect -15360 56090 -15140 56140
rect -15360 56020 -15350 56090
rect -15150 56020 -15140 56090
rect -15360 55980 -15140 56020
rect -15360 55910 -15350 55980
rect -15150 55910 -15140 55980
rect -15360 55860 -15140 55910
rect -14860 56090 -14640 56140
rect -14860 56020 -14850 56090
rect -14650 56020 -14640 56090
rect -14860 55980 -14640 56020
rect -14860 55910 -14850 55980
rect -14650 55910 -14640 55980
rect -14860 55860 -14640 55910
rect -14360 56090 -14140 56140
rect -14360 56020 -14350 56090
rect -14150 56020 -14140 56090
rect -14360 55980 -14140 56020
rect -14360 55910 -14350 55980
rect -14150 55910 -14140 55980
rect -14360 55860 -14140 55910
rect -13860 56090 -13640 56140
rect -13860 56020 -13850 56090
rect -13650 56020 -13640 56090
rect -13860 55980 -13640 56020
rect -13860 55910 -13850 55980
rect -13650 55910 -13640 55980
rect -13860 55860 -13640 55910
rect -13360 56090 -13140 56140
rect -13360 56020 -13350 56090
rect -13150 56020 -13140 56090
rect -13360 55980 -13140 56020
rect -13360 55910 -13350 55980
rect -13150 55910 -13140 55980
rect -13360 55860 -13140 55910
rect -12860 56090 -12640 56140
rect -12860 56020 -12850 56090
rect -12650 56020 -12640 56090
rect -12860 55980 -12640 56020
rect -12860 55910 -12850 55980
rect -12650 55910 -12640 55980
rect -12860 55860 -12640 55910
rect -12360 56090 -12140 56140
rect -12360 56020 -12350 56090
rect -12150 56020 -12140 56090
rect -12360 55980 -12140 56020
rect -12360 55910 -12350 55980
rect -12150 55910 -12140 55980
rect -12360 55860 -12140 55910
rect 96140 56090 96360 56140
rect 96140 56020 96150 56090
rect 96350 56020 96360 56090
rect 96140 55980 96360 56020
rect 96140 55910 96150 55980
rect 96350 55910 96360 55980
rect 96140 55860 96360 55910
rect 96640 56090 96860 56140
rect 96640 56020 96650 56090
rect 96850 56020 96860 56090
rect 96640 55980 96860 56020
rect 96640 55910 96650 55980
rect 96850 55910 96860 55980
rect 96640 55860 96860 55910
rect 97140 56090 97360 56140
rect 97140 56020 97150 56090
rect 97350 56020 97360 56090
rect 97140 55980 97360 56020
rect 97140 55910 97150 55980
rect 97350 55910 97360 55980
rect 97140 55860 97360 55910
rect 97640 56090 97860 56140
rect 97640 56020 97650 56090
rect 97850 56020 97860 56090
rect 97640 55980 97860 56020
rect 97640 55910 97650 55980
rect 97850 55910 97860 55980
rect 97640 55860 97860 55910
rect 98140 56090 98360 56140
rect 98140 56020 98150 56090
rect 98350 56020 98360 56090
rect 98140 55980 98360 56020
rect 98140 55910 98150 55980
rect 98350 55910 98360 55980
rect 98140 55860 98360 55910
rect 98640 56090 98860 56140
rect 98640 56020 98650 56090
rect 98850 56020 98860 56090
rect 98640 55980 98860 56020
rect 98640 55910 98650 55980
rect 98850 55910 98860 55980
rect 98640 55860 98860 55910
rect 99140 56090 99360 56140
rect 99140 56020 99150 56090
rect 99350 56020 99360 56090
rect 99140 55980 99360 56020
rect 99140 55910 99150 55980
rect 99350 55910 99360 55980
rect 99140 55860 99360 55910
rect 99640 56090 99860 56140
rect 99640 56020 99650 56090
rect 99850 56020 99860 56090
rect 99640 55980 99860 56020
rect 99640 55910 99650 55980
rect 99850 55910 99860 55980
rect 99640 55860 99860 55910
rect -16000 55850 -12000 55860
rect -16000 55650 -15980 55850
rect -15910 55650 -15590 55850
rect -15520 55650 -15480 55850
rect -15410 55650 -15090 55850
rect -15020 55650 -14980 55850
rect -14910 55650 -14590 55850
rect -14520 55650 -14480 55850
rect -14410 55650 -14090 55850
rect -14020 55650 -13980 55850
rect -13910 55650 -13590 55850
rect -13520 55650 -13480 55850
rect -13410 55650 -13090 55850
rect -13020 55650 -12980 55850
rect -12910 55650 -12590 55850
rect -12520 55650 -12480 55850
rect -12410 55650 -12090 55850
rect -12020 55650 -12000 55850
rect -16000 55640 -12000 55650
rect 96000 55850 100000 55860
rect 96000 55650 96020 55850
rect 96090 55650 96410 55850
rect 96480 55650 96520 55850
rect 96590 55650 96910 55850
rect 96980 55650 97020 55850
rect 97090 55650 97410 55850
rect 97480 55650 97520 55850
rect 97590 55650 97910 55850
rect 97980 55650 98020 55850
rect 98090 55650 98410 55850
rect 98480 55650 98520 55850
rect 98590 55650 98910 55850
rect 98980 55650 99020 55850
rect 99090 55650 99410 55850
rect 99480 55650 99520 55850
rect 99590 55650 99910 55850
rect 99980 55650 100000 55850
rect 96000 55640 100000 55650
rect -15860 55590 -15640 55640
rect -15860 55520 -15850 55590
rect -15650 55520 -15640 55590
rect -15860 55480 -15640 55520
rect -15860 55410 -15850 55480
rect -15650 55410 -15640 55480
rect -15860 55360 -15640 55410
rect -15360 55590 -15140 55640
rect -15360 55520 -15350 55590
rect -15150 55520 -15140 55590
rect -15360 55480 -15140 55520
rect -15360 55410 -15350 55480
rect -15150 55410 -15140 55480
rect -15360 55360 -15140 55410
rect -14860 55590 -14640 55640
rect -14860 55520 -14850 55590
rect -14650 55520 -14640 55590
rect -14860 55480 -14640 55520
rect -14860 55410 -14850 55480
rect -14650 55410 -14640 55480
rect -14860 55360 -14640 55410
rect -14360 55590 -14140 55640
rect -14360 55520 -14350 55590
rect -14150 55520 -14140 55590
rect -14360 55480 -14140 55520
rect -14360 55410 -14350 55480
rect -14150 55410 -14140 55480
rect -14360 55360 -14140 55410
rect -13860 55590 -13640 55640
rect -13860 55520 -13850 55590
rect -13650 55520 -13640 55590
rect -13860 55480 -13640 55520
rect -13860 55410 -13850 55480
rect -13650 55410 -13640 55480
rect -13860 55360 -13640 55410
rect -13360 55590 -13140 55640
rect -13360 55520 -13350 55590
rect -13150 55520 -13140 55590
rect -13360 55480 -13140 55520
rect -13360 55410 -13350 55480
rect -13150 55410 -13140 55480
rect -13360 55360 -13140 55410
rect -12860 55590 -12640 55640
rect -12860 55520 -12850 55590
rect -12650 55520 -12640 55590
rect -12860 55480 -12640 55520
rect -12860 55410 -12850 55480
rect -12650 55410 -12640 55480
rect -12860 55360 -12640 55410
rect -12360 55590 -12140 55640
rect -12360 55520 -12350 55590
rect -12150 55520 -12140 55590
rect -12360 55480 -12140 55520
rect -12360 55410 -12350 55480
rect -12150 55410 -12140 55480
rect -12360 55360 -12140 55410
rect 96140 55590 96360 55640
rect 96140 55520 96150 55590
rect 96350 55520 96360 55590
rect 96140 55480 96360 55520
rect 96140 55410 96150 55480
rect 96350 55410 96360 55480
rect 96140 55360 96360 55410
rect 96640 55590 96860 55640
rect 96640 55520 96650 55590
rect 96850 55520 96860 55590
rect 96640 55480 96860 55520
rect 96640 55410 96650 55480
rect 96850 55410 96860 55480
rect 96640 55360 96860 55410
rect 97140 55590 97360 55640
rect 97140 55520 97150 55590
rect 97350 55520 97360 55590
rect 97140 55480 97360 55520
rect 97140 55410 97150 55480
rect 97350 55410 97360 55480
rect 97140 55360 97360 55410
rect 97640 55590 97860 55640
rect 97640 55520 97650 55590
rect 97850 55520 97860 55590
rect 97640 55480 97860 55520
rect 97640 55410 97650 55480
rect 97850 55410 97860 55480
rect 97640 55360 97860 55410
rect 98140 55590 98360 55640
rect 98140 55520 98150 55590
rect 98350 55520 98360 55590
rect 98140 55480 98360 55520
rect 98140 55410 98150 55480
rect 98350 55410 98360 55480
rect 98140 55360 98360 55410
rect 98640 55590 98860 55640
rect 98640 55520 98650 55590
rect 98850 55520 98860 55590
rect 98640 55480 98860 55520
rect 98640 55410 98650 55480
rect 98850 55410 98860 55480
rect 98640 55360 98860 55410
rect 99140 55590 99360 55640
rect 99140 55520 99150 55590
rect 99350 55520 99360 55590
rect 99140 55480 99360 55520
rect 99140 55410 99150 55480
rect 99350 55410 99360 55480
rect 99140 55360 99360 55410
rect 99640 55590 99860 55640
rect 99640 55520 99650 55590
rect 99850 55520 99860 55590
rect 99640 55480 99860 55520
rect 99640 55410 99650 55480
rect 99850 55410 99860 55480
rect 99640 55360 99860 55410
rect -16000 55350 -12000 55360
rect -16000 55150 -15980 55350
rect -15910 55150 -15590 55350
rect -15520 55150 -15480 55350
rect -15410 55150 -15090 55350
rect -15020 55150 -14980 55350
rect -14910 55150 -14590 55350
rect -14520 55150 -14480 55350
rect -14410 55150 -14090 55350
rect -14020 55150 -13980 55350
rect -13910 55150 -13590 55350
rect -13520 55150 -13480 55350
rect -13410 55150 -13090 55350
rect -13020 55150 -12980 55350
rect -12910 55150 -12590 55350
rect -12520 55150 -12480 55350
rect -12410 55150 -12090 55350
rect -12020 55150 -12000 55350
rect -16000 55140 -12000 55150
rect 96000 55350 100000 55360
rect 96000 55150 96020 55350
rect 96090 55150 96410 55350
rect 96480 55150 96520 55350
rect 96590 55150 96910 55350
rect 96980 55150 97020 55350
rect 97090 55150 97410 55350
rect 97480 55150 97520 55350
rect 97590 55150 97910 55350
rect 97980 55150 98020 55350
rect 98090 55150 98410 55350
rect 98480 55150 98520 55350
rect 98590 55150 98910 55350
rect 98980 55150 99020 55350
rect 99090 55150 99410 55350
rect 99480 55150 99520 55350
rect 99590 55150 99910 55350
rect 99980 55150 100000 55350
rect 96000 55140 100000 55150
rect -15860 55090 -15640 55140
rect -15860 55020 -15850 55090
rect -15650 55020 -15640 55090
rect -15860 54980 -15640 55020
rect -15860 54910 -15850 54980
rect -15650 54910 -15640 54980
rect -15860 54860 -15640 54910
rect -15360 55090 -15140 55140
rect -15360 55020 -15350 55090
rect -15150 55020 -15140 55090
rect -15360 54980 -15140 55020
rect -15360 54910 -15350 54980
rect -15150 54910 -15140 54980
rect -15360 54860 -15140 54910
rect -14860 55090 -14640 55140
rect -14860 55020 -14850 55090
rect -14650 55020 -14640 55090
rect -14860 54980 -14640 55020
rect -14860 54910 -14850 54980
rect -14650 54910 -14640 54980
rect -14860 54860 -14640 54910
rect -14360 55090 -14140 55140
rect -14360 55020 -14350 55090
rect -14150 55020 -14140 55090
rect -14360 54980 -14140 55020
rect -14360 54910 -14350 54980
rect -14150 54910 -14140 54980
rect -14360 54860 -14140 54910
rect -13860 55090 -13640 55140
rect -13860 55020 -13850 55090
rect -13650 55020 -13640 55090
rect -13860 54980 -13640 55020
rect -13860 54910 -13850 54980
rect -13650 54910 -13640 54980
rect -13860 54860 -13640 54910
rect -13360 55090 -13140 55140
rect -13360 55020 -13350 55090
rect -13150 55020 -13140 55090
rect -13360 54980 -13140 55020
rect -13360 54910 -13350 54980
rect -13150 54910 -13140 54980
rect -13360 54860 -13140 54910
rect -12860 55090 -12640 55140
rect -12860 55020 -12850 55090
rect -12650 55020 -12640 55090
rect -12860 54980 -12640 55020
rect -12860 54910 -12850 54980
rect -12650 54910 -12640 54980
rect -12860 54860 -12640 54910
rect -12360 55090 -12140 55140
rect -12360 55020 -12350 55090
rect -12150 55020 -12140 55090
rect -12360 54980 -12140 55020
rect -12360 54910 -12350 54980
rect -12150 54910 -12140 54980
rect -12360 54860 -12140 54910
rect 96140 55090 96360 55140
rect 96140 55020 96150 55090
rect 96350 55020 96360 55090
rect 96140 54980 96360 55020
rect 96140 54910 96150 54980
rect 96350 54910 96360 54980
rect 96140 54860 96360 54910
rect 96640 55090 96860 55140
rect 96640 55020 96650 55090
rect 96850 55020 96860 55090
rect 96640 54980 96860 55020
rect 96640 54910 96650 54980
rect 96850 54910 96860 54980
rect 96640 54860 96860 54910
rect 97140 55090 97360 55140
rect 97140 55020 97150 55090
rect 97350 55020 97360 55090
rect 97140 54980 97360 55020
rect 97140 54910 97150 54980
rect 97350 54910 97360 54980
rect 97140 54860 97360 54910
rect 97640 55090 97860 55140
rect 97640 55020 97650 55090
rect 97850 55020 97860 55090
rect 97640 54980 97860 55020
rect 97640 54910 97650 54980
rect 97850 54910 97860 54980
rect 97640 54860 97860 54910
rect 98140 55090 98360 55140
rect 98140 55020 98150 55090
rect 98350 55020 98360 55090
rect 98140 54980 98360 55020
rect 98140 54910 98150 54980
rect 98350 54910 98360 54980
rect 98140 54860 98360 54910
rect 98640 55090 98860 55140
rect 98640 55020 98650 55090
rect 98850 55020 98860 55090
rect 98640 54980 98860 55020
rect 98640 54910 98650 54980
rect 98850 54910 98860 54980
rect 98640 54860 98860 54910
rect 99140 55090 99360 55140
rect 99140 55020 99150 55090
rect 99350 55020 99360 55090
rect 99140 54980 99360 55020
rect 99140 54910 99150 54980
rect 99350 54910 99360 54980
rect 99140 54860 99360 54910
rect 99640 55090 99860 55140
rect 99640 55020 99650 55090
rect 99850 55020 99860 55090
rect 99640 54980 99860 55020
rect 99640 54910 99650 54980
rect 99850 54910 99860 54980
rect 99640 54860 99860 54910
rect -16000 54850 -12000 54860
rect -16000 54650 -15980 54850
rect -15910 54650 -15590 54850
rect -15520 54650 -15480 54850
rect -15410 54650 -15090 54850
rect -15020 54650 -14980 54850
rect -14910 54650 -14590 54850
rect -14520 54650 -14480 54850
rect -14410 54650 -14090 54850
rect -14020 54650 -13980 54850
rect -13910 54650 -13590 54850
rect -13520 54650 -13480 54850
rect -13410 54650 -13090 54850
rect -13020 54650 -12980 54850
rect -12910 54650 -12590 54850
rect -12520 54650 -12480 54850
rect -12410 54650 -12090 54850
rect -12020 54650 -12000 54850
rect -16000 54640 -12000 54650
rect 96000 54850 100000 54860
rect 96000 54650 96020 54850
rect 96090 54650 96410 54850
rect 96480 54650 96520 54850
rect 96590 54650 96910 54850
rect 96980 54650 97020 54850
rect 97090 54650 97410 54850
rect 97480 54650 97520 54850
rect 97590 54650 97910 54850
rect 97980 54650 98020 54850
rect 98090 54650 98410 54850
rect 98480 54650 98520 54850
rect 98590 54650 98910 54850
rect 98980 54650 99020 54850
rect 99090 54650 99410 54850
rect 99480 54650 99520 54850
rect 99590 54650 99910 54850
rect 99980 54650 100000 54850
rect 96000 54640 100000 54650
rect -15860 54590 -15640 54640
rect -15860 54520 -15850 54590
rect -15650 54520 -15640 54590
rect -15860 54480 -15640 54520
rect -15860 54410 -15850 54480
rect -15650 54410 -15640 54480
rect -15860 54360 -15640 54410
rect -15360 54590 -15140 54640
rect -15360 54520 -15350 54590
rect -15150 54520 -15140 54590
rect -15360 54480 -15140 54520
rect -15360 54410 -15350 54480
rect -15150 54410 -15140 54480
rect -15360 54360 -15140 54410
rect -14860 54590 -14640 54640
rect -14860 54520 -14850 54590
rect -14650 54520 -14640 54590
rect -14860 54480 -14640 54520
rect -14860 54410 -14850 54480
rect -14650 54410 -14640 54480
rect -14860 54360 -14640 54410
rect -14360 54590 -14140 54640
rect -14360 54520 -14350 54590
rect -14150 54520 -14140 54590
rect -14360 54480 -14140 54520
rect -14360 54410 -14350 54480
rect -14150 54410 -14140 54480
rect -14360 54360 -14140 54410
rect -13860 54590 -13640 54640
rect -13860 54520 -13850 54590
rect -13650 54520 -13640 54590
rect -13860 54480 -13640 54520
rect -13860 54410 -13850 54480
rect -13650 54410 -13640 54480
rect -13860 54360 -13640 54410
rect -13360 54590 -13140 54640
rect -13360 54520 -13350 54590
rect -13150 54520 -13140 54590
rect -13360 54480 -13140 54520
rect -13360 54410 -13350 54480
rect -13150 54410 -13140 54480
rect -13360 54360 -13140 54410
rect -12860 54590 -12640 54640
rect -12860 54520 -12850 54590
rect -12650 54520 -12640 54590
rect -12860 54480 -12640 54520
rect -12860 54410 -12850 54480
rect -12650 54410 -12640 54480
rect -12860 54360 -12640 54410
rect -12360 54590 -12140 54640
rect -12360 54520 -12350 54590
rect -12150 54520 -12140 54590
rect -12360 54480 -12140 54520
rect -12360 54410 -12350 54480
rect -12150 54410 -12140 54480
rect -12360 54360 -12140 54410
rect 96140 54590 96360 54640
rect 96140 54520 96150 54590
rect 96350 54520 96360 54590
rect 96140 54480 96360 54520
rect 96140 54410 96150 54480
rect 96350 54410 96360 54480
rect 96140 54360 96360 54410
rect 96640 54590 96860 54640
rect 96640 54520 96650 54590
rect 96850 54520 96860 54590
rect 96640 54480 96860 54520
rect 96640 54410 96650 54480
rect 96850 54410 96860 54480
rect 96640 54360 96860 54410
rect 97140 54590 97360 54640
rect 97140 54520 97150 54590
rect 97350 54520 97360 54590
rect 97140 54480 97360 54520
rect 97140 54410 97150 54480
rect 97350 54410 97360 54480
rect 97140 54360 97360 54410
rect 97640 54590 97860 54640
rect 97640 54520 97650 54590
rect 97850 54520 97860 54590
rect 97640 54480 97860 54520
rect 97640 54410 97650 54480
rect 97850 54410 97860 54480
rect 97640 54360 97860 54410
rect 98140 54590 98360 54640
rect 98140 54520 98150 54590
rect 98350 54520 98360 54590
rect 98140 54480 98360 54520
rect 98140 54410 98150 54480
rect 98350 54410 98360 54480
rect 98140 54360 98360 54410
rect 98640 54590 98860 54640
rect 98640 54520 98650 54590
rect 98850 54520 98860 54590
rect 98640 54480 98860 54520
rect 98640 54410 98650 54480
rect 98850 54410 98860 54480
rect 98640 54360 98860 54410
rect 99140 54590 99360 54640
rect 99140 54520 99150 54590
rect 99350 54520 99360 54590
rect 99140 54480 99360 54520
rect 99140 54410 99150 54480
rect 99350 54410 99360 54480
rect 99140 54360 99360 54410
rect 99640 54590 99860 54640
rect 99640 54520 99650 54590
rect 99850 54520 99860 54590
rect 99640 54480 99860 54520
rect 99640 54410 99650 54480
rect 99850 54410 99860 54480
rect 99640 54360 99860 54410
rect -16000 54350 -12000 54360
rect -16000 54150 -15980 54350
rect -15910 54150 -15590 54350
rect -15520 54150 -15480 54350
rect -15410 54150 -15090 54350
rect -15020 54150 -14980 54350
rect -14910 54150 -14590 54350
rect -14520 54150 -14480 54350
rect -14410 54150 -14090 54350
rect -14020 54150 -13980 54350
rect -13910 54150 -13590 54350
rect -13520 54150 -13480 54350
rect -13410 54150 -13090 54350
rect -13020 54150 -12980 54350
rect -12910 54150 -12590 54350
rect -12520 54150 -12480 54350
rect -12410 54150 -12090 54350
rect -12020 54150 -12000 54350
rect -16000 54140 -12000 54150
rect 96000 54350 100000 54360
rect 96000 54150 96020 54350
rect 96090 54150 96410 54350
rect 96480 54150 96520 54350
rect 96590 54150 96910 54350
rect 96980 54150 97020 54350
rect 97090 54150 97410 54350
rect 97480 54150 97520 54350
rect 97590 54150 97910 54350
rect 97980 54150 98020 54350
rect 98090 54150 98410 54350
rect 98480 54150 98520 54350
rect 98590 54150 98910 54350
rect 98980 54150 99020 54350
rect 99090 54150 99410 54350
rect 99480 54150 99520 54350
rect 99590 54150 99910 54350
rect 99980 54150 100000 54350
rect 96000 54140 100000 54150
rect -15860 54090 -15640 54140
rect -15860 54020 -15850 54090
rect -15650 54020 -15640 54090
rect -15860 53980 -15640 54020
rect -15860 53910 -15850 53980
rect -15650 53910 -15640 53980
rect -15860 53860 -15640 53910
rect -15360 54090 -15140 54140
rect -15360 54020 -15350 54090
rect -15150 54020 -15140 54090
rect -15360 53980 -15140 54020
rect -15360 53910 -15350 53980
rect -15150 53910 -15140 53980
rect -15360 53860 -15140 53910
rect -14860 54090 -14640 54140
rect -14860 54020 -14850 54090
rect -14650 54020 -14640 54090
rect -14860 53980 -14640 54020
rect -14860 53910 -14850 53980
rect -14650 53910 -14640 53980
rect -14860 53860 -14640 53910
rect -14360 54090 -14140 54140
rect -14360 54020 -14350 54090
rect -14150 54020 -14140 54090
rect -14360 53980 -14140 54020
rect -14360 53910 -14350 53980
rect -14150 53910 -14140 53980
rect -14360 53860 -14140 53910
rect -13860 54090 -13640 54140
rect -13860 54020 -13850 54090
rect -13650 54020 -13640 54090
rect -13860 53980 -13640 54020
rect -13860 53910 -13850 53980
rect -13650 53910 -13640 53980
rect -13860 53860 -13640 53910
rect -13360 54090 -13140 54140
rect -13360 54020 -13350 54090
rect -13150 54020 -13140 54090
rect -13360 53980 -13140 54020
rect -13360 53910 -13350 53980
rect -13150 53910 -13140 53980
rect -13360 53860 -13140 53910
rect -12860 54090 -12640 54140
rect -12860 54020 -12850 54090
rect -12650 54020 -12640 54090
rect -12860 53980 -12640 54020
rect -12860 53910 -12850 53980
rect -12650 53910 -12640 53980
rect -12860 53860 -12640 53910
rect -12360 54090 -12140 54140
rect -12360 54020 -12350 54090
rect -12150 54020 -12140 54090
rect -12360 53980 -12140 54020
rect -12360 53910 -12350 53980
rect -12150 53910 -12140 53980
rect -12360 53860 -12140 53910
rect 96140 54090 96360 54140
rect 96140 54020 96150 54090
rect 96350 54020 96360 54090
rect 96140 53980 96360 54020
rect 96140 53910 96150 53980
rect 96350 53910 96360 53980
rect 96140 53860 96360 53910
rect 96640 54090 96860 54140
rect 96640 54020 96650 54090
rect 96850 54020 96860 54090
rect 96640 53980 96860 54020
rect 96640 53910 96650 53980
rect 96850 53910 96860 53980
rect 96640 53860 96860 53910
rect 97140 54090 97360 54140
rect 97140 54020 97150 54090
rect 97350 54020 97360 54090
rect 97140 53980 97360 54020
rect 97140 53910 97150 53980
rect 97350 53910 97360 53980
rect 97140 53860 97360 53910
rect 97640 54090 97860 54140
rect 97640 54020 97650 54090
rect 97850 54020 97860 54090
rect 97640 53980 97860 54020
rect 97640 53910 97650 53980
rect 97850 53910 97860 53980
rect 97640 53860 97860 53910
rect 98140 54090 98360 54140
rect 98140 54020 98150 54090
rect 98350 54020 98360 54090
rect 98140 53980 98360 54020
rect 98140 53910 98150 53980
rect 98350 53910 98360 53980
rect 98140 53860 98360 53910
rect 98640 54090 98860 54140
rect 98640 54020 98650 54090
rect 98850 54020 98860 54090
rect 98640 53980 98860 54020
rect 98640 53910 98650 53980
rect 98850 53910 98860 53980
rect 98640 53860 98860 53910
rect 99140 54090 99360 54140
rect 99140 54020 99150 54090
rect 99350 54020 99360 54090
rect 99140 53980 99360 54020
rect 99140 53910 99150 53980
rect 99350 53910 99360 53980
rect 99140 53860 99360 53910
rect 99640 54090 99860 54140
rect 99640 54020 99650 54090
rect 99850 54020 99860 54090
rect 99640 53980 99860 54020
rect 99640 53910 99650 53980
rect 99850 53910 99860 53980
rect 99640 53860 99860 53910
rect -16000 53850 -12000 53860
rect -16000 53650 -15980 53850
rect -15910 53650 -15590 53850
rect -15520 53650 -15480 53850
rect -15410 53650 -15090 53850
rect -15020 53650 -14980 53850
rect -14910 53650 -14590 53850
rect -14520 53650 -14480 53850
rect -14410 53650 -14090 53850
rect -14020 53650 -13980 53850
rect -13910 53650 -13590 53850
rect -13520 53650 -13480 53850
rect -13410 53650 -13090 53850
rect -13020 53650 -12980 53850
rect -12910 53650 -12590 53850
rect -12520 53650 -12480 53850
rect -12410 53650 -12090 53850
rect -12020 53650 -12000 53850
rect -16000 53640 -12000 53650
rect 96000 53850 100000 53860
rect 96000 53650 96020 53850
rect 96090 53650 96410 53850
rect 96480 53650 96520 53850
rect 96590 53650 96910 53850
rect 96980 53650 97020 53850
rect 97090 53650 97410 53850
rect 97480 53650 97520 53850
rect 97590 53650 97910 53850
rect 97980 53650 98020 53850
rect 98090 53650 98410 53850
rect 98480 53650 98520 53850
rect 98590 53650 98910 53850
rect 98980 53650 99020 53850
rect 99090 53650 99410 53850
rect 99480 53650 99520 53850
rect 99590 53650 99910 53850
rect 99980 53650 100000 53850
rect 96000 53640 100000 53650
rect -15860 53590 -15640 53640
rect -15860 53520 -15850 53590
rect -15650 53520 -15640 53590
rect -15860 53480 -15640 53520
rect -15860 53410 -15850 53480
rect -15650 53410 -15640 53480
rect -15860 53360 -15640 53410
rect -15360 53590 -15140 53640
rect -15360 53520 -15350 53590
rect -15150 53520 -15140 53590
rect -15360 53480 -15140 53520
rect -15360 53410 -15350 53480
rect -15150 53410 -15140 53480
rect -15360 53360 -15140 53410
rect -14860 53590 -14640 53640
rect -14860 53520 -14850 53590
rect -14650 53520 -14640 53590
rect -14860 53480 -14640 53520
rect -14860 53410 -14850 53480
rect -14650 53410 -14640 53480
rect -14860 53360 -14640 53410
rect -14360 53590 -14140 53640
rect -14360 53520 -14350 53590
rect -14150 53520 -14140 53590
rect -14360 53480 -14140 53520
rect -14360 53410 -14350 53480
rect -14150 53410 -14140 53480
rect -14360 53360 -14140 53410
rect -13860 53590 -13640 53640
rect -13860 53520 -13850 53590
rect -13650 53520 -13640 53590
rect -13860 53480 -13640 53520
rect -13860 53410 -13850 53480
rect -13650 53410 -13640 53480
rect -13860 53360 -13640 53410
rect -13360 53590 -13140 53640
rect -13360 53520 -13350 53590
rect -13150 53520 -13140 53590
rect -13360 53480 -13140 53520
rect -13360 53410 -13350 53480
rect -13150 53410 -13140 53480
rect -13360 53360 -13140 53410
rect -12860 53590 -12640 53640
rect -12860 53520 -12850 53590
rect -12650 53520 -12640 53590
rect -12860 53480 -12640 53520
rect -12860 53410 -12850 53480
rect -12650 53410 -12640 53480
rect -12860 53360 -12640 53410
rect -12360 53590 -12140 53640
rect -12360 53520 -12350 53590
rect -12150 53520 -12140 53590
rect -12360 53480 -12140 53520
rect -12360 53410 -12350 53480
rect -12150 53410 -12140 53480
rect -12360 53360 -12140 53410
rect 96140 53590 96360 53640
rect 96140 53520 96150 53590
rect 96350 53520 96360 53590
rect 96140 53480 96360 53520
rect 96140 53410 96150 53480
rect 96350 53410 96360 53480
rect 96140 53360 96360 53410
rect 96640 53590 96860 53640
rect 96640 53520 96650 53590
rect 96850 53520 96860 53590
rect 96640 53480 96860 53520
rect 96640 53410 96650 53480
rect 96850 53410 96860 53480
rect 96640 53360 96860 53410
rect 97140 53590 97360 53640
rect 97140 53520 97150 53590
rect 97350 53520 97360 53590
rect 97140 53480 97360 53520
rect 97140 53410 97150 53480
rect 97350 53410 97360 53480
rect 97140 53360 97360 53410
rect 97640 53590 97860 53640
rect 97640 53520 97650 53590
rect 97850 53520 97860 53590
rect 97640 53480 97860 53520
rect 97640 53410 97650 53480
rect 97850 53410 97860 53480
rect 97640 53360 97860 53410
rect 98140 53590 98360 53640
rect 98140 53520 98150 53590
rect 98350 53520 98360 53590
rect 98140 53480 98360 53520
rect 98140 53410 98150 53480
rect 98350 53410 98360 53480
rect 98140 53360 98360 53410
rect 98640 53590 98860 53640
rect 98640 53520 98650 53590
rect 98850 53520 98860 53590
rect 98640 53480 98860 53520
rect 98640 53410 98650 53480
rect 98850 53410 98860 53480
rect 98640 53360 98860 53410
rect 99140 53590 99360 53640
rect 99140 53520 99150 53590
rect 99350 53520 99360 53590
rect 99140 53480 99360 53520
rect 99140 53410 99150 53480
rect 99350 53410 99360 53480
rect 99140 53360 99360 53410
rect 99640 53590 99860 53640
rect 99640 53520 99650 53590
rect 99850 53520 99860 53590
rect 99640 53480 99860 53520
rect 99640 53410 99650 53480
rect 99850 53410 99860 53480
rect 99640 53360 99860 53410
rect -16000 53350 -12000 53360
rect -16000 53150 -15980 53350
rect -15910 53150 -15590 53350
rect -15520 53150 -15480 53350
rect -15410 53150 -15090 53350
rect -15020 53150 -14980 53350
rect -14910 53150 -14590 53350
rect -14520 53150 -14480 53350
rect -14410 53150 -14090 53350
rect -14020 53150 -13980 53350
rect -13910 53150 -13590 53350
rect -13520 53150 -13480 53350
rect -13410 53150 -13090 53350
rect -13020 53150 -12980 53350
rect -12910 53150 -12590 53350
rect -12520 53150 -12480 53350
rect -12410 53150 -12090 53350
rect -12020 53150 -12000 53350
rect -16000 53140 -12000 53150
rect 96000 53350 100000 53360
rect 96000 53150 96020 53350
rect 96090 53150 96410 53350
rect 96480 53150 96520 53350
rect 96590 53150 96910 53350
rect 96980 53150 97020 53350
rect 97090 53150 97410 53350
rect 97480 53150 97520 53350
rect 97590 53150 97910 53350
rect 97980 53150 98020 53350
rect 98090 53150 98410 53350
rect 98480 53150 98520 53350
rect 98590 53150 98910 53350
rect 98980 53150 99020 53350
rect 99090 53150 99410 53350
rect 99480 53150 99520 53350
rect 99590 53150 99910 53350
rect 99980 53150 100000 53350
rect 96000 53140 100000 53150
rect -15860 53090 -15640 53140
rect -15860 53020 -15850 53090
rect -15650 53020 -15640 53090
rect -15860 52980 -15640 53020
rect -15860 52910 -15850 52980
rect -15650 52910 -15640 52980
rect -15860 52860 -15640 52910
rect -15360 53090 -15140 53140
rect -15360 53020 -15350 53090
rect -15150 53020 -15140 53090
rect -15360 52980 -15140 53020
rect -15360 52910 -15350 52980
rect -15150 52910 -15140 52980
rect -15360 52860 -15140 52910
rect -14860 53090 -14640 53140
rect -14860 53020 -14850 53090
rect -14650 53020 -14640 53090
rect -14860 52980 -14640 53020
rect -14860 52910 -14850 52980
rect -14650 52910 -14640 52980
rect -14860 52860 -14640 52910
rect -14360 53090 -14140 53140
rect -14360 53020 -14350 53090
rect -14150 53020 -14140 53090
rect -14360 52980 -14140 53020
rect -14360 52910 -14350 52980
rect -14150 52910 -14140 52980
rect -14360 52860 -14140 52910
rect -13860 53090 -13640 53140
rect -13860 53020 -13850 53090
rect -13650 53020 -13640 53090
rect -13860 52980 -13640 53020
rect -13860 52910 -13850 52980
rect -13650 52910 -13640 52980
rect -13860 52860 -13640 52910
rect -13360 53090 -13140 53140
rect -13360 53020 -13350 53090
rect -13150 53020 -13140 53090
rect -13360 52980 -13140 53020
rect -13360 52910 -13350 52980
rect -13150 52910 -13140 52980
rect -13360 52860 -13140 52910
rect -12860 53090 -12640 53140
rect -12860 53020 -12850 53090
rect -12650 53020 -12640 53090
rect -12860 52980 -12640 53020
rect -12860 52910 -12850 52980
rect -12650 52910 -12640 52980
rect -12860 52860 -12640 52910
rect -12360 53090 -12140 53140
rect -12360 53020 -12350 53090
rect -12150 53020 -12140 53090
rect -12360 52980 -12140 53020
rect -12360 52910 -12350 52980
rect -12150 52910 -12140 52980
rect -12360 52860 -12140 52910
rect 96140 53090 96360 53140
rect 96140 53020 96150 53090
rect 96350 53020 96360 53090
rect 96140 52980 96360 53020
rect 96140 52910 96150 52980
rect 96350 52910 96360 52980
rect 96140 52860 96360 52910
rect 96640 53090 96860 53140
rect 96640 53020 96650 53090
rect 96850 53020 96860 53090
rect 96640 52980 96860 53020
rect 96640 52910 96650 52980
rect 96850 52910 96860 52980
rect 96640 52860 96860 52910
rect 97140 53090 97360 53140
rect 97140 53020 97150 53090
rect 97350 53020 97360 53090
rect 97140 52980 97360 53020
rect 97140 52910 97150 52980
rect 97350 52910 97360 52980
rect 97140 52860 97360 52910
rect 97640 53090 97860 53140
rect 97640 53020 97650 53090
rect 97850 53020 97860 53090
rect 97640 52980 97860 53020
rect 97640 52910 97650 52980
rect 97850 52910 97860 52980
rect 97640 52860 97860 52910
rect 98140 53090 98360 53140
rect 98140 53020 98150 53090
rect 98350 53020 98360 53090
rect 98140 52980 98360 53020
rect 98140 52910 98150 52980
rect 98350 52910 98360 52980
rect 98140 52860 98360 52910
rect 98640 53090 98860 53140
rect 98640 53020 98650 53090
rect 98850 53020 98860 53090
rect 98640 52980 98860 53020
rect 98640 52910 98650 52980
rect 98850 52910 98860 52980
rect 98640 52860 98860 52910
rect 99140 53090 99360 53140
rect 99140 53020 99150 53090
rect 99350 53020 99360 53090
rect 99140 52980 99360 53020
rect 99140 52910 99150 52980
rect 99350 52910 99360 52980
rect 99140 52860 99360 52910
rect 99640 53090 99860 53140
rect 99640 53020 99650 53090
rect 99850 53020 99860 53090
rect 99640 52980 99860 53020
rect 99640 52910 99650 52980
rect 99850 52910 99860 52980
rect 99640 52860 99860 52910
rect -16000 52850 -12000 52860
rect -16000 52650 -15980 52850
rect -15910 52650 -15590 52850
rect -15520 52650 -15480 52850
rect -15410 52650 -15090 52850
rect -15020 52650 -14980 52850
rect -14910 52650 -14590 52850
rect -14520 52650 -14480 52850
rect -14410 52650 -14090 52850
rect -14020 52650 -13980 52850
rect -13910 52650 -13590 52850
rect -13520 52650 -13480 52850
rect -13410 52650 -13090 52850
rect -13020 52650 -12980 52850
rect -12910 52650 -12590 52850
rect -12520 52650 -12480 52850
rect -12410 52650 -12090 52850
rect -12020 52650 -12000 52850
rect -16000 52640 -12000 52650
rect 96000 52850 100000 52860
rect 96000 52650 96020 52850
rect 96090 52650 96410 52850
rect 96480 52650 96520 52850
rect 96590 52650 96910 52850
rect 96980 52650 97020 52850
rect 97090 52650 97410 52850
rect 97480 52650 97520 52850
rect 97590 52650 97910 52850
rect 97980 52650 98020 52850
rect 98090 52650 98410 52850
rect 98480 52650 98520 52850
rect 98590 52650 98910 52850
rect 98980 52650 99020 52850
rect 99090 52650 99410 52850
rect 99480 52650 99520 52850
rect 99590 52650 99910 52850
rect 99980 52650 100000 52850
rect 96000 52640 100000 52650
rect -15860 52590 -15640 52640
rect -15860 52520 -15850 52590
rect -15650 52520 -15640 52590
rect -15860 52480 -15640 52520
rect -15860 52410 -15850 52480
rect -15650 52410 -15640 52480
rect -15860 52360 -15640 52410
rect -15360 52590 -15140 52640
rect -15360 52520 -15350 52590
rect -15150 52520 -15140 52590
rect -15360 52480 -15140 52520
rect -15360 52410 -15350 52480
rect -15150 52410 -15140 52480
rect -15360 52360 -15140 52410
rect -14860 52590 -14640 52640
rect -14860 52520 -14850 52590
rect -14650 52520 -14640 52590
rect -14860 52480 -14640 52520
rect -14860 52410 -14850 52480
rect -14650 52410 -14640 52480
rect -14860 52360 -14640 52410
rect -14360 52590 -14140 52640
rect -14360 52520 -14350 52590
rect -14150 52520 -14140 52590
rect -14360 52480 -14140 52520
rect -14360 52410 -14350 52480
rect -14150 52410 -14140 52480
rect -14360 52360 -14140 52410
rect -13860 52590 -13640 52640
rect -13860 52520 -13850 52590
rect -13650 52520 -13640 52590
rect -13860 52480 -13640 52520
rect -13860 52410 -13850 52480
rect -13650 52410 -13640 52480
rect -13860 52360 -13640 52410
rect -13360 52590 -13140 52640
rect -13360 52520 -13350 52590
rect -13150 52520 -13140 52590
rect -13360 52480 -13140 52520
rect -13360 52410 -13350 52480
rect -13150 52410 -13140 52480
rect -13360 52360 -13140 52410
rect -12860 52590 -12640 52640
rect -12860 52520 -12850 52590
rect -12650 52520 -12640 52590
rect -12860 52480 -12640 52520
rect -12860 52410 -12850 52480
rect -12650 52410 -12640 52480
rect -12860 52360 -12640 52410
rect -12360 52590 -12140 52640
rect -12360 52520 -12350 52590
rect -12150 52520 -12140 52590
rect -12360 52480 -12140 52520
rect -12360 52410 -12350 52480
rect -12150 52410 -12140 52480
rect -12360 52360 -12140 52410
rect 96140 52590 96360 52640
rect 96140 52520 96150 52590
rect 96350 52520 96360 52590
rect 96140 52480 96360 52520
rect 96140 52410 96150 52480
rect 96350 52410 96360 52480
rect 96140 52360 96360 52410
rect 96640 52590 96860 52640
rect 96640 52520 96650 52590
rect 96850 52520 96860 52590
rect 96640 52480 96860 52520
rect 96640 52410 96650 52480
rect 96850 52410 96860 52480
rect 96640 52360 96860 52410
rect 97140 52590 97360 52640
rect 97140 52520 97150 52590
rect 97350 52520 97360 52590
rect 97140 52480 97360 52520
rect 97140 52410 97150 52480
rect 97350 52410 97360 52480
rect 97140 52360 97360 52410
rect 97640 52590 97860 52640
rect 97640 52520 97650 52590
rect 97850 52520 97860 52590
rect 97640 52480 97860 52520
rect 97640 52410 97650 52480
rect 97850 52410 97860 52480
rect 97640 52360 97860 52410
rect 98140 52590 98360 52640
rect 98140 52520 98150 52590
rect 98350 52520 98360 52590
rect 98140 52480 98360 52520
rect 98140 52410 98150 52480
rect 98350 52410 98360 52480
rect 98140 52360 98360 52410
rect 98640 52590 98860 52640
rect 98640 52520 98650 52590
rect 98850 52520 98860 52590
rect 98640 52480 98860 52520
rect 98640 52410 98650 52480
rect 98850 52410 98860 52480
rect 98640 52360 98860 52410
rect 99140 52590 99360 52640
rect 99140 52520 99150 52590
rect 99350 52520 99360 52590
rect 99140 52480 99360 52520
rect 99140 52410 99150 52480
rect 99350 52410 99360 52480
rect 99140 52360 99360 52410
rect 99640 52590 99860 52640
rect 99640 52520 99650 52590
rect 99850 52520 99860 52590
rect 99640 52480 99860 52520
rect 99640 52410 99650 52480
rect 99850 52410 99860 52480
rect 99640 52360 99860 52410
rect -16000 52350 -12000 52360
rect -16000 52150 -15980 52350
rect -15910 52150 -15590 52350
rect -15520 52150 -15480 52350
rect -15410 52150 -15090 52350
rect -15020 52150 -14980 52350
rect -14910 52150 -14590 52350
rect -14520 52150 -14480 52350
rect -14410 52150 -14090 52350
rect -14020 52150 -13980 52350
rect -13910 52150 -13590 52350
rect -13520 52150 -13480 52350
rect -13410 52150 -13090 52350
rect -13020 52150 -12980 52350
rect -12910 52150 -12590 52350
rect -12520 52150 -12480 52350
rect -12410 52150 -12090 52350
rect -12020 52150 -12000 52350
rect -16000 52140 -12000 52150
rect 96000 52350 100000 52360
rect 96000 52150 96020 52350
rect 96090 52150 96410 52350
rect 96480 52150 96520 52350
rect 96590 52150 96910 52350
rect 96980 52150 97020 52350
rect 97090 52150 97410 52350
rect 97480 52150 97520 52350
rect 97590 52150 97910 52350
rect 97980 52150 98020 52350
rect 98090 52150 98410 52350
rect 98480 52150 98520 52350
rect 98590 52150 98910 52350
rect 98980 52150 99020 52350
rect 99090 52150 99410 52350
rect 99480 52150 99520 52350
rect 99590 52150 99910 52350
rect 99980 52150 100000 52350
rect 96000 52140 100000 52150
rect -15860 52090 -15640 52140
rect -15860 52020 -15850 52090
rect -15650 52020 -15640 52090
rect -15860 51980 -15640 52020
rect -15860 51910 -15850 51980
rect -15650 51910 -15640 51980
rect -15860 51860 -15640 51910
rect -15360 52090 -15140 52140
rect -15360 52020 -15350 52090
rect -15150 52020 -15140 52090
rect -15360 51980 -15140 52020
rect -15360 51910 -15350 51980
rect -15150 51910 -15140 51980
rect -15360 51860 -15140 51910
rect -14860 52090 -14640 52140
rect -14860 52020 -14850 52090
rect -14650 52020 -14640 52090
rect -14860 51980 -14640 52020
rect -14860 51910 -14850 51980
rect -14650 51910 -14640 51980
rect -14860 51860 -14640 51910
rect -14360 52090 -14140 52140
rect -14360 52020 -14350 52090
rect -14150 52020 -14140 52090
rect -14360 51980 -14140 52020
rect -14360 51910 -14350 51980
rect -14150 51910 -14140 51980
rect -14360 51860 -14140 51910
rect -13860 52090 -13640 52140
rect -13860 52020 -13850 52090
rect -13650 52020 -13640 52090
rect -13860 51980 -13640 52020
rect -13860 51910 -13850 51980
rect -13650 51910 -13640 51980
rect -13860 51860 -13640 51910
rect -13360 52090 -13140 52140
rect -13360 52020 -13350 52090
rect -13150 52020 -13140 52090
rect -13360 51980 -13140 52020
rect -13360 51910 -13350 51980
rect -13150 51910 -13140 51980
rect -13360 51860 -13140 51910
rect -12860 52090 -12640 52140
rect -12860 52020 -12850 52090
rect -12650 52020 -12640 52090
rect -12860 51980 -12640 52020
rect -12860 51910 -12850 51980
rect -12650 51910 -12640 51980
rect -12860 51860 -12640 51910
rect -12360 52090 -12140 52140
rect -12360 52020 -12350 52090
rect -12150 52020 -12140 52090
rect -12360 51980 -12140 52020
rect -12360 51910 -12350 51980
rect -12150 51910 -12140 51980
rect -12360 51860 -12140 51910
rect 96140 52090 96360 52140
rect 96140 52020 96150 52090
rect 96350 52020 96360 52090
rect 96140 51980 96360 52020
rect 96140 51910 96150 51980
rect 96350 51910 96360 51980
rect 96140 51860 96360 51910
rect 96640 52090 96860 52140
rect 96640 52020 96650 52090
rect 96850 52020 96860 52090
rect 96640 51980 96860 52020
rect 96640 51910 96650 51980
rect 96850 51910 96860 51980
rect 96640 51860 96860 51910
rect 97140 52090 97360 52140
rect 97140 52020 97150 52090
rect 97350 52020 97360 52090
rect 97140 51980 97360 52020
rect 97140 51910 97150 51980
rect 97350 51910 97360 51980
rect 97140 51860 97360 51910
rect 97640 52090 97860 52140
rect 97640 52020 97650 52090
rect 97850 52020 97860 52090
rect 97640 51980 97860 52020
rect 97640 51910 97650 51980
rect 97850 51910 97860 51980
rect 97640 51860 97860 51910
rect 98140 52090 98360 52140
rect 98140 52020 98150 52090
rect 98350 52020 98360 52090
rect 98140 51980 98360 52020
rect 98140 51910 98150 51980
rect 98350 51910 98360 51980
rect 98140 51860 98360 51910
rect 98640 52090 98860 52140
rect 98640 52020 98650 52090
rect 98850 52020 98860 52090
rect 98640 51980 98860 52020
rect 98640 51910 98650 51980
rect 98850 51910 98860 51980
rect 98640 51860 98860 51910
rect 99140 52090 99360 52140
rect 99140 52020 99150 52090
rect 99350 52020 99360 52090
rect 99140 51980 99360 52020
rect 99140 51910 99150 51980
rect 99350 51910 99360 51980
rect 99140 51860 99360 51910
rect 99640 52090 99860 52140
rect 99640 52020 99650 52090
rect 99850 52020 99860 52090
rect 99640 51980 99860 52020
rect 99640 51910 99650 51980
rect 99850 51910 99860 51980
rect 99640 51860 99860 51910
rect -16000 51850 -12000 51860
rect -16000 51650 -15980 51850
rect -15910 51650 -15590 51850
rect -15520 51650 -15480 51850
rect -15410 51650 -15090 51850
rect -15020 51650 -14980 51850
rect -14910 51650 -14590 51850
rect -14520 51650 -14480 51850
rect -14410 51650 -14090 51850
rect -14020 51650 -13980 51850
rect -13910 51650 -13590 51850
rect -13520 51650 -13480 51850
rect -13410 51650 -13090 51850
rect -13020 51650 -12980 51850
rect -12910 51650 -12590 51850
rect -12520 51650 -12480 51850
rect -12410 51650 -12090 51850
rect -12020 51650 -12000 51850
rect -16000 51640 -12000 51650
rect 96000 51850 100000 51860
rect 96000 51650 96020 51850
rect 96090 51650 96410 51850
rect 96480 51650 96520 51850
rect 96590 51650 96910 51850
rect 96980 51650 97020 51850
rect 97090 51650 97410 51850
rect 97480 51650 97520 51850
rect 97590 51650 97910 51850
rect 97980 51650 98020 51850
rect 98090 51650 98410 51850
rect 98480 51650 98520 51850
rect 98590 51650 98910 51850
rect 98980 51650 99020 51850
rect 99090 51650 99410 51850
rect 99480 51650 99520 51850
rect 99590 51650 99910 51850
rect 99980 51650 100000 51850
rect 96000 51640 100000 51650
rect -15860 51590 -15640 51640
rect -15860 51520 -15850 51590
rect -15650 51520 -15640 51590
rect -15860 51480 -15640 51520
rect -15860 51410 -15850 51480
rect -15650 51410 -15640 51480
rect -15860 51360 -15640 51410
rect -15360 51590 -15140 51640
rect -15360 51520 -15350 51590
rect -15150 51520 -15140 51590
rect -15360 51480 -15140 51520
rect -15360 51410 -15350 51480
rect -15150 51410 -15140 51480
rect -15360 51360 -15140 51410
rect -14860 51590 -14640 51640
rect -14860 51520 -14850 51590
rect -14650 51520 -14640 51590
rect -14860 51480 -14640 51520
rect -14860 51410 -14850 51480
rect -14650 51410 -14640 51480
rect -14860 51360 -14640 51410
rect -14360 51590 -14140 51640
rect -14360 51520 -14350 51590
rect -14150 51520 -14140 51590
rect -14360 51480 -14140 51520
rect -14360 51410 -14350 51480
rect -14150 51410 -14140 51480
rect -14360 51360 -14140 51410
rect -13860 51590 -13640 51640
rect -13860 51520 -13850 51590
rect -13650 51520 -13640 51590
rect -13860 51480 -13640 51520
rect -13860 51410 -13850 51480
rect -13650 51410 -13640 51480
rect -13860 51360 -13640 51410
rect -13360 51590 -13140 51640
rect -13360 51520 -13350 51590
rect -13150 51520 -13140 51590
rect -13360 51480 -13140 51520
rect -13360 51410 -13350 51480
rect -13150 51410 -13140 51480
rect -13360 51360 -13140 51410
rect -12860 51590 -12640 51640
rect -12860 51520 -12850 51590
rect -12650 51520 -12640 51590
rect -12860 51480 -12640 51520
rect -12860 51410 -12850 51480
rect -12650 51410 -12640 51480
rect -12860 51360 -12640 51410
rect -12360 51590 -12140 51640
rect -12360 51520 -12350 51590
rect -12150 51520 -12140 51590
rect -12360 51480 -12140 51520
rect -12360 51410 -12350 51480
rect -12150 51410 -12140 51480
rect -12360 51360 -12140 51410
rect 96140 51590 96360 51640
rect 96140 51520 96150 51590
rect 96350 51520 96360 51590
rect 96140 51480 96360 51520
rect 96140 51410 96150 51480
rect 96350 51410 96360 51480
rect 96140 51360 96360 51410
rect 96640 51590 96860 51640
rect 96640 51520 96650 51590
rect 96850 51520 96860 51590
rect 96640 51480 96860 51520
rect 96640 51410 96650 51480
rect 96850 51410 96860 51480
rect 96640 51360 96860 51410
rect 97140 51590 97360 51640
rect 97140 51520 97150 51590
rect 97350 51520 97360 51590
rect 97140 51480 97360 51520
rect 97140 51410 97150 51480
rect 97350 51410 97360 51480
rect 97140 51360 97360 51410
rect 97640 51590 97860 51640
rect 97640 51520 97650 51590
rect 97850 51520 97860 51590
rect 97640 51480 97860 51520
rect 97640 51410 97650 51480
rect 97850 51410 97860 51480
rect 97640 51360 97860 51410
rect 98140 51590 98360 51640
rect 98140 51520 98150 51590
rect 98350 51520 98360 51590
rect 98140 51480 98360 51520
rect 98140 51410 98150 51480
rect 98350 51410 98360 51480
rect 98140 51360 98360 51410
rect 98640 51590 98860 51640
rect 98640 51520 98650 51590
rect 98850 51520 98860 51590
rect 98640 51480 98860 51520
rect 98640 51410 98650 51480
rect 98850 51410 98860 51480
rect 98640 51360 98860 51410
rect 99140 51590 99360 51640
rect 99140 51520 99150 51590
rect 99350 51520 99360 51590
rect 99140 51480 99360 51520
rect 99140 51410 99150 51480
rect 99350 51410 99360 51480
rect 99140 51360 99360 51410
rect 99640 51590 99860 51640
rect 99640 51520 99650 51590
rect 99850 51520 99860 51590
rect 99640 51480 99860 51520
rect 99640 51410 99650 51480
rect 99850 51410 99860 51480
rect 99640 51360 99860 51410
rect -16000 51350 -12000 51360
rect -16000 51150 -15980 51350
rect -15910 51150 -15590 51350
rect -15520 51150 -15480 51350
rect -15410 51150 -15090 51350
rect -15020 51150 -14980 51350
rect -14910 51150 -14590 51350
rect -14520 51150 -14480 51350
rect -14410 51150 -14090 51350
rect -14020 51150 -13980 51350
rect -13910 51150 -13590 51350
rect -13520 51150 -13480 51350
rect -13410 51150 -13090 51350
rect -13020 51150 -12980 51350
rect -12910 51150 -12590 51350
rect -12520 51150 -12480 51350
rect -12410 51150 -12090 51350
rect -12020 51150 -12000 51350
rect -16000 51140 -12000 51150
rect 96000 51350 100000 51360
rect 96000 51150 96020 51350
rect 96090 51150 96410 51350
rect 96480 51150 96520 51350
rect 96590 51150 96910 51350
rect 96980 51150 97020 51350
rect 97090 51150 97410 51350
rect 97480 51150 97520 51350
rect 97590 51150 97910 51350
rect 97980 51150 98020 51350
rect 98090 51150 98410 51350
rect 98480 51150 98520 51350
rect 98590 51150 98910 51350
rect 98980 51150 99020 51350
rect 99090 51150 99410 51350
rect 99480 51150 99520 51350
rect 99590 51150 99910 51350
rect 99980 51150 100000 51350
rect 96000 51140 100000 51150
rect -15860 51090 -15640 51140
rect -15860 51020 -15850 51090
rect -15650 51020 -15640 51090
rect -15860 50980 -15640 51020
rect -15860 50910 -15850 50980
rect -15650 50910 -15640 50980
rect -15860 50860 -15640 50910
rect -15360 51090 -15140 51140
rect -15360 51020 -15350 51090
rect -15150 51020 -15140 51090
rect -15360 50980 -15140 51020
rect -15360 50910 -15350 50980
rect -15150 50910 -15140 50980
rect -15360 50860 -15140 50910
rect -14860 51090 -14640 51140
rect -14860 51020 -14850 51090
rect -14650 51020 -14640 51090
rect -14860 50980 -14640 51020
rect -14860 50910 -14850 50980
rect -14650 50910 -14640 50980
rect -14860 50860 -14640 50910
rect -14360 51090 -14140 51140
rect -14360 51020 -14350 51090
rect -14150 51020 -14140 51090
rect -14360 50980 -14140 51020
rect -14360 50910 -14350 50980
rect -14150 50910 -14140 50980
rect -14360 50860 -14140 50910
rect -13860 51090 -13640 51140
rect -13860 51020 -13850 51090
rect -13650 51020 -13640 51090
rect -13860 50980 -13640 51020
rect -13860 50910 -13850 50980
rect -13650 50910 -13640 50980
rect -13860 50860 -13640 50910
rect -13360 51090 -13140 51140
rect -13360 51020 -13350 51090
rect -13150 51020 -13140 51090
rect -13360 50980 -13140 51020
rect -13360 50910 -13350 50980
rect -13150 50910 -13140 50980
rect -13360 50860 -13140 50910
rect -12860 51090 -12640 51140
rect -12860 51020 -12850 51090
rect -12650 51020 -12640 51090
rect -12860 50980 -12640 51020
rect -12860 50910 -12850 50980
rect -12650 50910 -12640 50980
rect -12860 50860 -12640 50910
rect -12360 51090 -12140 51140
rect -12360 51020 -12350 51090
rect -12150 51020 -12140 51090
rect -12360 50980 -12140 51020
rect -12360 50910 -12350 50980
rect -12150 50910 -12140 50980
rect -12360 50860 -12140 50910
rect 96140 51090 96360 51140
rect 96140 51020 96150 51090
rect 96350 51020 96360 51090
rect 96140 50980 96360 51020
rect 96140 50910 96150 50980
rect 96350 50910 96360 50980
rect 96140 50860 96360 50910
rect 96640 51090 96860 51140
rect 96640 51020 96650 51090
rect 96850 51020 96860 51090
rect 96640 50980 96860 51020
rect 96640 50910 96650 50980
rect 96850 50910 96860 50980
rect 96640 50860 96860 50910
rect 97140 51090 97360 51140
rect 97140 51020 97150 51090
rect 97350 51020 97360 51090
rect 97140 50980 97360 51020
rect 97140 50910 97150 50980
rect 97350 50910 97360 50980
rect 97140 50860 97360 50910
rect 97640 51090 97860 51140
rect 97640 51020 97650 51090
rect 97850 51020 97860 51090
rect 97640 50980 97860 51020
rect 97640 50910 97650 50980
rect 97850 50910 97860 50980
rect 97640 50860 97860 50910
rect 98140 51090 98360 51140
rect 98140 51020 98150 51090
rect 98350 51020 98360 51090
rect 98140 50980 98360 51020
rect 98140 50910 98150 50980
rect 98350 50910 98360 50980
rect 98140 50860 98360 50910
rect 98640 51090 98860 51140
rect 98640 51020 98650 51090
rect 98850 51020 98860 51090
rect 98640 50980 98860 51020
rect 98640 50910 98650 50980
rect 98850 50910 98860 50980
rect 98640 50860 98860 50910
rect 99140 51090 99360 51140
rect 99140 51020 99150 51090
rect 99350 51020 99360 51090
rect 99140 50980 99360 51020
rect 99140 50910 99150 50980
rect 99350 50910 99360 50980
rect 99140 50860 99360 50910
rect 99640 51090 99860 51140
rect 99640 51020 99650 51090
rect 99850 51020 99860 51090
rect 99640 50980 99860 51020
rect 99640 50910 99650 50980
rect 99850 50910 99860 50980
rect 99640 50860 99860 50910
rect -16000 50850 -12000 50860
rect -16000 50650 -15980 50850
rect -15910 50650 -15590 50850
rect -15520 50650 -15480 50850
rect -15410 50650 -15090 50850
rect -15020 50650 -14980 50850
rect -14910 50650 -14590 50850
rect -14520 50650 -14480 50850
rect -14410 50650 -14090 50850
rect -14020 50650 -13980 50850
rect -13910 50650 -13590 50850
rect -13520 50650 -13480 50850
rect -13410 50650 -13090 50850
rect -13020 50650 -12980 50850
rect -12910 50650 -12590 50850
rect -12520 50650 -12480 50850
rect -12410 50650 -12090 50850
rect -12020 50650 -12000 50850
rect -16000 50640 -12000 50650
rect 96000 50850 100000 50860
rect 96000 50650 96020 50850
rect 96090 50650 96410 50850
rect 96480 50650 96520 50850
rect 96590 50650 96910 50850
rect 96980 50650 97020 50850
rect 97090 50650 97410 50850
rect 97480 50650 97520 50850
rect 97590 50650 97910 50850
rect 97980 50650 98020 50850
rect 98090 50650 98410 50850
rect 98480 50650 98520 50850
rect 98590 50650 98910 50850
rect 98980 50650 99020 50850
rect 99090 50650 99410 50850
rect 99480 50650 99520 50850
rect 99590 50650 99910 50850
rect 99980 50650 100000 50850
rect 96000 50640 100000 50650
rect -15860 50590 -15640 50640
rect -15860 50520 -15850 50590
rect -15650 50520 -15640 50590
rect -15860 50480 -15640 50520
rect -15860 50410 -15850 50480
rect -15650 50410 -15640 50480
rect -15860 50360 -15640 50410
rect -15360 50590 -15140 50640
rect -15360 50520 -15350 50590
rect -15150 50520 -15140 50590
rect -15360 50480 -15140 50520
rect -15360 50410 -15350 50480
rect -15150 50410 -15140 50480
rect -15360 50360 -15140 50410
rect -14860 50590 -14640 50640
rect -14860 50520 -14850 50590
rect -14650 50520 -14640 50590
rect -14860 50480 -14640 50520
rect -14860 50410 -14850 50480
rect -14650 50410 -14640 50480
rect -14860 50360 -14640 50410
rect -14360 50590 -14140 50640
rect -14360 50520 -14350 50590
rect -14150 50520 -14140 50590
rect -14360 50480 -14140 50520
rect -14360 50410 -14350 50480
rect -14150 50410 -14140 50480
rect -14360 50360 -14140 50410
rect -13860 50590 -13640 50640
rect -13860 50520 -13850 50590
rect -13650 50520 -13640 50590
rect -13860 50480 -13640 50520
rect -13860 50410 -13850 50480
rect -13650 50410 -13640 50480
rect -13860 50360 -13640 50410
rect -13360 50590 -13140 50640
rect -13360 50520 -13350 50590
rect -13150 50520 -13140 50590
rect -13360 50480 -13140 50520
rect -13360 50410 -13350 50480
rect -13150 50410 -13140 50480
rect -13360 50360 -13140 50410
rect -12860 50590 -12640 50640
rect -12860 50520 -12850 50590
rect -12650 50520 -12640 50590
rect -12860 50480 -12640 50520
rect -12860 50410 -12850 50480
rect -12650 50410 -12640 50480
rect -12860 50360 -12640 50410
rect -12360 50590 -12140 50640
rect -12360 50520 -12350 50590
rect -12150 50520 -12140 50590
rect -12360 50480 -12140 50520
rect -12360 50410 -12350 50480
rect -12150 50410 -12140 50480
rect -12360 50360 -12140 50410
rect 96140 50590 96360 50640
rect 96140 50520 96150 50590
rect 96350 50520 96360 50590
rect 96140 50480 96360 50520
rect 96140 50410 96150 50480
rect 96350 50410 96360 50480
rect 96140 50360 96360 50410
rect 96640 50590 96860 50640
rect 96640 50520 96650 50590
rect 96850 50520 96860 50590
rect 96640 50480 96860 50520
rect 96640 50410 96650 50480
rect 96850 50410 96860 50480
rect 96640 50360 96860 50410
rect 97140 50590 97360 50640
rect 97140 50520 97150 50590
rect 97350 50520 97360 50590
rect 97140 50480 97360 50520
rect 97140 50410 97150 50480
rect 97350 50410 97360 50480
rect 97140 50360 97360 50410
rect 97640 50590 97860 50640
rect 97640 50520 97650 50590
rect 97850 50520 97860 50590
rect 97640 50480 97860 50520
rect 97640 50410 97650 50480
rect 97850 50410 97860 50480
rect 97640 50360 97860 50410
rect 98140 50590 98360 50640
rect 98140 50520 98150 50590
rect 98350 50520 98360 50590
rect 98140 50480 98360 50520
rect 98140 50410 98150 50480
rect 98350 50410 98360 50480
rect 98140 50360 98360 50410
rect 98640 50590 98860 50640
rect 98640 50520 98650 50590
rect 98850 50520 98860 50590
rect 98640 50480 98860 50520
rect 98640 50410 98650 50480
rect 98850 50410 98860 50480
rect 98640 50360 98860 50410
rect 99140 50590 99360 50640
rect 99140 50520 99150 50590
rect 99350 50520 99360 50590
rect 99140 50480 99360 50520
rect 99140 50410 99150 50480
rect 99350 50410 99360 50480
rect 99140 50360 99360 50410
rect 99640 50590 99860 50640
rect 99640 50520 99650 50590
rect 99850 50520 99860 50590
rect 99640 50480 99860 50520
rect 99640 50410 99650 50480
rect 99850 50410 99860 50480
rect 99640 50360 99860 50410
rect -16000 50350 -12000 50360
rect -16000 50150 -15980 50350
rect -15910 50150 -15590 50350
rect -15520 50150 -15480 50350
rect -15410 50150 -15090 50350
rect -15020 50150 -14980 50350
rect -14910 50150 -14590 50350
rect -14520 50150 -14480 50350
rect -14410 50150 -14090 50350
rect -14020 50150 -13980 50350
rect -13910 50150 -13590 50350
rect -13520 50150 -13480 50350
rect -13410 50150 -13090 50350
rect -13020 50150 -12980 50350
rect -12910 50150 -12590 50350
rect -12520 50150 -12480 50350
rect -12410 50150 -12090 50350
rect -12020 50150 -12000 50350
rect -16000 50140 -12000 50150
rect 96000 50350 100000 50360
rect 96000 50150 96020 50350
rect 96090 50150 96410 50350
rect 96480 50150 96520 50350
rect 96590 50150 96910 50350
rect 96980 50150 97020 50350
rect 97090 50150 97410 50350
rect 97480 50150 97520 50350
rect 97590 50150 97910 50350
rect 97980 50150 98020 50350
rect 98090 50150 98410 50350
rect 98480 50150 98520 50350
rect 98590 50150 98910 50350
rect 98980 50150 99020 50350
rect 99090 50150 99410 50350
rect 99480 50150 99520 50350
rect 99590 50150 99910 50350
rect 99980 50150 100000 50350
rect 96000 50140 100000 50150
rect -15860 50090 -15640 50140
rect -15860 50020 -15850 50090
rect -15650 50020 -15640 50090
rect -15860 49980 -15640 50020
rect -15860 49910 -15850 49980
rect -15650 49910 -15640 49980
rect -15860 49860 -15640 49910
rect -15360 50090 -15140 50140
rect -15360 50020 -15350 50090
rect -15150 50020 -15140 50090
rect -15360 49980 -15140 50020
rect -15360 49910 -15350 49980
rect -15150 49910 -15140 49980
rect -15360 49860 -15140 49910
rect -14860 50090 -14640 50140
rect -14860 50020 -14850 50090
rect -14650 50020 -14640 50090
rect -14860 49980 -14640 50020
rect -14860 49910 -14850 49980
rect -14650 49910 -14640 49980
rect -14860 49860 -14640 49910
rect -14360 50090 -14140 50140
rect -14360 50020 -14350 50090
rect -14150 50020 -14140 50090
rect -14360 49980 -14140 50020
rect -14360 49910 -14350 49980
rect -14150 49910 -14140 49980
rect -14360 49860 -14140 49910
rect -13860 50090 -13640 50140
rect -13860 50020 -13850 50090
rect -13650 50020 -13640 50090
rect -13860 49980 -13640 50020
rect -13860 49910 -13850 49980
rect -13650 49910 -13640 49980
rect -13860 49860 -13640 49910
rect -13360 50090 -13140 50140
rect -13360 50020 -13350 50090
rect -13150 50020 -13140 50090
rect -13360 49980 -13140 50020
rect -13360 49910 -13350 49980
rect -13150 49910 -13140 49980
rect -13360 49860 -13140 49910
rect -12860 50090 -12640 50140
rect -12860 50020 -12850 50090
rect -12650 50020 -12640 50090
rect -12860 49980 -12640 50020
rect -12860 49910 -12850 49980
rect -12650 49910 -12640 49980
rect -12860 49860 -12640 49910
rect -12360 50090 -12140 50140
rect -12360 50020 -12350 50090
rect -12150 50020 -12140 50090
rect -12360 49980 -12140 50020
rect 96140 50090 96360 50140
rect 96140 50020 96150 50090
rect 96350 50020 96360 50090
rect 96140 50000 96360 50020
rect 96640 50090 96860 50140
rect 96640 50020 96650 50090
rect 96850 50020 96860 50090
rect 96640 50000 96860 50020
rect 97140 50090 97360 50140
rect 97140 50020 97150 50090
rect 97350 50020 97360 50090
rect 97140 50000 97360 50020
rect 97640 50090 97860 50140
rect 97640 50020 97650 50090
rect 97850 50020 97860 50090
rect 97640 50000 97860 50020
rect 98140 50090 98360 50140
rect 98140 50020 98150 50090
rect 98350 50020 98360 50090
rect 98140 50000 98360 50020
rect 98640 50090 98860 50140
rect 98640 50020 98650 50090
rect 98850 50020 98860 50090
rect 98640 50000 98860 50020
rect 99140 50090 99360 50140
rect 99140 50020 99150 50090
rect 99350 50020 99360 50090
rect 99140 50000 99360 50020
rect 99640 50090 99860 50140
rect 99640 50020 99650 50090
rect 99850 50020 99860 50090
rect 99640 50000 99860 50020
rect -12360 49910 -12350 49980
rect -12150 49910 -12140 49980
rect -12360 49860 -12140 49910
rect -16000 49850 -12000 49860
rect -16000 49650 -15980 49850
rect -15910 49650 -15590 49850
rect -15520 49650 -15480 49850
rect -15410 49650 -15090 49850
rect -15020 49650 -14980 49850
rect -14910 49650 -14590 49850
rect -14520 49650 -14480 49850
rect -14410 49650 -14090 49850
rect -14020 49650 -13980 49850
rect -13910 49650 -13590 49850
rect -13520 49650 -13480 49850
rect -13410 49650 -13090 49850
rect -13020 49650 -12980 49850
rect -12910 49650 -12590 49850
rect -12520 49650 -12480 49850
rect -12410 49650 -12090 49850
rect -12020 49650 -12000 49850
rect -16000 49640 -12000 49650
rect -15860 49590 -15640 49640
rect -15860 49520 -15850 49590
rect -15650 49520 -15640 49590
rect -15860 49480 -15640 49520
rect -15860 49410 -15850 49480
rect -15650 49410 -15640 49480
rect -15860 49360 -15640 49410
rect -15360 49590 -15140 49640
rect -15360 49520 -15350 49590
rect -15150 49520 -15140 49590
rect -15360 49480 -15140 49520
rect -15360 49410 -15350 49480
rect -15150 49410 -15140 49480
rect -15360 49360 -15140 49410
rect -14860 49590 -14640 49640
rect -14860 49520 -14850 49590
rect -14650 49520 -14640 49590
rect -14860 49480 -14640 49520
rect -14860 49410 -14850 49480
rect -14650 49410 -14640 49480
rect -14860 49360 -14640 49410
rect -14360 49590 -14140 49640
rect -14360 49520 -14350 49590
rect -14150 49520 -14140 49590
rect -14360 49480 -14140 49520
rect -14360 49410 -14350 49480
rect -14150 49410 -14140 49480
rect -14360 49360 -14140 49410
rect -13860 49590 -13640 49640
rect -13860 49520 -13850 49590
rect -13650 49520 -13640 49590
rect -13860 49480 -13640 49520
rect -13860 49410 -13850 49480
rect -13650 49410 -13640 49480
rect -13860 49360 -13640 49410
rect -13360 49590 -13140 49640
rect -13360 49520 -13350 49590
rect -13150 49520 -13140 49590
rect -13360 49480 -13140 49520
rect -13360 49410 -13350 49480
rect -13150 49410 -13140 49480
rect -13360 49360 -13140 49410
rect -12860 49590 -12640 49640
rect -12860 49520 -12850 49590
rect -12650 49520 -12640 49590
rect -12860 49480 -12640 49520
rect -12860 49410 -12850 49480
rect -12650 49410 -12640 49480
rect -12860 49360 -12640 49410
rect -12360 49590 -12140 49640
rect -12360 49520 -12350 49590
rect -12150 49520 -12140 49590
rect -12360 49480 -12140 49520
rect -12360 49410 -12350 49480
rect -12150 49410 -12140 49480
rect -12360 49360 -12140 49410
rect -16000 49350 -12000 49360
rect -16000 49150 -15980 49350
rect -15910 49150 -15590 49350
rect -15520 49150 -15480 49350
rect -15410 49150 -15090 49350
rect -15020 49150 -14980 49350
rect -14910 49150 -14590 49350
rect -14520 49150 -14480 49350
rect -14410 49150 -14090 49350
rect -14020 49150 -13980 49350
rect -13910 49150 -13590 49350
rect -13520 49150 -13480 49350
rect -13410 49150 -13090 49350
rect -13020 49150 -12980 49350
rect -12910 49150 -12590 49350
rect -12520 49150 -12480 49350
rect -12410 49150 -12090 49350
rect -12020 49150 -12000 49350
rect -16000 49140 -12000 49150
rect -15860 49090 -15640 49140
rect -15860 49020 -15850 49090
rect -15650 49020 -15640 49090
rect -15860 48980 -15640 49020
rect -15860 48910 -15850 48980
rect -15650 48910 -15640 48980
rect -15860 48860 -15640 48910
rect -15360 49090 -15140 49140
rect -15360 49020 -15350 49090
rect -15150 49020 -15140 49090
rect -15360 48980 -15140 49020
rect -15360 48910 -15350 48980
rect -15150 48910 -15140 48980
rect -15360 48860 -15140 48910
rect -14860 49090 -14640 49140
rect -14860 49020 -14850 49090
rect -14650 49020 -14640 49090
rect -14860 48980 -14640 49020
rect -14860 48910 -14850 48980
rect -14650 48910 -14640 48980
rect -14860 48860 -14640 48910
rect -14360 49090 -14140 49140
rect -14360 49020 -14350 49090
rect -14150 49020 -14140 49090
rect -14360 48980 -14140 49020
rect -14360 48910 -14350 48980
rect -14150 48910 -14140 48980
rect -14360 48860 -14140 48910
rect -13860 49090 -13640 49140
rect -13860 49020 -13850 49090
rect -13650 49020 -13640 49090
rect -13860 48980 -13640 49020
rect -13860 48910 -13850 48980
rect -13650 48910 -13640 48980
rect -13860 48860 -13640 48910
rect -13360 49090 -13140 49140
rect -13360 49020 -13350 49090
rect -13150 49020 -13140 49090
rect -13360 48980 -13140 49020
rect -13360 48910 -13350 48980
rect -13150 48910 -13140 48980
rect -13360 48860 -13140 48910
rect -12860 49090 -12640 49140
rect -12860 49020 -12850 49090
rect -12650 49020 -12640 49090
rect -12860 48980 -12640 49020
rect -12860 48910 -12850 48980
rect -12650 48910 -12640 48980
rect -12860 48860 -12640 48910
rect -12360 49090 -12140 49140
rect -12360 49020 -12350 49090
rect -12150 49020 -12140 49090
rect -12360 48980 -12140 49020
rect -12360 48910 -12350 48980
rect -12150 48910 -12140 48980
rect -12360 48860 -12140 48910
rect -16000 48850 -12000 48860
rect -16000 48650 -15980 48850
rect -15910 48650 -15590 48850
rect -15520 48650 -15480 48850
rect -15410 48650 -15090 48850
rect -15020 48650 -14980 48850
rect -14910 48650 -14590 48850
rect -14520 48650 -14480 48850
rect -14410 48650 -14090 48850
rect -14020 48650 -13980 48850
rect -13910 48650 -13590 48850
rect -13520 48650 -13480 48850
rect -13410 48650 -13090 48850
rect -13020 48650 -12980 48850
rect -12910 48650 -12590 48850
rect -12520 48650 -12480 48850
rect -12410 48650 -12090 48850
rect -12020 48650 -12000 48850
rect -16000 48640 -12000 48650
rect -15860 48590 -15640 48640
rect -15860 48520 -15850 48590
rect -15650 48520 -15640 48590
rect -15860 48480 -15640 48520
rect -15860 48410 -15850 48480
rect -15650 48410 -15640 48480
rect -15860 48360 -15640 48410
rect -15360 48590 -15140 48640
rect -15360 48520 -15350 48590
rect -15150 48520 -15140 48590
rect -15360 48480 -15140 48520
rect -15360 48410 -15350 48480
rect -15150 48410 -15140 48480
rect -15360 48360 -15140 48410
rect -14860 48590 -14640 48640
rect -14860 48520 -14850 48590
rect -14650 48520 -14640 48590
rect -14860 48480 -14640 48520
rect -14860 48410 -14850 48480
rect -14650 48410 -14640 48480
rect -14860 48360 -14640 48410
rect -14360 48590 -14140 48640
rect -14360 48520 -14350 48590
rect -14150 48520 -14140 48590
rect -14360 48480 -14140 48520
rect -14360 48410 -14350 48480
rect -14150 48410 -14140 48480
rect -14360 48360 -14140 48410
rect -13860 48590 -13640 48640
rect -13860 48520 -13850 48590
rect -13650 48520 -13640 48590
rect -13860 48480 -13640 48520
rect -13860 48410 -13850 48480
rect -13650 48410 -13640 48480
rect -13860 48360 -13640 48410
rect -13360 48590 -13140 48640
rect -13360 48520 -13350 48590
rect -13150 48520 -13140 48590
rect -13360 48480 -13140 48520
rect -13360 48410 -13350 48480
rect -13150 48410 -13140 48480
rect -13360 48360 -13140 48410
rect -12860 48590 -12640 48640
rect -12860 48520 -12850 48590
rect -12650 48520 -12640 48590
rect -12860 48480 -12640 48520
rect -12860 48410 -12850 48480
rect -12650 48410 -12640 48480
rect -12860 48360 -12640 48410
rect -12360 48590 -12140 48640
rect -12360 48520 -12350 48590
rect -12150 48520 -12140 48590
rect -12360 48480 -12140 48520
rect -12360 48410 -12350 48480
rect -12150 48410 -12140 48480
rect -12360 48360 -12140 48410
rect -16000 48350 -12000 48360
rect -16000 48150 -15980 48350
rect -15910 48150 -15590 48350
rect -15520 48150 -15480 48350
rect -15410 48150 -15090 48350
rect -15020 48150 -14980 48350
rect -14910 48150 -14590 48350
rect -14520 48150 -14480 48350
rect -14410 48150 -14090 48350
rect -14020 48150 -13980 48350
rect -13910 48150 -13590 48350
rect -13520 48150 -13480 48350
rect -13410 48150 -13090 48350
rect -13020 48150 -12980 48350
rect -12910 48150 -12590 48350
rect -12520 48150 -12480 48350
rect -12410 48150 -12090 48350
rect -12020 48150 -12000 48350
rect -16000 48140 -12000 48150
rect -15860 48090 -15640 48140
rect -15860 48020 -15850 48090
rect -15650 48020 -15640 48090
rect -15860 47980 -15640 48020
rect -15860 47910 -15850 47980
rect -15650 47910 -15640 47980
rect -15860 47860 -15640 47910
rect -15360 48090 -15140 48140
rect -15360 48020 -15350 48090
rect -15150 48020 -15140 48090
rect -15360 47980 -15140 48020
rect -15360 47910 -15350 47980
rect -15150 47910 -15140 47980
rect -15360 47860 -15140 47910
rect -14860 48090 -14640 48140
rect -14860 48020 -14850 48090
rect -14650 48020 -14640 48090
rect -14860 47980 -14640 48020
rect -14860 47910 -14850 47980
rect -14650 47910 -14640 47980
rect -14860 47860 -14640 47910
rect -14360 48090 -14140 48140
rect -14360 48020 -14350 48090
rect -14150 48020 -14140 48090
rect -14360 47980 -14140 48020
rect -14360 47910 -14350 47980
rect -14150 47910 -14140 47980
rect -14360 47860 -14140 47910
rect -13860 48090 -13640 48140
rect -13860 48020 -13850 48090
rect -13650 48020 -13640 48090
rect -13860 47980 -13640 48020
rect -13860 47910 -13850 47980
rect -13650 47910 -13640 47980
rect -13860 47860 -13640 47910
rect -13360 48090 -13140 48140
rect -13360 48020 -13350 48090
rect -13150 48020 -13140 48090
rect -13360 47980 -13140 48020
rect -13360 47910 -13350 47980
rect -13150 47910 -13140 47980
rect -13360 47860 -13140 47910
rect -12860 48090 -12640 48140
rect -12860 48020 -12850 48090
rect -12650 48020 -12640 48090
rect -12860 47980 -12640 48020
rect -12860 47910 -12850 47980
rect -12650 47910 -12640 47980
rect -12860 47860 -12640 47910
rect -12360 48090 -12140 48140
rect -12360 48020 -12350 48090
rect -12150 48020 -12140 48090
rect -12360 47980 -12140 48020
rect -12360 47910 -12350 47980
rect -12150 47910 -12140 47980
rect -12360 47860 -12140 47910
rect -16000 47850 -12000 47860
rect -16000 47650 -15980 47850
rect -15910 47650 -15590 47850
rect -15520 47650 -15480 47850
rect -15410 47650 -15090 47850
rect -15020 47650 -14980 47850
rect -14910 47650 -14590 47850
rect -14520 47650 -14480 47850
rect -14410 47650 -14090 47850
rect -14020 47650 -13980 47850
rect -13910 47650 -13590 47850
rect -13520 47650 -13480 47850
rect -13410 47650 -13090 47850
rect -13020 47650 -12980 47850
rect -12910 47650 -12590 47850
rect -12520 47650 -12480 47850
rect -12410 47650 -12090 47850
rect -12020 47650 -12000 47850
rect -16000 47640 -12000 47650
rect -15860 47590 -15640 47640
rect -15860 47520 -15850 47590
rect -15650 47520 -15640 47590
rect -15860 47480 -15640 47520
rect -15860 47410 -15850 47480
rect -15650 47410 -15640 47480
rect -15860 47360 -15640 47410
rect -15360 47590 -15140 47640
rect -15360 47520 -15350 47590
rect -15150 47520 -15140 47590
rect -15360 47480 -15140 47520
rect -15360 47410 -15350 47480
rect -15150 47410 -15140 47480
rect -15360 47360 -15140 47410
rect -14860 47590 -14640 47640
rect -14860 47520 -14850 47590
rect -14650 47520 -14640 47590
rect -14860 47480 -14640 47520
rect -14860 47410 -14850 47480
rect -14650 47410 -14640 47480
rect -14860 47360 -14640 47410
rect -14360 47590 -14140 47640
rect -14360 47520 -14350 47590
rect -14150 47520 -14140 47590
rect -14360 47480 -14140 47520
rect -14360 47410 -14350 47480
rect -14150 47410 -14140 47480
rect -14360 47360 -14140 47410
rect -13860 47590 -13640 47640
rect -13860 47520 -13850 47590
rect -13650 47520 -13640 47590
rect -13860 47480 -13640 47520
rect -13860 47410 -13850 47480
rect -13650 47410 -13640 47480
rect -13860 47360 -13640 47410
rect -13360 47590 -13140 47640
rect -13360 47520 -13350 47590
rect -13150 47520 -13140 47590
rect -13360 47480 -13140 47520
rect -13360 47410 -13350 47480
rect -13150 47410 -13140 47480
rect -13360 47360 -13140 47410
rect -12860 47590 -12640 47640
rect -12860 47520 -12850 47590
rect -12650 47520 -12640 47590
rect -12860 47480 -12640 47520
rect -12860 47410 -12850 47480
rect -12650 47410 -12640 47480
rect -12860 47360 -12640 47410
rect -12360 47590 -12140 47640
rect -12360 47520 -12350 47590
rect -12150 47520 -12140 47590
rect -12360 47480 -12140 47520
rect -12360 47410 -12350 47480
rect -12150 47410 -12140 47480
rect -12360 47360 -12140 47410
rect -16000 47350 -12000 47360
rect -16000 47150 -15980 47350
rect -15910 47150 -15590 47350
rect -15520 47150 -15480 47350
rect -15410 47150 -15090 47350
rect -15020 47150 -14980 47350
rect -14910 47150 -14590 47350
rect -14520 47150 -14480 47350
rect -14410 47150 -14090 47350
rect -14020 47150 -13980 47350
rect -13910 47150 -13590 47350
rect -13520 47150 -13480 47350
rect -13410 47150 -13090 47350
rect -13020 47150 -12980 47350
rect -12910 47150 -12590 47350
rect -12520 47150 -12480 47350
rect -12410 47150 -12090 47350
rect -12020 47150 -12000 47350
rect -16000 47140 -12000 47150
rect -15860 47090 -15640 47140
rect -15860 47020 -15850 47090
rect -15650 47020 -15640 47090
rect -15860 46980 -15640 47020
rect -15860 46910 -15850 46980
rect -15650 46910 -15640 46980
rect -15860 46860 -15640 46910
rect -15360 47090 -15140 47140
rect -15360 47020 -15350 47090
rect -15150 47020 -15140 47090
rect -15360 46980 -15140 47020
rect -15360 46910 -15350 46980
rect -15150 46910 -15140 46980
rect -15360 46860 -15140 46910
rect -14860 47090 -14640 47140
rect -14860 47020 -14850 47090
rect -14650 47020 -14640 47090
rect -14860 46980 -14640 47020
rect -14860 46910 -14850 46980
rect -14650 46910 -14640 46980
rect -14860 46860 -14640 46910
rect -14360 47090 -14140 47140
rect -14360 47020 -14350 47090
rect -14150 47020 -14140 47090
rect -14360 46980 -14140 47020
rect -14360 46910 -14350 46980
rect -14150 46910 -14140 46980
rect -14360 46860 -14140 46910
rect -13860 47090 -13640 47140
rect -13860 47020 -13850 47090
rect -13650 47020 -13640 47090
rect -13860 46980 -13640 47020
rect -13860 46910 -13850 46980
rect -13650 46910 -13640 46980
rect -13860 46860 -13640 46910
rect -13360 47090 -13140 47140
rect -13360 47020 -13350 47090
rect -13150 47020 -13140 47090
rect -13360 46980 -13140 47020
rect -13360 46910 -13350 46980
rect -13150 46910 -13140 46980
rect -13360 46860 -13140 46910
rect -12860 47090 -12640 47140
rect -12860 47020 -12850 47090
rect -12650 47020 -12640 47090
rect -12860 46980 -12640 47020
rect -12860 46910 -12850 46980
rect -12650 46910 -12640 46980
rect -12860 46860 -12640 46910
rect -12360 47090 -12140 47140
rect -12360 47020 -12350 47090
rect -12150 47020 -12140 47090
rect -12360 46980 -12140 47020
rect -12360 46910 -12350 46980
rect -12150 46910 -12140 46980
rect -12360 46860 -12140 46910
rect -16000 46850 -12000 46860
rect -16000 46650 -15980 46850
rect -15910 46650 -15590 46850
rect -15520 46650 -15480 46850
rect -15410 46650 -15090 46850
rect -15020 46650 -14980 46850
rect -14910 46650 -14590 46850
rect -14520 46650 -14480 46850
rect -14410 46650 -14090 46850
rect -14020 46650 -13980 46850
rect -13910 46650 -13590 46850
rect -13520 46650 -13480 46850
rect -13410 46650 -13090 46850
rect -13020 46650 -12980 46850
rect -12910 46650 -12590 46850
rect -12520 46650 -12480 46850
rect -12410 46650 -12090 46850
rect -12020 46650 -12000 46850
rect -16000 46640 -12000 46650
rect -15860 46590 -15640 46640
rect -15860 46520 -15850 46590
rect -15650 46520 -15640 46590
rect -15860 46480 -15640 46520
rect -15860 46410 -15850 46480
rect -15650 46410 -15640 46480
rect -15860 46360 -15640 46410
rect -15360 46590 -15140 46640
rect -15360 46520 -15350 46590
rect -15150 46520 -15140 46590
rect -15360 46480 -15140 46520
rect -15360 46410 -15350 46480
rect -15150 46410 -15140 46480
rect -15360 46360 -15140 46410
rect -14860 46590 -14640 46640
rect -14860 46520 -14850 46590
rect -14650 46520 -14640 46590
rect -14860 46480 -14640 46520
rect -14860 46410 -14850 46480
rect -14650 46410 -14640 46480
rect -14860 46360 -14640 46410
rect -14360 46590 -14140 46640
rect -14360 46520 -14350 46590
rect -14150 46520 -14140 46590
rect -14360 46480 -14140 46520
rect -14360 46410 -14350 46480
rect -14150 46410 -14140 46480
rect -14360 46360 -14140 46410
rect -13860 46590 -13640 46640
rect -13860 46520 -13850 46590
rect -13650 46520 -13640 46590
rect -13860 46480 -13640 46520
rect -13860 46410 -13850 46480
rect -13650 46410 -13640 46480
rect -13860 46360 -13640 46410
rect -13360 46590 -13140 46640
rect -13360 46520 -13350 46590
rect -13150 46520 -13140 46590
rect -13360 46480 -13140 46520
rect -13360 46410 -13350 46480
rect -13150 46410 -13140 46480
rect -13360 46360 -13140 46410
rect -12860 46590 -12640 46640
rect -12860 46520 -12850 46590
rect -12650 46520 -12640 46590
rect -12860 46480 -12640 46520
rect -12860 46410 -12850 46480
rect -12650 46410 -12640 46480
rect -12860 46360 -12640 46410
rect -12360 46590 -12140 46640
rect -12360 46520 -12350 46590
rect -12150 46520 -12140 46590
rect -12360 46480 -12140 46520
rect -12360 46410 -12350 46480
rect -12150 46410 -12140 46480
rect -12360 46360 -12140 46410
rect -16000 46350 -12000 46360
rect -16000 46150 -15980 46350
rect -15910 46150 -15590 46350
rect -15520 46150 -15480 46350
rect -15410 46150 -15090 46350
rect -15020 46150 -14980 46350
rect -14910 46150 -14590 46350
rect -14520 46150 -14480 46350
rect -14410 46150 -14090 46350
rect -14020 46150 -13980 46350
rect -13910 46150 -13590 46350
rect -13520 46150 -13480 46350
rect -13410 46150 -13090 46350
rect -13020 46150 -12980 46350
rect -12910 46150 -12590 46350
rect -12520 46150 -12480 46350
rect -12410 46150 -12090 46350
rect -12020 46150 -12000 46350
rect -16000 46140 -12000 46150
rect -15860 46090 -15640 46140
rect -15860 46020 -15850 46090
rect -15650 46020 -15640 46090
rect -15860 45980 -15640 46020
rect -15860 45910 -15850 45980
rect -15650 45910 -15640 45980
rect -15860 45860 -15640 45910
rect -15360 46090 -15140 46140
rect -15360 46020 -15350 46090
rect -15150 46020 -15140 46090
rect -15360 45980 -15140 46020
rect -15360 45910 -15350 45980
rect -15150 45910 -15140 45980
rect -15360 45860 -15140 45910
rect -14860 46090 -14640 46140
rect -14860 46020 -14850 46090
rect -14650 46020 -14640 46090
rect -14860 45980 -14640 46020
rect -14860 45910 -14850 45980
rect -14650 45910 -14640 45980
rect -14860 45860 -14640 45910
rect -14360 46090 -14140 46140
rect -14360 46020 -14350 46090
rect -14150 46020 -14140 46090
rect -14360 45980 -14140 46020
rect -14360 45910 -14350 45980
rect -14150 45910 -14140 45980
rect -14360 45860 -14140 45910
rect -13860 46090 -13640 46140
rect -13860 46020 -13850 46090
rect -13650 46020 -13640 46090
rect -13860 45980 -13640 46020
rect -13860 45910 -13850 45980
rect -13650 45910 -13640 45980
rect -13860 45860 -13640 45910
rect -13360 46090 -13140 46140
rect -13360 46020 -13350 46090
rect -13150 46020 -13140 46090
rect -13360 45980 -13140 46020
rect -13360 45910 -13350 45980
rect -13150 45910 -13140 45980
rect -13360 45860 -13140 45910
rect -12860 46090 -12640 46140
rect -12860 46020 -12850 46090
rect -12650 46020 -12640 46090
rect -12860 45980 -12640 46020
rect -12860 45910 -12850 45980
rect -12650 45910 -12640 45980
rect -12860 45860 -12640 45910
rect -12360 46090 -12140 46140
rect -12360 46020 -12350 46090
rect -12150 46020 -12140 46090
rect -12360 45980 -12140 46020
rect -12360 45910 -12350 45980
rect -12150 45910 -12140 45980
rect -12360 45860 -12140 45910
rect -16000 45850 -12000 45860
rect -16000 45650 -15980 45850
rect -15910 45650 -15590 45850
rect -15520 45650 -15480 45850
rect -15410 45650 -15090 45850
rect -15020 45650 -14980 45850
rect -14910 45650 -14590 45850
rect -14520 45650 -14480 45850
rect -14410 45650 -14090 45850
rect -14020 45650 -13980 45850
rect -13910 45650 -13590 45850
rect -13520 45650 -13480 45850
rect -13410 45650 -13090 45850
rect -13020 45650 -12980 45850
rect -12910 45650 -12590 45850
rect -12520 45650 -12480 45850
rect -12410 45650 -12090 45850
rect -12020 45650 -12000 45850
rect -16000 45640 -12000 45650
rect -15860 45590 -15640 45640
rect -15860 45520 -15850 45590
rect -15650 45520 -15640 45590
rect -15860 45480 -15640 45520
rect -15860 45410 -15850 45480
rect -15650 45410 -15640 45480
rect -15860 45360 -15640 45410
rect -15360 45590 -15140 45640
rect -15360 45520 -15350 45590
rect -15150 45520 -15140 45590
rect -15360 45480 -15140 45520
rect -15360 45410 -15350 45480
rect -15150 45410 -15140 45480
rect -15360 45360 -15140 45410
rect -14860 45590 -14640 45640
rect -14860 45520 -14850 45590
rect -14650 45520 -14640 45590
rect -14860 45480 -14640 45520
rect -14860 45410 -14850 45480
rect -14650 45410 -14640 45480
rect -14860 45360 -14640 45410
rect -14360 45590 -14140 45640
rect -14360 45520 -14350 45590
rect -14150 45520 -14140 45590
rect -14360 45480 -14140 45520
rect -14360 45410 -14350 45480
rect -14150 45410 -14140 45480
rect -14360 45360 -14140 45410
rect -13860 45590 -13640 45640
rect -13860 45520 -13850 45590
rect -13650 45520 -13640 45590
rect -13860 45480 -13640 45520
rect -13860 45410 -13850 45480
rect -13650 45410 -13640 45480
rect -13860 45360 -13640 45410
rect -13360 45590 -13140 45640
rect -13360 45520 -13350 45590
rect -13150 45520 -13140 45590
rect -13360 45480 -13140 45520
rect -13360 45410 -13350 45480
rect -13150 45410 -13140 45480
rect -13360 45360 -13140 45410
rect -12860 45590 -12640 45640
rect -12860 45520 -12850 45590
rect -12650 45520 -12640 45590
rect -12860 45480 -12640 45520
rect -12860 45410 -12850 45480
rect -12650 45410 -12640 45480
rect -12860 45360 -12640 45410
rect -12360 45590 -12140 45640
rect -12360 45520 -12350 45590
rect -12150 45520 -12140 45590
rect -12360 45480 -12140 45520
rect -12360 45410 -12350 45480
rect -12150 45410 -12140 45480
rect -12360 45360 -12140 45410
rect -16000 45350 -12000 45360
rect -16000 45150 -15980 45350
rect -15910 45150 -15590 45350
rect -15520 45150 -15480 45350
rect -15410 45150 -15090 45350
rect -15020 45150 -14980 45350
rect -14910 45150 -14590 45350
rect -14520 45150 -14480 45350
rect -14410 45150 -14090 45350
rect -14020 45150 -13980 45350
rect -13910 45150 -13590 45350
rect -13520 45150 -13480 45350
rect -13410 45150 -13090 45350
rect -13020 45150 -12980 45350
rect -12910 45150 -12590 45350
rect -12520 45150 -12480 45350
rect -12410 45150 -12090 45350
rect -12020 45150 -12000 45350
rect -16000 45140 -12000 45150
rect -15860 45090 -15640 45140
rect -15860 45020 -15850 45090
rect -15650 45020 -15640 45090
rect -15860 44980 -15640 45020
rect -15860 44910 -15850 44980
rect -15650 44910 -15640 44980
rect -15860 44860 -15640 44910
rect -15360 45090 -15140 45140
rect -15360 45020 -15350 45090
rect -15150 45020 -15140 45090
rect -15360 44980 -15140 45020
rect -15360 44910 -15350 44980
rect -15150 44910 -15140 44980
rect -15360 44860 -15140 44910
rect -14860 45090 -14640 45140
rect -14860 45020 -14850 45090
rect -14650 45020 -14640 45090
rect -14860 44980 -14640 45020
rect -14860 44910 -14850 44980
rect -14650 44910 -14640 44980
rect -14860 44860 -14640 44910
rect -14360 45090 -14140 45140
rect -14360 45020 -14350 45090
rect -14150 45020 -14140 45090
rect -14360 44980 -14140 45020
rect -14360 44910 -14350 44980
rect -14150 44910 -14140 44980
rect -14360 44860 -14140 44910
rect -13860 45090 -13640 45140
rect -13860 45020 -13850 45090
rect -13650 45020 -13640 45090
rect -13860 44980 -13640 45020
rect -13860 44910 -13850 44980
rect -13650 44910 -13640 44980
rect -13860 44860 -13640 44910
rect -13360 45090 -13140 45140
rect -13360 45020 -13350 45090
rect -13150 45020 -13140 45090
rect -13360 44980 -13140 45020
rect -13360 44910 -13350 44980
rect -13150 44910 -13140 44980
rect -13360 44860 -13140 44910
rect -12860 45090 -12640 45140
rect -12860 45020 -12850 45090
rect -12650 45020 -12640 45090
rect -12860 44980 -12640 45020
rect -12860 44910 -12850 44980
rect -12650 44910 -12640 44980
rect -12860 44860 -12640 44910
rect -12360 45090 -12140 45140
rect -12360 45020 -12350 45090
rect -12150 45020 -12140 45090
rect -12360 44980 -12140 45020
rect -12360 44910 -12350 44980
rect -12150 44910 -12140 44980
rect -12360 44860 -12140 44910
rect -16000 44850 -12000 44860
rect -16000 44650 -15980 44850
rect -15910 44650 -15590 44850
rect -15520 44650 -15480 44850
rect -15410 44650 -15090 44850
rect -15020 44650 -14980 44850
rect -14910 44650 -14590 44850
rect -14520 44650 -14480 44850
rect -14410 44650 -14090 44850
rect -14020 44650 -13980 44850
rect -13910 44650 -13590 44850
rect -13520 44650 -13480 44850
rect -13410 44650 -13090 44850
rect -13020 44650 -12980 44850
rect -12910 44650 -12590 44850
rect -12520 44650 -12480 44850
rect -12410 44650 -12090 44850
rect -12020 44650 -12000 44850
rect -16000 44640 -12000 44650
rect -15860 44590 -15640 44640
rect -15860 44520 -15850 44590
rect -15650 44520 -15640 44590
rect -15860 44480 -15640 44520
rect -15860 44410 -15850 44480
rect -15650 44410 -15640 44480
rect -15860 44360 -15640 44410
rect -15360 44590 -15140 44640
rect -15360 44520 -15350 44590
rect -15150 44520 -15140 44590
rect -15360 44480 -15140 44520
rect -15360 44410 -15350 44480
rect -15150 44410 -15140 44480
rect -15360 44360 -15140 44410
rect -14860 44590 -14640 44640
rect -14860 44520 -14850 44590
rect -14650 44520 -14640 44590
rect -14860 44480 -14640 44520
rect -14860 44410 -14850 44480
rect -14650 44410 -14640 44480
rect -14860 44360 -14640 44410
rect -14360 44590 -14140 44640
rect -14360 44520 -14350 44590
rect -14150 44520 -14140 44590
rect -14360 44480 -14140 44520
rect -14360 44410 -14350 44480
rect -14150 44410 -14140 44480
rect -14360 44360 -14140 44410
rect -13860 44590 -13640 44640
rect -13860 44520 -13850 44590
rect -13650 44520 -13640 44590
rect -13860 44480 -13640 44520
rect -13860 44410 -13850 44480
rect -13650 44410 -13640 44480
rect -13860 44360 -13640 44410
rect -13360 44590 -13140 44640
rect -13360 44520 -13350 44590
rect -13150 44520 -13140 44590
rect -13360 44480 -13140 44520
rect -13360 44410 -13350 44480
rect -13150 44410 -13140 44480
rect -13360 44360 -13140 44410
rect -12860 44590 -12640 44640
rect -12860 44520 -12850 44590
rect -12650 44520 -12640 44590
rect -12860 44480 -12640 44520
rect -12860 44410 -12850 44480
rect -12650 44410 -12640 44480
rect -12860 44360 -12640 44410
rect -12360 44590 -12140 44640
rect -12360 44520 -12350 44590
rect -12150 44520 -12140 44590
rect -12360 44480 -12140 44520
rect -12360 44410 -12350 44480
rect -12150 44410 -12140 44480
rect -12360 44360 -12140 44410
rect -16000 44350 -12000 44360
rect -16000 44150 -15980 44350
rect -15910 44150 -15590 44350
rect -15520 44150 -15480 44350
rect -15410 44150 -15090 44350
rect -15020 44150 -14980 44350
rect -14910 44150 -14590 44350
rect -14520 44150 -14480 44350
rect -14410 44150 -14090 44350
rect -14020 44150 -13980 44350
rect -13910 44150 -13590 44350
rect -13520 44150 -13480 44350
rect -13410 44150 -13090 44350
rect -13020 44150 -12980 44350
rect -12910 44150 -12590 44350
rect -12520 44150 -12480 44350
rect -12410 44150 -12090 44350
rect -12020 44150 -12000 44350
rect -16000 44140 -12000 44150
rect -15860 44090 -15640 44140
rect -15860 44020 -15850 44090
rect -15650 44020 -15640 44090
rect -15860 43980 -15640 44020
rect -15860 43910 -15850 43980
rect -15650 43910 -15640 43980
rect -15860 43860 -15640 43910
rect -15360 44090 -15140 44140
rect -15360 44020 -15350 44090
rect -15150 44020 -15140 44090
rect -15360 43980 -15140 44020
rect -15360 43910 -15350 43980
rect -15150 43910 -15140 43980
rect -15360 43860 -15140 43910
rect -14860 44090 -14640 44140
rect -14860 44020 -14850 44090
rect -14650 44020 -14640 44090
rect -14860 43980 -14640 44020
rect -14860 43910 -14850 43980
rect -14650 43910 -14640 43980
rect -14860 43860 -14640 43910
rect -14360 44090 -14140 44140
rect -14360 44020 -14350 44090
rect -14150 44020 -14140 44090
rect -14360 43980 -14140 44020
rect -14360 43910 -14350 43980
rect -14150 43910 -14140 43980
rect -14360 43860 -14140 43910
rect -13860 44090 -13640 44140
rect -13860 44020 -13850 44090
rect -13650 44020 -13640 44090
rect -13860 43980 -13640 44020
rect -13860 43910 -13850 43980
rect -13650 43910 -13640 43980
rect -13860 43860 -13640 43910
rect -13360 44090 -13140 44140
rect -13360 44020 -13350 44090
rect -13150 44020 -13140 44090
rect -13360 43980 -13140 44020
rect -13360 43910 -13350 43980
rect -13150 43910 -13140 43980
rect -13360 43860 -13140 43910
rect -12860 44090 -12640 44140
rect -12860 44020 -12850 44090
rect -12650 44020 -12640 44090
rect -12860 43980 -12640 44020
rect -12860 43910 -12850 43980
rect -12650 43910 -12640 43980
rect -12860 43860 -12640 43910
rect -12360 44090 -12140 44140
rect -12360 44020 -12350 44090
rect -12150 44020 -12140 44090
rect -12360 43980 -12140 44020
rect -12360 43910 -12350 43980
rect -12150 43910 -12140 43980
rect -12360 43860 -12140 43910
rect -16000 43850 -12000 43860
rect -16000 43650 -15980 43850
rect -15910 43650 -15590 43850
rect -15520 43650 -15480 43850
rect -15410 43650 -15090 43850
rect -15020 43650 -14980 43850
rect -14910 43650 -14590 43850
rect -14520 43650 -14480 43850
rect -14410 43650 -14090 43850
rect -14020 43650 -13980 43850
rect -13910 43650 -13590 43850
rect -13520 43650 -13480 43850
rect -13410 43650 -13090 43850
rect -13020 43650 -12980 43850
rect -12910 43650 -12590 43850
rect -12520 43650 -12480 43850
rect -12410 43650 -12090 43850
rect -12020 43650 -12000 43850
rect -16000 43640 -12000 43650
rect -15860 43590 -15640 43640
rect -15860 43520 -15850 43590
rect -15650 43520 -15640 43590
rect -15860 43480 -15640 43520
rect -15860 43410 -15850 43480
rect -15650 43410 -15640 43480
rect -15860 43360 -15640 43410
rect -15360 43590 -15140 43640
rect -15360 43520 -15350 43590
rect -15150 43520 -15140 43590
rect -15360 43480 -15140 43520
rect -15360 43410 -15350 43480
rect -15150 43410 -15140 43480
rect -15360 43360 -15140 43410
rect -14860 43590 -14640 43640
rect -14860 43520 -14850 43590
rect -14650 43520 -14640 43590
rect -14860 43480 -14640 43520
rect -14860 43410 -14850 43480
rect -14650 43410 -14640 43480
rect -14860 43360 -14640 43410
rect -14360 43590 -14140 43640
rect -14360 43520 -14350 43590
rect -14150 43520 -14140 43590
rect -14360 43480 -14140 43520
rect -14360 43410 -14350 43480
rect -14150 43410 -14140 43480
rect -14360 43360 -14140 43410
rect -13860 43590 -13640 43640
rect -13860 43520 -13850 43590
rect -13650 43520 -13640 43590
rect -13860 43480 -13640 43520
rect -13860 43410 -13850 43480
rect -13650 43410 -13640 43480
rect -13860 43360 -13640 43410
rect -13360 43590 -13140 43640
rect -13360 43520 -13350 43590
rect -13150 43520 -13140 43590
rect -13360 43480 -13140 43520
rect -13360 43410 -13350 43480
rect -13150 43410 -13140 43480
rect -13360 43360 -13140 43410
rect -12860 43590 -12640 43640
rect -12860 43520 -12850 43590
rect -12650 43520 -12640 43590
rect -12860 43480 -12640 43520
rect -12860 43410 -12850 43480
rect -12650 43410 -12640 43480
rect -12860 43360 -12640 43410
rect -12360 43590 -12140 43640
rect -12360 43520 -12350 43590
rect -12150 43520 -12140 43590
rect -12360 43480 -12140 43520
rect -12360 43410 -12350 43480
rect -12150 43410 -12140 43480
rect -12360 43360 -12140 43410
rect -16000 43350 -12000 43360
rect -16000 43150 -15980 43350
rect -15910 43150 -15590 43350
rect -15520 43150 -15480 43350
rect -15410 43150 -15090 43350
rect -15020 43150 -14980 43350
rect -14910 43150 -14590 43350
rect -14520 43150 -14480 43350
rect -14410 43150 -14090 43350
rect -14020 43150 -13980 43350
rect -13910 43150 -13590 43350
rect -13520 43150 -13480 43350
rect -13410 43150 -13090 43350
rect -13020 43150 -12980 43350
rect -12910 43150 -12590 43350
rect -12520 43150 -12480 43350
rect -12410 43150 -12090 43350
rect -12020 43150 -12000 43350
rect -16000 43140 -12000 43150
rect -15860 43090 -15640 43140
rect -15860 43020 -15850 43090
rect -15650 43020 -15640 43090
rect -15860 42980 -15640 43020
rect -15860 42910 -15850 42980
rect -15650 42910 -15640 42980
rect -15860 42860 -15640 42910
rect -15360 43090 -15140 43140
rect -15360 43020 -15350 43090
rect -15150 43020 -15140 43090
rect -15360 42980 -15140 43020
rect -15360 42910 -15350 42980
rect -15150 42910 -15140 42980
rect -15360 42860 -15140 42910
rect -14860 43090 -14640 43140
rect -14860 43020 -14850 43090
rect -14650 43020 -14640 43090
rect -14860 42980 -14640 43020
rect -14860 42910 -14850 42980
rect -14650 42910 -14640 42980
rect -14860 42860 -14640 42910
rect -14360 43090 -14140 43140
rect -14360 43020 -14350 43090
rect -14150 43020 -14140 43090
rect -14360 42980 -14140 43020
rect -14360 42910 -14350 42980
rect -14150 42910 -14140 42980
rect -14360 42860 -14140 42910
rect -13860 43090 -13640 43140
rect -13860 43020 -13850 43090
rect -13650 43020 -13640 43090
rect -13860 42980 -13640 43020
rect -13860 42910 -13850 42980
rect -13650 42910 -13640 42980
rect -13860 42860 -13640 42910
rect -13360 43090 -13140 43140
rect -13360 43020 -13350 43090
rect -13150 43020 -13140 43090
rect -13360 42980 -13140 43020
rect -13360 42910 -13350 42980
rect -13150 42910 -13140 42980
rect -13360 42860 -13140 42910
rect -12860 43090 -12640 43140
rect -12860 43020 -12850 43090
rect -12650 43020 -12640 43090
rect -12860 42980 -12640 43020
rect -12860 42910 -12850 42980
rect -12650 42910 -12640 42980
rect -12860 42860 -12640 42910
rect -12360 43090 -12140 43140
rect -12360 43020 -12350 43090
rect -12150 43020 -12140 43090
rect -12360 42980 -12140 43020
rect -12360 42910 -12350 42980
rect -12150 42910 -12140 42980
rect -12360 42860 -12140 42910
rect -16000 42850 -12000 42860
rect -16000 42650 -15980 42850
rect -15910 42650 -15590 42850
rect -15520 42650 -15480 42850
rect -15410 42650 -15090 42850
rect -15020 42650 -14980 42850
rect -14910 42650 -14590 42850
rect -14520 42650 -14480 42850
rect -14410 42650 -14090 42850
rect -14020 42650 -13980 42850
rect -13910 42650 -13590 42850
rect -13520 42650 -13480 42850
rect -13410 42650 -13090 42850
rect -13020 42650 -12980 42850
rect -12910 42650 -12590 42850
rect -12520 42650 -12480 42850
rect -12410 42650 -12090 42850
rect -12020 42650 -12000 42850
rect -16000 42640 -12000 42650
rect -15860 42590 -15640 42640
rect -15860 42520 -15850 42590
rect -15650 42520 -15640 42590
rect -15860 42480 -15640 42520
rect -15860 42410 -15850 42480
rect -15650 42410 -15640 42480
rect -15860 42360 -15640 42410
rect -15360 42590 -15140 42640
rect -15360 42520 -15350 42590
rect -15150 42520 -15140 42590
rect -15360 42480 -15140 42520
rect -15360 42410 -15350 42480
rect -15150 42410 -15140 42480
rect -15360 42360 -15140 42410
rect -14860 42590 -14640 42640
rect -14860 42520 -14850 42590
rect -14650 42520 -14640 42590
rect -14860 42480 -14640 42520
rect -14860 42410 -14850 42480
rect -14650 42410 -14640 42480
rect -14860 42360 -14640 42410
rect -14360 42590 -14140 42640
rect -14360 42520 -14350 42590
rect -14150 42520 -14140 42590
rect -14360 42480 -14140 42520
rect -14360 42410 -14350 42480
rect -14150 42410 -14140 42480
rect -14360 42360 -14140 42410
rect -13860 42590 -13640 42640
rect -13860 42520 -13850 42590
rect -13650 42520 -13640 42590
rect -13860 42480 -13640 42520
rect -13860 42410 -13850 42480
rect -13650 42410 -13640 42480
rect -13860 42360 -13640 42410
rect -13360 42590 -13140 42640
rect -13360 42520 -13350 42590
rect -13150 42520 -13140 42590
rect -13360 42480 -13140 42520
rect -13360 42410 -13350 42480
rect -13150 42410 -13140 42480
rect -13360 42360 -13140 42410
rect -12860 42590 -12640 42640
rect -12860 42520 -12850 42590
rect -12650 42520 -12640 42590
rect -12860 42480 -12640 42520
rect -12860 42410 -12850 42480
rect -12650 42410 -12640 42480
rect -12860 42360 -12640 42410
rect -12360 42590 -12140 42640
rect -12360 42520 -12350 42590
rect -12150 42520 -12140 42590
rect -12360 42480 -12140 42520
rect -12360 42410 -12350 42480
rect -12150 42410 -12140 42480
rect -12360 42360 -12140 42410
rect -16000 42350 -12000 42360
rect -16000 42150 -15980 42350
rect -15910 42150 -15590 42350
rect -15520 42150 -15480 42350
rect -15410 42150 -15090 42350
rect -15020 42150 -14980 42350
rect -14910 42150 -14590 42350
rect -14520 42150 -14480 42350
rect -14410 42150 -14090 42350
rect -14020 42150 -13980 42350
rect -13910 42150 -13590 42350
rect -13520 42150 -13480 42350
rect -13410 42150 -13090 42350
rect -13020 42150 -12980 42350
rect -12910 42150 -12590 42350
rect -12520 42150 -12480 42350
rect -12410 42150 -12090 42350
rect -12020 42150 -12000 42350
rect -16000 42140 -12000 42150
rect -15860 42090 -15640 42140
rect -15860 42020 -15850 42090
rect -15650 42020 -15640 42090
rect -15860 41980 -15640 42020
rect -15860 41910 -15850 41980
rect -15650 41910 -15640 41980
rect -15860 41860 -15640 41910
rect -15360 42090 -15140 42140
rect -15360 42020 -15350 42090
rect -15150 42020 -15140 42090
rect -15360 41980 -15140 42020
rect -15360 41910 -15350 41980
rect -15150 41910 -15140 41980
rect -15360 41860 -15140 41910
rect -14860 42090 -14640 42140
rect -14860 42020 -14850 42090
rect -14650 42020 -14640 42090
rect -14860 41980 -14640 42020
rect -14860 41910 -14850 41980
rect -14650 41910 -14640 41980
rect -14860 41860 -14640 41910
rect -14360 42090 -14140 42140
rect -14360 42020 -14350 42090
rect -14150 42020 -14140 42090
rect -14360 41980 -14140 42020
rect -14360 41910 -14350 41980
rect -14150 41910 -14140 41980
rect -14360 41860 -14140 41910
rect -13860 42090 -13640 42140
rect -13860 42020 -13850 42090
rect -13650 42020 -13640 42090
rect -13860 41980 -13640 42020
rect -13860 41910 -13850 41980
rect -13650 41910 -13640 41980
rect -13860 41860 -13640 41910
rect -13360 42090 -13140 42140
rect -13360 42020 -13350 42090
rect -13150 42020 -13140 42090
rect -13360 41980 -13140 42020
rect -13360 41910 -13350 41980
rect -13150 41910 -13140 41980
rect -13360 41860 -13140 41910
rect -12860 42090 -12640 42140
rect -12860 42020 -12850 42090
rect -12650 42020 -12640 42090
rect -12860 41980 -12640 42020
rect -12860 41910 -12850 41980
rect -12650 41910 -12640 41980
rect -12860 41860 -12640 41910
rect -12360 42090 -12140 42140
rect -12360 42020 -12350 42090
rect -12150 42020 -12140 42090
rect -12360 41980 -12140 42020
rect -12360 41910 -12350 41980
rect -12150 41910 -12140 41980
rect -12360 41860 -12140 41910
rect -11860 41980 -11640 42000
rect -11860 41910 -11850 41980
rect -11650 41910 -11640 41980
rect -11860 41860 -11640 41910
rect -11360 41980 -11140 42000
rect -11360 41910 -11350 41980
rect -11150 41910 -11140 41980
rect -11360 41860 -11140 41910
rect -10860 41980 -10640 42000
rect -10860 41910 -10850 41980
rect -10650 41910 -10640 41980
rect -10860 41860 -10640 41910
rect -10360 41980 -10140 42000
rect -10360 41910 -10350 41980
rect -10150 41910 -10140 41980
rect -10360 41860 -10140 41910
rect -9860 41980 -9640 42000
rect -9860 41910 -9850 41980
rect -9650 41910 -9640 41980
rect -9860 41860 -9640 41910
rect -9360 41980 -9140 42000
rect -9360 41910 -9350 41980
rect -9150 41910 -9140 41980
rect -9360 41860 -9140 41910
rect -8860 41980 -8640 42000
rect -8860 41910 -8850 41980
rect -8650 41910 -8640 41980
rect -8860 41860 -8640 41910
rect -8360 41980 -8140 42000
rect -8360 41910 -8350 41980
rect -8150 41910 -8140 41980
rect -8360 41860 -8140 41910
rect -7860 41980 -7640 42000
rect -7860 41910 -7850 41980
rect -7650 41910 -7640 41980
rect -7860 41860 -7640 41910
rect -7360 41980 -7140 42000
rect -7360 41910 -7350 41980
rect -7150 41910 -7140 41980
rect -7360 41860 -7140 41910
rect -6860 41980 -6640 42000
rect -6860 41910 -6850 41980
rect -6650 41910 -6640 41980
rect -6860 41860 -6640 41910
rect -6360 41980 -6140 42000
rect -6360 41910 -6350 41980
rect -6150 41910 -6140 41980
rect -6360 41860 -6140 41910
rect -5860 41980 -5640 42000
rect -5860 41910 -5850 41980
rect -5650 41910 -5640 41980
rect -5860 41860 -5640 41910
rect -5360 41980 -5140 42000
rect -5360 41910 -5350 41980
rect -5150 41910 -5140 41980
rect -5360 41860 -5140 41910
rect -4860 41980 -4640 42000
rect -4860 41910 -4850 41980
rect -4650 41910 -4640 41980
rect -4860 41860 -4640 41910
rect -4360 41980 -4140 42000
rect -4360 41910 -4350 41980
rect -4150 41910 -4140 41980
rect -4360 41860 -4140 41910
rect -3860 41980 -3640 42000
rect -3860 41910 -3850 41980
rect -3650 41910 -3640 41980
rect -3860 41860 -3640 41910
rect -3360 41980 -3140 42000
rect -3360 41910 -3350 41980
rect -3150 41910 -3140 41980
rect -3360 41860 -3140 41910
rect -2860 41980 -2640 42000
rect -2860 41910 -2850 41980
rect -2650 41910 -2640 41980
rect -2860 41860 -2640 41910
rect -2360 41980 -2140 42000
rect -2360 41910 -2350 41980
rect -2150 41910 -2140 41980
rect -2360 41860 -2140 41910
rect -1860 41980 -1640 42000
rect -1860 41910 -1850 41980
rect -1650 41910 -1640 41980
rect -1860 41860 -1640 41910
rect -1360 41980 -1140 42000
rect -1360 41910 -1350 41980
rect -1150 41910 -1140 41980
rect -1360 41860 -1140 41910
rect -860 41980 -640 42000
rect -860 41910 -850 41980
rect -650 41910 -640 41980
rect -860 41860 -640 41910
rect -360 41980 -140 42000
rect -360 41910 -350 41980
rect -150 41910 -140 41980
rect -360 41860 -140 41910
rect 140 41980 360 42000
rect 140 41910 150 41980
rect 350 41910 360 41980
rect 140 41860 360 41910
rect 640 41980 860 42000
rect 640 41910 650 41980
rect 850 41910 860 41980
rect 640 41860 860 41910
rect 1140 41980 1360 42000
rect 1140 41910 1150 41980
rect 1350 41910 1360 41980
rect 1140 41860 1360 41910
rect 1640 41980 1860 42000
rect 1640 41910 1650 41980
rect 1850 41910 1860 41980
rect 1640 41860 1860 41910
rect 2140 41980 2360 42000
rect 2140 41910 2150 41980
rect 2350 41910 2360 41980
rect 2140 41860 2360 41910
rect 2640 41980 2860 42000
rect 2640 41910 2650 41980
rect 2850 41910 2860 41980
rect 2640 41860 2860 41910
rect 3140 41980 3360 42000
rect 3140 41910 3150 41980
rect 3350 41910 3360 41980
rect 3140 41860 3360 41910
rect 3640 41980 3860 42000
rect 3640 41910 3650 41980
rect 3850 41910 3860 41980
rect 3640 41860 3860 41910
rect -16000 41850 4000 41860
rect -16000 41650 -15980 41850
rect -15910 41650 -15590 41850
rect -15520 41650 -15480 41850
rect -15410 41650 -15090 41850
rect -15020 41650 -14980 41850
rect -14910 41650 -14590 41850
rect -14520 41650 -14480 41850
rect -14410 41650 -14090 41850
rect -14020 41650 -13980 41850
rect -13910 41650 -13590 41850
rect -13520 41650 -13480 41850
rect -13410 41650 -13090 41850
rect -13020 41650 -12980 41850
rect -12910 41650 -12590 41850
rect -12520 41650 -12480 41850
rect -12410 41650 -12090 41850
rect -12020 41650 -11980 41850
rect -11910 41650 -11590 41850
rect -11520 41650 -11480 41850
rect -11410 41650 -11090 41850
rect -11020 41650 -10980 41850
rect -10910 41650 -10590 41850
rect -10520 41650 -10480 41850
rect -10410 41650 -10090 41850
rect -10020 41650 -9980 41850
rect -9910 41650 -9590 41850
rect -9520 41650 -9480 41850
rect -9410 41650 -9090 41850
rect -9020 41650 -8980 41850
rect -8910 41650 -8590 41850
rect -8520 41650 -8480 41850
rect -8410 41650 -8090 41850
rect -8020 41650 -7980 41850
rect -7910 41650 -7590 41850
rect -7520 41650 -7480 41850
rect -7410 41650 -7090 41850
rect -7020 41650 -6980 41850
rect -6910 41650 -6590 41850
rect -6520 41650 -6480 41850
rect -6410 41650 -6090 41850
rect -6020 41650 -5980 41850
rect -5910 41650 -5590 41850
rect -5520 41650 -5480 41850
rect -5410 41650 -5090 41850
rect -5020 41650 -4980 41850
rect -4910 41650 -4590 41850
rect -4520 41650 -4480 41850
rect -4410 41650 -4090 41850
rect -4020 41650 -3980 41850
rect -3910 41650 -3590 41850
rect -3520 41650 -3480 41850
rect -3410 41650 -3090 41850
rect -3020 41650 -2980 41850
rect -2910 41650 -2590 41850
rect -2520 41650 -2480 41850
rect -2410 41650 -2090 41850
rect -2020 41650 -1980 41850
rect -1910 41650 -1590 41850
rect -1520 41650 -1480 41850
rect -1410 41650 -1090 41850
rect -1020 41650 -980 41850
rect -910 41650 -590 41850
rect -520 41650 -480 41850
rect -410 41650 -90 41850
rect -20 41650 20 41850
rect 90 41650 410 41850
rect 480 41650 520 41850
rect 590 41650 910 41850
rect 980 41650 1020 41850
rect 1090 41650 1410 41850
rect 1480 41650 1520 41850
rect 1590 41650 1910 41850
rect 1980 41650 2020 41850
rect 2090 41650 2410 41850
rect 2480 41650 2520 41850
rect 2590 41650 2910 41850
rect 2980 41650 3020 41850
rect 3090 41650 3410 41850
rect 3480 41650 3520 41850
rect 3590 41650 3910 41850
rect 3980 41650 4000 41850
rect -16000 41640 4000 41650
rect -15860 41590 -15640 41640
rect -15860 41520 -15850 41590
rect -15650 41520 -15640 41590
rect -15860 41480 -15640 41520
rect -15860 41410 -15850 41480
rect -15650 41410 -15640 41480
rect -15860 41360 -15640 41410
rect -15360 41590 -15140 41640
rect -15360 41520 -15350 41590
rect -15150 41520 -15140 41590
rect -15360 41480 -15140 41520
rect -15360 41410 -15350 41480
rect -15150 41410 -15140 41480
rect -15360 41360 -15140 41410
rect -14860 41590 -14640 41640
rect -14860 41520 -14850 41590
rect -14650 41520 -14640 41590
rect -14860 41480 -14640 41520
rect -14860 41410 -14850 41480
rect -14650 41410 -14640 41480
rect -14860 41360 -14640 41410
rect -14360 41590 -14140 41640
rect -14360 41520 -14350 41590
rect -14150 41520 -14140 41590
rect -14360 41480 -14140 41520
rect -14360 41410 -14350 41480
rect -14150 41410 -14140 41480
rect -14360 41360 -14140 41410
rect -13860 41590 -13640 41640
rect -13860 41520 -13850 41590
rect -13650 41520 -13640 41590
rect -13860 41480 -13640 41520
rect -13860 41410 -13850 41480
rect -13650 41410 -13640 41480
rect -13860 41360 -13640 41410
rect -13360 41590 -13140 41640
rect -13360 41520 -13350 41590
rect -13150 41520 -13140 41590
rect -13360 41480 -13140 41520
rect -13360 41410 -13350 41480
rect -13150 41410 -13140 41480
rect -13360 41360 -13140 41410
rect -12860 41590 -12640 41640
rect -12860 41520 -12850 41590
rect -12650 41520 -12640 41590
rect -12860 41480 -12640 41520
rect -12860 41410 -12850 41480
rect -12650 41410 -12640 41480
rect -12860 41360 -12640 41410
rect -12360 41590 -12140 41640
rect -12360 41520 -12350 41590
rect -12150 41520 -12140 41590
rect -12360 41480 -12140 41520
rect -12360 41410 -12350 41480
rect -12150 41410 -12140 41480
rect -12360 41360 -12140 41410
rect -11860 41590 -11640 41640
rect -11860 41520 -11850 41590
rect -11650 41520 -11640 41590
rect -11860 41480 -11640 41520
rect -11860 41410 -11850 41480
rect -11650 41410 -11640 41480
rect -11860 41360 -11640 41410
rect -11360 41590 -11140 41640
rect -11360 41520 -11350 41590
rect -11150 41520 -11140 41590
rect -11360 41480 -11140 41520
rect -11360 41410 -11350 41480
rect -11150 41410 -11140 41480
rect -11360 41360 -11140 41410
rect -10860 41590 -10640 41640
rect -10860 41520 -10850 41590
rect -10650 41520 -10640 41590
rect -10860 41480 -10640 41520
rect -10860 41410 -10850 41480
rect -10650 41410 -10640 41480
rect -10860 41360 -10640 41410
rect -10360 41590 -10140 41640
rect -10360 41520 -10350 41590
rect -10150 41520 -10140 41590
rect -10360 41480 -10140 41520
rect -10360 41410 -10350 41480
rect -10150 41410 -10140 41480
rect -10360 41360 -10140 41410
rect -9860 41590 -9640 41640
rect -9860 41520 -9850 41590
rect -9650 41520 -9640 41590
rect -9860 41480 -9640 41520
rect -9860 41410 -9850 41480
rect -9650 41410 -9640 41480
rect -9860 41360 -9640 41410
rect -9360 41590 -9140 41640
rect -9360 41520 -9350 41590
rect -9150 41520 -9140 41590
rect -9360 41480 -9140 41520
rect -9360 41410 -9350 41480
rect -9150 41410 -9140 41480
rect -9360 41360 -9140 41410
rect -8860 41590 -8640 41640
rect -8860 41520 -8850 41590
rect -8650 41520 -8640 41590
rect -8860 41480 -8640 41520
rect -8860 41410 -8850 41480
rect -8650 41410 -8640 41480
rect -8860 41360 -8640 41410
rect -8360 41590 -8140 41640
rect -8360 41520 -8350 41590
rect -8150 41520 -8140 41590
rect -8360 41480 -8140 41520
rect -8360 41410 -8350 41480
rect -8150 41410 -8140 41480
rect -8360 41360 -8140 41410
rect -7860 41590 -7640 41640
rect -7860 41520 -7850 41590
rect -7650 41520 -7640 41590
rect -7860 41480 -7640 41520
rect -7860 41410 -7850 41480
rect -7650 41410 -7640 41480
rect -7860 41360 -7640 41410
rect -7360 41590 -7140 41640
rect -7360 41520 -7350 41590
rect -7150 41520 -7140 41590
rect -7360 41480 -7140 41520
rect -7360 41410 -7350 41480
rect -7150 41410 -7140 41480
rect -7360 41360 -7140 41410
rect -6860 41590 -6640 41640
rect -6860 41520 -6850 41590
rect -6650 41520 -6640 41590
rect -6860 41480 -6640 41520
rect -6860 41410 -6850 41480
rect -6650 41410 -6640 41480
rect -6860 41360 -6640 41410
rect -6360 41590 -6140 41640
rect -6360 41520 -6350 41590
rect -6150 41520 -6140 41590
rect -6360 41480 -6140 41520
rect -6360 41410 -6350 41480
rect -6150 41410 -6140 41480
rect -6360 41360 -6140 41410
rect -5860 41590 -5640 41640
rect -5860 41520 -5850 41590
rect -5650 41520 -5640 41590
rect -5860 41480 -5640 41520
rect -5860 41410 -5850 41480
rect -5650 41410 -5640 41480
rect -5860 41360 -5640 41410
rect -5360 41590 -5140 41640
rect -5360 41520 -5350 41590
rect -5150 41520 -5140 41590
rect -5360 41480 -5140 41520
rect -5360 41410 -5350 41480
rect -5150 41410 -5140 41480
rect -5360 41360 -5140 41410
rect -4860 41590 -4640 41640
rect -4860 41520 -4850 41590
rect -4650 41520 -4640 41590
rect -4860 41480 -4640 41520
rect -4860 41410 -4850 41480
rect -4650 41410 -4640 41480
rect -4860 41360 -4640 41410
rect -4360 41590 -4140 41640
rect -4360 41520 -4350 41590
rect -4150 41520 -4140 41590
rect -4360 41480 -4140 41520
rect -4360 41410 -4350 41480
rect -4150 41410 -4140 41480
rect -4360 41360 -4140 41410
rect -3860 41590 -3640 41640
rect -3860 41520 -3850 41590
rect -3650 41520 -3640 41590
rect -3860 41480 -3640 41520
rect -3860 41410 -3850 41480
rect -3650 41410 -3640 41480
rect -3860 41360 -3640 41410
rect -3360 41590 -3140 41640
rect -3360 41520 -3350 41590
rect -3150 41520 -3140 41590
rect -3360 41480 -3140 41520
rect -3360 41410 -3350 41480
rect -3150 41410 -3140 41480
rect -3360 41360 -3140 41410
rect -2860 41590 -2640 41640
rect -2860 41520 -2850 41590
rect -2650 41520 -2640 41590
rect -2860 41480 -2640 41520
rect -2860 41410 -2850 41480
rect -2650 41410 -2640 41480
rect -2860 41360 -2640 41410
rect -2360 41590 -2140 41640
rect -2360 41520 -2350 41590
rect -2150 41520 -2140 41590
rect -2360 41480 -2140 41520
rect -2360 41410 -2350 41480
rect -2150 41410 -2140 41480
rect -2360 41360 -2140 41410
rect -1860 41590 -1640 41640
rect -1860 41520 -1850 41590
rect -1650 41520 -1640 41590
rect -1860 41480 -1640 41520
rect -1860 41410 -1850 41480
rect -1650 41410 -1640 41480
rect -1860 41360 -1640 41410
rect -1360 41590 -1140 41640
rect -1360 41520 -1350 41590
rect -1150 41520 -1140 41590
rect -1360 41480 -1140 41520
rect -1360 41410 -1350 41480
rect -1150 41410 -1140 41480
rect -1360 41360 -1140 41410
rect -860 41590 -640 41640
rect -860 41520 -850 41590
rect -650 41520 -640 41590
rect -860 41480 -640 41520
rect -860 41410 -850 41480
rect -650 41410 -640 41480
rect -860 41360 -640 41410
rect -360 41590 -140 41640
rect -360 41520 -350 41590
rect -150 41520 -140 41590
rect -360 41480 -140 41520
rect -360 41410 -350 41480
rect -150 41410 -140 41480
rect -360 41360 -140 41410
rect 140 41590 360 41640
rect 140 41520 150 41590
rect 350 41520 360 41590
rect 140 41480 360 41520
rect 140 41410 150 41480
rect 350 41410 360 41480
rect 140 41360 360 41410
rect 640 41590 860 41640
rect 640 41520 650 41590
rect 850 41520 860 41590
rect 640 41480 860 41520
rect 640 41410 650 41480
rect 850 41410 860 41480
rect 640 41360 860 41410
rect 1140 41590 1360 41640
rect 1140 41520 1150 41590
rect 1350 41520 1360 41590
rect 1140 41480 1360 41520
rect 1140 41410 1150 41480
rect 1350 41410 1360 41480
rect 1140 41360 1360 41410
rect 1640 41590 1860 41640
rect 1640 41520 1650 41590
rect 1850 41520 1860 41590
rect 1640 41480 1860 41520
rect 1640 41410 1650 41480
rect 1850 41410 1860 41480
rect 1640 41360 1860 41410
rect 2140 41590 2360 41640
rect 2140 41520 2150 41590
rect 2350 41520 2360 41590
rect 2140 41480 2360 41520
rect 2140 41410 2150 41480
rect 2350 41410 2360 41480
rect 2140 41360 2360 41410
rect 2640 41590 2860 41640
rect 2640 41520 2650 41590
rect 2850 41520 2860 41590
rect 2640 41480 2860 41520
rect 2640 41410 2650 41480
rect 2850 41410 2860 41480
rect 2640 41360 2860 41410
rect 3140 41590 3360 41640
rect 3140 41520 3150 41590
rect 3350 41520 3360 41590
rect 3140 41480 3360 41520
rect 3140 41410 3150 41480
rect 3350 41410 3360 41480
rect 3140 41360 3360 41410
rect 3640 41590 3860 41640
rect 3640 41520 3650 41590
rect 3850 41520 3860 41590
rect 3640 41480 3860 41520
rect 3640 41410 3650 41480
rect 3850 41410 3860 41480
rect 3640 41360 3860 41410
rect -16000 41350 4000 41360
rect -16000 41150 -15980 41350
rect -15910 41150 -15590 41350
rect -15520 41150 -15480 41350
rect -15410 41150 -15090 41350
rect -15020 41150 -14980 41350
rect -14910 41150 -14590 41350
rect -14520 41150 -14480 41350
rect -14410 41150 -14090 41350
rect -14020 41150 -13980 41350
rect -13910 41150 -13590 41350
rect -13520 41150 -13480 41350
rect -13410 41150 -13090 41350
rect -13020 41150 -12980 41350
rect -12910 41150 -12590 41350
rect -12520 41150 -12480 41350
rect -12410 41150 -12090 41350
rect -12020 41150 -11980 41350
rect -11910 41150 -11590 41350
rect -11520 41150 -11480 41350
rect -11410 41150 -11090 41350
rect -11020 41150 -10980 41350
rect -10910 41150 -10590 41350
rect -10520 41150 -10480 41350
rect -10410 41150 -10090 41350
rect -10020 41150 -9980 41350
rect -9910 41150 -9590 41350
rect -9520 41150 -9480 41350
rect -9410 41150 -9090 41350
rect -9020 41150 -8980 41350
rect -8910 41150 -8590 41350
rect -8520 41150 -8480 41350
rect -8410 41150 -8090 41350
rect -8020 41150 -7980 41350
rect -7910 41150 -7590 41350
rect -7520 41150 -7480 41350
rect -7410 41150 -7090 41350
rect -7020 41150 -6980 41350
rect -6910 41150 -6590 41350
rect -6520 41150 -6480 41350
rect -6410 41150 -6090 41350
rect -6020 41150 -5980 41350
rect -5910 41150 -5590 41350
rect -5520 41150 -5480 41350
rect -5410 41150 -5090 41350
rect -5020 41150 -4980 41350
rect -4910 41150 -4590 41350
rect -4520 41150 -4480 41350
rect -4410 41150 -4090 41350
rect -4020 41150 -3980 41350
rect -3910 41150 -3590 41350
rect -3520 41150 -3480 41350
rect -3410 41150 -3090 41350
rect -3020 41150 -2980 41350
rect -2910 41150 -2590 41350
rect -2520 41150 -2480 41350
rect -2410 41150 -2090 41350
rect -2020 41150 -1980 41350
rect -1910 41150 -1590 41350
rect -1520 41150 -1480 41350
rect -1410 41150 -1090 41350
rect -1020 41150 -980 41350
rect -910 41150 -590 41350
rect -520 41150 -480 41350
rect -410 41150 -90 41350
rect -20 41150 20 41350
rect 90 41150 410 41350
rect 480 41150 520 41350
rect 590 41150 910 41350
rect 980 41150 1020 41350
rect 1090 41150 1410 41350
rect 1480 41150 1520 41350
rect 1590 41150 1910 41350
rect 1980 41150 2020 41350
rect 2090 41150 2410 41350
rect 2480 41150 2520 41350
rect 2590 41150 2910 41350
rect 2980 41150 3020 41350
rect 3090 41150 3410 41350
rect 3480 41150 3520 41350
rect 3590 41150 3910 41350
rect 3980 41150 4000 41350
rect -16000 41140 4000 41150
rect -15860 41090 -15640 41140
rect -15860 41020 -15850 41090
rect -15650 41020 -15640 41090
rect -15860 40980 -15640 41020
rect -15860 40910 -15850 40980
rect -15650 40910 -15640 40980
rect -15860 40860 -15640 40910
rect -15360 41090 -15140 41140
rect -15360 41020 -15350 41090
rect -15150 41020 -15140 41090
rect -15360 40980 -15140 41020
rect -15360 40910 -15350 40980
rect -15150 40910 -15140 40980
rect -15360 40860 -15140 40910
rect -14860 41090 -14640 41140
rect -14860 41020 -14850 41090
rect -14650 41020 -14640 41090
rect -14860 40980 -14640 41020
rect -14860 40910 -14850 40980
rect -14650 40910 -14640 40980
rect -14860 40860 -14640 40910
rect -14360 41090 -14140 41140
rect -14360 41020 -14350 41090
rect -14150 41020 -14140 41090
rect -14360 40980 -14140 41020
rect -14360 40910 -14350 40980
rect -14150 40910 -14140 40980
rect -14360 40860 -14140 40910
rect -13860 41090 -13640 41140
rect -13860 41020 -13850 41090
rect -13650 41020 -13640 41090
rect -13860 40980 -13640 41020
rect -13860 40910 -13850 40980
rect -13650 40910 -13640 40980
rect -13860 40860 -13640 40910
rect -13360 41090 -13140 41140
rect -13360 41020 -13350 41090
rect -13150 41020 -13140 41090
rect -13360 40980 -13140 41020
rect -13360 40910 -13350 40980
rect -13150 40910 -13140 40980
rect -13360 40860 -13140 40910
rect -12860 41090 -12640 41140
rect -12860 41020 -12850 41090
rect -12650 41020 -12640 41090
rect -12860 40980 -12640 41020
rect -12860 40910 -12850 40980
rect -12650 40910 -12640 40980
rect -12860 40860 -12640 40910
rect -12360 41090 -12140 41140
rect -12360 41020 -12350 41090
rect -12150 41020 -12140 41090
rect -12360 40980 -12140 41020
rect -12360 40910 -12350 40980
rect -12150 40910 -12140 40980
rect -12360 40860 -12140 40910
rect -11860 41090 -11640 41140
rect -11860 41020 -11850 41090
rect -11650 41020 -11640 41090
rect -11860 40980 -11640 41020
rect -11860 40910 -11850 40980
rect -11650 40910 -11640 40980
rect -11860 40860 -11640 40910
rect -11360 41090 -11140 41140
rect -11360 41020 -11350 41090
rect -11150 41020 -11140 41090
rect -11360 40980 -11140 41020
rect -11360 40910 -11350 40980
rect -11150 40910 -11140 40980
rect -11360 40860 -11140 40910
rect -10860 41090 -10640 41140
rect -10860 41020 -10850 41090
rect -10650 41020 -10640 41090
rect -10860 40980 -10640 41020
rect -10860 40910 -10850 40980
rect -10650 40910 -10640 40980
rect -10860 40860 -10640 40910
rect -10360 41090 -10140 41140
rect -10360 41020 -10350 41090
rect -10150 41020 -10140 41090
rect -10360 40980 -10140 41020
rect -10360 40910 -10350 40980
rect -10150 40910 -10140 40980
rect -10360 40860 -10140 40910
rect -9860 41090 -9640 41140
rect -9860 41020 -9850 41090
rect -9650 41020 -9640 41090
rect -9860 40980 -9640 41020
rect -9860 40910 -9850 40980
rect -9650 40910 -9640 40980
rect -9860 40860 -9640 40910
rect -9360 41090 -9140 41140
rect -9360 41020 -9350 41090
rect -9150 41020 -9140 41090
rect -9360 40980 -9140 41020
rect -9360 40910 -9350 40980
rect -9150 40910 -9140 40980
rect -9360 40860 -9140 40910
rect -8860 41090 -8640 41140
rect -8860 41020 -8850 41090
rect -8650 41020 -8640 41090
rect -8860 40980 -8640 41020
rect -8860 40910 -8850 40980
rect -8650 40910 -8640 40980
rect -8860 40860 -8640 40910
rect -8360 41090 -8140 41140
rect -8360 41020 -8350 41090
rect -8150 41020 -8140 41090
rect -8360 40980 -8140 41020
rect -8360 40910 -8350 40980
rect -8150 40910 -8140 40980
rect -8360 40860 -8140 40910
rect -7860 41090 -7640 41140
rect -7860 41020 -7850 41090
rect -7650 41020 -7640 41090
rect -7860 40980 -7640 41020
rect -7860 40910 -7850 40980
rect -7650 40910 -7640 40980
rect -7860 40860 -7640 40910
rect -7360 41090 -7140 41140
rect -7360 41020 -7350 41090
rect -7150 41020 -7140 41090
rect -7360 40980 -7140 41020
rect -7360 40910 -7350 40980
rect -7150 40910 -7140 40980
rect -7360 40860 -7140 40910
rect -6860 41090 -6640 41140
rect -6860 41020 -6850 41090
rect -6650 41020 -6640 41090
rect -6860 40980 -6640 41020
rect -6860 40910 -6850 40980
rect -6650 40910 -6640 40980
rect -6860 40860 -6640 40910
rect -6360 41090 -6140 41140
rect -6360 41020 -6350 41090
rect -6150 41020 -6140 41090
rect -6360 40980 -6140 41020
rect -6360 40910 -6350 40980
rect -6150 40910 -6140 40980
rect -6360 40860 -6140 40910
rect -5860 41090 -5640 41140
rect -5860 41020 -5850 41090
rect -5650 41020 -5640 41090
rect -5860 40980 -5640 41020
rect -5860 40910 -5850 40980
rect -5650 40910 -5640 40980
rect -5860 40860 -5640 40910
rect -5360 41090 -5140 41140
rect -5360 41020 -5350 41090
rect -5150 41020 -5140 41090
rect -5360 40980 -5140 41020
rect -5360 40910 -5350 40980
rect -5150 40910 -5140 40980
rect -5360 40860 -5140 40910
rect -4860 41090 -4640 41140
rect -4860 41020 -4850 41090
rect -4650 41020 -4640 41090
rect -4860 40980 -4640 41020
rect -4860 40910 -4850 40980
rect -4650 40910 -4640 40980
rect -4860 40860 -4640 40910
rect -4360 41090 -4140 41140
rect -4360 41020 -4350 41090
rect -4150 41020 -4140 41090
rect -4360 40980 -4140 41020
rect -4360 40910 -4350 40980
rect -4150 40910 -4140 40980
rect -4360 40860 -4140 40910
rect -3860 41090 -3640 41140
rect -3860 41020 -3850 41090
rect -3650 41020 -3640 41090
rect -3860 40980 -3640 41020
rect -3860 40910 -3850 40980
rect -3650 40910 -3640 40980
rect -3860 40860 -3640 40910
rect -3360 41090 -3140 41140
rect -3360 41020 -3350 41090
rect -3150 41020 -3140 41090
rect -3360 40980 -3140 41020
rect -3360 40910 -3350 40980
rect -3150 40910 -3140 40980
rect -3360 40860 -3140 40910
rect -2860 41090 -2640 41140
rect -2860 41020 -2850 41090
rect -2650 41020 -2640 41090
rect -2860 40980 -2640 41020
rect -2860 40910 -2850 40980
rect -2650 40910 -2640 40980
rect -2860 40860 -2640 40910
rect -2360 41090 -2140 41140
rect -2360 41020 -2350 41090
rect -2150 41020 -2140 41090
rect -2360 40980 -2140 41020
rect -2360 40910 -2350 40980
rect -2150 40910 -2140 40980
rect -2360 40860 -2140 40910
rect -1860 41090 -1640 41140
rect -1860 41020 -1850 41090
rect -1650 41020 -1640 41090
rect -1860 40980 -1640 41020
rect -1860 40910 -1850 40980
rect -1650 40910 -1640 40980
rect -1860 40860 -1640 40910
rect -1360 41090 -1140 41140
rect -1360 41020 -1350 41090
rect -1150 41020 -1140 41090
rect -1360 40980 -1140 41020
rect -1360 40910 -1350 40980
rect -1150 40910 -1140 40980
rect -1360 40860 -1140 40910
rect -860 41090 -640 41140
rect -860 41020 -850 41090
rect -650 41020 -640 41090
rect -860 40980 -640 41020
rect -860 40910 -850 40980
rect -650 40910 -640 40980
rect -860 40860 -640 40910
rect -360 41090 -140 41140
rect -360 41020 -350 41090
rect -150 41020 -140 41090
rect -360 40980 -140 41020
rect -360 40910 -350 40980
rect -150 40910 -140 40980
rect -360 40860 -140 40910
rect 140 41090 360 41140
rect 140 41020 150 41090
rect 350 41020 360 41090
rect 140 40980 360 41020
rect 140 40910 150 40980
rect 350 40910 360 40980
rect 140 40860 360 40910
rect 640 41090 860 41140
rect 640 41020 650 41090
rect 850 41020 860 41090
rect 640 40980 860 41020
rect 640 40910 650 40980
rect 850 40910 860 40980
rect 640 40860 860 40910
rect 1140 41090 1360 41140
rect 1140 41020 1150 41090
rect 1350 41020 1360 41090
rect 1140 40980 1360 41020
rect 1140 40910 1150 40980
rect 1350 40910 1360 40980
rect 1140 40860 1360 40910
rect 1640 41090 1860 41140
rect 1640 41020 1650 41090
rect 1850 41020 1860 41090
rect 1640 40980 1860 41020
rect 1640 40910 1650 40980
rect 1850 40910 1860 40980
rect 1640 40860 1860 40910
rect 2140 41090 2360 41140
rect 2140 41020 2150 41090
rect 2350 41020 2360 41090
rect 2140 40980 2360 41020
rect 2140 40910 2150 40980
rect 2350 40910 2360 40980
rect 2140 40860 2360 40910
rect 2640 41090 2860 41140
rect 2640 41020 2650 41090
rect 2850 41020 2860 41090
rect 2640 40980 2860 41020
rect 2640 40910 2650 40980
rect 2850 40910 2860 40980
rect 2640 40860 2860 40910
rect 3140 41090 3360 41140
rect 3140 41020 3150 41090
rect 3350 41020 3360 41090
rect 3140 40980 3360 41020
rect 3140 40910 3150 40980
rect 3350 40910 3360 40980
rect 3140 40860 3360 40910
rect 3640 41090 3860 41140
rect 3640 41020 3650 41090
rect 3850 41020 3860 41090
rect 3640 40980 3860 41020
rect 3640 40910 3650 40980
rect 3850 40910 3860 40980
rect 3640 40860 3860 40910
rect -16000 40850 4000 40860
rect -16000 40650 -15980 40850
rect -15910 40650 -15590 40850
rect -15520 40650 -15480 40850
rect -15410 40650 -15090 40850
rect -15020 40650 -14980 40850
rect -14910 40650 -14590 40850
rect -14520 40650 -14480 40850
rect -14410 40650 -14090 40850
rect -14020 40650 -13980 40850
rect -13910 40650 -13590 40850
rect -13520 40650 -13480 40850
rect -13410 40650 -13090 40850
rect -13020 40650 -12980 40850
rect -12910 40650 -12590 40850
rect -12520 40650 -12480 40850
rect -12410 40650 -12090 40850
rect -12020 40650 -11980 40850
rect -11910 40650 -11590 40850
rect -11520 40650 -11480 40850
rect -11410 40650 -11090 40850
rect -11020 40650 -10980 40850
rect -10910 40650 -10590 40850
rect -10520 40650 -10480 40850
rect -10410 40650 -10090 40850
rect -10020 40650 -9980 40850
rect -9910 40650 -9590 40850
rect -9520 40650 -9480 40850
rect -9410 40650 -9090 40850
rect -9020 40650 -8980 40850
rect -8910 40650 -8590 40850
rect -8520 40650 -8480 40850
rect -8410 40650 -8090 40850
rect -8020 40650 -7980 40850
rect -7910 40650 -7590 40850
rect -7520 40650 -7480 40850
rect -7410 40650 -7090 40850
rect -7020 40650 -6980 40850
rect -6910 40650 -6590 40850
rect -6520 40650 -6480 40850
rect -6410 40650 -6090 40850
rect -6020 40650 -5980 40850
rect -5910 40650 -5590 40850
rect -5520 40650 -5480 40850
rect -5410 40650 -5090 40850
rect -5020 40650 -4980 40850
rect -4910 40650 -4590 40850
rect -4520 40650 -4480 40850
rect -4410 40650 -4090 40850
rect -4020 40650 -3980 40850
rect -3910 40650 -3590 40850
rect -3520 40650 -3480 40850
rect -3410 40650 -3090 40850
rect -3020 40650 -2980 40850
rect -2910 40650 -2590 40850
rect -2520 40650 -2480 40850
rect -2410 40650 -2090 40850
rect -2020 40650 -1980 40850
rect -1910 40650 -1590 40850
rect -1520 40650 -1480 40850
rect -1410 40650 -1090 40850
rect -1020 40650 -980 40850
rect -910 40650 -590 40850
rect -520 40650 -480 40850
rect -410 40650 -90 40850
rect -20 40650 20 40850
rect 90 40650 410 40850
rect 480 40650 520 40850
rect 590 40650 910 40850
rect 980 40650 1020 40850
rect 1090 40650 1410 40850
rect 1480 40650 1520 40850
rect 1590 40650 1910 40850
rect 1980 40650 2020 40850
rect 2090 40650 2410 40850
rect 2480 40650 2520 40850
rect 2590 40650 2910 40850
rect 2980 40650 3020 40850
rect 3090 40650 3410 40850
rect 3480 40650 3520 40850
rect 3590 40650 3910 40850
rect 3980 40650 4000 40850
rect -16000 40640 4000 40650
rect -15860 40590 -15640 40640
rect -15860 40520 -15850 40590
rect -15650 40520 -15640 40590
rect -15860 40480 -15640 40520
rect -15860 40410 -15850 40480
rect -15650 40410 -15640 40480
rect -15860 40360 -15640 40410
rect -15360 40590 -15140 40640
rect -15360 40520 -15350 40590
rect -15150 40520 -15140 40590
rect -15360 40480 -15140 40520
rect -15360 40410 -15350 40480
rect -15150 40410 -15140 40480
rect -15360 40360 -15140 40410
rect -14860 40590 -14640 40640
rect -14860 40520 -14850 40590
rect -14650 40520 -14640 40590
rect -14860 40480 -14640 40520
rect -14860 40410 -14850 40480
rect -14650 40410 -14640 40480
rect -14860 40360 -14640 40410
rect -14360 40590 -14140 40640
rect -14360 40520 -14350 40590
rect -14150 40520 -14140 40590
rect -14360 40480 -14140 40520
rect -14360 40410 -14350 40480
rect -14150 40410 -14140 40480
rect -14360 40360 -14140 40410
rect -13860 40590 -13640 40640
rect -13860 40520 -13850 40590
rect -13650 40520 -13640 40590
rect -13860 40480 -13640 40520
rect -13860 40410 -13850 40480
rect -13650 40410 -13640 40480
rect -13860 40360 -13640 40410
rect -13360 40590 -13140 40640
rect -13360 40520 -13350 40590
rect -13150 40520 -13140 40590
rect -13360 40480 -13140 40520
rect -13360 40410 -13350 40480
rect -13150 40410 -13140 40480
rect -13360 40360 -13140 40410
rect -12860 40590 -12640 40640
rect -12860 40520 -12850 40590
rect -12650 40520 -12640 40590
rect -12860 40480 -12640 40520
rect -12860 40410 -12850 40480
rect -12650 40410 -12640 40480
rect -12860 40360 -12640 40410
rect -12360 40590 -12140 40640
rect -12360 40520 -12350 40590
rect -12150 40520 -12140 40590
rect -12360 40480 -12140 40520
rect -12360 40410 -12350 40480
rect -12150 40410 -12140 40480
rect -12360 40360 -12140 40410
rect -11860 40590 -11640 40640
rect -11860 40520 -11850 40590
rect -11650 40520 -11640 40590
rect -11860 40480 -11640 40520
rect -11860 40410 -11850 40480
rect -11650 40410 -11640 40480
rect -11860 40360 -11640 40410
rect -11360 40590 -11140 40640
rect -11360 40520 -11350 40590
rect -11150 40520 -11140 40590
rect -11360 40480 -11140 40520
rect -11360 40410 -11350 40480
rect -11150 40410 -11140 40480
rect -11360 40360 -11140 40410
rect -10860 40590 -10640 40640
rect -10860 40520 -10850 40590
rect -10650 40520 -10640 40590
rect -10860 40480 -10640 40520
rect -10860 40410 -10850 40480
rect -10650 40410 -10640 40480
rect -10860 40360 -10640 40410
rect -10360 40590 -10140 40640
rect -10360 40520 -10350 40590
rect -10150 40520 -10140 40590
rect -10360 40480 -10140 40520
rect -10360 40410 -10350 40480
rect -10150 40410 -10140 40480
rect -10360 40360 -10140 40410
rect -9860 40590 -9640 40640
rect -9860 40520 -9850 40590
rect -9650 40520 -9640 40590
rect -9860 40480 -9640 40520
rect -9860 40410 -9850 40480
rect -9650 40410 -9640 40480
rect -9860 40360 -9640 40410
rect -9360 40590 -9140 40640
rect -9360 40520 -9350 40590
rect -9150 40520 -9140 40590
rect -9360 40480 -9140 40520
rect -9360 40410 -9350 40480
rect -9150 40410 -9140 40480
rect -9360 40360 -9140 40410
rect -8860 40590 -8640 40640
rect -8860 40520 -8850 40590
rect -8650 40520 -8640 40590
rect -8860 40480 -8640 40520
rect -8860 40410 -8850 40480
rect -8650 40410 -8640 40480
rect -8860 40360 -8640 40410
rect -8360 40590 -8140 40640
rect -8360 40520 -8350 40590
rect -8150 40520 -8140 40590
rect -8360 40480 -8140 40520
rect -8360 40410 -8350 40480
rect -8150 40410 -8140 40480
rect -8360 40360 -8140 40410
rect -7860 40590 -7640 40640
rect -7860 40520 -7850 40590
rect -7650 40520 -7640 40590
rect -7860 40480 -7640 40520
rect -7860 40410 -7850 40480
rect -7650 40410 -7640 40480
rect -7860 40360 -7640 40410
rect -7360 40590 -7140 40640
rect -7360 40520 -7350 40590
rect -7150 40520 -7140 40590
rect -7360 40480 -7140 40520
rect -7360 40410 -7350 40480
rect -7150 40410 -7140 40480
rect -7360 40360 -7140 40410
rect -6860 40590 -6640 40640
rect -6860 40520 -6850 40590
rect -6650 40520 -6640 40590
rect -6860 40480 -6640 40520
rect -6860 40410 -6850 40480
rect -6650 40410 -6640 40480
rect -6860 40360 -6640 40410
rect -6360 40590 -6140 40640
rect -6360 40520 -6350 40590
rect -6150 40520 -6140 40590
rect -6360 40480 -6140 40520
rect -6360 40410 -6350 40480
rect -6150 40410 -6140 40480
rect -6360 40360 -6140 40410
rect -5860 40590 -5640 40640
rect -5860 40520 -5850 40590
rect -5650 40520 -5640 40590
rect -5860 40480 -5640 40520
rect -5860 40410 -5850 40480
rect -5650 40410 -5640 40480
rect -5860 40360 -5640 40410
rect -5360 40590 -5140 40640
rect -5360 40520 -5350 40590
rect -5150 40520 -5140 40590
rect -5360 40480 -5140 40520
rect -5360 40410 -5350 40480
rect -5150 40410 -5140 40480
rect -5360 40360 -5140 40410
rect -4860 40590 -4640 40640
rect -4860 40520 -4850 40590
rect -4650 40520 -4640 40590
rect -4860 40480 -4640 40520
rect -4860 40410 -4850 40480
rect -4650 40410 -4640 40480
rect -4860 40360 -4640 40410
rect -4360 40590 -4140 40640
rect -4360 40520 -4350 40590
rect -4150 40520 -4140 40590
rect -4360 40480 -4140 40520
rect -4360 40410 -4350 40480
rect -4150 40410 -4140 40480
rect -4360 40360 -4140 40410
rect -3860 40590 -3640 40640
rect -3860 40520 -3850 40590
rect -3650 40520 -3640 40590
rect -3860 40480 -3640 40520
rect -3860 40410 -3850 40480
rect -3650 40410 -3640 40480
rect -3860 40360 -3640 40410
rect -3360 40590 -3140 40640
rect -3360 40520 -3350 40590
rect -3150 40520 -3140 40590
rect -3360 40480 -3140 40520
rect -3360 40410 -3350 40480
rect -3150 40410 -3140 40480
rect -3360 40360 -3140 40410
rect -2860 40590 -2640 40640
rect -2860 40520 -2850 40590
rect -2650 40520 -2640 40590
rect -2860 40480 -2640 40520
rect -2860 40410 -2850 40480
rect -2650 40410 -2640 40480
rect -2860 40360 -2640 40410
rect -2360 40590 -2140 40640
rect -2360 40520 -2350 40590
rect -2150 40520 -2140 40590
rect -2360 40480 -2140 40520
rect -2360 40410 -2350 40480
rect -2150 40410 -2140 40480
rect -2360 40360 -2140 40410
rect -1860 40590 -1640 40640
rect -1860 40520 -1850 40590
rect -1650 40520 -1640 40590
rect -1860 40480 -1640 40520
rect -1860 40410 -1850 40480
rect -1650 40410 -1640 40480
rect -1860 40360 -1640 40410
rect -1360 40590 -1140 40640
rect -1360 40520 -1350 40590
rect -1150 40520 -1140 40590
rect -1360 40480 -1140 40520
rect -1360 40410 -1350 40480
rect -1150 40410 -1140 40480
rect -1360 40360 -1140 40410
rect -860 40590 -640 40640
rect -860 40520 -850 40590
rect -650 40520 -640 40590
rect -860 40480 -640 40520
rect -860 40410 -850 40480
rect -650 40410 -640 40480
rect -860 40360 -640 40410
rect -360 40590 -140 40640
rect -360 40520 -350 40590
rect -150 40520 -140 40590
rect -360 40480 -140 40520
rect -360 40410 -350 40480
rect -150 40410 -140 40480
rect -360 40360 -140 40410
rect 140 40590 360 40640
rect 140 40520 150 40590
rect 350 40520 360 40590
rect 140 40480 360 40520
rect 140 40410 150 40480
rect 350 40410 360 40480
rect 140 40360 360 40410
rect 640 40590 860 40640
rect 640 40520 650 40590
rect 850 40520 860 40590
rect 640 40480 860 40520
rect 640 40410 650 40480
rect 850 40410 860 40480
rect 640 40360 860 40410
rect 1140 40590 1360 40640
rect 1140 40520 1150 40590
rect 1350 40520 1360 40590
rect 1140 40480 1360 40520
rect 1140 40410 1150 40480
rect 1350 40410 1360 40480
rect 1140 40360 1360 40410
rect 1640 40590 1860 40640
rect 1640 40520 1650 40590
rect 1850 40520 1860 40590
rect 1640 40480 1860 40520
rect 1640 40410 1650 40480
rect 1850 40410 1860 40480
rect 1640 40360 1860 40410
rect 2140 40590 2360 40640
rect 2140 40520 2150 40590
rect 2350 40520 2360 40590
rect 2140 40480 2360 40520
rect 2140 40410 2150 40480
rect 2350 40410 2360 40480
rect 2140 40360 2360 40410
rect 2640 40590 2860 40640
rect 2640 40520 2650 40590
rect 2850 40520 2860 40590
rect 2640 40480 2860 40520
rect 2640 40410 2650 40480
rect 2850 40410 2860 40480
rect 2640 40360 2860 40410
rect 3140 40590 3360 40640
rect 3140 40520 3150 40590
rect 3350 40520 3360 40590
rect 3140 40480 3360 40520
rect 3140 40410 3150 40480
rect 3350 40410 3360 40480
rect 3140 40360 3360 40410
rect 3640 40590 3860 40640
rect 3640 40520 3650 40590
rect 3850 40520 3860 40590
rect 3640 40480 3860 40520
rect 3640 40410 3650 40480
rect 3850 40410 3860 40480
rect 3640 40360 3860 40410
rect -16000 40350 4000 40360
rect -16000 40150 -15980 40350
rect -15910 40150 -15590 40350
rect -15520 40150 -15480 40350
rect -15410 40150 -15090 40350
rect -15020 40150 -14980 40350
rect -14910 40150 -14590 40350
rect -14520 40150 -14480 40350
rect -14410 40150 -14090 40350
rect -14020 40150 -13980 40350
rect -13910 40150 -13590 40350
rect -13520 40150 -13480 40350
rect -13410 40150 -13090 40350
rect -13020 40150 -12980 40350
rect -12910 40150 -12590 40350
rect -12520 40150 -12480 40350
rect -12410 40150 -12090 40350
rect -12020 40150 -11980 40350
rect -11910 40150 -11590 40350
rect -11520 40150 -11480 40350
rect -11410 40150 -11090 40350
rect -11020 40150 -10980 40350
rect -10910 40150 -10590 40350
rect -10520 40150 -10480 40350
rect -10410 40150 -10090 40350
rect -10020 40150 -9980 40350
rect -9910 40150 -9590 40350
rect -9520 40150 -9480 40350
rect -9410 40150 -9090 40350
rect -9020 40150 -8980 40350
rect -8910 40150 -8590 40350
rect -8520 40150 -8480 40350
rect -8410 40150 -8090 40350
rect -8020 40150 -7980 40350
rect -7910 40150 -7590 40350
rect -7520 40150 -7480 40350
rect -7410 40150 -7090 40350
rect -7020 40150 -6980 40350
rect -6910 40150 -6590 40350
rect -6520 40150 -6480 40350
rect -6410 40150 -6090 40350
rect -6020 40150 -5980 40350
rect -5910 40150 -5590 40350
rect -5520 40150 -5480 40350
rect -5410 40150 -5090 40350
rect -5020 40150 -4980 40350
rect -4910 40150 -4590 40350
rect -4520 40150 -4480 40350
rect -4410 40150 -4090 40350
rect -4020 40150 -3980 40350
rect -3910 40150 -3590 40350
rect -3520 40150 -3480 40350
rect -3410 40150 -3090 40350
rect -3020 40150 -2980 40350
rect -2910 40150 -2590 40350
rect -2520 40150 -2480 40350
rect -2410 40150 -2090 40350
rect -2020 40150 -1980 40350
rect -1910 40150 -1590 40350
rect -1520 40150 -1480 40350
rect -1410 40150 -1090 40350
rect -1020 40150 -980 40350
rect -910 40150 -590 40350
rect -520 40150 -480 40350
rect -410 40150 -90 40350
rect -20 40150 20 40350
rect 90 40150 410 40350
rect 480 40150 520 40350
rect 590 40150 910 40350
rect 980 40150 1020 40350
rect 1090 40150 1410 40350
rect 1480 40150 1520 40350
rect 1590 40150 1910 40350
rect 1980 40150 2020 40350
rect 2090 40150 2410 40350
rect 2480 40150 2520 40350
rect 2590 40150 2910 40350
rect 2980 40150 3020 40350
rect 3090 40150 3410 40350
rect 3480 40150 3520 40350
rect 3590 40150 3910 40350
rect 3980 40150 4000 40350
rect -16000 40140 4000 40150
rect -15860 40090 -15640 40140
rect -15860 40020 -15850 40090
rect -15650 40020 -15640 40090
rect -27860 39980 -27640 40000
rect -27860 39910 -27850 39980
rect -27650 39910 -27640 39980
rect -27860 39860 -27640 39910
rect -27360 39980 -27140 40000
rect -27360 39910 -27350 39980
rect -27150 39910 -27140 39980
rect -27360 39860 -27140 39910
rect -26860 39980 -26640 40000
rect -26860 39910 -26850 39980
rect -26650 39910 -26640 39980
rect -26860 39860 -26640 39910
rect -26360 39980 -26140 40000
rect -26360 39910 -26350 39980
rect -26150 39910 -26140 39980
rect -26360 39860 -26140 39910
rect -25860 39980 -25640 40000
rect -25860 39910 -25850 39980
rect -25650 39910 -25640 39980
rect -25860 39860 -25640 39910
rect -25360 39980 -25140 40000
rect -25360 39910 -25350 39980
rect -25150 39910 -25140 39980
rect -25360 39860 -25140 39910
rect -24860 39980 -24640 40000
rect -24860 39910 -24850 39980
rect -24650 39910 -24640 39980
rect -24860 39860 -24640 39910
rect -24360 39980 -24140 40000
rect -24360 39910 -24350 39980
rect -24150 39910 -24140 39980
rect -24360 39860 -24140 39910
rect -23860 39980 -23640 40000
rect -23860 39910 -23850 39980
rect -23650 39910 -23640 39980
rect -23860 39860 -23640 39910
rect -23360 39980 -23140 40000
rect -23360 39910 -23350 39980
rect -23150 39910 -23140 39980
rect -23360 39860 -23140 39910
rect -22860 39980 -22640 40000
rect -22860 39910 -22850 39980
rect -22650 39910 -22640 39980
rect -22860 39860 -22640 39910
rect -22360 39980 -22140 40000
rect -22360 39910 -22350 39980
rect -22150 39910 -22140 39980
rect -22360 39860 -22140 39910
rect -21860 39980 -21640 40000
rect -21860 39910 -21850 39980
rect -21650 39910 -21640 39980
rect -21860 39860 -21640 39910
rect -21360 39980 -21140 40000
rect -21360 39910 -21350 39980
rect -21150 39910 -21140 39980
rect -21360 39860 -21140 39910
rect -20860 39980 -20640 40000
rect -20860 39910 -20850 39980
rect -20650 39910 -20640 39980
rect -20860 39860 -20640 39910
rect -20360 39980 -20140 40000
rect -20360 39910 -20350 39980
rect -20150 39910 -20140 39980
rect -20360 39860 -20140 39910
rect -19860 39980 -19640 40000
rect -19860 39910 -19850 39980
rect -19650 39910 -19640 39980
rect -19860 39860 -19640 39910
rect -19360 39980 -19140 40000
rect -19360 39910 -19350 39980
rect -19150 39910 -19140 39980
rect -19360 39860 -19140 39910
rect -18860 39980 -18640 40000
rect -18860 39910 -18850 39980
rect -18650 39910 -18640 39980
rect -18860 39860 -18640 39910
rect -18360 39980 -18140 40000
rect -18360 39910 -18350 39980
rect -18150 39910 -18140 39980
rect -18360 39860 -18140 39910
rect -17860 39980 -17640 40000
rect -17860 39910 -17850 39980
rect -17650 39910 -17640 39980
rect -17860 39860 -17640 39910
rect -17360 39980 -17140 40000
rect -17360 39910 -17350 39980
rect -17150 39910 -17140 39980
rect -17360 39860 -17140 39910
rect -16860 39980 -16640 40000
rect -16860 39910 -16850 39980
rect -16650 39910 -16640 39980
rect -16860 39860 -16640 39910
rect -16360 39980 -16140 40000
rect -16360 39910 -16350 39980
rect -16150 39910 -16140 39980
rect -16360 39860 -16140 39910
rect -15860 39980 -15640 40020
rect -15860 39910 -15850 39980
rect -15650 39910 -15640 39980
rect -15860 39860 -15640 39910
rect -15360 40090 -15140 40140
rect -15360 40020 -15350 40090
rect -15150 40020 -15140 40090
rect -15360 39980 -15140 40020
rect -15360 39910 -15350 39980
rect -15150 39910 -15140 39980
rect -15360 39860 -15140 39910
rect -14860 40090 -14640 40140
rect -14860 40020 -14850 40090
rect -14650 40020 -14640 40090
rect -14860 39980 -14640 40020
rect -14860 39910 -14850 39980
rect -14650 39910 -14640 39980
rect -14860 39860 -14640 39910
rect -14360 40090 -14140 40140
rect -14360 40020 -14350 40090
rect -14150 40020 -14140 40090
rect -14360 39980 -14140 40020
rect -14360 39910 -14350 39980
rect -14150 39910 -14140 39980
rect -14360 39860 -14140 39910
rect -13860 40090 -13640 40140
rect -13860 40020 -13850 40090
rect -13650 40020 -13640 40090
rect -13860 39980 -13640 40020
rect -13860 39910 -13850 39980
rect -13650 39910 -13640 39980
rect -13860 39860 -13640 39910
rect -13360 40090 -13140 40140
rect -13360 40020 -13350 40090
rect -13150 40020 -13140 40090
rect -13360 39980 -13140 40020
rect -13360 39910 -13350 39980
rect -13150 39910 -13140 39980
rect -13360 39860 -13140 39910
rect -12860 40090 -12640 40140
rect -12860 40020 -12850 40090
rect -12650 40020 -12640 40090
rect -12860 39980 -12640 40020
rect -12860 39910 -12850 39980
rect -12650 39910 -12640 39980
rect -12860 39860 -12640 39910
rect -12360 40090 -12140 40140
rect -12360 40020 -12350 40090
rect -12150 40020 -12140 40090
rect -12360 39980 -12140 40020
rect -12360 39910 -12350 39980
rect -12150 39910 -12140 39980
rect -12360 39860 -12140 39910
rect -11860 40090 -11640 40140
rect -11860 40020 -11850 40090
rect -11650 40020 -11640 40090
rect -11860 39980 -11640 40020
rect -11860 39910 -11850 39980
rect -11650 39910 -11640 39980
rect -11860 39860 -11640 39910
rect -11360 40090 -11140 40140
rect -11360 40020 -11350 40090
rect -11150 40020 -11140 40090
rect -11360 39980 -11140 40020
rect -11360 39910 -11350 39980
rect -11150 39910 -11140 39980
rect -11360 39860 -11140 39910
rect -10860 40090 -10640 40140
rect -10860 40020 -10850 40090
rect -10650 40020 -10640 40090
rect -10860 39980 -10640 40020
rect -10860 39910 -10850 39980
rect -10650 39910 -10640 39980
rect -10860 39860 -10640 39910
rect -10360 40090 -10140 40140
rect -10360 40020 -10350 40090
rect -10150 40020 -10140 40090
rect -10360 39980 -10140 40020
rect -10360 39910 -10350 39980
rect -10150 39910 -10140 39980
rect -10360 39860 -10140 39910
rect -9860 40090 -9640 40140
rect -9860 40020 -9850 40090
rect -9650 40020 -9640 40090
rect -9860 39980 -9640 40020
rect -9860 39910 -9850 39980
rect -9650 39910 -9640 39980
rect -9860 39860 -9640 39910
rect -9360 40090 -9140 40140
rect -9360 40020 -9350 40090
rect -9150 40020 -9140 40090
rect -9360 39980 -9140 40020
rect -9360 39910 -9350 39980
rect -9150 39910 -9140 39980
rect -9360 39860 -9140 39910
rect -8860 40090 -8640 40140
rect -8860 40020 -8850 40090
rect -8650 40020 -8640 40090
rect -8860 39980 -8640 40020
rect -8860 39910 -8850 39980
rect -8650 39910 -8640 39980
rect -8860 39860 -8640 39910
rect -8360 40090 -8140 40140
rect -8360 40020 -8350 40090
rect -8150 40020 -8140 40090
rect -8360 39980 -8140 40020
rect -8360 39910 -8350 39980
rect -8150 39910 -8140 39980
rect -8360 39860 -8140 39910
rect -7860 40090 -7640 40140
rect -7860 40020 -7850 40090
rect -7650 40020 -7640 40090
rect -7860 39980 -7640 40020
rect -7860 39910 -7850 39980
rect -7650 39910 -7640 39980
rect -7860 39860 -7640 39910
rect -7360 40090 -7140 40140
rect -7360 40020 -7350 40090
rect -7150 40020 -7140 40090
rect -7360 39980 -7140 40020
rect -7360 39910 -7350 39980
rect -7150 39910 -7140 39980
rect -7360 39860 -7140 39910
rect -6860 40090 -6640 40140
rect -6860 40020 -6850 40090
rect -6650 40020 -6640 40090
rect -6860 39980 -6640 40020
rect -6860 39910 -6850 39980
rect -6650 39910 -6640 39980
rect -6860 39860 -6640 39910
rect -6360 40090 -6140 40140
rect -6360 40020 -6350 40090
rect -6150 40020 -6140 40090
rect -6360 39980 -6140 40020
rect -6360 39910 -6350 39980
rect -6150 39910 -6140 39980
rect -6360 39860 -6140 39910
rect -5860 40090 -5640 40140
rect -5860 40020 -5850 40090
rect -5650 40020 -5640 40090
rect -5860 39980 -5640 40020
rect -5860 39910 -5850 39980
rect -5650 39910 -5640 39980
rect -5860 39860 -5640 39910
rect -5360 40090 -5140 40140
rect -5360 40020 -5350 40090
rect -5150 40020 -5140 40090
rect -5360 39980 -5140 40020
rect -5360 39910 -5350 39980
rect -5150 39910 -5140 39980
rect -5360 39860 -5140 39910
rect -4860 40090 -4640 40140
rect -4860 40020 -4850 40090
rect -4650 40020 -4640 40090
rect -4860 39980 -4640 40020
rect -4860 39910 -4850 39980
rect -4650 39910 -4640 39980
rect -4860 39860 -4640 39910
rect -4360 40090 -4140 40140
rect -4360 40020 -4350 40090
rect -4150 40020 -4140 40090
rect -4360 39980 -4140 40020
rect -4360 39910 -4350 39980
rect -4150 39910 -4140 39980
rect -4360 39860 -4140 39910
rect -3860 40090 -3640 40140
rect -3860 40020 -3850 40090
rect -3650 40020 -3640 40090
rect -3860 39980 -3640 40020
rect -3860 39910 -3850 39980
rect -3650 39910 -3640 39980
rect -3860 39860 -3640 39910
rect -3360 40090 -3140 40140
rect -3360 40020 -3350 40090
rect -3150 40020 -3140 40090
rect -3360 39980 -3140 40020
rect -3360 39910 -3350 39980
rect -3150 39910 -3140 39980
rect -3360 39860 -3140 39910
rect -2860 40090 -2640 40140
rect -2860 40020 -2850 40090
rect -2650 40020 -2640 40090
rect -2860 39980 -2640 40020
rect -2860 39910 -2850 39980
rect -2650 39910 -2640 39980
rect -2860 39860 -2640 39910
rect -2360 40090 -2140 40140
rect -2360 40020 -2350 40090
rect -2150 40020 -2140 40090
rect -2360 39980 -2140 40020
rect -2360 39910 -2350 39980
rect -2150 39910 -2140 39980
rect -2360 39860 -2140 39910
rect -1860 40090 -1640 40140
rect -1860 40020 -1850 40090
rect -1650 40020 -1640 40090
rect -1860 39980 -1640 40020
rect -1860 39910 -1850 39980
rect -1650 39910 -1640 39980
rect -1860 39860 -1640 39910
rect -1360 40090 -1140 40140
rect -1360 40020 -1350 40090
rect -1150 40020 -1140 40090
rect -1360 39980 -1140 40020
rect -1360 39910 -1350 39980
rect -1150 39910 -1140 39980
rect -1360 39860 -1140 39910
rect -860 40090 -640 40140
rect -860 40020 -850 40090
rect -650 40020 -640 40090
rect -860 39980 -640 40020
rect -860 39910 -850 39980
rect -650 39910 -640 39980
rect -860 39860 -640 39910
rect -360 40090 -140 40140
rect -360 40020 -350 40090
rect -150 40020 -140 40090
rect -360 39980 -140 40020
rect -360 39910 -350 39980
rect -150 39910 -140 39980
rect -360 39860 -140 39910
rect 140 40090 360 40140
rect 140 40020 150 40090
rect 350 40020 360 40090
rect 140 39980 360 40020
rect 140 39910 150 39980
rect 350 39910 360 39980
rect 140 39860 360 39910
rect 640 40090 860 40140
rect 640 40020 650 40090
rect 850 40020 860 40090
rect 640 39980 860 40020
rect 640 39910 650 39980
rect 850 39910 860 39980
rect 640 39860 860 39910
rect 1140 40090 1360 40140
rect 1140 40020 1150 40090
rect 1350 40020 1360 40090
rect 1140 39980 1360 40020
rect 1140 39910 1150 39980
rect 1350 39910 1360 39980
rect 1140 39860 1360 39910
rect 1640 40090 1860 40140
rect 1640 40020 1650 40090
rect 1850 40020 1860 40090
rect 1640 39980 1860 40020
rect 1640 39910 1650 39980
rect 1850 39910 1860 39980
rect 1640 39860 1860 39910
rect 2140 40090 2360 40140
rect 2140 40020 2150 40090
rect 2350 40020 2360 40090
rect 2140 39980 2360 40020
rect 2140 39910 2150 39980
rect 2350 39910 2360 39980
rect 2140 39860 2360 39910
rect 2640 40090 2860 40140
rect 2640 40020 2650 40090
rect 2850 40020 2860 40090
rect 2640 39980 2860 40020
rect 2640 39910 2650 39980
rect 2850 39910 2860 39980
rect 2640 39860 2860 39910
rect 3140 40090 3360 40140
rect 3140 40020 3150 40090
rect 3350 40020 3360 40090
rect 3140 39980 3360 40020
rect 3140 39910 3150 39980
rect 3350 39910 3360 39980
rect 3140 39860 3360 39910
rect 3640 40090 3860 40140
rect 3640 40020 3650 40090
rect 3850 40020 3860 40090
rect 3640 39980 3860 40020
rect 3640 39910 3650 39980
rect 3850 39910 3860 39980
rect 3640 39860 3860 39910
rect -28000 39850 4000 39860
rect -28000 39650 -27980 39850
rect -27910 39650 -27590 39850
rect -27520 39650 -27480 39850
rect -27410 39650 -27090 39850
rect -27020 39650 -26980 39850
rect -26910 39650 -26590 39850
rect -26520 39650 -26480 39850
rect -26410 39650 -26090 39850
rect -26020 39650 -25980 39850
rect -25910 39650 -25590 39850
rect -25520 39650 -25480 39850
rect -25410 39650 -25090 39850
rect -25020 39650 -24980 39850
rect -24910 39650 -24590 39850
rect -24520 39650 -24480 39850
rect -24410 39650 -24090 39850
rect -24020 39650 -23980 39850
rect -23910 39650 -23590 39850
rect -23520 39650 -23480 39850
rect -23410 39650 -23090 39850
rect -23020 39650 -22980 39850
rect -22910 39650 -22590 39850
rect -22520 39650 -22480 39850
rect -22410 39650 -22090 39850
rect -22020 39650 -21980 39850
rect -21910 39650 -21590 39850
rect -21520 39650 -21480 39850
rect -21410 39650 -21090 39850
rect -21020 39650 -20980 39850
rect -20910 39650 -20590 39850
rect -20520 39650 -20480 39850
rect -20410 39650 -20090 39850
rect -20020 39650 -19980 39850
rect -19910 39650 -19590 39850
rect -19520 39650 -19480 39850
rect -19410 39650 -19090 39850
rect -19020 39650 -18980 39850
rect -18910 39650 -18590 39850
rect -18520 39650 -18480 39850
rect -18410 39650 -18090 39850
rect -18020 39650 -17980 39850
rect -17910 39650 -17590 39850
rect -17520 39650 -17480 39850
rect -17410 39650 -17090 39850
rect -17020 39650 -16980 39850
rect -16910 39650 -16590 39850
rect -16520 39650 -16480 39850
rect -16410 39650 -16090 39850
rect -16020 39650 -15980 39850
rect -15910 39650 -15590 39850
rect -15520 39650 -15480 39850
rect -15410 39650 -15090 39850
rect -15020 39650 -14980 39850
rect -14910 39650 -14590 39850
rect -14520 39650 -14480 39850
rect -14410 39650 -14090 39850
rect -14020 39650 -13980 39850
rect -13910 39650 -13590 39850
rect -13520 39650 -13480 39850
rect -13410 39650 -13090 39850
rect -13020 39650 -12980 39850
rect -12910 39650 -12590 39850
rect -12520 39650 -12480 39850
rect -12410 39650 -12090 39850
rect -12020 39650 -11980 39850
rect -11910 39650 -11590 39850
rect -11520 39650 -11480 39850
rect -11410 39650 -11090 39850
rect -11020 39650 -10980 39850
rect -10910 39650 -10590 39850
rect -10520 39650 -10480 39850
rect -10410 39650 -10090 39850
rect -10020 39650 -9980 39850
rect -9910 39650 -9590 39850
rect -9520 39650 -9480 39850
rect -9410 39650 -9090 39850
rect -9020 39650 -8980 39850
rect -8910 39650 -8590 39850
rect -8520 39650 -8480 39850
rect -8410 39650 -8090 39850
rect -8020 39650 -7980 39850
rect -7910 39650 -7590 39850
rect -7520 39650 -7480 39850
rect -7410 39650 -7090 39850
rect -7020 39650 -6980 39850
rect -6910 39650 -6590 39850
rect -6520 39650 -6480 39850
rect -6410 39650 -6090 39850
rect -6020 39650 -5980 39850
rect -5910 39650 -5590 39850
rect -5520 39650 -5480 39850
rect -5410 39650 -5090 39850
rect -5020 39650 -4980 39850
rect -4910 39650 -4590 39850
rect -4520 39650 -4480 39850
rect -4410 39650 -4090 39850
rect -4020 39650 -3980 39850
rect -3910 39650 -3590 39850
rect -3520 39650 -3480 39850
rect -3410 39650 -3090 39850
rect -3020 39650 -2980 39850
rect -2910 39650 -2590 39850
rect -2520 39650 -2480 39850
rect -2410 39650 -2090 39850
rect -2020 39650 -1980 39850
rect -1910 39650 -1590 39850
rect -1520 39650 -1480 39850
rect -1410 39650 -1090 39850
rect -1020 39650 -980 39850
rect -910 39650 -590 39850
rect -520 39650 -480 39850
rect -410 39650 -90 39850
rect -20 39650 20 39850
rect 90 39650 410 39850
rect 480 39650 520 39850
rect 590 39650 910 39850
rect 980 39650 1020 39850
rect 1090 39650 1410 39850
rect 1480 39650 1520 39850
rect 1590 39650 1910 39850
rect 1980 39650 2020 39850
rect 2090 39650 2410 39850
rect 2480 39650 2520 39850
rect 2590 39650 2910 39850
rect 2980 39650 3020 39850
rect 3090 39650 3410 39850
rect 3480 39650 3520 39850
rect 3590 39650 3910 39850
rect 3980 39650 4000 39850
rect -28000 39640 4000 39650
rect -27860 39590 -27640 39640
rect -27860 39520 -27850 39590
rect -27650 39520 -27640 39590
rect -27860 39480 -27640 39520
rect -27860 39410 -27850 39480
rect -27650 39410 -27640 39480
rect -27860 39360 -27640 39410
rect -27360 39590 -27140 39640
rect -27360 39520 -27350 39590
rect -27150 39520 -27140 39590
rect -27360 39480 -27140 39520
rect -27360 39410 -27350 39480
rect -27150 39410 -27140 39480
rect -27360 39360 -27140 39410
rect -26860 39590 -26640 39640
rect -26860 39520 -26850 39590
rect -26650 39520 -26640 39590
rect -26860 39480 -26640 39520
rect -26860 39410 -26850 39480
rect -26650 39410 -26640 39480
rect -26860 39360 -26640 39410
rect -26360 39590 -26140 39640
rect -26360 39520 -26350 39590
rect -26150 39520 -26140 39590
rect -26360 39480 -26140 39520
rect -26360 39410 -26350 39480
rect -26150 39410 -26140 39480
rect -26360 39360 -26140 39410
rect -25860 39590 -25640 39640
rect -25860 39520 -25850 39590
rect -25650 39520 -25640 39590
rect -25860 39480 -25640 39520
rect -25860 39410 -25850 39480
rect -25650 39410 -25640 39480
rect -25860 39360 -25640 39410
rect -25360 39590 -25140 39640
rect -25360 39520 -25350 39590
rect -25150 39520 -25140 39590
rect -25360 39480 -25140 39520
rect -25360 39410 -25350 39480
rect -25150 39410 -25140 39480
rect -25360 39360 -25140 39410
rect -24860 39590 -24640 39640
rect -24860 39520 -24850 39590
rect -24650 39520 -24640 39590
rect -24860 39480 -24640 39520
rect -24860 39410 -24850 39480
rect -24650 39410 -24640 39480
rect -24860 39360 -24640 39410
rect -24360 39590 -24140 39640
rect -24360 39520 -24350 39590
rect -24150 39520 -24140 39590
rect -24360 39480 -24140 39520
rect -24360 39410 -24350 39480
rect -24150 39410 -24140 39480
rect -24360 39360 -24140 39410
rect -23860 39590 -23640 39640
rect -23860 39520 -23850 39590
rect -23650 39520 -23640 39590
rect -23860 39480 -23640 39520
rect -23860 39410 -23850 39480
rect -23650 39410 -23640 39480
rect -23860 39360 -23640 39410
rect -23360 39590 -23140 39640
rect -23360 39520 -23350 39590
rect -23150 39520 -23140 39590
rect -23360 39480 -23140 39520
rect -23360 39410 -23350 39480
rect -23150 39410 -23140 39480
rect -23360 39360 -23140 39410
rect -22860 39590 -22640 39640
rect -22860 39520 -22850 39590
rect -22650 39520 -22640 39590
rect -22860 39480 -22640 39520
rect -22860 39410 -22850 39480
rect -22650 39410 -22640 39480
rect -22860 39360 -22640 39410
rect -22360 39590 -22140 39640
rect -22360 39520 -22350 39590
rect -22150 39520 -22140 39590
rect -22360 39480 -22140 39520
rect -22360 39410 -22350 39480
rect -22150 39410 -22140 39480
rect -22360 39360 -22140 39410
rect -21860 39590 -21640 39640
rect -21860 39520 -21850 39590
rect -21650 39520 -21640 39590
rect -21860 39480 -21640 39520
rect -21860 39410 -21850 39480
rect -21650 39410 -21640 39480
rect -21860 39360 -21640 39410
rect -21360 39590 -21140 39640
rect -21360 39520 -21350 39590
rect -21150 39520 -21140 39590
rect -21360 39480 -21140 39520
rect -21360 39410 -21350 39480
rect -21150 39410 -21140 39480
rect -21360 39360 -21140 39410
rect -20860 39590 -20640 39640
rect -20860 39520 -20850 39590
rect -20650 39520 -20640 39590
rect -20860 39480 -20640 39520
rect -20860 39410 -20850 39480
rect -20650 39410 -20640 39480
rect -20860 39360 -20640 39410
rect -20360 39590 -20140 39640
rect -20360 39520 -20350 39590
rect -20150 39520 -20140 39590
rect -20360 39480 -20140 39520
rect -20360 39410 -20350 39480
rect -20150 39410 -20140 39480
rect -20360 39360 -20140 39410
rect -19860 39590 -19640 39640
rect -19860 39520 -19850 39590
rect -19650 39520 -19640 39590
rect -19860 39480 -19640 39520
rect -19860 39410 -19850 39480
rect -19650 39410 -19640 39480
rect -19860 39360 -19640 39410
rect -19360 39590 -19140 39640
rect -19360 39520 -19350 39590
rect -19150 39520 -19140 39590
rect -19360 39480 -19140 39520
rect -19360 39410 -19350 39480
rect -19150 39410 -19140 39480
rect -19360 39360 -19140 39410
rect -18860 39590 -18640 39640
rect -18860 39520 -18850 39590
rect -18650 39520 -18640 39590
rect -18860 39480 -18640 39520
rect -18860 39410 -18850 39480
rect -18650 39410 -18640 39480
rect -18860 39360 -18640 39410
rect -18360 39590 -18140 39640
rect -18360 39520 -18350 39590
rect -18150 39520 -18140 39590
rect -18360 39480 -18140 39520
rect -18360 39410 -18350 39480
rect -18150 39410 -18140 39480
rect -18360 39360 -18140 39410
rect -17860 39590 -17640 39640
rect -17860 39520 -17850 39590
rect -17650 39520 -17640 39590
rect -17860 39480 -17640 39520
rect -17860 39410 -17850 39480
rect -17650 39410 -17640 39480
rect -17860 39360 -17640 39410
rect -17360 39590 -17140 39640
rect -17360 39520 -17350 39590
rect -17150 39520 -17140 39590
rect -17360 39480 -17140 39520
rect -17360 39410 -17350 39480
rect -17150 39410 -17140 39480
rect -17360 39360 -17140 39410
rect -16860 39590 -16640 39640
rect -16860 39520 -16850 39590
rect -16650 39520 -16640 39590
rect -16860 39480 -16640 39520
rect -16860 39410 -16850 39480
rect -16650 39410 -16640 39480
rect -16860 39360 -16640 39410
rect -16360 39590 -16140 39640
rect -16360 39520 -16350 39590
rect -16150 39520 -16140 39590
rect -16360 39480 -16140 39520
rect -16360 39410 -16350 39480
rect -16150 39410 -16140 39480
rect -16360 39360 -16140 39410
rect -15860 39590 -15640 39640
rect -15860 39520 -15850 39590
rect -15650 39520 -15640 39590
rect -15860 39480 -15640 39520
rect -15860 39410 -15850 39480
rect -15650 39410 -15640 39480
rect -15860 39360 -15640 39410
rect -15360 39590 -15140 39640
rect -15360 39520 -15350 39590
rect -15150 39520 -15140 39590
rect -15360 39480 -15140 39520
rect -15360 39410 -15350 39480
rect -15150 39410 -15140 39480
rect -15360 39360 -15140 39410
rect -14860 39590 -14640 39640
rect -14860 39520 -14850 39590
rect -14650 39520 -14640 39590
rect -14860 39480 -14640 39520
rect -14860 39410 -14850 39480
rect -14650 39410 -14640 39480
rect -14860 39360 -14640 39410
rect -14360 39590 -14140 39640
rect -14360 39520 -14350 39590
rect -14150 39520 -14140 39590
rect -14360 39480 -14140 39520
rect -14360 39410 -14350 39480
rect -14150 39410 -14140 39480
rect -14360 39360 -14140 39410
rect -13860 39590 -13640 39640
rect -13860 39520 -13850 39590
rect -13650 39520 -13640 39590
rect -13860 39480 -13640 39520
rect -13860 39410 -13850 39480
rect -13650 39410 -13640 39480
rect -13860 39360 -13640 39410
rect -13360 39590 -13140 39640
rect -13360 39520 -13350 39590
rect -13150 39520 -13140 39590
rect -13360 39480 -13140 39520
rect -13360 39410 -13350 39480
rect -13150 39410 -13140 39480
rect -13360 39360 -13140 39410
rect -12860 39590 -12640 39640
rect -12860 39520 -12850 39590
rect -12650 39520 -12640 39590
rect -12860 39480 -12640 39520
rect -12860 39410 -12850 39480
rect -12650 39410 -12640 39480
rect -12860 39360 -12640 39410
rect -12360 39590 -12140 39640
rect -12360 39520 -12350 39590
rect -12150 39520 -12140 39590
rect -12360 39480 -12140 39520
rect -12360 39410 -12350 39480
rect -12150 39410 -12140 39480
rect -12360 39360 -12140 39410
rect -11860 39590 -11640 39640
rect -11860 39520 -11850 39590
rect -11650 39520 -11640 39590
rect -11860 39480 -11640 39520
rect -11860 39410 -11850 39480
rect -11650 39410 -11640 39480
rect -11860 39360 -11640 39410
rect -11360 39590 -11140 39640
rect -11360 39520 -11350 39590
rect -11150 39520 -11140 39590
rect -11360 39480 -11140 39520
rect -11360 39410 -11350 39480
rect -11150 39410 -11140 39480
rect -11360 39360 -11140 39410
rect -10860 39590 -10640 39640
rect -10860 39520 -10850 39590
rect -10650 39520 -10640 39590
rect -10860 39480 -10640 39520
rect -10860 39410 -10850 39480
rect -10650 39410 -10640 39480
rect -10860 39360 -10640 39410
rect -10360 39590 -10140 39640
rect -10360 39520 -10350 39590
rect -10150 39520 -10140 39590
rect -10360 39480 -10140 39520
rect -10360 39410 -10350 39480
rect -10150 39410 -10140 39480
rect -10360 39360 -10140 39410
rect -9860 39590 -9640 39640
rect -9860 39520 -9850 39590
rect -9650 39520 -9640 39590
rect -9860 39480 -9640 39520
rect -9860 39410 -9850 39480
rect -9650 39410 -9640 39480
rect -9860 39360 -9640 39410
rect -9360 39590 -9140 39640
rect -9360 39520 -9350 39590
rect -9150 39520 -9140 39590
rect -9360 39480 -9140 39520
rect -9360 39410 -9350 39480
rect -9150 39410 -9140 39480
rect -9360 39360 -9140 39410
rect -8860 39590 -8640 39640
rect -8860 39520 -8850 39590
rect -8650 39520 -8640 39590
rect -8860 39480 -8640 39520
rect -8860 39410 -8850 39480
rect -8650 39410 -8640 39480
rect -8860 39360 -8640 39410
rect -8360 39590 -8140 39640
rect -8360 39520 -8350 39590
rect -8150 39520 -8140 39590
rect -8360 39480 -8140 39520
rect -8360 39410 -8350 39480
rect -8150 39410 -8140 39480
rect -8360 39360 -8140 39410
rect -7860 39590 -7640 39640
rect -7860 39520 -7850 39590
rect -7650 39520 -7640 39590
rect -7860 39480 -7640 39520
rect -7860 39410 -7850 39480
rect -7650 39410 -7640 39480
rect -7860 39360 -7640 39410
rect -7360 39590 -7140 39640
rect -7360 39520 -7350 39590
rect -7150 39520 -7140 39590
rect -7360 39480 -7140 39520
rect -7360 39410 -7350 39480
rect -7150 39410 -7140 39480
rect -7360 39360 -7140 39410
rect -6860 39590 -6640 39640
rect -6860 39520 -6850 39590
rect -6650 39520 -6640 39590
rect -6860 39480 -6640 39520
rect -6860 39410 -6850 39480
rect -6650 39410 -6640 39480
rect -6860 39360 -6640 39410
rect -6360 39590 -6140 39640
rect -6360 39520 -6350 39590
rect -6150 39520 -6140 39590
rect -6360 39480 -6140 39520
rect -6360 39410 -6350 39480
rect -6150 39410 -6140 39480
rect -6360 39360 -6140 39410
rect -5860 39590 -5640 39640
rect -5860 39520 -5850 39590
rect -5650 39520 -5640 39590
rect -5860 39480 -5640 39520
rect -5860 39410 -5850 39480
rect -5650 39410 -5640 39480
rect -5860 39360 -5640 39410
rect -5360 39590 -5140 39640
rect -5360 39520 -5350 39590
rect -5150 39520 -5140 39590
rect -5360 39480 -5140 39520
rect -5360 39410 -5350 39480
rect -5150 39410 -5140 39480
rect -5360 39360 -5140 39410
rect -4860 39590 -4640 39640
rect -4860 39520 -4850 39590
rect -4650 39520 -4640 39590
rect -4860 39480 -4640 39520
rect -4860 39410 -4850 39480
rect -4650 39410 -4640 39480
rect -4860 39360 -4640 39410
rect -4360 39590 -4140 39640
rect -4360 39520 -4350 39590
rect -4150 39520 -4140 39590
rect -4360 39480 -4140 39520
rect -4360 39410 -4350 39480
rect -4150 39410 -4140 39480
rect -4360 39360 -4140 39410
rect -3860 39590 -3640 39640
rect -3860 39520 -3850 39590
rect -3650 39520 -3640 39590
rect -3860 39480 -3640 39520
rect -3860 39410 -3850 39480
rect -3650 39410 -3640 39480
rect -3860 39360 -3640 39410
rect -3360 39590 -3140 39640
rect -3360 39520 -3350 39590
rect -3150 39520 -3140 39590
rect -3360 39480 -3140 39520
rect -3360 39410 -3350 39480
rect -3150 39410 -3140 39480
rect -3360 39360 -3140 39410
rect -2860 39590 -2640 39640
rect -2860 39520 -2850 39590
rect -2650 39520 -2640 39590
rect -2860 39480 -2640 39520
rect -2860 39410 -2850 39480
rect -2650 39410 -2640 39480
rect -2860 39360 -2640 39410
rect -2360 39590 -2140 39640
rect -2360 39520 -2350 39590
rect -2150 39520 -2140 39590
rect -2360 39480 -2140 39520
rect -2360 39410 -2350 39480
rect -2150 39410 -2140 39480
rect -2360 39360 -2140 39410
rect -1860 39590 -1640 39640
rect -1860 39520 -1850 39590
rect -1650 39520 -1640 39590
rect -1860 39480 -1640 39520
rect -1860 39410 -1850 39480
rect -1650 39410 -1640 39480
rect -1860 39360 -1640 39410
rect -1360 39590 -1140 39640
rect -1360 39520 -1350 39590
rect -1150 39520 -1140 39590
rect -1360 39480 -1140 39520
rect -1360 39410 -1350 39480
rect -1150 39410 -1140 39480
rect -1360 39360 -1140 39410
rect -860 39590 -640 39640
rect -860 39520 -850 39590
rect -650 39520 -640 39590
rect -860 39480 -640 39520
rect -860 39410 -850 39480
rect -650 39410 -640 39480
rect -860 39360 -640 39410
rect -360 39590 -140 39640
rect -360 39520 -350 39590
rect -150 39520 -140 39590
rect -360 39480 -140 39520
rect -360 39410 -350 39480
rect -150 39410 -140 39480
rect -360 39360 -140 39410
rect 140 39590 360 39640
rect 140 39520 150 39590
rect 350 39520 360 39590
rect 140 39480 360 39520
rect 140 39410 150 39480
rect 350 39410 360 39480
rect 140 39360 360 39410
rect 640 39590 860 39640
rect 640 39520 650 39590
rect 850 39520 860 39590
rect 640 39480 860 39520
rect 640 39410 650 39480
rect 850 39410 860 39480
rect 640 39360 860 39410
rect 1140 39590 1360 39640
rect 1140 39520 1150 39590
rect 1350 39520 1360 39590
rect 1140 39480 1360 39520
rect 1140 39410 1150 39480
rect 1350 39410 1360 39480
rect 1140 39360 1360 39410
rect 1640 39590 1860 39640
rect 1640 39520 1650 39590
rect 1850 39520 1860 39590
rect 1640 39480 1860 39520
rect 1640 39410 1650 39480
rect 1850 39410 1860 39480
rect 1640 39360 1860 39410
rect 2140 39590 2360 39640
rect 2140 39520 2150 39590
rect 2350 39520 2360 39590
rect 2140 39480 2360 39520
rect 2140 39410 2150 39480
rect 2350 39410 2360 39480
rect 2140 39360 2360 39410
rect 2640 39590 2860 39640
rect 2640 39520 2650 39590
rect 2850 39520 2860 39590
rect 2640 39480 2860 39520
rect 2640 39410 2650 39480
rect 2850 39410 2860 39480
rect 2640 39360 2860 39410
rect 3140 39590 3360 39640
rect 3140 39520 3150 39590
rect 3350 39520 3360 39590
rect 3140 39480 3360 39520
rect 3140 39410 3150 39480
rect 3350 39410 3360 39480
rect 3140 39360 3360 39410
rect 3640 39590 3860 39640
rect 3640 39520 3650 39590
rect 3850 39520 3860 39590
rect 3640 39480 3860 39520
rect 3640 39410 3650 39480
rect 3850 39410 3860 39480
rect 3640 39360 3860 39410
rect -28000 39350 4000 39360
rect -28000 39150 -27980 39350
rect -27910 39150 -27590 39350
rect -27520 39150 -27480 39350
rect -27410 39150 -27090 39350
rect -27020 39150 -26980 39350
rect -26910 39150 -26590 39350
rect -26520 39150 -26480 39350
rect -26410 39150 -26090 39350
rect -26020 39150 -25980 39350
rect -25910 39150 -25590 39350
rect -25520 39150 -25480 39350
rect -25410 39150 -25090 39350
rect -25020 39150 -24980 39350
rect -24910 39150 -24590 39350
rect -24520 39150 -24480 39350
rect -24410 39150 -24090 39350
rect -24020 39150 -23980 39350
rect -23910 39150 -23590 39350
rect -23520 39150 -23480 39350
rect -23410 39150 -23090 39350
rect -23020 39150 -22980 39350
rect -22910 39150 -22590 39350
rect -22520 39150 -22480 39350
rect -22410 39150 -22090 39350
rect -22020 39150 -21980 39350
rect -21910 39150 -21590 39350
rect -21520 39150 -21480 39350
rect -21410 39150 -21090 39350
rect -21020 39150 -20980 39350
rect -20910 39150 -20590 39350
rect -20520 39150 -20480 39350
rect -20410 39150 -20090 39350
rect -20020 39150 -19980 39350
rect -19910 39150 -19590 39350
rect -19520 39150 -19480 39350
rect -19410 39150 -19090 39350
rect -19020 39150 -18980 39350
rect -18910 39150 -18590 39350
rect -18520 39150 -18480 39350
rect -18410 39150 -18090 39350
rect -18020 39150 -17980 39350
rect -17910 39150 -17590 39350
rect -17520 39150 -17480 39350
rect -17410 39150 -17090 39350
rect -17020 39150 -16980 39350
rect -16910 39150 -16590 39350
rect -16520 39150 -16480 39350
rect -16410 39150 -16090 39350
rect -16020 39150 -15980 39350
rect -15910 39150 -15590 39350
rect -15520 39150 -15480 39350
rect -15410 39150 -15090 39350
rect -15020 39150 -14980 39350
rect -14910 39150 -14590 39350
rect -14520 39150 -14480 39350
rect -14410 39150 -14090 39350
rect -14020 39150 -13980 39350
rect -13910 39150 -13590 39350
rect -13520 39150 -13480 39350
rect -13410 39150 -13090 39350
rect -13020 39150 -12980 39350
rect -12910 39150 -12590 39350
rect -12520 39150 -12480 39350
rect -12410 39150 -12090 39350
rect -12020 39150 -11980 39350
rect -11910 39150 -11590 39350
rect -11520 39150 -11480 39350
rect -11410 39150 -11090 39350
rect -11020 39150 -10980 39350
rect -10910 39150 -10590 39350
rect -10520 39150 -10480 39350
rect -10410 39150 -10090 39350
rect -10020 39150 -9980 39350
rect -9910 39150 -9590 39350
rect -9520 39150 -9480 39350
rect -9410 39150 -9090 39350
rect -9020 39150 -8980 39350
rect -8910 39150 -8590 39350
rect -8520 39150 -8480 39350
rect -8410 39150 -8090 39350
rect -8020 39150 -7980 39350
rect -7910 39150 -7590 39350
rect -7520 39150 -7480 39350
rect -7410 39150 -7090 39350
rect -7020 39150 -6980 39350
rect -6910 39150 -6590 39350
rect -6520 39150 -6480 39350
rect -6410 39150 -6090 39350
rect -6020 39150 -5980 39350
rect -5910 39150 -5590 39350
rect -5520 39150 -5480 39350
rect -5410 39150 -5090 39350
rect -5020 39150 -4980 39350
rect -4910 39150 -4590 39350
rect -4520 39150 -4480 39350
rect -4410 39150 -4090 39350
rect -4020 39150 -3980 39350
rect -3910 39150 -3590 39350
rect -3520 39150 -3480 39350
rect -3410 39150 -3090 39350
rect -3020 39150 -2980 39350
rect -2910 39150 -2590 39350
rect -2520 39150 -2480 39350
rect -2410 39150 -2090 39350
rect -2020 39150 -1980 39350
rect -1910 39150 -1590 39350
rect -1520 39150 -1480 39350
rect -1410 39150 -1090 39350
rect -1020 39150 -980 39350
rect -910 39150 -590 39350
rect -520 39150 -480 39350
rect -410 39150 -90 39350
rect -20 39150 20 39350
rect 90 39150 410 39350
rect 480 39150 520 39350
rect 590 39150 910 39350
rect 980 39150 1020 39350
rect 1090 39150 1410 39350
rect 1480 39150 1520 39350
rect 1590 39150 1910 39350
rect 1980 39150 2020 39350
rect 2090 39150 2410 39350
rect 2480 39150 2520 39350
rect 2590 39150 2910 39350
rect 2980 39150 3020 39350
rect 3090 39150 3410 39350
rect 3480 39150 3520 39350
rect 3590 39150 3910 39350
rect 3980 39150 4000 39350
rect -28000 39140 4000 39150
rect -27860 39090 -27640 39140
rect -27860 39020 -27850 39090
rect -27650 39020 -27640 39090
rect -27860 38980 -27640 39020
rect -27860 38910 -27850 38980
rect -27650 38910 -27640 38980
rect -27860 38860 -27640 38910
rect -27360 39090 -27140 39140
rect -27360 39020 -27350 39090
rect -27150 39020 -27140 39090
rect -27360 38980 -27140 39020
rect -27360 38910 -27350 38980
rect -27150 38910 -27140 38980
rect -27360 38860 -27140 38910
rect -26860 39090 -26640 39140
rect -26860 39020 -26850 39090
rect -26650 39020 -26640 39090
rect -26860 38980 -26640 39020
rect -26860 38910 -26850 38980
rect -26650 38910 -26640 38980
rect -26860 38860 -26640 38910
rect -26360 39090 -26140 39140
rect -26360 39020 -26350 39090
rect -26150 39020 -26140 39090
rect -26360 38980 -26140 39020
rect -26360 38910 -26350 38980
rect -26150 38910 -26140 38980
rect -26360 38860 -26140 38910
rect -25860 39090 -25640 39140
rect -25860 39020 -25850 39090
rect -25650 39020 -25640 39090
rect -25860 38980 -25640 39020
rect -25860 38910 -25850 38980
rect -25650 38910 -25640 38980
rect -25860 38860 -25640 38910
rect -25360 39090 -25140 39140
rect -25360 39020 -25350 39090
rect -25150 39020 -25140 39090
rect -25360 38980 -25140 39020
rect -25360 38910 -25350 38980
rect -25150 38910 -25140 38980
rect -25360 38860 -25140 38910
rect -24860 39090 -24640 39140
rect -24860 39020 -24850 39090
rect -24650 39020 -24640 39090
rect -24860 38980 -24640 39020
rect -24860 38910 -24850 38980
rect -24650 38910 -24640 38980
rect -24860 38860 -24640 38910
rect -24360 39090 -24140 39140
rect -24360 39020 -24350 39090
rect -24150 39020 -24140 39090
rect -24360 38980 -24140 39020
rect -24360 38910 -24350 38980
rect -24150 38910 -24140 38980
rect -24360 38860 -24140 38910
rect -23860 39090 -23640 39140
rect -23860 39020 -23850 39090
rect -23650 39020 -23640 39090
rect -23860 38980 -23640 39020
rect -23860 38910 -23850 38980
rect -23650 38910 -23640 38980
rect -23860 38860 -23640 38910
rect -23360 39090 -23140 39140
rect -23360 39020 -23350 39090
rect -23150 39020 -23140 39090
rect -23360 38980 -23140 39020
rect -23360 38910 -23350 38980
rect -23150 38910 -23140 38980
rect -23360 38860 -23140 38910
rect -22860 39090 -22640 39140
rect -22860 39020 -22850 39090
rect -22650 39020 -22640 39090
rect -22860 38980 -22640 39020
rect -22860 38910 -22850 38980
rect -22650 38910 -22640 38980
rect -22860 38860 -22640 38910
rect -22360 39090 -22140 39140
rect -22360 39020 -22350 39090
rect -22150 39020 -22140 39090
rect -22360 38980 -22140 39020
rect -22360 38910 -22350 38980
rect -22150 38910 -22140 38980
rect -22360 38860 -22140 38910
rect -21860 39090 -21640 39140
rect -21860 39020 -21850 39090
rect -21650 39020 -21640 39090
rect -21860 38980 -21640 39020
rect -21860 38910 -21850 38980
rect -21650 38910 -21640 38980
rect -21860 38860 -21640 38910
rect -21360 39090 -21140 39140
rect -21360 39020 -21350 39090
rect -21150 39020 -21140 39090
rect -21360 38980 -21140 39020
rect -21360 38910 -21350 38980
rect -21150 38910 -21140 38980
rect -21360 38860 -21140 38910
rect -20860 39090 -20640 39140
rect -20860 39020 -20850 39090
rect -20650 39020 -20640 39090
rect -20860 38980 -20640 39020
rect -20860 38910 -20850 38980
rect -20650 38910 -20640 38980
rect -20860 38860 -20640 38910
rect -20360 39090 -20140 39140
rect -20360 39020 -20350 39090
rect -20150 39020 -20140 39090
rect -20360 38980 -20140 39020
rect -20360 38910 -20350 38980
rect -20150 38910 -20140 38980
rect -20360 38860 -20140 38910
rect -19860 39090 -19640 39140
rect -19860 39020 -19850 39090
rect -19650 39020 -19640 39090
rect -19860 38980 -19640 39020
rect -19860 38910 -19850 38980
rect -19650 38910 -19640 38980
rect -19860 38860 -19640 38910
rect -19360 39090 -19140 39140
rect -19360 39020 -19350 39090
rect -19150 39020 -19140 39090
rect -19360 38980 -19140 39020
rect -19360 38910 -19350 38980
rect -19150 38910 -19140 38980
rect -19360 38860 -19140 38910
rect -18860 39090 -18640 39140
rect -18860 39020 -18850 39090
rect -18650 39020 -18640 39090
rect -18860 38980 -18640 39020
rect -18860 38910 -18850 38980
rect -18650 38910 -18640 38980
rect -18860 38860 -18640 38910
rect -18360 39090 -18140 39140
rect -18360 39020 -18350 39090
rect -18150 39020 -18140 39090
rect -18360 38980 -18140 39020
rect -18360 38910 -18350 38980
rect -18150 38910 -18140 38980
rect -18360 38860 -18140 38910
rect -17860 39090 -17640 39140
rect -17860 39020 -17850 39090
rect -17650 39020 -17640 39090
rect -17860 38980 -17640 39020
rect -17860 38910 -17850 38980
rect -17650 38910 -17640 38980
rect -17860 38860 -17640 38910
rect -17360 39090 -17140 39140
rect -17360 39020 -17350 39090
rect -17150 39020 -17140 39090
rect -17360 38980 -17140 39020
rect -17360 38910 -17350 38980
rect -17150 38910 -17140 38980
rect -17360 38860 -17140 38910
rect -16860 39090 -16640 39140
rect -16860 39020 -16850 39090
rect -16650 39020 -16640 39090
rect -16860 38980 -16640 39020
rect -16860 38910 -16850 38980
rect -16650 38910 -16640 38980
rect -16860 38860 -16640 38910
rect -16360 39090 -16140 39140
rect -16360 39020 -16350 39090
rect -16150 39020 -16140 39090
rect -16360 38980 -16140 39020
rect -16360 38910 -16350 38980
rect -16150 38910 -16140 38980
rect -16360 38860 -16140 38910
rect -15860 39090 -15640 39140
rect -15860 39020 -15850 39090
rect -15650 39020 -15640 39090
rect -15860 38980 -15640 39020
rect -15860 38910 -15850 38980
rect -15650 38910 -15640 38980
rect -15860 38860 -15640 38910
rect -15360 39090 -15140 39140
rect -15360 39020 -15350 39090
rect -15150 39020 -15140 39090
rect -15360 38980 -15140 39020
rect -15360 38910 -15350 38980
rect -15150 38910 -15140 38980
rect -15360 38860 -15140 38910
rect -14860 39090 -14640 39140
rect -14860 39020 -14850 39090
rect -14650 39020 -14640 39090
rect -14860 38980 -14640 39020
rect -14860 38910 -14850 38980
rect -14650 38910 -14640 38980
rect -14860 38860 -14640 38910
rect -14360 39090 -14140 39140
rect -14360 39020 -14350 39090
rect -14150 39020 -14140 39090
rect -14360 38980 -14140 39020
rect -14360 38910 -14350 38980
rect -14150 38910 -14140 38980
rect -14360 38860 -14140 38910
rect -13860 39090 -13640 39140
rect -13860 39020 -13850 39090
rect -13650 39020 -13640 39090
rect -13860 38980 -13640 39020
rect -13860 38910 -13850 38980
rect -13650 38910 -13640 38980
rect -13860 38860 -13640 38910
rect -13360 39090 -13140 39140
rect -13360 39020 -13350 39090
rect -13150 39020 -13140 39090
rect -13360 38980 -13140 39020
rect -13360 38910 -13350 38980
rect -13150 38910 -13140 38980
rect -13360 38860 -13140 38910
rect -12860 39090 -12640 39140
rect -12860 39020 -12850 39090
rect -12650 39020 -12640 39090
rect -12860 38980 -12640 39020
rect -12860 38910 -12850 38980
rect -12650 38910 -12640 38980
rect -12860 38860 -12640 38910
rect -12360 39090 -12140 39140
rect -12360 39020 -12350 39090
rect -12150 39020 -12140 39090
rect -12360 38980 -12140 39020
rect -12360 38910 -12350 38980
rect -12150 38910 -12140 38980
rect -12360 38860 -12140 38910
rect -11860 39090 -11640 39140
rect -11860 39020 -11850 39090
rect -11650 39020 -11640 39090
rect -11860 38980 -11640 39020
rect -11860 38910 -11850 38980
rect -11650 38910 -11640 38980
rect -11860 38860 -11640 38910
rect -11360 39090 -11140 39140
rect -11360 39020 -11350 39090
rect -11150 39020 -11140 39090
rect -11360 38980 -11140 39020
rect -11360 38910 -11350 38980
rect -11150 38910 -11140 38980
rect -11360 38860 -11140 38910
rect -10860 39090 -10640 39140
rect -10860 39020 -10850 39090
rect -10650 39020 -10640 39090
rect -10860 38980 -10640 39020
rect -10860 38910 -10850 38980
rect -10650 38910 -10640 38980
rect -10860 38860 -10640 38910
rect -10360 39090 -10140 39140
rect -10360 39020 -10350 39090
rect -10150 39020 -10140 39090
rect -10360 38980 -10140 39020
rect -10360 38910 -10350 38980
rect -10150 38910 -10140 38980
rect -10360 38860 -10140 38910
rect -9860 39090 -9640 39140
rect -9860 39020 -9850 39090
rect -9650 39020 -9640 39090
rect -9860 38980 -9640 39020
rect -9860 38910 -9850 38980
rect -9650 38910 -9640 38980
rect -9860 38860 -9640 38910
rect -9360 39090 -9140 39140
rect -9360 39020 -9350 39090
rect -9150 39020 -9140 39090
rect -9360 38980 -9140 39020
rect -9360 38910 -9350 38980
rect -9150 38910 -9140 38980
rect -9360 38860 -9140 38910
rect -8860 39090 -8640 39140
rect -8860 39020 -8850 39090
rect -8650 39020 -8640 39090
rect -8860 38980 -8640 39020
rect -8860 38910 -8850 38980
rect -8650 38910 -8640 38980
rect -8860 38860 -8640 38910
rect -8360 39090 -8140 39140
rect -8360 39020 -8350 39090
rect -8150 39020 -8140 39090
rect -8360 38980 -8140 39020
rect -8360 38910 -8350 38980
rect -8150 38910 -8140 38980
rect -8360 38860 -8140 38910
rect -7860 39090 -7640 39140
rect -7860 39020 -7850 39090
rect -7650 39020 -7640 39090
rect -7860 38980 -7640 39020
rect -7860 38910 -7850 38980
rect -7650 38910 -7640 38980
rect -7860 38860 -7640 38910
rect -7360 39090 -7140 39140
rect -7360 39020 -7350 39090
rect -7150 39020 -7140 39090
rect -7360 38980 -7140 39020
rect -7360 38910 -7350 38980
rect -7150 38910 -7140 38980
rect -7360 38860 -7140 38910
rect -6860 39090 -6640 39140
rect -6860 39020 -6850 39090
rect -6650 39020 -6640 39090
rect -6860 38980 -6640 39020
rect -6860 38910 -6850 38980
rect -6650 38910 -6640 38980
rect -6860 38860 -6640 38910
rect -6360 39090 -6140 39140
rect -6360 39020 -6350 39090
rect -6150 39020 -6140 39090
rect -6360 38980 -6140 39020
rect -6360 38910 -6350 38980
rect -6150 38910 -6140 38980
rect -6360 38860 -6140 38910
rect -5860 39090 -5640 39140
rect -5860 39020 -5850 39090
rect -5650 39020 -5640 39090
rect -5860 38980 -5640 39020
rect -5860 38910 -5850 38980
rect -5650 38910 -5640 38980
rect -5860 38860 -5640 38910
rect -5360 39090 -5140 39140
rect -5360 39020 -5350 39090
rect -5150 39020 -5140 39090
rect -5360 38980 -5140 39020
rect -5360 38910 -5350 38980
rect -5150 38910 -5140 38980
rect -5360 38860 -5140 38910
rect -4860 39090 -4640 39140
rect -4860 39020 -4850 39090
rect -4650 39020 -4640 39090
rect -4860 38980 -4640 39020
rect -4860 38910 -4850 38980
rect -4650 38910 -4640 38980
rect -4860 38860 -4640 38910
rect -4360 39090 -4140 39140
rect -4360 39020 -4350 39090
rect -4150 39020 -4140 39090
rect -4360 38980 -4140 39020
rect -4360 38910 -4350 38980
rect -4150 38910 -4140 38980
rect -4360 38860 -4140 38910
rect -3860 39090 -3640 39140
rect -3860 39020 -3850 39090
rect -3650 39020 -3640 39090
rect -3860 38980 -3640 39020
rect -3860 38910 -3850 38980
rect -3650 38910 -3640 38980
rect -3860 38860 -3640 38910
rect -3360 39090 -3140 39140
rect -3360 39020 -3350 39090
rect -3150 39020 -3140 39090
rect -3360 38980 -3140 39020
rect -3360 38910 -3350 38980
rect -3150 38910 -3140 38980
rect -3360 38860 -3140 38910
rect -2860 39090 -2640 39140
rect -2860 39020 -2850 39090
rect -2650 39020 -2640 39090
rect -2860 38980 -2640 39020
rect -2860 38910 -2850 38980
rect -2650 38910 -2640 38980
rect -2860 38860 -2640 38910
rect -2360 39090 -2140 39140
rect -2360 39020 -2350 39090
rect -2150 39020 -2140 39090
rect -2360 38980 -2140 39020
rect -2360 38910 -2350 38980
rect -2150 38910 -2140 38980
rect -2360 38860 -2140 38910
rect -1860 39090 -1640 39140
rect -1860 39020 -1850 39090
rect -1650 39020 -1640 39090
rect -1860 38980 -1640 39020
rect -1860 38910 -1850 38980
rect -1650 38910 -1640 38980
rect -1860 38860 -1640 38910
rect -1360 39090 -1140 39140
rect -1360 39020 -1350 39090
rect -1150 39020 -1140 39090
rect -1360 38980 -1140 39020
rect -1360 38910 -1350 38980
rect -1150 38910 -1140 38980
rect -1360 38860 -1140 38910
rect -860 39090 -640 39140
rect -860 39020 -850 39090
rect -650 39020 -640 39090
rect -860 38980 -640 39020
rect -860 38910 -850 38980
rect -650 38910 -640 38980
rect -860 38860 -640 38910
rect -360 39090 -140 39140
rect -360 39020 -350 39090
rect -150 39020 -140 39090
rect -360 38980 -140 39020
rect -360 38910 -350 38980
rect -150 38910 -140 38980
rect -360 38860 -140 38910
rect 140 39090 360 39140
rect 140 39020 150 39090
rect 350 39020 360 39090
rect 140 38980 360 39020
rect 140 38910 150 38980
rect 350 38910 360 38980
rect 140 38860 360 38910
rect 640 39090 860 39140
rect 640 39020 650 39090
rect 850 39020 860 39090
rect 640 38980 860 39020
rect 640 38910 650 38980
rect 850 38910 860 38980
rect 640 38860 860 38910
rect 1140 39090 1360 39140
rect 1140 39020 1150 39090
rect 1350 39020 1360 39090
rect 1140 38980 1360 39020
rect 1140 38910 1150 38980
rect 1350 38910 1360 38980
rect 1140 38860 1360 38910
rect 1640 39090 1860 39140
rect 1640 39020 1650 39090
rect 1850 39020 1860 39090
rect 1640 38980 1860 39020
rect 1640 38910 1650 38980
rect 1850 38910 1860 38980
rect 1640 38860 1860 38910
rect 2140 39090 2360 39140
rect 2140 39020 2150 39090
rect 2350 39020 2360 39090
rect 2140 38980 2360 39020
rect 2140 38910 2150 38980
rect 2350 38910 2360 38980
rect 2140 38860 2360 38910
rect 2640 39090 2860 39140
rect 2640 39020 2650 39090
rect 2850 39020 2860 39090
rect 2640 38980 2860 39020
rect 2640 38910 2650 38980
rect 2850 38910 2860 38980
rect 2640 38860 2860 38910
rect 3140 39090 3360 39140
rect 3140 39020 3150 39090
rect 3350 39020 3360 39090
rect 3140 38980 3360 39020
rect 3140 38910 3150 38980
rect 3350 38910 3360 38980
rect 3140 38860 3360 38910
rect 3640 39090 3860 39140
rect 3640 39020 3650 39090
rect 3850 39020 3860 39090
rect 3640 38980 3860 39020
rect 3640 38910 3650 38980
rect 3850 38910 3860 38980
rect 3640 38860 3860 38910
rect -28000 38850 4000 38860
rect -28000 38650 -27980 38850
rect -27910 38650 -27590 38850
rect -27520 38650 -27480 38850
rect -27410 38650 -27090 38850
rect -27020 38650 -26980 38850
rect -26910 38650 -26590 38850
rect -26520 38650 -26480 38850
rect -26410 38650 -26090 38850
rect -26020 38650 -25980 38850
rect -25910 38650 -25590 38850
rect -25520 38650 -25480 38850
rect -25410 38650 -25090 38850
rect -25020 38650 -24980 38850
rect -24910 38650 -24590 38850
rect -24520 38650 -24480 38850
rect -24410 38650 -24090 38850
rect -24020 38650 -23980 38850
rect -23910 38650 -23590 38850
rect -23520 38650 -23480 38850
rect -23410 38650 -23090 38850
rect -23020 38650 -22980 38850
rect -22910 38650 -22590 38850
rect -22520 38650 -22480 38850
rect -22410 38650 -22090 38850
rect -22020 38650 -21980 38850
rect -21910 38650 -21590 38850
rect -21520 38650 -21480 38850
rect -21410 38650 -21090 38850
rect -21020 38650 -20980 38850
rect -20910 38650 -20590 38850
rect -20520 38650 -20480 38850
rect -20410 38650 -20090 38850
rect -20020 38650 -19980 38850
rect -19910 38650 -19590 38850
rect -19520 38650 -19480 38850
rect -19410 38650 -19090 38850
rect -19020 38650 -18980 38850
rect -18910 38650 -18590 38850
rect -18520 38650 -18480 38850
rect -18410 38650 -18090 38850
rect -18020 38650 -17980 38850
rect -17910 38650 -17590 38850
rect -17520 38650 -17480 38850
rect -17410 38650 -17090 38850
rect -17020 38650 -16980 38850
rect -16910 38650 -16590 38850
rect -16520 38650 -16480 38850
rect -16410 38650 -16090 38850
rect -16020 38650 -15980 38850
rect -15910 38650 -15590 38850
rect -15520 38650 -15480 38850
rect -15410 38650 -15090 38850
rect -15020 38650 -14980 38850
rect -14910 38650 -14590 38850
rect -14520 38650 -14480 38850
rect -14410 38650 -14090 38850
rect -14020 38650 -13980 38850
rect -13910 38650 -13590 38850
rect -13520 38650 -13480 38850
rect -13410 38650 -13090 38850
rect -13020 38650 -12980 38850
rect -12910 38650 -12590 38850
rect -12520 38650 -12480 38850
rect -12410 38650 -12090 38850
rect -12020 38650 -11980 38850
rect -11910 38650 -11590 38850
rect -11520 38650 -11480 38850
rect -11410 38650 -11090 38850
rect -11020 38650 -10980 38850
rect -10910 38650 -10590 38850
rect -10520 38650 -10480 38850
rect -10410 38650 -10090 38850
rect -10020 38650 -9980 38850
rect -9910 38650 -9590 38850
rect -9520 38650 -9480 38850
rect -9410 38650 -9090 38850
rect -9020 38650 -8980 38850
rect -8910 38650 -8590 38850
rect -8520 38650 -8480 38850
rect -8410 38650 -8090 38850
rect -8020 38650 -7980 38850
rect -7910 38650 -7590 38850
rect -7520 38650 -7480 38850
rect -7410 38650 -7090 38850
rect -7020 38650 -6980 38850
rect -6910 38650 -6590 38850
rect -6520 38650 -6480 38850
rect -6410 38650 -6090 38850
rect -6020 38650 -5980 38850
rect -5910 38650 -5590 38850
rect -5520 38650 -5480 38850
rect -5410 38650 -5090 38850
rect -5020 38650 -4980 38850
rect -4910 38650 -4590 38850
rect -4520 38650 -4480 38850
rect -4410 38650 -4090 38850
rect -4020 38650 -3980 38850
rect -3910 38650 -3590 38850
rect -3520 38650 -3480 38850
rect -3410 38650 -3090 38850
rect -3020 38650 -2980 38850
rect -2910 38650 -2590 38850
rect -2520 38650 -2480 38850
rect -2410 38650 -2090 38850
rect -2020 38650 -1980 38850
rect -1910 38650 -1590 38850
rect -1520 38650 -1480 38850
rect -1410 38650 -1090 38850
rect -1020 38650 -980 38850
rect -910 38650 -590 38850
rect -520 38650 -480 38850
rect -410 38650 -90 38850
rect -20 38650 20 38850
rect 90 38650 410 38850
rect 480 38650 520 38850
rect 590 38650 910 38850
rect 980 38650 1020 38850
rect 1090 38650 1410 38850
rect 1480 38650 1520 38850
rect 1590 38650 1910 38850
rect 1980 38650 2020 38850
rect 2090 38650 2410 38850
rect 2480 38650 2520 38850
rect 2590 38650 2910 38850
rect 2980 38650 3020 38850
rect 3090 38650 3410 38850
rect 3480 38650 3520 38850
rect 3590 38650 3910 38850
rect 3980 38650 4000 38850
rect -28000 38640 4000 38650
rect -27860 38590 -27640 38640
rect -27860 38520 -27850 38590
rect -27650 38520 -27640 38590
rect -27860 38480 -27640 38520
rect -27860 38410 -27850 38480
rect -27650 38410 -27640 38480
rect -27860 38360 -27640 38410
rect -27360 38590 -27140 38640
rect -27360 38520 -27350 38590
rect -27150 38520 -27140 38590
rect -27360 38480 -27140 38520
rect -27360 38410 -27350 38480
rect -27150 38410 -27140 38480
rect -27360 38360 -27140 38410
rect -26860 38590 -26640 38640
rect -26860 38520 -26850 38590
rect -26650 38520 -26640 38590
rect -26860 38480 -26640 38520
rect -26860 38410 -26850 38480
rect -26650 38410 -26640 38480
rect -26860 38360 -26640 38410
rect -26360 38590 -26140 38640
rect -26360 38520 -26350 38590
rect -26150 38520 -26140 38590
rect -26360 38480 -26140 38520
rect -26360 38410 -26350 38480
rect -26150 38410 -26140 38480
rect -26360 38360 -26140 38410
rect -25860 38590 -25640 38640
rect -25860 38520 -25850 38590
rect -25650 38520 -25640 38590
rect -25860 38480 -25640 38520
rect -25860 38410 -25850 38480
rect -25650 38410 -25640 38480
rect -25860 38360 -25640 38410
rect -25360 38590 -25140 38640
rect -25360 38520 -25350 38590
rect -25150 38520 -25140 38590
rect -25360 38480 -25140 38520
rect -25360 38410 -25350 38480
rect -25150 38410 -25140 38480
rect -25360 38360 -25140 38410
rect -24860 38590 -24640 38640
rect -24860 38520 -24850 38590
rect -24650 38520 -24640 38590
rect -24860 38480 -24640 38520
rect -24860 38410 -24850 38480
rect -24650 38410 -24640 38480
rect -24860 38360 -24640 38410
rect -24360 38590 -24140 38640
rect -24360 38520 -24350 38590
rect -24150 38520 -24140 38590
rect -24360 38480 -24140 38520
rect -24360 38410 -24350 38480
rect -24150 38410 -24140 38480
rect -24360 38360 -24140 38410
rect -23860 38590 -23640 38640
rect -23860 38520 -23850 38590
rect -23650 38520 -23640 38590
rect -23860 38480 -23640 38520
rect -23860 38410 -23850 38480
rect -23650 38410 -23640 38480
rect -23860 38360 -23640 38410
rect -23360 38590 -23140 38640
rect -23360 38520 -23350 38590
rect -23150 38520 -23140 38590
rect -23360 38480 -23140 38520
rect -23360 38410 -23350 38480
rect -23150 38410 -23140 38480
rect -23360 38360 -23140 38410
rect -22860 38590 -22640 38640
rect -22860 38520 -22850 38590
rect -22650 38520 -22640 38590
rect -22860 38480 -22640 38520
rect -22860 38410 -22850 38480
rect -22650 38410 -22640 38480
rect -22860 38360 -22640 38410
rect -22360 38590 -22140 38640
rect -22360 38520 -22350 38590
rect -22150 38520 -22140 38590
rect -22360 38480 -22140 38520
rect -22360 38410 -22350 38480
rect -22150 38410 -22140 38480
rect -22360 38360 -22140 38410
rect -21860 38590 -21640 38640
rect -21860 38520 -21850 38590
rect -21650 38520 -21640 38590
rect -21860 38480 -21640 38520
rect -21860 38410 -21850 38480
rect -21650 38410 -21640 38480
rect -21860 38360 -21640 38410
rect -21360 38590 -21140 38640
rect -21360 38520 -21350 38590
rect -21150 38520 -21140 38590
rect -21360 38480 -21140 38520
rect -21360 38410 -21350 38480
rect -21150 38410 -21140 38480
rect -21360 38360 -21140 38410
rect -20860 38590 -20640 38640
rect -20860 38520 -20850 38590
rect -20650 38520 -20640 38590
rect -20860 38480 -20640 38520
rect -20860 38410 -20850 38480
rect -20650 38410 -20640 38480
rect -20860 38360 -20640 38410
rect -20360 38590 -20140 38640
rect -20360 38520 -20350 38590
rect -20150 38520 -20140 38590
rect -20360 38480 -20140 38520
rect -20360 38410 -20350 38480
rect -20150 38410 -20140 38480
rect -20360 38360 -20140 38410
rect -19860 38590 -19640 38640
rect -19860 38520 -19850 38590
rect -19650 38520 -19640 38590
rect -19860 38480 -19640 38520
rect -19860 38410 -19850 38480
rect -19650 38410 -19640 38480
rect -19860 38360 -19640 38410
rect -19360 38590 -19140 38640
rect -19360 38520 -19350 38590
rect -19150 38520 -19140 38590
rect -19360 38480 -19140 38520
rect -19360 38410 -19350 38480
rect -19150 38410 -19140 38480
rect -19360 38360 -19140 38410
rect -18860 38590 -18640 38640
rect -18860 38520 -18850 38590
rect -18650 38520 -18640 38590
rect -18860 38480 -18640 38520
rect -18860 38410 -18850 38480
rect -18650 38410 -18640 38480
rect -18860 38360 -18640 38410
rect -18360 38590 -18140 38640
rect -18360 38520 -18350 38590
rect -18150 38520 -18140 38590
rect -18360 38480 -18140 38520
rect -18360 38410 -18350 38480
rect -18150 38410 -18140 38480
rect -18360 38360 -18140 38410
rect -17860 38590 -17640 38640
rect -17860 38520 -17850 38590
rect -17650 38520 -17640 38590
rect -17860 38480 -17640 38520
rect -17860 38410 -17850 38480
rect -17650 38410 -17640 38480
rect -17860 38360 -17640 38410
rect -17360 38590 -17140 38640
rect -17360 38520 -17350 38590
rect -17150 38520 -17140 38590
rect -17360 38480 -17140 38520
rect -17360 38410 -17350 38480
rect -17150 38410 -17140 38480
rect -17360 38360 -17140 38410
rect -16860 38590 -16640 38640
rect -16860 38520 -16850 38590
rect -16650 38520 -16640 38590
rect -16860 38480 -16640 38520
rect -16860 38410 -16850 38480
rect -16650 38410 -16640 38480
rect -16860 38360 -16640 38410
rect -16360 38590 -16140 38640
rect -16360 38520 -16350 38590
rect -16150 38520 -16140 38590
rect -16360 38480 -16140 38520
rect -16360 38410 -16350 38480
rect -16150 38410 -16140 38480
rect -16360 38360 -16140 38410
rect -15860 38590 -15640 38640
rect -15860 38520 -15850 38590
rect -15650 38520 -15640 38590
rect -15860 38480 -15640 38520
rect -15860 38410 -15850 38480
rect -15650 38410 -15640 38480
rect -15860 38360 -15640 38410
rect -15360 38590 -15140 38640
rect -15360 38520 -15350 38590
rect -15150 38520 -15140 38590
rect -15360 38480 -15140 38520
rect -15360 38410 -15350 38480
rect -15150 38410 -15140 38480
rect -15360 38360 -15140 38410
rect -14860 38590 -14640 38640
rect -14860 38520 -14850 38590
rect -14650 38520 -14640 38590
rect -14860 38480 -14640 38520
rect -14860 38410 -14850 38480
rect -14650 38410 -14640 38480
rect -14860 38360 -14640 38410
rect -14360 38590 -14140 38640
rect -14360 38520 -14350 38590
rect -14150 38520 -14140 38590
rect -14360 38480 -14140 38520
rect -14360 38410 -14350 38480
rect -14150 38410 -14140 38480
rect -14360 38360 -14140 38410
rect -13860 38590 -13640 38640
rect -13860 38520 -13850 38590
rect -13650 38520 -13640 38590
rect -13860 38480 -13640 38520
rect -13860 38410 -13850 38480
rect -13650 38410 -13640 38480
rect -13860 38360 -13640 38410
rect -13360 38590 -13140 38640
rect -13360 38520 -13350 38590
rect -13150 38520 -13140 38590
rect -13360 38480 -13140 38520
rect -13360 38410 -13350 38480
rect -13150 38410 -13140 38480
rect -13360 38360 -13140 38410
rect -12860 38590 -12640 38640
rect -12860 38520 -12850 38590
rect -12650 38520 -12640 38590
rect -12860 38480 -12640 38520
rect -12860 38410 -12850 38480
rect -12650 38410 -12640 38480
rect -12860 38360 -12640 38410
rect -12360 38590 -12140 38640
rect -12360 38520 -12350 38590
rect -12150 38520 -12140 38590
rect -12360 38480 -12140 38520
rect -12360 38410 -12350 38480
rect -12150 38410 -12140 38480
rect -12360 38360 -12140 38410
rect -11860 38590 -11640 38640
rect -11860 38520 -11850 38590
rect -11650 38520 -11640 38590
rect -11860 38480 -11640 38520
rect -11860 38410 -11850 38480
rect -11650 38410 -11640 38480
rect -11860 38360 -11640 38410
rect -11360 38590 -11140 38640
rect -11360 38520 -11350 38590
rect -11150 38520 -11140 38590
rect -11360 38480 -11140 38520
rect -11360 38410 -11350 38480
rect -11150 38410 -11140 38480
rect -11360 38360 -11140 38410
rect -10860 38590 -10640 38640
rect -10860 38520 -10850 38590
rect -10650 38520 -10640 38590
rect -10860 38480 -10640 38520
rect -10860 38410 -10850 38480
rect -10650 38410 -10640 38480
rect -10860 38360 -10640 38410
rect -10360 38590 -10140 38640
rect -10360 38520 -10350 38590
rect -10150 38520 -10140 38590
rect -10360 38480 -10140 38520
rect -10360 38410 -10350 38480
rect -10150 38410 -10140 38480
rect -10360 38360 -10140 38410
rect -9860 38590 -9640 38640
rect -9860 38520 -9850 38590
rect -9650 38520 -9640 38590
rect -9860 38480 -9640 38520
rect -9860 38410 -9850 38480
rect -9650 38410 -9640 38480
rect -9860 38360 -9640 38410
rect -9360 38590 -9140 38640
rect -9360 38520 -9350 38590
rect -9150 38520 -9140 38590
rect -9360 38480 -9140 38520
rect -9360 38410 -9350 38480
rect -9150 38410 -9140 38480
rect -9360 38360 -9140 38410
rect -8860 38590 -8640 38640
rect -8860 38520 -8850 38590
rect -8650 38520 -8640 38590
rect -8860 38480 -8640 38520
rect -8860 38410 -8850 38480
rect -8650 38410 -8640 38480
rect -8860 38360 -8640 38410
rect -8360 38590 -8140 38640
rect -8360 38520 -8350 38590
rect -8150 38520 -8140 38590
rect -8360 38480 -8140 38520
rect -8360 38410 -8350 38480
rect -8150 38410 -8140 38480
rect -8360 38360 -8140 38410
rect -7860 38590 -7640 38640
rect -7860 38520 -7850 38590
rect -7650 38520 -7640 38590
rect -7860 38480 -7640 38520
rect -7860 38410 -7850 38480
rect -7650 38410 -7640 38480
rect -7860 38360 -7640 38410
rect -7360 38590 -7140 38640
rect -7360 38520 -7350 38590
rect -7150 38520 -7140 38590
rect -7360 38480 -7140 38520
rect -7360 38410 -7350 38480
rect -7150 38410 -7140 38480
rect -7360 38360 -7140 38410
rect -6860 38590 -6640 38640
rect -6860 38520 -6850 38590
rect -6650 38520 -6640 38590
rect -6860 38480 -6640 38520
rect -6860 38410 -6850 38480
rect -6650 38410 -6640 38480
rect -6860 38360 -6640 38410
rect -6360 38590 -6140 38640
rect -6360 38520 -6350 38590
rect -6150 38520 -6140 38590
rect -6360 38480 -6140 38520
rect -6360 38410 -6350 38480
rect -6150 38410 -6140 38480
rect -6360 38360 -6140 38410
rect -5860 38590 -5640 38640
rect -5860 38520 -5850 38590
rect -5650 38520 -5640 38590
rect -5860 38480 -5640 38520
rect -5860 38410 -5850 38480
rect -5650 38410 -5640 38480
rect -5860 38360 -5640 38410
rect -5360 38590 -5140 38640
rect -5360 38520 -5350 38590
rect -5150 38520 -5140 38590
rect -5360 38480 -5140 38520
rect -5360 38410 -5350 38480
rect -5150 38410 -5140 38480
rect -5360 38360 -5140 38410
rect -4860 38590 -4640 38640
rect -4860 38520 -4850 38590
rect -4650 38520 -4640 38590
rect -4860 38480 -4640 38520
rect -4860 38410 -4850 38480
rect -4650 38410 -4640 38480
rect -4860 38360 -4640 38410
rect -4360 38590 -4140 38640
rect -4360 38520 -4350 38590
rect -4150 38520 -4140 38590
rect -4360 38480 -4140 38520
rect -4360 38410 -4350 38480
rect -4150 38410 -4140 38480
rect -4360 38360 -4140 38410
rect -3860 38590 -3640 38640
rect -3860 38520 -3850 38590
rect -3650 38520 -3640 38590
rect -3860 38480 -3640 38520
rect -3860 38410 -3850 38480
rect -3650 38410 -3640 38480
rect -3860 38360 -3640 38410
rect -3360 38590 -3140 38640
rect -3360 38520 -3350 38590
rect -3150 38520 -3140 38590
rect -3360 38480 -3140 38520
rect -3360 38410 -3350 38480
rect -3150 38410 -3140 38480
rect -3360 38360 -3140 38410
rect -2860 38590 -2640 38640
rect -2860 38520 -2850 38590
rect -2650 38520 -2640 38590
rect -2860 38480 -2640 38520
rect -2860 38410 -2850 38480
rect -2650 38410 -2640 38480
rect -2860 38360 -2640 38410
rect -2360 38590 -2140 38640
rect -2360 38520 -2350 38590
rect -2150 38520 -2140 38590
rect -2360 38480 -2140 38520
rect -2360 38410 -2350 38480
rect -2150 38410 -2140 38480
rect -2360 38360 -2140 38410
rect -1860 38590 -1640 38640
rect -1860 38520 -1850 38590
rect -1650 38520 -1640 38590
rect -1860 38480 -1640 38520
rect -1860 38410 -1850 38480
rect -1650 38410 -1640 38480
rect -1860 38360 -1640 38410
rect -1360 38590 -1140 38640
rect -1360 38520 -1350 38590
rect -1150 38520 -1140 38590
rect -1360 38480 -1140 38520
rect -1360 38410 -1350 38480
rect -1150 38410 -1140 38480
rect -1360 38360 -1140 38410
rect -860 38590 -640 38640
rect -860 38520 -850 38590
rect -650 38520 -640 38590
rect -860 38480 -640 38520
rect -860 38410 -850 38480
rect -650 38410 -640 38480
rect -860 38360 -640 38410
rect -360 38590 -140 38640
rect -360 38520 -350 38590
rect -150 38520 -140 38590
rect -360 38480 -140 38520
rect -360 38410 -350 38480
rect -150 38410 -140 38480
rect -360 38360 -140 38410
rect 140 38590 360 38640
rect 140 38520 150 38590
rect 350 38520 360 38590
rect 140 38480 360 38520
rect 140 38410 150 38480
rect 350 38410 360 38480
rect 140 38360 360 38410
rect 640 38590 860 38640
rect 640 38520 650 38590
rect 850 38520 860 38590
rect 640 38480 860 38520
rect 640 38410 650 38480
rect 850 38410 860 38480
rect 640 38360 860 38410
rect 1140 38590 1360 38640
rect 1140 38520 1150 38590
rect 1350 38520 1360 38590
rect 1140 38480 1360 38520
rect 1140 38410 1150 38480
rect 1350 38410 1360 38480
rect 1140 38360 1360 38410
rect 1640 38590 1860 38640
rect 1640 38520 1650 38590
rect 1850 38520 1860 38590
rect 1640 38480 1860 38520
rect 1640 38410 1650 38480
rect 1850 38410 1860 38480
rect 1640 38360 1860 38410
rect 2140 38590 2360 38640
rect 2140 38520 2150 38590
rect 2350 38520 2360 38590
rect 2140 38480 2360 38520
rect 2140 38410 2150 38480
rect 2350 38410 2360 38480
rect 2140 38360 2360 38410
rect 2640 38590 2860 38640
rect 2640 38520 2650 38590
rect 2850 38520 2860 38590
rect 2640 38480 2860 38520
rect 2640 38410 2650 38480
rect 2850 38410 2860 38480
rect 2640 38360 2860 38410
rect 3140 38590 3360 38640
rect 3140 38520 3150 38590
rect 3350 38520 3360 38590
rect 3140 38480 3360 38520
rect 3140 38410 3150 38480
rect 3350 38410 3360 38480
rect 3140 38360 3360 38410
rect 3640 38590 3860 38640
rect 3640 38520 3650 38590
rect 3850 38520 3860 38590
rect 3640 38480 3860 38520
rect 3640 38410 3650 38480
rect 3850 38410 3860 38480
rect 3640 38360 3860 38410
rect -28000 38350 4000 38360
rect -28000 38150 -27980 38350
rect -27910 38150 -27590 38350
rect -27520 38150 -27480 38350
rect -27410 38150 -27090 38350
rect -27020 38150 -26980 38350
rect -26910 38150 -26590 38350
rect -26520 38150 -26480 38350
rect -26410 38150 -26090 38350
rect -26020 38150 -25980 38350
rect -25910 38150 -25590 38350
rect -25520 38150 -25480 38350
rect -25410 38150 -25090 38350
rect -25020 38150 -24980 38350
rect -24910 38150 -24590 38350
rect -24520 38150 -24480 38350
rect -24410 38150 -24090 38350
rect -24020 38150 -23980 38350
rect -23910 38150 -23590 38350
rect -23520 38150 -23480 38350
rect -23410 38150 -23090 38350
rect -23020 38150 -22980 38350
rect -22910 38150 -22590 38350
rect -22520 38150 -22480 38350
rect -22410 38150 -22090 38350
rect -22020 38150 -21980 38350
rect -21910 38150 -21590 38350
rect -21520 38150 -21480 38350
rect -21410 38150 -21090 38350
rect -21020 38150 -20980 38350
rect -20910 38150 -20590 38350
rect -20520 38150 -20480 38350
rect -20410 38150 -20090 38350
rect -20020 38150 -19980 38350
rect -19910 38150 -19590 38350
rect -19520 38150 -19480 38350
rect -19410 38150 -19090 38350
rect -19020 38150 -18980 38350
rect -18910 38150 -18590 38350
rect -18520 38150 -18480 38350
rect -18410 38150 -18090 38350
rect -18020 38150 -17980 38350
rect -17910 38150 -17590 38350
rect -17520 38150 -17480 38350
rect -17410 38150 -17090 38350
rect -17020 38150 -16980 38350
rect -16910 38150 -16590 38350
rect -16520 38150 -16480 38350
rect -16410 38150 -16090 38350
rect -16020 38150 -15980 38350
rect -15910 38150 -15590 38350
rect -15520 38150 -15480 38350
rect -15410 38150 -15090 38350
rect -15020 38150 -14980 38350
rect -14910 38150 -14590 38350
rect -14520 38150 -14480 38350
rect -14410 38150 -14090 38350
rect -14020 38150 -13980 38350
rect -13910 38150 -13590 38350
rect -13520 38150 -13480 38350
rect -13410 38150 -13090 38350
rect -13020 38150 -12980 38350
rect -12910 38150 -12590 38350
rect -12520 38150 -12480 38350
rect -12410 38150 -12090 38350
rect -12020 38150 -11980 38350
rect -11910 38150 -11590 38350
rect -11520 38150 -11480 38350
rect -11410 38150 -11090 38350
rect -11020 38150 -10980 38350
rect -10910 38150 -10590 38350
rect -10520 38150 -10480 38350
rect -10410 38150 -10090 38350
rect -10020 38150 -9980 38350
rect -9910 38150 -9590 38350
rect -9520 38150 -9480 38350
rect -9410 38150 -9090 38350
rect -9020 38150 -8980 38350
rect -8910 38150 -8590 38350
rect -8520 38150 -8480 38350
rect -8410 38150 -8090 38350
rect -8020 38150 -7980 38350
rect -7910 38150 -7590 38350
rect -7520 38150 -7480 38350
rect -7410 38150 -7090 38350
rect -7020 38150 -6980 38350
rect -6910 38150 -6590 38350
rect -6520 38150 -6480 38350
rect -6410 38150 -6090 38350
rect -6020 38150 -5980 38350
rect -5910 38150 -5590 38350
rect -5520 38150 -5480 38350
rect -5410 38150 -5090 38350
rect -5020 38150 -4980 38350
rect -4910 38150 -4590 38350
rect -4520 38150 -4480 38350
rect -4410 38150 -4090 38350
rect -4020 38150 -3980 38350
rect -3910 38150 -3590 38350
rect -3520 38150 -3480 38350
rect -3410 38150 -3090 38350
rect -3020 38150 -2980 38350
rect -2910 38150 -2590 38350
rect -2520 38150 -2480 38350
rect -2410 38150 -2090 38350
rect -2020 38150 -1980 38350
rect -1910 38150 -1590 38350
rect -1520 38150 -1480 38350
rect -1410 38150 -1090 38350
rect -1020 38150 -980 38350
rect -910 38150 -590 38350
rect -520 38150 -480 38350
rect -410 38150 -90 38350
rect -20 38150 20 38350
rect 90 38150 410 38350
rect 480 38150 520 38350
rect 590 38150 910 38350
rect 980 38150 1020 38350
rect 1090 38150 1410 38350
rect 1480 38150 1520 38350
rect 1590 38150 1910 38350
rect 1980 38150 2020 38350
rect 2090 38150 2410 38350
rect 2480 38150 2520 38350
rect 2590 38150 2910 38350
rect 2980 38150 3020 38350
rect 3090 38150 3410 38350
rect 3480 38150 3520 38350
rect 3590 38150 3910 38350
rect 3980 38150 4000 38350
rect -28000 38140 4000 38150
rect -27860 38090 -27640 38140
rect -27860 38020 -27850 38090
rect -27650 38020 -27640 38090
rect -27860 38000 -27640 38020
rect -27360 38090 -27140 38140
rect -27360 38020 -27350 38090
rect -27150 38020 -27140 38090
rect -27360 38000 -27140 38020
rect -26860 38090 -26640 38140
rect -26860 38020 -26850 38090
rect -26650 38020 -26640 38090
rect -26860 38000 -26640 38020
rect -26360 38090 -26140 38140
rect -26360 38020 -26350 38090
rect -26150 38020 -26140 38090
rect -26360 38000 -26140 38020
rect -25860 38090 -25640 38140
rect -25860 38020 -25850 38090
rect -25650 38020 -25640 38090
rect -25860 38000 -25640 38020
rect -25360 38090 -25140 38140
rect -25360 38020 -25350 38090
rect -25150 38020 -25140 38090
rect -25360 38000 -25140 38020
rect -24860 38090 -24640 38140
rect -24860 38020 -24850 38090
rect -24650 38020 -24640 38090
rect -24860 38000 -24640 38020
rect -24360 38090 -24140 38140
rect -24360 38020 -24350 38090
rect -24150 38020 -24140 38090
rect -24360 38000 -24140 38020
rect -23860 38090 -23640 38140
rect -23860 38020 -23850 38090
rect -23650 38020 -23640 38090
rect -23860 38000 -23640 38020
rect -23360 38090 -23140 38140
rect -23360 38020 -23350 38090
rect -23150 38020 -23140 38090
rect -23360 38000 -23140 38020
rect -22860 38090 -22640 38140
rect -22860 38020 -22850 38090
rect -22650 38020 -22640 38090
rect -22860 38000 -22640 38020
rect -22360 38090 -22140 38140
rect -22360 38020 -22350 38090
rect -22150 38020 -22140 38090
rect -22360 38000 -22140 38020
rect -21860 38090 -21640 38140
rect -21860 38020 -21850 38090
rect -21650 38020 -21640 38090
rect -21860 38000 -21640 38020
rect -21360 38090 -21140 38140
rect -21360 38020 -21350 38090
rect -21150 38020 -21140 38090
rect -21360 38000 -21140 38020
rect -20860 38090 -20640 38140
rect -20860 38020 -20850 38090
rect -20650 38020 -20640 38090
rect -20860 38000 -20640 38020
rect -20360 38090 -20140 38140
rect -20360 38020 -20350 38090
rect -20150 38020 -20140 38090
rect -20360 38000 -20140 38020
rect -19860 38090 -19640 38140
rect -19860 38020 -19850 38090
rect -19650 38020 -19640 38090
rect -19860 38000 -19640 38020
rect -19360 38090 -19140 38140
rect -19360 38020 -19350 38090
rect -19150 38020 -19140 38090
rect -19360 38000 -19140 38020
rect -18860 38090 -18640 38140
rect -18860 38020 -18850 38090
rect -18650 38020 -18640 38090
rect -18860 38000 -18640 38020
rect -18360 38090 -18140 38140
rect -18360 38020 -18350 38090
rect -18150 38020 -18140 38090
rect -18360 38000 -18140 38020
rect -17860 38090 -17640 38140
rect -17860 38020 -17850 38090
rect -17650 38020 -17640 38090
rect -17860 38000 -17640 38020
rect -17360 38090 -17140 38140
rect -17360 38020 -17350 38090
rect -17150 38020 -17140 38090
rect -17360 38000 -17140 38020
rect -16860 38090 -16640 38140
rect -16860 38020 -16850 38090
rect -16650 38020 -16640 38090
rect -16860 38000 -16640 38020
rect -16360 38090 -16140 38140
rect -16360 38020 -16350 38090
rect -16150 38020 -16140 38090
rect -16360 38000 -16140 38020
rect -15860 38090 -15640 38140
rect -15860 38020 -15850 38090
rect -15650 38020 -15640 38090
rect -15860 38000 -15640 38020
rect -15360 38090 -15140 38140
rect -15360 38020 -15350 38090
rect -15150 38020 -15140 38090
rect -15360 38000 -15140 38020
rect -14860 38090 -14640 38140
rect -14860 38020 -14850 38090
rect -14650 38020 -14640 38090
rect -14860 38000 -14640 38020
rect -14360 38090 -14140 38140
rect -14360 38020 -14350 38090
rect -14150 38020 -14140 38090
rect -14360 38000 -14140 38020
rect -13860 38090 -13640 38140
rect -13860 38020 -13850 38090
rect -13650 38020 -13640 38090
rect -13860 38000 -13640 38020
rect -13360 38090 -13140 38140
rect -13360 38020 -13350 38090
rect -13150 38020 -13140 38090
rect -13360 38000 -13140 38020
rect -12860 38090 -12640 38140
rect -12860 38020 -12850 38090
rect -12650 38020 -12640 38090
rect -12860 38000 -12640 38020
rect -12360 38090 -12140 38140
rect -12360 38020 -12350 38090
rect -12150 38020 -12140 38090
rect -12360 38000 -12140 38020
rect -11860 38090 -11640 38140
rect -11860 38020 -11850 38090
rect -11650 38020 -11640 38090
rect -11860 38000 -11640 38020
rect -11360 38090 -11140 38140
rect -11360 38020 -11350 38090
rect -11150 38020 -11140 38090
rect -11360 38000 -11140 38020
rect -10860 38090 -10640 38140
rect -10860 38020 -10850 38090
rect -10650 38020 -10640 38090
rect -10860 38000 -10640 38020
rect -10360 38090 -10140 38140
rect -10360 38020 -10350 38090
rect -10150 38020 -10140 38090
rect -10360 38000 -10140 38020
rect -9860 38090 -9640 38140
rect -9860 38020 -9850 38090
rect -9650 38020 -9640 38090
rect -9860 38000 -9640 38020
rect -9360 38090 -9140 38140
rect -9360 38020 -9350 38090
rect -9150 38020 -9140 38090
rect -9360 38000 -9140 38020
rect -8860 38090 -8640 38140
rect -8860 38020 -8850 38090
rect -8650 38020 -8640 38090
rect -8860 38000 -8640 38020
rect -8360 38090 -8140 38140
rect -8360 38020 -8350 38090
rect -8150 38020 -8140 38090
rect -8360 38000 -8140 38020
rect -7860 38090 -7640 38140
rect -7860 38020 -7850 38090
rect -7650 38020 -7640 38090
rect -7860 38000 -7640 38020
rect -7360 38090 -7140 38140
rect -7360 38020 -7350 38090
rect -7150 38020 -7140 38090
rect -7360 38000 -7140 38020
rect -6860 38090 -6640 38140
rect -6860 38020 -6850 38090
rect -6650 38020 -6640 38090
rect -6860 38000 -6640 38020
rect -6360 38090 -6140 38140
rect -6360 38020 -6350 38090
rect -6150 38020 -6140 38090
rect -6360 38000 -6140 38020
rect -5860 38090 -5640 38140
rect -5860 38020 -5850 38090
rect -5650 38020 -5640 38090
rect -5860 38000 -5640 38020
rect -5360 38090 -5140 38140
rect -5360 38020 -5350 38090
rect -5150 38020 -5140 38090
rect -5360 38000 -5140 38020
rect -4860 38090 -4640 38140
rect -4860 38020 -4850 38090
rect -4650 38020 -4640 38090
rect -4860 38000 -4640 38020
rect -4360 38090 -4140 38140
rect -4360 38020 -4350 38090
rect -4150 38020 -4140 38090
rect -4360 38000 -4140 38020
rect -3860 38090 -3640 38140
rect -3860 38020 -3850 38090
rect -3650 38020 -3640 38090
rect -3860 38000 -3640 38020
rect -3360 38090 -3140 38140
rect -3360 38020 -3350 38090
rect -3150 38020 -3140 38090
rect -3360 38000 -3140 38020
rect -2860 38090 -2640 38140
rect -2860 38020 -2850 38090
rect -2650 38020 -2640 38090
rect -2860 38000 -2640 38020
rect -2360 38090 -2140 38140
rect -2360 38020 -2350 38090
rect -2150 38020 -2140 38090
rect -2360 38000 -2140 38020
rect -1860 38090 -1640 38140
rect -1860 38020 -1850 38090
rect -1650 38020 -1640 38090
rect -1860 38000 -1640 38020
rect -1360 38090 -1140 38140
rect -1360 38020 -1350 38090
rect -1150 38020 -1140 38090
rect -1360 38000 -1140 38020
rect -860 38090 -640 38140
rect -860 38020 -850 38090
rect -650 38020 -640 38090
rect -860 38000 -640 38020
rect -360 38090 -140 38140
rect -360 38020 -350 38090
rect -150 38020 -140 38090
rect -360 38000 -140 38020
rect 140 38090 360 38140
rect 140 38020 150 38090
rect 350 38020 360 38090
rect 140 38000 360 38020
rect 640 38090 860 38140
rect 640 38020 650 38090
rect 850 38020 860 38090
rect 640 38000 860 38020
rect 1140 38090 1360 38140
rect 1140 38020 1150 38090
rect 1350 38020 1360 38090
rect 1140 38000 1360 38020
rect 1640 38090 1860 38140
rect 1640 38020 1650 38090
rect 1850 38020 1860 38090
rect 1640 38000 1860 38020
rect 2140 38090 2360 38140
rect 2140 38020 2150 38090
rect 2350 38020 2360 38090
rect 2140 38000 2360 38020
rect 2640 38090 2860 38140
rect 2640 38020 2650 38090
rect 2850 38020 2860 38090
rect 2640 38000 2860 38020
rect 3140 38090 3360 38140
rect 3140 38020 3150 38090
rect 3350 38020 3360 38090
rect 3140 38000 3360 38020
rect 3640 38090 3860 38140
rect 3640 38020 3650 38090
rect 3850 38020 3860 38090
rect 3640 38000 3860 38020
rect 17800 36190 18400 36200
rect 17800 35810 17810 36190
rect 18390 35810 18400 36190
rect 17800 35800 18400 35810
rect 17800 35600 26800 35800
rect 17000 35590 17600 35600
rect 17000 35210 17010 35590
rect 17590 35400 17600 35590
rect 17590 35210 26400 35400
rect 17000 35200 26400 35210
rect 17000 34990 26000 35000
rect 17000 34610 17010 34990
rect 17590 34800 26000 34990
rect 17590 34610 17600 34800
rect 17000 34600 17600 34610
rect 17800 34400 25600 34600
rect 17800 34390 18400 34400
rect 17800 34010 17810 34390
rect 18390 34010 18400 34390
rect 17800 34000 18400 34010
rect 14600 33780 15200 33800
rect 14600 33220 14620 33780
rect 15180 33220 15200 33780
rect 14600 33200 15200 33220
rect 14800 31200 15200 33200
rect 25400 32200 25600 34400
rect 25800 32200 26000 34800
rect 26200 32200 26400 35200
rect 26600 32200 26800 35600
rect 15000 15800 15200 31200
rect 15000 15600 20700 15800
rect 20500 13400 20700 15600
rect 20500 13200 24500 13400
rect 24300 12900 24500 13200
rect 128140 10980 128360 11000
rect 128140 10910 128150 10980
rect 128350 10910 128360 10980
rect 128140 10860 128360 10910
rect 128640 10980 128860 11000
rect 128640 10910 128650 10980
rect 128850 10910 128860 10980
rect 128640 10860 128860 10910
rect 129140 10980 129360 11000
rect 129140 10910 129150 10980
rect 129350 10910 129360 10980
rect 129140 10860 129360 10910
rect 129640 10980 129860 11000
rect 129640 10910 129650 10980
rect 129850 10910 129860 10980
rect 129640 10860 129860 10910
rect 130140 10980 130360 11000
rect 130140 10910 130150 10980
rect 130350 10910 130360 10980
rect 130140 10860 130360 10910
rect 130640 10980 130860 11000
rect 130640 10910 130650 10980
rect 130850 10910 130860 10980
rect 130640 10860 130860 10910
rect 131140 10980 131360 11000
rect 131140 10910 131150 10980
rect 131350 10910 131360 10980
rect 131140 10860 131360 10910
rect 131640 10980 131860 11000
rect 131640 10910 131650 10980
rect 131850 10910 131860 10980
rect 131640 10860 131860 10910
rect 132140 10980 132360 11000
rect 132140 10910 132150 10980
rect 132350 10910 132360 10980
rect 132140 10860 132360 10910
rect 132640 10980 132860 11000
rect 132640 10910 132650 10980
rect 132850 10910 132860 10980
rect 132640 10860 132860 10910
rect 133140 10980 133360 11000
rect 133140 10910 133150 10980
rect 133350 10910 133360 10980
rect 133140 10860 133360 10910
rect 133640 10980 133860 11000
rect 133640 10910 133650 10980
rect 133850 10910 133860 10980
rect 133640 10860 133860 10910
rect 134140 10980 134360 11000
rect 134140 10910 134150 10980
rect 134350 10910 134360 10980
rect 134140 10860 134360 10910
rect 134640 10980 134860 11000
rect 134640 10910 134650 10980
rect 134850 10910 134860 10980
rect 134640 10860 134860 10910
rect 135140 10980 135360 11000
rect 135140 10910 135150 10980
rect 135350 10910 135360 10980
rect 135140 10860 135360 10910
rect 135640 10980 135860 11000
rect 135640 10910 135650 10980
rect 135850 10910 135860 10980
rect 135640 10860 135860 10910
rect 136140 10980 136360 11000
rect 136140 10910 136150 10980
rect 136350 10910 136360 10980
rect 136140 10860 136360 10910
rect 136640 10980 136860 11000
rect 136640 10910 136650 10980
rect 136850 10910 136860 10980
rect 136640 10860 136860 10910
rect 137140 10980 137360 11000
rect 137140 10910 137150 10980
rect 137350 10910 137360 10980
rect 137140 10860 137360 10910
rect 137640 10980 137860 11000
rect 137640 10910 137650 10980
rect 137850 10910 137860 10980
rect 137640 10860 137860 10910
rect 138140 10980 138360 11000
rect 138140 10910 138150 10980
rect 138350 10910 138360 10980
rect 138140 10860 138360 10910
rect 138640 10980 138860 11000
rect 138640 10910 138650 10980
rect 138850 10910 138860 10980
rect 138640 10860 138860 10910
rect 139140 10980 139360 11000
rect 139140 10910 139150 10980
rect 139350 10910 139360 10980
rect 139140 10860 139360 10910
rect 139640 10980 139860 11000
rect 139640 10910 139650 10980
rect 139850 10910 139860 10980
rect 139640 10860 139860 10910
rect 128000 10850 140000 10860
rect 128000 10650 128020 10850
rect 128090 10650 128410 10850
rect 128480 10650 128520 10850
rect 128590 10650 128910 10850
rect 128980 10650 129020 10850
rect 129090 10650 129410 10850
rect 129480 10650 129520 10850
rect 129590 10650 129910 10850
rect 129980 10650 130020 10850
rect 130090 10650 130410 10850
rect 130480 10650 130520 10850
rect 130590 10650 130910 10850
rect 130980 10650 131020 10850
rect 131090 10650 131410 10850
rect 131480 10650 131520 10850
rect 131590 10650 131910 10850
rect 131980 10650 132020 10850
rect 132090 10650 132410 10850
rect 132480 10650 132520 10850
rect 132590 10650 132910 10850
rect 132980 10650 133020 10850
rect 133090 10650 133410 10850
rect 133480 10650 133520 10850
rect 133590 10650 133910 10850
rect 133980 10650 134020 10850
rect 134090 10650 134410 10850
rect 134480 10650 134520 10850
rect 134590 10650 134910 10850
rect 134980 10650 135020 10850
rect 135090 10650 135410 10850
rect 135480 10650 135520 10850
rect 135590 10650 135910 10850
rect 135980 10650 136020 10850
rect 136090 10650 136410 10850
rect 136480 10650 136520 10850
rect 136590 10650 136910 10850
rect 136980 10650 137020 10850
rect 137090 10650 137410 10850
rect 137480 10650 137520 10850
rect 137590 10650 137910 10850
rect 137980 10650 138020 10850
rect 138090 10650 138410 10850
rect 138480 10650 138520 10850
rect 138590 10650 138910 10850
rect 138980 10650 139020 10850
rect 139090 10650 139410 10850
rect 139480 10650 139520 10850
rect 139590 10650 139910 10850
rect 139980 10650 140000 10850
rect 128000 10640 140000 10650
rect 128140 10590 128360 10640
rect 128140 10520 128150 10590
rect 128350 10520 128360 10590
rect 128140 10480 128360 10520
rect 128140 10410 128150 10480
rect 128350 10410 128360 10480
rect 128140 10360 128360 10410
rect 128640 10590 128860 10640
rect 128640 10520 128650 10590
rect 128850 10520 128860 10590
rect 128640 10480 128860 10520
rect 128640 10410 128650 10480
rect 128850 10410 128860 10480
rect 128640 10360 128860 10410
rect 129140 10590 129360 10640
rect 129140 10520 129150 10590
rect 129350 10520 129360 10590
rect 129140 10480 129360 10520
rect 129140 10410 129150 10480
rect 129350 10410 129360 10480
rect 129140 10360 129360 10410
rect 129640 10590 129860 10640
rect 129640 10520 129650 10590
rect 129850 10520 129860 10590
rect 129640 10480 129860 10520
rect 129640 10410 129650 10480
rect 129850 10410 129860 10480
rect 129640 10360 129860 10410
rect 130140 10590 130360 10640
rect 130140 10520 130150 10590
rect 130350 10520 130360 10590
rect 130140 10480 130360 10520
rect 130140 10410 130150 10480
rect 130350 10410 130360 10480
rect 130140 10360 130360 10410
rect 130640 10590 130860 10640
rect 130640 10520 130650 10590
rect 130850 10520 130860 10590
rect 130640 10480 130860 10520
rect 130640 10410 130650 10480
rect 130850 10410 130860 10480
rect 130640 10360 130860 10410
rect 131140 10590 131360 10640
rect 131140 10520 131150 10590
rect 131350 10520 131360 10590
rect 131140 10480 131360 10520
rect 131140 10410 131150 10480
rect 131350 10410 131360 10480
rect 131140 10360 131360 10410
rect 131640 10590 131860 10640
rect 131640 10520 131650 10590
rect 131850 10520 131860 10590
rect 131640 10480 131860 10520
rect 131640 10410 131650 10480
rect 131850 10410 131860 10480
rect 131640 10360 131860 10410
rect 132140 10590 132360 10640
rect 132140 10520 132150 10590
rect 132350 10520 132360 10590
rect 132140 10480 132360 10520
rect 132140 10410 132150 10480
rect 132350 10410 132360 10480
rect 132140 10360 132360 10410
rect 132640 10590 132860 10640
rect 132640 10520 132650 10590
rect 132850 10520 132860 10590
rect 132640 10480 132860 10520
rect 132640 10410 132650 10480
rect 132850 10410 132860 10480
rect 132640 10360 132860 10410
rect 133140 10590 133360 10640
rect 133140 10520 133150 10590
rect 133350 10520 133360 10590
rect 133140 10480 133360 10520
rect 133140 10410 133150 10480
rect 133350 10410 133360 10480
rect 133140 10360 133360 10410
rect 133640 10590 133860 10640
rect 133640 10520 133650 10590
rect 133850 10520 133860 10590
rect 133640 10480 133860 10520
rect 133640 10410 133650 10480
rect 133850 10410 133860 10480
rect 133640 10360 133860 10410
rect 134140 10590 134360 10640
rect 134140 10520 134150 10590
rect 134350 10520 134360 10590
rect 134140 10480 134360 10520
rect 134140 10410 134150 10480
rect 134350 10410 134360 10480
rect 134140 10360 134360 10410
rect 134640 10590 134860 10640
rect 134640 10520 134650 10590
rect 134850 10520 134860 10590
rect 134640 10480 134860 10520
rect 134640 10410 134650 10480
rect 134850 10410 134860 10480
rect 134640 10360 134860 10410
rect 135140 10590 135360 10640
rect 135140 10520 135150 10590
rect 135350 10520 135360 10590
rect 135140 10480 135360 10520
rect 135140 10410 135150 10480
rect 135350 10410 135360 10480
rect 135140 10360 135360 10410
rect 135640 10590 135860 10640
rect 135640 10520 135650 10590
rect 135850 10520 135860 10590
rect 135640 10480 135860 10520
rect 135640 10410 135650 10480
rect 135850 10410 135860 10480
rect 135640 10360 135860 10410
rect 136140 10590 136360 10640
rect 136140 10520 136150 10590
rect 136350 10520 136360 10590
rect 136140 10480 136360 10520
rect 136140 10410 136150 10480
rect 136350 10410 136360 10480
rect 136140 10360 136360 10410
rect 136640 10590 136860 10640
rect 136640 10520 136650 10590
rect 136850 10520 136860 10590
rect 136640 10480 136860 10520
rect 136640 10410 136650 10480
rect 136850 10410 136860 10480
rect 136640 10360 136860 10410
rect 137140 10590 137360 10640
rect 137140 10520 137150 10590
rect 137350 10520 137360 10590
rect 137140 10480 137360 10520
rect 137140 10410 137150 10480
rect 137350 10410 137360 10480
rect 137140 10360 137360 10410
rect 137640 10590 137860 10640
rect 137640 10520 137650 10590
rect 137850 10520 137860 10590
rect 137640 10480 137860 10520
rect 137640 10410 137650 10480
rect 137850 10410 137860 10480
rect 137640 10360 137860 10410
rect 138140 10590 138360 10640
rect 138140 10520 138150 10590
rect 138350 10520 138360 10590
rect 138140 10480 138360 10520
rect 138140 10410 138150 10480
rect 138350 10410 138360 10480
rect 138140 10360 138360 10410
rect 138640 10590 138860 10640
rect 138640 10520 138650 10590
rect 138850 10520 138860 10590
rect 138640 10480 138860 10520
rect 138640 10410 138650 10480
rect 138850 10410 138860 10480
rect 138640 10360 138860 10410
rect 139140 10590 139360 10640
rect 139140 10520 139150 10590
rect 139350 10520 139360 10590
rect 139140 10480 139360 10520
rect 139140 10410 139150 10480
rect 139350 10410 139360 10480
rect 139140 10360 139360 10410
rect 139640 10590 139860 10640
rect 139640 10520 139650 10590
rect 139850 10520 139860 10590
rect 139640 10480 139860 10520
rect 139640 10410 139650 10480
rect 139850 10410 139860 10480
rect 139640 10360 139860 10410
rect 128000 10350 140000 10360
rect 128000 10150 128020 10350
rect 128090 10150 128410 10350
rect 128480 10150 128520 10350
rect 128590 10150 128910 10350
rect 128980 10150 129020 10350
rect 129090 10150 129410 10350
rect 129480 10150 129520 10350
rect 129590 10150 129910 10350
rect 129980 10150 130020 10350
rect 130090 10150 130410 10350
rect 130480 10150 130520 10350
rect 130590 10150 130910 10350
rect 130980 10150 131020 10350
rect 131090 10150 131410 10350
rect 131480 10150 131520 10350
rect 131590 10150 131910 10350
rect 131980 10150 132020 10350
rect 132090 10150 132410 10350
rect 132480 10150 132520 10350
rect 132590 10150 132910 10350
rect 132980 10150 133020 10350
rect 133090 10150 133410 10350
rect 133480 10150 133520 10350
rect 133590 10150 133910 10350
rect 133980 10150 134020 10350
rect 134090 10150 134410 10350
rect 134480 10150 134520 10350
rect 134590 10150 134910 10350
rect 134980 10150 135020 10350
rect 135090 10150 135410 10350
rect 135480 10150 135520 10350
rect 135590 10150 135910 10350
rect 135980 10150 136020 10350
rect 136090 10150 136410 10350
rect 136480 10150 136520 10350
rect 136590 10150 136910 10350
rect 136980 10150 137020 10350
rect 137090 10150 137410 10350
rect 137480 10150 137520 10350
rect 137590 10150 137910 10350
rect 137980 10150 138020 10350
rect 138090 10150 138410 10350
rect 138480 10150 138520 10350
rect 138590 10150 138910 10350
rect 138980 10150 139020 10350
rect 139090 10150 139410 10350
rect 139480 10150 139520 10350
rect 139590 10150 139910 10350
rect 139980 10150 140000 10350
rect 128000 10140 140000 10150
rect 128140 10090 128360 10140
rect 128140 10020 128150 10090
rect 128350 10020 128360 10090
rect 128140 9980 128360 10020
rect 128140 9910 128150 9980
rect 128350 9910 128360 9980
rect 128140 9860 128360 9910
rect 128640 10090 128860 10140
rect 128640 10020 128650 10090
rect 128850 10020 128860 10090
rect 128640 9980 128860 10020
rect 128640 9910 128650 9980
rect 128850 9910 128860 9980
rect 128640 9860 128860 9910
rect 129140 10090 129360 10140
rect 129140 10020 129150 10090
rect 129350 10020 129360 10090
rect 129140 9980 129360 10020
rect 129140 9910 129150 9980
rect 129350 9910 129360 9980
rect 129140 9860 129360 9910
rect 129640 10090 129860 10140
rect 129640 10020 129650 10090
rect 129850 10020 129860 10090
rect 129640 9980 129860 10020
rect 129640 9910 129650 9980
rect 129850 9910 129860 9980
rect 129640 9860 129860 9910
rect 130140 10090 130360 10140
rect 130140 10020 130150 10090
rect 130350 10020 130360 10090
rect 130140 9980 130360 10020
rect 130140 9910 130150 9980
rect 130350 9910 130360 9980
rect 130140 9860 130360 9910
rect 130640 10090 130860 10140
rect 130640 10020 130650 10090
rect 130850 10020 130860 10090
rect 130640 9980 130860 10020
rect 130640 9910 130650 9980
rect 130850 9910 130860 9980
rect 130640 9860 130860 9910
rect 131140 10090 131360 10140
rect 131140 10020 131150 10090
rect 131350 10020 131360 10090
rect 131140 9980 131360 10020
rect 131140 9910 131150 9980
rect 131350 9910 131360 9980
rect 131140 9860 131360 9910
rect 131640 10090 131860 10140
rect 131640 10020 131650 10090
rect 131850 10020 131860 10090
rect 131640 9980 131860 10020
rect 131640 9910 131650 9980
rect 131850 9910 131860 9980
rect 131640 9860 131860 9910
rect 132140 10090 132360 10140
rect 132140 10020 132150 10090
rect 132350 10020 132360 10090
rect 132140 9980 132360 10020
rect 132140 9910 132150 9980
rect 132350 9910 132360 9980
rect 132140 9860 132360 9910
rect 132640 10090 132860 10140
rect 132640 10020 132650 10090
rect 132850 10020 132860 10090
rect 132640 9980 132860 10020
rect 132640 9910 132650 9980
rect 132850 9910 132860 9980
rect 132640 9860 132860 9910
rect 133140 10090 133360 10140
rect 133140 10020 133150 10090
rect 133350 10020 133360 10090
rect 133140 9980 133360 10020
rect 133140 9910 133150 9980
rect 133350 9910 133360 9980
rect 133140 9860 133360 9910
rect 133640 10090 133860 10140
rect 133640 10020 133650 10090
rect 133850 10020 133860 10090
rect 133640 9980 133860 10020
rect 133640 9910 133650 9980
rect 133850 9910 133860 9980
rect 133640 9860 133860 9910
rect 134140 10090 134360 10140
rect 134140 10020 134150 10090
rect 134350 10020 134360 10090
rect 134140 9980 134360 10020
rect 134140 9910 134150 9980
rect 134350 9910 134360 9980
rect 134140 9860 134360 9910
rect 134640 10090 134860 10140
rect 134640 10020 134650 10090
rect 134850 10020 134860 10090
rect 134640 9980 134860 10020
rect 134640 9910 134650 9980
rect 134850 9910 134860 9980
rect 134640 9860 134860 9910
rect 135140 10090 135360 10140
rect 135140 10020 135150 10090
rect 135350 10020 135360 10090
rect 135140 9980 135360 10020
rect 135140 9910 135150 9980
rect 135350 9910 135360 9980
rect 135140 9860 135360 9910
rect 135640 10090 135860 10140
rect 135640 10020 135650 10090
rect 135850 10020 135860 10090
rect 135640 9980 135860 10020
rect 135640 9910 135650 9980
rect 135850 9910 135860 9980
rect 135640 9860 135860 9910
rect 136140 10090 136360 10140
rect 136140 10020 136150 10090
rect 136350 10020 136360 10090
rect 136140 9980 136360 10020
rect 136140 9910 136150 9980
rect 136350 9910 136360 9980
rect 136140 9860 136360 9910
rect 136640 10090 136860 10140
rect 136640 10020 136650 10090
rect 136850 10020 136860 10090
rect 136640 9980 136860 10020
rect 136640 9910 136650 9980
rect 136850 9910 136860 9980
rect 136640 9860 136860 9910
rect 137140 10090 137360 10140
rect 137140 10020 137150 10090
rect 137350 10020 137360 10090
rect 137140 9980 137360 10020
rect 137140 9910 137150 9980
rect 137350 9910 137360 9980
rect 137140 9860 137360 9910
rect 137640 10090 137860 10140
rect 137640 10020 137650 10090
rect 137850 10020 137860 10090
rect 137640 9980 137860 10020
rect 137640 9910 137650 9980
rect 137850 9910 137860 9980
rect 137640 9860 137860 9910
rect 138140 10090 138360 10140
rect 138140 10020 138150 10090
rect 138350 10020 138360 10090
rect 138140 9980 138360 10020
rect 138140 9910 138150 9980
rect 138350 9910 138360 9980
rect 138140 9860 138360 9910
rect 138640 10090 138860 10140
rect 138640 10020 138650 10090
rect 138850 10020 138860 10090
rect 138640 9980 138860 10020
rect 138640 9910 138650 9980
rect 138850 9910 138860 9980
rect 138640 9860 138860 9910
rect 139140 10090 139360 10140
rect 139140 10020 139150 10090
rect 139350 10020 139360 10090
rect 139140 9980 139360 10020
rect 139140 9910 139150 9980
rect 139350 9910 139360 9980
rect 139140 9860 139360 9910
rect 139640 10090 139860 10140
rect 139640 10020 139650 10090
rect 139850 10020 139860 10090
rect 139640 9980 139860 10020
rect 139640 9910 139650 9980
rect 139850 9910 139860 9980
rect 139640 9860 139860 9910
rect 128000 9850 140000 9860
rect 128000 9650 128020 9850
rect 128090 9650 128410 9850
rect 128480 9650 128520 9850
rect 128590 9650 128910 9850
rect 128980 9650 129020 9850
rect 129090 9650 129410 9850
rect 129480 9650 129520 9850
rect 129590 9650 129910 9850
rect 129980 9650 130020 9850
rect 130090 9650 130410 9850
rect 130480 9650 130520 9850
rect 130590 9650 130910 9850
rect 130980 9650 131020 9850
rect 131090 9650 131410 9850
rect 131480 9650 131520 9850
rect 131590 9650 131910 9850
rect 131980 9650 132020 9850
rect 132090 9650 132410 9850
rect 132480 9650 132520 9850
rect 132590 9650 132910 9850
rect 132980 9650 133020 9850
rect 133090 9650 133410 9850
rect 133480 9650 133520 9850
rect 133590 9650 133910 9850
rect 133980 9650 134020 9850
rect 134090 9650 134410 9850
rect 134480 9650 134520 9850
rect 134590 9650 134910 9850
rect 134980 9650 135020 9850
rect 135090 9650 135410 9850
rect 135480 9650 135520 9850
rect 135590 9650 135910 9850
rect 135980 9650 136020 9850
rect 136090 9650 136410 9850
rect 136480 9650 136520 9850
rect 136590 9650 136910 9850
rect 136980 9650 137020 9850
rect 137090 9650 137410 9850
rect 137480 9650 137520 9850
rect 137590 9650 137910 9850
rect 137980 9650 138020 9850
rect 138090 9650 138410 9850
rect 138480 9650 138520 9850
rect 138590 9650 138910 9850
rect 138980 9650 139020 9850
rect 139090 9650 139410 9850
rect 139480 9650 139520 9850
rect 139590 9650 139910 9850
rect 139980 9650 140000 9850
rect 128000 9640 140000 9650
rect 128140 9590 128360 9640
rect 128140 9520 128150 9590
rect 128350 9520 128360 9590
rect 128140 9480 128360 9520
rect 128140 9410 128150 9480
rect 128350 9410 128360 9480
rect 128140 9360 128360 9410
rect 128640 9590 128860 9640
rect 128640 9520 128650 9590
rect 128850 9520 128860 9590
rect 128640 9480 128860 9520
rect 128640 9410 128650 9480
rect 128850 9410 128860 9480
rect 128640 9360 128860 9410
rect 129140 9590 129360 9640
rect 129140 9520 129150 9590
rect 129350 9520 129360 9590
rect 129140 9480 129360 9520
rect 129140 9410 129150 9480
rect 129350 9410 129360 9480
rect 129140 9360 129360 9410
rect 129640 9590 129860 9640
rect 129640 9520 129650 9590
rect 129850 9520 129860 9590
rect 129640 9480 129860 9520
rect 129640 9410 129650 9480
rect 129850 9410 129860 9480
rect 129640 9360 129860 9410
rect 130140 9590 130360 9640
rect 130140 9520 130150 9590
rect 130350 9520 130360 9590
rect 130140 9480 130360 9520
rect 130140 9410 130150 9480
rect 130350 9410 130360 9480
rect 130140 9360 130360 9410
rect 130640 9590 130860 9640
rect 130640 9520 130650 9590
rect 130850 9520 130860 9590
rect 130640 9480 130860 9520
rect 130640 9410 130650 9480
rect 130850 9410 130860 9480
rect 130640 9360 130860 9410
rect 131140 9590 131360 9640
rect 131140 9520 131150 9590
rect 131350 9520 131360 9590
rect 131140 9480 131360 9520
rect 131140 9410 131150 9480
rect 131350 9410 131360 9480
rect 131140 9360 131360 9410
rect 131640 9590 131860 9640
rect 131640 9520 131650 9590
rect 131850 9520 131860 9590
rect 131640 9480 131860 9520
rect 131640 9410 131650 9480
rect 131850 9410 131860 9480
rect 131640 9360 131860 9410
rect 132140 9590 132360 9640
rect 132140 9520 132150 9590
rect 132350 9520 132360 9590
rect 132140 9480 132360 9520
rect 132140 9410 132150 9480
rect 132350 9410 132360 9480
rect 132140 9360 132360 9410
rect 132640 9590 132860 9640
rect 132640 9520 132650 9590
rect 132850 9520 132860 9590
rect 132640 9480 132860 9520
rect 132640 9410 132650 9480
rect 132850 9410 132860 9480
rect 132640 9360 132860 9410
rect 133140 9590 133360 9640
rect 133140 9520 133150 9590
rect 133350 9520 133360 9590
rect 133140 9480 133360 9520
rect 133140 9410 133150 9480
rect 133350 9410 133360 9480
rect 133140 9360 133360 9410
rect 133640 9590 133860 9640
rect 133640 9520 133650 9590
rect 133850 9520 133860 9590
rect 133640 9480 133860 9520
rect 133640 9410 133650 9480
rect 133850 9410 133860 9480
rect 133640 9360 133860 9410
rect 134140 9590 134360 9640
rect 134140 9520 134150 9590
rect 134350 9520 134360 9590
rect 134140 9480 134360 9520
rect 134140 9410 134150 9480
rect 134350 9410 134360 9480
rect 134140 9360 134360 9410
rect 134640 9590 134860 9640
rect 134640 9520 134650 9590
rect 134850 9520 134860 9590
rect 134640 9480 134860 9520
rect 134640 9410 134650 9480
rect 134850 9410 134860 9480
rect 134640 9360 134860 9410
rect 135140 9590 135360 9640
rect 135140 9520 135150 9590
rect 135350 9520 135360 9590
rect 135140 9480 135360 9520
rect 135140 9410 135150 9480
rect 135350 9410 135360 9480
rect 135140 9360 135360 9410
rect 135640 9590 135860 9640
rect 135640 9520 135650 9590
rect 135850 9520 135860 9590
rect 135640 9480 135860 9520
rect 135640 9410 135650 9480
rect 135850 9410 135860 9480
rect 135640 9360 135860 9410
rect 136140 9590 136360 9640
rect 136140 9520 136150 9590
rect 136350 9520 136360 9590
rect 136140 9480 136360 9520
rect 136140 9410 136150 9480
rect 136350 9410 136360 9480
rect 136140 9360 136360 9410
rect 136640 9590 136860 9640
rect 136640 9520 136650 9590
rect 136850 9520 136860 9590
rect 136640 9480 136860 9520
rect 136640 9410 136650 9480
rect 136850 9410 136860 9480
rect 136640 9360 136860 9410
rect 137140 9590 137360 9640
rect 137140 9520 137150 9590
rect 137350 9520 137360 9590
rect 137140 9480 137360 9520
rect 137140 9410 137150 9480
rect 137350 9410 137360 9480
rect 137140 9360 137360 9410
rect 137640 9590 137860 9640
rect 137640 9520 137650 9590
rect 137850 9520 137860 9590
rect 137640 9480 137860 9520
rect 137640 9410 137650 9480
rect 137850 9410 137860 9480
rect 137640 9360 137860 9410
rect 138140 9590 138360 9640
rect 138140 9520 138150 9590
rect 138350 9520 138360 9590
rect 138140 9480 138360 9520
rect 138140 9410 138150 9480
rect 138350 9410 138360 9480
rect 138140 9360 138360 9410
rect 138640 9590 138860 9640
rect 138640 9520 138650 9590
rect 138850 9520 138860 9590
rect 138640 9480 138860 9520
rect 138640 9410 138650 9480
rect 138850 9410 138860 9480
rect 138640 9360 138860 9410
rect 139140 9590 139360 9640
rect 139140 9520 139150 9590
rect 139350 9520 139360 9590
rect 139140 9480 139360 9520
rect 139140 9410 139150 9480
rect 139350 9410 139360 9480
rect 139140 9360 139360 9410
rect 139640 9590 139860 9640
rect 139640 9520 139650 9590
rect 139850 9520 139860 9590
rect 139640 9480 139860 9520
rect 139640 9410 139650 9480
rect 139850 9410 139860 9480
rect 139640 9360 139860 9410
rect 128000 9350 140000 9360
rect 128000 9150 128020 9350
rect 128090 9150 128410 9350
rect 128480 9150 128520 9350
rect 128590 9150 128910 9350
rect 128980 9150 129020 9350
rect 129090 9150 129410 9350
rect 129480 9150 129520 9350
rect 129590 9150 129910 9350
rect 129980 9150 130020 9350
rect 130090 9150 130410 9350
rect 130480 9150 130520 9350
rect 130590 9150 130910 9350
rect 130980 9150 131020 9350
rect 131090 9150 131410 9350
rect 131480 9150 131520 9350
rect 131590 9150 131910 9350
rect 131980 9150 132020 9350
rect 132090 9150 132410 9350
rect 132480 9150 132520 9350
rect 132590 9150 132910 9350
rect 132980 9150 133020 9350
rect 133090 9150 133410 9350
rect 133480 9150 133520 9350
rect 133590 9150 133910 9350
rect 133980 9150 134020 9350
rect 134090 9150 134410 9350
rect 134480 9150 134520 9350
rect 134590 9150 134910 9350
rect 134980 9150 135020 9350
rect 135090 9150 135410 9350
rect 135480 9150 135520 9350
rect 135590 9150 135910 9350
rect 135980 9150 136020 9350
rect 136090 9150 136410 9350
rect 136480 9150 136520 9350
rect 136590 9150 136910 9350
rect 136980 9150 137020 9350
rect 137090 9150 137410 9350
rect 137480 9150 137520 9350
rect 137590 9150 137910 9350
rect 137980 9150 138020 9350
rect 138090 9150 138410 9350
rect 138480 9150 138520 9350
rect 138590 9150 138910 9350
rect 138980 9150 139020 9350
rect 139090 9150 139410 9350
rect 139480 9150 139520 9350
rect 139590 9150 139910 9350
rect 139980 9150 140000 9350
rect 128000 9140 140000 9150
rect 128140 9090 128360 9140
rect 128140 9020 128150 9090
rect 128350 9020 128360 9090
rect 128140 8980 128360 9020
rect 128140 8910 128150 8980
rect 128350 8910 128360 8980
rect 128140 8860 128360 8910
rect 128640 9090 128860 9140
rect 128640 9020 128650 9090
rect 128850 9020 128860 9090
rect 128640 8980 128860 9020
rect 128640 8910 128650 8980
rect 128850 8910 128860 8980
rect 128640 8860 128860 8910
rect 129140 9090 129360 9140
rect 129140 9020 129150 9090
rect 129350 9020 129360 9090
rect 129140 8980 129360 9020
rect 129140 8910 129150 8980
rect 129350 8910 129360 8980
rect 129140 8860 129360 8910
rect 129640 9090 129860 9140
rect 129640 9020 129650 9090
rect 129850 9020 129860 9090
rect 129640 8980 129860 9020
rect 129640 8910 129650 8980
rect 129850 8910 129860 8980
rect 129640 8860 129860 8910
rect 130140 9090 130360 9140
rect 130140 9020 130150 9090
rect 130350 9020 130360 9090
rect 130140 8980 130360 9020
rect 130140 8910 130150 8980
rect 130350 8910 130360 8980
rect 130140 8860 130360 8910
rect 130640 9090 130860 9140
rect 130640 9020 130650 9090
rect 130850 9020 130860 9090
rect 130640 8980 130860 9020
rect 130640 8910 130650 8980
rect 130850 8910 130860 8980
rect 130640 8860 130860 8910
rect 131140 9090 131360 9140
rect 131140 9020 131150 9090
rect 131350 9020 131360 9090
rect 131140 8980 131360 9020
rect 131140 8910 131150 8980
rect 131350 8910 131360 8980
rect 131140 8860 131360 8910
rect 131640 9090 131860 9140
rect 131640 9020 131650 9090
rect 131850 9020 131860 9090
rect 131640 8980 131860 9020
rect 131640 8910 131650 8980
rect 131850 8910 131860 8980
rect 131640 8860 131860 8910
rect 132140 9090 132360 9140
rect 132140 9020 132150 9090
rect 132350 9020 132360 9090
rect 132140 8980 132360 9020
rect 132140 8910 132150 8980
rect 132350 8910 132360 8980
rect 132140 8860 132360 8910
rect 132640 9090 132860 9140
rect 132640 9020 132650 9090
rect 132850 9020 132860 9090
rect 132640 8980 132860 9020
rect 132640 8910 132650 8980
rect 132850 8910 132860 8980
rect 132640 8860 132860 8910
rect 133140 9090 133360 9140
rect 133140 9020 133150 9090
rect 133350 9020 133360 9090
rect 133140 8980 133360 9020
rect 133140 8910 133150 8980
rect 133350 8910 133360 8980
rect 133140 8860 133360 8910
rect 133640 9090 133860 9140
rect 133640 9020 133650 9090
rect 133850 9020 133860 9090
rect 133640 8980 133860 9020
rect 133640 8910 133650 8980
rect 133850 8910 133860 8980
rect 133640 8860 133860 8910
rect 134140 9090 134360 9140
rect 134140 9020 134150 9090
rect 134350 9020 134360 9090
rect 134140 8980 134360 9020
rect 134140 8910 134150 8980
rect 134350 8910 134360 8980
rect 134140 8860 134360 8910
rect 134640 9090 134860 9140
rect 134640 9020 134650 9090
rect 134850 9020 134860 9090
rect 134640 8980 134860 9020
rect 134640 8910 134650 8980
rect 134850 8910 134860 8980
rect 134640 8860 134860 8910
rect 135140 9090 135360 9140
rect 135140 9020 135150 9090
rect 135350 9020 135360 9090
rect 135140 8980 135360 9020
rect 135140 8910 135150 8980
rect 135350 8910 135360 8980
rect 135140 8860 135360 8910
rect 135640 9090 135860 9140
rect 135640 9020 135650 9090
rect 135850 9020 135860 9090
rect 135640 8980 135860 9020
rect 135640 8910 135650 8980
rect 135850 8910 135860 8980
rect 135640 8860 135860 8910
rect 136140 9090 136360 9140
rect 136140 9020 136150 9090
rect 136350 9020 136360 9090
rect 136140 8980 136360 9020
rect 136140 8910 136150 8980
rect 136350 8910 136360 8980
rect 136140 8860 136360 8910
rect 136640 9090 136860 9140
rect 136640 9020 136650 9090
rect 136850 9020 136860 9090
rect 136640 8980 136860 9020
rect 136640 8910 136650 8980
rect 136850 8910 136860 8980
rect 136640 8860 136860 8910
rect 137140 9090 137360 9140
rect 137140 9020 137150 9090
rect 137350 9020 137360 9090
rect 137140 8980 137360 9020
rect 137140 8910 137150 8980
rect 137350 8910 137360 8980
rect 137140 8860 137360 8910
rect 137640 9090 137860 9140
rect 137640 9020 137650 9090
rect 137850 9020 137860 9090
rect 137640 8980 137860 9020
rect 137640 8910 137650 8980
rect 137850 8910 137860 8980
rect 137640 8860 137860 8910
rect 138140 9090 138360 9140
rect 138140 9020 138150 9090
rect 138350 9020 138360 9090
rect 138140 8980 138360 9020
rect 138140 8910 138150 8980
rect 138350 8910 138360 8980
rect 138140 8860 138360 8910
rect 138640 9090 138860 9140
rect 138640 9020 138650 9090
rect 138850 9020 138860 9090
rect 138640 8980 138860 9020
rect 138640 8910 138650 8980
rect 138850 8910 138860 8980
rect 138640 8860 138860 8910
rect 139140 9090 139360 9140
rect 139140 9020 139150 9090
rect 139350 9020 139360 9090
rect 139140 8980 139360 9020
rect 139140 8910 139150 8980
rect 139350 8910 139360 8980
rect 139140 8860 139360 8910
rect 139640 9090 139860 9140
rect 139640 9020 139650 9090
rect 139850 9020 139860 9090
rect 139640 8980 139860 9020
rect 139640 8910 139650 8980
rect 139850 8910 139860 8980
rect 139640 8860 139860 8910
rect 128000 8850 140000 8860
rect 128000 8650 128020 8850
rect 128090 8650 128410 8850
rect 128480 8650 128520 8850
rect 128590 8650 128910 8850
rect 128980 8650 129020 8850
rect 129090 8650 129410 8850
rect 129480 8650 129520 8850
rect 129590 8650 129910 8850
rect 129980 8650 130020 8850
rect 130090 8650 130410 8850
rect 130480 8650 130520 8850
rect 130590 8650 130910 8850
rect 130980 8650 131020 8850
rect 131090 8650 131410 8850
rect 131480 8650 131520 8850
rect 131590 8650 131910 8850
rect 131980 8650 132020 8850
rect 132090 8650 132410 8850
rect 132480 8650 132520 8850
rect 132590 8650 132910 8850
rect 132980 8650 133020 8850
rect 133090 8650 133410 8850
rect 133480 8650 133520 8850
rect 133590 8650 133910 8850
rect 133980 8650 134020 8850
rect 134090 8650 134410 8850
rect 134480 8650 134520 8850
rect 134590 8650 134910 8850
rect 134980 8650 135020 8850
rect 135090 8650 135410 8850
rect 135480 8650 135520 8850
rect 135590 8650 135910 8850
rect 135980 8650 136020 8850
rect 136090 8650 136410 8850
rect 136480 8650 136520 8850
rect 136590 8650 136910 8850
rect 136980 8650 137020 8850
rect 137090 8650 137410 8850
rect 137480 8650 137520 8850
rect 137590 8650 137910 8850
rect 137980 8650 138020 8850
rect 138090 8650 138410 8850
rect 138480 8650 138520 8850
rect 138590 8650 138910 8850
rect 138980 8650 139020 8850
rect 139090 8650 139410 8850
rect 139480 8650 139520 8850
rect 139590 8650 139910 8850
rect 139980 8650 140000 8850
rect 128000 8640 140000 8650
rect 128140 8590 128360 8640
rect 128140 8520 128150 8590
rect 128350 8520 128360 8590
rect 128140 8480 128360 8520
rect 128140 8410 128150 8480
rect 128350 8410 128360 8480
rect 128140 8360 128360 8410
rect 128640 8590 128860 8640
rect 128640 8520 128650 8590
rect 128850 8520 128860 8590
rect 128640 8480 128860 8520
rect 128640 8410 128650 8480
rect 128850 8410 128860 8480
rect 128640 8360 128860 8410
rect 129140 8590 129360 8640
rect 129140 8520 129150 8590
rect 129350 8520 129360 8590
rect 129140 8480 129360 8520
rect 129140 8410 129150 8480
rect 129350 8410 129360 8480
rect 129140 8360 129360 8410
rect 129640 8590 129860 8640
rect 129640 8520 129650 8590
rect 129850 8520 129860 8590
rect 129640 8480 129860 8520
rect 129640 8410 129650 8480
rect 129850 8410 129860 8480
rect 129640 8360 129860 8410
rect 130140 8590 130360 8640
rect 130140 8520 130150 8590
rect 130350 8520 130360 8590
rect 130140 8480 130360 8520
rect 130140 8410 130150 8480
rect 130350 8410 130360 8480
rect 130140 8360 130360 8410
rect 130640 8590 130860 8640
rect 130640 8520 130650 8590
rect 130850 8520 130860 8590
rect 130640 8480 130860 8520
rect 130640 8410 130650 8480
rect 130850 8410 130860 8480
rect 130640 8360 130860 8410
rect 131140 8590 131360 8640
rect 131140 8520 131150 8590
rect 131350 8520 131360 8590
rect 131140 8480 131360 8520
rect 131140 8410 131150 8480
rect 131350 8410 131360 8480
rect 131140 8360 131360 8410
rect 131640 8590 131860 8640
rect 131640 8520 131650 8590
rect 131850 8520 131860 8590
rect 131640 8480 131860 8520
rect 131640 8410 131650 8480
rect 131850 8410 131860 8480
rect 131640 8360 131860 8410
rect 132140 8590 132360 8640
rect 132140 8520 132150 8590
rect 132350 8520 132360 8590
rect 132140 8480 132360 8520
rect 132140 8410 132150 8480
rect 132350 8410 132360 8480
rect 132140 8360 132360 8410
rect 132640 8590 132860 8640
rect 132640 8520 132650 8590
rect 132850 8520 132860 8590
rect 132640 8480 132860 8520
rect 132640 8410 132650 8480
rect 132850 8410 132860 8480
rect 132640 8360 132860 8410
rect 133140 8590 133360 8640
rect 133140 8520 133150 8590
rect 133350 8520 133360 8590
rect 133140 8480 133360 8520
rect 133140 8410 133150 8480
rect 133350 8410 133360 8480
rect 133140 8360 133360 8410
rect 133640 8590 133860 8640
rect 133640 8520 133650 8590
rect 133850 8520 133860 8590
rect 133640 8480 133860 8520
rect 133640 8410 133650 8480
rect 133850 8410 133860 8480
rect 133640 8360 133860 8410
rect 134140 8590 134360 8640
rect 134140 8520 134150 8590
rect 134350 8520 134360 8590
rect 134140 8480 134360 8520
rect 134140 8410 134150 8480
rect 134350 8410 134360 8480
rect 134140 8360 134360 8410
rect 134640 8590 134860 8640
rect 134640 8520 134650 8590
rect 134850 8520 134860 8590
rect 134640 8480 134860 8520
rect 134640 8410 134650 8480
rect 134850 8410 134860 8480
rect 134640 8360 134860 8410
rect 135140 8590 135360 8640
rect 135140 8520 135150 8590
rect 135350 8520 135360 8590
rect 135140 8480 135360 8520
rect 135140 8410 135150 8480
rect 135350 8410 135360 8480
rect 135140 8360 135360 8410
rect 135640 8590 135860 8640
rect 135640 8520 135650 8590
rect 135850 8520 135860 8590
rect 135640 8480 135860 8520
rect 135640 8410 135650 8480
rect 135850 8410 135860 8480
rect 135640 8360 135860 8410
rect 136140 8590 136360 8640
rect 136140 8520 136150 8590
rect 136350 8520 136360 8590
rect 136140 8480 136360 8520
rect 136140 8410 136150 8480
rect 136350 8410 136360 8480
rect 136140 8360 136360 8410
rect 136640 8590 136860 8640
rect 136640 8520 136650 8590
rect 136850 8520 136860 8590
rect 136640 8480 136860 8520
rect 136640 8410 136650 8480
rect 136850 8410 136860 8480
rect 136640 8360 136860 8410
rect 137140 8590 137360 8640
rect 137140 8520 137150 8590
rect 137350 8520 137360 8590
rect 137140 8480 137360 8520
rect 137140 8410 137150 8480
rect 137350 8410 137360 8480
rect 137140 8360 137360 8410
rect 137640 8590 137860 8640
rect 137640 8520 137650 8590
rect 137850 8520 137860 8590
rect 137640 8480 137860 8520
rect 137640 8410 137650 8480
rect 137850 8410 137860 8480
rect 137640 8360 137860 8410
rect 138140 8590 138360 8640
rect 138140 8520 138150 8590
rect 138350 8520 138360 8590
rect 138140 8480 138360 8520
rect 138140 8410 138150 8480
rect 138350 8410 138360 8480
rect 138140 8360 138360 8410
rect 138640 8590 138860 8640
rect 138640 8520 138650 8590
rect 138850 8520 138860 8590
rect 138640 8480 138860 8520
rect 138640 8410 138650 8480
rect 138850 8410 138860 8480
rect 138640 8360 138860 8410
rect 139140 8590 139360 8640
rect 139140 8520 139150 8590
rect 139350 8520 139360 8590
rect 139140 8480 139360 8520
rect 139140 8410 139150 8480
rect 139350 8410 139360 8480
rect 139140 8360 139360 8410
rect 139640 8590 139860 8640
rect 139640 8520 139650 8590
rect 139850 8520 139860 8590
rect 139640 8480 139860 8520
rect 139640 8410 139650 8480
rect 139850 8410 139860 8480
rect 139640 8360 139860 8410
rect 128000 8350 140000 8360
rect 128000 8150 128020 8350
rect 128090 8150 128410 8350
rect 128480 8150 128520 8350
rect 128590 8150 128910 8350
rect 128980 8150 129020 8350
rect 129090 8150 129410 8350
rect 129480 8150 129520 8350
rect 129590 8150 129910 8350
rect 129980 8150 130020 8350
rect 130090 8150 130410 8350
rect 130480 8150 130520 8350
rect 130590 8150 130910 8350
rect 130980 8150 131020 8350
rect 131090 8150 131410 8350
rect 131480 8150 131520 8350
rect 131590 8150 131910 8350
rect 131980 8150 132020 8350
rect 132090 8150 132410 8350
rect 132480 8150 132520 8350
rect 132590 8150 132910 8350
rect 132980 8150 133020 8350
rect 133090 8150 133410 8350
rect 133480 8150 133520 8350
rect 133590 8150 133910 8350
rect 133980 8150 134020 8350
rect 134090 8150 134410 8350
rect 134480 8150 134520 8350
rect 134590 8150 134910 8350
rect 134980 8150 135020 8350
rect 135090 8150 135410 8350
rect 135480 8150 135520 8350
rect 135590 8150 135910 8350
rect 135980 8150 136020 8350
rect 136090 8150 136410 8350
rect 136480 8150 136520 8350
rect 136590 8150 136910 8350
rect 136980 8150 137020 8350
rect 137090 8150 137410 8350
rect 137480 8150 137520 8350
rect 137590 8150 137910 8350
rect 137980 8150 138020 8350
rect 138090 8150 138410 8350
rect 138480 8150 138520 8350
rect 138590 8150 138910 8350
rect 138980 8150 139020 8350
rect 139090 8150 139410 8350
rect 139480 8150 139520 8350
rect 139590 8150 139910 8350
rect 139980 8150 140000 8350
rect 128000 8140 140000 8150
rect 128140 8090 128360 8140
rect 128140 8020 128150 8090
rect 128350 8020 128360 8090
rect 128140 7980 128360 8020
rect 128140 7910 128150 7980
rect 128350 7910 128360 7980
rect 128140 7860 128360 7910
rect 128640 8090 128860 8140
rect 128640 8020 128650 8090
rect 128850 8020 128860 8090
rect 128640 7980 128860 8020
rect 128640 7910 128650 7980
rect 128850 7910 128860 7980
rect 128640 7860 128860 7910
rect 129140 8090 129360 8140
rect 129140 8020 129150 8090
rect 129350 8020 129360 8090
rect 129140 7980 129360 8020
rect 129140 7910 129150 7980
rect 129350 7910 129360 7980
rect 129140 7860 129360 7910
rect 129640 8090 129860 8140
rect 129640 8020 129650 8090
rect 129850 8020 129860 8090
rect 129640 7980 129860 8020
rect 129640 7910 129650 7980
rect 129850 7910 129860 7980
rect 129640 7860 129860 7910
rect 130140 8090 130360 8140
rect 130140 8020 130150 8090
rect 130350 8020 130360 8090
rect 130140 7980 130360 8020
rect 130140 7910 130150 7980
rect 130350 7910 130360 7980
rect 130140 7860 130360 7910
rect 130640 8090 130860 8140
rect 130640 8020 130650 8090
rect 130850 8020 130860 8090
rect 130640 7980 130860 8020
rect 130640 7910 130650 7980
rect 130850 7910 130860 7980
rect 130640 7860 130860 7910
rect 131140 8090 131360 8140
rect 131140 8020 131150 8090
rect 131350 8020 131360 8090
rect 131140 7980 131360 8020
rect 131140 7910 131150 7980
rect 131350 7910 131360 7980
rect 131140 7860 131360 7910
rect 131640 8090 131860 8140
rect 131640 8020 131650 8090
rect 131850 8020 131860 8090
rect 131640 7980 131860 8020
rect 131640 7910 131650 7980
rect 131850 7910 131860 7980
rect 131640 7860 131860 7910
rect 132140 8090 132360 8140
rect 132140 8020 132150 8090
rect 132350 8020 132360 8090
rect 132140 7980 132360 8020
rect 132140 7910 132150 7980
rect 132350 7910 132360 7980
rect 132140 7860 132360 7910
rect 132640 8090 132860 8140
rect 132640 8020 132650 8090
rect 132850 8020 132860 8090
rect 132640 7980 132860 8020
rect 132640 7910 132650 7980
rect 132850 7910 132860 7980
rect 132640 7860 132860 7910
rect 133140 8090 133360 8140
rect 133140 8020 133150 8090
rect 133350 8020 133360 8090
rect 133140 7980 133360 8020
rect 133140 7910 133150 7980
rect 133350 7910 133360 7980
rect 133140 7860 133360 7910
rect 133640 8090 133860 8140
rect 133640 8020 133650 8090
rect 133850 8020 133860 8090
rect 133640 7980 133860 8020
rect 133640 7910 133650 7980
rect 133850 7910 133860 7980
rect 133640 7860 133860 7910
rect 134140 8090 134360 8140
rect 134140 8020 134150 8090
rect 134350 8020 134360 8090
rect 134140 7980 134360 8020
rect 134140 7910 134150 7980
rect 134350 7910 134360 7980
rect 134140 7860 134360 7910
rect 134640 8090 134860 8140
rect 134640 8020 134650 8090
rect 134850 8020 134860 8090
rect 134640 7980 134860 8020
rect 134640 7910 134650 7980
rect 134850 7910 134860 7980
rect 134640 7860 134860 7910
rect 135140 8090 135360 8140
rect 135140 8020 135150 8090
rect 135350 8020 135360 8090
rect 135140 7980 135360 8020
rect 135140 7910 135150 7980
rect 135350 7910 135360 7980
rect 135140 7860 135360 7910
rect 135640 8090 135860 8140
rect 135640 8020 135650 8090
rect 135850 8020 135860 8090
rect 135640 7980 135860 8020
rect 135640 7910 135650 7980
rect 135850 7910 135860 7980
rect 135640 7860 135860 7910
rect 136140 8090 136360 8140
rect 136140 8020 136150 8090
rect 136350 8020 136360 8090
rect 136140 7980 136360 8020
rect 136140 7910 136150 7980
rect 136350 7910 136360 7980
rect 136140 7860 136360 7910
rect 136640 8090 136860 8140
rect 136640 8020 136650 8090
rect 136850 8020 136860 8090
rect 136640 7980 136860 8020
rect 136640 7910 136650 7980
rect 136850 7910 136860 7980
rect 136640 7860 136860 7910
rect 137140 8090 137360 8140
rect 137140 8020 137150 8090
rect 137350 8020 137360 8090
rect 137140 7980 137360 8020
rect 137140 7910 137150 7980
rect 137350 7910 137360 7980
rect 137140 7860 137360 7910
rect 137640 8090 137860 8140
rect 137640 8020 137650 8090
rect 137850 8020 137860 8090
rect 137640 7980 137860 8020
rect 137640 7910 137650 7980
rect 137850 7910 137860 7980
rect 137640 7860 137860 7910
rect 138140 8090 138360 8140
rect 138140 8020 138150 8090
rect 138350 8020 138360 8090
rect 138140 7980 138360 8020
rect 138140 7910 138150 7980
rect 138350 7910 138360 7980
rect 138140 7860 138360 7910
rect 138640 8090 138860 8140
rect 138640 8020 138650 8090
rect 138850 8020 138860 8090
rect 138640 7980 138860 8020
rect 138640 7910 138650 7980
rect 138850 7910 138860 7980
rect 138640 7860 138860 7910
rect 139140 8090 139360 8140
rect 139140 8020 139150 8090
rect 139350 8020 139360 8090
rect 139140 7980 139360 8020
rect 139140 7910 139150 7980
rect 139350 7910 139360 7980
rect 139140 7860 139360 7910
rect 139640 8090 139860 8140
rect 139640 8020 139650 8090
rect 139850 8020 139860 8090
rect 139640 7980 139860 8020
rect 139640 7910 139650 7980
rect 139850 7910 139860 7980
rect 139640 7860 139860 7910
rect 128000 7850 140000 7860
rect 128000 7650 128020 7850
rect 128090 7650 128410 7850
rect 128480 7650 128520 7850
rect 128590 7650 128910 7850
rect 128980 7650 129020 7850
rect 129090 7650 129410 7850
rect 129480 7650 129520 7850
rect 129590 7650 129910 7850
rect 129980 7650 130020 7850
rect 130090 7650 130410 7850
rect 130480 7650 130520 7850
rect 130590 7650 130910 7850
rect 130980 7650 131020 7850
rect 131090 7650 131410 7850
rect 131480 7650 131520 7850
rect 131590 7650 131910 7850
rect 131980 7650 132020 7850
rect 132090 7650 132410 7850
rect 132480 7650 132520 7850
rect 132590 7650 132910 7850
rect 132980 7650 133020 7850
rect 133090 7650 133410 7850
rect 133480 7650 133520 7850
rect 133590 7650 133910 7850
rect 133980 7650 134020 7850
rect 134090 7650 134410 7850
rect 134480 7650 134520 7850
rect 134590 7650 134910 7850
rect 134980 7650 135020 7850
rect 135090 7650 135410 7850
rect 135480 7650 135520 7850
rect 135590 7650 135910 7850
rect 135980 7650 136020 7850
rect 136090 7650 136410 7850
rect 136480 7650 136520 7850
rect 136590 7650 136910 7850
rect 136980 7650 137020 7850
rect 137090 7650 137410 7850
rect 137480 7650 137520 7850
rect 137590 7650 137910 7850
rect 137980 7650 138020 7850
rect 138090 7650 138410 7850
rect 138480 7650 138520 7850
rect 138590 7650 138910 7850
rect 138980 7650 139020 7850
rect 139090 7650 139410 7850
rect 139480 7650 139520 7850
rect 139590 7650 139910 7850
rect 139980 7650 140000 7850
rect 128000 7640 140000 7650
rect 128140 7590 128360 7640
rect 128140 7520 128150 7590
rect 128350 7520 128360 7590
rect 128140 7480 128360 7520
rect 128140 7410 128150 7480
rect 128350 7410 128360 7480
rect 128140 7360 128360 7410
rect 128640 7590 128860 7640
rect 128640 7520 128650 7590
rect 128850 7520 128860 7590
rect 128640 7480 128860 7520
rect 128640 7410 128650 7480
rect 128850 7410 128860 7480
rect 128640 7360 128860 7410
rect 129140 7590 129360 7640
rect 129140 7520 129150 7590
rect 129350 7520 129360 7590
rect 129140 7480 129360 7520
rect 129140 7410 129150 7480
rect 129350 7410 129360 7480
rect 129140 7360 129360 7410
rect 129640 7590 129860 7640
rect 129640 7520 129650 7590
rect 129850 7520 129860 7590
rect 129640 7480 129860 7520
rect 129640 7410 129650 7480
rect 129850 7410 129860 7480
rect 129640 7360 129860 7410
rect 130140 7590 130360 7640
rect 130140 7520 130150 7590
rect 130350 7520 130360 7590
rect 130140 7480 130360 7520
rect 130140 7410 130150 7480
rect 130350 7410 130360 7480
rect 130140 7360 130360 7410
rect 130640 7590 130860 7640
rect 130640 7520 130650 7590
rect 130850 7520 130860 7590
rect 130640 7480 130860 7520
rect 130640 7410 130650 7480
rect 130850 7410 130860 7480
rect 130640 7360 130860 7410
rect 131140 7590 131360 7640
rect 131140 7520 131150 7590
rect 131350 7520 131360 7590
rect 131140 7480 131360 7520
rect 131140 7410 131150 7480
rect 131350 7410 131360 7480
rect 131140 7360 131360 7410
rect 131640 7590 131860 7640
rect 131640 7520 131650 7590
rect 131850 7520 131860 7590
rect 131640 7480 131860 7520
rect 131640 7410 131650 7480
rect 131850 7410 131860 7480
rect 131640 7360 131860 7410
rect 132140 7590 132360 7640
rect 132140 7520 132150 7590
rect 132350 7520 132360 7590
rect 132140 7480 132360 7520
rect 132140 7410 132150 7480
rect 132350 7410 132360 7480
rect 132140 7360 132360 7410
rect 132640 7590 132860 7640
rect 132640 7520 132650 7590
rect 132850 7520 132860 7590
rect 132640 7480 132860 7520
rect 132640 7410 132650 7480
rect 132850 7410 132860 7480
rect 132640 7360 132860 7410
rect 133140 7590 133360 7640
rect 133140 7520 133150 7590
rect 133350 7520 133360 7590
rect 133140 7480 133360 7520
rect 133140 7410 133150 7480
rect 133350 7410 133360 7480
rect 133140 7360 133360 7410
rect 133640 7590 133860 7640
rect 133640 7520 133650 7590
rect 133850 7520 133860 7590
rect 133640 7480 133860 7520
rect 133640 7410 133650 7480
rect 133850 7410 133860 7480
rect 133640 7360 133860 7410
rect 134140 7590 134360 7640
rect 134140 7520 134150 7590
rect 134350 7520 134360 7590
rect 134140 7480 134360 7520
rect 134140 7410 134150 7480
rect 134350 7410 134360 7480
rect 134140 7360 134360 7410
rect 134640 7590 134860 7640
rect 134640 7520 134650 7590
rect 134850 7520 134860 7590
rect 134640 7480 134860 7520
rect 134640 7410 134650 7480
rect 134850 7410 134860 7480
rect 134640 7360 134860 7410
rect 135140 7590 135360 7640
rect 135140 7520 135150 7590
rect 135350 7520 135360 7590
rect 135140 7480 135360 7520
rect 135140 7410 135150 7480
rect 135350 7410 135360 7480
rect 135140 7360 135360 7410
rect 135640 7590 135860 7640
rect 135640 7520 135650 7590
rect 135850 7520 135860 7590
rect 135640 7480 135860 7520
rect 135640 7410 135650 7480
rect 135850 7410 135860 7480
rect 135640 7360 135860 7410
rect 136140 7590 136360 7640
rect 136140 7520 136150 7590
rect 136350 7520 136360 7590
rect 136140 7480 136360 7520
rect 136140 7410 136150 7480
rect 136350 7410 136360 7480
rect 136140 7360 136360 7410
rect 136640 7590 136860 7640
rect 136640 7520 136650 7590
rect 136850 7520 136860 7590
rect 136640 7480 136860 7520
rect 136640 7410 136650 7480
rect 136850 7410 136860 7480
rect 136640 7360 136860 7410
rect 137140 7590 137360 7640
rect 137140 7520 137150 7590
rect 137350 7520 137360 7590
rect 137140 7480 137360 7520
rect 137140 7410 137150 7480
rect 137350 7410 137360 7480
rect 137140 7360 137360 7410
rect 137640 7590 137860 7640
rect 137640 7520 137650 7590
rect 137850 7520 137860 7590
rect 137640 7480 137860 7520
rect 137640 7410 137650 7480
rect 137850 7410 137860 7480
rect 137640 7360 137860 7410
rect 138140 7590 138360 7640
rect 138140 7520 138150 7590
rect 138350 7520 138360 7590
rect 138140 7480 138360 7520
rect 138140 7410 138150 7480
rect 138350 7410 138360 7480
rect 138140 7360 138360 7410
rect 138640 7590 138860 7640
rect 138640 7520 138650 7590
rect 138850 7520 138860 7590
rect 138640 7480 138860 7520
rect 138640 7410 138650 7480
rect 138850 7410 138860 7480
rect 138640 7360 138860 7410
rect 139140 7590 139360 7640
rect 139140 7520 139150 7590
rect 139350 7520 139360 7590
rect 139140 7480 139360 7520
rect 139140 7410 139150 7480
rect 139350 7410 139360 7480
rect 139140 7360 139360 7410
rect 139640 7590 139860 7640
rect 139640 7520 139650 7590
rect 139850 7520 139860 7590
rect 139640 7480 139860 7520
rect 139640 7410 139650 7480
rect 139850 7410 139860 7480
rect 139640 7360 139860 7410
rect 128000 7350 140000 7360
rect 128000 7150 128020 7350
rect 128090 7150 128410 7350
rect 128480 7150 128520 7350
rect 128590 7150 128910 7350
rect 128980 7150 129020 7350
rect 129090 7150 129410 7350
rect 129480 7150 129520 7350
rect 129590 7150 129910 7350
rect 129980 7150 130020 7350
rect 130090 7150 130410 7350
rect 130480 7150 130520 7350
rect 130590 7150 130910 7350
rect 130980 7150 131020 7350
rect 131090 7150 131410 7350
rect 131480 7150 131520 7350
rect 131590 7150 131910 7350
rect 131980 7150 132020 7350
rect 132090 7150 132410 7350
rect 132480 7150 132520 7350
rect 132590 7150 132910 7350
rect 132980 7150 133020 7350
rect 133090 7150 133410 7350
rect 133480 7150 133520 7350
rect 133590 7150 133910 7350
rect 133980 7150 134020 7350
rect 134090 7150 134410 7350
rect 134480 7150 134520 7350
rect 134590 7150 134910 7350
rect 134980 7150 135020 7350
rect 135090 7150 135410 7350
rect 135480 7150 135520 7350
rect 135590 7150 135910 7350
rect 135980 7150 136020 7350
rect 136090 7150 136410 7350
rect 136480 7150 136520 7350
rect 136590 7150 136910 7350
rect 136980 7150 137020 7350
rect 137090 7150 137410 7350
rect 137480 7150 137520 7350
rect 137590 7150 137910 7350
rect 137980 7150 138020 7350
rect 138090 7150 138410 7350
rect 138480 7150 138520 7350
rect 138590 7150 138910 7350
rect 138980 7150 139020 7350
rect 139090 7150 139410 7350
rect 139480 7150 139520 7350
rect 139590 7150 139910 7350
rect 139980 7150 140000 7350
rect 128000 7140 140000 7150
rect 128140 7090 128360 7140
rect 128140 7020 128150 7090
rect 128350 7020 128360 7090
rect 128140 6980 128360 7020
rect 128140 6910 128150 6980
rect 128350 6910 128360 6980
rect 128140 6860 128360 6910
rect 128640 7090 128860 7140
rect 128640 7020 128650 7090
rect 128850 7020 128860 7090
rect 128640 6980 128860 7020
rect 128640 6910 128650 6980
rect 128850 6910 128860 6980
rect 128640 6860 128860 6910
rect 129140 7090 129360 7140
rect 129140 7020 129150 7090
rect 129350 7020 129360 7090
rect 129140 6980 129360 7020
rect 129140 6910 129150 6980
rect 129350 6910 129360 6980
rect 129140 6860 129360 6910
rect 129640 7090 129860 7140
rect 129640 7020 129650 7090
rect 129850 7020 129860 7090
rect 129640 6980 129860 7020
rect 129640 6910 129650 6980
rect 129850 6910 129860 6980
rect 129640 6860 129860 6910
rect 130140 7090 130360 7140
rect 130140 7020 130150 7090
rect 130350 7020 130360 7090
rect 130140 6980 130360 7020
rect 130140 6910 130150 6980
rect 130350 6910 130360 6980
rect 130140 6860 130360 6910
rect 130640 7090 130860 7140
rect 130640 7020 130650 7090
rect 130850 7020 130860 7090
rect 130640 6980 130860 7020
rect 130640 6910 130650 6980
rect 130850 6910 130860 6980
rect 130640 6860 130860 6910
rect 131140 7090 131360 7140
rect 131140 7020 131150 7090
rect 131350 7020 131360 7090
rect 131140 6980 131360 7020
rect 131140 6910 131150 6980
rect 131350 6910 131360 6980
rect 131140 6860 131360 6910
rect 131640 7090 131860 7140
rect 131640 7020 131650 7090
rect 131850 7020 131860 7090
rect 131640 6980 131860 7020
rect 131640 6910 131650 6980
rect 131850 6910 131860 6980
rect 131640 6860 131860 6910
rect 132140 7090 132360 7140
rect 132140 7020 132150 7090
rect 132350 7020 132360 7090
rect 132140 6980 132360 7020
rect 132140 6910 132150 6980
rect 132350 6910 132360 6980
rect 132140 6860 132360 6910
rect 132640 7090 132860 7140
rect 132640 7020 132650 7090
rect 132850 7020 132860 7090
rect 132640 6980 132860 7020
rect 132640 6910 132650 6980
rect 132850 6910 132860 6980
rect 132640 6860 132860 6910
rect 133140 7090 133360 7140
rect 133140 7020 133150 7090
rect 133350 7020 133360 7090
rect 133140 6980 133360 7020
rect 133140 6910 133150 6980
rect 133350 6910 133360 6980
rect 133140 6860 133360 6910
rect 133640 7090 133860 7140
rect 133640 7020 133650 7090
rect 133850 7020 133860 7090
rect 133640 6980 133860 7020
rect 133640 6910 133650 6980
rect 133850 6910 133860 6980
rect 133640 6860 133860 6910
rect 134140 7090 134360 7140
rect 134140 7020 134150 7090
rect 134350 7020 134360 7090
rect 134140 6980 134360 7020
rect 134140 6910 134150 6980
rect 134350 6910 134360 6980
rect 134140 6860 134360 6910
rect 134640 7090 134860 7140
rect 134640 7020 134650 7090
rect 134850 7020 134860 7090
rect 134640 6980 134860 7020
rect 134640 6910 134650 6980
rect 134850 6910 134860 6980
rect 134640 6860 134860 6910
rect 135140 7090 135360 7140
rect 135140 7020 135150 7090
rect 135350 7020 135360 7090
rect 135140 6980 135360 7020
rect 135140 6910 135150 6980
rect 135350 6910 135360 6980
rect 135140 6860 135360 6910
rect 135640 7090 135860 7140
rect 135640 7020 135650 7090
rect 135850 7020 135860 7090
rect 135640 6980 135860 7020
rect 135640 6910 135650 6980
rect 135850 6910 135860 6980
rect 135640 6860 135860 6910
rect 136140 7090 136360 7140
rect 136140 7020 136150 7090
rect 136350 7020 136360 7090
rect 136140 6980 136360 7020
rect 136140 6910 136150 6980
rect 136350 6910 136360 6980
rect 136140 6860 136360 6910
rect 136640 7090 136860 7140
rect 136640 7020 136650 7090
rect 136850 7020 136860 7090
rect 136640 6980 136860 7020
rect 136640 6910 136650 6980
rect 136850 6910 136860 6980
rect 136640 6860 136860 6910
rect 137140 7090 137360 7140
rect 137140 7020 137150 7090
rect 137350 7020 137360 7090
rect 137140 6980 137360 7020
rect 137140 6910 137150 6980
rect 137350 6910 137360 6980
rect 137140 6860 137360 6910
rect 137640 7090 137860 7140
rect 137640 7020 137650 7090
rect 137850 7020 137860 7090
rect 137640 6980 137860 7020
rect 137640 6910 137650 6980
rect 137850 6910 137860 6980
rect 137640 6860 137860 6910
rect 138140 7090 138360 7140
rect 138140 7020 138150 7090
rect 138350 7020 138360 7090
rect 138140 6980 138360 7020
rect 138140 6910 138150 6980
rect 138350 6910 138360 6980
rect 138140 6860 138360 6910
rect 138640 7090 138860 7140
rect 138640 7020 138650 7090
rect 138850 7020 138860 7090
rect 138640 6980 138860 7020
rect 138640 6910 138650 6980
rect 138850 6910 138860 6980
rect 138640 6860 138860 6910
rect 139140 7090 139360 7140
rect 139140 7020 139150 7090
rect 139350 7020 139360 7090
rect 139140 6980 139360 7020
rect 139140 6910 139150 6980
rect 139350 6910 139360 6980
rect 139140 6860 139360 6910
rect 139640 7090 139860 7140
rect 139640 7020 139650 7090
rect 139850 7020 139860 7090
rect 139640 6980 139860 7020
rect 139640 6910 139650 6980
rect 139850 6910 139860 6980
rect 139640 6860 139860 6910
rect 128000 6850 140000 6860
rect 128000 6650 128020 6850
rect 128090 6650 128410 6850
rect 128480 6650 128520 6850
rect 128590 6650 128910 6850
rect 128980 6650 129020 6850
rect 129090 6650 129410 6850
rect 129480 6650 129520 6850
rect 129590 6650 129910 6850
rect 129980 6650 130020 6850
rect 130090 6650 130410 6850
rect 130480 6650 130520 6850
rect 130590 6650 130910 6850
rect 130980 6650 131020 6850
rect 131090 6650 131410 6850
rect 131480 6650 131520 6850
rect 131590 6650 131910 6850
rect 131980 6650 132020 6850
rect 132090 6650 132410 6850
rect 132480 6650 132520 6850
rect 132590 6650 132910 6850
rect 132980 6650 133020 6850
rect 133090 6650 133410 6850
rect 133480 6650 133520 6850
rect 133590 6650 133910 6850
rect 133980 6650 134020 6850
rect 134090 6650 134410 6850
rect 134480 6650 134520 6850
rect 134590 6650 134910 6850
rect 134980 6650 135020 6850
rect 135090 6650 135410 6850
rect 135480 6650 135520 6850
rect 135590 6650 135910 6850
rect 135980 6650 136020 6850
rect 136090 6650 136410 6850
rect 136480 6650 136520 6850
rect 136590 6650 136910 6850
rect 136980 6650 137020 6850
rect 137090 6650 137410 6850
rect 137480 6650 137520 6850
rect 137590 6650 137910 6850
rect 137980 6650 138020 6850
rect 138090 6650 138410 6850
rect 138480 6650 138520 6850
rect 138590 6650 138910 6850
rect 138980 6650 139020 6850
rect 139090 6650 139410 6850
rect 139480 6650 139520 6850
rect 139590 6650 139910 6850
rect 139980 6650 140000 6850
rect 128000 6640 140000 6650
rect 128140 6590 128360 6640
rect 128140 6520 128150 6590
rect 128350 6520 128360 6590
rect 128140 6480 128360 6520
rect 128140 6410 128150 6480
rect 128350 6410 128360 6480
rect 128140 6360 128360 6410
rect 128640 6590 128860 6640
rect 128640 6520 128650 6590
rect 128850 6520 128860 6590
rect 128640 6480 128860 6520
rect 128640 6410 128650 6480
rect 128850 6410 128860 6480
rect 128640 6360 128860 6410
rect 129140 6590 129360 6640
rect 129140 6520 129150 6590
rect 129350 6520 129360 6590
rect 129140 6480 129360 6520
rect 129140 6410 129150 6480
rect 129350 6410 129360 6480
rect 129140 6360 129360 6410
rect 129640 6590 129860 6640
rect 129640 6520 129650 6590
rect 129850 6520 129860 6590
rect 129640 6480 129860 6520
rect 129640 6410 129650 6480
rect 129850 6410 129860 6480
rect 129640 6360 129860 6410
rect 130140 6590 130360 6640
rect 130140 6520 130150 6590
rect 130350 6520 130360 6590
rect 130140 6480 130360 6520
rect 130140 6410 130150 6480
rect 130350 6410 130360 6480
rect 130140 6360 130360 6410
rect 130640 6590 130860 6640
rect 130640 6520 130650 6590
rect 130850 6520 130860 6590
rect 130640 6480 130860 6520
rect 130640 6410 130650 6480
rect 130850 6410 130860 6480
rect 130640 6360 130860 6410
rect 131140 6590 131360 6640
rect 131140 6520 131150 6590
rect 131350 6520 131360 6590
rect 131140 6480 131360 6520
rect 131140 6410 131150 6480
rect 131350 6410 131360 6480
rect 131140 6360 131360 6410
rect 131640 6590 131860 6640
rect 131640 6520 131650 6590
rect 131850 6520 131860 6590
rect 131640 6480 131860 6520
rect 131640 6410 131650 6480
rect 131850 6410 131860 6480
rect 131640 6360 131860 6410
rect 132140 6590 132360 6640
rect 132140 6520 132150 6590
rect 132350 6520 132360 6590
rect 132140 6480 132360 6520
rect 132140 6410 132150 6480
rect 132350 6410 132360 6480
rect 132140 6360 132360 6410
rect 132640 6590 132860 6640
rect 132640 6520 132650 6590
rect 132850 6520 132860 6590
rect 132640 6480 132860 6520
rect 132640 6410 132650 6480
rect 132850 6410 132860 6480
rect 132640 6360 132860 6410
rect 133140 6590 133360 6640
rect 133140 6520 133150 6590
rect 133350 6520 133360 6590
rect 133140 6480 133360 6520
rect 133140 6410 133150 6480
rect 133350 6410 133360 6480
rect 133140 6360 133360 6410
rect 133640 6590 133860 6640
rect 133640 6520 133650 6590
rect 133850 6520 133860 6590
rect 133640 6480 133860 6520
rect 133640 6410 133650 6480
rect 133850 6410 133860 6480
rect 133640 6360 133860 6410
rect 134140 6590 134360 6640
rect 134140 6520 134150 6590
rect 134350 6520 134360 6590
rect 134140 6480 134360 6520
rect 134140 6410 134150 6480
rect 134350 6410 134360 6480
rect 134140 6360 134360 6410
rect 134640 6590 134860 6640
rect 134640 6520 134650 6590
rect 134850 6520 134860 6590
rect 134640 6480 134860 6520
rect 134640 6410 134650 6480
rect 134850 6410 134860 6480
rect 134640 6360 134860 6410
rect 135140 6590 135360 6640
rect 135140 6520 135150 6590
rect 135350 6520 135360 6590
rect 135140 6480 135360 6520
rect 135140 6410 135150 6480
rect 135350 6410 135360 6480
rect 135140 6360 135360 6410
rect 135640 6590 135860 6640
rect 135640 6520 135650 6590
rect 135850 6520 135860 6590
rect 135640 6480 135860 6520
rect 135640 6410 135650 6480
rect 135850 6410 135860 6480
rect 135640 6360 135860 6410
rect 136140 6590 136360 6640
rect 136140 6520 136150 6590
rect 136350 6520 136360 6590
rect 136140 6480 136360 6520
rect 136140 6410 136150 6480
rect 136350 6410 136360 6480
rect 136140 6360 136360 6410
rect 136640 6590 136860 6640
rect 136640 6520 136650 6590
rect 136850 6520 136860 6590
rect 136640 6480 136860 6520
rect 136640 6410 136650 6480
rect 136850 6410 136860 6480
rect 136640 6360 136860 6410
rect 137140 6590 137360 6640
rect 137140 6520 137150 6590
rect 137350 6520 137360 6590
rect 137140 6480 137360 6520
rect 137140 6410 137150 6480
rect 137350 6410 137360 6480
rect 137140 6360 137360 6410
rect 137640 6590 137860 6640
rect 137640 6520 137650 6590
rect 137850 6520 137860 6590
rect 137640 6480 137860 6520
rect 137640 6410 137650 6480
rect 137850 6410 137860 6480
rect 137640 6360 137860 6410
rect 138140 6590 138360 6640
rect 138140 6520 138150 6590
rect 138350 6520 138360 6590
rect 138140 6480 138360 6520
rect 138140 6410 138150 6480
rect 138350 6410 138360 6480
rect 138140 6360 138360 6410
rect 138640 6590 138860 6640
rect 138640 6520 138650 6590
rect 138850 6520 138860 6590
rect 138640 6480 138860 6520
rect 138640 6410 138650 6480
rect 138850 6410 138860 6480
rect 138640 6360 138860 6410
rect 139140 6590 139360 6640
rect 139140 6520 139150 6590
rect 139350 6520 139360 6590
rect 139140 6480 139360 6520
rect 139140 6410 139150 6480
rect 139350 6410 139360 6480
rect 139140 6360 139360 6410
rect 139640 6590 139860 6640
rect 139640 6520 139650 6590
rect 139850 6520 139860 6590
rect 139640 6480 139860 6520
rect 139640 6410 139650 6480
rect 139850 6410 139860 6480
rect 139640 6360 139860 6410
rect 128000 6350 140000 6360
rect 128000 6150 128020 6350
rect 128090 6150 128410 6350
rect 128480 6150 128520 6350
rect 128590 6150 128910 6350
rect 128980 6150 129020 6350
rect 129090 6150 129410 6350
rect 129480 6150 129520 6350
rect 129590 6150 129910 6350
rect 129980 6150 130020 6350
rect 130090 6150 130410 6350
rect 130480 6150 130520 6350
rect 130590 6150 130910 6350
rect 130980 6150 131020 6350
rect 131090 6150 131410 6350
rect 131480 6150 131520 6350
rect 131590 6150 131910 6350
rect 131980 6150 132020 6350
rect 132090 6150 132410 6350
rect 132480 6150 132520 6350
rect 132590 6150 132910 6350
rect 132980 6150 133020 6350
rect 133090 6150 133410 6350
rect 133480 6150 133520 6350
rect 133590 6150 133910 6350
rect 133980 6150 134020 6350
rect 134090 6150 134410 6350
rect 134480 6150 134520 6350
rect 134590 6150 134910 6350
rect 134980 6150 135020 6350
rect 135090 6150 135410 6350
rect 135480 6150 135520 6350
rect 135590 6150 135910 6350
rect 135980 6150 136020 6350
rect 136090 6150 136410 6350
rect 136480 6150 136520 6350
rect 136590 6150 136910 6350
rect 136980 6150 137020 6350
rect 137090 6150 137410 6350
rect 137480 6150 137520 6350
rect 137590 6150 137910 6350
rect 137980 6150 138020 6350
rect 138090 6150 138410 6350
rect 138480 6150 138520 6350
rect 138590 6150 138910 6350
rect 138980 6150 139020 6350
rect 139090 6150 139410 6350
rect 139480 6150 139520 6350
rect 139590 6150 139910 6350
rect 139980 6150 140000 6350
rect 128000 6140 140000 6150
rect 128140 6090 128360 6140
rect 128140 6020 128150 6090
rect 128350 6020 128360 6090
rect 128140 6000 128360 6020
rect 128640 6090 128860 6140
rect 128640 6020 128650 6090
rect 128850 6020 128860 6090
rect 128640 6000 128860 6020
rect 129140 6090 129360 6140
rect 129140 6020 129150 6090
rect 129350 6020 129360 6090
rect 129140 6000 129360 6020
rect 129640 6090 129860 6140
rect 129640 6020 129650 6090
rect 129850 6020 129860 6090
rect 129640 6000 129860 6020
rect 130140 6090 130360 6140
rect 130140 6020 130150 6090
rect 130350 6020 130360 6090
rect 130140 6000 130360 6020
rect 130640 6090 130860 6140
rect 130640 6020 130650 6090
rect 130850 6020 130860 6090
rect 130640 6000 130860 6020
rect 131140 6090 131360 6140
rect 131140 6020 131150 6090
rect 131350 6020 131360 6090
rect 131140 6000 131360 6020
rect 131640 6090 131860 6140
rect 131640 6020 131650 6090
rect 131850 6020 131860 6090
rect 131640 6000 131860 6020
rect 132140 6090 132360 6140
rect 132140 6020 132150 6090
rect 132350 6020 132360 6090
rect 132140 6000 132360 6020
rect 132640 6090 132860 6140
rect 132640 6020 132650 6090
rect 132850 6020 132860 6090
rect 132640 6000 132860 6020
rect 133140 6090 133360 6140
rect 133140 6020 133150 6090
rect 133350 6020 133360 6090
rect 133140 6000 133360 6020
rect 133640 6090 133860 6140
rect 133640 6020 133650 6090
rect 133850 6020 133860 6090
rect 133640 6000 133860 6020
rect 134140 6090 134360 6140
rect 134140 6020 134150 6090
rect 134350 6020 134360 6090
rect 134140 6000 134360 6020
rect 134640 6090 134860 6140
rect 134640 6020 134650 6090
rect 134850 6020 134860 6090
rect 134640 6000 134860 6020
rect 135140 6090 135360 6140
rect 135140 6020 135150 6090
rect 135350 6020 135360 6090
rect 135140 6000 135360 6020
rect 135640 6090 135860 6140
rect 135640 6020 135650 6090
rect 135850 6020 135860 6090
rect 135640 6000 135860 6020
rect 136140 6090 136360 6140
rect 136140 6020 136150 6090
rect 136350 6020 136360 6090
rect 136140 5980 136360 6020
rect 136140 5910 136150 5980
rect 136350 5910 136360 5980
rect 136140 5860 136360 5910
rect 136640 6090 136860 6140
rect 136640 6020 136650 6090
rect 136850 6020 136860 6090
rect 136640 5980 136860 6020
rect 136640 5910 136650 5980
rect 136850 5910 136860 5980
rect 136640 5860 136860 5910
rect 137140 6090 137360 6140
rect 137140 6020 137150 6090
rect 137350 6020 137360 6090
rect 137140 5980 137360 6020
rect 137140 5910 137150 5980
rect 137350 5910 137360 5980
rect 137140 5860 137360 5910
rect 137640 6090 137860 6140
rect 137640 6020 137650 6090
rect 137850 6020 137860 6090
rect 137640 5980 137860 6020
rect 137640 5910 137650 5980
rect 137850 5910 137860 5980
rect 137640 5860 137860 5910
rect 138140 6090 138360 6140
rect 138140 6020 138150 6090
rect 138350 6020 138360 6090
rect 138140 5980 138360 6020
rect 138140 5910 138150 5980
rect 138350 5910 138360 5980
rect 138140 5860 138360 5910
rect 138640 6090 138860 6140
rect 138640 6020 138650 6090
rect 138850 6020 138860 6090
rect 138640 5980 138860 6020
rect 138640 5910 138650 5980
rect 138850 5910 138860 5980
rect 138640 5860 138860 5910
rect 139140 6090 139360 6140
rect 139140 6020 139150 6090
rect 139350 6020 139360 6090
rect 139140 5980 139360 6020
rect 139140 5910 139150 5980
rect 139350 5910 139360 5980
rect 139140 5860 139360 5910
rect 139640 6090 139860 6140
rect 139640 6020 139650 6090
rect 139850 6020 139860 6090
rect 139640 5980 139860 6020
rect 139640 5910 139650 5980
rect 139850 5910 139860 5980
rect 139640 5860 139860 5910
rect 136000 5850 140000 5860
rect 136000 5650 136020 5850
rect 136090 5650 136410 5850
rect 136480 5650 136520 5850
rect 136590 5650 136910 5850
rect 136980 5650 137020 5850
rect 137090 5650 137410 5850
rect 137480 5650 137520 5850
rect 137590 5650 137910 5850
rect 137980 5650 138020 5850
rect 138090 5650 138410 5850
rect 138480 5650 138520 5850
rect 138590 5650 138910 5850
rect 138980 5650 139020 5850
rect 139090 5650 139410 5850
rect 139480 5650 139520 5850
rect 139590 5650 139910 5850
rect 139980 5650 140000 5850
rect 136000 5640 140000 5650
rect 136140 5590 136360 5640
rect 136140 5520 136150 5590
rect 136350 5520 136360 5590
rect 136140 5480 136360 5520
rect 136140 5410 136150 5480
rect 136350 5410 136360 5480
rect 136140 5360 136360 5410
rect 136640 5590 136860 5640
rect 136640 5520 136650 5590
rect 136850 5520 136860 5590
rect 136640 5480 136860 5520
rect 136640 5410 136650 5480
rect 136850 5410 136860 5480
rect 136640 5360 136860 5410
rect 137140 5590 137360 5640
rect 137140 5520 137150 5590
rect 137350 5520 137360 5590
rect 137140 5480 137360 5520
rect 137140 5410 137150 5480
rect 137350 5410 137360 5480
rect 137140 5360 137360 5410
rect 137640 5590 137860 5640
rect 137640 5520 137650 5590
rect 137850 5520 137860 5590
rect 137640 5480 137860 5520
rect 137640 5410 137650 5480
rect 137850 5410 137860 5480
rect 137640 5360 137860 5410
rect 138140 5590 138360 5640
rect 138140 5520 138150 5590
rect 138350 5520 138360 5590
rect 138140 5480 138360 5520
rect 138140 5410 138150 5480
rect 138350 5410 138360 5480
rect 138140 5360 138360 5410
rect 138640 5590 138860 5640
rect 138640 5520 138650 5590
rect 138850 5520 138860 5590
rect 138640 5480 138860 5520
rect 138640 5410 138650 5480
rect 138850 5410 138860 5480
rect 138640 5360 138860 5410
rect 139140 5590 139360 5640
rect 139140 5520 139150 5590
rect 139350 5520 139360 5590
rect 139140 5480 139360 5520
rect 139140 5410 139150 5480
rect 139350 5410 139360 5480
rect 139140 5360 139360 5410
rect 139640 5590 139860 5640
rect 139640 5520 139650 5590
rect 139850 5520 139860 5590
rect 139640 5480 139860 5520
rect 139640 5410 139650 5480
rect 139850 5410 139860 5480
rect 139640 5360 139860 5410
rect 136000 5350 140000 5360
rect 136000 5150 136020 5350
rect 136090 5150 136410 5350
rect 136480 5150 136520 5350
rect 136590 5150 136910 5350
rect 136980 5150 137020 5350
rect 137090 5150 137410 5350
rect 137480 5150 137520 5350
rect 137590 5150 137910 5350
rect 137980 5150 138020 5350
rect 138090 5150 138410 5350
rect 138480 5150 138520 5350
rect 138590 5150 138910 5350
rect 138980 5150 139020 5350
rect 139090 5150 139410 5350
rect 139480 5150 139520 5350
rect 139590 5150 139910 5350
rect 139980 5150 140000 5350
rect 136000 5140 140000 5150
rect 136140 5090 136360 5140
rect 136140 5020 136150 5090
rect 136350 5020 136360 5090
rect 136140 4980 136360 5020
rect 136140 4910 136150 4980
rect 136350 4910 136360 4980
rect 136140 4860 136360 4910
rect 136640 5090 136860 5140
rect 136640 5020 136650 5090
rect 136850 5020 136860 5090
rect 136640 4980 136860 5020
rect 136640 4910 136650 4980
rect 136850 4910 136860 4980
rect 136640 4860 136860 4910
rect 137140 5090 137360 5140
rect 137140 5020 137150 5090
rect 137350 5020 137360 5090
rect 137140 4980 137360 5020
rect 137140 4910 137150 4980
rect 137350 4910 137360 4980
rect 137140 4860 137360 4910
rect 137640 5090 137860 5140
rect 137640 5020 137650 5090
rect 137850 5020 137860 5090
rect 137640 4980 137860 5020
rect 137640 4910 137650 4980
rect 137850 4910 137860 4980
rect 137640 4860 137860 4910
rect 138140 5090 138360 5140
rect 138140 5020 138150 5090
rect 138350 5020 138360 5090
rect 138140 4980 138360 5020
rect 138140 4910 138150 4980
rect 138350 4910 138360 4980
rect 138140 4860 138360 4910
rect 138640 5090 138860 5140
rect 138640 5020 138650 5090
rect 138850 5020 138860 5090
rect 138640 4980 138860 5020
rect 138640 4910 138650 4980
rect 138850 4910 138860 4980
rect 138640 4860 138860 4910
rect 139140 5090 139360 5140
rect 139140 5020 139150 5090
rect 139350 5020 139360 5090
rect 139140 4980 139360 5020
rect 139140 4910 139150 4980
rect 139350 4910 139360 4980
rect 139140 4860 139360 4910
rect 139640 5090 139860 5140
rect 139640 5020 139650 5090
rect 139850 5020 139860 5090
rect 139640 4980 139860 5020
rect 139640 4910 139650 4980
rect 139850 4910 139860 4980
rect 139640 4860 139860 4910
rect 136000 4850 140000 4860
rect 136000 4650 136020 4850
rect 136090 4650 136410 4850
rect 136480 4650 136520 4850
rect 136590 4650 136910 4850
rect 136980 4650 137020 4850
rect 137090 4650 137410 4850
rect 137480 4650 137520 4850
rect 137590 4650 137910 4850
rect 137980 4650 138020 4850
rect 138090 4650 138410 4850
rect 138480 4650 138520 4850
rect 138590 4650 138910 4850
rect 138980 4650 139020 4850
rect 139090 4650 139410 4850
rect 139480 4650 139520 4850
rect 139590 4650 139910 4850
rect 139980 4650 140000 4850
rect 136000 4640 140000 4650
rect 136140 4590 136360 4640
rect 136140 4520 136150 4590
rect 136350 4520 136360 4590
rect 136140 4480 136360 4520
rect 136140 4410 136150 4480
rect 136350 4410 136360 4480
rect 136140 4360 136360 4410
rect 136640 4590 136860 4640
rect 136640 4520 136650 4590
rect 136850 4520 136860 4590
rect 136640 4480 136860 4520
rect 136640 4410 136650 4480
rect 136850 4410 136860 4480
rect 136640 4360 136860 4410
rect 137140 4590 137360 4640
rect 137140 4520 137150 4590
rect 137350 4520 137360 4590
rect 137140 4480 137360 4520
rect 137140 4410 137150 4480
rect 137350 4410 137360 4480
rect 137140 4360 137360 4410
rect 137640 4590 137860 4640
rect 137640 4520 137650 4590
rect 137850 4520 137860 4590
rect 137640 4480 137860 4520
rect 137640 4410 137650 4480
rect 137850 4410 137860 4480
rect 137640 4360 137860 4410
rect 138140 4590 138360 4640
rect 138140 4520 138150 4590
rect 138350 4520 138360 4590
rect 138140 4480 138360 4520
rect 138140 4410 138150 4480
rect 138350 4410 138360 4480
rect 138140 4360 138360 4410
rect 138640 4590 138860 4640
rect 138640 4520 138650 4590
rect 138850 4520 138860 4590
rect 138640 4480 138860 4520
rect 138640 4410 138650 4480
rect 138850 4410 138860 4480
rect 138640 4360 138860 4410
rect 139140 4590 139360 4640
rect 139140 4520 139150 4590
rect 139350 4520 139360 4590
rect 139140 4480 139360 4520
rect 139140 4410 139150 4480
rect 139350 4410 139360 4480
rect 139140 4360 139360 4410
rect 139640 4590 139860 4640
rect 139640 4520 139650 4590
rect 139850 4520 139860 4590
rect 139640 4480 139860 4520
rect 139640 4410 139650 4480
rect 139850 4410 139860 4480
rect 139640 4360 139860 4410
rect 136000 4350 140000 4360
rect 136000 4150 136020 4350
rect 136090 4150 136410 4350
rect 136480 4150 136520 4350
rect 136590 4150 136910 4350
rect 136980 4150 137020 4350
rect 137090 4150 137410 4350
rect 137480 4150 137520 4350
rect 137590 4150 137910 4350
rect 137980 4150 138020 4350
rect 138090 4150 138410 4350
rect 138480 4150 138520 4350
rect 138590 4150 138910 4350
rect 138980 4150 139020 4350
rect 139090 4150 139410 4350
rect 139480 4150 139520 4350
rect 139590 4150 139910 4350
rect 139980 4150 140000 4350
rect 136000 4140 140000 4150
rect 136140 4090 136360 4140
rect 136140 4020 136150 4090
rect 136350 4020 136360 4090
rect 136140 3980 136360 4020
rect 136140 3910 136150 3980
rect 136350 3910 136360 3980
rect 136140 3860 136360 3910
rect 136640 4090 136860 4140
rect 136640 4020 136650 4090
rect 136850 4020 136860 4090
rect 136640 3980 136860 4020
rect 136640 3910 136650 3980
rect 136850 3910 136860 3980
rect 136640 3860 136860 3910
rect 137140 4090 137360 4140
rect 137140 4020 137150 4090
rect 137350 4020 137360 4090
rect 137140 3980 137360 4020
rect 137140 3910 137150 3980
rect 137350 3910 137360 3980
rect 137140 3860 137360 3910
rect 137640 4090 137860 4140
rect 137640 4020 137650 4090
rect 137850 4020 137860 4090
rect 137640 3980 137860 4020
rect 137640 3910 137650 3980
rect 137850 3910 137860 3980
rect 137640 3860 137860 3910
rect 138140 4090 138360 4140
rect 138140 4020 138150 4090
rect 138350 4020 138360 4090
rect 138140 3980 138360 4020
rect 138140 3910 138150 3980
rect 138350 3910 138360 3980
rect 138140 3860 138360 3910
rect 138640 4090 138860 4140
rect 138640 4020 138650 4090
rect 138850 4020 138860 4090
rect 138640 3980 138860 4020
rect 138640 3910 138650 3980
rect 138850 3910 138860 3980
rect 138640 3860 138860 3910
rect 139140 4090 139360 4140
rect 139140 4020 139150 4090
rect 139350 4020 139360 4090
rect 139140 3980 139360 4020
rect 139140 3910 139150 3980
rect 139350 3910 139360 3980
rect 139140 3860 139360 3910
rect 139640 4090 139860 4140
rect 139640 4020 139650 4090
rect 139850 4020 139860 4090
rect 139640 3980 139860 4020
rect 139640 3910 139650 3980
rect 139850 3910 139860 3980
rect 139640 3860 139860 3910
rect 136000 3850 140000 3860
rect 136000 3650 136020 3850
rect 136090 3650 136410 3850
rect 136480 3650 136520 3850
rect 136590 3650 136910 3850
rect 136980 3650 137020 3850
rect 137090 3650 137410 3850
rect 137480 3650 137520 3850
rect 137590 3650 137910 3850
rect 137980 3650 138020 3850
rect 138090 3650 138410 3850
rect 138480 3650 138520 3850
rect 138590 3650 138910 3850
rect 138980 3650 139020 3850
rect 139090 3650 139410 3850
rect 139480 3650 139520 3850
rect 139590 3650 139910 3850
rect 139980 3650 140000 3850
rect 136000 3640 140000 3650
rect 136140 3590 136360 3640
rect 136140 3520 136150 3590
rect 136350 3520 136360 3590
rect 136140 3480 136360 3520
rect 136140 3410 136150 3480
rect 136350 3410 136360 3480
rect 136140 3360 136360 3410
rect 136640 3590 136860 3640
rect 136640 3520 136650 3590
rect 136850 3520 136860 3590
rect 136640 3480 136860 3520
rect 136640 3410 136650 3480
rect 136850 3410 136860 3480
rect 136640 3360 136860 3410
rect 137140 3590 137360 3640
rect 137140 3520 137150 3590
rect 137350 3520 137360 3590
rect 137140 3480 137360 3520
rect 137140 3410 137150 3480
rect 137350 3410 137360 3480
rect 137140 3360 137360 3410
rect 137640 3590 137860 3640
rect 137640 3520 137650 3590
rect 137850 3520 137860 3590
rect 137640 3480 137860 3520
rect 137640 3410 137650 3480
rect 137850 3410 137860 3480
rect 137640 3360 137860 3410
rect 138140 3590 138360 3640
rect 138140 3520 138150 3590
rect 138350 3520 138360 3590
rect 138140 3480 138360 3520
rect 138140 3410 138150 3480
rect 138350 3410 138360 3480
rect 138140 3360 138360 3410
rect 138640 3590 138860 3640
rect 138640 3520 138650 3590
rect 138850 3520 138860 3590
rect 138640 3480 138860 3520
rect 138640 3410 138650 3480
rect 138850 3410 138860 3480
rect 138640 3360 138860 3410
rect 139140 3590 139360 3640
rect 139140 3520 139150 3590
rect 139350 3520 139360 3590
rect 139140 3480 139360 3520
rect 139140 3410 139150 3480
rect 139350 3410 139360 3480
rect 139140 3360 139360 3410
rect 139640 3590 139860 3640
rect 139640 3520 139650 3590
rect 139850 3520 139860 3590
rect 139640 3480 139860 3520
rect 139640 3410 139650 3480
rect 139850 3410 139860 3480
rect 139640 3360 139860 3410
rect 136000 3350 140000 3360
rect 136000 3150 136020 3350
rect 136090 3150 136410 3350
rect 136480 3150 136520 3350
rect 136590 3150 136910 3350
rect 136980 3150 137020 3350
rect 137090 3150 137410 3350
rect 137480 3150 137520 3350
rect 137590 3150 137910 3350
rect 137980 3150 138020 3350
rect 138090 3150 138410 3350
rect 138480 3150 138520 3350
rect 138590 3150 138910 3350
rect 138980 3150 139020 3350
rect 139090 3150 139410 3350
rect 139480 3150 139520 3350
rect 139590 3150 139910 3350
rect 139980 3150 140000 3350
rect 136000 3140 140000 3150
rect 136140 3090 136360 3140
rect 136140 3020 136150 3090
rect 136350 3020 136360 3090
rect 136140 2980 136360 3020
rect 136140 2910 136150 2980
rect 136350 2910 136360 2980
rect 136140 2860 136360 2910
rect 136640 3090 136860 3140
rect 136640 3020 136650 3090
rect 136850 3020 136860 3090
rect 136640 2980 136860 3020
rect 136640 2910 136650 2980
rect 136850 2910 136860 2980
rect 136640 2860 136860 2910
rect 137140 3090 137360 3140
rect 137140 3020 137150 3090
rect 137350 3020 137360 3090
rect 137140 2980 137360 3020
rect 137140 2910 137150 2980
rect 137350 2910 137360 2980
rect 137140 2860 137360 2910
rect 137640 3090 137860 3140
rect 137640 3020 137650 3090
rect 137850 3020 137860 3090
rect 137640 2980 137860 3020
rect 137640 2910 137650 2980
rect 137850 2910 137860 2980
rect 137640 2860 137860 2910
rect 138140 3090 138360 3140
rect 138140 3020 138150 3090
rect 138350 3020 138360 3090
rect 138140 2980 138360 3020
rect 138140 2910 138150 2980
rect 138350 2910 138360 2980
rect 138140 2860 138360 2910
rect 138640 3090 138860 3140
rect 138640 3020 138650 3090
rect 138850 3020 138860 3090
rect 138640 2980 138860 3020
rect 138640 2910 138650 2980
rect 138850 2910 138860 2980
rect 138640 2860 138860 2910
rect 139140 3090 139360 3140
rect 139140 3020 139150 3090
rect 139350 3020 139360 3090
rect 139140 2980 139360 3020
rect 139140 2910 139150 2980
rect 139350 2910 139360 2980
rect 139140 2860 139360 2910
rect 139640 3090 139860 3140
rect 139640 3020 139650 3090
rect 139850 3020 139860 3090
rect 139640 2980 139860 3020
rect 139640 2910 139650 2980
rect 139850 2910 139860 2980
rect 139640 2860 139860 2910
rect 136000 2850 140000 2860
rect 136000 2650 136020 2850
rect 136090 2650 136410 2850
rect 136480 2650 136520 2850
rect 136590 2650 136910 2850
rect 136980 2650 137020 2850
rect 137090 2650 137410 2850
rect 137480 2650 137520 2850
rect 137590 2650 137910 2850
rect 137980 2650 138020 2850
rect 138090 2650 138410 2850
rect 138480 2650 138520 2850
rect 138590 2650 138910 2850
rect 138980 2650 139020 2850
rect 139090 2650 139410 2850
rect 139480 2650 139520 2850
rect 139590 2650 139910 2850
rect 139980 2650 140000 2850
rect 136000 2640 140000 2650
rect 136140 2590 136360 2640
rect 136140 2520 136150 2590
rect 136350 2520 136360 2590
rect 136140 2480 136360 2520
rect 136140 2410 136150 2480
rect 136350 2410 136360 2480
rect 136140 2360 136360 2410
rect 136640 2590 136860 2640
rect 136640 2520 136650 2590
rect 136850 2520 136860 2590
rect 136640 2480 136860 2520
rect 136640 2410 136650 2480
rect 136850 2410 136860 2480
rect 136640 2360 136860 2410
rect 137140 2590 137360 2640
rect 137140 2520 137150 2590
rect 137350 2520 137360 2590
rect 137140 2480 137360 2520
rect 137140 2410 137150 2480
rect 137350 2410 137360 2480
rect 137140 2360 137360 2410
rect 137640 2590 137860 2640
rect 137640 2520 137650 2590
rect 137850 2520 137860 2590
rect 137640 2480 137860 2520
rect 137640 2410 137650 2480
rect 137850 2410 137860 2480
rect 137640 2360 137860 2410
rect 138140 2590 138360 2640
rect 138140 2520 138150 2590
rect 138350 2520 138360 2590
rect 138140 2480 138360 2520
rect 138140 2410 138150 2480
rect 138350 2410 138360 2480
rect 138140 2360 138360 2410
rect 138640 2590 138860 2640
rect 138640 2520 138650 2590
rect 138850 2520 138860 2590
rect 138640 2480 138860 2520
rect 138640 2410 138650 2480
rect 138850 2410 138860 2480
rect 138640 2360 138860 2410
rect 139140 2590 139360 2640
rect 139140 2520 139150 2590
rect 139350 2520 139360 2590
rect 139140 2480 139360 2520
rect 139140 2410 139150 2480
rect 139350 2410 139360 2480
rect 139140 2360 139360 2410
rect 139640 2590 139860 2640
rect 139640 2520 139650 2590
rect 139850 2520 139860 2590
rect 139640 2480 139860 2520
rect 139640 2410 139650 2480
rect 139850 2410 139860 2480
rect 139640 2360 139860 2410
rect 136000 2350 140000 2360
rect 136000 2150 136020 2350
rect 136090 2150 136410 2350
rect 136480 2150 136520 2350
rect 136590 2150 136910 2350
rect 136980 2150 137020 2350
rect 137090 2150 137410 2350
rect 137480 2150 137520 2350
rect 137590 2150 137910 2350
rect 137980 2150 138020 2350
rect 138090 2150 138410 2350
rect 138480 2150 138520 2350
rect 138590 2150 138910 2350
rect 138980 2150 139020 2350
rect 139090 2150 139410 2350
rect 139480 2150 139520 2350
rect 139590 2150 139910 2350
rect 139980 2150 140000 2350
rect 136000 2140 140000 2150
rect 136140 2090 136360 2140
rect 136140 2020 136150 2090
rect 136350 2020 136360 2090
rect 136140 1980 136360 2020
rect 136140 1910 136150 1980
rect 136350 1910 136360 1980
rect 136140 1860 136360 1910
rect 136640 2090 136860 2140
rect 136640 2020 136650 2090
rect 136850 2020 136860 2090
rect 136640 1980 136860 2020
rect 136640 1910 136650 1980
rect 136850 1910 136860 1980
rect 136640 1860 136860 1910
rect 137140 2090 137360 2140
rect 137140 2020 137150 2090
rect 137350 2020 137360 2090
rect 137140 1980 137360 2020
rect 137140 1910 137150 1980
rect 137350 1910 137360 1980
rect 137140 1860 137360 1910
rect 137640 2090 137860 2140
rect 137640 2020 137650 2090
rect 137850 2020 137860 2090
rect 137640 1980 137860 2020
rect 137640 1910 137650 1980
rect 137850 1910 137860 1980
rect 137640 1860 137860 1910
rect 138140 2090 138360 2140
rect 138140 2020 138150 2090
rect 138350 2020 138360 2090
rect 138140 1980 138360 2020
rect 138140 1910 138150 1980
rect 138350 1910 138360 1980
rect 138140 1860 138360 1910
rect 138640 2090 138860 2140
rect 138640 2020 138650 2090
rect 138850 2020 138860 2090
rect 138640 1980 138860 2020
rect 138640 1910 138650 1980
rect 138850 1910 138860 1980
rect 138640 1860 138860 1910
rect 139140 2090 139360 2140
rect 139140 2020 139150 2090
rect 139350 2020 139360 2090
rect 139140 1980 139360 2020
rect 139140 1910 139150 1980
rect 139350 1910 139360 1980
rect 139140 1860 139360 1910
rect 139640 2090 139860 2140
rect 139640 2020 139650 2090
rect 139850 2020 139860 2090
rect 139640 1980 139860 2020
rect 139640 1910 139650 1980
rect 139850 1910 139860 1980
rect 139640 1860 139860 1910
rect 136000 1850 140000 1860
rect 136000 1650 136020 1850
rect 136090 1650 136410 1850
rect 136480 1650 136520 1850
rect 136590 1650 136910 1850
rect 136980 1650 137020 1850
rect 137090 1650 137410 1850
rect 137480 1650 137520 1850
rect 137590 1650 137910 1850
rect 137980 1650 138020 1850
rect 138090 1650 138410 1850
rect 138480 1650 138520 1850
rect 138590 1650 138910 1850
rect 138980 1650 139020 1850
rect 139090 1650 139410 1850
rect 139480 1650 139520 1850
rect 139590 1650 139910 1850
rect 139980 1650 140000 1850
rect 136000 1640 140000 1650
rect 136140 1590 136360 1640
rect 136140 1520 136150 1590
rect 136350 1520 136360 1590
rect 136140 1480 136360 1520
rect 136140 1410 136150 1480
rect 136350 1410 136360 1480
rect 136140 1360 136360 1410
rect 136640 1590 136860 1640
rect 136640 1520 136650 1590
rect 136850 1520 136860 1590
rect 136640 1480 136860 1520
rect 136640 1410 136650 1480
rect 136850 1410 136860 1480
rect 136640 1360 136860 1410
rect 137140 1590 137360 1640
rect 137140 1520 137150 1590
rect 137350 1520 137360 1590
rect 137140 1480 137360 1520
rect 137140 1410 137150 1480
rect 137350 1410 137360 1480
rect 137140 1360 137360 1410
rect 137640 1590 137860 1640
rect 137640 1520 137650 1590
rect 137850 1520 137860 1590
rect 137640 1480 137860 1520
rect 137640 1410 137650 1480
rect 137850 1410 137860 1480
rect 137640 1360 137860 1410
rect 138140 1590 138360 1640
rect 138140 1520 138150 1590
rect 138350 1520 138360 1590
rect 138140 1480 138360 1520
rect 138140 1410 138150 1480
rect 138350 1410 138360 1480
rect 138140 1360 138360 1410
rect 138640 1590 138860 1640
rect 138640 1520 138650 1590
rect 138850 1520 138860 1590
rect 138640 1480 138860 1520
rect 138640 1410 138650 1480
rect 138850 1410 138860 1480
rect 138640 1360 138860 1410
rect 139140 1590 139360 1640
rect 139140 1520 139150 1590
rect 139350 1520 139360 1590
rect 139140 1480 139360 1520
rect 139140 1410 139150 1480
rect 139350 1410 139360 1480
rect 139140 1360 139360 1410
rect 139640 1590 139860 1640
rect 139640 1520 139650 1590
rect 139850 1520 139860 1590
rect 139640 1480 139860 1520
rect 139640 1410 139650 1480
rect 139850 1410 139860 1480
rect 139640 1360 139860 1410
rect 136000 1350 140000 1360
rect 136000 1150 136020 1350
rect 136090 1150 136410 1350
rect 136480 1150 136520 1350
rect 136590 1150 136910 1350
rect 136980 1150 137020 1350
rect 137090 1150 137410 1350
rect 137480 1150 137520 1350
rect 137590 1150 137910 1350
rect 137980 1150 138020 1350
rect 138090 1150 138410 1350
rect 138480 1150 138520 1350
rect 138590 1150 138910 1350
rect 138980 1150 139020 1350
rect 139090 1150 139410 1350
rect 139480 1150 139520 1350
rect 139590 1150 139910 1350
rect 139980 1150 140000 1350
rect 136000 1140 140000 1150
rect 136140 1090 136360 1140
rect 136140 1020 136150 1090
rect 136350 1020 136360 1090
rect 136140 980 136360 1020
rect 136140 910 136150 980
rect 136350 910 136360 980
rect 136140 860 136360 910
rect 136640 1090 136860 1140
rect 136640 1020 136650 1090
rect 136850 1020 136860 1090
rect 136640 980 136860 1020
rect 136640 910 136650 980
rect 136850 910 136860 980
rect 136640 860 136860 910
rect 137140 1090 137360 1140
rect 137140 1020 137150 1090
rect 137350 1020 137360 1090
rect 137140 980 137360 1020
rect 137140 910 137150 980
rect 137350 910 137360 980
rect 137140 860 137360 910
rect 137640 1090 137860 1140
rect 137640 1020 137650 1090
rect 137850 1020 137860 1090
rect 137640 980 137860 1020
rect 137640 910 137650 980
rect 137850 910 137860 980
rect 137640 860 137860 910
rect 138140 1090 138360 1140
rect 138140 1020 138150 1090
rect 138350 1020 138360 1090
rect 138140 980 138360 1020
rect 138140 910 138150 980
rect 138350 910 138360 980
rect 138140 860 138360 910
rect 138640 1090 138860 1140
rect 138640 1020 138650 1090
rect 138850 1020 138860 1090
rect 138640 980 138860 1020
rect 138640 910 138650 980
rect 138850 910 138860 980
rect 138640 860 138860 910
rect 139140 1090 139360 1140
rect 139140 1020 139150 1090
rect 139350 1020 139360 1090
rect 139140 980 139360 1020
rect 139140 910 139150 980
rect 139350 910 139360 980
rect 139140 860 139360 910
rect 139640 1090 139860 1140
rect 139640 1020 139650 1090
rect 139850 1020 139860 1090
rect 139640 980 139860 1020
rect 139640 910 139650 980
rect 139850 910 139860 980
rect 139640 860 139860 910
rect 136000 850 140000 860
rect 136000 650 136020 850
rect 136090 650 136410 850
rect 136480 650 136520 850
rect 136590 650 136910 850
rect 136980 650 137020 850
rect 137090 650 137410 850
rect 137480 650 137520 850
rect 137590 650 137910 850
rect 137980 650 138020 850
rect 138090 650 138410 850
rect 138480 650 138520 850
rect 138590 650 138910 850
rect 138980 650 139020 850
rect 139090 650 139410 850
rect 139480 650 139520 850
rect 139590 650 139910 850
rect 139980 650 140000 850
rect 136000 640 140000 650
rect 136140 590 136360 640
rect 136140 520 136150 590
rect 136350 520 136360 590
rect 136140 480 136360 520
rect 136140 410 136150 480
rect 136350 410 136360 480
rect 136140 360 136360 410
rect 136640 590 136860 640
rect 136640 520 136650 590
rect 136850 520 136860 590
rect 136640 480 136860 520
rect 136640 410 136650 480
rect 136850 410 136860 480
rect 136640 360 136860 410
rect 137140 590 137360 640
rect 137140 520 137150 590
rect 137350 520 137360 590
rect 137140 480 137360 520
rect 137140 410 137150 480
rect 137350 410 137360 480
rect 137140 360 137360 410
rect 137640 590 137860 640
rect 137640 520 137650 590
rect 137850 520 137860 590
rect 137640 480 137860 520
rect 137640 410 137650 480
rect 137850 410 137860 480
rect 137640 360 137860 410
rect 138140 590 138360 640
rect 138140 520 138150 590
rect 138350 520 138360 590
rect 138140 480 138360 520
rect 138140 410 138150 480
rect 138350 410 138360 480
rect 138140 360 138360 410
rect 138640 590 138860 640
rect 138640 520 138650 590
rect 138850 520 138860 590
rect 138640 480 138860 520
rect 138640 410 138650 480
rect 138850 410 138860 480
rect 138640 360 138860 410
rect 139140 590 139360 640
rect 139140 520 139150 590
rect 139350 520 139360 590
rect 139140 480 139360 520
rect 139140 410 139150 480
rect 139350 410 139360 480
rect 139140 360 139360 410
rect 139640 590 139860 640
rect 139640 520 139650 590
rect 139850 520 139860 590
rect 139640 480 139860 520
rect 139640 410 139650 480
rect 139850 410 139860 480
rect 139640 360 139860 410
rect 136000 350 140000 360
rect 136000 150 136020 350
rect 136090 150 136410 350
rect 136480 150 136520 350
rect 136590 150 136910 350
rect 136980 150 137020 350
rect 137090 150 137410 350
rect 137480 150 137520 350
rect 137590 150 137910 350
rect 137980 150 138020 350
rect 138090 150 138410 350
rect 138480 150 138520 350
rect 138590 150 138910 350
rect 138980 150 139020 350
rect 139090 150 139410 350
rect 139480 150 139520 350
rect 139590 150 139910 350
rect 139980 150 140000 350
rect 136000 140 140000 150
rect 136140 90 136360 140
rect 136140 20 136150 90
rect 136350 20 136360 90
rect 136140 -20 136360 20
rect 136140 -90 136150 -20
rect 136350 -90 136360 -20
rect 136140 -140 136360 -90
rect 136640 90 136860 140
rect 136640 20 136650 90
rect 136850 20 136860 90
rect 136640 -20 136860 20
rect 136640 -90 136650 -20
rect 136850 -90 136860 -20
rect 136640 -140 136860 -90
rect 137140 90 137360 140
rect 137140 20 137150 90
rect 137350 20 137360 90
rect 137140 -20 137360 20
rect 137140 -90 137150 -20
rect 137350 -90 137360 -20
rect 137140 -140 137360 -90
rect 137640 90 137860 140
rect 137640 20 137650 90
rect 137850 20 137860 90
rect 137640 -20 137860 20
rect 137640 -90 137650 -20
rect 137850 -90 137860 -20
rect 137640 -140 137860 -90
rect 138140 90 138360 140
rect 138140 20 138150 90
rect 138350 20 138360 90
rect 138140 -20 138360 20
rect 138140 -90 138150 -20
rect 138350 -90 138360 -20
rect 138140 -140 138360 -90
rect 138640 90 138860 140
rect 138640 20 138650 90
rect 138850 20 138860 90
rect 138640 -20 138860 20
rect 138640 -90 138650 -20
rect 138850 -90 138860 -20
rect 138640 -140 138860 -90
rect 139140 90 139360 140
rect 139140 20 139150 90
rect 139350 20 139360 90
rect 139140 -20 139360 20
rect 139140 -90 139150 -20
rect 139350 -90 139360 -20
rect 139140 -140 139360 -90
rect 139640 90 139860 140
rect 139640 20 139650 90
rect 139850 20 139860 90
rect 139640 -20 139860 20
rect 139640 -90 139650 -20
rect 139850 -90 139860 -20
rect 139640 -140 139860 -90
rect 136000 -150 140000 -140
rect 136000 -350 136020 -150
rect 136090 -350 136410 -150
rect 136480 -350 136520 -150
rect 136590 -350 136910 -150
rect 136980 -350 137020 -150
rect 137090 -350 137410 -150
rect 137480 -350 137520 -150
rect 137590 -350 137910 -150
rect 137980 -350 138020 -150
rect 138090 -350 138410 -150
rect 138480 -350 138520 -150
rect 138590 -350 138910 -150
rect 138980 -350 139020 -150
rect 139090 -350 139410 -150
rect 139480 -350 139520 -150
rect 139590 -350 139910 -150
rect 139980 -350 140000 -150
rect 136000 -360 140000 -350
rect 136140 -410 136360 -360
rect 136140 -480 136150 -410
rect 136350 -480 136360 -410
rect 136140 -520 136360 -480
rect 136140 -590 136150 -520
rect 136350 -590 136360 -520
rect 136140 -640 136360 -590
rect 136640 -410 136860 -360
rect 136640 -480 136650 -410
rect 136850 -480 136860 -410
rect 136640 -520 136860 -480
rect 136640 -590 136650 -520
rect 136850 -590 136860 -520
rect 136640 -640 136860 -590
rect 137140 -410 137360 -360
rect 137140 -480 137150 -410
rect 137350 -480 137360 -410
rect 137140 -520 137360 -480
rect 137140 -590 137150 -520
rect 137350 -590 137360 -520
rect 137140 -640 137360 -590
rect 137640 -410 137860 -360
rect 137640 -480 137650 -410
rect 137850 -480 137860 -410
rect 137640 -520 137860 -480
rect 137640 -590 137650 -520
rect 137850 -590 137860 -520
rect 137640 -640 137860 -590
rect 138140 -410 138360 -360
rect 138140 -480 138150 -410
rect 138350 -480 138360 -410
rect 138140 -520 138360 -480
rect 138140 -590 138150 -520
rect 138350 -590 138360 -520
rect 138140 -640 138360 -590
rect 138640 -410 138860 -360
rect 138640 -480 138650 -410
rect 138850 -480 138860 -410
rect 138640 -520 138860 -480
rect 138640 -590 138650 -520
rect 138850 -590 138860 -520
rect 138640 -640 138860 -590
rect 139140 -410 139360 -360
rect 139140 -480 139150 -410
rect 139350 -480 139360 -410
rect 139140 -520 139360 -480
rect 139140 -590 139150 -520
rect 139350 -590 139360 -520
rect 139140 -640 139360 -590
rect 139640 -410 139860 -360
rect 139640 -480 139650 -410
rect 139850 -480 139860 -410
rect 139640 -520 139860 -480
rect 139640 -590 139650 -520
rect 139850 -590 139860 -520
rect 139640 -640 139860 -590
rect 136000 -650 140000 -640
rect 136000 -850 136020 -650
rect 136090 -850 136410 -650
rect 136480 -850 136520 -650
rect 136590 -850 136910 -650
rect 136980 -850 137020 -650
rect 137090 -850 137410 -650
rect 137480 -850 137520 -650
rect 137590 -850 137910 -650
rect 137980 -850 138020 -650
rect 138090 -850 138410 -650
rect 138480 -850 138520 -650
rect 138590 -850 138910 -650
rect 138980 -850 139020 -650
rect 139090 -850 139410 -650
rect 139480 -850 139520 -650
rect 139590 -850 139910 -650
rect 139980 -850 140000 -650
rect 136000 -860 140000 -850
rect 136140 -910 136360 -860
rect 136140 -980 136150 -910
rect 136350 -980 136360 -910
rect 136140 -1020 136360 -980
rect 136140 -1090 136150 -1020
rect 136350 -1090 136360 -1020
rect 136140 -1140 136360 -1090
rect 136640 -910 136860 -860
rect 136640 -980 136650 -910
rect 136850 -980 136860 -910
rect 136640 -1020 136860 -980
rect 136640 -1090 136650 -1020
rect 136850 -1090 136860 -1020
rect 136640 -1140 136860 -1090
rect 137140 -910 137360 -860
rect 137140 -980 137150 -910
rect 137350 -980 137360 -910
rect 137140 -1020 137360 -980
rect 137140 -1090 137150 -1020
rect 137350 -1090 137360 -1020
rect 137140 -1140 137360 -1090
rect 137640 -910 137860 -860
rect 137640 -980 137650 -910
rect 137850 -980 137860 -910
rect 137640 -1020 137860 -980
rect 137640 -1090 137650 -1020
rect 137850 -1090 137860 -1020
rect 137640 -1140 137860 -1090
rect 138140 -910 138360 -860
rect 138140 -980 138150 -910
rect 138350 -980 138360 -910
rect 138140 -1020 138360 -980
rect 138140 -1090 138150 -1020
rect 138350 -1090 138360 -1020
rect 138140 -1140 138360 -1090
rect 138640 -910 138860 -860
rect 138640 -980 138650 -910
rect 138850 -980 138860 -910
rect 138640 -1020 138860 -980
rect 138640 -1090 138650 -1020
rect 138850 -1090 138860 -1020
rect 138640 -1140 138860 -1090
rect 139140 -910 139360 -860
rect 139140 -980 139150 -910
rect 139350 -980 139360 -910
rect 139140 -1020 139360 -980
rect 139140 -1090 139150 -1020
rect 139350 -1090 139360 -1020
rect 139140 -1140 139360 -1090
rect 139640 -910 139860 -860
rect 139640 -980 139650 -910
rect 139850 -980 139860 -910
rect 139640 -1020 139860 -980
rect 139640 -1090 139650 -1020
rect 139850 -1090 139860 -1020
rect 139640 -1140 139860 -1090
rect 136000 -1150 140000 -1140
rect 136000 -1350 136020 -1150
rect 136090 -1350 136410 -1150
rect 136480 -1350 136520 -1150
rect 136590 -1350 136910 -1150
rect 136980 -1350 137020 -1150
rect 137090 -1350 137410 -1150
rect 137480 -1350 137520 -1150
rect 137590 -1350 137910 -1150
rect 137980 -1350 138020 -1150
rect 138090 -1350 138410 -1150
rect 138480 -1350 138520 -1150
rect 138590 -1350 138910 -1150
rect 138980 -1350 139020 -1150
rect 139090 -1350 139410 -1150
rect 139480 -1350 139520 -1150
rect 139590 -1350 139910 -1150
rect 139980 -1350 140000 -1150
rect 136000 -1360 140000 -1350
rect 136140 -1410 136360 -1360
rect 136140 -1480 136150 -1410
rect 136350 -1480 136360 -1410
rect 136140 -1520 136360 -1480
rect 136140 -1590 136150 -1520
rect 136350 -1590 136360 -1520
rect 136140 -1640 136360 -1590
rect 136640 -1410 136860 -1360
rect 136640 -1480 136650 -1410
rect 136850 -1480 136860 -1410
rect 136640 -1520 136860 -1480
rect 136640 -1590 136650 -1520
rect 136850 -1590 136860 -1520
rect 136640 -1640 136860 -1590
rect 137140 -1410 137360 -1360
rect 137140 -1480 137150 -1410
rect 137350 -1480 137360 -1410
rect 137140 -1520 137360 -1480
rect 137140 -1590 137150 -1520
rect 137350 -1590 137360 -1520
rect 137140 -1640 137360 -1590
rect 137640 -1410 137860 -1360
rect 137640 -1480 137650 -1410
rect 137850 -1480 137860 -1410
rect 137640 -1520 137860 -1480
rect 137640 -1590 137650 -1520
rect 137850 -1590 137860 -1520
rect 137640 -1640 137860 -1590
rect 138140 -1410 138360 -1360
rect 138140 -1480 138150 -1410
rect 138350 -1480 138360 -1410
rect 138140 -1520 138360 -1480
rect 138140 -1590 138150 -1520
rect 138350 -1590 138360 -1520
rect 138140 -1640 138360 -1590
rect 138640 -1410 138860 -1360
rect 138640 -1480 138650 -1410
rect 138850 -1480 138860 -1410
rect 138640 -1520 138860 -1480
rect 138640 -1590 138650 -1520
rect 138850 -1590 138860 -1520
rect 138640 -1640 138860 -1590
rect 139140 -1410 139360 -1360
rect 139140 -1480 139150 -1410
rect 139350 -1480 139360 -1410
rect 139140 -1520 139360 -1480
rect 139140 -1590 139150 -1520
rect 139350 -1590 139360 -1520
rect 139140 -1640 139360 -1590
rect 139640 -1410 139860 -1360
rect 139640 -1480 139650 -1410
rect 139850 -1480 139860 -1410
rect 139640 -1520 139860 -1480
rect 139640 -1590 139650 -1520
rect 139850 -1590 139860 -1520
rect 139640 -1640 139860 -1590
rect 136000 -1650 140000 -1640
rect 136000 -1850 136020 -1650
rect 136090 -1850 136410 -1650
rect 136480 -1850 136520 -1650
rect 136590 -1850 136910 -1650
rect 136980 -1850 137020 -1650
rect 137090 -1850 137410 -1650
rect 137480 -1850 137520 -1650
rect 137590 -1850 137910 -1650
rect 137980 -1850 138020 -1650
rect 138090 -1850 138410 -1650
rect 138480 -1850 138520 -1650
rect 138590 -1850 138910 -1650
rect 138980 -1850 139020 -1650
rect 139090 -1850 139410 -1650
rect 139480 -1850 139520 -1650
rect 139590 -1850 139910 -1650
rect 139980 -1850 140000 -1650
rect 136000 -1860 140000 -1850
rect 136140 -1910 136360 -1860
rect 136140 -1980 136150 -1910
rect 136350 -1980 136360 -1910
rect 136140 -2000 136360 -1980
rect 136640 -1910 136860 -1860
rect 136640 -1980 136650 -1910
rect 136850 -1980 136860 -1910
rect 136640 -2000 136860 -1980
rect 137140 -1910 137360 -1860
rect 137140 -1980 137150 -1910
rect 137350 -1980 137360 -1910
rect 137140 -2000 137360 -1980
rect 137640 -1910 137860 -1860
rect 137640 -1980 137650 -1910
rect 137850 -1980 137860 -1910
rect 137640 -2000 137860 -1980
rect 138140 -1910 138360 -1860
rect 138140 -1980 138150 -1910
rect 138350 -1980 138360 -1910
rect 138140 -2000 138360 -1980
rect 138640 -1910 138860 -1860
rect 138640 -1980 138650 -1910
rect 138850 -1980 138860 -1910
rect 138640 -2000 138860 -1980
rect 139140 -1910 139360 -1860
rect 139140 -1980 139150 -1910
rect 139350 -1980 139360 -1910
rect 139140 -2000 139360 -1980
rect 139640 -1910 139860 -1860
rect 139640 -1980 139650 -1910
rect 139850 -1980 139860 -1910
rect 139640 -2000 139860 -1980
<< via2 >>
rect 17810 35810 18390 36190
rect 17010 35210 17590 35590
rect 17010 34610 17590 34990
rect 17810 34010 18390 34390
rect 14620 33220 15180 33780
<< metal3 >>
rect -11800 135600 -11600 139800
rect -5600 136600 -5400 139600
rect 600 137600 800 139600
rect 6800 138600 7000 139600
rect 6800 137800 8600 138600
rect 600 136800 7600 137600
rect -5600 135800 6600 136600
rect -11800 135595 -11204 135600
rect 3800 135595 5600 135600
rect -11800 134804 5600 135595
rect 3800 134800 5600 134804
rect -37000 129800 -20000 131000
rect -37000 125000 -16000 129800
rect -28000 118000 -16000 125000
rect -14000 129000 2000 129200
rect -14000 125000 -1200 129000
rect 1800 125000 2000 129000
rect -14000 124800 2000 125000
rect -14000 124000 2000 124200
rect -14000 120000 -1200 124000
rect 1800 120000 2000 124000
rect -14000 119800 2000 120000
rect -14000 119000 2000 119200
rect -14000 115000 -1200 119000
rect 1800 115000 2000 119000
rect -14000 114800 2000 115000
rect -14000 114000 2000 114200
rect -14000 110000 -1200 114000
rect 1800 110000 2000 114000
rect -14000 109800 2000 110000
rect -14000 109000 2000 109200
rect -14000 105000 -1200 109000
rect 1800 105000 2000 109000
rect -14000 104800 2000 105000
rect -14000 104000 2000 104200
rect -14000 100000 -1200 104000
rect 1800 100000 2000 104000
rect -14000 99800 2000 100000
rect -15800 48036 -15400 96600
rect 4800 96400 5600 134800
rect -15200 96000 5600 96400
rect -37000 46900 -32000 47000
rect -37000 40100 -35900 46900
rect -32100 40100 -32000 46900
rect -37000 40000 -32000 40100
rect -15200 39200 -14800 96000
rect 5800 95800 6600 135800
rect -14600 95400 6600 95800
rect -14600 39800 -14200 95400
rect 6800 95200 7600 136800
rect -14000 94800 7600 95200
rect -14000 40400 -13600 94800
rect 7800 94600 8600 137800
rect -13400 94200 8600 94600
rect -13400 41000 -13000 94200
rect 96200 49300 96600 86000
rect 96800 49500 97200 86000
rect 97400 49700 97800 86000
rect 98000 49900 98400 86000
rect 98600 50100 99000 86000
rect 98600 50000 100980 50100
rect 98000 49800 100240 49900
rect 97400 49600 99880 49700
rect 96800 49400 99040 49500
rect 96200 49200 98680 49300
rect 98500 49100 98680 49200
rect 98860 49100 99040 49400
rect 99700 49100 99880 49600
rect 100060 49100 100240 49800
rect 100800 49100 100980 50000
rect 92200 46000 97500 46400
rect -13400 40600 11600 41000
rect -14000 40000 11000 40400
rect -14600 39400 10400 39800
rect -15200 39199 -13800 39200
rect 9400 39199 9800 39200
rect -15200 38802 9800 39199
rect -15200 38800 -13800 38802
rect -28600 38200 9200 38600
rect -28600 32400 -28200 38200
rect 8800 35800 9200 38200
rect 9400 36400 9800 38802
rect 10000 37000 10400 39400
rect 10600 37600 11000 40000
rect 11200 38200 11600 40600
rect 11200 37800 14400 38200
rect 10600 37200 13800 37600
rect 10000 36600 13200 37000
rect 9400 36000 12600 36400
rect 8800 35400 12000 35800
rect 11600 33800 12000 35400
rect 12200 34400 12600 36000
rect 12800 35000 13200 36600
rect 13400 35600 13800 37200
rect 14000 36200 14400 37800
rect 14000 36190 18400 36200
rect 14000 35810 17810 36190
rect 18390 35810 18400 36190
rect 14000 35800 18400 35810
rect 13400 35590 17600 35600
rect 13400 35210 17010 35590
rect 17590 35210 17600 35590
rect 13400 35200 17600 35210
rect 12800 34990 17600 35000
rect 12800 34610 17010 34990
rect 17590 34610 17600 34990
rect 12800 34600 17600 34610
rect 12200 34390 18400 34400
rect 12200 34010 17810 34390
rect 18390 34010 18400 34390
rect 12200 34000 18400 34010
rect 11600 33780 15200 33800
rect 11600 33400 14620 33780
rect 14600 33220 14620 33400
rect 15180 33220 15200 33780
rect 14600 33200 15200 33220
rect 92200 27600 92800 46000
rect 97000 45280 97400 45300
rect 97000 45000 97020 45280
rect 89400 27000 92800 27600
rect 93200 44600 97020 45000
rect 89400 23400 90200 27000
rect 93200 26800 93800 44600
rect 97000 44020 97020 44600
rect 97380 44020 97400 45280
rect 97000 44000 97400 44020
rect 91600 26200 93800 26800
rect 91600 23400 92400 26200
rect 89000 22600 90200 23400
rect 91300 22600 92500 23400
rect 89800 5600 90600 12400
rect 90800 6800 91600 12400
rect 103400 8000 113800 8200
rect 103400 6800 103600 8000
rect 90800 6400 103600 6800
rect 113600 6400 113800 8000
rect 90800 5800 113800 6400
rect 89800 5000 113800 5600
rect 89800 4600 103600 5000
rect 103400 3400 103600 4600
rect 113600 3400 113800 5000
rect 103400 3200 113800 3400
<< via3 >>
rect -1200 125000 1800 129000
rect -1200 120000 1800 124000
rect -1200 115000 1800 119000
rect -1200 110000 1800 114000
rect -1200 105000 1800 109000
rect -1200 100000 1800 104000
rect -35900 40100 -32100 46900
rect 97020 44020 97380 45280
rect 103600 6400 113600 8000
rect 103600 3400 113600 5000
<< mimcap >>
rect -13800 128800 -2200 129000
rect -13800 125200 -13600 128800
rect -2400 125200 -2200 128800
rect -13800 125000 -2200 125200
rect -13800 123800 -2200 124000
rect -13800 120200 -13600 123800
rect -2400 120200 -2200 123800
rect -13800 120000 -2200 120200
rect -13800 118800 -2200 119000
rect -13800 115200 -13600 118800
rect -2400 115200 -2200 118800
rect -13800 115000 -2200 115200
rect -13800 113800 -2200 114000
rect -13800 110200 -13600 113800
rect -2400 110200 -2200 113800
rect -13800 110000 -2200 110200
rect -13800 108800 -2200 109000
rect -13800 105200 -13600 108800
rect -2400 105200 -2200 108800
rect -13800 105000 -2200 105200
rect -13800 103800 -2200 104000
rect -13800 100200 -13600 103800
rect -2400 100200 -2200 103800
rect -13800 100000 -2200 100200
<< mimcapcontact >>
rect -13600 125200 -2400 128800
rect -13600 120200 -2400 123800
rect -13600 115200 -2400 118800
rect -13600 110200 -2400 113800
rect -13600 105200 -2400 108800
rect -13600 100200 -2400 103800
<< metal4 >>
rect -31800 138000 -24400 140000
rect -35200 137800 -24000 138000
rect -35200 131800 -35000 137800
rect -24200 131800 -24000 137800
rect -35200 131600 -24000 131800
rect -14000 129000 -2000 129200
rect -16000 128800 -2000 129000
rect -16000 125200 -13600 128800
rect -2400 125200 -2000 128800
rect -16000 125000 -2000 125200
rect -14000 124800 -2000 125000
rect -1400 129000 2000 129200
rect -1400 125000 -1200 129000
rect 1800 125000 2000 129000
rect -1400 124800 2000 125000
rect -14000 124000 -2000 124200
rect -16000 123800 -2000 124000
rect -16000 120200 -13600 123800
rect -2400 120200 -2000 123800
rect -16000 120000 -2000 120200
rect -14000 119800 -2000 120000
rect -1400 124000 2000 124200
rect -1400 120000 -1200 124000
rect 1800 120000 2000 124000
rect -1400 119800 2000 120000
rect -14000 119000 -2000 119200
rect -16000 118800 -2000 119000
rect -16000 115200 -13600 118800
rect -2400 115200 -2000 118800
rect -16000 115000 -2000 115200
rect -14000 114800 -2000 115000
rect -1400 119000 2000 119200
rect -1400 115000 -1200 119000
rect 1800 115000 2000 119000
rect -1400 114800 2000 115000
rect -14000 114000 -2000 114200
rect -16000 113800 -2000 114000
rect -16000 110200 -13600 113800
rect -2400 110200 -2000 113800
rect -16000 110000 -2000 110200
rect -14000 109800 -2000 110000
rect -1400 114000 2000 114200
rect -1400 110000 -1200 114000
rect 1800 110000 2000 114000
rect -1400 109800 2000 110000
rect -14000 109000 -2000 109200
rect -16000 108800 -2000 109000
rect -16000 105200 -13600 108800
rect -2400 105200 -2000 108800
rect -16000 105000 -2000 105200
rect -14000 104800 -2000 105000
rect -1400 109000 2000 109200
rect -1400 105000 -1200 109000
rect 1800 105000 2000 109000
rect -1400 104800 2000 105000
rect -14000 104000 -2000 104200
rect -16000 103800 -2000 104000
rect -16000 100200 -13600 103800
rect -2400 100200 -2000 103800
rect -16000 100000 -2000 100200
rect -14000 99800 -2000 100000
rect -1400 104000 2000 104200
rect -1400 100000 -1200 104000
rect 1800 100000 2000 104000
rect -1400 99800 2000 100000
rect 100000 52000 102000 53000
rect 96000 50000 106000 52000
rect -36000 46900 -32000 47000
rect -36000 40100 -35900 46900
rect -32100 40100 -32000 46900
rect 97000 45280 97400 45300
rect 97000 44020 97020 45280
rect 97380 44020 97400 45280
rect 97000 44000 97400 44020
rect -36000 40000 -32000 40100
rect 96000 40000 106000 41000
rect -36600 39200 -36200 39400
rect -35600 39200 -34600 39400
rect -34200 39200 -33200 39400
rect -36800 39000 -36000 39200
rect -35600 39000 -34400 39200
rect -37000 38800 -35800 39000
rect -37000 37800 -36600 38800
rect -36200 37800 -35800 38800
rect -35600 38200 -35200 39000
rect -34800 38200 -34400 39000
rect -35600 38000 -34400 38200
rect -34200 39000 -33000 39200
rect -34200 38200 -33800 39000
rect -33400 38200 -33000 39000
rect -34200 38000 -33000 38200
rect -32800 39000 -31600 39400
rect -35600 37800 -34600 38000
rect -34200 37800 -33200 38000
rect -32800 37800 -32400 39000
rect -31400 38800 -31000 39400
rect -30600 39200 -30200 39400
rect -30800 38800 -30200 39200
rect -31400 38400 -30200 38800
rect -31400 38000 -30800 38400
rect -31400 37800 -31000 38000
rect -30600 37800 -30200 38400
rect -30000 39000 -29600 39400
rect -29200 39000 -28800 39400
rect -30000 38600 -28800 39000
rect -30000 38200 -29600 38600
rect -29200 38200 -28800 38600
rect -30000 38000 -28800 38200
rect -29800 37800 -29000 38000
rect 40000 28000 46000 34000
rect 41000 18600 53400 25400
rect 86400 22600 87300 24200
rect 94000 24100 100000 26000
rect 93700 23000 100000 24100
rect 93700 22600 94600 23000
rect 86400 22500 87400 22600
rect 86400 21900 86500 22500
rect 87300 21900 87400 22500
rect 86400 21800 87400 21900
rect 93700 22500 94700 22600
rect 93700 21900 93800 22500
rect 94600 21900 94700 22500
rect 93700 21800 94700 21900
rect 94800 19800 99000 19900
rect 86200 17300 86600 19500
rect 94800 16100 96100 19800
rect 36200 13800 40000 14000
rect 32000 9800 36000 10000
rect 14000 2600 18000 2800
rect 14000 400 14200 2600
rect 17800 400 18000 2600
rect 14000 200 18000 400
rect 32000 200 32200 9800
rect 34800 200 36000 9800
rect 38600 200 40000 13800
rect 96000 13300 96100 16100
rect 98900 13300 99000 19800
rect 96000 13100 99000 13300
rect 103200 8000 120200 9000
rect 103200 7000 103600 8000
rect 103400 6400 103600 7000
rect 113600 6400 120200 8000
rect 103400 6200 120200 6400
rect 113200 6000 120200 6200
rect 103400 5000 113800 5200
rect 103400 4000 103600 5000
rect 103200 3400 103600 4000
rect 113600 3400 116200 5000
rect 103200 2000 116200 3400
rect 32000 0 40000 200
rect 113200 -10000 116200 2000
rect 117200 -5000 120200 6000
rect 117200 -8000 132000 -5000
rect 113200 -13000 132000 -10000
rect 35600 -22600 36000 -22200
rect 36400 -22400 36800 -22200
rect 36200 -22600 36800 -22400
rect 35600 -23000 36600 -22600
rect 37000 -22800 37400 -22200
rect 38600 -22400 39600 -22200
rect 38400 -22600 39600 -22400
rect 35600 -23400 36000 -23000
rect 36400 -23400 36800 -23000
rect 35600 -23600 36800 -23400
rect 37000 -23200 38000 -22800
rect 37000 -23400 37400 -23200
rect 38400 -23400 38800 -22600
rect 39200 -22800 39600 -22600
rect 39000 -23000 39600 -22800
rect 39800 -22800 40200 -22200
rect 40600 -22400 41000 -22200
rect 40400 -22800 41000 -22400
rect 39800 -23200 41000 -22800
rect 39200 -23400 39600 -23200
rect 35600 -23800 36600 -23600
rect 37000 -23800 38200 -23400
rect 38400 -23600 39600 -23400
rect 39800 -23600 40400 -23200
rect 38600 -23800 39400 -23600
rect 39800 -23800 40200 -23600
rect 40600 -23800 41000 -23200
rect 41200 -22400 42200 -22200
rect 41200 -22600 42400 -22400
rect 41200 -23400 41600 -22600
rect 42000 -23400 42400 -22600
rect 41200 -23600 42400 -23400
rect 41200 -23800 42200 -23600
<< via4 >>
rect -35000 131800 -24200 137800
rect -1200 125000 1800 129000
rect -1200 120000 1800 124000
rect -1200 115000 1800 119000
rect -1200 110000 1800 114000
rect -1200 105000 1800 109000
rect -1200 100000 1800 104000
rect -35900 40100 -32100 46900
rect 86500 21900 87300 22500
rect 93800 21900 94600 22500
rect 14200 400 17800 2600
rect 32200 200 34800 9800
rect 36000 200 38600 13800
rect 96100 13300 98900 19800
<< mimcap2 >>
rect -13800 128800 -2200 129000
rect -13800 125200 -13600 128800
rect -2400 125200 -2200 128800
rect -13800 125000 -2200 125200
rect -13800 123800 -2200 124000
rect -13800 120200 -13600 123800
rect -2400 120200 -2200 123800
rect -13800 120000 -2200 120200
rect -13800 118800 -2200 119000
rect -13800 115200 -13600 118800
rect -2400 115200 -2200 118800
rect -13800 115000 -2200 115200
rect -13800 113800 -2200 114000
rect -13800 110200 -13600 113800
rect -2400 110200 -2200 113800
rect -13800 110000 -2200 110200
rect -13800 108800 -2200 109000
rect -13800 105200 -13600 108800
rect -2400 105200 -2200 108800
rect -13800 105000 -2200 105200
rect -13800 103800 -2200 104000
rect -13800 100200 -13600 103800
rect -2400 100200 -2200 103800
rect -13800 100000 -2200 100200
rect 41200 25000 53200 25200
rect 41200 19000 41400 25000
rect 53000 19000 53200 25000
rect 41200 18800 53200 19000
<< mimcap2contact >>
rect -13600 125200 -2400 128800
rect -13600 120200 -2400 123800
rect -13600 115200 -2400 118800
rect -13600 110200 -2400 113800
rect -13600 105200 -2400 108800
rect -13600 100200 -2400 103800
rect 41400 19000 53000 25000
<< metal5 >>
rect -36000 137800 -23000 138000
rect -36000 131800 -35000 137800
rect -24200 131800 -23000 137800
rect -36000 126000 -23000 131800
rect -14000 129000 2000 129200
rect -14000 128800 -1200 129000
rect -14000 125200 -13600 128800
rect -2400 125200 -1200 128800
rect -14000 125000 -1200 125200
rect 1800 125000 2000 129000
rect -14000 124800 2000 125000
rect -1400 124200 2000 124800
rect -14000 124000 2000 124200
rect -14000 123800 -1200 124000
rect -14000 120200 -13600 123800
rect -2400 120200 -1200 123800
rect -14000 120000 -1200 120200
rect 1800 120000 2000 124000
rect -14000 119800 2000 120000
rect -1400 119200 2000 119800
rect -14000 119000 2000 119200
rect -14000 118800 -1200 119000
rect -14000 115200 -13600 118800
rect -2400 115200 -1200 118800
rect -14000 115000 -1200 115200
rect 1800 115000 2000 119000
rect -14000 114800 2000 115000
rect -1400 114200 2000 114800
rect -14000 114000 2000 114200
rect -14000 113800 -1200 114000
rect -14000 110200 -13600 113800
rect -2400 110200 -1200 113800
rect -14000 110000 -1200 110200
rect 1800 110000 2000 114000
rect -14000 109800 2000 110000
rect -1400 109200 2000 109800
rect -14000 109000 2000 109200
rect -14000 108800 -1200 109000
rect -14000 105200 -13600 108800
rect -2400 105200 -1200 108800
rect -14000 105000 -1200 105200
rect 1800 105000 2000 109000
rect -14000 104800 2000 105000
rect -1400 104200 2000 104800
rect -14000 104000 2000 104200
rect -14000 103800 -1200 104000
rect -14000 100200 -13600 103800
rect -2400 100200 -1200 103800
rect -14000 100000 -1200 100200
rect 1800 100000 2000 104000
rect -14000 99800 2000 100000
rect -1400 95000 2000 99800
rect -27000 91000 76000 95000
rect -27000 90000 -23000 91000
rect -22000 90000 -18000 91000
rect -1400 90000 2000 91000
rect 60000 90000 64000 91000
rect 66000 90000 70000 91000
rect 72000 90000 76000 91000
rect -27000 86000 76000 90000
rect -27000 78000 -23000 86000
rect -22000 78000 -18000 86000
rect -27000 74000 -18000 78000
rect -27000 66000 -23000 74000
rect -22000 66000 -18000 74000
rect -27000 62000 -18000 66000
rect -27000 54000 -23000 62000
rect -22000 54000 -18000 62000
rect -27000 50000 -18000 54000
rect -27000 47000 -23000 50000
rect -22000 47000 -18000 50000
rect -36000 46900 -32000 47000
rect -36000 40100 -35900 46900
rect -32100 46000 -32000 46900
rect -27000 46000 -18000 47000
rect -32100 41000 -18000 46000
rect 60000 84000 64000 86000
rect 66000 84000 70000 86000
rect 72000 84000 76000 86000
rect 60000 80000 76000 84000
rect 60000 76000 64000 80000
rect 66000 76000 70000 80000
rect 72000 76000 76000 80000
rect 60000 72000 76000 76000
rect 60000 68000 64000 72000
rect 66000 68000 70000 72000
rect 72000 68000 76000 72000
rect 60000 64000 76000 68000
rect 60000 60000 64000 64000
rect 66000 60000 70000 64000
rect 72000 60000 76000 64000
rect 60000 56000 76000 60000
rect 60000 52000 64000 56000
rect 66000 52000 70000 56000
rect 72000 52000 76000 56000
rect 60000 48400 102000 52000
rect 60000 48000 97000 48400
rect 101600 48000 102000 48400
rect 60000 44000 64000 48000
rect 66000 44000 70000 48000
rect 72000 44000 76000 48000
rect -32100 40100 -32000 41000
rect -36000 40000 -32000 40100
rect 60000 40000 76000 44000
rect 56000 36000 64000 40000
rect 66000 36000 70000 40000
rect 72000 36000 76000 40000
rect 56000 34000 76000 36000
rect 40000 32000 76000 34000
rect 40000 28000 62000 32000
rect 41000 25000 54800 25400
rect 41000 19000 41400 25000
rect 53000 21200 54800 25000
rect 86400 22500 87400 22600
rect 86400 21900 86500 22500
rect 87300 21900 87400 22500
rect 86400 21800 87400 21900
rect 93700 22500 94700 22600
rect 93700 21900 93800 22500
rect 94600 21900 94700 22500
rect 93700 21800 94700 21900
rect 53000 19200 65400 21200
rect 96000 19800 99000 19900
rect 53000 19000 54800 19200
rect 41000 18600 54800 19000
rect 14000 2600 18000 2800
rect 14000 400 14200 2600
rect 17800 400 18000 2600
rect 14000 -12000 18000 400
rect 96000 13300 96100 19800
rect 98900 13300 99000 19800
rect 96000 12000 99000 13300
rect 96000 -11000 100600 12000
use MIXER_5G_core  MIXER_5G_core_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/MIXER
timestamp 1659323209
transform 0 -1 90200 1 0 13460
box -1160 -4800 9880 3800
use OSC_5GHz_1  OSC_5GHz_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/OSC
timestamp 1661649873
transform 1 0 86000 0 -1 52000
box 10000 -21000 68022 34000
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501465
transform 1 0 -4000 0 1 77700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_1
timestamp 1659501465
transform 1 0 -4000 0 1 75700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_2
timestamp 1659501465
transform 1 0 -4000 0 1 73700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_3
timestamp 1659501465
transform 1 0 -4000 0 1 71700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_4
timestamp 1659501465
transform 1 0 -4000 0 1 63700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_5
timestamp 1659501465
transform 1 0 -4000 0 1 65700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_6
timestamp 1659501465
transform 1 0 -4000 0 1 67700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_7
timestamp 1659501465
transform 1 0 -4000 0 1 69700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_8
timestamp 1659501465
transform 1 0 -4000 0 1 55700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_9
timestamp 1659501465
transform 1 0 -4000 0 1 57700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_10
timestamp 1659501465
transform 1 0 -4000 0 1 59700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_11
timestamp 1659501465
transform 1 0 -4000 0 1 61700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_12
timestamp 1659501465
transform 1 0 -4000 0 1 47700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_13
timestamp 1659501465
transform 1 0 -4000 0 1 49700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_14
timestamp 1659501465
transform 1 0 -4000 0 1 51700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_15
timestamp 1659501465
transform 1 0 -4000 0 1 53700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_16
timestamp 1659501465
transform 1 0 120000 0 1 15700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_17
timestamp 1659501465
transform 1 0 116000 0 1 19700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_18
timestamp 1659501465
transform 1 0 112000 0 1 23700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_19
timestamp 1659501465
transform 1 0 108000 0 1 31700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_20
timestamp 1659501465
transform 1 0 108000 0 1 33700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_21
timestamp 1659501465
transform 1 0 108000 0 1 35700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_22
timestamp 1659501465
transform 1 0 108000 0 1 37700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_23
timestamp 1659501465
transform 1 0 104000 0 1 39700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_24
timestamp 1659501465
transform 1 0 102000 0 1 39700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_25
timestamp 1659501465
transform 1 0 100000 0 1 39700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_26
timestamp 1659501465
transform 1 0 98000 0 1 39700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_27
timestamp 1659501465
transform 1 0 96000 0 1 39700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_28
timestamp 1659501465
transform 1 0 86000 0 1 25700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_29
timestamp 1659501465
transform 1 0 88000 0 1 29700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_30
timestamp 1659501465
transform 1 0 90000 0 1 29700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_31
timestamp 1659501465
transform 1 0 94000 0 1 27700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_32
timestamp 1659501465
transform 1 0 94000 0 1 29700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_33
timestamp 1659501465
transform 1 0 94000 0 1 31700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_34
timestamp 1659501465
transform 1 0 94000 0 1 33700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_35
timestamp 1659501465
transform 1 0 94000 0 1 35700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_36
timestamp 1659501465
transform 1 0 94000 0 1 37700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_37
timestamp 1659501465
transform 1 0 150000 0 1 15700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_38
timestamp 1659501465
transform 1 0 154000 0 1 19700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_39
timestamp 1659501465
transform 1 0 158000 0 1 23700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_40
timestamp 1659501465
transform 1 0 158000 0 1 69700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_41
timestamp 1659501465
transform 1 0 54000 0 1 43700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_42
timestamp 1659501465
transform 1 0 50000 0 1 39700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_43
timestamp 1659501465
transform 1 0 54000 0 1 73700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_44
timestamp 1659501465
transform 1 0 50000 0 1 77700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_45
timestamp 1659501465
transform 1 0 46000 0 1 81700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_46
timestamp 1659501465
transform 1 0 42000 0 1 85700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_47
timestamp 1659501465
transform 1 0 8000 0 1 85700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_48
timestamp 1659501465
transform 1 0 4000 0 1 81700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_49
timestamp 1659501465
transform 1 0 -2000 0 1 77700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_50
timestamp 1659501465
transform 1 0 0 0 1 77700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_51
timestamp 1659501465
transform 1 0 -2000 0 1 75700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_52
timestamp 1659501465
transform 1 0 -2000 0 1 47700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_53
timestamp 1659501465
transform 1 0 0 0 1 43700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_54
timestamp 1659501465
transform 1 0 -24000 0 1 3700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_55
timestamp 1659501465
transform 1 0 0 0 1 45700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_56
timestamp 1659501465
transform 1 0 2000 0 1 43700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_57
timestamp 1659501465
transform 1 0 -24000 0 1 1700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_58
timestamp 1659501465
transform 1 0 -24000 0 1 -300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_59
timestamp 1659501465
transform 1 0 -22000 0 1 29700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_60
timestamp 1659501465
transform 1 0 -18000 0 1 33700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_61
timestamp 1659501465
transform 1 0 -14000 0 1 37700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_62
timestamp 1659501465
transform 1 0 -22000 0 1 3700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_63
timestamp 1659501465
transform 1 0 -18000 0 1 -300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_64
timestamp 1659501465
transform 1 0 -12000 0 1 -4300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_65
timestamp 1659501465
transform 1 0 10000 0 1 -4300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_66
timestamp 1659501465
transform 1 0 8000 0 1 -4300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_67
timestamp 1659501465
transform 1 0 10000 0 1 -2300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_68
timestamp 1659501465
transform 1 0 60000 0 1 25700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_69
timestamp 1659501465
transform 1 0 64000 0 1 29700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_70
timestamp 1659501465
transform 1 0 82000 0 1 29700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_71
timestamp 1659501465
transform 1 0 64000 0 1 7700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_72
timestamp 1659501465
transform 1 0 104000 0 1 -300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_73
timestamp 1659501465
transform 1 0 68000 0 1 3700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_74
timestamp 1659501465
transform 1 0 84000 0 1 3700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_75
timestamp 1659501465
transform 1 0 86000 0 1 3700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_76
timestamp 1659501465
transform 1 0 86000 0 1 5700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_77
timestamp 1659501465
transform 1 0 46000 0 1 35700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_78
timestamp 1659501465
transform 1 0 -24000 0 1 5700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_79
timestamp 1659501465
transform 1 0 -24000 0 1 7700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_80
timestamp 1659501465
transform 1 0 -24000 0 1 9700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_81
timestamp 1659501465
transform 1 0 -24000 0 1 11700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_82
timestamp 1659501465
transform 1 0 -24000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_83
timestamp 1659501465
transform 1 0 -24000 0 1 15700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_84
timestamp 1659501465
transform 1 0 -24000 0 1 17700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_85
timestamp 1659501465
transform 1 0 -24000 0 1 19700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_86
timestamp 1659501465
transform 1 0 -24000 0 1 21700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_87
timestamp 1659501465
transform 1 0 -24000 0 1 23700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_88
timestamp 1659501465
transform 1 0 -24000 0 1 25700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_89
timestamp 1659501465
transform 1 0 -24000 0 1 27700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_90
timestamp 1659501465
transform 1 0 -24000 0 1 29700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_91
timestamp 1659501465
transform 1 0 -20000 0 1 31700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_92
timestamp 1659501465
transform 1 0 -20000 0 1 33700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_93
timestamp 1659501465
transform 1 0 -16000 0 1 35700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_94
timestamp 1659501465
transform 1 0 -16000 0 1 37700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_95
timestamp 1659501465
transform 1 0 106000 0 1 -300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_96
timestamp 1659501465
transform 1 0 108000 0 1 -300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_97
timestamp 1659501465
transform 1 0 110000 0 1 -300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_98
timestamp 1659501465
transform 1 0 104000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_99
timestamp 1659501465
transform 1 0 106000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_100
timestamp 1659501465
transform 1 0 108000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_101
timestamp 1659501465
transform 1 0 110000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_102
timestamp 1659501465
transform 1 0 112000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_103
timestamp 1659501465
transform 1 0 114000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_104
timestamp 1659501465
transform 1 0 116000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_105
timestamp 1659501465
transform 1 0 118000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_106
timestamp 1659501465
transform 1 0 120000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_107
timestamp 1659501465
transform 1 0 122000 0 1 13700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_108
timestamp 1659501465
transform 1 0 122000 0 1 11700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_109
timestamp 1659501465
transform 1 0 92000 0 1 1700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_110
timestamp 1659501465
transform 1 0 92000 0 1 -300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_111
timestamp 1659501465
transform 1 0 92000 0 1 -2300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_112
timestamp 1659501465
transform 1 0 92000 0 1 -4300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_113
timestamp 1659501465
transform 1 0 92000 0 1 -6300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_114
timestamp 1659501465
transform 1 0 92000 0 1 -8300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_115
timestamp 1659501465
transform 1 0 92000 0 1 -10300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_116
timestamp 1659501465
transform 1 0 92000 0 1 -12300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_117
timestamp 1659501465
transform 1 0 154000 0 1 73700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_118
timestamp 1659501465
transform 1 0 150000 0 1 77700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_119
timestamp 1659501465
transform 1 0 120000 0 1 77700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_120
timestamp 1659501465
transform 1 0 116000 0 1 73700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_121
timestamp 1659501465
transform 1 0 112000 0 1 69700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_122
timestamp 1659501465
transform 1 0 108000 0 1 65700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_123
timestamp 1659501465
transform 1 0 122000 0 1 77700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_124
timestamp 1659501465
transform 1 0 100000 0 1 57700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_125
timestamp 1659501465
transform 1 0 100000 0 1 55700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_126
timestamp 1659501465
transform 1 0 100000 0 1 53700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_127
timestamp 1659501465
transform 1 0 100000 0 1 52700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_128
timestamp 1659501465
transform 1 0 -20000 0 1 41700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_129
timestamp 1659501465
transform 1 0 -18000 0 1 41700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_130
timestamp 1659501465
transform 1 0 -24000 0 1 41700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_131
timestamp 1659501465
transform 1 0 -22000 0 1 41700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_132
timestamp 1659501465
transform 1 0 -28000 0 1 41700
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_133
timestamp 1659501465
transform 1 0 -26000 0 1 41700
box 0 -1700 2000 300
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501637
transform 1 0 56000 0 1 10000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_1
timestamp 1659501637
transform 1 0 56000 0 1 14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_2
timestamp 1659501637
transform 1 0 56000 0 1 22000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_3
timestamp 1659501637
transform 1 0 60000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_4
timestamp 1659501637
transform 1 0 64000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_5
timestamp 1659501637
transform 1 0 60000 0 1 26000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_6
timestamp 1659501637
transform 1 0 56000 0 1 42000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_7
timestamp 1659501637
transform 1 0 56000 0 1 46000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_8
timestamp 1659501637
transform 1 0 56000 0 1 50000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_9
timestamp 1659501637
transform 1 0 56000 0 1 54000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_10
timestamp 1659501637
transform 1 0 56000 0 1 58000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_11
timestamp 1659501637
transform 1 0 56000 0 1 62000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_12
timestamp 1659501637
transform 1 0 56000 0 1 66000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_13
timestamp 1659501637
transform 1 0 56000 0 1 70000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_14
timestamp 1659501637
transform 1 0 112000 0 1 14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_15
timestamp 1659501637
transform 1 0 52000 0 1 78000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_16
timestamp 1659501637
transform 1 0 52000 0 1 74000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_17
timestamp 1659501637
transform 1 0 48000 0 1 78000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_18
timestamp 1659501637
transform 1 0 44000 0 1 82000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_19
timestamp 1659501637
transform 1 0 0 0 1 82000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_20
timestamp 1659501637
transform 1 0 0 0 1 78000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_21
timestamp 1659501637
transform 1 0 56000 0 1 74000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_22
timestamp 1659501637
transform 1 0 56000 0 1 78000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_23
timestamp 1659501637
transform 1 0 56000 0 1 82000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_24
timestamp 1659501637
transform 1 0 56000 0 1 86000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_25
timestamp 1659501637
transform 1 0 52000 0 1 90000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_26
timestamp 1659501637
transform 1 0 48000 0 1 90000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_27
timestamp 1659501637
transform 1 0 4000 0 1 82000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_28
timestamp 1659501637
transform 1 0 -12000 0 1 78000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_29
timestamp 1659501637
transform 1 0 -12000 0 1 82000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_30
timestamp 1659501637
transform 1 0 -12000 0 1 86000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_31
timestamp 1659501637
transform 1 0 -12000 0 1 90000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_32
timestamp 1659501637
transform 1 0 -28000 0 1 42000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_33
timestamp 1659501637
transform 1 0 -4000 0 1 42000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_34
timestamp 1659501637
transform 1 0 116000 0 1 14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_35
timestamp 1659501637
transform 1 0 112000 0 1 18000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_36
timestamp 1659501637
transform 1 0 128000 0 1 6000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_37
timestamp 1659501637
transform 1 0 -20000 0 1 34000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_38
timestamp 1659501637
transform 1 0 -22000 0 1 -2000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_39
timestamp 1659501637
transform 1 0 -16000 0 1 -14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_40
timestamp 1659501637
transform 1 0 -20000 0 1 -14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_41
timestamp 1659501637
transform 1 0 -28000 0 1 -14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_42
timestamp 1659501637
transform 1 0 -24000 0 1 -14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_43
timestamp 1659501637
transform 1 0 36000 0 1 -14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_44
timestamp 1659501637
transform 1 0 36000 0 1 -10000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_45
timestamp 1659501637
transform 1 0 36000 0 1 -6000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_46
timestamp 1659501637
transform 1 0 36000 0 1 -2000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_47
timestamp 1659501637
transform 1 0 60000 0 1 10000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_48
timestamp 1659501637
transform 1 0 36000 0 1 10000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_49
timestamp 1659501637
transform 1 0 36000 0 1 14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_50
timestamp 1659501637
transform 1 0 48000 0 1 26000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_51
timestamp 1659501637
transform 1 0 48000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_52
timestamp 1659501637
transform 1 0 48000 0 1 34000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_53
timestamp 1659501637
transform 1 0 68000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_54
timestamp 1659501637
transform 1 0 44000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_55
timestamp 1659501637
transform 1 0 132000 0 1 6000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_56
timestamp 1659501637
transform 1 0 92000 0 1 54000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_57
timestamp 1659501637
transform 1 0 128000 0 1 10000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_58
timestamp 1659501637
transform 1 0 132000 0 1 10000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_59
timestamp 1659501637
transform 1 0 92000 0 1 50000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_60
timestamp 1659501637
transform 1 0 96000 0 1 26000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_61
timestamp 1659501637
transform 1 0 100000 0 1 26000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_62
timestamp 1659501637
transform 1 0 100000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_63
timestamp 1659501637
transform 1 0 104000 0 1 26000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_64
timestamp 1659501637
transform 1 0 104000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_65
timestamp 1659501637
transform 1 0 108000 0 1 26000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_66
timestamp 1659501637
transform 1 0 104000 0 1 34000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_67
timestamp 1659501637
transform 1 0 100000 0 1 34000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_68
timestamp 1659501637
transform 1 0 96000 0 1 34000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_69
timestamp 1659501637
transform 1 0 84000 0 1 26000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_70
timestamp 1659501637
transform 1 0 72000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_71
timestamp 1659501637
transform 1 0 76000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_72
timestamp 1659501637
transform 1 0 80000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_73
timestamp 1659501637
transform 1 0 84000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_74
timestamp 1659501637
transform 1 0 88000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_75
timestamp 1659501637
transform 1 0 64000 0 1 2000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_76
timestamp 1659501637
transform 1 0 56000 0 1 90000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_77
timestamp 1659501637
transform 1 0 -20000 0 1 106000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_78
timestamp 1659501637
transform 1 0 104000 0 1 22000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_79
timestamp 1659501637
transform 1 0 96000 0 1 30000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_80
timestamp 1659501637
transform 1 0 108000 0 1 22000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_81
timestamp 1659501637
transform 1 0 100000 0 1 22000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_82
timestamp 1659501637
transform 1 0 44000 0 1 26000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_83
timestamp 1659501637
transform 1 0 -20000 0 1 42000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_84
timestamp 1659501637
transform 1 0 -20000 0 1 46000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_85
timestamp 1659501637
transform 1 0 -12000 0 1 42000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_86
timestamp 1659501637
transform 1 0 -8000 0 1 42000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_87
timestamp 1659501637
transform 1 0 -20000 0 1 102000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_88
timestamp 1659501637
transform 1 0 156000 0 1 14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_89
timestamp 1659501637
transform 1 0 102000 0 1 50000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_90
timestamp 1659501637
transform 1 0 102000 0 1 54000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_91
timestamp 1659501637
transform 1 0 156000 0 1 18000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_92
timestamp 1659501637
transform 1 0 152000 0 1 14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_93
timestamp 1659501637
transform 1 0 104000 0 1 -6000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_94
timestamp 1659501637
transform 1 0 108000 0 1 -6000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_95
timestamp 1659501637
transform 1 0 88000 0 1 -2000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_96
timestamp 1659501637
transform 1 0 88000 0 1 -6000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_97
timestamp 1659501637
transform 1 0 88000 0 1 -10000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_98
timestamp 1659501637
transform 1 0 -28000 0 1 -2000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_99
timestamp 1659501637
transform 1 0 -28000 0 1 2000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_100
timestamp 1659501637
transform 1 0 -28000 0 1 6000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_101
timestamp 1659501637
transform 1 0 -28000 0 1 10000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_102
timestamp 1659501637
transform 1 0 -28000 0 1 14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_103
timestamp 1659501637
transform 1 0 -28000 0 1 18000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_104
timestamp 1659501637
transform 1 0 -28000 0 1 22000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_105
timestamp 1659501637
transform 1 0 -28000 0 1 26000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_106
timestamp 1659501637
transform 1 0 156000 0 1 70000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_107
timestamp 1659501637
transform 1 0 152000 0 1 74000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_108
timestamp 1659501637
transform 1 0 60000 0 1 14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_109
timestamp 1659501637
transform 1 0 88000 0 1 -14000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_110
timestamp 1659501637
transform 1 0 124000 0 1 10000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_111
timestamp 1659501637
transform 1 0 124000 0 1 6000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_112
timestamp 1659501637
transform 1 0 124000 0 1 2000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_113
timestamp 1659501637
transform 1 0 124000 0 1 -2000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_114
timestamp 1659501637
transform 1 0 -20000 0 1 50000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_115
timestamp 1659501637
transform 1 0 -20000 0 1 54000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_116
timestamp 1659501637
transform 1 0 -20000 0 1 58000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_117
timestamp 1659501637
transform 1 0 -20000 0 1 62000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_118
timestamp 1659501637
transform 1 0 -20000 0 1 66000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_119
timestamp 1659501637
transform 1 0 -20000 0 1 70000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_120
timestamp 1659501637
transform 1 0 -20000 0 1 74000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_121
timestamp 1659501637
transform 1 0 -20000 0 1 78000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_122
timestamp 1659501637
transform 1 0 -20000 0 1 82000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_123
timestamp 1659501637
transform 1 0 -20000 0 1 86000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_124
timestamp 1659501637
transform 1 0 -20000 0 1 90000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_125
timestamp 1659501637
transform 1 0 112000 0 1 74000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_126
timestamp 1659501637
transform 1 0 104000 0 1 66000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_127
timestamp 1659501637
transform 1 0 100000 0 1 62000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_128
timestamp 1659501637
transform 1 0 156000 0 1 74000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_129
timestamp 1659501637
transform 1 0 100000 0 1 58000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_130
timestamp 1659501637
transform 1 0 104000 0 1 58000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_131
timestamp 1659501637
transform 1 0 104000 0 1 62000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_132
timestamp 1659501637
transform 1 0 108000 0 1 66000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_133
timestamp 1659501637
transform 1 0 112000 0 1 70000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_134
timestamp 1659501637
transform 1 0 116000 0 1 74000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_135
timestamp 1659501637
transform 1 0 100000 0 1 66000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_136
timestamp 1659501637
transform 1 0 100000 0 1 70000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_137
timestamp 1659501637
transform 1 0 100000 0 1 74000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_138
timestamp 1659501637
transform 1 0 100000 0 1 78000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_139
timestamp 1659501637
transform 1 0 100000 0 1 82000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_140
timestamp 1659501637
transform 1 0 -20000 0 1 98000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_141
timestamp 1659501637
transform 1 0 -20000 0 1 94000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_142
timestamp 1659501637
transform 1 0 -20000 0 1 122000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_143
timestamp 1659501637
transform 1 0 -20000 0 1 118000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_144
timestamp 1659501637
transform 1 0 -20000 0 1 114000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_145
timestamp 1659501637
transform 1 0 -20000 0 1 110000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_146
timestamp 1659501637
transform 1 0 -20000 0 1 126000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_147
timestamp 1659501637
transform 1 0 -24000 0 1 42000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660792292
transform 1 0 40000 0 1 -6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_1
timestamp 1660792292
transform 1 0 48000 0 1 -6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_2
timestamp 1660792292
transform 1 0 40000 0 1 2000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_3
timestamp 1660792292
transform 1 0 48000 0 1 2000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_4
timestamp 1660792292
transform 1 0 40000 0 1 10000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_5
timestamp 1660792292
transform 1 0 48000 0 1 10000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_6
timestamp 1660792292
transform 1 0 56000 0 1 -6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_7
timestamp 1660792292
transform 1 0 64000 0 1 -6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_8
timestamp 1660792292
transform 1 0 72000 0 1 -6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_9
timestamp 1660792292
transform 1 0 80000 0 1 -6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_10
timestamp 1660792292
transform 1 0 80000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_11
timestamp 1660792292
transform 1 0 72000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_12
timestamp 1660792292
transform 1 0 64000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_13
timestamp 1660792292
transform 1 0 56000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_14
timestamp 1660792292
transform 1 0 48000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_15
timestamp 1660792292
transform 1 0 40000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_16
timestamp 1660792292
transform 1 0 56000 0 1 2000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_17
timestamp 1660792292
transform 1 0 52000 0 1 26000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_18
timestamp 1660792292
transform 1 0 52000 0 1 34000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_19
timestamp 1660792292
transform 1 0 60000 0 1 34000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_20
timestamp 1660792292
transform 1 0 84000 0 1 34000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_21
timestamp 1660792292
transform 1 0 68000 0 1 34000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_22
timestamp 1660792292
transform 1 0 76000 0 1 34000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_23
timestamp 1660792292
transform 1 0 60000 0 1 42000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_24
timestamp 1660792292
transform 1 0 68000 0 1 42000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_25
timestamp 1660792292
transform 1 0 76000 0 1 42000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_26
timestamp 1660792292
transform 1 0 48000 0 1 82000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_27
timestamp 1660792292
transform 1 0 84000 0 1 42000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_28
timestamp 1660792292
transform 1 0 60000 0 1 50000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_29
timestamp 1660792292
transform 1 0 68000 0 1 50000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_30
timestamp 1660792292
transform 1 0 76000 0 1 50000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_31
timestamp 1660792292
transform 1 0 84000 0 1 50000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_32
timestamp 1660792292
transform 1 0 60000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_33
timestamp 1660792292
transform 1 0 40000 0 1 86000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_34
timestamp 1660792292
transform 1 0 32000 0 1 86000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_35
timestamp 1660792292
transform 1 0 24000 0 1 86000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_36
timestamp 1660792292
transform 1 0 16000 0 1 86000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_37
timestamp 1660792292
transform 1 0 8000 0 1 86000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_38
timestamp 1660792292
transform 1 0 0 0 1 86000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_39
timestamp 1660792292
transform 1 0 -8000 0 1 86000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_40
timestamp 1660792292
transform 1 0 -8000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_41
timestamp 1660792292
transform 1 0 -12000 0 1 70000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_42
timestamp 1660792292
transform 1 0 -12000 0 1 62000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_43
timestamp 1660792292
transform 1 0 -12000 0 1 54000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_44
timestamp 1660792292
transform 1 0 -12000 0 1 46000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_45
timestamp 1660792292
transform 1 0 104000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_47
timestamp 1660792292
transform 1 0 -28000 0 1 30000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_48
timestamp 1660792292
transform 1 0 60000 0 1 86000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_49
timestamp 1660792292
transform 1 0 60000 0 1 70000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_50
timestamp 1660792292
transform 1 0 60000 0 1 62000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_51
timestamp 1660792292
transform 1 0 60000 0 1 58000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_52
timestamp 1660792292
transform 1 0 -28000 0 1 94000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_53
timestamp 1660792292
transform 1 0 -28000 0 1 86000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_54
timestamp 1660792292
transform 1 0 -28000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_55
timestamp 1660792292
transform 1 0 -28000 0 1 70000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_56
timestamp 1660792292
transform 1 0 -28000 0 1 62000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_57
timestamp 1660792292
transform 1 0 -28000 0 1 54000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_58
timestamp 1660792292
transform 1 0 -28000 0 1 46000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_59
timestamp 1660792292
transform 1 0 136000 0 1 6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_60
timestamp 1660792292
transform 1 0 144000 0 1 6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_61
timestamp 1660792292
transform 1 0 152000 0 1 6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_62
timestamp 1660792292
transform 1 0 160000 0 1 6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_63
timestamp 1660792292
transform 1 0 160000 0 1 14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_64
timestamp 1660792292
transform 1 0 160000 0 1 30000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_65
timestamp 1660792292
transform 1 0 -28000 0 1 -10000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_66
timestamp 1660792292
transform 1 0 -20000 0 1 -10000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_67
timestamp 1660792292
transform 1 0 -12000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_68
timestamp 1660792292
transform 1 0 -4000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_69
timestamp 1660792292
transform 1 0 4000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_70
timestamp 1660792292
transform 1 0 20000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_71
timestamp 1660792292
transform 1 0 28000 0 1 -14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_72
timestamp 1660792292
transform 1 0 20000 0 1 -6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_73
timestamp 1660792292
transform 1 0 28000 0 1 -6000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_74
timestamp 1660792292
transform 1 0 32000 0 1 2000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_75
timestamp 1660792292
transform 1 0 160000 0 1 22000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_76
timestamp 1660792292
transform 1 0 160000 0 1 46000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_77
timestamp 1660792292
transform 1 0 160000 0 1 38000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_78
timestamp 1660792292
transform 1 0 160000 0 1 62000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_79
timestamp 1660792292
transform 1 0 160000 0 1 54000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_80
timestamp 1660792292
transform 1 0 160000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_81
timestamp 1660792292
transform 1 0 160000 0 1 70000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_82
timestamp 1660792292
transform 1 0 152000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_83
timestamp 1660792292
transform 1 0 144000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_84
timestamp 1660792292
transform 1 0 136000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_85
timestamp 1660792292
transform 1 0 128000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_86
timestamp 1660792292
transform 1 0 120000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_87
timestamp 1660792292
transform 1 0 104000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_88
timestamp 1660792292
transform 1 0 112000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_89
timestamp 1660792292
transform 1 0 -28000 0 1 102000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_90
timestamp 1660792292
transform 1 0 -28000 0 1 110000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_91
timestamp 1660792292
transform 1 0 104000 0 1 14000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_92
timestamp 1660792292
transform 1 0 -28000 0 1 118000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_93
timestamp 1660792292
transform 1 0 104000 0 1 70000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_94
timestamp 1660792292
transform 1 0 88000 0 1 62000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_95
timestamp 1660792292
transform 1 0 88000 0 1 70000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_96
timestamp 1660792292
transform 1 0 128000 0 1 -2000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_97
timestamp 1660792292
transform 1 0 88000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_98
timestamp 1660792292
transform 1 0 80000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_99
timestamp 1660792292
transform 1 0 68000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_100
timestamp 1660792292
transform 1 0 72000 0 1 78000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_101
timestamp 1660792292
transform 1 0 68000 0 1 70000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_102
timestamp 1660792292
transform 1 0 72000 0 1 70000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_103
timestamp 1660792292
transform 1 0 80000 0 1 70000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_104
timestamp 1660792292
transform 1 0 68000 0 1 62000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_105
timestamp 1660792292
transform 1 0 72000 0 1 62000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_106
timestamp 1660792292
transform 1 0 80000 0 1 62000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_107
timestamp 1660792292
transform 1 0 68000 0 1 58000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_108
timestamp 1660792292
transform 1 0 72000 0 1 58000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_109
timestamp 1660792292
transform 1 0 80000 0 1 58000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_110
timestamp 1660792292
transform 1 0 88000 0 1 58000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_111
timestamp 1660792292
transform 1 0 136000 0 1 -2000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_112
timestamp 1660792292
transform 1 0 144000 0 1 -2000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_113
timestamp 1660792292
transform 1 0 152000 0 1 -2000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_114
timestamp 1660792292
transform 1 0 160000 0 1 -2000
box 0 0 8000 8000
use lna_complete_2  lna_complete_2_1 ~/openmpw/Project-Yatsuhashi-Chip1/mag/LNA
timestamp 1662004902
transform -1 0 20100 0 1 13800
box -31800 -16200 37700 70200
use octal_ind_0p700n_5GHz_1  octal_ind_0p700n_5GHz_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1661738380
transform -1 0 54600 0 -1 -4600
box -33800 -32500 -8800 -10100
<< end >>
