magic
tech sky130B
magscale 1 2
timestamp 1659838778
<< error_p >>
rect -1386 617 -1328 623
rect -1268 617 -1210 623
rect -1150 617 -1092 623
rect -1032 617 -974 623
rect -914 617 -856 623
rect -796 617 -738 623
rect -678 617 -620 623
rect -560 617 -502 623
rect -442 617 -384 623
rect -324 617 -266 623
rect -206 617 -148 623
rect -88 617 -30 623
rect 30 617 88 623
rect 148 617 206 623
rect 266 617 324 623
rect 384 617 442 623
rect 502 617 560 623
rect 620 617 678 623
rect 738 617 796 623
rect 856 617 914 623
rect 974 617 1032 623
rect 1092 617 1150 623
rect 1210 617 1268 623
rect 1328 617 1386 623
rect -1386 583 -1374 617
rect -1268 583 -1256 617
rect -1150 583 -1138 617
rect -1032 583 -1020 617
rect -914 583 -902 617
rect -796 583 -784 617
rect -678 583 -666 617
rect -560 583 -548 617
rect -442 583 -430 617
rect -324 583 -312 617
rect -206 583 -194 617
rect -88 583 -76 617
rect 30 583 42 617
rect 148 583 160 617
rect 266 583 278 617
rect 384 583 396 617
rect 502 583 514 617
rect 620 583 632 617
rect 738 583 750 617
rect 856 583 868 617
rect 974 583 986 617
rect 1092 583 1104 617
rect 1210 583 1222 617
rect 1328 583 1340 617
rect -1386 577 -1328 583
rect -1268 577 -1210 583
rect -1150 577 -1092 583
rect -1032 577 -974 583
rect -914 577 -856 583
rect -796 577 -738 583
rect -678 577 -620 583
rect -560 577 -502 583
rect -442 577 -384 583
rect -324 577 -266 583
rect -206 577 -148 583
rect -88 577 -30 583
rect 30 577 88 583
rect 148 577 206 583
rect 266 577 324 583
rect 384 577 442 583
rect 502 577 560 583
rect 620 577 678 583
rect 738 577 796 583
rect 856 577 914 583
rect 974 577 1032 583
rect 1092 577 1150 583
rect 1210 577 1268 583
rect 1328 577 1386 583
rect -1386 289 -1328 295
rect -1268 289 -1210 295
rect -1150 289 -1092 295
rect -1032 289 -974 295
rect -914 289 -856 295
rect -796 289 -738 295
rect -678 289 -620 295
rect -560 289 -502 295
rect -442 289 -384 295
rect -324 289 -266 295
rect -206 289 -148 295
rect -88 289 -30 295
rect 30 289 88 295
rect 148 289 206 295
rect 266 289 324 295
rect 384 289 442 295
rect 502 289 560 295
rect 620 289 678 295
rect 738 289 796 295
rect 856 289 914 295
rect 974 289 1032 295
rect 1092 289 1150 295
rect 1210 289 1268 295
rect 1328 289 1386 295
rect -1386 255 -1374 289
rect -1268 255 -1256 289
rect -1150 255 -1138 289
rect -1032 255 -1020 289
rect -914 255 -902 289
rect -796 255 -784 289
rect -678 255 -666 289
rect -560 255 -548 289
rect -442 255 -430 289
rect -324 255 -312 289
rect -206 255 -194 289
rect -88 255 -76 289
rect 30 255 42 289
rect 148 255 160 289
rect 266 255 278 289
rect 384 255 396 289
rect 502 255 514 289
rect 620 255 632 289
rect 738 255 750 289
rect 856 255 868 289
rect 974 255 986 289
rect 1092 255 1104 289
rect 1210 255 1222 289
rect 1328 255 1340 289
rect -1386 249 -1328 255
rect -1268 249 -1210 255
rect -1150 249 -1092 255
rect -1032 249 -974 255
rect -914 249 -856 255
rect -796 249 -738 255
rect -678 249 -620 255
rect -560 249 -502 255
rect -442 249 -384 255
rect -324 249 -266 255
rect -206 249 -148 255
rect -88 249 -30 255
rect 30 249 88 255
rect 148 249 206 255
rect 266 249 324 255
rect 384 249 442 255
rect 502 249 560 255
rect 620 249 678 255
rect 738 249 796 255
rect 856 249 914 255
rect 974 249 1032 255
rect 1092 249 1150 255
rect 1210 249 1268 255
rect 1328 249 1386 255
rect -1386 181 -1328 187
rect -1268 181 -1210 187
rect -1150 181 -1092 187
rect -1032 181 -974 187
rect -914 181 -856 187
rect -796 181 -738 187
rect -678 181 -620 187
rect -560 181 -502 187
rect -442 181 -384 187
rect -324 181 -266 187
rect -206 181 -148 187
rect -88 181 -30 187
rect 30 181 88 187
rect 148 181 206 187
rect 266 181 324 187
rect 384 181 442 187
rect 502 181 560 187
rect 620 181 678 187
rect 738 181 796 187
rect 856 181 914 187
rect 974 181 1032 187
rect 1092 181 1150 187
rect 1210 181 1268 187
rect 1328 181 1386 187
rect -1386 147 -1374 181
rect -1268 147 -1256 181
rect -1150 147 -1138 181
rect -1032 147 -1020 181
rect -914 147 -902 181
rect -796 147 -784 181
rect -678 147 -666 181
rect -560 147 -548 181
rect -442 147 -430 181
rect -324 147 -312 181
rect -206 147 -194 181
rect -88 147 -76 181
rect 30 147 42 181
rect 148 147 160 181
rect 266 147 278 181
rect 384 147 396 181
rect 502 147 514 181
rect 620 147 632 181
rect 738 147 750 181
rect 856 147 868 181
rect 974 147 986 181
rect 1092 147 1104 181
rect 1210 147 1222 181
rect 1328 147 1340 181
rect -1386 141 -1328 147
rect -1268 141 -1210 147
rect -1150 141 -1092 147
rect -1032 141 -974 147
rect -914 141 -856 147
rect -796 141 -738 147
rect -678 141 -620 147
rect -560 141 -502 147
rect -442 141 -384 147
rect -324 141 -266 147
rect -206 141 -148 147
rect -88 141 -30 147
rect 30 141 88 147
rect 148 141 206 147
rect 266 141 324 147
rect 384 141 442 147
rect 502 141 560 147
rect 620 141 678 147
rect 738 141 796 147
rect 856 141 914 147
rect 974 141 1032 147
rect 1092 141 1150 147
rect 1210 141 1268 147
rect 1328 141 1386 147
rect -1386 -147 -1328 -141
rect -1268 -147 -1210 -141
rect -1150 -147 -1092 -141
rect -1032 -147 -974 -141
rect -914 -147 -856 -141
rect -796 -147 -738 -141
rect -678 -147 -620 -141
rect -560 -147 -502 -141
rect -442 -147 -384 -141
rect -324 -147 -266 -141
rect -206 -147 -148 -141
rect -88 -147 -30 -141
rect 30 -147 88 -141
rect 148 -147 206 -141
rect 266 -147 324 -141
rect 384 -147 442 -141
rect 502 -147 560 -141
rect 620 -147 678 -141
rect 738 -147 796 -141
rect 856 -147 914 -141
rect 974 -147 1032 -141
rect 1092 -147 1150 -141
rect 1210 -147 1268 -141
rect 1328 -147 1386 -141
rect -1386 -181 -1374 -147
rect -1268 -181 -1256 -147
rect -1150 -181 -1138 -147
rect -1032 -181 -1020 -147
rect -914 -181 -902 -147
rect -796 -181 -784 -147
rect -678 -181 -666 -147
rect -560 -181 -548 -147
rect -442 -181 -430 -147
rect -324 -181 -312 -147
rect -206 -181 -194 -147
rect -88 -181 -76 -147
rect 30 -181 42 -147
rect 148 -181 160 -147
rect 266 -181 278 -147
rect 384 -181 396 -147
rect 502 -181 514 -147
rect 620 -181 632 -147
rect 738 -181 750 -147
rect 856 -181 868 -147
rect 974 -181 986 -147
rect 1092 -181 1104 -147
rect 1210 -181 1222 -147
rect 1328 -181 1340 -147
rect -1386 -187 -1328 -181
rect -1268 -187 -1210 -181
rect -1150 -187 -1092 -181
rect -1032 -187 -974 -181
rect -914 -187 -856 -181
rect -796 -187 -738 -181
rect -678 -187 -620 -181
rect -560 -187 -502 -181
rect -442 -187 -384 -181
rect -324 -187 -266 -181
rect -206 -187 -148 -181
rect -88 -187 -30 -181
rect 30 -187 88 -181
rect 148 -187 206 -181
rect 266 -187 324 -181
rect 384 -187 442 -181
rect 502 -187 560 -181
rect 620 -187 678 -181
rect 738 -187 796 -181
rect 856 -187 914 -181
rect 974 -187 1032 -181
rect 1092 -187 1150 -181
rect 1210 -187 1268 -181
rect 1328 -187 1386 -181
rect -1386 -255 -1328 -249
rect -1268 -255 -1210 -249
rect -1150 -255 -1092 -249
rect -1032 -255 -974 -249
rect -914 -255 -856 -249
rect -796 -255 -738 -249
rect -678 -255 -620 -249
rect -560 -255 -502 -249
rect -442 -255 -384 -249
rect -324 -255 -266 -249
rect -206 -255 -148 -249
rect -88 -255 -30 -249
rect 30 -255 88 -249
rect 148 -255 206 -249
rect 266 -255 324 -249
rect 384 -255 442 -249
rect 502 -255 560 -249
rect 620 -255 678 -249
rect 738 -255 796 -249
rect 856 -255 914 -249
rect 974 -255 1032 -249
rect 1092 -255 1150 -249
rect 1210 -255 1268 -249
rect 1328 -255 1386 -249
rect -1386 -289 -1374 -255
rect -1268 -289 -1256 -255
rect -1150 -289 -1138 -255
rect -1032 -289 -1020 -255
rect -914 -289 -902 -255
rect -796 -289 -784 -255
rect -678 -289 -666 -255
rect -560 -289 -548 -255
rect -442 -289 -430 -255
rect -324 -289 -312 -255
rect -206 -289 -194 -255
rect -88 -289 -76 -255
rect 30 -289 42 -255
rect 148 -289 160 -255
rect 266 -289 278 -255
rect 384 -289 396 -255
rect 502 -289 514 -255
rect 620 -289 632 -255
rect 738 -289 750 -255
rect 856 -289 868 -255
rect 974 -289 986 -255
rect 1092 -289 1104 -255
rect 1210 -289 1222 -255
rect 1328 -289 1340 -255
rect -1386 -295 -1328 -289
rect -1268 -295 -1210 -289
rect -1150 -295 -1092 -289
rect -1032 -295 -974 -289
rect -914 -295 -856 -289
rect -796 -295 -738 -289
rect -678 -295 -620 -289
rect -560 -295 -502 -289
rect -442 -295 -384 -289
rect -324 -295 -266 -289
rect -206 -295 -148 -289
rect -88 -295 -30 -289
rect 30 -295 88 -289
rect 148 -295 206 -289
rect 266 -295 324 -289
rect 384 -295 442 -289
rect 502 -295 560 -289
rect 620 -295 678 -289
rect 738 -295 796 -289
rect 856 -295 914 -289
rect 974 -295 1032 -289
rect 1092 -295 1150 -289
rect 1210 -295 1268 -289
rect 1328 -295 1386 -289
rect -1386 -583 -1328 -577
rect -1268 -583 -1210 -577
rect -1150 -583 -1092 -577
rect -1032 -583 -974 -577
rect -914 -583 -856 -577
rect -796 -583 -738 -577
rect -678 -583 -620 -577
rect -560 -583 -502 -577
rect -442 -583 -384 -577
rect -324 -583 -266 -577
rect -206 -583 -148 -577
rect -88 -583 -30 -577
rect 30 -583 88 -577
rect 148 -583 206 -577
rect 266 -583 324 -577
rect 384 -583 442 -577
rect 502 -583 560 -577
rect 620 -583 678 -577
rect 738 -583 796 -577
rect 856 -583 914 -577
rect 974 -583 1032 -577
rect 1092 -583 1150 -577
rect 1210 -583 1268 -577
rect 1328 -583 1386 -577
rect -1386 -617 -1374 -583
rect -1268 -617 -1256 -583
rect -1150 -617 -1138 -583
rect -1032 -617 -1020 -583
rect -914 -617 -902 -583
rect -796 -617 -784 -583
rect -678 -617 -666 -583
rect -560 -617 -548 -583
rect -442 -617 -430 -583
rect -324 -617 -312 -583
rect -206 -617 -194 -583
rect -88 -617 -76 -583
rect 30 -617 42 -583
rect 148 -617 160 -583
rect 266 -617 278 -583
rect 384 -617 396 -583
rect 502 -617 514 -583
rect 620 -617 632 -583
rect 738 -617 750 -583
rect 856 -617 868 -583
rect 974 -617 986 -583
rect 1092 -617 1104 -583
rect 1210 -617 1222 -583
rect 1328 -617 1340 -583
rect -1386 -623 -1328 -617
rect -1268 -623 -1210 -617
rect -1150 -623 -1092 -617
rect -1032 -623 -974 -617
rect -914 -623 -856 -617
rect -796 -623 -738 -617
rect -678 -623 -620 -617
rect -560 -623 -502 -617
rect -442 -623 -384 -617
rect -324 -623 -266 -617
rect -206 -623 -148 -617
rect -88 -623 -30 -617
rect 30 -623 88 -617
rect 148 -623 206 -617
rect 266 -623 324 -617
rect 384 -623 442 -617
rect 502 -623 560 -617
rect 620 -623 678 -617
rect 738 -623 796 -617
rect 856 -623 914 -617
rect 974 -623 1032 -617
rect 1092 -623 1150 -617
rect 1210 -623 1268 -617
rect 1328 -623 1386 -617
<< nwell >>
rect -1583 -755 1583 755
<< pmos >>
rect -1387 336 -1327 536
rect -1269 336 -1209 536
rect -1151 336 -1091 536
rect -1033 336 -973 536
rect -915 336 -855 536
rect -797 336 -737 536
rect -679 336 -619 536
rect -561 336 -501 536
rect -443 336 -383 536
rect -325 336 -265 536
rect -207 336 -147 536
rect -89 336 -29 536
rect 29 336 89 536
rect 147 336 207 536
rect 265 336 325 536
rect 383 336 443 536
rect 501 336 561 536
rect 619 336 679 536
rect 737 336 797 536
rect 855 336 915 536
rect 973 336 1033 536
rect 1091 336 1151 536
rect 1209 336 1269 536
rect 1327 336 1387 536
rect -1387 -100 -1327 100
rect -1269 -100 -1209 100
rect -1151 -100 -1091 100
rect -1033 -100 -973 100
rect -915 -100 -855 100
rect -797 -100 -737 100
rect -679 -100 -619 100
rect -561 -100 -501 100
rect -443 -100 -383 100
rect -325 -100 -265 100
rect -207 -100 -147 100
rect -89 -100 -29 100
rect 29 -100 89 100
rect 147 -100 207 100
rect 265 -100 325 100
rect 383 -100 443 100
rect 501 -100 561 100
rect 619 -100 679 100
rect 737 -100 797 100
rect 855 -100 915 100
rect 973 -100 1033 100
rect 1091 -100 1151 100
rect 1209 -100 1269 100
rect 1327 -100 1387 100
rect -1387 -536 -1327 -336
rect -1269 -536 -1209 -336
rect -1151 -536 -1091 -336
rect -1033 -536 -973 -336
rect -915 -536 -855 -336
rect -797 -536 -737 -336
rect -679 -536 -619 -336
rect -561 -536 -501 -336
rect -443 -536 -383 -336
rect -325 -536 -265 -336
rect -207 -536 -147 -336
rect -89 -536 -29 -336
rect 29 -536 89 -336
rect 147 -536 207 -336
rect 265 -536 325 -336
rect 383 -536 443 -336
rect 501 -536 561 -336
rect 619 -536 679 -336
rect 737 -536 797 -336
rect 855 -536 915 -336
rect 973 -536 1033 -336
rect 1091 -536 1151 -336
rect 1209 -536 1269 -336
rect 1327 -536 1387 -336
<< pdiff >>
rect -1445 524 -1387 536
rect -1445 348 -1433 524
rect -1399 348 -1387 524
rect -1445 336 -1387 348
rect -1327 524 -1269 536
rect -1327 348 -1315 524
rect -1281 348 -1269 524
rect -1327 336 -1269 348
rect -1209 524 -1151 536
rect -1209 348 -1197 524
rect -1163 348 -1151 524
rect -1209 336 -1151 348
rect -1091 524 -1033 536
rect -1091 348 -1079 524
rect -1045 348 -1033 524
rect -1091 336 -1033 348
rect -973 524 -915 536
rect -973 348 -961 524
rect -927 348 -915 524
rect -973 336 -915 348
rect -855 524 -797 536
rect -855 348 -843 524
rect -809 348 -797 524
rect -855 336 -797 348
rect -737 524 -679 536
rect -737 348 -725 524
rect -691 348 -679 524
rect -737 336 -679 348
rect -619 524 -561 536
rect -619 348 -607 524
rect -573 348 -561 524
rect -619 336 -561 348
rect -501 524 -443 536
rect -501 348 -489 524
rect -455 348 -443 524
rect -501 336 -443 348
rect -383 524 -325 536
rect -383 348 -371 524
rect -337 348 -325 524
rect -383 336 -325 348
rect -265 524 -207 536
rect -265 348 -253 524
rect -219 348 -207 524
rect -265 336 -207 348
rect -147 524 -89 536
rect -147 348 -135 524
rect -101 348 -89 524
rect -147 336 -89 348
rect -29 524 29 536
rect -29 348 -17 524
rect 17 348 29 524
rect -29 336 29 348
rect 89 524 147 536
rect 89 348 101 524
rect 135 348 147 524
rect 89 336 147 348
rect 207 524 265 536
rect 207 348 219 524
rect 253 348 265 524
rect 207 336 265 348
rect 325 524 383 536
rect 325 348 337 524
rect 371 348 383 524
rect 325 336 383 348
rect 443 524 501 536
rect 443 348 455 524
rect 489 348 501 524
rect 443 336 501 348
rect 561 524 619 536
rect 561 348 573 524
rect 607 348 619 524
rect 561 336 619 348
rect 679 524 737 536
rect 679 348 691 524
rect 725 348 737 524
rect 679 336 737 348
rect 797 524 855 536
rect 797 348 809 524
rect 843 348 855 524
rect 797 336 855 348
rect 915 524 973 536
rect 915 348 927 524
rect 961 348 973 524
rect 915 336 973 348
rect 1033 524 1091 536
rect 1033 348 1045 524
rect 1079 348 1091 524
rect 1033 336 1091 348
rect 1151 524 1209 536
rect 1151 348 1163 524
rect 1197 348 1209 524
rect 1151 336 1209 348
rect 1269 524 1327 536
rect 1269 348 1281 524
rect 1315 348 1327 524
rect 1269 336 1327 348
rect 1387 524 1445 536
rect 1387 348 1399 524
rect 1433 348 1445 524
rect 1387 336 1445 348
rect -1445 88 -1387 100
rect -1445 -88 -1433 88
rect -1399 -88 -1387 88
rect -1445 -100 -1387 -88
rect -1327 88 -1269 100
rect -1327 -88 -1315 88
rect -1281 -88 -1269 88
rect -1327 -100 -1269 -88
rect -1209 88 -1151 100
rect -1209 -88 -1197 88
rect -1163 -88 -1151 88
rect -1209 -100 -1151 -88
rect -1091 88 -1033 100
rect -1091 -88 -1079 88
rect -1045 -88 -1033 88
rect -1091 -100 -1033 -88
rect -973 88 -915 100
rect -973 -88 -961 88
rect -927 -88 -915 88
rect -973 -100 -915 -88
rect -855 88 -797 100
rect -855 -88 -843 88
rect -809 -88 -797 88
rect -855 -100 -797 -88
rect -737 88 -679 100
rect -737 -88 -725 88
rect -691 -88 -679 88
rect -737 -100 -679 -88
rect -619 88 -561 100
rect -619 -88 -607 88
rect -573 -88 -561 88
rect -619 -100 -561 -88
rect -501 88 -443 100
rect -501 -88 -489 88
rect -455 -88 -443 88
rect -501 -100 -443 -88
rect -383 88 -325 100
rect -383 -88 -371 88
rect -337 -88 -325 88
rect -383 -100 -325 -88
rect -265 88 -207 100
rect -265 -88 -253 88
rect -219 -88 -207 88
rect -265 -100 -207 -88
rect -147 88 -89 100
rect -147 -88 -135 88
rect -101 -88 -89 88
rect -147 -100 -89 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 89 88 147 100
rect 89 -88 101 88
rect 135 -88 147 88
rect 89 -100 147 -88
rect 207 88 265 100
rect 207 -88 219 88
rect 253 -88 265 88
rect 207 -100 265 -88
rect 325 88 383 100
rect 325 -88 337 88
rect 371 -88 383 88
rect 325 -100 383 -88
rect 443 88 501 100
rect 443 -88 455 88
rect 489 -88 501 88
rect 443 -100 501 -88
rect 561 88 619 100
rect 561 -88 573 88
rect 607 -88 619 88
rect 561 -100 619 -88
rect 679 88 737 100
rect 679 -88 691 88
rect 725 -88 737 88
rect 679 -100 737 -88
rect 797 88 855 100
rect 797 -88 809 88
rect 843 -88 855 88
rect 797 -100 855 -88
rect 915 88 973 100
rect 915 -88 927 88
rect 961 -88 973 88
rect 915 -100 973 -88
rect 1033 88 1091 100
rect 1033 -88 1045 88
rect 1079 -88 1091 88
rect 1033 -100 1091 -88
rect 1151 88 1209 100
rect 1151 -88 1163 88
rect 1197 -88 1209 88
rect 1151 -100 1209 -88
rect 1269 88 1327 100
rect 1269 -88 1281 88
rect 1315 -88 1327 88
rect 1269 -100 1327 -88
rect 1387 88 1445 100
rect 1387 -88 1399 88
rect 1433 -88 1445 88
rect 1387 -100 1445 -88
rect -1445 -348 -1387 -336
rect -1445 -524 -1433 -348
rect -1399 -524 -1387 -348
rect -1445 -536 -1387 -524
rect -1327 -348 -1269 -336
rect -1327 -524 -1315 -348
rect -1281 -524 -1269 -348
rect -1327 -536 -1269 -524
rect -1209 -348 -1151 -336
rect -1209 -524 -1197 -348
rect -1163 -524 -1151 -348
rect -1209 -536 -1151 -524
rect -1091 -348 -1033 -336
rect -1091 -524 -1079 -348
rect -1045 -524 -1033 -348
rect -1091 -536 -1033 -524
rect -973 -348 -915 -336
rect -973 -524 -961 -348
rect -927 -524 -915 -348
rect -973 -536 -915 -524
rect -855 -348 -797 -336
rect -855 -524 -843 -348
rect -809 -524 -797 -348
rect -855 -536 -797 -524
rect -737 -348 -679 -336
rect -737 -524 -725 -348
rect -691 -524 -679 -348
rect -737 -536 -679 -524
rect -619 -348 -561 -336
rect -619 -524 -607 -348
rect -573 -524 -561 -348
rect -619 -536 -561 -524
rect -501 -348 -443 -336
rect -501 -524 -489 -348
rect -455 -524 -443 -348
rect -501 -536 -443 -524
rect -383 -348 -325 -336
rect -383 -524 -371 -348
rect -337 -524 -325 -348
rect -383 -536 -325 -524
rect -265 -348 -207 -336
rect -265 -524 -253 -348
rect -219 -524 -207 -348
rect -265 -536 -207 -524
rect -147 -348 -89 -336
rect -147 -524 -135 -348
rect -101 -524 -89 -348
rect -147 -536 -89 -524
rect -29 -348 29 -336
rect -29 -524 -17 -348
rect 17 -524 29 -348
rect -29 -536 29 -524
rect 89 -348 147 -336
rect 89 -524 101 -348
rect 135 -524 147 -348
rect 89 -536 147 -524
rect 207 -348 265 -336
rect 207 -524 219 -348
rect 253 -524 265 -348
rect 207 -536 265 -524
rect 325 -348 383 -336
rect 325 -524 337 -348
rect 371 -524 383 -348
rect 325 -536 383 -524
rect 443 -348 501 -336
rect 443 -524 455 -348
rect 489 -524 501 -348
rect 443 -536 501 -524
rect 561 -348 619 -336
rect 561 -524 573 -348
rect 607 -524 619 -348
rect 561 -536 619 -524
rect 679 -348 737 -336
rect 679 -524 691 -348
rect 725 -524 737 -348
rect 679 -536 737 -524
rect 797 -348 855 -336
rect 797 -524 809 -348
rect 843 -524 855 -348
rect 797 -536 855 -524
rect 915 -348 973 -336
rect 915 -524 927 -348
rect 961 -524 973 -348
rect 915 -536 973 -524
rect 1033 -348 1091 -336
rect 1033 -524 1045 -348
rect 1079 -524 1091 -348
rect 1033 -536 1091 -524
rect 1151 -348 1209 -336
rect 1151 -524 1163 -348
rect 1197 -524 1209 -348
rect 1151 -536 1209 -524
rect 1269 -348 1327 -336
rect 1269 -524 1281 -348
rect 1315 -524 1327 -348
rect 1269 -536 1327 -524
rect 1387 -348 1445 -336
rect 1387 -524 1399 -348
rect 1433 -524 1445 -348
rect 1387 -536 1445 -524
<< pdiffc >>
rect -1433 348 -1399 524
rect -1315 348 -1281 524
rect -1197 348 -1163 524
rect -1079 348 -1045 524
rect -961 348 -927 524
rect -843 348 -809 524
rect -725 348 -691 524
rect -607 348 -573 524
rect -489 348 -455 524
rect -371 348 -337 524
rect -253 348 -219 524
rect -135 348 -101 524
rect -17 348 17 524
rect 101 348 135 524
rect 219 348 253 524
rect 337 348 371 524
rect 455 348 489 524
rect 573 348 607 524
rect 691 348 725 524
rect 809 348 843 524
rect 927 348 961 524
rect 1045 348 1079 524
rect 1163 348 1197 524
rect 1281 348 1315 524
rect 1399 348 1433 524
rect -1433 -88 -1399 88
rect -1315 -88 -1281 88
rect -1197 -88 -1163 88
rect -1079 -88 -1045 88
rect -961 -88 -927 88
rect -843 -88 -809 88
rect -725 -88 -691 88
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
rect 691 -88 725 88
rect 809 -88 843 88
rect 927 -88 961 88
rect 1045 -88 1079 88
rect 1163 -88 1197 88
rect 1281 -88 1315 88
rect 1399 -88 1433 88
rect -1433 -524 -1399 -348
rect -1315 -524 -1281 -348
rect -1197 -524 -1163 -348
rect -1079 -524 -1045 -348
rect -961 -524 -927 -348
rect -843 -524 -809 -348
rect -725 -524 -691 -348
rect -607 -524 -573 -348
rect -489 -524 -455 -348
rect -371 -524 -337 -348
rect -253 -524 -219 -348
rect -135 -524 -101 -348
rect -17 -524 17 -348
rect 101 -524 135 -348
rect 219 -524 253 -348
rect 337 -524 371 -348
rect 455 -524 489 -348
rect 573 -524 607 -348
rect 691 -524 725 -348
rect 809 -524 843 -348
rect 927 -524 961 -348
rect 1045 -524 1079 -348
rect 1163 -524 1197 -348
rect 1281 -524 1315 -348
rect 1399 -524 1433 -348
<< nsubdiff >>
rect -1547 685 -1451 719
rect 1451 685 1547 719
rect -1547 623 -1513 685
rect 1513 623 1547 685
rect -1547 -685 -1513 -623
rect 1513 -685 1547 -623
rect -1547 -719 -1451 -685
rect 1451 -719 1547 -685
<< nsubdiffcont >>
rect -1451 685 1451 719
rect -1547 -623 -1513 623
rect 1513 -623 1547 623
rect -1451 -719 1451 -685
<< poly >>
rect -1390 617 -1324 633
rect -1390 583 -1374 617
rect -1340 583 -1324 617
rect -1390 567 -1324 583
rect -1272 617 -1206 633
rect -1272 583 -1256 617
rect -1222 583 -1206 617
rect -1272 567 -1206 583
rect -1154 617 -1088 633
rect -1154 583 -1138 617
rect -1104 583 -1088 617
rect -1154 567 -1088 583
rect -1036 617 -970 633
rect -1036 583 -1020 617
rect -986 583 -970 617
rect -1036 567 -970 583
rect -918 617 -852 633
rect -918 583 -902 617
rect -868 583 -852 617
rect -918 567 -852 583
rect -800 617 -734 633
rect -800 583 -784 617
rect -750 583 -734 617
rect -800 567 -734 583
rect -682 617 -616 633
rect -682 583 -666 617
rect -632 583 -616 617
rect -682 567 -616 583
rect -564 617 -498 633
rect -564 583 -548 617
rect -514 583 -498 617
rect -564 567 -498 583
rect -446 617 -380 633
rect -446 583 -430 617
rect -396 583 -380 617
rect -446 567 -380 583
rect -328 617 -262 633
rect -328 583 -312 617
rect -278 583 -262 617
rect -328 567 -262 583
rect -210 617 -144 633
rect -210 583 -194 617
rect -160 583 -144 617
rect -210 567 -144 583
rect -92 617 -26 633
rect -92 583 -76 617
rect -42 583 -26 617
rect -92 567 -26 583
rect 26 617 92 633
rect 26 583 42 617
rect 76 583 92 617
rect 26 567 92 583
rect 144 617 210 633
rect 144 583 160 617
rect 194 583 210 617
rect 144 567 210 583
rect 262 617 328 633
rect 262 583 278 617
rect 312 583 328 617
rect 262 567 328 583
rect 380 617 446 633
rect 380 583 396 617
rect 430 583 446 617
rect 380 567 446 583
rect 498 617 564 633
rect 498 583 514 617
rect 548 583 564 617
rect 498 567 564 583
rect 616 617 682 633
rect 616 583 632 617
rect 666 583 682 617
rect 616 567 682 583
rect 734 617 800 633
rect 734 583 750 617
rect 784 583 800 617
rect 734 567 800 583
rect 852 617 918 633
rect 852 583 868 617
rect 902 583 918 617
rect 852 567 918 583
rect 970 617 1036 633
rect 970 583 986 617
rect 1020 583 1036 617
rect 970 567 1036 583
rect 1088 617 1154 633
rect 1088 583 1104 617
rect 1138 583 1154 617
rect 1088 567 1154 583
rect 1206 617 1272 633
rect 1206 583 1222 617
rect 1256 583 1272 617
rect 1206 567 1272 583
rect 1324 617 1390 633
rect 1324 583 1340 617
rect 1374 583 1390 617
rect 1324 567 1390 583
rect -1387 536 -1327 567
rect -1269 536 -1209 567
rect -1151 536 -1091 567
rect -1033 536 -973 567
rect -915 536 -855 567
rect -797 536 -737 567
rect -679 536 -619 567
rect -561 536 -501 567
rect -443 536 -383 567
rect -325 536 -265 567
rect -207 536 -147 567
rect -89 536 -29 567
rect 29 536 89 567
rect 147 536 207 567
rect 265 536 325 567
rect 383 536 443 567
rect 501 536 561 567
rect 619 536 679 567
rect 737 536 797 567
rect 855 536 915 567
rect 973 536 1033 567
rect 1091 536 1151 567
rect 1209 536 1269 567
rect 1327 536 1387 567
rect -1387 305 -1327 336
rect -1269 305 -1209 336
rect -1151 305 -1091 336
rect -1033 305 -973 336
rect -915 305 -855 336
rect -797 305 -737 336
rect -679 305 -619 336
rect -561 305 -501 336
rect -443 305 -383 336
rect -325 305 -265 336
rect -207 305 -147 336
rect -89 305 -29 336
rect 29 305 89 336
rect 147 305 207 336
rect 265 305 325 336
rect 383 305 443 336
rect 501 305 561 336
rect 619 305 679 336
rect 737 305 797 336
rect 855 305 915 336
rect 973 305 1033 336
rect 1091 305 1151 336
rect 1209 305 1269 336
rect 1327 305 1387 336
rect -1390 289 -1324 305
rect -1390 255 -1374 289
rect -1340 255 -1324 289
rect -1390 239 -1324 255
rect -1272 289 -1206 305
rect -1272 255 -1256 289
rect -1222 255 -1206 289
rect -1272 239 -1206 255
rect -1154 289 -1088 305
rect -1154 255 -1138 289
rect -1104 255 -1088 289
rect -1154 239 -1088 255
rect -1036 289 -970 305
rect -1036 255 -1020 289
rect -986 255 -970 289
rect -1036 239 -970 255
rect -918 289 -852 305
rect -918 255 -902 289
rect -868 255 -852 289
rect -918 239 -852 255
rect -800 289 -734 305
rect -800 255 -784 289
rect -750 255 -734 289
rect -800 239 -734 255
rect -682 289 -616 305
rect -682 255 -666 289
rect -632 255 -616 289
rect -682 239 -616 255
rect -564 289 -498 305
rect -564 255 -548 289
rect -514 255 -498 289
rect -564 239 -498 255
rect -446 289 -380 305
rect -446 255 -430 289
rect -396 255 -380 289
rect -446 239 -380 255
rect -328 289 -262 305
rect -328 255 -312 289
rect -278 255 -262 289
rect -328 239 -262 255
rect -210 289 -144 305
rect -210 255 -194 289
rect -160 255 -144 289
rect -210 239 -144 255
rect -92 289 -26 305
rect -92 255 -76 289
rect -42 255 -26 289
rect -92 239 -26 255
rect 26 289 92 305
rect 26 255 42 289
rect 76 255 92 289
rect 26 239 92 255
rect 144 289 210 305
rect 144 255 160 289
rect 194 255 210 289
rect 144 239 210 255
rect 262 289 328 305
rect 262 255 278 289
rect 312 255 328 289
rect 262 239 328 255
rect 380 289 446 305
rect 380 255 396 289
rect 430 255 446 289
rect 380 239 446 255
rect 498 289 564 305
rect 498 255 514 289
rect 548 255 564 289
rect 498 239 564 255
rect 616 289 682 305
rect 616 255 632 289
rect 666 255 682 289
rect 616 239 682 255
rect 734 289 800 305
rect 734 255 750 289
rect 784 255 800 289
rect 734 239 800 255
rect 852 289 918 305
rect 852 255 868 289
rect 902 255 918 289
rect 852 239 918 255
rect 970 289 1036 305
rect 970 255 986 289
rect 1020 255 1036 289
rect 970 239 1036 255
rect 1088 289 1154 305
rect 1088 255 1104 289
rect 1138 255 1154 289
rect 1088 239 1154 255
rect 1206 289 1272 305
rect 1206 255 1222 289
rect 1256 255 1272 289
rect 1206 239 1272 255
rect 1324 289 1390 305
rect 1324 255 1340 289
rect 1374 255 1390 289
rect 1324 239 1390 255
rect -1390 181 -1324 197
rect -1390 147 -1374 181
rect -1340 147 -1324 181
rect -1390 131 -1324 147
rect -1272 181 -1206 197
rect -1272 147 -1256 181
rect -1222 147 -1206 181
rect -1272 131 -1206 147
rect -1154 181 -1088 197
rect -1154 147 -1138 181
rect -1104 147 -1088 181
rect -1154 131 -1088 147
rect -1036 181 -970 197
rect -1036 147 -1020 181
rect -986 147 -970 181
rect -1036 131 -970 147
rect -918 181 -852 197
rect -918 147 -902 181
rect -868 147 -852 181
rect -918 131 -852 147
rect -800 181 -734 197
rect -800 147 -784 181
rect -750 147 -734 181
rect -800 131 -734 147
rect -682 181 -616 197
rect -682 147 -666 181
rect -632 147 -616 181
rect -682 131 -616 147
rect -564 181 -498 197
rect -564 147 -548 181
rect -514 147 -498 181
rect -564 131 -498 147
rect -446 181 -380 197
rect -446 147 -430 181
rect -396 147 -380 181
rect -446 131 -380 147
rect -328 181 -262 197
rect -328 147 -312 181
rect -278 147 -262 181
rect -328 131 -262 147
rect -210 181 -144 197
rect -210 147 -194 181
rect -160 147 -144 181
rect -210 131 -144 147
rect -92 181 -26 197
rect -92 147 -76 181
rect -42 147 -26 181
rect -92 131 -26 147
rect 26 181 92 197
rect 26 147 42 181
rect 76 147 92 181
rect 26 131 92 147
rect 144 181 210 197
rect 144 147 160 181
rect 194 147 210 181
rect 144 131 210 147
rect 262 181 328 197
rect 262 147 278 181
rect 312 147 328 181
rect 262 131 328 147
rect 380 181 446 197
rect 380 147 396 181
rect 430 147 446 181
rect 380 131 446 147
rect 498 181 564 197
rect 498 147 514 181
rect 548 147 564 181
rect 498 131 564 147
rect 616 181 682 197
rect 616 147 632 181
rect 666 147 682 181
rect 616 131 682 147
rect 734 181 800 197
rect 734 147 750 181
rect 784 147 800 181
rect 734 131 800 147
rect 852 181 918 197
rect 852 147 868 181
rect 902 147 918 181
rect 852 131 918 147
rect 970 181 1036 197
rect 970 147 986 181
rect 1020 147 1036 181
rect 970 131 1036 147
rect 1088 181 1154 197
rect 1088 147 1104 181
rect 1138 147 1154 181
rect 1088 131 1154 147
rect 1206 181 1272 197
rect 1206 147 1222 181
rect 1256 147 1272 181
rect 1206 131 1272 147
rect 1324 181 1390 197
rect 1324 147 1340 181
rect 1374 147 1390 181
rect 1324 131 1390 147
rect -1387 100 -1327 131
rect -1269 100 -1209 131
rect -1151 100 -1091 131
rect -1033 100 -973 131
rect -915 100 -855 131
rect -797 100 -737 131
rect -679 100 -619 131
rect -561 100 -501 131
rect -443 100 -383 131
rect -325 100 -265 131
rect -207 100 -147 131
rect -89 100 -29 131
rect 29 100 89 131
rect 147 100 207 131
rect 265 100 325 131
rect 383 100 443 131
rect 501 100 561 131
rect 619 100 679 131
rect 737 100 797 131
rect 855 100 915 131
rect 973 100 1033 131
rect 1091 100 1151 131
rect 1209 100 1269 131
rect 1327 100 1387 131
rect -1387 -131 -1327 -100
rect -1269 -131 -1209 -100
rect -1151 -131 -1091 -100
rect -1033 -131 -973 -100
rect -915 -131 -855 -100
rect -797 -131 -737 -100
rect -679 -131 -619 -100
rect -561 -131 -501 -100
rect -443 -131 -383 -100
rect -325 -131 -265 -100
rect -207 -131 -147 -100
rect -89 -131 -29 -100
rect 29 -131 89 -100
rect 147 -131 207 -100
rect 265 -131 325 -100
rect 383 -131 443 -100
rect 501 -131 561 -100
rect 619 -131 679 -100
rect 737 -131 797 -100
rect 855 -131 915 -100
rect 973 -131 1033 -100
rect 1091 -131 1151 -100
rect 1209 -131 1269 -100
rect 1327 -131 1387 -100
rect -1390 -147 -1324 -131
rect -1390 -181 -1374 -147
rect -1340 -181 -1324 -147
rect -1390 -197 -1324 -181
rect -1272 -147 -1206 -131
rect -1272 -181 -1256 -147
rect -1222 -181 -1206 -147
rect -1272 -197 -1206 -181
rect -1154 -147 -1088 -131
rect -1154 -181 -1138 -147
rect -1104 -181 -1088 -147
rect -1154 -197 -1088 -181
rect -1036 -147 -970 -131
rect -1036 -181 -1020 -147
rect -986 -181 -970 -147
rect -1036 -197 -970 -181
rect -918 -147 -852 -131
rect -918 -181 -902 -147
rect -868 -181 -852 -147
rect -918 -197 -852 -181
rect -800 -147 -734 -131
rect -800 -181 -784 -147
rect -750 -181 -734 -147
rect -800 -197 -734 -181
rect -682 -147 -616 -131
rect -682 -181 -666 -147
rect -632 -181 -616 -147
rect -682 -197 -616 -181
rect -564 -147 -498 -131
rect -564 -181 -548 -147
rect -514 -181 -498 -147
rect -564 -197 -498 -181
rect -446 -147 -380 -131
rect -446 -181 -430 -147
rect -396 -181 -380 -147
rect -446 -197 -380 -181
rect -328 -147 -262 -131
rect -328 -181 -312 -147
rect -278 -181 -262 -147
rect -328 -197 -262 -181
rect -210 -147 -144 -131
rect -210 -181 -194 -147
rect -160 -181 -144 -147
rect -210 -197 -144 -181
rect -92 -147 -26 -131
rect -92 -181 -76 -147
rect -42 -181 -26 -147
rect -92 -197 -26 -181
rect 26 -147 92 -131
rect 26 -181 42 -147
rect 76 -181 92 -147
rect 26 -197 92 -181
rect 144 -147 210 -131
rect 144 -181 160 -147
rect 194 -181 210 -147
rect 144 -197 210 -181
rect 262 -147 328 -131
rect 262 -181 278 -147
rect 312 -181 328 -147
rect 262 -197 328 -181
rect 380 -147 446 -131
rect 380 -181 396 -147
rect 430 -181 446 -147
rect 380 -197 446 -181
rect 498 -147 564 -131
rect 498 -181 514 -147
rect 548 -181 564 -147
rect 498 -197 564 -181
rect 616 -147 682 -131
rect 616 -181 632 -147
rect 666 -181 682 -147
rect 616 -197 682 -181
rect 734 -147 800 -131
rect 734 -181 750 -147
rect 784 -181 800 -147
rect 734 -197 800 -181
rect 852 -147 918 -131
rect 852 -181 868 -147
rect 902 -181 918 -147
rect 852 -197 918 -181
rect 970 -147 1036 -131
rect 970 -181 986 -147
rect 1020 -181 1036 -147
rect 970 -197 1036 -181
rect 1088 -147 1154 -131
rect 1088 -181 1104 -147
rect 1138 -181 1154 -147
rect 1088 -197 1154 -181
rect 1206 -147 1272 -131
rect 1206 -181 1222 -147
rect 1256 -181 1272 -147
rect 1206 -197 1272 -181
rect 1324 -147 1390 -131
rect 1324 -181 1340 -147
rect 1374 -181 1390 -147
rect 1324 -197 1390 -181
rect -1390 -255 -1324 -239
rect -1390 -289 -1374 -255
rect -1340 -289 -1324 -255
rect -1390 -305 -1324 -289
rect -1272 -255 -1206 -239
rect -1272 -289 -1256 -255
rect -1222 -289 -1206 -255
rect -1272 -305 -1206 -289
rect -1154 -255 -1088 -239
rect -1154 -289 -1138 -255
rect -1104 -289 -1088 -255
rect -1154 -305 -1088 -289
rect -1036 -255 -970 -239
rect -1036 -289 -1020 -255
rect -986 -289 -970 -255
rect -1036 -305 -970 -289
rect -918 -255 -852 -239
rect -918 -289 -902 -255
rect -868 -289 -852 -255
rect -918 -305 -852 -289
rect -800 -255 -734 -239
rect -800 -289 -784 -255
rect -750 -289 -734 -255
rect -800 -305 -734 -289
rect -682 -255 -616 -239
rect -682 -289 -666 -255
rect -632 -289 -616 -255
rect -682 -305 -616 -289
rect -564 -255 -498 -239
rect -564 -289 -548 -255
rect -514 -289 -498 -255
rect -564 -305 -498 -289
rect -446 -255 -380 -239
rect -446 -289 -430 -255
rect -396 -289 -380 -255
rect -446 -305 -380 -289
rect -328 -255 -262 -239
rect -328 -289 -312 -255
rect -278 -289 -262 -255
rect -328 -305 -262 -289
rect -210 -255 -144 -239
rect -210 -289 -194 -255
rect -160 -289 -144 -255
rect -210 -305 -144 -289
rect -92 -255 -26 -239
rect -92 -289 -76 -255
rect -42 -289 -26 -255
rect -92 -305 -26 -289
rect 26 -255 92 -239
rect 26 -289 42 -255
rect 76 -289 92 -255
rect 26 -305 92 -289
rect 144 -255 210 -239
rect 144 -289 160 -255
rect 194 -289 210 -255
rect 144 -305 210 -289
rect 262 -255 328 -239
rect 262 -289 278 -255
rect 312 -289 328 -255
rect 262 -305 328 -289
rect 380 -255 446 -239
rect 380 -289 396 -255
rect 430 -289 446 -255
rect 380 -305 446 -289
rect 498 -255 564 -239
rect 498 -289 514 -255
rect 548 -289 564 -255
rect 498 -305 564 -289
rect 616 -255 682 -239
rect 616 -289 632 -255
rect 666 -289 682 -255
rect 616 -305 682 -289
rect 734 -255 800 -239
rect 734 -289 750 -255
rect 784 -289 800 -255
rect 734 -305 800 -289
rect 852 -255 918 -239
rect 852 -289 868 -255
rect 902 -289 918 -255
rect 852 -305 918 -289
rect 970 -255 1036 -239
rect 970 -289 986 -255
rect 1020 -289 1036 -255
rect 970 -305 1036 -289
rect 1088 -255 1154 -239
rect 1088 -289 1104 -255
rect 1138 -289 1154 -255
rect 1088 -305 1154 -289
rect 1206 -255 1272 -239
rect 1206 -289 1222 -255
rect 1256 -289 1272 -255
rect 1206 -305 1272 -289
rect 1324 -255 1390 -239
rect 1324 -289 1340 -255
rect 1374 -289 1390 -255
rect 1324 -305 1390 -289
rect -1387 -336 -1327 -305
rect -1269 -336 -1209 -305
rect -1151 -336 -1091 -305
rect -1033 -336 -973 -305
rect -915 -336 -855 -305
rect -797 -336 -737 -305
rect -679 -336 -619 -305
rect -561 -336 -501 -305
rect -443 -336 -383 -305
rect -325 -336 -265 -305
rect -207 -336 -147 -305
rect -89 -336 -29 -305
rect 29 -336 89 -305
rect 147 -336 207 -305
rect 265 -336 325 -305
rect 383 -336 443 -305
rect 501 -336 561 -305
rect 619 -336 679 -305
rect 737 -336 797 -305
rect 855 -336 915 -305
rect 973 -336 1033 -305
rect 1091 -336 1151 -305
rect 1209 -336 1269 -305
rect 1327 -336 1387 -305
rect -1387 -567 -1327 -536
rect -1269 -567 -1209 -536
rect -1151 -567 -1091 -536
rect -1033 -567 -973 -536
rect -915 -567 -855 -536
rect -797 -567 -737 -536
rect -679 -567 -619 -536
rect -561 -567 -501 -536
rect -443 -567 -383 -536
rect -325 -567 -265 -536
rect -207 -567 -147 -536
rect -89 -567 -29 -536
rect 29 -567 89 -536
rect 147 -567 207 -536
rect 265 -567 325 -536
rect 383 -567 443 -536
rect 501 -567 561 -536
rect 619 -567 679 -536
rect 737 -567 797 -536
rect 855 -567 915 -536
rect 973 -567 1033 -536
rect 1091 -567 1151 -536
rect 1209 -567 1269 -536
rect 1327 -567 1387 -536
rect -1390 -583 -1324 -567
rect -1390 -617 -1374 -583
rect -1340 -617 -1324 -583
rect -1390 -633 -1324 -617
rect -1272 -583 -1206 -567
rect -1272 -617 -1256 -583
rect -1222 -617 -1206 -583
rect -1272 -633 -1206 -617
rect -1154 -583 -1088 -567
rect -1154 -617 -1138 -583
rect -1104 -617 -1088 -583
rect -1154 -633 -1088 -617
rect -1036 -583 -970 -567
rect -1036 -617 -1020 -583
rect -986 -617 -970 -583
rect -1036 -633 -970 -617
rect -918 -583 -852 -567
rect -918 -617 -902 -583
rect -868 -617 -852 -583
rect -918 -633 -852 -617
rect -800 -583 -734 -567
rect -800 -617 -784 -583
rect -750 -617 -734 -583
rect -800 -633 -734 -617
rect -682 -583 -616 -567
rect -682 -617 -666 -583
rect -632 -617 -616 -583
rect -682 -633 -616 -617
rect -564 -583 -498 -567
rect -564 -617 -548 -583
rect -514 -617 -498 -583
rect -564 -633 -498 -617
rect -446 -583 -380 -567
rect -446 -617 -430 -583
rect -396 -617 -380 -583
rect -446 -633 -380 -617
rect -328 -583 -262 -567
rect -328 -617 -312 -583
rect -278 -617 -262 -583
rect -328 -633 -262 -617
rect -210 -583 -144 -567
rect -210 -617 -194 -583
rect -160 -617 -144 -583
rect -210 -633 -144 -617
rect -92 -583 -26 -567
rect -92 -617 -76 -583
rect -42 -617 -26 -583
rect -92 -633 -26 -617
rect 26 -583 92 -567
rect 26 -617 42 -583
rect 76 -617 92 -583
rect 26 -633 92 -617
rect 144 -583 210 -567
rect 144 -617 160 -583
rect 194 -617 210 -583
rect 144 -633 210 -617
rect 262 -583 328 -567
rect 262 -617 278 -583
rect 312 -617 328 -583
rect 262 -633 328 -617
rect 380 -583 446 -567
rect 380 -617 396 -583
rect 430 -617 446 -583
rect 380 -633 446 -617
rect 498 -583 564 -567
rect 498 -617 514 -583
rect 548 -617 564 -583
rect 498 -633 564 -617
rect 616 -583 682 -567
rect 616 -617 632 -583
rect 666 -617 682 -583
rect 616 -633 682 -617
rect 734 -583 800 -567
rect 734 -617 750 -583
rect 784 -617 800 -583
rect 734 -633 800 -617
rect 852 -583 918 -567
rect 852 -617 868 -583
rect 902 -617 918 -583
rect 852 -633 918 -617
rect 970 -583 1036 -567
rect 970 -617 986 -583
rect 1020 -617 1036 -583
rect 970 -633 1036 -617
rect 1088 -583 1154 -567
rect 1088 -617 1104 -583
rect 1138 -617 1154 -583
rect 1088 -633 1154 -617
rect 1206 -583 1272 -567
rect 1206 -617 1222 -583
rect 1256 -617 1272 -583
rect 1206 -633 1272 -617
rect 1324 -583 1390 -567
rect 1324 -617 1340 -583
rect 1374 -617 1390 -583
rect 1324 -633 1390 -617
<< polycont >>
rect -1374 583 -1340 617
rect -1256 583 -1222 617
rect -1138 583 -1104 617
rect -1020 583 -986 617
rect -902 583 -868 617
rect -784 583 -750 617
rect -666 583 -632 617
rect -548 583 -514 617
rect -430 583 -396 617
rect -312 583 -278 617
rect -194 583 -160 617
rect -76 583 -42 617
rect 42 583 76 617
rect 160 583 194 617
rect 278 583 312 617
rect 396 583 430 617
rect 514 583 548 617
rect 632 583 666 617
rect 750 583 784 617
rect 868 583 902 617
rect 986 583 1020 617
rect 1104 583 1138 617
rect 1222 583 1256 617
rect 1340 583 1374 617
rect -1374 255 -1340 289
rect -1256 255 -1222 289
rect -1138 255 -1104 289
rect -1020 255 -986 289
rect -902 255 -868 289
rect -784 255 -750 289
rect -666 255 -632 289
rect -548 255 -514 289
rect -430 255 -396 289
rect -312 255 -278 289
rect -194 255 -160 289
rect -76 255 -42 289
rect 42 255 76 289
rect 160 255 194 289
rect 278 255 312 289
rect 396 255 430 289
rect 514 255 548 289
rect 632 255 666 289
rect 750 255 784 289
rect 868 255 902 289
rect 986 255 1020 289
rect 1104 255 1138 289
rect 1222 255 1256 289
rect 1340 255 1374 289
rect -1374 147 -1340 181
rect -1256 147 -1222 181
rect -1138 147 -1104 181
rect -1020 147 -986 181
rect -902 147 -868 181
rect -784 147 -750 181
rect -666 147 -632 181
rect -548 147 -514 181
rect -430 147 -396 181
rect -312 147 -278 181
rect -194 147 -160 181
rect -76 147 -42 181
rect 42 147 76 181
rect 160 147 194 181
rect 278 147 312 181
rect 396 147 430 181
rect 514 147 548 181
rect 632 147 666 181
rect 750 147 784 181
rect 868 147 902 181
rect 986 147 1020 181
rect 1104 147 1138 181
rect 1222 147 1256 181
rect 1340 147 1374 181
rect -1374 -181 -1340 -147
rect -1256 -181 -1222 -147
rect -1138 -181 -1104 -147
rect -1020 -181 -986 -147
rect -902 -181 -868 -147
rect -784 -181 -750 -147
rect -666 -181 -632 -147
rect -548 -181 -514 -147
rect -430 -181 -396 -147
rect -312 -181 -278 -147
rect -194 -181 -160 -147
rect -76 -181 -42 -147
rect 42 -181 76 -147
rect 160 -181 194 -147
rect 278 -181 312 -147
rect 396 -181 430 -147
rect 514 -181 548 -147
rect 632 -181 666 -147
rect 750 -181 784 -147
rect 868 -181 902 -147
rect 986 -181 1020 -147
rect 1104 -181 1138 -147
rect 1222 -181 1256 -147
rect 1340 -181 1374 -147
rect -1374 -289 -1340 -255
rect -1256 -289 -1222 -255
rect -1138 -289 -1104 -255
rect -1020 -289 -986 -255
rect -902 -289 -868 -255
rect -784 -289 -750 -255
rect -666 -289 -632 -255
rect -548 -289 -514 -255
rect -430 -289 -396 -255
rect -312 -289 -278 -255
rect -194 -289 -160 -255
rect -76 -289 -42 -255
rect 42 -289 76 -255
rect 160 -289 194 -255
rect 278 -289 312 -255
rect 396 -289 430 -255
rect 514 -289 548 -255
rect 632 -289 666 -255
rect 750 -289 784 -255
rect 868 -289 902 -255
rect 986 -289 1020 -255
rect 1104 -289 1138 -255
rect 1222 -289 1256 -255
rect 1340 -289 1374 -255
rect -1374 -617 -1340 -583
rect -1256 -617 -1222 -583
rect -1138 -617 -1104 -583
rect -1020 -617 -986 -583
rect -902 -617 -868 -583
rect -784 -617 -750 -583
rect -666 -617 -632 -583
rect -548 -617 -514 -583
rect -430 -617 -396 -583
rect -312 -617 -278 -583
rect -194 -617 -160 -583
rect -76 -617 -42 -583
rect 42 -617 76 -583
rect 160 -617 194 -583
rect 278 -617 312 -583
rect 396 -617 430 -583
rect 514 -617 548 -583
rect 632 -617 666 -583
rect 750 -617 784 -583
rect 868 -617 902 -583
rect 986 -617 1020 -583
rect 1104 -617 1138 -583
rect 1222 -617 1256 -583
rect 1340 -617 1374 -583
<< locali >>
rect -1547 685 -1451 719
rect 1451 685 1547 719
rect -1547 623 -1513 685
rect 1513 623 1547 685
rect -1390 583 -1374 617
rect -1340 583 -1324 617
rect -1272 583 -1256 617
rect -1222 583 -1206 617
rect -1154 583 -1138 617
rect -1104 583 -1088 617
rect -1036 583 -1020 617
rect -986 583 -970 617
rect -918 583 -902 617
rect -868 583 -852 617
rect -800 583 -784 617
rect -750 583 -734 617
rect -682 583 -666 617
rect -632 583 -616 617
rect -564 583 -548 617
rect -514 583 -498 617
rect -446 583 -430 617
rect -396 583 -380 617
rect -328 583 -312 617
rect -278 583 -262 617
rect -210 583 -194 617
rect -160 583 -144 617
rect -92 583 -76 617
rect -42 583 -26 617
rect 26 583 42 617
rect 76 583 92 617
rect 144 583 160 617
rect 194 583 210 617
rect 262 583 278 617
rect 312 583 328 617
rect 380 583 396 617
rect 430 583 446 617
rect 498 583 514 617
rect 548 583 564 617
rect 616 583 632 617
rect 666 583 682 617
rect 734 583 750 617
rect 784 583 800 617
rect 852 583 868 617
rect 902 583 918 617
rect 970 583 986 617
rect 1020 583 1036 617
rect 1088 583 1104 617
rect 1138 583 1154 617
rect 1206 583 1222 617
rect 1256 583 1272 617
rect 1324 583 1340 617
rect 1374 583 1390 617
rect -1433 524 -1399 540
rect -1433 332 -1399 348
rect -1315 524 -1281 540
rect -1315 332 -1281 348
rect -1197 524 -1163 540
rect -1197 332 -1163 348
rect -1079 524 -1045 540
rect -1079 332 -1045 348
rect -961 524 -927 540
rect -961 332 -927 348
rect -843 524 -809 540
rect -843 332 -809 348
rect -725 524 -691 540
rect -725 332 -691 348
rect -607 524 -573 540
rect -607 332 -573 348
rect -489 524 -455 540
rect -489 332 -455 348
rect -371 524 -337 540
rect -371 332 -337 348
rect -253 524 -219 540
rect -253 332 -219 348
rect -135 524 -101 540
rect -135 332 -101 348
rect -17 524 17 540
rect -17 332 17 348
rect 101 524 135 540
rect 101 332 135 348
rect 219 524 253 540
rect 219 332 253 348
rect 337 524 371 540
rect 337 332 371 348
rect 455 524 489 540
rect 455 332 489 348
rect 573 524 607 540
rect 573 332 607 348
rect 691 524 725 540
rect 691 332 725 348
rect 809 524 843 540
rect 809 332 843 348
rect 927 524 961 540
rect 927 332 961 348
rect 1045 524 1079 540
rect 1045 332 1079 348
rect 1163 524 1197 540
rect 1163 332 1197 348
rect 1281 524 1315 540
rect 1281 332 1315 348
rect 1399 524 1433 540
rect 1399 332 1433 348
rect -1390 255 -1374 289
rect -1340 255 -1324 289
rect -1272 255 -1256 289
rect -1222 255 -1206 289
rect -1154 255 -1138 289
rect -1104 255 -1088 289
rect -1036 255 -1020 289
rect -986 255 -970 289
rect -918 255 -902 289
rect -868 255 -852 289
rect -800 255 -784 289
rect -750 255 -734 289
rect -682 255 -666 289
rect -632 255 -616 289
rect -564 255 -548 289
rect -514 255 -498 289
rect -446 255 -430 289
rect -396 255 -380 289
rect -328 255 -312 289
rect -278 255 -262 289
rect -210 255 -194 289
rect -160 255 -144 289
rect -92 255 -76 289
rect -42 255 -26 289
rect 26 255 42 289
rect 76 255 92 289
rect 144 255 160 289
rect 194 255 210 289
rect 262 255 278 289
rect 312 255 328 289
rect 380 255 396 289
rect 430 255 446 289
rect 498 255 514 289
rect 548 255 564 289
rect 616 255 632 289
rect 666 255 682 289
rect 734 255 750 289
rect 784 255 800 289
rect 852 255 868 289
rect 902 255 918 289
rect 970 255 986 289
rect 1020 255 1036 289
rect 1088 255 1104 289
rect 1138 255 1154 289
rect 1206 255 1222 289
rect 1256 255 1272 289
rect 1324 255 1340 289
rect 1374 255 1390 289
rect -1390 147 -1374 181
rect -1340 147 -1324 181
rect -1272 147 -1256 181
rect -1222 147 -1206 181
rect -1154 147 -1138 181
rect -1104 147 -1088 181
rect -1036 147 -1020 181
rect -986 147 -970 181
rect -918 147 -902 181
rect -868 147 -852 181
rect -800 147 -784 181
rect -750 147 -734 181
rect -682 147 -666 181
rect -632 147 -616 181
rect -564 147 -548 181
rect -514 147 -498 181
rect -446 147 -430 181
rect -396 147 -380 181
rect -328 147 -312 181
rect -278 147 -262 181
rect -210 147 -194 181
rect -160 147 -144 181
rect -92 147 -76 181
rect -42 147 -26 181
rect 26 147 42 181
rect 76 147 92 181
rect 144 147 160 181
rect 194 147 210 181
rect 262 147 278 181
rect 312 147 328 181
rect 380 147 396 181
rect 430 147 446 181
rect 498 147 514 181
rect 548 147 564 181
rect 616 147 632 181
rect 666 147 682 181
rect 734 147 750 181
rect 784 147 800 181
rect 852 147 868 181
rect 902 147 918 181
rect 970 147 986 181
rect 1020 147 1036 181
rect 1088 147 1104 181
rect 1138 147 1154 181
rect 1206 147 1222 181
rect 1256 147 1272 181
rect 1324 147 1340 181
rect 1374 147 1390 181
rect -1433 88 -1399 104
rect -1433 -104 -1399 -88
rect -1315 88 -1281 104
rect -1315 -104 -1281 -88
rect -1197 88 -1163 104
rect -1197 -104 -1163 -88
rect -1079 88 -1045 104
rect -1079 -104 -1045 -88
rect -961 88 -927 104
rect -961 -104 -927 -88
rect -843 88 -809 104
rect -843 -104 -809 -88
rect -725 88 -691 104
rect -725 -104 -691 -88
rect -607 88 -573 104
rect -607 -104 -573 -88
rect -489 88 -455 104
rect -489 -104 -455 -88
rect -371 88 -337 104
rect -371 -104 -337 -88
rect -253 88 -219 104
rect -253 -104 -219 -88
rect -135 88 -101 104
rect -135 -104 -101 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 101 88 135 104
rect 101 -104 135 -88
rect 219 88 253 104
rect 219 -104 253 -88
rect 337 88 371 104
rect 337 -104 371 -88
rect 455 88 489 104
rect 455 -104 489 -88
rect 573 88 607 104
rect 573 -104 607 -88
rect 691 88 725 104
rect 691 -104 725 -88
rect 809 88 843 104
rect 809 -104 843 -88
rect 927 88 961 104
rect 927 -104 961 -88
rect 1045 88 1079 104
rect 1045 -104 1079 -88
rect 1163 88 1197 104
rect 1163 -104 1197 -88
rect 1281 88 1315 104
rect 1281 -104 1315 -88
rect 1399 88 1433 104
rect 1399 -104 1433 -88
rect -1390 -181 -1374 -147
rect -1340 -181 -1324 -147
rect -1272 -181 -1256 -147
rect -1222 -181 -1206 -147
rect -1154 -181 -1138 -147
rect -1104 -181 -1088 -147
rect -1036 -181 -1020 -147
rect -986 -181 -970 -147
rect -918 -181 -902 -147
rect -868 -181 -852 -147
rect -800 -181 -784 -147
rect -750 -181 -734 -147
rect -682 -181 -666 -147
rect -632 -181 -616 -147
rect -564 -181 -548 -147
rect -514 -181 -498 -147
rect -446 -181 -430 -147
rect -396 -181 -380 -147
rect -328 -181 -312 -147
rect -278 -181 -262 -147
rect -210 -181 -194 -147
rect -160 -181 -144 -147
rect -92 -181 -76 -147
rect -42 -181 -26 -147
rect 26 -181 42 -147
rect 76 -181 92 -147
rect 144 -181 160 -147
rect 194 -181 210 -147
rect 262 -181 278 -147
rect 312 -181 328 -147
rect 380 -181 396 -147
rect 430 -181 446 -147
rect 498 -181 514 -147
rect 548 -181 564 -147
rect 616 -181 632 -147
rect 666 -181 682 -147
rect 734 -181 750 -147
rect 784 -181 800 -147
rect 852 -181 868 -147
rect 902 -181 918 -147
rect 970 -181 986 -147
rect 1020 -181 1036 -147
rect 1088 -181 1104 -147
rect 1138 -181 1154 -147
rect 1206 -181 1222 -147
rect 1256 -181 1272 -147
rect 1324 -181 1340 -147
rect 1374 -181 1390 -147
rect -1390 -289 -1374 -255
rect -1340 -289 -1324 -255
rect -1272 -289 -1256 -255
rect -1222 -289 -1206 -255
rect -1154 -289 -1138 -255
rect -1104 -289 -1088 -255
rect -1036 -289 -1020 -255
rect -986 -289 -970 -255
rect -918 -289 -902 -255
rect -868 -289 -852 -255
rect -800 -289 -784 -255
rect -750 -289 -734 -255
rect -682 -289 -666 -255
rect -632 -289 -616 -255
rect -564 -289 -548 -255
rect -514 -289 -498 -255
rect -446 -289 -430 -255
rect -396 -289 -380 -255
rect -328 -289 -312 -255
rect -278 -289 -262 -255
rect -210 -289 -194 -255
rect -160 -289 -144 -255
rect -92 -289 -76 -255
rect -42 -289 -26 -255
rect 26 -289 42 -255
rect 76 -289 92 -255
rect 144 -289 160 -255
rect 194 -289 210 -255
rect 262 -289 278 -255
rect 312 -289 328 -255
rect 380 -289 396 -255
rect 430 -289 446 -255
rect 498 -289 514 -255
rect 548 -289 564 -255
rect 616 -289 632 -255
rect 666 -289 682 -255
rect 734 -289 750 -255
rect 784 -289 800 -255
rect 852 -289 868 -255
rect 902 -289 918 -255
rect 970 -289 986 -255
rect 1020 -289 1036 -255
rect 1088 -289 1104 -255
rect 1138 -289 1154 -255
rect 1206 -289 1222 -255
rect 1256 -289 1272 -255
rect 1324 -289 1340 -255
rect 1374 -289 1390 -255
rect -1433 -348 -1399 -332
rect -1433 -540 -1399 -524
rect -1315 -348 -1281 -332
rect -1315 -540 -1281 -524
rect -1197 -348 -1163 -332
rect -1197 -540 -1163 -524
rect -1079 -348 -1045 -332
rect -1079 -540 -1045 -524
rect -961 -348 -927 -332
rect -961 -540 -927 -524
rect -843 -348 -809 -332
rect -843 -540 -809 -524
rect -725 -348 -691 -332
rect -725 -540 -691 -524
rect -607 -348 -573 -332
rect -607 -540 -573 -524
rect -489 -348 -455 -332
rect -489 -540 -455 -524
rect -371 -348 -337 -332
rect -371 -540 -337 -524
rect -253 -348 -219 -332
rect -253 -540 -219 -524
rect -135 -348 -101 -332
rect -135 -540 -101 -524
rect -17 -348 17 -332
rect -17 -540 17 -524
rect 101 -348 135 -332
rect 101 -540 135 -524
rect 219 -348 253 -332
rect 219 -540 253 -524
rect 337 -348 371 -332
rect 337 -540 371 -524
rect 455 -348 489 -332
rect 455 -540 489 -524
rect 573 -348 607 -332
rect 573 -540 607 -524
rect 691 -348 725 -332
rect 691 -540 725 -524
rect 809 -348 843 -332
rect 809 -540 843 -524
rect 927 -348 961 -332
rect 927 -540 961 -524
rect 1045 -348 1079 -332
rect 1045 -540 1079 -524
rect 1163 -348 1197 -332
rect 1163 -540 1197 -524
rect 1281 -348 1315 -332
rect 1281 -540 1315 -524
rect 1399 -348 1433 -332
rect 1399 -540 1433 -524
rect -1390 -617 -1374 -583
rect -1340 -617 -1324 -583
rect -1272 -617 -1256 -583
rect -1222 -617 -1206 -583
rect -1154 -617 -1138 -583
rect -1104 -617 -1088 -583
rect -1036 -617 -1020 -583
rect -986 -617 -970 -583
rect -918 -617 -902 -583
rect -868 -617 -852 -583
rect -800 -617 -784 -583
rect -750 -617 -734 -583
rect -682 -617 -666 -583
rect -632 -617 -616 -583
rect -564 -617 -548 -583
rect -514 -617 -498 -583
rect -446 -617 -430 -583
rect -396 -617 -380 -583
rect -328 -617 -312 -583
rect -278 -617 -262 -583
rect -210 -617 -194 -583
rect -160 -617 -144 -583
rect -92 -617 -76 -583
rect -42 -617 -26 -583
rect 26 -617 42 -583
rect 76 -617 92 -583
rect 144 -617 160 -583
rect 194 -617 210 -583
rect 262 -617 278 -583
rect 312 -617 328 -583
rect 380 -617 396 -583
rect 430 -617 446 -583
rect 498 -617 514 -583
rect 548 -617 564 -583
rect 616 -617 632 -583
rect 666 -617 682 -583
rect 734 -617 750 -583
rect 784 -617 800 -583
rect 852 -617 868 -583
rect 902 -617 918 -583
rect 970 -617 986 -583
rect 1020 -617 1036 -583
rect 1088 -617 1104 -583
rect 1138 -617 1154 -583
rect 1206 -617 1222 -583
rect 1256 -617 1272 -583
rect 1324 -617 1340 -583
rect 1374 -617 1390 -583
rect -1547 -685 -1513 -623
rect 1513 -685 1547 -623
rect -1547 -719 -1451 -685
rect 1451 -719 1547 -685
<< viali >>
rect -1374 583 -1340 617
rect -1256 583 -1222 617
rect -1138 583 -1104 617
rect -1020 583 -986 617
rect -902 583 -868 617
rect -784 583 -750 617
rect -666 583 -632 617
rect -548 583 -514 617
rect -430 583 -396 617
rect -312 583 -278 617
rect -194 583 -160 617
rect -76 583 -42 617
rect 42 583 76 617
rect 160 583 194 617
rect 278 583 312 617
rect 396 583 430 617
rect 514 583 548 617
rect 632 583 666 617
rect 750 583 784 617
rect 868 583 902 617
rect 986 583 1020 617
rect 1104 583 1138 617
rect 1222 583 1256 617
rect 1340 583 1374 617
rect -1433 348 -1399 524
rect -1315 348 -1281 524
rect -1197 348 -1163 524
rect -1079 348 -1045 524
rect -961 348 -927 524
rect -843 348 -809 524
rect -725 348 -691 524
rect -607 348 -573 524
rect -489 348 -455 524
rect -371 348 -337 524
rect -253 348 -219 524
rect -135 348 -101 524
rect -17 348 17 524
rect 101 348 135 524
rect 219 348 253 524
rect 337 348 371 524
rect 455 348 489 524
rect 573 348 607 524
rect 691 348 725 524
rect 809 348 843 524
rect 927 348 961 524
rect 1045 348 1079 524
rect 1163 348 1197 524
rect 1281 348 1315 524
rect 1399 348 1433 524
rect -1374 255 -1340 289
rect -1256 255 -1222 289
rect -1138 255 -1104 289
rect -1020 255 -986 289
rect -902 255 -868 289
rect -784 255 -750 289
rect -666 255 -632 289
rect -548 255 -514 289
rect -430 255 -396 289
rect -312 255 -278 289
rect -194 255 -160 289
rect -76 255 -42 289
rect 42 255 76 289
rect 160 255 194 289
rect 278 255 312 289
rect 396 255 430 289
rect 514 255 548 289
rect 632 255 666 289
rect 750 255 784 289
rect 868 255 902 289
rect 986 255 1020 289
rect 1104 255 1138 289
rect 1222 255 1256 289
rect 1340 255 1374 289
rect -1374 147 -1340 181
rect -1256 147 -1222 181
rect -1138 147 -1104 181
rect -1020 147 -986 181
rect -902 147 -868 181
rect -784 147 -750 181
rect -666 147 -632 181
rect -548 147 -514 181
rect -430 147 -396 181
rect -312 147 -278 181
rect -194 147 -160 181
rect -76 147 -42 181
rect 42 147 76 181
rect 160 147 194 181
rect 278 147 312 181
rect 396 147 430 181
rect 514 147 548 181
rect 632 147 666 181
rect 750 147 784 181
rect 868 147 902 181
rect 986 147 1020 181
rect 1104 147 1138 181
rect 1222 147 1256 181
rect 1340 147 1374 181
rect -1433 -88 -1399 88
rect -1315 -88 -1281 88
rect -1197 -88 -1163 88
rect -1079 -88 -1045 88
rect -961 -88 -927 88
rect -843 -88 -809 88
rect -725 -88 -691 88
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
rect 691 -88 725 88
rect 809 -88 843 88
rect 927 -88 961 88
rect 1045 -88 1079 88
rect 1163 -88 1197 88
rect 1281 -88 1315 88
rect 1399 -88 1433 88
rect -1374 -181 -1340 -147
rect -1256 -181 -1222 -147
rect -1138 -181 -1104 -147
rect -1020 -181 -986 -147
rect -902 -181 -868 -147
rect -784 -181 -750 -147
rect -666 -181 -632 -147
rect -548 -181 -514 -147
rect -430 -181 -396 -147
rect -312 -181 -278 -147
rect -194 -181 -160 -147
rect -76 -181 -42 -147
rect 42 -181 76 -147
rect 160 -181 194 -147
rect 278 -181 312 -147
rect 396 -181 430 -147
rect 514 -181 548 -147
rect 632 -181 666 -147
rect 750 -181 784 -147
rect 868 -181 902 -147
rect 986 -181 1020 -147
rect 1104 -181 1138 -147
rect 1222 -181 1256 -147
rect 1340 -181 1374 -147
rect -1374 -289 -1340 -255
rect -1256 -289 -1222 -255
rect -1138 -289 -1104 -255
rect -1020 -289 -986 -255
rect -902 -289 -868 -255
rect -784 -289 -750 -255
rect -666 -289 -632 -255
rect -548 -289 -514 -255
rect -430 -289 -396 -255
rect -312 -289 -278 -255
rect -194 -289 -160 -255
rect -76 -289 -42 -255
rect 42 -289 76 -255
rect 160 -289 194 -255
rect 278 -289 312 -255
rect 396 -289 430 -255
rect 514 -289 548 -255
rect 632 -289 666 -255
rect 750 -289 784 -255
rect 868 -289 902 -255
rect 986 -289 1020 -255
rect 1104 -289 1138 -255
rect 1222 -289 1256 -255
rect 1340 -289 1374 -255
rect -1433 -524 -1399 -348
rect -1315 -524 -1281 -348
rect -1197 -524 -1163 -348
rect -1079 -524 -1045 -348
rect -961 -524 -927 -348
rect -843 -524 -809 -348
rect -725 -524 -691 -348
rect -607 -524 -573 -348
rect -489 -524 -455 -348
rect -371 -524 -337 -348
rect -253 -524 -219 -348
rect -135 -524 -101 -348
rect -17 -524 17 -348
rect 101 -524 135 -348
rect 219 -524 253 -348
rect 337 -524 371 -348
rect 455 -524 489 -348
rect 573 -524 607 -348
rect 691 -524 725 -348
rect 809 -524 843 -348
rect 927 -524 961 -348
rect 1045 -524 1079 -348
rect 1163 -524 1197 -348
rect 1281 -524 1315 -348
rect 1399 -524 1433 -348
rect -1374 -617 -1340 -583
rect -1256 -617 -1222 -583
rect -1138 -617 -1104 -583
rect -1020 -617 -986 -583
rect -902 -617 -868 -583
rect -784 -617 -750 -583
rect -666 -617 -632 -583
rect -548 -617 -514 -583
rect -430 -617 -396 -583
rect -312 -617 -278 -583
rect -194 -617 -160 -583
rect -76 -617 -42 -583
rect 42 -617 76 -583
rect 160 -617 194 -583
rect 278 -617 312 -583
rect 396 -617 430 -583
rect 514 -617 548 -583
rect 632 -617 666 -583
rect 750 -617 784 -583
rect 868 -617 902 -583
rect 986 -617 1020 -583
rect 1104 -617 1138 -583
rect 1222 -617 1256 -583
rect 1340 -617 1374 -583
<< metal1 >>
rect -1386 617 -1328 623
rect -1386 583 -1374 617
rect -1340 583 -1328 617
rect -1386 577 -1328 583
rect -1268 617 -1210 623
rect -1268 583 -1256 617
rect -1222 583 -1210 617
rect -1268 577 -1210 583
rect -1150 617 -1092 623
rect -1150 583 -1138 617
rect -1104 583 -1092 617
rect -1150 577 -1092 583
rect -1032 617 -974 623
rect -1032 583 -1020 617
rect -986 583 -974 617
rect -1032 577 -974 583
rect -914 617 -856 623
rect -914 583 -902 617
rect -868 583 -856 617
rect -914 577 -856 583
rect -796 617 -738 623
rect -796 583 -784 617
rect -750 583 -738 617
rect -796 577 -738 583
rect -678 617 -620 623
rect -678 583 -666 617
rect -632 583 -620 617
rect -678 577 -620 583
rect -560 617 -502 623
rect -560 583 -548 617
rect -514 583 -502 617
rect -560 577 -502 583
rect -442 617 -384 623
rect -442 583 -430 617
rect -396 583 -384 617
rect -442 577 -384 583
rect -324 617 -266 623
rect -324 583 -312 617
rect -278 583 -266 617
rect -324 577 -266 583
rect -206 617 -148 623
rect -206 583 -194 617
rect -160 583 -148 617
rect -206 577 -148 583
rect -88 617 -30 623
rect -88 583 -76 617
rect -42 583 -30 617
rect -88 577 -30 583
rect 30 617 88 623
rect 30 583 42 617
rect 76 583 88 617
rect 30 577 88 583
rect 148 617 206 623
rect 148 583 160 617
rect 194 583 206 617
rect 148 577 206 583
rect 266 617 324 623
rect 266 583 278 617
rect 312 583 324 617
rect 266 577 324 583
rect 384 617 442 623
rect 384 583 396 617
rect 430 583 442 617
rect 384 577 442 583
rect 502 617 560 623
rect 502 583 514 617
rect 548 583 560 617
rect 502 577 560 583
rect 620 617 678 623
rect 620 583 632 617
rect 666 583 678 617
rect 620 577 678 583
rect 738 617 796 623
rect 738 583 750 617
rect 784 583 796 617
rect 738 577 796 583
rect 856 617 914 623
rect 856 583 868 617
rect 902 583 914 617
rect 856 577 914 583
rect 974 617 1032 623
rect 974 583 986 617
rect 1020 583 1032 617
rect 974 577 1032 583
rect 1092 617 1150 623
rect 1092 583 1104 617
rect 1138 583 1150 617
rect 1092 577 1150 583
rect 1210 617 1268 623
rect 1210 583 1222 617
rect 1256 583 1268 617
rect 1210 577 1268 583
rect 1328 617 1386 623
rect 1328 583 1340 617
rect 1374 583 1386 617
rect 1328 577 1386 583
rect -1439 524 -1393 536
rect -1439 348 -1433 524
rect -1399 348 -1393 524
rect -1439 336 -1393 348
rect -1321 524 -1275 536
rect -1321 348 -1315 524
rect -1281 348 -1275 524
rect -1321 336 -1275 348
rect -1203 524 -1157 536
rect -1203 348 -1197 524
rect -1163 348 -1157 524
rect -1203 336 -1157 348
rect -1085 524 -1039 536
rect -1085 348 -1079 524
rect -1045 348 -1039 524
rect -1085 336 -1039 348
rect -967 524 -921 536
rect -967 348 -961 524
rect -927 348 -921 524
rect -967 336 -921 348
rect -849 524 -803 536
rect -849 348 -843 524
rect -809 348 -803 524
rect -849 336 -803 348
rect -731 524 -685 536
rect -731 348 -725 524
rect -691 348 -685 524
rect -731 336 -685 348
rect -613 524 -567 536
rect -613 348 -607 524
rect -573 348 -567 524
rect -613 336 -567 348
rect -495 524 -449 536
rect -495 348 -489 524
rect -455 348 -449 524
rect -495 336 -449 348
rect -377 524 -331 536
rect -377 348 -371 524
rect -337 348 -331 524
rect -377 336 -331 348
rect -259 524 -213 536
rect -259 348 -253 524
rect -219 348 -213 524
rect -259 336 -213 348
rect -141 524 -95 536
rect -141 348 -135 524
rect -101 348 -95 524
rect -141 336 -95 348
rect -23 524 23 536
rect -23 348 -17 524
rect 17 348 23 524
rect -23 336 23 348
rect 95 524 141 536
rect 95 348 101 524
rect 135 348 141 524
rect 95 336 141 348
rect 213 524 259 536
rect 213 348 219 524
rect 253 348 259 524
rect 213 336 259 348
rect 331 524 377 536
rect 331 348 337 524
rect 371 348 377 524
rect 331 336 377 348
rect 449 524 495 536
rect 449 348 455 524
rect 489 348 495 524
rect 449 336 495 348
rect 567 524 613 536
rect 567 348 573 524
rect 607 348 613 524
rect 567 336 613 348
rect 685 524 731 536
rect 685 348 691 524
rect 725 348 731 524
rect 685 336 731 348
rect 803 524 849 536
rect 803 348 809 524
rect 843 348 849 524
rect 803 336 849 348
rect 921 524 967 536
rect 921 348 927 524
rect 961 348 967 524
rect 921 336 967 348
rect 1039 524 1085 536
rect 1039 348 1045 524
rect 1079 348 1085 524
rect 1039 336 1085 348
rect 1157 524 1203 536
rect 1157 348 1163 524
rect 1197 348 1203 524
rect 1157 336 1203 348
rect 1275 524 1321 536
rect 1275 348 1281 524
rect 1315 348 1321 524
rect 1275 336 1321 348
rect 1393 524 1439 536
rect 1393 348 1399 524
rect 1433 348 1439 524
rect 1393 336 1439 348
rect -1386 289 -1328 295
rect -1386 255 -1374 289
rect -1340 255 -1328 289
rect -1386 249 -1328 255
rect -1268 289 -1210 295
rect -1268 255 -1256 289
rect -1222 255 -1210 289
rect -1268 249 -1210 255
rect -1150 289 -1092 295
rect -1150 255 -1138 289
rect -1104 255 -1092 289
rect -1150 249 -1092 255
rect -1032 289 -974 295
rect -1032 255 -1020 289
rect -986 255 -974 289
rect -1032 249 -974 255
rect -914 289 -856 295
rect -914 255 -902 289
rect -868 255 -856 289
rect -914 249 -856 255
rect -796 289 -738 295
rect -796 255 -784 289
rect -750 255 -738 289
rect -796 249 -738 255
rect -678 289 -620 295
rect -678 255 -666 289
rect -632 255 -620 289
rect -678 249 -620 255
rect -560 289 -502 295
rect -560 255 -548 289
rect -514 255 -502 289
rect -560 249 -502 255
rect -442 289 -384 295
rect -442 255 -430 289
rect -396 255 -384 289
rect -442 249 -384 255
rect -324 289 -266 295
rect -324 255 -312 289
rect -278 255 -266 289
rect -324 249 -266 255
rect -206 289 -148 295
rect -206 255 -194 289
rect -160 255 -148 289
rect -206 249 -148 255
rect -88 289 -30 295
rect -88 255 -76 289
rect -42 255 -30 289
rect -88 249 -30 255
rect 30 289 88 295
rect 30 255 42 289
rect 76 255 88 289
rect 30 249 88 255
rect 148 289 206 295
rect 148 255 160 289
rect 194 255 206 289
rect 148 249 206 255
rect 266 289 324 295
rect 266 255 278 289
rect 312 255 324 289
rect 266 249 324 255
rect 384 289 442 295
rect 384 255 396 289
rect 430 255 442 289
rect 384 249 442 255
rect 502 289 560 295
rect 502 255 514 289
rect 548 255 560 289
rect 502 249 560 255
rect 620 289 678 295
rect 620 255 632 289
rect 666 255 678 289
rect 620 249 678 255
rect 738 289 796 295
rect 738 255 750 289
rect 784 255 796 289
rect 738 249 796 255
rect 856 289 914 295
rect 856 255 868 289
rect 902 255 914 289
rect 856 249 914 255
rect 974 289 1032 295
rect 974 255 986 289
rect 1020 255 1032 289
rect 974 249 1032 255
rect 1092 289 1150 295
rect 1092 255 1104 289
rect 1138 255 1150 289
rect 1092 249 1150 255
rect 1210 289 1268 295
rect 1210 255 1222 289
rect 1256 255 1268 289
rect 1210 249 1268 255
rect 1328 289 1386 295
rect 1328 255 1340 289
rect 1374 255 1386 289
rect 1328 249 1386 255
rect -1386 181 -1328 187
rect -1386 147 -1374 181
rect -1340 147 -1328 181
rect -1386 141 -1328 147
rect -1268 181 -1210 187
rect -1268 147 -1256 181
rect -1222 147 -1210 181
rect -1268 141 -1210 147
rect -1150 181 -1092 187
rect -1150 147 -1138 181
rect -1104 147 -1092 181
rect -1150 141 -1092 147
rect -1032 181 -974 187
rect -1032 147 -1020 181
rect -986 147 -974 181
rect -1032 141 -974 147
rect -914 181 -856 187
rect -914 147 -902 181
rect -868 147 -856 181
rect -914 141 -856 147
rect -796 181 -738 187
rect -796 147 -784 181
rect -750 147 -738 181
rect -796 141 -738 147
rect -678 181 -620 187
rect -678 147 -666 181
rect -632 147 -620 181
rect -678 141 -620 147
rect -560 181 -502 187
rect -560 147 -548 181
rect -514 147 -502 181
rect -560 141 -502 147
rect -442 181 -384 187
rect -442 147 -430 181
rect -396 147 -384 181
rect -442 141 -384 147
rect -324 181 -266 187
rect -324 147 -312 181
rect -278 147 -266 181
rect -324 141 -266 147
rect -206 181 -148 187
rect -206 147 -194 181
rect -160 147 -148 181
rect -206 141 -148 147
rect -88 181 -30 187
rect -88 147 -76 181
rect -42 147 -30 181
rect -88 141 -30 147
rect 30 181 88 187
rect 30 147 42 181
rect 76 147 88 181
rect 30 141 88 147
rect 148 181 206 187
rect 148 147 160 181
rect 194 147 206 181
rect 148 141 206 147
rect 266 181 324 187
rect 266 147 278 181
rect 312 147 324 181
rect 266 141 324 147
rect 384 181 442 187
rect 384 147 396 181
rect 430 147 442 181
rect 384 141 442 147
rect 502 181 560 187
rect 502 147 514 181
rect 548 147 560 181
rect 502 141 560 147
rect 620 181 678 187
rect 620 147 632 181
rect 666 147 678 181
rect 620 141 678 147
rect 738 181 796 187
rect 738 147 750 181
rect 784 147 796 181
rect 738 141 796 147
rect 856 181 914 187
rect 856 147 868 181
rect 902 147 914 181
rect 856 141 914 147
rect 974 181 1032 187
rect 974 147 986 181
rect 1020 147 1032 181
rect 974 141 1032 147
rect 1092 181 1150 187
rect 1092 147 1104 181
rect 1138 147 1150 181
rect 1092 141 1150 147
rect 1210 181 1268 187
rect 1210 147 1222 181
rect 1256 147 1268 181
rect 1210 141 1268 147
rect 1328 181 1386 187
rect 1328 147 1340 181
rect 1374 147 1386 181
rect 1328 141 1386 147
rect -1439 88 -1393 100
rect -1439 -88 -1433 88
rect -1399 -88 -1393 88
rect -1439 -100 -1393 -88
rect -1321 88 -1275 100
rect -1321 -88 -1315 88
rect -1281 -88 -1275 88
rect -1321 -100 -1275 -88
rect -1203 88 -1157 100
rect -1203 -88 -1197 88
rect -1163 -88 -1157 88
rect -1203 -100 -1157 -88
rect -1085 88 -1039 100
rect -1085 -88 -1079 88
rect -1045 -88 -1039 88
rect -1085 -100 -1039 -88
rect -967 88 -921 100
rect -967 -88 -961 88
rect -927 -88 -921 88
rect -967 -100 -921 -88
rect -849 88 -803 100
rect -849 -88 -843 88
rect -809 -88 -803 88
rect -849 -100 -803 -88
rect -731 88 -685 100
rect -731 -88 -725 88
rect -691 -88 -685 88
rect -731 -100 -685 -88
rect -613 88 -567 100
rect -613 -88 -607 88
rect -573 -88 -567 88
rect -613 -100 -567 -88
rect -495 88 -449 100
rect -495 -88 -489 88
rect -455 -88 -449 88
rect -495 -100 -449 -88
rect -377 88 -331 100
rect -377 -88 -371 88
rect -337 -88 -331 88
rect -377 -100 -331 -88
rect -259 88 -213 100
rect -259 -88 -253 88
rect -219 -88 -213 88
rect -259 -100 -213 -88
rect -141 88 -95 100
rect -141 -88 -135 88
rect -101 -88 -95 88
rect -141 -100 -95 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 95 88 141 100
rect 95 -88 101 88
rect 135 -88 141 88
rect 95 -100 141 -88
rect 213 88 259 100
rect 213 -88 219 88
rect 253 -88 259 88
rect 213 -100 259 -88
rect 331 88 377 100
rect 331 -88 337 88
rect 371 -88 377 88
rect 331 -100 377 -88
rect 449 88 495 100
rect 449 -88 455 88
rect 489 -88 495 88
rect 449 -100 495 -88
rect 567 88 613 100
rect 567 -88 573 88
rect 607 -88 613 88
rect 567 -100 613 -88
rect 685 88 731 100
rect 685 -88 691 88
rect 725 -88 731 88
rect 685 -100 731 -88
rect 803 88 849 100
rect 803 -88 809 88
rect 843 -88 849 88
rect 803 -100 849 -88
rect 921 88 967 100
rect 921 -88 927 88
rect 961 -88 967 88
rect 921 -100 967 -88
rect 1039 88 1085 100
rect 1039 -88 1045 88
rect 1079 -88 1085 88
rect 1039 -100 1085 -88
rect 1157 88 1203 100
rect 1157 -88 1163 88
rect 1197 -88 1203 88
rect 1157 -100 1203 -88
rect 1275 88 1321 100
rect 1275 -88 1281 88
rect 1315 -88 1321 88
rect 1275 -100 1321 -88
rect 1393 88 1439 100
rect 1393 -88 1399 88
rect 1433 -88 1439 88
rect 1393 -100 1439 -88
rect -1386 -147 -1328 -141
rect -1386 -181 -1374 -147
rect -1340 -181 -1328 -147
rect -1386 -187 -1328 -181
rect -1268 -147 -1210 -141
rect -1268 -181 -1256 -147
rect -1222 -181 -1210 -147
rect -1268 -187 -1210 -181
rect -1150 -147 -1092 -141
rect -1150 -181 -1138 -147
rect -1104 -181 -1092 -147
rect -1150 -187 -1092 -181
rect -1032 -147 -974 -141
rect -1032 -181 -1020 -147
rect -986 -181 -974 -147
rect -1032 -187 -974 -181
rect -914 -147 -856 -141
rect -914 -181 -902 -147
rect -868 -181 -856 -147
rect -914 -187 -856 -181
rect -796 -147 -738 -141
rect -796 -181 -784 -147
rect -750 -181 -738 -147
rect -796 -187 -738 -181
rect -678 -147 -620 -141
rect -678 -181 -666 -147
rect -632 -181 -620 -147
rect -678 -187 -620 -181
rect -560 -147 -502 -141
rect -560 -181 -548 -147
rect -514 -181 -502 -147
rect -560 -187 -502 -181
rect -442 -147 -384 -141
rect -442 -181 -430 -147
rect -396 -181 -384 -147
rect -442 -187 -384 -181
rect -324 -147 -266 -141
rect -324 -181 -312 -147
rect -278 -181 -266 -147
rect -324 -187 -266 -181
rect -206 -147 -148 -141
rect -206 -181 -194 -147
rect -160 -181 -148 -147
rect -206 -187 -148 -181
rect -88 -147 -30 -141
rect -88 -181 -76 -147
rect -42 -181 -30 -147
rect -88 -187 -30 -181
rect 30 -147 88 -141
rect 30 -181 42 -147
rect 76 -181 88 -147
rect 30 -187 88 -181
rect 148 -147 206 -141
rect 148 -181 160 -147
rect 194 -181 206 -147
rect 148 -187 206 -181
rect 266 -147 324 -141
rect 266 -181 278 -147
rect 312 -181 324 -147
rect 266 -187 324 -181
rect 384 -147 442 -141
rect 384 -181 396 -147
rect 430 -181 442 -147
rect 384 -187 442 -181
rect 502 -147 560 -141
rect 502 -181 514 -147
rect 548 -181 560 -147
rect 502 -187 560 -181
rect 620 -147 678 -141
rect 620 -181 632 -147
rect 666 -181 678 -147
rect 620 -187 678 -181
rect 738 -147 796 -141
rect 738 -181 750 -147
rect 784 -181 796 -147
rect 738 -187 796 -181
rect 856 -147 914 -141
rect 856 -181 868 -147
rect 902 -181 914 -147
rect 856 -187 914 -181
rect 974 -147 1032 -141
rect 974 -181 986 -147
rect 1020 -181 1032 -147
rect 974 -187 1032 -181
rect 1092 -147 1150 -141
rect 1092 -181 1104 -147
rect 1138 -181 1150 -147
rect 1092 -187 1150 -181
rect 1210 -147 1268 -141
rect 1210 -181 1222 -147
rect 1256 -181 1268 -147
rect 1210 -187 1268 -181
rect 1328 -147 1386 -141
rect 1328 -181 1340 -147
rect 1374 -181 1386 -147
rect 1328 -187 1386 -181
rect -1386 -255 -1328 -249
rect -1386 -289 -1374 -255
rect -1340 -289 -1328 -255
rect -1386 -295 -1328 -289
rect -1268 -255 -1210 -249
rect -1268 -289 -1256 -255
rect -1222 -289 -1210 -255
rect -1268 -295 -1210 -289
rect -1150 -255 -1092 -249
rect -1150 -289 -1138 -255
rect -1104 -289 -1092 -255
rect -1150 -295 -1092 -289
rect -1032 -255 -974 -249
rect -1032 -289 -1020 -255
rect -986 -289 -974 -255
rect -1032 -295 -974 -289
rect -914 -255 -856 -249
rect -914 -289 -902 -255
rect -868 -289 -856 -255
rect -914 -295 -856 -289
rect -796 -255 -738 -249
rect -796 -289 -784 -255
rect -750 -289 -738 -255
rect -796 -295 -738 -289
rect -678 -255 -620 -249
rect -678 -289 -666 -255
rect -632 -289 -620 -255
rect -678 -295 -620 -289
rect -560 -255 -502 -249
rect -560 -289 -548 -255
rect -514 -289 -502 -255
rect -560 -295 -502 -289
rect -442 -255 -384 -249
rect -442 -289 -430 -255
rect -396 -289 -384 -255
rect -442 -295 -384 -289
rect -324 -255 -266 -249
rect -324 -289 -312 -255
rect -278 -289 -266 -255
rect -324 -295 -266 -289
rect -206 -255 -148 -249
rect -206 -289 -194 -255
rect -160 -289 -148 -255
rect -206 -295 -148 -289
rect -88 -255 -30 -249
rect -88 -289 -76 -255
rect -42 -289 -30 -255
rect -88 -295 -30 -289
rect 30 -255 88 -249
rect 30 -289 42 -255
rect 76 -289 88 -255
rect 30 -295 88 -289
rect 148 -255 206 -249
rect 148 -289 160 -255
rect 194 -289 206 -255
rect 148 -295 206 -289
rect 266 -255 324 -249
rect 266 -289 278 -255
rect 312 -289 324 -255
rect 266 -295 324 -289
rect 384 -255 442 -249
rect 384 -289 396 -255
rect 430 -289 442 -255
rect 384 -295 442 -289
rect 502 -255 560 -249
rect 502 -289 514 -255
rect 548 -289 560 -255
rect 502 -295 560 -289
rect 620 -255 678 -249
rect 620 -289 632 -255
rect 666 -289 678 -255
rect 620 -295 678 -289
rect 738 -255 796 -249
rect 738 -289 750 -255
rect 784 -289 796 -255
rect 738 -295 796 -289
rect 856 -255 914 -249
rect 856 -289 868 -255
rect 902 -289 914 -255
rect 856 -295 914 -289
rect 974 -255 1032 -249
rect 974 -289 986 -255
rect 1020 -289 1032 -255
rect 974 -295 1032 -289
rect 1092 -255 1150 -249
rect 1092 -289 1104 -255
rect 1138 -289 1150 -255
rect 1092 -295 1150 -289
rect 1210 -255 1268 -249
rect 1210 -289 1222 -255
rect 1256 -289 1268 -255
rect 1210 -295 1268 -289
rect 1328 -255 1386 -249
rect 1328 -289 1340 -255
rect 1374 -289 1386 -255
rect 1328 -295 1386 -289
rect -1439 -348 -1393 -336
rect -1439 -524 -1433 -348
rect -1399 -524 -1393 -348
rect -1439 -536 -1393 -524
rect -1321 -348 -1275 -336
rect -1321 -524 -1315 -348
rect -1281 -524 -1275 -348
rect -1321 -536 -1275 -524
rect -1203 -348 -1157 -336
rect -1203 -524 -1197 -348
rect -1163 -524 -1157 -348
rect -1203 -536 -1157 -524
rect -1085 -348 -1039 -336
rect -1085 -524 -1079 -348
rect -1045 -524 -1039 -348
rect -1085 -536 -1039 -524
rect -967 -348 -921 -336
rect -967 -524 -961 -348
rect -927 -524 -921 -348
rect -967 -536 -921 -524
rect -849 -348 -803 -336
rect -849 -524 -843 -348
rect -809 -524 -803 -348
rect -849 -536 -803 -524
rect -731 -348 -685 -336
rect -731 -524 -725 -348
rect -691 -524 -685 -348
rect -731 -536 -685 -524
rect -613 -348 -567 -336
rect -613 -524 -607 -348
rect -573 -524 -567 -348
rect -613 -536 -567 -524
rect -495 -348 -449 -336
rect -495 -524 -489 -348
rect -455 -524 -449 -348
rect -495 -536 -449 -524
rect -377 -348 -331 -336
rect -377 -524 -371 -348
rect -337 -524 -331 -348
rect -377 -536 -331 -524
rect -259 -348 -213 -336
rect -259 -524 -253 -348
rect -219 -524 -213 -348
rect -259 -536 -213 -524
rect -141 -348 -95 -336
rect -141 -524 -135 -348
rect -101 -524 -95 -348
rect -141 -536 -95 -524
rect -23 -348 23 -336
rect -23 -524 -17 -348
rect 17 -524 23 -348
rect -23 -536 23 -524
rect 95 -348 141 -336
rect 95 -524 101 -348
rect 135 -524 141 -348
rect 95 -536 141 -524
rect 213 -348 259 -336
rect 213 -524 219 -348
rect 253 -524 259 -348
rect 213 -536 259 -524
rect 331 -348 377 -336
rect 331 -524 337 -348
rect 371 -524 377 -348
rect 331 -536 377 -524
rect 449 -348 495 -336
rect 449 -524 455 -348
rect 489 -524 495 -348
rect 449 -536 495 -524
rect 567 -348 613 -336
rect 567 -524 573 -348
rect 607 -524 613 -348
rect 567 -536 613 -524
rect 685 -348 731 -336
rect 685 -524 691 -348
rect 725 -524 731 -348
rect 685 -536 731 -524
rect 803 -348 849 -336
rect 803 -524 809 -348
rect 843 -524 849 -348
rect 803 -536 849 -524
rect 921 -348 967 -336
rect 921 -524 927 -348
rect 961 -524 967 -348
rect 921 -536 967 -524
rect 1039 -348 1085 -336
rect 1039 -524 1045 -348
rect 1079 -524 1085 -348
rect 1039 -536 1085 -524
rect 1157 -348 1203 -336
rect 1157 -524 1163 -348
rect 1197 -524 1203 -348
rect 1157 -536 1203 -524
rect 1275 -348 1321 -336
rect 1275 -524 1281 -348
rect 1315 -524 1321 -348
rect 1275 -536 1321 -524
rect 1393 -348 1439 -336
rect 1393 -524 1399 -348
rect 1433 -524 1439 -348
rect 1393 -536 1439 -524
rect -1386 -583 -1328 -577
rect -1386 -617 -1374 -583
rect -1340 -617 -1328 -583
rect -1386 -623 -1328 -617
rect -1268 -583 -1210 -577
rect -1268 -617 -1256 -583
rect -1222 -617 -1210 -583
rect -1268 -623 -1210 -617
rect -1150 -583 -1092 -577
rect -1150 -617 -1138 -583
rect -1104 -617 -1092 -583
rect -1150 -623 -1092 -617
rect -1032 -583 -974 -577
rect -1032 -617 -1020 -583
rect -986 -617 -974 -583
rect -1032 -623 -974 -617
rect -914 -583 -856 -577
rect -914 -617 -902 -583
rect -868 -617 -856 -583
rect -914 -623 -856 -617
rect -796 -583 -738 -577
rect -796 -617 -784 -583
rect -750 -617 -738 -583
rect -796 -623 -738 -617
rect -678 -583 -620 -577
rect -678 -617 -666 -583
rect -632 -617 -620 -583
rect -678 -623 -620 -617
rect -560 -583 -502 -577
rect -560 -617 -548 -583
rect -514 -617 -502 -583
rect -560 -623 -502 -617
rect -442 -583 -384 -577
rect -442 -617 -430 -583
rect -396 -617 -384 -583
rect -442 -623 -384 -617
rect -324 -583 -266 -577
rect -324 -617 -312 -583
rect -278 -617 -266 -583
rect -324 -623 -266 -617
rect -206 -583 -148 -577
rect -206 -617 -194 -583
rect -160 -617 -148 -583
rect -206 -623 -148 -617
rect -88 -583 -30 -577
rect -88 -617 -76 -583
rect -42 -617 -30 -583
rect -88 -623 -30 -617
rect 30 -583 88 -577
rect 30 -617 42 -583
rect 76 -617 88 -583
rect 30 -623 88 -617
rect 148 -583 206 -577
rect 148 -617 160 -583
rect 194 -617 206 -583
rect 148 -623 206 -617
rect 266 -583 324 -577
rect 266 -617 278 -583
rect 312 -617 324 -583
rect 266 -623 324 -617
rect 384 -583 442 -577
rect 384 -617 396 -583
rect 430 -617 442 -583
rect 384 -623 442 -617
rect 502 -583 560 -577
rect 502 -617 514 -583
rect 548 -617 560 -583
rect 502 -623 560 -617
rect 620 -583 678 -577
rect 620 -617 632 -583
rect 666 -617 678 -583
rect 620 -623 678 -617
rect 738 -583 796 -577
rect 738 -617 750 -583
rect 784 -617 796 -583
rect 738 -623 796 -617
rect 856 -583 914 -577
rect 856 -617 868 -583
rect 902 -617 914 -583
rect 856 -623 914 -617
rect 974 -583 1032 -577
rect 974 -617 986 -583
rect 1020 -617 1032 -583
rect 974 -623 1032 -617
rect 1092 -583 1150 -577
rect 1092 -617 1104 -583
rect 1138 -617 1150 -583
rect 1092 -623 1150 -617
rect 1210 -583 1268 -577
rect 1210 -617 1222 -583
rect 1256 -617 1268 -583
rect 1210 -623 1268 -617
rect 1328 -583 1386 -577
rect 1328 -617 1340 -583
rect 1374 -617 1386 -583
rect 1328 -623 1386 -617
<< properties >>
string FIXED_BBOX -1530 -702 1530 702
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.3 m 3 nf 24 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
