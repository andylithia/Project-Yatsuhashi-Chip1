magic
tech sky130B
timestamp 1658895968
<< metal1 >>
rect -40 1090 100 1110
rect -40 1050 0 1090
rect 60 1050 100 1090
rect -40 1030 100 1050
rect -40 990 0 1030
rect 60 990 100 1030
rect -40 970 100 990
rect -40 930 0 970
rect 60 930 100 970
rect -40 910 100 930
rect -40 870 0 910
rect 60 870 100 910
rect -40 850 100 870
rect -40 810 0 850
rect 60 810 100 850
rect -40 790 100 810
rect -40 750 0 790
rect 60 750 100 790
rect -40 730 100 750
rect -40 690 0 730
rect 60 690 100 730
rect -40 670 100 690
rect -40 630 0 670
rect 60 630 100 670
rect -40 610 100 630
rect -40 570 0 610
rect 60 570 100 610
rect -40 550 100 570
rect -40 510 0 550
rect 60 510 100 550
rect -40 490 100 510
rect -40 450 0 490
rect 60 450 100 490
rect -40 430 100 450
rect -40 390 0 430
rect 60 390 100 430
rect -40 370 100 390
rect -40 330 0 370
rect 60 330 100 370
rect -40 310 100 330
rect -40 270 0 310
rect 60 270 100 310
rect -40 250 100 270
rect -40 210 0 250
rect 60 210 100 250
rect -40 190 100 210
rect -40 150 0 190
rect 60 150 100 190
rect -40 110 100 150
rect 200 1090 340 1110
rect 200 1050 240 1090
rect 300 1050 340 1090
rect 200 1030 340 1050
rect 200 990 240 1030
rect 300 990 340 1030
rect 200 970 340 990
rect 200 930 240 970
rect 300 930 340 970
rect 200 910 340 930
rect 200 870 240 910
rect 300 870 340 910
rect 200 850 340 870
rect 200 810 240 850
rect 300 810 340 850
rect 200 790 340 810
rect 200 750 240 790
rect 300 750 340 790
rect 200 730 340 750
rect 200 690 240 730
rect 300 690 340 730
rect 200 670 340 690
rect 200 630 240 670
rect 300 630 340 670
rect 200 610 340 630
rect 200 570 240 610
rect 300 570 340 610
rect 200 550 340 570
rect 200 510 240 550
rect 300 510 340 550
rect 200 490 340 510
rect 200 450 240 490
rect 300 450 340 490
rect 200 430 340 450
rect 200 390 240 430
rect 300 390 340 430
rect 200 370 340 390
rect 200 330 240 370
rect 300 330 340 370
rect 200 310 340 330
rect 200 270 240 310
rect 300 270 340 310
rect 200 250 340 270
rect 200 210 240 250
rect 300 210 340 250
rect 200 190 340 210
rect 200 150 240 190
rect 300 150 340 190
rect 200 110 340 150
rect 440 1090 580 1110
rect 440 1050 480 1090
rect 540 1050 580 1090
rect 440 1030 580 1050
rect 440 990 480 1030
rect 540 990 580 1030
rect 440 970 580 990
rect 440 930 480 970
rect 540 930 580 970
rect 440 910 580 930
rect 440 870 480 910
rect 540 870 580 910
rect 440 850 580 870
rect 440 810 480 850
rect 540 810 580 850
rect 440 790 580 810
rect 440 750 480 790
rect 540 750 580 790
rect 440 730 580 750
rect 440 690 480 730
rect 540 690 580 730
rect 440 670 580 690
rect 440 630 480 670
rect 540 630 580 670
rect 440 610 580 630
rect 440 570 480 610
rect 540 570 580 610
rect 440 550 580 570
rect 440 510 480 550
rect 540 510 580 550
rect 440 490 580 510
rect 440 450 480 490
rect 540 450 580 490
rect 440 430 580 450
rect 440 390 480 430
rect 540 390 580 430
rect 440 370 580 390
rect 440 330 480 370
rect 540 330 580 370
rect 440 310 580 330
rect 440 270 480 310
rect 540 270 580 310
rect 440 250 580 270
rect 440 210 480 250
rect 540 210 580 250
rect 440 190 580 210
rect 440 150 480 190
rect 540 150 580 190
rect 440 110 580 150
rect 690 1090 830 1110
rect 690 1050 730 1090
rect 790 1050 830 1090
rect 690 1030 830 1050
rect 690 990 730 1030
rect 790 990 830 1030
rect 690 970 830 990
rect 690 930 730 970
rect 790 930 830 970
rect 690 910 830 930
rect 690 870 730 910
rect 790 870 830 910
rect 690 850 830 870
rect 690 810 730 850
rect 790 810 830 850
rect 690 790 830 810
rect 690 750 730 790
rect 790 750 830 790
rect 690 730 830 750
rect 690 690 730 730
rect 790 690 830 730
rect 690 670 830 690
rect 690 630 730 670
rect 790 630 830 670
rect 690 610 830 630
rect 690 570 730 610
rect 790 570 830 610
rect 690 550 830 570
rect 690 510 730 550
rect 790 510 830 550
rect 690 490 830 510
rect 690 450 730 490
rect 790 450 830 490
rect 690 430 830 450
rect 690 390 730 430
rect 790 390 830 430
rect 690 370 830 390
rect 690 330 730 370
rect 790 330 830 370
rect 690 310 830 330
rect 690 270 730 310
rect 790 270 830 310
rect 690 250 830 270
rect 690 210 730 250
rect 790 210 830 250
rect 690 190 830 210
rect 690 150 730 190
rect 790 150 830 190
rect 690 110 830 150
rect 930 1090 1070 1110
rect 930 1050 970 1090
rect 1030 1050 1070 1090
rect 930 1030 1070 1050
rect 930 990 970 1030
rect 1030 990 1070 1030
rect 930 970 1070 990
rect 930 930 970 970
rect 1030 930 1070 970
rect 930 910 1070 930
rect 930 870 970 910
rect 1030 870 1070 910
rect 930 850 1070 870
rect 930 810 970 850
rect 1030 810 1070 850
rect 930 790 1070 810
rect 930 750 970 790
rect 1030 750 1070 790
rect 930 730 1070 750
rect 930 690 970 730
rect 1030 690 1070 730
rect 930 670 1070 690
rect 930 630 970 670
rect 1030 630 1070 670
rect 930 610 1070 630
rect 930 570 970 610
rect 1030 570 1070 610
rect 930 550 1070 570
rect 930 510 970 550
rect 1030 510 1070 550
rect 930 490 1070 510
rect 930 450 970 490
rect 1030 450 1070 490
rect 930 430 1070 450
rect 930 390 970 430
rect 1030 390 1070 430
rect 930 370 1070 390
rect 930 330 970 370
rect 1030 330 1070 370
rect 930 310 1070 330
rect 930 270 970 310
rect 1030 270 1070 310
rect 930 250 1070 270
rect 930 210 970 250
rect 1030 210 1070 250
rect 930 190 1070 210
rect 930 150 970 190
rect 1030 150 1070 190
rect 930 110 1070 150
rect 1170 1090 1310 1110
rect 1170 1050 1210 1090
rect 1270 1050 1310 1090
rect 1170 1030 1310 1050
rect 1170 990 1210 1030
rect 1270 990 1310 1030
rect 1170 970 1310 990
rect 1170 930 1210 970
rect 1270 930 1310 970
rect 1170 910 1310 930
rect 1170 870 1210 910
rect 1270 870 1310 910
rect 1170 850 1310 870
rect 1170 810 1210 850
rect 1270 810 1310 850
rect 1170 790 1310 810
rect 1170 750 1210 790
rect 1270 750 1310 790
rect 1170 730 1310 750
rect 1170 690 1210 730
rect 1270 690 1310 730
rect 1170 670 1310 690
rect 1170 630 1210 670
rect 1270 630 1310 670
rect 1170 610 1310 630
rect 1170 570 1210 610
rect 1270 570 1310 610
rect 1170 550 1310 570
rect 1170 510 1210 550
rect 1270 510 1310 550
rect 1170 490 1310 510
rect 1170 450 1210 490
rect 1270 450 1310 490
rect 1170 430 1310 450
rect 1170 390 1210 430
rect 1270 390 1310 430
rect 1170 370 1310 390
rect 1170 330 1210 370
rect 1270 330 1310 370
rect 1170 310 1310 330
rect 1170 270 1210 310
rect 1270 270 1310 310
rect 1170 250 1310 270
rect 1170 210 1210 250
rect 1270 210 1310 250
rect 1170 190 1310 210
rect 1170 150 1210 190
rect 1270 150 1310 190
rect 1170 110 1310 150
rect 1410 1090 1550 1110
rect 1410 1050 1450 1090
rect 1510 1050 1550 1090
rect 1410 1030 1550 1050
rect 1410 990 1450 1030
rect 1510 990 1550 1030
rect 1410 970 1550 990
rect 1410 930 1450 970
rect 1510 930 1550 970
rect 1410 910 1550 930
rect 1410 870 1450 910
rect 1510 870 1550 910
rect 1410 850 1550 870
rect 1410 810 1450 850
rect 1510 810 1550 850
rect 1410 790 1550 810
rect 1410 750 1450 790
rect 1510 750 1550 790
rect 1410 730 1550 750
rect 1410 690 1450 730
rect 1510 690 1550 730
rect 1410 670 1550 690
rect 1410 630 1450 670
rect 1510 630 1550 670
rect 1410 610 1550 630
rect 1410 570 1450 610
rect 1510 570 1550 610
rect 1410 550 1550 570
rect 1410 510 1450 550
rect 1510 510 1550 550
rect 1410 490 1550 510
rect 1410 450 1450 490
rect 1510 450 1550 490
rect 1410 430 1550 450
rect 1410 390 1450 430
rect 1510 390 1550 430
rect 1410 370 1550 390
rect 1410 330 1450 370
rect 1510 330 1550 370
rect 1410 310 1550 330
rect 1410 270 1450 310
rect 1510 270 1550 310
rect 1410 250 1550 270
rect 1410 210 1450 250
rect 1510 210 1550 250
rect 1410 190 1550 210
rect 1410 150 1450 190
rect 1510 150 1550 190
rect 1410 110 1550 150
rect 1660 1090 1800 1110
rect 1660 1050 1700 1090
rect 1760 1050 1800 1090
rect 1660 1030 1800 1050
rect 1660 990 1700 1030
rect 1760 990 1800 1030
rect 1660 970 1800 990
rect 1660 930 1700 970
rect 1760 930 1800 970
rect 1660 910 1800 930
rect 1660 870 1700 910
rect 1760 870 1800 910
rect 1660 850 1800 870
rect 1660 810 1700 850
rect 1760 810 1800 850
rect 1660 790 1800 810
rect 1660 750 1700 790
rect 1760 750 1800 790
rect 1660 730 1800 750
rect 1660 690 1700 730
rect 1760 690 1800 730
rect 1660 670 1800 690
rect 1660 630 1700 670
rect 1760 630 1800 670
rect 1660 610 1800 630
rect 1660 570 1700 610
rect 1760 570 1800 610
rect 1660 550 1800 570
rect 1660 510 1700 550
rect 1760 510 1800 550
rect 1660 490 1800 510
rect 1660 450 1700 490
rect 1760 450 1800 490
rect 1660 430 1800 450
rect 1660 390 1700 430
rect 1760 390 1800 430
rect 1660 370 1800 390
rect 1660 330 1700 370
rect 1760 330 1800 370
rect 1660 310 1800 330
rect 1660 270 1700 310
rect 1760 270 1800 310
rect 1660 250 1800 270
rect 1660 210 1700 250
rect 1760 210 1800 250
rect 1660 190 1800 210
rect 1660 150 1700 190
rect 1760 150 1800 190
rect 1660 110 1800 150
rect 1900 1090 2040 1110
rect 1900 1050 1940 1090
rect 2000 1050 2040 1090
rect 1900 1030 2040 1050
rect 1900 990 1940 1030
rect 2000 990 2040 1030
rect 1900 970 2040 990
rect 1900 930 1940 970
rect 2000 930 2040 970
rect 1900 910 2040 930
rect 1900 870 1940 910
rect 2000 870 2040 910
rect 1900 850 2040 870
rect 1900 810 1940 850
rect 2000 810 2040 850
rect 1900 790 2040 810
rect 1900 750 1940 790
rect 2000 750 2040 790
rect 1900 730 2040 750
rect 1900 690 1940 730
rect 2000 690 2040 730
rect 1900 670 2040 690
rect 1900 630 1940 670
rect 2000 630 2040 670
rect 1900 610 2040 630
rect 1900 570 1940 610
rect 2000 570 2040 610
rect 1900 550 2040 570
rect 1900 510 1940 550
rect 2000 510 2040 550
rect 1900 490 2040 510
rect 1900 450 1940 490
rect 2000 450 2040 490
rect 1900 430 2040 450
rect 1900 390 1940 430
rect 2000 390 2040 430
rect 1900 370 2040 390
rect 1900 330 1940 370
rect 2000 330 2040 370
rect 1900 310 2040 330
rect 1900 270 1940 310
rect 2000 270 2040 310
rect 1900 250 2040 270
rect 1900 210 1940 250
rect 2000 210 2040 250
rect 1900 190 2040 210
rect 1900 150 1940 190
rect 2000 150 2040 190
rect 1900 110 2040 150
rect 2140 1090 2280 1110
rect 2140 1050 2180 1090
rect 2240 1050 2280 1090
rect 2140 1030 2280 1050
rect 2140 990 2180 1030
rect 2240 990 2280 1030
rect 2140 970 2280 990
rect 2140 930 2180 970
rect 2240 930 2280 970
rect 2140 910 2280 930
rect 2140 870 2180 910
rect 2240 870 2280 910
rect 2140 850 2280 870
rect 2140 810 2180 850
rect 2240 810 2280 850
rect 2140 790 2280 810
rect 2140 750 2180 790
rect 2240 750 2280 790
rect 2140 730 2280 750
rect 2140 690 2180 730
rect 2240 690 2280 730
rect 2140 670 2280 690
rect 2140 630 2180 670
rect 2240 630 2280 670
rect 2140 610 2280 630
rect 2140 570 2180 610
rect 2240 570 2280 610
rect 2140 550 2280 570
rect 2140 510 2180 550
rect 2240 510 2280 550
rect 2140 490 2280 510
rect 2140 450 2180 490
rect 2240 450 2280 490
rect 2140 430 2280 450
rect 2140 390 2180 430
rect 2240 390 2280 430
rect 2140 370 2280 390
rect 2140 330 2180 370
rect 2240 330 2280 370
rect 2140 310 2280 330
rect 2140 270 2180 310
rect 2240 270 2280 310
rect 2140 250 2280 270
rect 2140 210 2180 250
rect 2240 210 2280 250
rect 2140 190 2280 210
rect 2140 150 2180 190
rect 2240 150 2280 190
rect 2140 110 2280 150
rect 2390 1090 2530 1110
rect 2390 1050 2420 1090
rect 2480 1050 2530 1090
rect 2390 1030 2530 1050
rect 2390 990 2420 1030
rect 2480 990 2530 1030
rect 2390 970 2530 990
rect 2390 930 2420 970
rect 2480 930 2530 970
rect 2390 910 2530 930
rect 2390 870 2420 910
rect 2480 870 2530 910
rect 2390 850 2530 870
rect 2390 810 2420 850
rect 2480 810 2530 850
rect 2390 790 2530 810
rect 2390 750 2420 790
rect 2480 750 2530 790
rect 2390 730 2530 750
rect 2390 690 2420 730
rect 2480 690 2530 730
rect 2390 670 2530 690
rect 2390 630 2420 670
rect 2480 630 2530 670
rect 2390 610 2530 630
rect 2390 570 2420 610
rect 2480 570 2530 610
rect 2390 550 2530 570
rect 2390 510 2420 550
rect 2480 510 2530 550
rect 2390 490 2530 510
rect 2390 450 2420 490
rect 2480 450 2530 490
rect 2390 430 2530 450
rect 2390 390 2420 430
rect 2480 390 2530 430
rect 2390 370 2530 390
rect 2390 330 2420 370
rect 2480 330 2530 370
rect 2390 310 2530 330
rect 2390 270 2420 310
rect 2480 270 2530 310
rect 2390 250 2530 270
rect 2390 210 2420 250
rect 2480 210 2530 250
rect 2390 190 2530 210
rect 2390 150 2420 190
rect 2480 150 2530 190
rect 2390 110 2530 150
rect 2630 1090 2770 1110
rect 2630 1050 2670 1090
rect 2730 1050 2770 1090
rect 2630 1030 2770 1050
rect 2630 990 2670 1030
rect 2730 990 2770 1030
rect 2630 970 2770 990
rect 2630 930 2670 970
rect 2730 930 2770 970
rect 2630 910 2770 930
rect 2630 870 2670 910
rect 2730 870 2770 910
rect 2630 850 2770 870
rect 2630 810 2670 850
rect 2730 810 2770 850
rect 2630 790 2770 810
rect 2630 750 2670 790
rect 2730 750 2770 790
rect 2630 730 2770 750
rect 2630 690 2670 730
rect 2730 690 2770 730
rect 2630 670 2770 690
rect 2630 630 2670 670
rect 2730 630 2770 670
rect 2630 610 2770 630
rect 2630 570 2670 610
rect 2730 570 2770 610
rect 2630 550 2770 570
rect 2630 510 2670 550
rect 2730 510 2770 550
rect 2630 490 2770 510
rect 2630 450 2670 490
rect 2730 450 2770 490
rect 2630 430 2770 450
rect 2630 390 2670 430
rect 2730 390 2770 430
rect 2630 370 2770 390
rect 2630 330 2670 370
rect 2730 330 2770 370
rect 2630 310 2770 330
rect 2630 270 2670 310
rect 2730 270 2770 310
rect 2630 250 2770 270
rect 2630 210 2670 250
rect 2730 210 2770 250
rect 2630 190 2770 210
rect 2630 150 2670 190
rect 2730 150 2770 190
rect 2630 110 2770 150
rect 2870 1090 3010 1110
rect 2870 1050 2900 1090
rect 2960 1050 3010 1090
rect 2870 1030 3010 1050
rect 2870 990 2900 1030
rect 2960 990 3010 1030
rect 2870 970 3010 990
rect 2870 930 2900 970
rect 2960 930 3010 970
rect 2870 910 3010 930
rect 2870 870 2900 910
rect 2960 870 3010 910
rect 2870 850 3010 870
rect 2870 810 2900 850
rect 2960 810 3010 850
rect 2870 790 3010 810
rect 2870 750 2900 790
rect 2960 750 3010 790
rect 2870 730 3010 750
rect 2870 690 2900 730
rect 2960 690 3010 730
rect 2870 670 3010 690
rect 2870 630 2900 670
rect 2960 630 3010 670
rect 2870 610 3010 630
rect 2870 570 2900 610
rect 2960 570 3010 610
rect 2870 550 3010 570
rect 2870 510 2900 550
rect 2960 510 3010 550
rect 2870 490 3010 510
rect 2870 450 2900 490
rect 2960 450 3010 490
rect 2870 430 3010 450
rect 2870 390 2900 430
rect 2960 390 3010 430
rect 2870 370 3010 390
rect 2870 330 2900 370
rect 2960 330 3010 370
rect 2870 310 3010 330
rect 2870 270 2900 310
rect 2960 270 3010 310
rect 2870 250 3010 270
rect 2870 210 2900 250
rect 2960 210 3010 250
rect 2870 190 3010 210
rect 2870 150 2900 190
rect 2960 150 3010 190
rect 2870 110 3010 150
<< via1 >>
rect 0 1050 60 1090
rect 0 990 60 1030
rect 0 930 60 970
rect 0 870 60 910
rect 0 810 60 850
rect 0 750 60 790
rect 0 690 60 730
rect 0 630 60 670
rect 0 570 60 610
rect 0 510 60 550
rect 0 450 60 490
rect 0 390 60 430
rect 0 330 60 370
rect 0 270 60 310
rect 0 210 60 250
rect 0 150 60 190
rect 240 1050 300 1090
rect 240 990 300 1030
rect 240 930 300 970
rect 240 870 300 910
rect 240 810 300 850
rect 240 750 300 790
rect 240 690 300 730
rect 240 630 300 670
rect 240 570 300 610
rect 240 510 300 550
rect 240 450 300 490
rect 240 390 300 430
rect 240 330 300 370
rect 240 270 300 310
rect 240 210 300 250
rect 240 150 300 190
rect 480 1050 540 1090
rect 480 990 540 1030
rect 480 930 540 970
rect 480 870 540 910
rect 480 810 540 850
rect 480 750 540 790
rect 480 690 540 730
rect 480 630 540 670
rect 480 570 540 610
rect 480 510 540 550
rect 480 450 540 490
rect 480 390 540 430
rect 480 330 540 370
rect 480 270 540 310
rect 480 210 540 250
rect 480 150 540 190
rect 730 1050 790 1090
rect 730 990 790 1030
rect 730 930 790 970
rect 730 870 790 910
rect 730 810 790 850
rect 730 750 790 790
rect 730 690 790 730
rect 730 630 790 670
rect 730 570 790 610
rect 730 510 790 550
rect 730 450 790 490
rect 730 390 790 430
rect 730 330 790 370
rect 730 270 790 310
rect 730 210 790 250
rect 730 150 790 190
rect 970 1050 1030 1090
rect 970 990 1030 1030
rect 970 930 1030 970
rect 970 870 1030 910
rect 970 810 1030 850
rect 970 750 1030 790
rect 970 690 1030 730
rect 970 630 1030 670
rect 970 570 1030 610
rect 970 510 1030 550
rect 970 450 1030 490
rect 970 390 1030 430
rect 970 330 1030 370
rect 970 270 1030 310
rect 970 210 1030 250
rect 970 150 1030 190
rect 1210 1050 1270 1090
rect 1210 990 1270 1030
rect 1210 930 1270 970
rect 1210 870 1270 910
rect 1210 810 1270 850
rect 1210 750 1270 790
rect 1210 690 1270 730
rect 1210 630 1270 670
rect 1210 570 1270 610
rect 1210 510 1270 550
rect 1210 450 1270 490
rect 1210 390 1270 430
rect 1210 330 1270 370
rect 1210 270 1270 310
rect 1210 210 1270 250
rect 1210 150 1270 190
rect 1450 1050 1510 1090
rect 1450 990 1510 1030
rect 1450 930 1510 970
rect 1450 870 1510 910
rect 1450 810 1510 850
rect 1450 750 1510 790
rect 1450 690 1510 730
rect 1450 630 1510 670
rect 1450 570 1510 610
rect 1450 510 1510 550
rect 1450 450 1510 490
rect 1450 390 1510 430
rect 1450 330 1510 370
rect 1450 270 1510 310
rect 1450 210 1510 250
rect 1450 150 1510 190
rect 1700 1050 1760 1090
rect 1700 990 1760 1030
rect 1700 930 1760 970
rect 1700 870 1760 910
rect 1700 810 1760 850
rect 1700 750 1760 790
rect 1700 690 1760 730
rect 1700 630 1760 670
rect 1700 570 1760 610
rect 1700 510 1760 550
rect 1700 450 1760 490
rect 1700 390 1760 430
rect 1700 330 1760 370
rect 1700 270 1760 310
rect 1700 210 1760 250
rect 1700 150 1760 190
rect 1940 1050 2000 1090
rect 1940 990 2000 1030
rect 1940 930 2000 970
rect 1940 870 2000 910
rect 1940 810 2000 850
rect 1940 750 2000 790
rect 1940 690 2000 730
rect 1940 630 2000 670
rect 1940 570 2000 610
rect 1940 510 2000 550
rect 1940 450 2000 490
rect 1940 390 2000 430
rect 1940 330 2000 370
rect 1940 270 2000 310
rect 1940 210 2000 250
rect 1940 150 2000 190
rect 2180 1050 2240 1090
rect 2180 990 2240 1030
rect 2180 930 2240 970
rect 2180 870 2240 910
rect 2180 810 2240 850
rect 2180 750 2240 790
rect 2180 690 2240 730
rect 2180 630 2240 670
rect 2180 570 2240 610
rect 2180 510 2240 550
rect 2180 450 2240 490
rect 2180 390 2240 430
rect 2180 330 2240 370
rect 2180 270 2240 310
rect 2180 210 2240 250
rect 2180 150 2240 190
rect 2420 1050 2480 1090
rect 2420 990 2480 1030
rect 2420 930 2480 970
rect 2420 870 2480 910
rect 2420 810 2480 850
rect 2420 750 2480 790
rect 2420 690 2480 730
rect 2420 630 2480 670
rect 2420 570 2480 610
rect 2420 510 2480 550
rect 2420 450 2480 490
rect 2420 390 2480 430
rect 2420 330 2480 370
rect 2420 270 2480 310
rect 2420 210 2480 250
rect 2420 150 2480 190
rect 2670 1050 2730 1090
rect 2670 990 2730 1030
rect 2670 930 2730 970
rect 2670 870 2730 910
rect 2670 810 2730 850
rect 2670 750 2730 790
rect 2670 690 2730 730
rect 2670 630 2730 670
rect 2670 570 2730 610
rect 2670 510 2730 550
rect 2670 450 2730 490
rect 2670 390 2730 430
rect 2670 330 2730 370
rect 2670 270 2730 310
rect 2670 210 2730 250
rect 2670 150 2730 190
rect 2900 1050 2960 1090
rect 2900 990 2960 1030
rect 2900 930 2960 970
rect 2900 870 2960 910
rect 2900 810 2960 850
rect 2900 750 2960 790
rect 2900 690 2960 730
rect 2900 630 2960 670
rect 2900 570 2960 610
rect 2900 510 2960 550
rect 2900 450 2960 490
rect 2900 390 2960 430
rect 2900 330 2960 370
rect 2900 270 2960 310
rect 2900 210 2960 250
rect 2900 150 2960 190
<< metal2 >>
rect 1410 1180 1550 1250
rect 50 1130 2890 1180
rect -40 1090 100 1110
rect -40 1050 0 1090
rect 60 1050 100 1090
rect -40 1030 100 1050
rect -40 990 0 1030
rect 60 990 100 1030
rect -40 970 100 990
rect -40 930 0 970
rect 60 930 100 970
rect -40 910 100 930
rect -40 870 0 910
rect 60 870 100 910
rect -40 850 100 870
rect -40 810 0 850
rect 60 810 100 850
rect -40 790 100 810
rect -40 750 0 790
rect 60 750 100 790
rect -40 730 100 750
rect -40 690 0 730
rect 60 690 100 730
rect -40 670 100 690
rect -40 630 0 670
rect 60 630 100 670
rect -40 610 100 630
rect -40 570 0 610
rect 60 570 100 610
rect -40 550 100 570
rect -40 510 0 550
rect 60 510 100 550
rect -40 490 100 510
rect -40 450 0 490
rect 60 450 100 490
rect -40 430 100 450
rect -40 390 0 430
rect 60 390 100 430
rect -40 370 100 390
rect -40 330 0 370
rect 60 330 100 370
rect -40 310 100 330
rect -40 270 0 310
rect 60 270 100 310
rect -40 250 100 270
rect -40 210 0 250
rect 60 210 100 250
rect -40 190 100 210
rect -40 150 0 190
rect 60 150 100 190
rect -40 110 100 150
rect 200 1090 340 1110
rect 200 1050 240 1090
rect 300 1050 340 1090
rect 200 1030 340 1050
rect 200 990 240 1030
rect 300 990 340 1030
rect 200 970 340 990
rect 200 930 240 970
rect 300 930 340 970
rect 200 910 340 930
rect 200 870 240 910
rect 300 870 340 910
rect 200 850 340 870
rect 200 810 240 850
rect 300 810 340 850
rect 200 790 340 810
rect 200 750 240 790
rect 300 750 340 790
rect 200 730 340 750
rect 200 690 240 730
rect 300 690 340 730
rect 200 670 340 690
rect 200 630 240 670
rect 300 630 340 670
rect 200 610 340 630
rect 200 570 240 610
rect 300 570 340 610
rect 200 550 340 570
rect 200 510 240 550
rect 300 510 340 550
rect 200 490 340 510
rect 200 450 240 490
rect 300 450 340 490
rect 200 430 340 450
rect 200 390 240 430
rect 300 390 340 430
rect 200 370 340 390
rect 200 330 240 370
rect 300 330 340 370
rect 200 310 340 330
rect 200 270 240 310
rect 300 270 340 310
rect 200 250 340 270
rect 200 210 240 250
rect 300 210 340 250
rect 200 190 340 210
rect 200 150 240 190
rect 300 150 340 190
rect 200 110 340 150
rect 440 1090 580 1110
rect 440 1050 480 1090
rect 540 1050 580 1090
rect 440 1030 580 1050
rect 440 990 480 1030
rect 540 990 580 1030
rect 440 970 580 990
rect 440 930 480 970
rect 540 930 580 970
rect 440 910 580 930
rect 440 870 480 910
rect 540 870 580 910
rect 440 850 580 870
rect 440 810 480 850
rect 540 810 580 850
rect 440 790 580 810
rect 440 750 480 790
rect 540 750 580 790
rect 440 730 580 750
rect 440 690 480 730
rect 540 690 580 730
rect 440 670 580 690
rect 440 630 480 670
rect 540 630 580 670
rect 440 610 580 630
rect 440 570 480 610
rect 540 570 580 610
rect 440 550 580 570
rect 440 510 480 550
rect 540 510 580 550
rect 440 490 580 510
rect 440 450 480 490
rect 540 450 580 490
rect 440 430 580 450
rect 440 390 480 430
rect 540 390 580 430
rect 440 370 580 390
rect 440 330 480 370
rect 540 330 580 370
rect 440 310 580 330
rect 440 270 480 310
rect 540 270 580 310
rect 440 250 580 270
rect 440 210 480 250
rect 540 210 580 250
rect 440 190 580 210
rect 440 150 480 190
rect 540 150 580 190
rect 440 110 580 150
rect 680 1090 820 1110
rect 680 1050 730 1090
rect 790 1050 820 1090
rect 680 1030 820 1050
rect 680 990 730 1030
rect 790 990 820 1030
rect 680 970 820 990
rect 680 930 730 970
rect 790 930 820 970
rect 680 910 820 930
rect 680 870 730 910
rect 790 870 820 910
rect 680 850 820 870
rect 680 810 730 850
rect 790 810 820 850
rect 680 790 820 810
rect 680 750 730 790
rect 790 750 820 790
rect 680 730 820 750
rect 680 690 730 730
rect 790 690 820 730
rect 680 670 820 690
rect 680 630 730 670
rect 790 630 820 670
rect 680 610 820 630
rect 680 570 730 610
rect 790 570 820 610
rect 680 550 820 570
rect 680 510 730 550
rect 790 510 820 550
rect 680 490 820 510
rect 680 450 730 490
rect 790 450 820 490
rect 680 430 820 450
rect 680 390 730 430
rect 790 390 820 430
rect 680 370 820 390
rect 680 330 730 370
rect 790 330 820 370
rect 680 310 820 330
rect 680 270 730 310
rect 790 270 820 310
rect 680 250 820 270
rect 680 210 730 250
rect 790 210 820 250
rect 680 190 820 210
rect 680 150 730 190
rect 790 150 820 190
rect 680 110 820 150
rect 930 1090 1070 1110
rect 930 1050 970 1090
rect 1030 1050 1070 1090
rect 930 1030 1070 1050
rect 930 990 970 1030
rect 1030 990 1070 1030
rect 930 970 1070 990
rect 930 930 970 970
rect 1030 930 1070 970
rect 930 910 1070 930
rect 930 870 970 910
rect 1030 870 1070 910
rect 930 850 1070 870
rect 930 810 970 850
rect 1030 810 1070 850
rect 930 790 1070 810
rect 930 750 970 790
rect 1030 750 1070 790
rect 930 730 1070 750
rect 930 690 970 730
rect 1030 690 1070 730
rect 930 670 1070 690
rect 930 630 970 670
rect 1030 630 1070 670
rect 930 610 1070 630
rect 930 570 970 610
rect 1030 570 1070 610
rect 930 550 1070 570
rect 930 510 970 550
rect 1030 510 1070 550
rect 930 490 1070 510
rect 930 450 970 490
rect 1030 450 1070 490
rect 930 430 1070 450
rect 930 390 970 430
rect 1030 390 1070 430
rect 930 370 1070 390
rect 930 330 970 370
rect 1030 330 1070 370
rect 930 310 1070 330
rect 930 270 970 310
rect 1030 270 1070 310
rect 930 250 1070 270
rect 930 210 970 250
rect 1030 210 1070 250
rect 930 190 1070 210
rect 930 150 970 190
rect 1030 150 1070 190
rect 930 110 1070 150
rect 1170 1090 1310 1110
rect 1170 1050 1210 1090
rect 1270 1050 1310 1090
rect 1170 1030 1310 1050
rect 1170 990 1210 1030
rect 1270 990 1310 1030
rect 1170 970 1310 990
rect 1170 930 1210 970
rect 1270 930 1310 970
rect 1170 910 1310 930
rect 1170 870 1210 910
rect 1270 870 1310 910
rect 1170 850 1310 870
rect 1170 810 1210 850
rect 1270 810 1310 850
rect 1170 790 1310 810
rect 1170 750 1210 790
rect 1270 750 1310 790
rect 1170 730 1310 750
rect 1170 690 1210 730
rect 1270 690 1310 730
rect 1170 670 1310 690
rect 1170 630 1210 670
rect 1270 630 1310 670
rect 1170 610 1310 630
rect 1170 570 1210 610
rect 1270 570 1310 610
rect 1170 550 1310 570
rect 1170 510 1210 550
rect 1270 510 1310 550
rect 1170 490 1310 510
rect 1170 450 1210 490
rect 1270 450 1310 490
rect 1170 430 1310 450
rect 1170 390 1210 430
rect 1270 390 1310 430
rect 1170 370 1310 390
rect 1170 330 1210 370
rect 1270 330 1310 370
rect 1170 310 1310 330
rect 1170 270 1210 310
rect 1270 270 1310 310
rect 1170 250 1310 270
rect 1170 210 1210 250
rect 1270 210 1310 250
rect 1170 190 1310 210
rect 1170 150 1210 190
rect 1270 150 1310 190
rect 1170 110 1310 150
rect 1410 1090 1550 1130
rect 1410 1050 1450 1090
rect 1510 1050 1550 1090
rect 1410 1030 1550 1050
rect 1410 990 1450 1030
rect 1510 990 1550 1030
rect 1410 970 1550 990
rect 1410 930 1450 970
rect 1510 930 1550 970
rect 1410 910 1550 930
rect 1410 870 1450 910
rect 1510 870 1550 910
rect 1410 850 1550 870
rect 1410 810 1450 850
rect 1510 810 1550 850
rect 1410 790 1550 810
rect 1410 750 1450 790
rect 1510 750 1550 790
rect 1410 730 1550 750
rect 1410 690 1450 730
rect 1510 690 1550 730
rect 1410 670 1550 690
rect 1410 630 1450 670
rect 1510 630 1550 670
rect 1410 610 1550 630
rect 1410 570 1450 610
rect 1510 570 1550 610
rect 1410 550 1550 570
rect 1410 510 1450 550
rect 1510 510 1550 550
rect 1410 490 1550 510
rect 1410 450 1450 490
rect 1510 450 1550 490
rect 1410 430 1550 450
rect 1410 390 1450 430
rect 1510 390 1550 430
rect 1410 370 1550 390
rect 1410 330 1450 370
rect 1510 330 1550 370
rect 1410 310 1550 330
rect 1410 270 1450 310
rect 1510 270 1550 310
rect 1410 250 1550 270
rect 1410 210 1450 250
rect 1510 210 1550 250
rect 1410 190 1550 210
rect 1410 150 1450 190
rect 1510 150 1550 190
rect 1410 90 1550 150
rect 1660 1090 1800 1110
rect 1660 1050 1700 1090
rect 1760 1050 1800 1090
rect 1660 1030 1800 1050
rect 1660 990 1700 1030
rect 1760 990 1800 1030
rect 1660 970 1800 990
rect 1660 930 1700 970
rect 1760 930 1800 970
rect 1660 910 1800 930
rect 1660 870 1700 910
rect 1760 870 1800 910
rect 1660 850 1800 870
rect 1660 810 1700 850
rect 1760 810 1800 850
rect 1660 790 1800 810
rect 1660 750 1700 790
rect 1760 750 1800 790
rect 1660 730 1800 750
rect 1660 690 1700 730
rect 1760 690 1800 730
rect 1660 670 1800 690
rect 1660 630 1700 670
rect 1760 630 1800 670
rect 1660 610 1800 630
rect 1660 570 1700 610
rect 1760 570 1800 610
rect 1660 550 1800 570
rect 1660 510 1700 550
rect 1760 510 1800 550
rect 1660 490 1800 510
rect 1660 450 1700 490
rect 1760 450 1800 490
rect 1660 430 1800 450
rect 1660 390 1700 430
rect 1760 390 1800 430
rect 1660 370 1800 390
rect 1660 330 1700 370
rect 1760 330 1800 370
rect 1660 310 1800 330
rect 1660 270 1700 310
rect 1760 270 1800 310
rect 1660 250 1800 270
rect 1660 210 1700 250
rect 1760 210 1800 250
rect 1660 190 1800 210
rect 1660 150 1700 190
rect 1760 150 1800 190
rect 1660 110 1800 150
rect 1900 1090 2040 1110
rect 1900 1050 1940 1090
rect 2000 1050 2040 1090
rect 1900 1030 2040 1050
rect 1900 990 1940 1030
rect 2000 990 2040 1030
rect 1900 970 2040 990
rect 1900 930 1940 970
rect 2000 930 2040 970
rect 1900 910 2040 930
rect 1900 870 1940 910
rect 2000 870 2040 910
rect 1900 850 2040 870
rect 1900 810 1940 850
rect 2000 810 2040 850
rect 1900 790 2040 810
rect 1900 750 1940 790
rect 2000 750 2040 790
rect 1900 730 2040 750
rect 1900 690 1940 730
rect 2000 690 2040 730
rect 1900 670 2040 690
rect 1900 630 1940 670
rect 2000 630 2040 670
rect 1900 610 2040 630
rect 1900 570 1940 610
rect 2000 570 2040 610
rect 1900 550 2040 570
rect 1900 510 1940 550
rect 2000 510 2040 550
rect 1900 490 2040 510
rect 1900 450 1940 490
rect 2000 450 2040 490
rect 1900 430 2040 450
rect 1900 390 1940 430
rect 2000 390 2040 430
rect 1900 370 2040 390
rect 1900 330 1940 370
rect 2000 330 2040 370
rect 1900 310 2040 330
rect 1900 270 1940 310
rect 2000 270 2040 310
rect 1900 250 2040 270
rect 1900 210 1940 250
rect 2000 210 2040 250
rect 1900 190 2040 210
rect 1900 150 1940 190
rect 2000 150 2040 190
rect 1900 110 2040 150
rect 2140 1090 2280 1110
rect 2140 1050 2180 1090
rect 2240 1050 2280 1090
rect 2140 1030 2280 1050
rect 2140 990 2180 1030
rect 2240 990 2280 1030
rect 2140 970 2280 990
rect 2140 930 2180 970
rect 2240 930 2280 970
rect 2140 910 2280 930
rect 2140 870 2180 910
rect 2240 870 2280 910
rect 2140 850 2280 870
rect 2140 810 2180 850
rect 2240 810 2280 850
rect 2140 790 2280 810
rect 2140 750 2180 790
rect 2240 750 2280 790
rect 2140 730 2280 750
rect 2140 690 2180 730
rect 2240 690 2280 730
rect 2140 670 2280 690
rect 2140 630 2180 670
rect 2240 630 2280 670
rect 2140 610 2280 630
rect 2140 570 2180 610
rect 2240 570 2280 610
rect 2140 550 2280 570
rect 2140 510 2180 550
rect 2240 510 2280 550
rect 2140 490 2280 510
rect 2140 450 2180 490
rect 2240 450 2280 490
rect 2140 430 2280 450
rect 2140 390 2180 430
rect 2240 390 2280 430
rect 2140 370 2280 390
rect 2140 330 2180 370
rect 2240 330 2280 370
rect 2140 310 2280 330
rect 2140 270 2180 310
rect 2240 270 2280 310
rect 2140 250 2280 270
rect 2140 210 2180 250
rect 2240 210 2280 250
rect 2140 190 2280 210
rect 2140 150 2180 190
rect 2240 150 2280 190
rect 2140 110 2280 150
rect 2380 1090 2520 1110
rect 2380 1050 2420 1090
rect 2480 1050 2520 1090
rect 2380 1030 2520 1050
rect 2380 990 2420 1030
rect 2480 990 2520 1030
rect 2380 970 2520 990
rect 2380 930 2420 970
rect 2480 930 2520 970
rect 2380 910 2520 930
rect 2380 870 2420 910
rect 2480 870 2520 910
rect 2380 850 2520 870
rect 2380 810 2420 850
rect 2480 810 2520 850
rect 2380 790 2520 810
rect 2380 750 2420 790
rect 2480 750 2520 790
rect 2380 730 2520 750
rect 2380 690 2420 730
rect 2480 690 2520 730
rect 2380 670 2520 690
rect 2380 630 2420 670
rect 2480 630 2520 670
rect 2380 610 2520 630
rect 2380 570 2420 610
rect 2480 570 2520 610
rect 2380 550 2520 570
rect 2380 510 2420 550
rect 2480 510 2520 550
rect 2380 490 2520 510
rect 2380 450 2420 490
rect 2480 450 2520 490
rect 2380 430 2520 450
rect 2380 390 2420 430
rect 2480 390 2520 430
rect 2380 370 2520 390
rect 2380 330 2420 370
rect 2480 330 2520 370
rect 2380 310 2520 330
rect 2380 270 2420 310
rect 2480 270 2520 310
rect 2380 250 2520 270
rect 2380 210 2420 250
rect 2480 210 2520 250
rect 2380 190 2520 210
rect 2380 150 2420 190
rect 2480 150 2520 190
rect 2380 110 2520 150
rect 2630 1090 2770 1110
rect 2630 1050 2670 1090
rect 2730 1050 2770 1090
rect 2630 1030 2770 1050
rect 2630 990 2670 1030
rect 2730 990 2770 1030
rect 2630 970 2770 990
rect 2630 930 2670 970
rect 2730 930 2770 970
rect 2630 910 2770 930
rect 2630 870 2670 910
rect 2730 870 2770 910
rect 2630 850 2770 870
rect 2630 810 2670 850
rect 2730 810 2770 850
rect 2630 790 2770 810
rect 2630 750 2670 790
rect 2730 750 2770 790
rect 2630 730 2770 750
rect 2630 690 2670 730
rect 2730 690 2770 730
rect 2630 670 2770 690
rect 2630 630 2670 670
rect 2730 630 2770 670
rect 2630 610 2770 630
rect 2630 570 2670 610
rect 2730 570 2770 610
rect 2630 550 2770 570
rect 2630 510 2670 550
rect 2730 510 2770 550
rect 2630 490 2770 510
rect 2630 450 2670 490
rect 2730 450 2770 490
rect 2630 430 2770 450
rect 2630 390 2670 430
rect 2730 390 2770 430
rect 2630 370 2770 390
rect 2630 330 2670 370
rect 2730 330 2770 370
rect 2630 310 2770 330
rect 2630 270 2670 310
rect 2730 270 2770 310
rect 2630 250 2770 270
rect 2630 210 2670 250
rect 2730 210 2770 250
rect 2630 190 2770 210
rect 2630 150 2670 190
rect 2730 150 2770 190
rect 2630 110 2770 150
rect 2870 1090 3010 1110
rect 2870 1050 2900 1090
rect 2960 1050 3010 1090
rect 2870 1030 3010 1050
rect 2870 990 2900 1030
rect 2960 990 3010 1030
rect 2870 970 3010 990
rect 2870 930 2900 970
rect 2960 930 3010 970
rect 2870 910 3010 930
rect 2870 870 2900 910
rect 2960 870 3010 910
rect 2870 850 3010 870
rect 2870 810 2900 850
rect 2960 810 3010 850
rect 2870 790 3010 810
rect 2870 750 2900 790
rect 2960 750 3010 790
rect 2870 730 3010 750
rect 2870 690 2900 730
rect 2960 690 3010 730
rect 2870 670 3010 690
rect 2870 630 2900 670
rect 2960 630 3010 670
rect 2870 610 3010 630
rect 2870 570 2900 610
rect 2960 570 3010 610
rect 2870 550 3010 570
rect 2870 510 2900 550
rect 2960 510 3010 550
rect 2870 490 3010 510
rect 2870 450 2900 490
rect 2960 450 3010 490
rect 2870 430 3010 450
rect 2870 390 2900 430
rect 2960 390 3010 430
rect 2870 370 3010 390
rect 2870 330 2900 370
rect 2960 330 3010 370
rect 2870 310 3010 330
rect 2870 270 2900 310
rect 2960 270 3010 310
rect 2870 250 3010 270
rect 2870 210 2900 250
rect 2960 210 3010 250
rect 2870 190 3010 210
rect 2870 150 2900 190
rect 2960 150 3010 190
rect 2870 110 3010 150
rect 90 40 2930 90
<< via2 >>
rect 0 1050 60 1090
rect 0 990 60 1030
rect 0 930 60 970
rect 0 870 60 910
rect 0 810 60 850
rect 0 750 60 790
rect 0 690 60 730
rect 0 630 60 670
rect 0 570 60 610
rect 0 510 60 550
rect 0 450 60 490
rect 0 390 60 430
rect 0 330 60 370
rect 0 270 60 310
rect 0 210 60 250
rect 0 150 60 190
rect 240 1050 300 1090
rect 240 990 300 1030
rect 240 930 300 970
rect 240 870 300 910
rect 240 810 300 850
rect 240 750 300 790
rect 240 690 300 730
rect 240 630 300 670
rect 240 570 300 610
rect 240 510 300 550
rect 240 450 300 490
rect 240 390 300 430
rect 240 330 300 370
rect 240 270 300 310
rect 240 210 300 250
rect 240 150 300 190
rect 480 1050 540 1090
rect 480 990 540 1030
rect 480 930 540 970
rect 480 870 540 910
rect 480 810 540 850
rect 480 750 540 790
rect 480 690 540 730
rect 480 630 540 670
rect 480 570 540 610
rect 480 510 540 550
rect 480 450 540 490
rect 480 390 540 430
rect 480 330 540 370
rect 480 270 540 310
rect 480 210 540 250
rect 480 150 540 190
rect 730 1050 790 1090
rect 730 990 790 1030
rect 730 930 790 970
rect 730 870 790 910
rect 730 810 790 850
rect 730 750 790 790
rect 730 690 790 730
rect 730 630 790 670
rect 730 570 790 610
rect 730 510 790 550
rect 730 450 790 490
rect 730 390 790 430
rect 730 330 790 370
rect 730 270 790 310
rect 730 210 790 250
rect 730 150 790 190
rect 970 1050 1030 1090
rect 970 990 1030 1030
rect 970 930 1030 970
rect 970 870 1030 910
rect 970 810 1030 850
rect 970 750 1030 790
rect 970 690 1030 730
rect 970 630 1030 670
rect 970 570 1030 610
rect 970 510 1030 550
rect 970 450 1030 490
rect 970 390 1030 430
rect 970 330 1030 370
rect 970 270 1030 310
rect 970 210 1030 250
rect 970 150 1030 190
rect 1210 1050 1270 1090
rect 1210 990 1270 1030
rect 1210 930 1270 970
rect 1210 870 1270 910
rect 1210 810 1270 850
rect 1210 750 1270 790
rect 1210 690 1270 730
rect 1210 630 1270 670
rect 1210 570 1270 610
rect 1210 510 1270 550
rect 1210 450 1270 490
rect 1210 390 1270 430
rect 1210 330 1270 370
rect 1210 270 1270 310
rect 1210 210 1270 250
rect 1210 150 1270 190
rect 1700 1050 1760 1090
rect 1700 990 1760 1030
rect 1700 930 1760 970
rect 1700 870 1760 910
rect 1700 810 1760 850
rect 1700 750 1760 790
rect 1700 690 1760 730
rect 1700 630 1760 670
rect 1700 570 1760 610
rect 1700 510 1760 550
rect 1700 450 1760 490
rect 1700 390 1760 430
rect 1700 330 1760 370
rect 1700 270 1760 310
rect 1700 210 1760 250
rect 1700 150 1760 190
rect 1940 1050 2000 1090
rect 1940 990 2000 1030
rect 1940 930 2000 970
rect 1940 870 2000 910
rect 1940 810 2000 850
rect 1940 750 2000 790
rect 1940 690 2000 730
rect 1940 630 2000 670
rect 1940 570 2000 610
rect 1940 510 2000 550
rect 1940 450 2000 490
rect 1940 390 2000 430
rect 1940 330 2000 370
rect 1940 270 2000 310
rect 1940 210 2000 250
rect 1940 150 2000 190
rect 2180 1050 2240 1090
rect 2180 990 2240 1030
rect 2180 930 2240 970
rect 2180 870 2240 910
rect 2180 810 2240 850
rect 2180 750 2240 790
rect 2180 690 2240 730
rect 2180 630 2240 670
rect 2180 570 2240 610
rect 2180 510 2240 550
rect 2180 450 2240 490
rect 2180 390 2240 430
rect 2180 330 2240 370
rect 2180 270 2240 310
rect 2180 210 2240 250
rect 2180 150 2240 190
rect 2420 1050 2480 1090
rect 2420 990 2480 1030
rect 2420 930 2480 970
rect 2420 870 2480 910
rect 2420 810 2480 850
rect 2420 750 2480 790
rect 2420 690 2480 730
rect 2420 630 2480 670
rect 2420 570 2480 610
rect 2420 510 2480 550
rect 2420 450 2480 490
rect 2420 390 2480 430
rect 2420 330 2480 370
rect 2420 270 2480 310
rect 2420 210 2480 250
rect 2420 150 2480 190
rect 2670 1050 2730 1090
rect 2670 990 2730 1030
rect 2670 930 2730 970
rect 2670 870 2730 910
rect 2670 810 2730 850
rect 2670 750 2730 790
rect 2670 690 2730 730
rect 2670 630 2730 670
rect 2670 570 2730 610
rect 2670 510 2730 550
rect 2670 450 2730 490
rect 2670 390 2730 430
rect 2670 330 2730 370
rect 2670 270 2730 310
rect 2670 210 2730 250
rect 2670 150 2730 190
rect 2900 1050 2960 1090
rect 2900 990 2960 1030
rect 2900 930 2960 970
rect 2900 870 2960 910
rect 2900 810 2960 850
rect 2900 750 2960 790
rect 2900 690 2960 730
rect 2900 630 2960 670
rect 2900 570 2960 610
rect 2900 510 2960 550
rect 2900 450 2960 490
rect 2900 390 2960 430
rect 2900 330 2960 370
rect 2900 270 2960 310
rect 2900 210 2960 250
rect 2900 150 2960 190
<< metal3 >>
rect -40 1150 3010 1210
rect -40 1090 100 1150
rect -40 1050 0 1090
rect 60 1050 100 1090
rect -40 1030 100 1050
rect -40 990 0 1030
rect 60 990 100 1030
rect -40 970 100 990
rect -40 930 0 970
rect 60 930 100 970
rect -40 910 100 930
rect -40 870 0 910
rect 60 870 100 910
rect -40 850 100 870
rect -40 810 0 850
rect 60 810 100 850
rect -40 790 100 810
rect -40 750 0 790
rect 60 750 100 790
rect -40 730 100 750
rect -40 690 0 730
rect 60 690 100 730
rect -40 670 100 690
rect -40 630 0 670
rect 60 630 100 670
rect -40 610 100 630
rect -40 570 0 610
rect 60 570 100 610
rect -40 550 100 570
rect -40 510 0 550
rect 60 510 100 550
rect -40 490 100 510
rect -40 450 0 490
rect 60 450 100 490
rect -40 430 100 450
rect -40 390 0 430
rect 60 390 100 430
rect -40 370 100 390
rect -40 330 0 370
rect 60 330 100 370
rect -40 310 100 330
rect -40 270 0 310
rect 60 270 100 310
rect -40 250 100 270
rect -40 210 0 250
rect 60 210 100 250
rect -40 190 100 210
rect -40 150 0 190
rect 60 150 100 190
rect -40 110 100 150
rect 200 1090 340 1110
rect 200 1050 240 1090
rect 300 1050 340 1090
rect 200 1030 340 1050
rect 200 990 240 1030
rect 300 990 340 1030
rect 200 970 340 990
rect 200 930 240 970
rect 300 930 340 970
rect 200 910 340 930
rect 200 870 240 910
rect 300 870 340 910
rect 200 850 340 870
rect 200 810 240 850
rect 300 810 340 850
rect 200 790 340 810
rect 200 750 240 790
rect 300 750 340 790
rect 200 730 340 750
rect 200 690 240 730
rect 300 690 340 730
rect 200 670 340 690
rect 200 630 240 670
rect 300 630 340 670
rect 200 610 340 630
rect 200 570 240 610
rect 300 570 340 610
rect 200 550 340 570
rect 200 510 240 550
rect 300 510 340 550
rect 200 490 340 510
rect 200 450 240 490
rect 300 450 340 490
rect 200 430 340 450
rect 200 390 240 430
rect 300 390 340 430
rect 200 370 340 390
rect 200 330 240 370
rect 300 330 340 370
rect 200 310 340 330
rect 200 270 240 310
rect 300 270 340 310
rect 200 250 340 270
rect 200 210 240 250
rect 300 210 340 250
rect 200 190 340 210
rect 200 150 240 190
rect 300 150 340 190
rect 200 10 340 150
rect 440 1090 580 1150
rect 440 1050 480 1090
rect 540 1050 580 1090
rect 440 1030 580 1050
rect 440 990 480 1030
rect 540 990 580 1030
rect 440 970 580 990
rect 440 930 480 970
rect 540 930 580 970
rect 440 910 580 930
rect 440 870 480 910
rect 540 870 580 910
rect 440 850 580 870
rect 440 810 480 850
rect 540 810 580 850
rect 440 790 580 810
rect 440 750 480 790
rect 540 750 580 790
rect 440 730 580 750
rect 440 690 480 730
rect 540 690 580 730
rect 440 670 580 690
rect 440 630 480 670
rect 540 630 580 670
rect 440 610 580 630
rect 440 570 480 610
rect 540 570 580 610
rect 440 550 580 570
rect 440 510 480 550
rect 540 510 580 550
rect 440 490 580 510
rect 440 450 480 490
rect 540 450 580 490
rect 440 430 580 450
rect 440 390 480 430
rect 540 390 580 430
rect 440 370 580 390
rect 440 330 480 370
rect 540 330 580 370
rect 440 310 580 330
rect 440 270 480 310
rect 540 270 580 310
rect 440 250 580 270
rect 440 210 480 250
rect 540 210 580 250
rect 440 190 580 210
rect 440 150 480 190
rect 540 150 580 190
rect 440 110 580 150
rect 680 1090 820 1110
rect 680 1050 730 1090
rect 790 1050 820 1090
rect 680 1030 820 1050
rect 680 990 730 1030
rect 790 990 820 1030
rect 680 970 820 990
rect 680 930 730 970
rect 790 930 820 970
rect 680 910 820 930
rect 680 870 730 910
rect 790 870 820 910
rect 680 850 820 870
rect 680 810 730 850
rect 790 810 820 850
rect 680 790 820 810
rect 680 750 730 790
rect 790 750 820 790
rect 680 730 820 750
rect 680 690 730 730
rect 790 690 820 730
rect 680 670 820 690
rect 680 630 730 670
rect 790 630 820 670
rect 680 610 820 630
rect 680 570 730 610
rect 790 570 820 610
rect 680 550 820 570
rect 680 510 730 550
rect 790 510 820 550
rect 680 490 820 510
rect 680 450 730 490
rect 790 450 820 490
rect 680 430 820 450
rect 680 390 730 430
rect 790 390 820 430
rect 680 370 820 390
rect 680 330 730 370
rect 790 330 820 370
rect 680 310 820 330
rect 680 270 730 310
rect 790 270 820 310
rect 680 250 820 270
rect 680 210 730 250
rect 790 210 820 250
rect 680 190 820 210
rect 680 150 730 190
rect 790 150 820 190
rect 680 10 820 150
rect 930 1090 1070 1150
rect 930 1050 970 1090
rect 1030 1050 1070 1090
rect 930 1030 1070 1050
rect 930 990 970 1030
rect 1030 990 1070 1030
rect 930 970 1070 990
rect 930 930 970 970
rect 1030 930 1070 970
rect 930 910 1070 930
rect 930 870 970 910
rect 1030 870 1070 910
rect 930 850 1070 870
rect 930 810 970 850
rect 1030 810 1070 850
rect 930 790 1070 810
rect 930 750 970 790
rect 1030 750 1070 790
rect 930 730 1070 750
rect 930 690 970 730
rect 1030 690 1070 730
rect 930 670 1070 690
rect 930 630 970 670
rect 1030 630 1070 670
rect 930 610 1070 630
rect 930 570 970 610
rect 1030 570 1070 610
rect 930 550 1070 570
rect 930 510 970 550
rect 1030 510 1070 550
rect 930 490 1070 510
rect 930 450 970 490
rect 1030 450 1070 490
rect 930 430 1070 450
rect 930 390 970 430
rect 1030 390 1070 430
rect 930 370 1070 390
rect 930 330 970 370
rect 1030 330 1070 370
rect 930 310 1070 330
rect 930 270 970 310
rect 1030 270 1070 310
rect 930 250 1070 270
rect 930 210 970 250
rect 1030 210 1070 250
rect 930 190 1070 210
rect 930 150 970 190
rect 1030 150 1070 190
rect 930 110 1070 150
rect 1170 1090 1310 1110
rect 1170 1050 1210 1090
rect 1270 1050 1310 1090
rect 1170 1030 1310 1050
rect 1170 990 1210 1030
rect 1270 990 1310 1030
rect 1170 970 1310 990
rect 1170 930 1210 970
rect 1270 930 1310 970
rect 1170 910 1310 930
rect 1170 870 1210 910
rect 1270 870 1310 910
rect 1170 850 1310 870
rect 1170 810 1210 850
rect 1270 810 1310 850
rect 1170 790 1310 810
rect 1170 750 1210 790
rect 1270 750 1310 790
rect 1170 730 1310 750
rect 1170 690 1210 730
rect 1270 690 1310 730
rect 1170 670 1310 690
rect 1170 630 1210 670
rect 1270 630 1310 670
rect 1170 610 1310 630
rect 1170 570 1210 610
rect 1270 570 1310 610
rect 1170 550 1310 570
rect 1170 510 1210 550
rect 1270 510 1310 550
rect 1170 490 1310 510
rect 1170 450 1210 490
rect 1270 450 1310 490
rect 1170 430 1310 450
rect 1170 390 1210 430
rect 1270 390 1310 430
rect 1170 370 1310 390
rect 1170 330 1210 370
rect 1270 330 1310 370
rect 1170 310 1310 330
rect 1170 270 1210 310
rect 1270 270 1310 310
rect 1170 250 1310 270
rect 1170 210 1210 250
rect 1270 210 1310 250
rect 1170 190 1310 210
rect 1170 150 1210 190
rect 1270 150 1310 190
rect 1170 10 1310 150
rect 1660 1090 1800 1110
rect 1660 1050 1700 1090
rect 1760 1050 1800 1090
rect 1660 1030 1800 1050
rect 1660 990 1700 1030
rect 1760 990 1800 1030
rect 1660 970 1800 990
rect 1660 930 1700 970
rect 1760 930 1800 970
rect 1660 910 1800 930
rect 1660 870 1700 910
rect 1760 870 1800 910
rect 1660 850 1800 870
rect 1660 810 1700 850
rect 1760 810 1800 850
rect 1660 790 1800 810
rect 1660 750 1700 790
rect 1760 750 1800 790
rect 1660 730 1800 750
rect 1660 690 1700 730
rect 1760 690 1800 730
rect 1660 670 1800 690
rect 1660 630 1700 670
rect 1760 630 1800 670
rect 1660 610 1800 630
rect 1660 570 1700 610
rect 1760 570 1800 610
rect 1660 550 1800 570
rect 1660 510 1700 550
rect 1760 510 1800 550
rect 1660 490 1800 510
rect 1660 450 1700 490
rect 1760 450 1800 490
rect 1660 430 1800 450
rect 1660 390 1700 430
rect 1760 390 1800 430
rect 1660 370 1800 390
rect 1660 330 1700 370
rect 1760 330 1800 370
rect 1660 310 1800 330
rect 1660 270 1700 310
rect 1760 270 1800 310
rect 1660 250 1800 270
rect 1660 210 1700 250
rect 1760 210 1800 250
rect 1660 190 1800 210
rect 1660 150 1700 190
rect 1760 150 1800 190
rect 1660 10 1800 150
rect 1900 1090 2040 1150
rect 1900 1050 1940 1090
rect 2000 1050 2040 1090
rect 1900 1030 2040 1050
rect 1900 990 1940 1030
rect 2000 990 2040 1030
rect 1900 970 2040 990
rect 1900 930 1940 970
rect 2000 930 2040 970
rect 1900 910 2040 930
rect 1900 870 1940 910
rect 2000 870 2040 910
rect 1900 850 2040 870
rect 1900 810 1940 850
rect 2000 810 2040 850
rect 1900 790 2040 810
rect 1900 750 1940 790
rect 2000 750 2040 790
rect 1900 730 2040 750
rect 1900 690 1940 730
rect 2000 690 2040 730
rect 1900 670 2040 690
rect 1900 630 1940 670
rect 2000 630 2040 670
rect 1900 610 2040 630
rect 1900 570 1940 610
rect 2000 570 2040 610
rect 1900 550 2040 570
rect 1900 510 1940 550
rect 2000 510 2040 550
rect 1900 490 2040 510
rect 1900 450 1940 490
rect 2000 450 2040 490
rect 1900 430 2040 450
rect 1900 390 1940 430
rect 2000 390 2040 430
rect 1900 370 2040 390
rect 1900 330 1940 370
rect 2000 330 2040 370
rect 1900 310 2040 330
rect 1900 270 1940 310
rect 2000 270 2040 310
rect 1900 250 2040 270
rect 1900 210 1940 250
rect 2000 210 2040 250
rect 1900 190 2040 210
rect 1900 150 1940 190
rect 2000 150 2040 190
rect 1900 110 2040 150
rect 2140 1090 2280 1110
rect 2140 1050 2180 1090
rect 2240 1050 2280 1090
rect 2140 1030 2280 1050
rect 2140 990 2180 1030
rect 2240 990 2280 1030
rect 2140 970 2280 990
rect 2140 930 2180 970
rect 2240 930 2280 970
rect 2140 910 2280 930
rect 2140 870 2180 910
rect 2240 870 2280 910
rect 2140 850 2280 870
rect 2140 810 2180 850
rect 2240 810 2280 850
rect 2140 790 2280 810
rect 2140 750 2180 790
rect 2240 750 2280 790
rect 2140 730 2280 750
rect 2140 690 2180 730
rect 2240 690 2280 730
rect 2140 670 2280 690
rect 2140 630 2180 670
rect 2240 630 2280 670
rect 2140 610 2280 630
rect 2140 570 2180 610
rect 2240 570 2280 610
rect 2140 550 2280 570
rect 2140 510 2180 550
rect 2240 510 2280 550
rect 2140 490 2280 510
rect 2140 450 2180 490
rect 2240 450 2280 490
rect 2140 430 2280 450
rect 2140 390 2180 430
rect 2240 390 2280 430
rect 2140 370 2280 390
rect 2140 330 2180 370
rect 2240 330 2280 370
rect 2140 310 2280 330
rect 2140 270 2180 310
rect 2240 270 2280 310
rect 2140 250 2280 270
rect 2140 210 2180 250
rect 2240 210 2280 250
rect 2140 190 2280 210
rect 2140 150 2180 190
rect 2240 150 2280 190
rect 2140 10 2280 150
rect 2380 1090 2520 1150
rect 2380 1050 2420 1090
rect 2480 1050 2520 1090
rect 2380 1030 2520 1050
rect 2380 990 2420 1030
rect 2480 990 2520 1030
rect 2380 970 2520 990
rect 2380 930 2420 970
rect 2480 930 2520 970
rect 2380 910 2520 930
rect 2380 870 2420 910
rect 2480 870 2520 910
rect 2380 850 2520 870
rect 2380 810 2420 850
rect 2480 810 2520 850
rect 2380 790 2520 810
rect 2380 750 2420 790
rect 2480 750 2520 790
rect 2380 730 2520 750
rect 2380 690 2420 730
rect 2480 690 2520 730
rect 2380 670 2520 690
rect 2380 630 2420 670
rect 2480 630 2520 670
rect 2380 610 2520 630
rect 2380 570 2420 610
rect 2480 570 2520 610
rect 2380 550 2520 570
rect 2380 510 2420 550
rect 2480 510 2520 550
rect 2380 490 2520 510
rect 2380 450 2420 490
rect 2480 450 2520 490
rect 2380 430 2520 450
rect 2380 390 2420 430
rect 2480 390 2520 430
rect 2380 370 2520 390
rect 2380 330 2420 370
rect 2480 330 2520 370
rect 2380 310 2520 330
rect 2380 270 2420 310
rect 2480 270 2520 310
rect 2380 250 2520 270
rect 2380 210 2420 250
rect 2480 210 2520 250
rect 2380 190 2520 210
rect 2380 150 2420 190
rect 2480 150 2520 190
rect 2380 110 2520 150
rect 2630 1090 2770 1110
rect 2630 1050 2670 1090
rect 2730 1050 2770 1090
rect 2630 1030 2770 1050
rect 2630 990 2670 1030
rect 2730 990 2770 1030
rect 2630 970 2770 990
rect 2630 930 2670 970
rect 2730 930 2770 970
rect 2630 910 2770 930
rect 2630 870 2670 910
rect 2730 870 2770 910
rect 2630 850 2770 870
rect 2630 810 2670 850
rect 2730 810 2770 850
rect 2630 790 2770 810
rect 2630 750 2670 790
rect 2730 750 2770 790
rect 2630 730 2770 750
rect 2630 690 2670 730
rect 2730 690 2770 730
rect 2630 670 2770 690
rect 2630 630 2670 670
rect 2730 630 2770 670
rect 2630 610 2770 630
rect 2630 570 2670 610
rect 2730 570 2770 610
rect 2630 550 2770 570
rect 2630 510 2670 550
rect 2730 510 2770 550
rect 2630 490 2770 510
rect 2630 450 2670 490
rect 2730 450 2770 490
rect 2630 430 2770 450
rect 2630 390 2670 430
rect 2730 390 2770 430
rect 2630 370 2770 390
rect 2630 330 2670 370
rect 2730 330 2770 370
rect 2630 310 2770 330
rect 2630 270 2670 310
rect 2730 270 2770 310
rect 2630 250 2770 270
rect 2630 210 2670 250
rect 2730 210 2770 250
rect 2630 190 2770 210
rect 2630 150 2670 190
rect 2730 150 2770 190
rect 2630 10 2770 150
rect 2870 1090 3010 1150
rect 2870 1050 2900 1090
rect 2960 1050 3010 1090
rect 2870 1030 3010 1050
rect 2870 990 2900 1030
rect 2960 990 3010 1030
rect 2870 970 3010 990
rect 2870 930 2900 970
rect 2960 930 3010 970
rect 2870 910 3010 930
rect 2870 870 2900 910
rect 2960 870 3010 910
rect 2870 850 3010 870
rect 2870 810 2900 850
rect 2960 810 3010 850
rect 2870 790 3010 810
rect 2870 750 2900 790
rect 2960 750 3010 790
rect 2870 730 3010 750
rect 2870 690 2900 730
rect 2960 690 3010 730
rect 2870 670 3010 690
rect 2870 630 2900 670
rect 2960 630 3010 670
rect 2870 610 3010 630
rect 2870 570 2900 610
rect 2960 570 3010 610
rect 2870 550 3010 570
rect 2870 510 2900 550
rect 2960 510 3010 550
rect 2870 490 3010 510
rect 2870 450 2900 490
rect 2960 450 3010 490
rect 2870 430 3010 450
rect 2870 390 2900 430
rect 2960 390 3010 430
rect 2870 370 3010 390
rect 2870 330 2900 370
rect 2960 330 3010 370
rect 2870 310 3010 330
rect 2870 270 2900 310
rect 2960 270 3010 310
rect 2870 250 3010 270
rect 2870 210 2900 250
rect 2960 210 3010 250
rect 2870 190 3010 210
rect 2870 150 2900 190
rect 2960 150 3010 190
rect 2870 110 3010 150
rect 200 -90 2770 10
use sky130_fd_pr__pfet_01v8_1um_10um_mult2  sky130_fd_pr__pfet_01v8_1um_10um_mult2_0
timestamp 1658894429
transform 1 0 2430 0 1 0
box 0 0 539 1219
use sky130_fd_pr__pfet_01v8_1um_10um_mult10  sky130_fd_pr__pfet_01v8_1um_10um_mult10_0
timestamp 1658894606
transform 1 0 0 0 1 0
box 0 0 2483 1219
<< labels >>
rlabel metal2 1410 1220 1550 1250 1 IREF
rlabel metal3 200 -90 2770 10 1 VDD
rlabel metal3 -40 1150 3010 1210 1 IOUT
<< end >>
