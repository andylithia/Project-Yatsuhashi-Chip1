magic
tech sky130A
timestamp 1659151574
use OSC_5GHz_1  OSC_5GHz_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/OSC
timestamp 1659147692
transform 0 1 22200 -1 0 1500
box -2250 -4200 12500 6000
use lna_complete_1  lna_complete_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/LNA
timestamp 1659151574
transform -1 0 6050 0 -1 11730
box -15400 -13600 6050 11720
use lna_complete_1  lna_complete_1_1
timestamp 1659151574
transform 1 0 40400 0 -1 11730
box -15400 -13600 6050 11720
<< end >>
