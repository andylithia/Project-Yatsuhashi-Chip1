magic
tech sky130A
timestamp 1659502258
use MIXER_5G_complete  MIXER_5G_complete_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/MIXER
timestamp 1659501813
transform 1 0 4687 0 1 11510
box -4700 -11500 28800 15800
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501465
transform 1 0 3000 0 1 13850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_1
timestamp 1659501465
transform 1 0 2000 0 1 13850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_2
timestamp 1659501465
transform 1 0 0 0 1 12850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_3
timestamp 1659501465
transform 1 0 1000 0 1 12850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_4
timestamp 1659501465
transform 1 0 16000 0 1 6850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_5
timestamp 1659501465
transform 1 0 18000 0 1 4850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_6
timestamp 1659501465
transform 1 0 20000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_7
timestamp 1659501465
transform 1 0 21000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_8
timestamp 1659501465
transform 1 0 22000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_9
timestamp 1659501465
transform 1 0 23000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_10
timestamp 1659501465
transform 1 0 24000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_11
timestamp 1659501465
transform 1 0 25000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_12
timestamp 1659501465
transform 1 0 26000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_13
timestamp 1659501465
transform 1 0 27000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_14
timestamp 1659501465
transform 1 0 28000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_15
timestamp 1659501465
transform 1 0 29000 0 1 2850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_16
timestamp 1659501465
transform 1 0 31000 0 1 4850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_17
timestamp 1659501465
transform 1 0 33000 0 1 6850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_18
timestamp 1659501465
transform 1 0 35000 0 1 8850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_19
timestamp 1659501465
transform 1 0 35000 0 1 19850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_20
timestamp 1659501465
transform 1 0 35000 0 1 18850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_21
timestamp 1659501465
transform 1 0 35000 0 1 17850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_22
timestamp 1659501465
transform 1 0 35000 0 1 16850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_23
timestamp 1659501465
transform 1 0 35000 0 1 15850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_24
timestamp 1659501465
transform 1 0 35000 0 1 14850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_25
timestamp 1659501465
transform 1 0 35000 0 1 13850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_26
timestamp 1659501465
transform 1 0 35000 0 1 12850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_27
timestamp 1659501465
transform 1 0 35000 0 1 11850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_28
timestamp 1659501465
transform 1 0 35000 0 1 10850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_29
timestamp 1659501465
transform 1 0 35000 0 1 9850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_30
timestamp 1659501465
transform 1 0 34000 0 1 19850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_31
timestamp 1659501465
transform 1 0 33000 0 1 20850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_32
timestamp 1659501465
transform 1 0 33000 0 1 21850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_33
timestamp 1659501465
transform 1 0 32000 0 1 21850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_34
timestamp 1659501465
transform 1 0 31000 0 1 22850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_35
timestamp 1659501465
transform 1 0 31000 0 1 23850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_36
timestamp 1659501465
transform 1 0 30000 0 1 23850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_37
timestamp 1659501465
transform 1 0 18000 0 1 23850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_38
timestamp 1659501465
transform 1 0 16000 0 1 21850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_39
timestamp 1659501465
transform 1 0 13000 0 1 25850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_40
timestamp 1659501465
transform 1 0 12000 0 1 26850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_41
timestamp 1659501465
transform 1 0 11000 0 1 27850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_42
timestamp 1659501465
transform 1 0 12000 0 1 27850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_43
timestamp 1659501465
transform 1 0 13000 0 1 27850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_44
timestamp 1659501465
transform 1 0 13000 0 1 26850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_45
timestamp 1659501465
transform 1 0 13000 0 1 850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_46
timestamp 1659501465
transform 1 0 12000 0 1 850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_47
timestamp 1659501465
transform 1 0 11000 0 1 -150
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_48
timestamp 1659501465
transform 1 0 10000 0 1 -1150
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_49
timestamp 1659501465
transform 1 0 11000 0 1 -1150
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_50
timestamp 1659501465
transform 1 0 12000 0 1 -1150
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_51
timestamp 1659501465
transform 1 0 13000 0 1 -1150
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_52
timestamp 1659501465
transform 1 0 12000 0 1 -150
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_53
timestamp 1659501465
transform 1 0 13000 0 1 -150
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_54
timestamp 1659501465
transform 1 0 13000 0 1 1850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_55
timestamp 1659501465
transform 1 0 -21000 0 1 3850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_56
timestamp 1659501465
transform 1 0 14000 0 1 10850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_57
timestamp 1659501465
transform 1 0 15000 0 1 10850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_58
timestamp 1659501465
transform 1 0 13000 0 1 10850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_59
timestamp 1659501465
transform 1 0 12000 0 1 10850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_60
timestamp 1659501465
transform 1 0 13000 0 1 9850
box 0 -850 1000 150
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_61
timestamp 1659501465
transform 1 0 12000 0 1 16850
box 0 -850 1000 150
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501637
transform 1 0 0 0 1 13000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_1
timestamp 1659501637
transform 1 0 13000 0 1 16000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_2
timestamp 1659501637
transform 1 0 14000 0 1 18000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_3
timestamp 1659501637
transform 1 0 14000 0 1 20000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_4
timestamp 1659501637
transform 1 0 14000 0 1 22000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_5
timestamp 1659501637
transform 1 0 14000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_6
timestamp 1659501637
transform 1 0 14000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_7
timestamp 1659501637
transform 1 0 16000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_8
timestamp 1659501637
transform 1 0 16000 0 1 22000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_9
timestamp 1659501637
transform 1 0 16000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_10
timestamp 1659501637
transform 1 0 18000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_11
timestamp 1659501637
transform 1 0 18000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_12
timestamp 1659501637
transform 1 0 20000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_13
timestamp 1659501637
transform 1 0 20000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_14
timestamp 1659501637
transform 1 0 22000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_15
timestamp 1659501637
transform 1 0 24000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_16
timestamp 1659501637
transform 1 0 26000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_17
timestamp 1659501637
transform 1 0 22000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_18
timestamp 1659501637
transform 1 0 24000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_19
timestamp 1659501637
transform 1 0 26000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_20
timestamp 1659501637
transform 1 0 28000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_21
timestamp 1659501637
transform 1 0 28000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_22
timestamp 1659501637
transform 1 0 14000 0 1 6000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_23
timestamp 1659501637
transform 1 0 14000 0 1 4000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_24
timestamp 1659501637
transform 1 0 14000 0 1 2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_25
timestamp 1659501637
transform 1 0 14000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_26
timestamp 1659501637
transform 1 0 16000 0 1 2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_27
timestamp 1659501637
transform 1 0 16000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_28
timestamp 1659501637
transform 1 0 14000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_29
timestamp 1659501637
transform 1 0 16000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_30
timestamp 1659501637
transform 1 0 18000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_31
timestamp 1659501637
transform 1 0 20000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_32
timestamp 1659501637
transform 1 0 22000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_33
timestamp 1659501637
transform 1 0 24000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_34
timestamp 1659501637
transform 1 0 26000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_35
timestamp 1659501637
transform 1 0 28000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_36
timestamp 1659501637
transform 1 0 30000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_37
timestamp 1659501637
transform 1 0 32000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_38
timestamp 1659501637
transform 1 0 34000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_39
timestamp 1659501637
transform 1 0 30000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_40
timestamp 1659501637
transform 1 0 32000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_41
timestamp 1659501637
transform 1 0 34000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_42
timestamp 1659501637
transform 1 0 36000 0 1 24000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_43
timestamp 1659501637
transform 1 0 36000 0 1 -2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_44
timestamp 1659501637
transform 1 0 36000 0 1 22000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_45
timestamp 1659501637
transform 1 0 36000 0 1 20000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_46
timestamp 1659501637
transform 1 0 36000 0 1 18000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_47
timestamp 1659501637
transform 1 0 36000 0 1 16000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_48
timestamp 1659501637
transform 1 0 36000 0 1 14000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_49
timestamp 1659501637
transform 1 0 36000 0 1 12000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_50
timestamp 1659501637
transform 1 0 36000 0 1 10000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_51
timestamp 1659501637
transform 1 0 36000 0 1 8000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_52
timestamp 1659501637
transform 1 0 36000 0 1 6000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_53
timestamp 1659501637
transform 1 0 36000 0 1 4000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_54
timestamp 1659501637
transform 1 0 34000 0 1 4000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_55
timestamp 1659501637
transform 1 0 34000 0 1 22000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_56
timestamp 1659501637
transform 1 0 34000 0 1 20000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_57
timestamp 1659501637
transform 1 0 32000 0 1 22000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_58
timestamp 1659501637
transform 1 0 34000 0 1 6000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_59
timestamp 1659501637
transform 1 0 32000 0 1 4000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_60
timestamp 1659501637
transform 1 0 30000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_61
timestamp 1659501637
transform 1 0 32000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_62
timestamp 1659501637
transform 1 0 34000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_63
timestamp 1659501637
transform 1 0 36000 0 1 26000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_64
timestamp 1659501637
transform 1 0 16000 0 1 4000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_65
timestamp 1659501637
transform 1 0 18000 0 1 2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_66
timestamp 1659501637
transform 1 0 18000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_67
timestamp 1659501637
transform 1 0 20000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_68
timestamp 1659501637
transform 1 0 22000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_69
timestamp 1659501637
transform 1 0 24000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_70
timestamp 1659501637
transform 1 0 26000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_71
timestamp 1659501637
transform 1 0 28000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_72
timestamp 1659501637
transform 1 0 30000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_73
timestamp 1659501637
transform 1 0 32000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_74
timestamp 1659501637
transform 1 0 34000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_75
timestamp 1659501637
transform 1 0 36000 0 1 0
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_76
timestamp 1659501637
transform 1 0 32000 0 1 2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_77
timestamp 1659501637
transform 1 0 34000 0 1 2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_78
timestamp 1659501637
transform 1 0 36000 0 1 2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_79
timestamp 1659501637
transform 1 0 30000 0 1 2000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_80
timestamp 1659501637
transform 1 0 14000 0 1 8000
box 0 0 2000 2000
<< end >>
