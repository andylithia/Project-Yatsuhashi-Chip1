magic
tech sky130B
timestamp 1660792292
<< metal1 >>
rect 0 3990 4000 4000
rect 0 3955 75 3990
rect 175 3955 325 3990
rect 425 3955 575 3990
rect 675 3955 825 3990
rect 925 3955 1075 3990
rect 1175 3955 1325 3990
rect 1425 3955 1575 3990
rect 1675 3955 1825 3990
rect 1925 3955 2075 3990
rect 2175 3955 2325 3990
rect 2425 3955 2575 3990
rect 2675 3955 2825 3990
rect 2925 3955 3075 3990
rect 3175 3955 3325 3990
rect 3425 3955 3575 3990
rect 3675 3955 3825 3990
rect 3925 3955 4000 3990
rect 0 3950 4000 3955
rect 0 3940 60 3950
rect 190 3940 310 3950
rect 440 3940 560 3950
rect 690 3940 810 3950
rect 940 3940 1060 3950
rect 1190 3940 1310 3950
rect 1440 3940 1560 3950
rect 1690 3940 1810 3950
rect 1940 3940 2060 3950
rect 2190 3940 2310 3950
rect 2440 3940 2560 3950
rect 2690 3940 2810 3950
rect 2940 3940 3060 3950
rect 3190 3940 3310 3950
rect 3440 3940 3560 3950
rect 3690 3940 3810 3950
rect 3940 3940 4000 3950
rect 0 3925 50 3940
rect 0 3825 10 3925
rect 45 3825 50 3925
rect 0 3810 50 3825
rect 200 3925 300 3940
rect 200 3825 205 3925
rect 240 3825 260 3925
rect 295 3825 300 3925
rect 200 3810 300 3825
rect 450 3925 550 3940
rect 450 3825 455 3925
rect 490 3825 510 3925
rect 545 3825 550 3925
rect 450 3810 550 3825
rect 700 3925 800 3940
rect 700 3825 705 3925
rect 740 3825 760 3925
rect 795 3825 800 3925
rect 700 3810 800 3825
rect 950 3925 1050 3940
rect 950 3825 955 3925
rect 990 3825 1010 3925
rect 1045 3825 1050 3925
rect 950 3810 1050 3825
rect 1200 3925 1300 3940
rect 1200 3825 1205 3925
rect 1240 3825 1260 3925
rect 1295 3825 1300 3925
rect 1200 3810 1300 3825
rect 1450 3925 1550 3940
rect 1450 3825 1455 3925
rect 1490 3825 1510 3925
rect 1545 3825 1550 3925
rect 1450 3810 1550 3825
rect 1700 3925 1800 3940
rect 1700 3825 1705 3925
rect 1740 3825 1760 3925
rect 1795 3825 1800 3925
rect 1700 3810 1800 3825
rect 1950 3925 2050 3940
rect 1950 3825 1955 3925
rect 1990 3825 2010 3925
rect 2045 3825 2050 3925
rect 1950 3810 2050 3825
rect 2200 3925 2300 3940
rect 2200 3825 2205 3925
rect 2240 3825 2260 3925
rect 2295 3825 2300 3925
rect 2200 3810 2300 3825
rect 2450 3925 2550 3940
rect 2450 3825 2455 3925
rect 2490 3825 2510 3925
rect 2545 3825 2550 3925
rect 2450 3810 2550 3825
rect 2700 3925 2800 3940
rect 2700 3825 2705 3925
rect 2740 3825 2760 3925
rect 2795 3825 2800 3925
rect 2700 3810 2800 3825
rect 2950 3925 3050 3940
rect 2950 3825 2955 3925
rect 2990 3825 3010 3925
rect 3045 3825 3050 3925
rect 2950 3810 3050 3825
rect 3200 3925 3300 3940
rect 3200 3825 3205 3925
rect 3240 3825 3260 3925
rect 3295 3825 3300 3925
rect 3200 3810 3300 3825
rect 3450 3925 3550 3940
rect 3450 3825 3455 3925
rect 3490 3825 3510 3925
rect 3545 3825 3550 3925
rect 3450 3810 3550 3825
rect 3700 3925 3800 3940
rect 3700 3825 3705 3925
rect 3740 3825 3760 3925
rect 3795 3825 3800 3925
rect 3700 3810 3800 3825
rect 3950 3925 4000 3940
rect 3950 3825 3955 3925
rect 3990 3825 4000 3925
rect 3950 3810 4000 3825
rect 0 3800 60 3810
rect 190 3800 310 3810
rect 440 3800 560 3810
rect 690 3800 810 3810
rect 940 3800 1060 3810
rect 1190 3800 1310 3810
rect 1440 3800 1560 3810
rect 1690 3800 1810 3810
rect 1940 3800 2060 3810
rect 2190 3800 2310 3810
rect 2440 3800 2560 3810
rect 2690 3800 2810 3810
rect 2940 3800 3060 3810
rect 3190 3800 3310 3810
rect 3440 3800 3560 3810
rect 3690 3800 3810 3810
rect 3940 3800 4000 3810
rect 0 3795 4000 3800
rect 0 3760 75 3795
rect 175 3760 325 3795
rect 425 3760 575 3795
rect 675 3760 825 3795
rect 925 3760 1075 3795
rect 1175 3760 1325 3795
rect 1425 3760 1575 3795
rect 1675 3760 1825 3795
rect 1925 3760 2075 3795
rect 2175 3760 2325 3795
rect 2425 3760 2575 3795
rect 2675 3760 2825 3795
rect 2925 3760 3075 3795
rect 3175 3760 3325 3795
rect 3425 3760 3575 3795
rect 3675 3760 3825 3795
rect 3925 3760 4000 3795
rect 0 3740 4000 3760
rect 0 3705 75 3740
rect 175 3705 325 3740
rect 425 3705 575 3740
rect 675 3705 825 3740
rect 925 3705 1075 3740
rect 1175 3705 1325 3740
rect 1425 3705 1575 3740
rect 1675 3705 1825 3740
rect 1925 3705 2075 3740
rect 2175 3705 2325 3740
rect 2425 3705 2575 3740
rect 2675 3705 2825 3740
rect 2925 3705 3075 3740
rect 3175 3705 3325 3740
rect 3425 3705 3575 3740
rect 3675 3705 3825 3740
rect 3925 3705 4000 3740
rect 0 3700 4000 3705
rect 0 3690 60 3700
rect 190 3690 310 3700
rect 440 3690 560 3700
rect 690 3690 810 3700
rect 940 3690 1060 3700
rect 1190 3690 1310 3700
rect 1440 3690 1560 3700
rect 1690 3690 1810 3700
rect 1940 3690 2060 3700
rect 2190 3690 2310 3700
rect 2440 3690 2560 3700
rect 2690 3690 2810 3700
rect 2940 3690 3060 3700
rect 3190 3690 3310 3700
rect 3440 3690 3560 3700
rect 3690 3690 3810 3700
rect 3940 3690 4000 3700
rect 0 3675 50 3690
rect 0 3575 10 3675
rect 45 3575 50 3675
rect 0 3560 50 3575
rect 200 3675 300 3690
rect 200 3575 205 3675
rect 240 3575 260 3675
rect 295 3575 300 3675
rect 200 3560 300 3575
rect 450 3675 550 3690
rect 450 3575 455 3675
rect 490 3575 510 3675
rect 545 3575 550 3675
rect 450 3560 550 3575
rect 700 3675 800 3690
rect 700 3575 705 3675
rect 740 3575 760 3675
rect 795 3575 800 3675
rect 700 3560 800 3575
rect 950 3675 1050 3690
rect 950 3575 955 3675
rect 990 3575 1010 3675
rect 1045 3575 1050 3675
rect 950 3560 1050 3575
rect 1200 3675 1300 3690
rect 1200 3575 1205 3675
rect 1240 3575 1260 3675
rect 1295 3575 1300 3675
rect 1200 3560 1300 3575
rect 1450 3675 1550 3690
rect 1450 3575 1455 3675
rect 1490 3575 1510 3675
rect 1545 3575 1550 3675
rect 1450 3560 1550 3575
rect 1700 3675 1800 3690
rect 1700 3575 1705 3675
rect 1740 3575 1760 3675
rect 1795 3575 1800 3675
rect 1700 3560 1800 3575
rect 1950 3675 2050 3690
rect 1950 3575 1955 3675
rect 1990 3575 2010 3675
rect 2045 3575 2050 3675
rect 1950 3560 2050 3575
rect 2200 3675 2300 3690
rect 2200 3575 2205 3675
rect 2240 3575 2260 3675
rect 2295 3575 2300 3675
rect 2200 3560 2300 3575
rect 2450 3675 2550 3690
rect 2450 3575 2455 3675
rect 2490 3575 2510 3675
rect 2545 3575 2550 3675
rect 2450 3560 2550 3575
rect 2700 3675 2800 3690
rect 2700 3575 2705 3675
rect 2740 3575 2760 3675
rect 2795 3575 2800 3675
rect 2700 3560 2800 3575
rect 2950 3675 3050 3690
rect 2950 3575 2955 3675
rect 2990 3575 3010 3675
rect 3045 3575 3050 3675
rect 2950 3560 3050 3575
rect 3200 3675 3300 3690
rect 3200 3575 3205 3675
rect 3240 3575 3260 3675
rect 3295 3575 3300 3675
rect 3200 3560 3300 3575
rect 3450 3675 3550 3690
rect 3450 3575 3455 3675
rect 3490 3575 3510 3675
rect 3545 3575 3550 3675
rect 3450 3560 3550 3575
rect 3700 3675 3800 3690
rect 3700 3575 3705 3675
rect 3740 3575 3760 3675
rect 3795 3575 3800 3675
rect 3700 3560 3800 3575
rect 3950 3675 4000 3690
rect 3950 3575 3955 3675
rect 3990 3575 4000 3675
rect 3950 3560 4000 3575
rect 0 3550 60 3560
rect 190 3550 310 3560
rect 440 3550 560 3560
rect 690 3550 810 3560
rect 940 3550 1060 3560
rect 1190 3550 1310 3560
rect 1440 3550 1560 3560
rect 1690 3550 1810 3560
rect 1940 3550 2060 3560
rect 2190 3550 2310 3560
rect 2440 3550 2560 3560
rect 2690 3550 2810 3560
rect 2940 3550 3060 3560
rect 3190 3550 3310 3560
rect 3440 3550 3560 3560
rect 3690 3550 3810 3560
rect 3940 3550 4000 3560
rect 0 3545 4000 3550
rect 0 3510 75 3545
rect 175 3510 325 3545
rect 425 3510 575 3545
rect 675 3510 825 3545
rect 925 3510 1075 3545
rect 1175 3510 1325 3545
rect 1425 3510 1575 3545
rect 1675 3510 1825 3545
rect 1925 3510 2075 3545
rect 2175 3510 2325 3545
rect 2425 3510 2575 3545
rect 2675 3510 2825 3545
rect 2925 3510 3075 3545
rect 3175 3510 3325 3545
rect 3425 3510 3575 3545
rect 3675 3510 3825 3545
rect 3925 3510 4000 3545
rect 0 3490 4000 3510
rect 0 3455 75 3490
rect 175 3455 325 3490
rect 425 3455 575 3490
rect 675 3455 825 3490
rect 925 3455 1075 3490
rect 1175 3455 1325 3490
rect 1425 3455 1575 3490
rect 1675 3455 1825 3490
rect 1925 3455 2075 3490
rect 2175 3455 2325 3490
rect 2425 3455 2575 3490
rect 2675 3455 2825 3490
rect 2925 3455 3075 3490
rect 3175 3455 3325 3490
rect 3425 3455 3575 3490
rect 3675 3455 3825 3490
rect 3925 3455 4000 3490
rect 0 3450 4000 3455
rect 0 3440 60 3450
rect 190 3440 310 3450
rect 440 3440 560 3450
rect 690 3440 810 3450
rect 940 3440 1060 3450
rect 1190 3440 1310 3450
rect 1440 3440 1560 3450
rect 1690 3440 1810 3450
rect 1940 3440 2060 3450
rect 2190 3440 2310 3450
rect 2440 3440 2560 3450
rect 2690 3440 2810 3450
rect 2940 3440 3060 3450
rect 3190 3440 3310 3450
rect 3440 3440 3560 3450
rect 3690 3440 3810 3450
rect 3940 3440 4000 3450
rect 0 3425 50 3440
rect 0 3325 10 3425
rect 45 3325 50 3425
rect 0 3310 50 3325
rect 200 3425 300 3440
rect 200 3325 205 3425
rect 240 3325 260 3425
rect 295 3325 300 3425
rect 200 3310 300 3325
rect 450 3425 550 3440
rect 450 3325 455 3425
rect 490 3325 510 3425
rect 545 3325 550 3425
rect 450 3310 550 3325
rect 700 3425 800 3440
rect 700 3325 705 3425
rect 740 3325 760 3425
rect 795 3325 800 3425
rect 700 3310 800 3325
rect 950 3425 1050 3440
rect 950 3325 955 3425
rect 990 3325 1010 3425
rect 1045 3325 1050 3425
rect 950 3310 1050 3325
rect 1200 3425 1300 3440
rect 1200 3325 1205 3425
rect 1240 3325 1260 3425
rect 1295 3325 1300 3425
rect 1200 3310 1300 3325
rect 1450 3425 1550 3440
rect 1450 3325 1455 3425
rect 1490 3325 1510 3425
rect 1545 3325 1550 3425
rect 1450 3310 1550 3325
rect 1700 3425 1800 3440
rect 1700 3325 1705 3425
rect 1740 3325 1760 3425
rect 1795 3325 1800 3425
rect 1700 3310 1800 3325
rect 1950 3425 2050 3440
rect 1950 3325 1955 3425
rect 1990 3325 2010 3425
rect 2045 3325 2050 3425
rect 1950 3310 2050 3325
rect 2200 3425 2300 3440
rect 2200 3325 2205 3425
rect 2240 3325 2260 3425
rect 2295 3325 2300 3425
rect 2200 3310 2300 3325
rect 2450 3425 2550 3440
rect 2450 3325 2455 3425
rect 2490 3325 2510 3425
rect 2545 3325 2550 3425
rect 2450 3310 2550 3325
rect 2700 3425 2800 3440
rect 2700 3325 2705 3425
rect 2740 3325 2760 3425
rect 2795 3325 2800 3425
rect 2700 3310 2800 3325
rect 2950 3425 3050 3440
rect 2950 3325 2955 3425
rect 2990 3325 3010 3425
rect 3045 3325 3050 3425
rect 2950 3310 3050 3325
rect 3200 3425 3300 3440
rect 3200 3325 3205 3425
rect 3240 3325 3260 3425
rect 3295 3325 3300 3425
rect 3200 3310 3300 3325
rect 3450 3425 3550 3440
rect 3450 3325 3455 3425
rect 3490 3325 3510 3425
rect 3545 3325 3550 3425
rect 3450 3310 3550 3325
rect 3700 3425 3800 3440
rect 3700 3325 3705 3425
rect 3740 3325 3760 3425
rect 3795 3325 3800 3425
rect 3700 3310 3800 3325
rect 3950 3425 4000 3440
rect 3950 3325 3955 3425
rect 3990 3325 4000 3425
rect 3950 3310 4000 3325
rect 0 3300 60 3310
rect 190 3300 310 3310
rect 440 3300 560 3310
rect 690 3300 810 3310
rect 940 3300 1060 3310
rect 1190 3300 1310 3310
rect 1440 3300 1560 3310
rect 1690 3300 1810 3310
rect 1940 3300 2060 3310
rect 2190 3300 2310 3310
rect 2440 3300 2560 3310
rect 2690 3300 2810 3310
rect 2940 3300 3060 3310
rect 3190 3300 3310 3310
rect 3440 3300 3560 3310
rect 3690 3300 3810 3310
rect 3940 3300 4000 3310
rect 0 3295 4000 3300
rect 0 3260 75 3295
rect 175 3260 325 3295
rect 425 3260 575 3295
rect 675 3260 825 3295
rect 925 3260 1075 3295
rect 1175 3260 1325 3295
rect 1425 3260 1575 3295
rect 1675 3260 1825 3295
rect 1925 3260 2075 3295
rect 2175 3260 2325 3295
rect 2425 3260 2575 3295
rect 2675 3260 2825 3295
rect 2925 3260 3075 3295
rect 3175 3260 3325 3295
rect 3425 3260 3575 3295
rect 3675 3260 3825 3295
rect 3925 3260 4000 3295
rect 0 3240 4000 3260
rect 0 3205 75 3240
rect 175 3205 325 3240
rect 425 3205 575 3240
rect 675 3205 825 3240
rect 925 3205 1075 3240
rect 1175 3205 1325 3240
rect 1425 3205 1575 3240
rect 1675 3205 1825 3240
rect 1925 3205 2075 3240
rect 2175 3205 2325 3240
rect 2425 3205 2575 3240
rect 2675 3205 2825 3240
rect 2925 3205 3075 3240
rect 3175 3205 3325 3240
rect 3425 3205 3575 3240
rect 3675 3205 3825 3240
rect 3925 3205 4000 3240
rect 0 3200 4000 3205
rect 0 3190 60 3200
rect 190 3190 310 3200
rect 440 3190 560 3200
rect 690 3190 810 3200
rect 940 3190 1060 3200
rect 1190 3190 1310 3200
rect 1440 3190 1560 3200
rect 1690 3190 1810 3200
rect 1940 3190 2060 3200
rect 2190 3190 2310 3200
rect 2440 3190 2560 3200
rect 2690 3190 2810 3200
rect 2940 3190 3060 3200
rect 3190 3190 3310 3200
rect 3440 3190 3560 3200
rect 3690 3190 3810 3200
rect 3940 3190 4000 3200
rect 0 3175 50 3190
rect 0 3075 10 3175
rect 45 3075 50 3175
rect 0 3060 50 3075
rect 200 3175 300 3190
rect 200 3075 205 3175
rect 240 3075 260 3175
rect 295 3075 300 3175
rect 200 3060 300 3075
rect 450 3175 550 3190
rect 450 3075 455 3175
rect 490 3075 510 3175
rect 545 3075 550 3175
rect 450 3060 550 3075
rect 700 3175 800 3190
rect 700 3075 705 3175
rect 740 3075 760 3175
rect 795 3075 800 3175
rect 700 3060 800 3075
rect 950 3175 1050 3190
rect 950 3075 955 3175
rect 990 3075 1010 3175
rect 1045 3075 1050 3175
rect 950 3060 1050 3075
rect 1200 3175 1300 3190
rect 1200 3075 1205 3175
rect 1240 3075 1260 3175
rect 1295 3075 1300 3175
rect 1200 3060 1300 3075
rect 1450 3175 1550 3190
rect 1450 3075 1455 3175
rect 1490 3075 1510 3175
rect 1545 3075 1550 3175
rect 1450 3060 1550 3075
rect 1700 3175 1800 3190
rect 1700 3075 1705 3175
rect 1740 3075 1760 3175
rect 1795 3075 1800 3175
rect 1700 3060 1800 3075
rect 1950 3175 2050 3190
rect 1950 3075 1955 3175
rect 1990 3075 2010 3175
rect 2045 3075 2050 3175
rect 1950 3060 2050 3075
rect 2200 3175 2300 3190
rect 2200 3075 2205 3175
rect 2240 3075 2260 3175
rect 2295 3075 2300 3175
rect 2200 3060 2300 3075
rect 2450 3175 2550 3190
rect 2450 3075 2455 3175
rect 2490 3075 2510 3175
rect 2545 3075 2550 3175
rect 2450 3060 2550 3075
rect 2700 3175 2800 3190
rect 2700 3075 2705 3175
rect 2740 3075 2760 3175
rect 2795 3075 2800 3175
rect 2700 3060 2800 3075
rect 2950 3175 3050 3190
rect 2950 3075 2955 3175
rect 2990 3075 3010 3175
rect 3045 3075 3050 3175
rect 2950 3060 3050 3075
rect 3200 3175 3300 3190
rect 3200 3075 3205 3175
rect 3240 3075 3260 3175
rect 3295 3075 3300 3175
rect 3200 3060 3300 3075
rect 3450 3175 3550 3190
rect 3450 3075 3455 3175
rect 3490 3075 3510 3175
rect 3545 3075 3550 3175
rect 3450 3060 3550 3075
rect 3700 3175 3800 3190
rect 3700 3075 3705 3175
rect 3740 3075 3760 3175
rect 3795 3075 3800 3175
rect 3700 3060 3800 3075
rect 3950 3175 4000 3190
rect 3950 3075 3955 3175
rect 3990 3075 4000 3175
rect 3950 3060 4000 3075
rect 0 3050 60 3060
rect 190 3050 310 3060
rect 440 3050 560 3060
rect 690 3050 810 3060
rect 940 3050 1060 3060
rect 1190 3050 1310 3060
rect 1440 3050 1560 3060
rect 1690 3050 1810 3060
rect 1940 3050 2060 3060
rect 2190 3050 2310 3060
rect 2440 3050 2560 3060
rect 2690 3050 2810 3060
rect 2940 3050 3060 3060
rect 3190 3050 3310 3060
rect 3440 3050 3560 3060
rect 3690 3050 3810 3060
rect 3940 3050 4000 3060
rect 0 3045 4000 3050
rect 0 3010 75 3045
rect 175 3010 325 3045
rect 425 3010 575 3045
rect 675 3010 825 3045
rect 925 3010 1075 3045
rect 1175 3010 1325 3045
rect 1425 3010 1575 3045
rect 1675 3010 1825 3045
rect 1925 3010 2075 3045
rect 2175 3010 2325 3045
rect 2425 3010 2575 3045
rect 2675 3010 2825 3045
rect 2925 3010 3075 3045
rect 3175 3010 3325 3045
rect 3425 3010 3575 3045
rect 3675 3010 3825 3045
rect 3925 3010 4000 3045
rect 0 2990 4000 3010
rect 0 2955 75 2990
rect 175 2955 325 2990
rect 425 2955 575 2990
rect 675 2955 825 2990
rect 925 2955 1075 2990
rect 1175 2955 1325 2990
rect 1425 2955 1575 2990
rect 1675 2955 1825 2990
rect 1925 2955 2075 2990
rect 2175 2955 2325 2990
rect 2425 2955 2575 2990
rect 2675 2955 2825 2990
rect 2925 2955 3075 2990
rect 3175 2955 3325 2990
rect 3425 2955 3575 2990
rect 3675 2955 3825 2990
rect 3925 2955 4000 2990
rect 0 2950 4000 2955
rect 0 2940 60 2950
rect 190 2940 310 2950
rect 440 2940 560 2950
rect 690 2940 810 2950
rect 940 2940 1060 2950
rect 1190 2940 1310 2950
rect 1440 2940 1560 2950
rect 1690 2940 1810 2950
rect 1940 2940 2060 2950
rect 2190 2940 2310 2950
rect 2440 2940 2560 2950
rect 2690 2940 2810 2950
rect 2940 2940 3060 2950
rect 3190 2940 3310 2950
rect 3440 2940 3560 2950
rect 3690 2940 3810 2950
rect 3940 2940 4000 2950
rect 0 2925 50 2940
rect 0 2825 10 2925
rect 45 2825 50 2925
rect 0 2810 50 2825
rect 200 2925 300 2940
rect 200 2825 205 2925
rect 240 2825 260 2925
rect 295 2825 300 2925
rect 200 2810 300 2825
rect 450 2925 550 2940
rect 450 2825 455 2925
rect 490 2825 510 2925
rect 545 2825 550 2925
rect 450 2810 550 2825
rect 700 2925 800 2940
rect 700 2825 705 2925
rect 740 2825 760 2925
rect 795 2825 800 2925
rect 700 2810 800 2825
rect 950 2925 1050 2940
rect 950 2825 955 2925
rect 990 2825 1010 2925
rect 1045 2825 1050 2925
rect 950 2810 1050 2825
rect 1200 2925 1300 2940
rect 1200 2825 1205 2925
rect 1240 2825 1260 2925
rect 1295 2825 1300 2925
rect 1200 2810 1300 2825
rect 1450 2925 1550 2940
rect 1450 2825 1455 2925
rect 1490 2825 1510 2925
rect 1545 2825 1550 2925
rect 1450 2810 1550 2825
rect 1700 2925 1800 2940
rect 1700 2825 1705 2925
rect 1740 2825 1760 2925
rect 1795 2825 1800 2925
rect 1700 2810 1800 2825
rect 1950 2925 2050 2940
rect 1950 2825 1955 2925
rect 1990 2825 2010 2925
rect 2045 2825 2050 2925
rect 1950 2810 2050 2825
rect 2200 2925 2300 2940
rect 2200 2825 2205 2925
rect 2240 2825 2260 2925
rect 2295 2825 2300 2925
rect 2200 2810 2300 2825
rect 2450 2925 2550 2940
rect 2450 2825 2455 2925
rect 2490 2825 2510 2925
rect 2545 2825 2550 2925
rect 2450 2810 2550 2825
rect 2700 2925 2800 2940
rect 2700 2825 2705 2925
rect 2740 2825 2760 2925
rect 2795 2825 2800 2925
rect 2700 2810 2800 2825
rect 2950 2925 3050 2940
rect 2950 2825 2955 2925
rect 2990 2825 3010 2925
rect 3045 2825 3050 2925
rect 2950 2810 3050 2825
rect 3200 2925 3300 2940
rect 3200 2825 3205 2925
rect 3240 2825 3260 2925
rect 3295 2825 3300 2925
rect 3200 2810 3300 2825
rect 3450 2925 3550 2940
rect 3450 2825 3455 2925
rect 3490 2825 3510 2925
rect 3545 2825 3550 2925
rect 3450 2810 3550 2825
rect 3700 2925 3800 2940
rect 3700 2825 3705 2925
rect 3740 2825 3760 2925
rect 3795 2825 3800 2925
rect 3700 2810 3800 2825
rect 3950 2925 4000 2940
rect 3950 2825 3955 2925
rect 3990 2825 4000 2925
rect 3950 2810 4000 2825
rect 0 2800 60 2810
rect 190 2800 310 2810
rect 440 2800 560 2810
rect 690 2800 810 2810
rect 940 2800 1060 2810
rect 1190 2800 1310 2810
rect 1440 2800 1560 2810
rect 1690 2800 1810 2810
rect 1940 2800 2060 2810
rect 2190 2800 2310 2810
rect 2440 2800 2560 2810
rect 2690 2800 2810 2810
rect 2940 2800 3060 2810
rect 3190 2800 3310 2810
rect 3440 2800 3560 2810
rect 3690 2800 3810 2810
rect 3940 2800 4000 2810
rect 0 2795 4000 2800
rect 0 2760 75 2795
rect 175 2760 325 2795
rect 425 2760 575 2795
rect 675 2760 825 2795
rect 925 2760 1075 2795
rect 1175 2760 1325 2795
rect 1425 2760 1575 2795
rect 1675 2760 1825 2795
rect 1925 2760 2075 2795
rect 2175 2760 2325 2795
rect 2425 2760 2575 2795
rect 2675 2760 2825 2795
rect 2925 2760 3075 2795
rect 3175 2760 3325 2795
rect 3425 2760 3575 2795
rect 3675 2760 3825 2795
rect 3925 2760 4000 2795
rect 0 2740 4000 2760
rect 0 2705 75 2740
rect 175 2705 325 2740
rect 425 2705 575 2740
rect 675 2705 825 2740
rect 925 2705 1075 2740
rect 1175 2705 1325 2740
rect 1425 2705 1575 2740
rect 1675 2705 1825 2740
rect 1925 2705 2075 2740
rect 2175 2705 2325 2740
rect 2425 2705 2575 2740
rect 2675 2705 2825 2740
rect 2925 2705 3075 2740
rect 3175 2705 3325 2740
rect 3425 2705 3575 2740
rect 3675 2705 3825 2740
rect 3925 2705 4000 2740
rect 0 2700 4000 2705
rect 0 2690 60 2700
rect 190 2690 310 2700
rect 440 2690 560 2700
rect 690 2690 810 2700
rect 940 2690 1060 2700
rect 1190 2690 1310 2700
rect 1440 2690 1560 2700
rect 1690 2690 1810 2700
rect 1940 2690 2060 2700
rect 2190 2690 2310 2700
rect 2440 2690 2560 2700
rect 2690 2690 2810 2700
rect 2940 2690 3060 2700
rect 3190 2690 3310 2700
rect 3440 2690 3560 2700
rect 3690 2690 3810 2700
rect 3940 2690 4000 2700
rect 0 2675 50 2690
rect 0 2575 10 2675
rect 45 2575 50 2675
rect 0 2560 50 2575
rect 200 2675 300 2690
rect 200 2575 205 2675
rect 240 2575 260 2675
rect 295 2575 300 2675
rect 200 2560 300 2575
rect 450 2675 550 2690
rect 450 2575 455 2675
rect 490 2575 510 2675
rect 545 2575 550 2675
rect 450 2560 550 2575
rect 700 2675 800 2690
rect 700 2575 705 2675
rect 740 2575 760 2675
rect 795 2575 800 2675
rect 700 2560 800 2575
rect 950 2675 1050 2690
rect 950 2575 955 2675
rect 990 2575 1010 2675
rect 1045 2575 1050 2675
rect 950 2560 1050 2575
rect 1200 2675 1300 2690
rect 1200 2575 1205 2675
rect 1240 2575 1260 2675
rect 1295 2575 1300 2675
rect 1200 2560 1300 2575
rect 1450 2675 1550 2690
rect 1450 2575 1455 2675
rect 1490 2575 1510 2675
rect 1545 2575 1550 2675
rect 1450 2560 1550 2575
rect 1700 2675 1800 2690
rect 1700 2575 1705 2675
rect 1740 2575 1760 2675
rect 1795 2575 1800 2675
rect 1700 2560 1800 2575
rect 1950 2675 2050 2690
rect 1950 2575 1955 2675
rect 1990 2575 2010 2675
rect 2045 2575 2050 2675
rect 1950 2560 2050 2575
rect 2200 2675 2300 2690
rect 2200 2575 2205 2675
rect 2240 2575 2260 2675
rect 2295 2575 2300 2675
rect 2200 2560 2300 2575
rect 2450 2675 2550 2690
rect 2450 2575 2455 2675
rect 2490 2575 2510 2675
rect 2545 2575 2550 2675
rect 2450 2560 2550 2575
rect 2700 2675 2800 2690
rect 2700 2575 2705 2675
rect 2740 2575 2760 2675
rect 2795 2575 2800 2675
rect 2700 2560 2800 2575
rect 2950 2675 3050 2690
rect 2950 2575 2955 2675
rect 2990 2575 3010 2675
rect 3045 2575 3050 2675
rect 2950 2560 3050 2575
rect 3200 2675 3300 2690
rect 3200 2575 3205 2675
rect 3240 2575 3260 2675
rect 3295 2575 3300 2675
rect 3200 2560 3300 2575
rect 3450 2675 3550 2690
rect 3450 2575 3455 2675
rect 3490 2575 3510 2675
rect 3545 2575 3550 2675
rect 3450 2560 3550 2575
rect 3700 2675 3800 2690
rect 3700 2575 3705 2675
rect 3740 2575 3760 2675
rect 3795 2575 3800 2675
rect 3700 2560 3800 2575
rect 3950 2675 4000 2690
rect 3950 2575 3955 2675
rect 3990 2575 4000 2675
rect 3950 2560 4000 2575
rect 0 2550 60 2560
rect 190 2550 310 2560
rect 440 2550 560 2560
rect 690 2550 810 2560
rect 940 2550 1060 2560
rect 1190 2550 1310 2560
rect 1440 2550 1560 2560
rect 1690 2550 1810 2560
rect 1940 2550 2060 2560
rect 2190 2550 2310 2560
rect 2440 2550 2560 2560
rect 2690 2550 2810 2560
rect 2940 2550 3060 2560
rect 3190 2550 3310 2560
rect 3440 2550 3560 2560
rect 3690 2550 3810 2560
rect 3940 2550 4000 2560
rect 0 2545 4000 2550
rect 0 2510 75 2545
rect 175 2510 325 2545
rect 425 2510 575 2545
rect 675 2510 825 2545
rect 925 2510 1075 2545
rect 1175 2510 1325 2545
rect 1425 2510 1575 2545
rect 1675 2510 1825 2545
rect 1925 2510 2075 2545
rect 2175 2510 2325 2545
rect 2425 2510 2575 2545
rect 2675 2510 2825 2545
rect 2925 2510 3075 2545
rect 3175 2510 3325 2545
rect 3425 2510 3575 2545
rect 3675 2510 3825 2545
rect 3925 2510 4000 2545
rect 0 2490 4000 2510
rect 0 2455 75 2490
rect 175 2455 325 2490
rect 425 2455 575 2490
rect 675 2455 825 2490
rect 925 2455 1075 2490
rect 1175 2455 1325 2490
rect 1425 2455 1575 2490
rect 1675 2455 1825 2490
rect 1925 2455 2075 2490
rect 2175 2455 2325 2490
rect 2425 2455 2575 2490
rect 2675 2455 2825 2490
rect 2925 2455 3075 2490
rect 3175 2455 3325 2490
rect 3425 2455 3575 2490
rect 3675 2455 3825 2490
rect 3925 2455 4000 2490
rect 0 2450 4000 2455
rect 0 2440 60 2450
rect 190 2440 310 2450
rect 440 2440 560 2450
rect 690 2440 810 2450
rect 940 2440 1060 2450
rect 1190 2440 1310 2450
rect 1440 2440 1560 2450
rect 1690 2440 1810 2450
rect 1940 2440 2060 2450
rect 2190 2440 2310 2450
rect 2440 2440 2560 2450
rect 2690 2440 2810 2450
rect 2940 2440 3060 2450
rect 3190 2440 3310 2450
rect 3440 2440 3560 2450
rect 3690 2440 3810 2450
rect 3940 2440 4000 2450
rect 0 2425 50 2440
rect 0 2325 10 2425
rect 45 2325 50 2425
rect 0 2310 50 2325
rect 200 2425 300 2440
rect 200 2325 205 2425
rect 240 2325 260 2425
rect 295 2325 300 2425
rect 200 2310 300 2325
rect 450 2425 550 2440
rect 450 2325 455 2425
rect 490 2325 510 2425
rect 545 2325 550 2425
rect 450 2310 550 2325
rect 700 2425 800 2440
rect 700 2325 705 2425
rect 740 2325 760 2425
rect 795 2325 800 2425
rect 700 2310 800 2325
rect 950 2425 1050 2440
rect 950 2325 955 2425
rect 990 2325 1010 2425
rect 1045 2325 1050 2425
rect 950 2310 1050 2325
rect 1200 2425 1300 2440
rect 1200 2325 1205 2425
rect 1240 2325 1260 2425
rect 1295 2325 1300 2425
rect 1200 2310 1300 2325
rect 1450 2425 1550 2440
rect 1450 2325 1455 2425
rect 1490 2325 1510 2425
rect 1545 2325 1550 2425
rect 1450 2310 1550 2325
rect 1700 2425 1800 2440
rect 1700 2325 1705 2425
rect 1740 2325 1760 2425
rect 1795 2325 1800 2425
rect 1700 2310 1800 2325
rect 1950 2425 2050 2440
rect 1950 2325 1955 2425
rect 1990 2325 2010 2425
rect 2045 2325 2050 2425
rect 1950 2310 2050 2325
rect 2200 2425 2300 2440
rect 2200 2325 2205 2425
rect 2240 2325 2260 2425
rect 2295 2325 2300 2425
rect 2200 2310 2300 2325
rect 2450 2425 2550 2440
rect 2450 2325 2455 2425
rect 2490 2325 2510 2425
rect 2545 2325 2550 2425
rect 2450 2310 2550 2325
rect 2700 2425 2800 2440
rect 2700 2325 2705 2425
rect 2740 2325 2760 2425
rect 2795 2325 2800 2425
rect 2700 2310 2800 2325
rect 2950 2425 3050 2440
rect 2950 2325 2955 2425
rect 2990 2325 3010 2425
rect 3045 2325 3050 2425
rect 2950 2310 3050 2325
rect 3200 2425 3300 2440
rect 3200 2325 3205 2425
rect 3240 2325 3260 2425
rect 3295 2325 3300 2425
rect 3200 2310 3300 2325
rect 3450 2425 3550 2440
rect 3450 2325 3455 2425
rect 3490 2325 3510 2425
rect 3545 2325 3550 2425
rect 3450 2310 3550 2325
rect 3700 2425 3800 2440
rect 3700 2325 3705 2425
rect 3740 2325 3760 2425
rect 3795 2325 3800 2425
rect 3700 2310 3800 2325
rect 3950 2425 4000 2440
rect 3950 2325 3955 2425
rect 3990 2325 4000 2425
rect 3950 2310 4000 2325
rect 0 2300 60 2310
rect 190 2300 310 2310
rect 440 2300 560 2310
rect 690 2300 810 2310
rect 940 2300 1060 2310
rect 1190 2300 1310 2310
rect 1440 2300 1560 2310
rect 1690 2300 1810 2310
rect 1940 2300 2060 2310
rect 2190 2300 2310 2310
rect 2440 2300 2560 2310
rect 2690 2300 2810 2310
rect 2940 2300 3060 2310
rect 3190 2300 3310 2310
rect 3440 2300 3560 2310
rect 3690 2300 3810 2310
rect 3940 2300 4000 2310
rect 0 2295 4000 2300
rect 0 2260 75 2295
rect 175 2260 325 2295
rect 425 2260 575 2295
rect 675 2260 825 2295
rect 925 2260 1075 2295
rect 1175 2260 1325 2295
rect 1425 2260 1575 2295
rect 1675 2260 1825 2295
rect 1925 2260 2075 2295
rect 2175 2260 2325 2295
rect 2425 2260 2575 2295
rect 2675 2260 2825 2295
rect 2925 2260 3075 2295
rect 3175 2260 3325 2295
rect 3425 2260 3575 2295
rect 3675 2260 3825 2295
rect 3925 2260 4000 2295
rect 0 2240 4000 2260
rect 0 2205 75 2240
rect 175 2205 325 2240
rect 425 2205 575 2240
rect 675 2205 825 2240
rect 925 2205 1075 2240
rect 1175 2205 1325 2240
rect 1425 2205 1575 2240
rect 1675 2205 1825 2240
rect 1925 2205 2075 2240
rect 2175 2205 2325 2240
rect 2425 2205 2575 2240
rect 2675 2205 2825 2240
rect 2925 2205 3075 2240
rect 3175 2205 3325 2240
rect 3425 2205 3575 2240
rect 3675 2205 3825 2240
rect 3925 2205 4000 2240
rect 0 2200 4000 2205
rect 0 2190 60 2200
rect 190 2190 310 2200
rect 440 2190 560 2200
rect 690 2190 810 2200
rect 940 2190 1060 2200
rect 1190 2190 1310 2200
rect 1440 2190 1560 2200
rect 1690 2190 1810 2200
rect 1940 2190 2060 2200
rect 2190 2190 2310 2200
rect 2440 2190 2560 2200
rect 2690 2190 2810 2200
rect 2940 2190 3060 2200
rect 3190 2190 3310 2200
rect 3440 2190 3560 2200
rect 3690 2190 3810 2200
rect 3940 2190 4000 2200
rect 0 2175 50 2190
rect 0 2075 10 2175
rect 45 2075 50 2175
rect 0 2060 50 2075
rect 200 2175 300 2190
rect 200 2075 205 2175
rect 240 2075 260 2175
rect 295 2075 300 2175
rect 200 2060 300 2075
rect 450 2175 550 2190
rect 450 2075 455 2175
rect 490 2075 510 2175
rect 545 2075 550 2175
rect 450 2060 550 2075
rect 700 2175 800 2190
rect 700 2075 705 2175
rect 740 2075 760 2175
rect 795 2075 800 2175
rect 700 2060 800 2075
rect 950 2175 1050 2190
rect 950 2075 955 2175
rect 990 2075 1010 2175
rect 1045 2075 1050 2175
rect 950 2060 1050 2075
rect 1200 2175 1300 2190
rect 1200 2075 1205 2175
rect 1240 2075 1260 2175
rect 1295 2075 1300 2175
rect 1200 2060 1300 2075
rect 1450 2175 1550 2190
rect 1450 2075 1455 2175
rect 1490 2075 1510 2175
rect 1545 2075 1550 2175
rect 1450 2060 1550 2075
rect 1700 2175 1800 2190
rect 1700 2075 1705 2175
rect 1740 2075 1760 2175
rect 1795 2075 1800 2175
rect 1700 2060 1800 2075
rect 1950 2175 2050 2190
rect 1950 2075 1955 2175
rect 1990 2075 2010 2175
rect 2045 2075 2050 2175
rect 1950 2060 2050 2075
rect 2200 2175 2300 2190
rect 2200 2075 2205 2175
rect 2240 2075 2260 2175
rect 2295 2075 2300 2175
rect 2200 2060 2300 2075
rect 2450 2175 2550 2190
rect 2450 2075 2455 2175
rect 2490 2075 2510 2175
rect 2545 2075 2550 2175
rect 2450 2060 2550 2075
rect 2700 2175 2800 2190
rect 2700 2075 2705 2175
rect 2740 2075 2760 2175
rect 2795 2075 2800 2175
rect 2700 2060 2800 2075
rect 2950 2175 3050 2190
rect 2950 2075 2955 2175
rect 2990 2075 3010 2175
rect 3045 2075 3050 2175
rect 2950 2060 3050 2075
rect 3200 2175 3300 2190
rect 3200 2075 3205 2175
rect 3240 2075 3260 2175
rect 3295 2075 3300 2175
rect 3200 2060 3300 2075
rect 3450 2175 3550 2190
rect 3450 2075 3455 2175
rect 3490 2075 3510 2175
rect 3545 2075 3550 2175
rect 3450 2060 3550 2075
rect 3700 2175 3800 2190
rect 3700 2075 3705 2175
rect 3740 2075 3760 2175
rect 3795 2075 3800 2175
rect 3700 2060 3800 2075
rect 3950 2175 4000 2190
rect 3950 2075 3955 2175
rect 3990 2075 4000 2175
rect 3950 2060 4000 2075
rect 0 2050 60 2060
rect 190 2050 310 2060
rect 440 2050 560 2060
rect 690 2050 810 2060
rect 940 2050 1060 2060
rect 1190 2050 1310 2060
rect 1440 2050 1560 2060
rect 1690 2050 1810 2060
rect 1940 2050 2060 2060
rect 2190 2050 2310 2060
rect 2440 2050 2560 2060
rect 2690 2050 2810 2060
rect 2940 2050 3060 2060
rect 3190 2050 3310 2060
rect 3440 2050 3560 2060
rect 3690 2050 3810 2060
rect 3940 2050 4000 2060
rect 0 2045 4000 2050
rect 0 2010 75 2045
rect 175 2010 325 2045
rect 425 2010 575 2045
rect 675 2010 825 2045
rect 925 2010 1075 2045
rect 1175 2010 1325 2045
rect 1425 2010 1575 2045
rect 1675 2010 1825 2045
rect 1925 2010 2075 2045
rect 2175 2010 2325 2045
rect 2425 2010 2575 2045
rect 2675 2010 2825 2045
rect 2925 2010 3075 2045
rect 3175 2010 3325 2045
rect 3425 2010 3575 2045
rect 3675 2010 3825 2045
rect 3925 2010 4000 2045
rect 0 1990 4000 2010
rect 0 1955 75 1990
rect 175 1955 325 1990
rect 425 1955 575 1990
rect 675 1955 825 1990
rect 925 1955 1075 1990
rect 1175 1955 1325 1990
rect 1425 1955 1575 1990
rect 1675 1955 1825 1990
rect 1925 1955 2075 1990
rect 2175 1955 2325 1990
rect 2425 1955 2575 1990
rect 2675 1955 2825 1990
rect 2925 1955 3075 1990
rect 3175 1955 3325 1990
rect 3425 1955 3575 1990
rect 3675 1955 3825 1990
rect 3925 1955 4000 1990
rect 0 1950 4000 1955
rect 0 1940 60 1950
rect 190 1940 310 1950
rect 440 1940 560 1950
rect 690 1940 810 1950
rect 940 1940 1060 1950
rect 1190 1940 1310 1950
rect 1440 1940 1560 1950
rect 1690 1940 1810 1950
rect 1940 1940 2060 1950
rect 2190 1940 2310 1950
rect 2440 1940 2560 1950
rect 2690 1940 2810 1950
rect 2940 1940 3060 1950
rect 3190 1940 3310 1950
rect 3440 1940 3560 1950
rect 3690 1940 3810 1950
rect 3940 1940 4000 1950
rect 0 1925 50 1940
rect 0 1825 10 1925
rect 45 1825 50 1925
rect 0 1810 50 1825
rect 200 1925 300 1940
rect 200 1825 205 1925
rect 240 1825 260 1925
rect 295 1825 300 1925
rect 200 1810 300 1825
rect 450 1925 550 1940
rect 450 1825 455 1925
rect 490 1825 510 1925
rect 545 1825 550 1925
rect 450 1810 550 1825
rect 700 1925 800 1940
rect 700 1825 705 1925
rect 740 1825 760 1925
rect 795 1825 800 1925
rect 700 1810 800 1825
rect 950 1925 1050 1940
rect 950 1825 955 1925
rect 990 1825 1010 1925
rect 1045 1825 1050 1925
rect 950 1810 1050 1825
rect 1200 1925 1300 1940
rect 1200 1825 1205 1925
rect 1240 1825 1260 1925
rect 1295 1825 1300 1925
rect 1200 1810 1300 1825
rect 1450 1925 1550 1940
rect 1450 1825 1455 1925
rect 1490 1825 1510 1925
rect 1545 1825 1550 1925
rect 1450 1810 1550 1825
rect 1700 1925 1800 1940
rect 1700 1825 1705 1925
rect 1740 1825 1760 1925
rect 1795 1825 1800 1925
rect 1700 1810 1800 1825
rect 1950 1925 2050 1940
rect 1950 1825 1955 1925
rect 1990 1825 2010 1925
rect 2045 1825 2050 1925
rect 1950 1810 2050 1825
rect 2200 1925 2300 1940
rect 2200 1825 2205 1925
rect 2240 1825 2260 1925
rect 2295 1825 2300 1925
rect 2200 1810 2300 1825
rect 2450 1925 2550 1940
rect 2450 1825 2455 1925
rect 2490 1825 2510 1925
rect 2545 1825 2550 1925
rect 2450 1810 2550 1825
rect 2700 1925 2800 1940
rect 2700 1825 2705 1925
rect 2740 1825 2760 1925
rect 2795 1825 2800 1925
rect 2700 1810 2800 1825
rect 2950 1925 3050 1940
rect 2950 1825 2955 1925
rect 2990 1825 3010 1925
rect 3045 1825 3050 1925
rect 2950 1810 3050 1825
rect 3200 1925 3300 1940
rect 3200 1825 3205 1925
rect 3240 1825 3260 1925
rect 3295 1825 3300 1925
rect 3200 1810 3300 1825
rect 3450 1925 3550 1940
rect 3450 1825 3455 1925
rect 3490 1825 3510 1925
rect 3545 1825 3550 1925
rect 3450 1810 3550 1825
rect 3700 1925 3800 1940
rect 3700 1825 3705 1925
rect 3740 1825 3760 1925
rect 3795 1825 3800 1925
rect 3700 1810 3800 1825
rect 3950 1925 4000 1940
rect 3950 1825 3955 1925
rect 3990 1825 4000 1925
rect 3950 1810 4000 1825
rect 0 1800 60 1810
rect 190 1800 310 1810
rect 440 1800 560 1810
rect 690 1800 810 1810
rect 940 1800 1060 1810
rect 1190 1800 1310 1810
rect 1440 1800 1560 1810
rect 1690 1800 1810 1810
rect 1940 1800 2060 1810
rect 2190 1800 2310 1810
rect 2440 1800 2560 1810
rect 2690 1800 2810 1810
rect 2940 1800 3060 1810
rect 3190 1800 3310 1810
rect 3440 1800 3560 1810
rect 3690 1800 3810 1810
rect 3940 1800 4000 1810
rect 0 1795 4000 1800
rect 0 1760 75 1795
rect 175 1760 325 1795
rect 425 1760 575 1795
rect 675 1760 825 1795
rect 925 1760 1075 1795
rect 1175 1760 1325 1795
rect 1425 1760 1575 1795
rect 1675 1760 1825 1795
rect 1925 1760 2075 1795
rect 2175 1760 2325 1795
rect 2425 1760 2575 1795
rect 2675 1760 2825 1795
rect 2925 1760 3075 1795
rect 3175 1760 3325 1795
rect 3425 1760 3575 1795
rect 3675 1760 3825 1795
rect 3925 1760 4000 1795
rect 0 1740 4000 1760
rect 0 1705 75 1740
rect 175 1705 325 1740
rect 425 1705 575 1740
rect 675 1705 825 1740
rect 925 1705 1075 1740
rect 1175 1705 1325 1740
rect 1425 1705 1575 1740
rect 1675 1705 1825 1740
rect 1925 1705 2075 1740
rect 2175 1705 2325 1740
rect 2425 1705 2575 1740
rect 2675 1705 2825 1740
rect 2925 1705 3075 1740
rect 3175 1705 3325 1740
rect 3425 1705 3575 1740
rect 3675 1705 3825 1740
rect 3925 1705 4000 1740
rect 0 1700 4000 1705
rect 0 1690 60 1700
rect 190 1690 310 1700
rect 440 1690 560 1700
rect 690 1690 810 1700
rect 940 1690 1060 1700
rect 1190 1690 1310 1700
rect 1440 1690 1560 1700
rect 1690 1690 1810 1700
rect 1940 1690 2060 1700
rect 2190 1690 2310 1700
rect 2440 1690 2560 1700
rect 2690 1690 2810 1700
rect 2940 1690 3060 1700
rect 3190 1690 3310 1700
rect 3440 1690 3560 1700
rect 3690 1690 3810 1700
rect 3940 1690 4000 1700
rect 0 1675 50 1690
rect 0 1575 10 1675
rect 45 1575 50 1675
rect 0 1560 50 1575
rect 200 1675 300 1690
rect 200 1575 205 1675
rect 240 1575 260 1675
rect 295 1575 300 1675
rect 200 1560 300 1575
rect 450 1675 550 1690
rect 450 1575 455 1675
rect 490 1575 510 1675
rect 545 1575 550 1675
rect 450 1560 550 1575
rect 700 1675 800 1690
rect 700 1575 705 1675
rect 740 1575 760 1675
rect 795 1575 800 1675
rect 700 1560 800 1575
rect 950 1675 1050 1690
rect 950 1575 955 1675
rect 990 1575 1010 1675
rect 1045 1575 1050 1675
rect 950 1560 1050 1575
rect 1200 1675 1300 1690
rect 1200 1575 1205 1675
rect 1240 1575 1260 1675
rect 1295 1575 1300 1675
rect 1200 1560 1300 1575
rect 1450 1675 1550 1690
rect 1450 1575 1455 1675
rect 1490 1575 1510 1675
rect 1545 1575 1550 1675
rect 1450 1560 1550 1575
rect 1700 1675 1800 1690
rect 1700 1575 1705 1675
rect 1740 1575 1760 1675
rect 1795 1575 1800 1675
rect 1700 1560 1800 1575
rect 1950 1675 2050 1690
rect 1950 1575 1955 1675
rect 1990 1575 2010 1675
rect 2045 1575 2050 1675
rect 1950 1560 2050 1575
rect 2200 1675 2300 1690
rect 2200 1575 2205 1675
rect 2240 1575 2260 1675
rect 2295 1575 2300 1675
rect 2200 1560 2300 1575
rect 2450 1675 2550 1690
rect 2450 1575 2455 1675
rect 2490 1575 2510 1675
rect 2545 1575 2550 1675
rect 2450 1560 2550 1575
rect 2700 1675 2800 1690
rect 2700 1575 2705 1675
rect 2740 1575 2760 1675
rect 2795 1575 2800 1675
rect 2700 1560 2800 1575
rect 2950 1675 3050 1690
rect 2950 1575 2955 1675
rect 2990 1575 3010 1675
rect 3045 1575 3050 1675
rect 2950 1560 3050 1575
rect 3200 1675 3300 1690
rect 3200 1575 3205 1675
rect 3240 1575 3260 1675
rect 3295 1575 3300 1675
rect 3200 1560 3300 1575
rect 3450 1675 3550 1690
rect 3450 1575 3455 1675
rect 3490 1575 3510 1675
rect 3545 1575 3550 1675
rect 3450 1560 3550 1575
rect 3700 1675 3800 1690
rect 3700 1575 3705 1675
rect 3740 1575 3760 1675
rect 3795 1575 3800 1675
rect 3700 1560 3800 1575
rect 3950 1675 4000 1690
rect 3950 1575 3955 1675
rect 3990 1575 4000 1675
rect 3950 1560 4000 1575
rect 0 1550 60 1560
rect 190 1550 310 1560
rect 440 1550 560 1560
rect 690 1550 810 1560
rect 940 1550 1060 1560
rect 1190 1550 1310 1560
rect 1440 1550 1560 1560
rect 1690 1550 1810 1560
rect 1940 1550 2060 1560
rect 2190 1550 2310 1560
rect 2440 1550 2560 1560
rect 2690 1550 2810 1560
rect 2940 1550 3060 1560
rect 3190 1550 3310 1560
rect 3440 1550 3560 1560
rect 3690 1550 3810 1560
rect 3940 1550 4000 1560
rect 0 1545 4000 1550
rect 0 1510 75 1545
rect 175 1510 325 1545
rect 425 1510 575 1545
rect 675 1510 825 1545
rect 925 1510 1075 1545
rect 1175 1510 1325 1545
rect 1425 1510 1575 1545
rect 1675 1510 1825 1545
rect 1925 1510 2075 1545
rect 2175 1510 2325 1545
rect 2425 1510 2575 1545
rect 2675 1510 2825 1545
rect 2925 1510 3075 1545
rect 3175 1510 3325 1545
rect 3425 1510 3575 1545
rect 3675 1510 3825 1545
rect 3925 1510 4000 1545
rect 0 1490 4000 1510
rect 0 1455 75 1490
rect 175 1455 325 1490
rect 425 1455 575 1490
rect 675 1455 825 1490
rect 925 1455 1075 1490
rect 1175 1455 1325 1490
rect 1425 1455 1575 1490
rect 1675 1455 1825 1490
rect 1925 1455 2075 1490
rect 2175 1455 2325 1490
rect 2425 1455 2575 1490
rect 2675 1455 2825 1490
rect 2925 1455 3075 1490
rect 3175 1455 3325 1490
rect 3425 1455 3575 1490
rect 3675 1455 3825 1490
rect 3925 1455 4000 1490
rect 0 1450 4000 1455
rect 0 1440 60 1450
rect 190 1440 310 1450
rect 440 1440 560 1450
rect 690 1440 810 1450
rect 940 1440 1060 1450
rect 1190 1440 1310 1450
rect 1440 1440 1560 1450
rect 1690 1440 1810 1450
rect 1940 1440 2060 1450
rect 2190 1440 2310 1450
rect 2440 1440 2560 1450
rect 2690 1440 2810 1450
rect 2940 1440 3060 1450
rect 3190 1440 3310 1450
rect 3440 1440 3560 1450
rect 3690 1440 3810 1450
rect 3940 1440 4000 1450
rect 0 1425 50 1440
rect 0 1325 10 1425
rect 45 1325 50 1425
rect 0 1310 50 1325
rect 200 1425 300 1440
rect 200 1325 205 1425
rect 240 1325 260 1425
rect 295 1325 300 1425
rect 200 1310 300 1325
rect 450 1425 550 1440
rect 450 1325 455 1425
rect 490 1325 510 1425
rect 545 1325 550 1425
rect 450 1310 550 1325
rect 700 1425 800 1440
rect 700 1325 705 1425
rect 740 1325 760 1425
rect 795 1325 800 1425
rect 700 1310 800 1325
rect 950 1425 1050 1440
rect 950 1325 955 1425
rect 990 1325 1010 1425
rect 1045 1325 1050 1425
rect 950 1310 1050 1325
rect 1200 1425 1300 1440
rect 1200 1325 1205 1425
rect 1240 1325 1260 1425
rect 1295 1325 1300 1425
rect 1200 1310 1300 1325
rect 1450 1425 1550 1440
rect 1450 1325 1455 1425
rect 1490 1325 1510 1425
rect 1545 1325 1550 1425
rect 1450 1310 1550 1325
rect 1700 1425 1800 1440
rect 1700 1325 1705 1425
rect 1740 1325 1760 1425
rect 1795 1325 1800 1425
rect 1700 1310 1800 1325
rect 1950 1425 2050 1440
rect 1950 1325 1955 1425
rect 1990 1325 2010 1425
rect 2045 1325 2050 1425
rect 1950 1310 2050 1325
rect 2200 1425 2300 1440
rect 2200 1325 2205 1425
rect 2240 1325 2260 1425
rect 2295 1325 2300 1425
rect 2200 1310 2300 1325
rect 2450 1425 2550 1440
rect 2450 1325 2455 1425
rect 2490 1325 2510 1425
rect 2545 1325 2550 1425
rect 2450 1310 2550 1325
rect 2700 1425 2800 1440
rect 2700 1325 2705 1425
rect 2740 1325 2760 1425
rect 2795 1325 2800 1425
rect 2700 1310 2800 1325
rect 2950 1425 3050 1440
rect 2950 1325 2955 1425
rect 2990 1325 3010 1425
rect 3045 1325 3050 1425
rect 2950 1310 3050 1325
rect 3200 1425 3300 1440
rect 3200 1325 3205 1425
rect 3240 1325 3260 1425
rect 3295 1325 3300 1425
rect 3200 1310 3300 1325
rect 3450 1425 3550 1440
rect 3450 1325 3455 1425
rect 3490 1325 3510 1425
rect 3545 1325 3550 1425
rect 3450 1310 3550 1325
rect 3700 1425 3800 1440
rect 3700 1325 3705 1425
rect 3740 1325 3760 1425
rect 3795 1325 3800 1425
rect 3700 1310 3800 1325
rect 3950 1425 4000 1440
rect 3950 1325 3955 1425
rect 3990 1325 4000 1425
rect 3950 1310 4000 1325
rect 0 1300 60 1310
rect 190 1300 310 1310
rect 440 1300 560 1310
rect 690 1300 810 1310
rect 940 1300 1060 1310
rect 1190 1300 1310 1310
rect 1440 1300 1560 1310
rect 1690 1300 1810 1310
rect 1940 1300 2060 1310
rect 2190 1300 2310 1310
rect 2440 1300 2560 1310
rect 2690 1300 2810 1310
rect 2940 1300 3060 1310
rect 3190 1300 3310 1310
rect 3440 1300 3560 1310
rect 3690 1300 3810 1310
rect 3940 1300 4000 1310
rect 0 1295 4000 1300
rect 0 1260 75 1295
rect 175 1260 325 1295
rect 425 1260 575 1295
rect 675 1260 825 1295
rect 925 1260 1075 1295
rect 1175 1260 1325 1295
rect 1425 1260 1575 1295
rect 1675 1260 1825 1295
rect 1925 1260 2075 1295
rect 2175 1260 2325 1295
rect 2425 1260 2575 1295
rect 2675 1260 2825 1295
rect 2925 1260 3075 1295
rect 3175 1260 3325 1295
rect 3425 1260 3575 1295
rect 3675 1260 3825 1295
rect 3925 1260 4000 1295
rect 0 1240 4000 1260
rect 0 1205 75 1240
rect 175 1205 325 1240
rect 425 1205 575 1240
rect 675 1205 825 1240
rect 925 1205 1075 1240
rect 1175 1205 1325 1240
rect 1425 1205 1575 1240
rect 1675 1205 1825 1240
rect 1925 1205 2075 1240
rect 2175 1205 2325 1240
rect 2425 1205 2575 1240
rect 2675 1205 2825 1240
rect 2925 1205 3075 1240
rect 3175 1205 3325 1240
rect 3425 1205 3575 1240
rect 3675 1205 3825 1240
rect 3925 1205 4000 1240
rect 0 1200 4000 1205
rect 0 1190 60 1200
rect 190 1190 310 1200
rect 440 1190 560 1200
rect 690 1190 810 1200
rect 940 1190 1060 1200
rect 1190 1190 1310 1200
rect 1440 1190 1560 1200
rect 1690 1190 1810 1200
rect 1940 1190 2060 1200
rect 2190 1190 2310 1200
rect 2440 1190 2560 1200
rect 2690 1190 2810 1200
rect 2940 1190 3060 1200
rect 3190 1190 3310 1200
rect 3440 1190 3560 1200
rect 3690 1190 3810 1200
rect 3940 1190 4000 1200
rect 0 1175 50 1190
rect 0 1075 10 1175
rect 45 1075 50 1175
rect 0 1060 50 1075
rect 200 1175 300 1190
rect 200 1075 205 1175
rect 240 1075 260 1175
rect 295 1075 300 1175
rect 200 1060 300 1075
rect 450 1175 550 1190
rect 450 1075 455 1175
rect 490 1075 510 1175
rect 545 1075 550 1175
rect 450 1060 550 1075
rect 700 1175 800 1190
rect 700 1075 705 1175
rect 740 1075 760 1175
rect 795 1075 800 1175
rect 700 1060 800 1075
rect 950 1175 1050 1190
rect 950 1075 955 1175
rect 990 1075 1010 1175
rect 1045 1075 1050 1175
rect 950 1060 1050 1075
rect 1200 1175 1300 1190
rect 1200 1075 1205 1175
rect 1240 1075 1260 1175
rect 1295 1075 1300 1175
rect 1200 1060 1300 1075
rect 1450 1175 1550 1190
rect 1450 1075 1455 1175
rect 1490 1075 1510 1175
rect 1545 1075 1550 1175
rect 1450 1060 1550 1075
rect 1700 1175 1800 1190
rect 1700 1075 1705 1175
rect 1740 1075 1760 1175
rect 1795 1075 1800 1175
rect 1700 1060 1800 1075
rect 1950 1175 2050 1190
rect 1950 1075 1955 1175
rect 1990 1075 2010 1175
rect 2045 1075 2050 1175
rect 1950 1060 2050 1075
rect 2200 1175 2300 1190
rect 2200 1075 2205 1175
rect 2240 1075 2260 1175
rect 2295 1075 2300 1175
rect 2200 1060 2300 1075
rect 2450 1175 2550 1190
rect 2450 1075 2455 1175
rect 2490 1075 2510 1175
rect 2545 1075 2550 1175
rect 2450 1060 2550 1075
rect 2700 1175 2800 1190
rect 2700 1075 2705 1175
rect 2740 1075 2760 1175
rect 2795 1075 2800 1175
rect 2700 1060 2800 1075
rect 2950 1175 3050 1190
rect 2950 1075 2955 1175
rect 2990 1075 3010 1175
rect 3045 1075 3050 1175
rect 2950 1060 3050 1075
rect 3200 1175 3300 1190
rect 3200 1075 3205 1175
rect 3240 1075 3260 1175
rect 3295 1075 3300 1175
rect 3200 1060 3300 1075
rect 3450 1175 3550 1190
rect 3450 1075 3455 1175
rect 3490 1075 3510 1175
rect 3545 1075 3550 1175
rect 3450 1060 3550 1075
rect 3700 1175 3800 1190
rect 3700 1075 3705 1175
rect 3740 1075 3760 1175
rect 3795 1075 3800 1175
rect 3700 1060 3800 1075
rect 3950 1175 4000 1190
rect 3950 1075 3955 1175
rect 3990 1075 4000 1175
rect 3950 1060 4000 1075
rect 0 1050 60 1060
rect 190 1050 310 1060
rect 440 1050 560 1060
rect 690 1050 810 1060
rect 940 1050 1060 1060
rect 1190 1050 1310 1060
rect 1440 1050 1560 1060
rect 1690 1050 1810 1060
rect 1940 1050 2060 1060
rect 2190 1050 2310 1060
rect 2440 1050 2560 1060
rect 2690 1050 2810 1060
rect 2940 1050 3060 1060
rect 3190 1050 3310 1060
rect 3440 1050 3560 1060
rect 3690 1050 3810 1060
rect 3940 1050 4000 1060
rect 0 1045 4000 1050
rect 0 1010 75 1045
rect 175 1010 325 1045
rect 425 1010 575 1045
rect 675 1010 825 1045
rect 925 1010 1075 1045
rect 1175 1010 1325 1045
rect 1425 1010 1575 1045
rect 1675 1010 1825 1045
rect 1925 1010 2075 1045
rect 2175 1010 2325 1045
rect 2425 1010 2575 1045
rect 2675 1010 2825 1045
rect 2925 1010 3075 1045
rect 3175 1010 3325 1045
rect 3425 1010 3575 1045
rect 3675 1010 3825 1045
rect 3925 1010 4000 1045
rect 0 990 4000 1010
rect 0 955 75 990
rect 175 955 325 990
rect 425 955 575 990
rect 675 955 825 990
rect 925 955 1075 990
rect 1175 955 1325 990
rect 1425 955 1575 990
rect 1675 955 1825 990
rect 1925 955 2075 990
rect 2175 955 2325 990
rect 2425 955 2575 990
rect 2675 955 2825 990
rect 2925 955 3075 990
rect 3175 955 3325 990
rect 3425 955 3575 990
rect 3675 955 3825 990
rect 3925 955 4000 990
rect 0 950 4000 955
rect 0 940 60 950
rect 190 940 310 950
rect 440 940 560 950
rect 690 940 810 950
rect 940 940 1060 950
rect 1190 940 1310 950
rect 1440 940 1560 950
rect 1690 940 1810 950
rect 1940 940 2060 950
rect 2190 940 2310 950
rect 2440 940 2560 950
rect 2690 940 2810 950
rect 2940 940 3060 950
rect 3190 940 3310 950
rect 3440 940 3560 950
rect 3690 940 3810 950
rect 3940 940 4000 950
rect 0 925 50 940
rect 0 825 10 925
rect 45 825 50 925
rect 0 810 50 825
rect 200 925 300 940
rect 200 825 205 925
rect 240 825 260 925
rect 295 825 300 925
rect 200 810 300 825
rect 450 925 550 940
rect 450 825 455 925
rect 490 825 510 925
rect 545 825 550 925
rect 450 810 550 825
rect 700 925 800 940
rect 700 825 705 925
rect 740 825 760 925
rect 795 825 800 925
rect 700 810 800 825
rect 950 925 1050 940
rect 950 825 955 925
rect 990 825 1010 925
rect 1045 825 1050 925
rect 950 810 1050 825
rect 1200 925 1300 940
rect 1200 825 1205 925
rect 1240 825 1260 925
rect 1295 825 1300 925
rect 1200 810 1300 825
rect 1450 925 1550 940
rect 1450 825 1455 925
rect 1490 825 1510 925
rect 1545 825 1550 925
rect 1450 810 1550 825
rect 1700 925 1800 940
rect 1700 825 1705 925
rect 1740 825 1760 925
rect 1795 825 1800 925
rect 1700 810 1800 825
rect 1950 925 2050 940
rect 1950 825 1955 925
rect 1990 825 2010 925
rect 2045 825 2050 925
rect 1950 810 2050 825
rect 2200 925 2300 940
rect 2200 825 2205 925
rect 2240 825 2260 925
rect 2295 825 2300 925
rect 2200 810 2300 825
rect 2450 925 2550 940
rect 2450 825 2455 925
rect 2490 825 2510 925
rect 2545 825 2550 925
rect 2450 810 2550 825
rect 2700 925 2800 940
rect 2700 825 2705 925
rect 2740 825 2760 925
rect 2795 825 2800 925
rect 2700 810 2800 825
rect 2950 925 3050 940
rect 2950 825 2955 925
rect 2990 825 3010 925
rect 3045 825 3050 925
rect 2950 810 3050 825
rect 3200 925 3300 940
rect 3200 825 3205 925
rect 3240 825 3260 925
rect 3295 825 3300 925
rect 3200 810 3300 825
rect 3450 925 3550 940
rect 3450 825 3455 925
rect 3490 825 3510 925
rect 3545 825 3550 925
rect 3450 810 3550 825
rect 3700 925 3800 940
rect 3700 825 3705 925
rect 3740 825 3760 925
rect 3795 825 3800 925
rect 3700 810 3800 825
rect 3950 925 4000 940
rect 3950 825 3955 925
rect 3990 825 4000 925
rect 3950 810 4000 825
rect 0 800 60 810
rect 190 800 310 810
rect 440 800 560 810
rect 690 800 810 810
rect 940 800 1060 810
rect 1190 800 1310 810
rect 1440 800 1560 810
rect 1690 800 1810 810
rect 1940 800 2060 810
rect 2190 800 2310 810
rect 2440 800 2560 810
rect 2690 800 2810 810
rect 2940 800 3060 810
rect 3190 800 3310 810
rect 3440 800 3560 810
rect 3690 800 3810 810
rect 3940 800 4000 810
rect 0 795 4000 800
rect 0 760 75 795
rect 175 760 325 795
rect 425 760 575 795
rect 675 760 825 795
rect 925 760 1075 795
rect 1175 760 1325 795
rect 1425 760 1575 795
rect 1675 760 1825 795
rect 1925 760 2075 795
rect 2175 760 2325 795
rect 2425 760 2575 795
rect 2675 760 2825 795
rect 2925 760 3075 795
rect 3175 760 3325 795
rect 3425 760 3575 795
rect 3675 760 3825 795
rect 3925 760 4000 795
rect 0 740 4000 760
rect 0 705 75 740
rect 175 705 325 740
rect 425 705 575 740
rect 675 705 825 740
rect 925 705 1075 740
rect 1175 705 1325 740
rect 1425 705 1575 740
rect 1675 705 1825 740
rect 1925 705 2075 740
rect 2175 705 2325 740
rect 2425 705 2575 740
rect 2675 705 2825 740
rect 2925 705 3075 740
rect 3175 705 3325 740
rect 3425 705 3575 740
rect 3675 705 3825 740
rect 3925 705 4000 740
rect 0 700 4000 705
rect 0 690 60 700
rect 190 690 310 700
rect 440 690 560 700
rect 690 690 810 700
rect 940 690 1060 700
rect 1190 690 1310 700
rect 1440 690 1560 700
rect 1690 690 1810 700
rect 1940 690 2060 700
rect 2190 690 2310 700
rect 2440 690 2560 700
rect 2690 690 2810 700
rect 2940 690 3060 700
rect 3190 690 3310 700
rect 3440 690 3560 700
rect 3690 690 3810 700
rect 3940 690 4000 700
rect 0 675 50 690
rect 0 575 10 675
rect 45 575 50 675
rect 0 560 50 575
rect 200 675 300 690
rect 200 575 205 675
rect 240 575 260 675
rect 295 575 300 675
rect 200 560 300 575
rect 450 675 550 690
rect 450 575 455 675
rect 490 575 510 675
rect 545 575 550 675
rect 450 560 550 575
rect 700 675 800 690
rect 700 575 705 675
rect 740 575 760 675
rect 795 575 800 675
rect 700 560 800 575
rect 950 675 1050 690
rect 950 575 955 675
rect 990 575 1010 675
rect 1045 575 1050 675
rect 950 560 1050 575
rect 1200 675 1300 690
rect 1200 575 1205 675
rect 1240 575 1260 675
rect 1295 575 1300 675
rect 1200 560 1300 575
rect 1450 675 1550 690
rect 1450 575 1455 675
rect 1490 575 1510 675
rect 1545 575 1550 675
rect 1450 560 1550 575
rect 1700 675 1800 690
rect 1700 575 1705 675
rect 1740 575 1760 675
rect 1795 575 1800 675
rect 1700 560 1800 575
rect 1950 675 2050 690
rect 1950 575 1955 675
rect 1990 575 2010 675
rect 2045 575 2050 675
rect 1950 560 2050 575
rect 2200 675 2300 690
rect 2200 575 2205 675
rect 2240 575 2260 675
rect 2295 575 2300 675
rect 2200 560 2300 575
rect 2450 675 2550 690
rect 2450 575 2455 675
rect 2490 575 2510 675
rect 2545 575 2550 675
rect 2450 560 2550 575
rect 2700 675 2800 690
rect 2700 575 2705 675
rect 2740 575 2760 675
rect 2795 575 2800 675
rect 2700 560 2800 575
rect 2950 675 3050 690
rect 2950 575 2955 675
rect 2990 575 3010 675
rect 3045 575 3050 675
rect 2950 560 3050 575
rect 3200 675 3300 690
rect 3200 575 3205 675
rect 3240 575 3260 675
rect 3295 575 3300 675
rect 3200 560 3300 575
rect 3450 675 3550 690
rect 3450 575 3455 675
rect 3490 575 3510 675
rect 3545 575 3550 675
rect 3450 560 3550 575
rect 3700 675 3800 690
rect 3700 575 3705 675
rect 3740 575 3760 675
rect 3795 575 3800 675
rect 3700 560 3800 575
rect 3950 675 4000 690
rect 3950 575 3955 675
rect 3990 575 4000 675
rect 3950 560 4000 575
rect 0 550 60 560
rect 190 550 310 560
rect 440 550 560 560
rect 690 550 810 560
rect 940 550 1060 560
rect 1190 550 1310 560
rect 1440 550 1560 560
rect 1690 550 1810 560
rect 1940 550 2060 560
rect 2190 550 2310 560
rect 2440 550 2560 560
rect 2690 550 2810 560
rect 2940 550 3060 560
rect 3190 550 3310 560
rect 3440 550 3560 560
rect 3690 550 3810 560
rect 3940 550 4000 560
rect 0 545 4000 550
rect 0 510 75 545
rect 175 510 325 545
rect 425 510 575 545
rect 675 510 825 545
rect 925 510 1075 545
rect 1175 510 1325 545
rect 1425 510 1575 545
rect 1675 510 1825 545
rect 1925 510 2075 545
rect 2175 510 2325 545
rect 2425 510 2575 545
rect 2675 510 2825 545
rect 2925 510 3075 545
rect 3175 510 3325 545
rect 3425 510 3575 545
rect 3675 510 3825 545
rect 3925 510 4000 545
rect 0 490 4000 510
rect 0 455 75 490
rect 175 455 325 490
rect 425 455 575 490
rect 675 455 825 490
rect 925 455 1075 490
rect 1175 455 1325 490
rect 1425 455 1575 490
rect 1675 455 1825 490
rect 1925 455 2075 490
rect 2175 455 2325 490
rect 2425 455 2575 490
rect 2675 455 2825 490
rect 2925 455 3075 490
rect 3175 455 3325 490
rect 3425 455 3575 490
rect 3675 455 3825 490
rect 3925 455 4000 490
rect 0 450 4000 455
rect 0 440 60 450
rect 190 440 310 450
rect 440 440 560 450
rect 690 440 810 450
rect 940 440 1060 450
rect 1190 440 1310 450
rect 1440 440 1560 450
rect 1690 440 1810 450
rect 1940 440 2060 450
rect 2190 440 2310 450
rect 2440 440 2560 450
rect 2690 440 2810 450
rect 2940 440 3060 450
rect 3190 440 3310 450
rect 3440 440 3560 450
rect 3690 440 3810 450
rect 3940 440 4000 450
rect 0 425 50 440
rect 0 325 10 425
rect 45 325 50 425
rect 0 310 50 325
rect 200 425 300 440
rect 200 325 205 425
rect 240 325 260 425
rect 295 325 300 425
rect 200 310 300 325
rect 450 425 550 440
rect 450 325 455 425
rect 490 325 510 425
rect 545 325 550 425
rect 450 310 550 325
rect 700 425 800 440
rect 700 325 705 425
rect 740 325 760 425
rect 795 325 800 425
rect 700 310 800 325
rect 950 425 1050 440
rect 950 325 955 425
rect 990 325 1010 425
rect 1045 325 1050 425
rect 950 310 1050 325
rect 1200 425 1300 440
rect 1200 325 1205 425
rect 1240 325 1260 425
rect 1295 325 1300 425
rect 1200 310 1300 325
rect 1450 425 1550 440
rect 1450 325 1455 425
rect 1490 325 1510 425
rect 1545 325 1550 425
rect 1450 310 1550 325
rect 1700 425 1800 440
rect 1700 325 1705 425
rect 1740 325 1760 425
rect 1795 325 1800 425
rect 1700 310 1800 325
rect 1950 425 2050 440
rect 1950 325 1955 425
rect 1990 325 2010 425
rect 2045 325 2050 425
rect 1950 310 2050 325
rect 2200 425 2300 440
rect 2200 325 2205 425
rect 2240 325 2260 425
rect 2295 325 2300 425
rect 2200 310 2300 325
rect 2450 425 2550 440
rect 2450 325 2455 425
rect 2490 325 2510 425
rect 2545 325 2550 425
rect 2450 310 2550 325
rect 2700 425 2800 440
rect 2700 325 2705 425
rect 2740 325 2760 425
rect 2795 325 2800 425
rect 2700 310 2800 325
rect 2950 425 3050 440
rect 2950 325 2955 425
rect 2990 325 3010 425
rect 3045 325 3050 425
rect 2950 310 3050 325
rect 3200 425 3300 440
rect 3200 325 3205 425
rect 3240 325 3260 425
rect 3295 325 3300 425
rect 3200 310 3300 325
rect 3450 425 3550 440
rect 3450 325 3455 425
rect 3490 325 3510 425
rect 3545 325 3550 425
rect 3450 310 3550 325
rect 3700 425 3800 440
rect 3700 325 3705 425
rect 3740 325 3760 425
rect 3795 325 3800 425
rect 3700 310 3800 325
rect 3950 425 4000 440
rect 3950 325 3955 425
rect 3990 325 4000 425
rect 3950 310 4000 325
rect 0 300 60 310
rect 190 300 310 310
rect 440 300 560 310
rect 690 300 810 310
rect 940 300 1060 310
rect 1190 300 1310 310
rect 1440 300 1560 310
rect 1690 300 1810 310
rect 1940 300 2060 310
rect 2190 300 2310 310
rect 2440 300 2560 310
rect 2690 300 2810 310
rect 2940 300 3060 310
rect 3190 300 3310 310
rect 3440 300 3560 310
rect 3690 300 3810 310
rect 3940 300 4000 310
rect 0 295 4000 300
rect 0 260 75 295
rect 175 260 325 295
rect 425 260 575 295
rect 675 260 825 295
rect 925 260 1075 295
rect 1175 260 1325 295
rect 1425 260 1575 295
rect 1675 260 1825 295
rect 1925 260 2075 295
rect 2175 260 2325 295
rect 2425 260 2575 295
rect 2675 260 2825 295
rect 2925 260 3075 295
rect 3175 260 3325 295
rect 3425 260 3575 295
rect 3675 260 3825 295
rect 3925 260 4000 295
rect 0 240 4000 260
rect 0 205 75 240
rect 175 205 325 240
rect 425 205 575 240
rect 675 205 825 240
rect 925 205 1075 240
rect 1175 205 1325 240
rect 1425 205 1575 240
rect 1675 205 1825 240
rect 1925 205 2075 240
rect 2175 205 2325 240
rect 2425 205 2575 240
rect 2675 205 2825 240
rect 2925 205 3075 240
rect 3175 205 3325 240
rect 3425 205 3575 240
rect 3675 205 3825 240
rect 3925 205 4000 240
rect 0 200 4000 205
rect 0 190 60 200
rect 190 190 310 200
rect 440 190 560 200
rect 690 190 810 200
rect 940 190 1060 200
rect 1190 190 1310 200
rect 1440 190 1560 200
rect 1690 190 1810 200
rect 1940 190 2060 200
rect 2190 190 2310 200
rect 2440 190 2560 200
rect 2690 190 2810 200
rect 2940 190 3060 200
rect 3190 190 3310 200
rect 3440 190 3560 200
rect 3690 190 3810 200
rect 3940 190 4000 200
rect 0 175 50 190
rect 0 75 10 175
rect 45 75 50 175
rect 0 60 50 75
rect 200 175 300 190
rect 200 75 205 175
rect 240 75 260 175
rect 295 75 300 175
rect 200 60 300 75
rect 450 175 550 190
rect 450 75 455 175
rect 490 75 510 175
rect 545 75 550 175
rect 450 60 550 75
rect 700 175 800 190
rect 700 75 705 175
rect 740 75 760 175
rect 795 75 800 175
rect 700 60 800 75
rect 950 175 1050 190
rect 950 75 955 175
rect 990 75 1010 175
rect 1045 75 1050 175
rect 950 60 1050 75
rect 1200 175 1300 190
rect 1200 75 1205 175
rect 1240 75 1260 175
rect 1295 75 1300 175
rect 1200 60 1300 75
rect 1450 175 1550 190
rect 1450 75 1455 175
rect 1490 75 1510 175
rect 1545 75 1550 175
rect 1450 60 1550 75
rect 1700 175 1800 190
rect 1700 75 1705 175
rect 1740 75 1760 175
rect 1795 75 1800 175
rect 1700 60 1800 75
rect 1950 175 2050 190
rect 1950 75 1955 175
rect 1990 75 2010 175
rect 2045 75 2050 175
rect 1950 60 2050 75
rect 2200 175 2300 190
rect 2200 75 2205 175
rect 2240 75 2260 175
rect 2295 75 2300 175
rect 2200 60 2300 75
rect 2450 175 2550 190
rect 2450 75 2455 175
rect 2490 75 2510 175
rect 2545 75 2550 175
rect 2450 60 2550 75
rect 2700 175 2800 190
rect 2700 75 2705 175
rect 2740 75 2760 175
rect 2795 75 2800 175
rect 2700 60 2800 75
rect 2950 175 3050 190
rect 2950 75 2955 175
rect 2990 75 3010 175
rect 3045 75 3050 175
rect 2950 60 3050 75
rect 3200 175 3300 190
rect 3200 75 3205 175
rect 3240 75 3260 175
rect 3295 75 3300 175
rect 3200 60 3300 75
rect 3450 175 3550 190
rect 3450 75 3455 175
rect 3490 75 3510 175
rect 3545 75 3550 175
rect 3450 60 3550 75
rect 3700 175 3800 190
rect 3700 75 3705 175
rect 3740 75 3760 175
rect 3795 75 3800 175
rect 3700 60 3800 75
rect 3950 175 4000 190
rect 3950 75 3955 175
rect 3990 75 4000 175
rect 3950 60 4000 75
rect 0 50 60 60
rect 190 50 310 60
rect 440 50 560 60
rect 690 50 810 60
rect 940 50 1060 60
rect 1190 50 1310 60
rect 1440 50 1560 60
rect 1690 50 1810 60
rect 1940 50 2060 60
rect 2190 50 2310 60
rect 2440 50 2560 60
rect 2690 50 2810 60
rect 2940 50 3060 60
rect 3190 50 3310 60
rect 3440 50 3560 60
rect 3690 50 3810 60
rect 3940 50 4000 60
rect 0 45 4000 50
rect 0 10 75 45
rect 175 10 325 45
rect 425 10 575 45
rect 675 10 825 45
rect 925 10 1075 45
rect 1175 10 1325 45
rect 1425 10 1575 45
rect 1675 10 1825 45
rect 1925 10 2075 45
rect 2175 10 2325 45
rect 2425 10 2575 45
rect 2675 10 2825 45
rect 2925 10 3075 45
rect 3175 10 3325 45
rect 3425 10 3575 45
rect 3675 10 3825 45
rect 3925 10 4000 45
rect 0 0 4000 10
<< via1 >>
rect 75 3955 175 3990
rect 325 3955 425 3990
rect 575 3955 675 3990
rect 825 3955 925 3990
rect 1075 3955 1175 3990
rect 1325 3955 1425 3990
rect 1575 3955 1675 3990
rect 1825 3955 1925 3990
rect 2075 3955 2175 3990
rect 2325 3955 2425 3990
rect 2575 3955 2675 3990
rect 2825 3955 2925 3990
rect 3075 3955 3175 3990
rect 3325 3955 3425 3990
rect 3575 3955 3675 3990
rect 3825 3955 3925 3990
rect 10 3825 45 3925
rect 205 3825 240 3925
rect 260 3825 295 3925
rect 455 3825 490 3925
rect 510 3825 545 3925
rect 705 3825 740 3925
rect 760 3825 795 3925
rect 955 3825 990 3925
rect 1010 3825 1045 3925
rect 1205 3825 1240 3925
rect 1260 3825 1295 3925
rect 1455 3825 1490 3925
rect 1510 3825 1545 3925
rect 1705 3825 1740 3925
rect 1760 3825 1795 3925
rect 1955 3825 1990 3925
rect 2010 3825 2045 3925
rect 2205 3825 2240 3925
rect 2260 3825 2295 3925
rect 2455 3825 2490 3925
rect 2510 3825 2545 3925
rect 2705 3825 2740 3925
rect 2760 3825 2795 3925
rect 2955 3825 2990 3925
rect 3010 3825 3045 3925
rect 3205 3825 3240 3925
rect 3260 3825 3295 3925
rect 3455 3825 3490 3925
rect 3510 3825 3545 3925
rect 3705 3825 3740 3925
rect 3760 3825 3795 3925
rect 3955 3825 3990 3925
rect 75 3760 175 3795
rect 325 3760 425 3795
rect 575 3760 675 3795
rect 825 3760 925 3795
rect 1075 3760 1175 3795
rect 1325 3760 1425 3795
rect 1575 3760 1675 3795
rect 1825 3760 1925 3795
rect 2075 3760 2175 3795
rect 2325 3760 2425 3795
rect 2575 3760 2675 3795
rect 2825 3760 2925 3795
rect 3075 3760 3175 3795
rect 3325 3760 3425 3795
rect 3575 3760 3675 3795
rect 3825 3760 3925 3795
rect 75 3705 175 3740
rect 325 3705 425 3740
rect 575 3705 675 3740
rect 825 3705 925 3740
rect 1075 3705 1175 3740
rect 1325 3705 1425 3740
rect 1575 3705 1675 3740
rect 1825 3705 1925 3740
rect 2075 3705 2175 3740
rect 2325 3705 2425 3740
rect 2575 3705 2675 3740
rect 2825 3705 2925 3740
rect 3075 3705 3175 3740
rect 3325 3705 3425 3740
rect 3575 3705 3675 3740
rect 3825 3705 3925 3740
rect 10 3575 45 3675
rect 205 3575 240 3675
rect 260 3575 295 3675
rect 455 3575 490 3675
rect 510 3575 545 3675
rect 705 3575 740 3675
rect 760 3575 795 3675
rect 955 3575 990 3675
rect 1010 3575 1045 3675
rect 1205 3575 1240 3675
rect 1260 3575 1295 3675
rect 1455 3575 1490 3675
rect 1510 3575 1545 3675
rect 1705 3575 1740 3675
rect 1760 3575 1795 3675
rect 1955 3575 1990 3675
rect 2010 3575 2045 3675
rect 2205 3575 2240 3675
rect 2260 3575 2295 3675
rect 2455 3575 2490 3675
rect 2510 3575 2545 3675
rect 2705 3575 2740 3675
rect 2760 3575 2795 3675
rect 2955 3575 2990 3675
rect 3010 3575 3045 3675
rect 3205 3575 3240 3675
rect 3260 3575 3295 3675
rect 3455 3575 3490 3675
rect 3510 3575 3545 3675
rect 3705 3575 3740 3675
rect 3760 3575 3795 3675
rect 3955 3575 3990 3675
rect 75 3510 175 3545
rect 325 3510 425 3545
rect 575 3510 675 3545
rect 825 3510 925 3545
rect 1075 3510 1175 3545
rect 1325 3510 1425 3545
rect 1575 3510 1675 3545
rect 1825 3510 1925 3545
rect 2075 3510 2175 3545
rect 2325 3510 2425 3545
rect 2575 3510 2675 3545
rect 2825 3510 2925 3545
rect 3075 3510 3175 3545
rect 3325 3510 3425 3545
rect 3575 3510 3675 3545
rect 3825 3510 3925 3545
rect 75 3455 175 3490
rect 325 3455 425 3490
rect 575 3455 675 3490
rect 825 3455 925 3490
rect 1075 3455 1175 3490
rect 1325 3455 1425 3490
rect 1575 3455 1675 3490
rect 1825 3455 1925 3490
rect 2075 3455 2175 3490
rect 2325 3455 2425 3490
rect 2575 3455 2675 3490
rect 2825 3455 2925 3490
rect 3075 3455 3175 3490
rect 3325 3455 3425 3490
rect 3575 3455 3675 3490
rect 3825 3455 3925 3490
rect 10 3325 45 3425
rect 205 3325 240 3425
rect 260 3325 295 3425
rect 455 3325 490 3425
rect 510 3325 545 3425
rect 705 3325 740 3425
rect 760 3325 795 3425
rect 955 3325 990 3425
rect 1010 3325 1045 3425
rect 1205 3325 1240 3425
rect 1260 3325 1295 3425
rect 1455 3325 1490 3425
rect 1510 3325 1545 3425
rect 1705 3325 1740 3425
rect 1760 3325 1795 3425
rect 1955 3325 1990 3425
rect 2010 3325 2045 3425
rect 2205 3325 2240 3425
rect 2260 3325 2295 3425
rect 2455 3325 2490 3425
rect 2510 3325 2545 3425
rect 2705 3325 2740 3425
rect 2760 3325 2795 3425
rect 2955 3325 2990 3425
rect 3010 3325 3045 3425
rect 3205 3325 3240 3425
rect 3260 3325 3295 3425
rect 3455 3325 3490 3425
rect 3510 3325 3545 3425
rect 3705 3325 3740 3425
rect 3760 3325 3795 3425
rect 3955 3325 3990 3425
rect 75 3260 175 3295
rect 325 3260 425 3295
rect 575 3260 675 3295
rect 825 3260 925 3295
rect 1075 3260 1175 3295
rect 1325 3260 1425 3295
rect 1575 3260 1675 3295
rect 1825 3260 1925 3295
rect 2075 3260 2175 3295
rect 2325 3260 2425 3295
rect 2575 3260 2675 3295
rect 2825 3260 2925 3295
rect 3075 3260 3175 3295
rect 3325 3260 3425 3295
rect 3575 3260 3675 3295
rect 3825 3260 3925 3295
rect 75 3205 175 3240
rect 325 3205 425 3240
rect 575 3205 675 3240
rect 825 3205 925 3240
rect 1075 3205 1175 3240
rect 1325 3205 1425 3240
rect 1575 3205 1675 3240
rect 1825 3205 1925 3240
rect 2075 3205 2175 3240
rect 2325 3205 2425 3240
rect 2575 3205 2675 3240
rect 2825 3205 2925 3240
rect 3075 3205 3175 3240
rect 3325 3205 3425 3240
rect 3575 3205 3675 3240
rect 3825 3205 3925 3240
rect 10 3075 45 3175
rect 205 3075 240 3175
rect 260 3075 295 3175
rect 455 3075 490 3175
rect 510 3075 545 3175
rect 705 3075 740 3175
rect 760 3075 795 3175
rect 955 3075 990 3175
rect 1010 3075 1045 3175
rect 1205 3075 1240 3175
rect 1260 3075 1295 3175
rect 1455 3075 1490 3175
rect 1510 3075 1545 3175
rect 1705 3075 1740 3175
rect 1760 3075 1795 3175
rect 1955 3075 1990 3175
rect 2010 3075 2045 3175
rect 2205 3075 2240 3175
rect 2260 3075 2295 3175
rect 2455 3075 2490 3175
rect 2510 3075 2545 3175
rect 2705 3075 2740 3175
rect 2760 3075 2795 3175
rect 2955 3075 2990 3175
rect 3010 3075 3045 3175
rect 3205 3075 3240 3175
rect 3260 3075 3295 3175
rect 3455 3075 3490 3175
rect 3510 3075 3545 3175
rect 3705 3075 3740 3175
rect 3760 3075 3795 3175
rect 3955 3075 3990 3175
rect 75 3010 175 3045
rect 325 3010 425 3045
rect 575 3010 675 3045
rect 825 3010 925 3045
rect 1075 3010 1175 3045
rect 1325 3010 1425 3045
rect 1575 3010 1675 3045
rect 1825 3010 1925 3045
rect 2075 3010 2175 3045
rect 2325 3010 2425 3045
rect 2575 3010 2675 3045
rect 2825 3010 2925 3045
rect 3075 3010 3175 3045
rect 3325 3010 3425 3045
rect 3575 3010 3675 3045
rect 3825 3010 3925 3045
rect 75 2955 175 2990
rect 325 2955 425 2990
rect 575 2955 675 2990
rect 825 2955 925 2990
rect 1075 2955 1175 2990
rect 1325 2955 1425 2990
rect 1575 2955 1675 2990
rect 1825 2955 1925 2990
rect 2075 2955 2175 2990
rect 2325 2955 2425 2990
rect 2575 2955 2675 2990
rect 2825 2955 2925 2990
rect 3075 2955 3175 2990
rect 3325 2955 3425 2990
rect 3575 2955 3675 2990
rect 3825 2955 3925 2990
rect 10 2825 45 2925
rect 205 2825 240 2925
rect 260 2825 295 2925
rect 455 2825 490 2925
rect 510 2825 545 2925
rect 705 2825 740 2925
rect 760 2825 795 2925
rect 955 2825 990 2925
rect 1010 2825 1045 2925
rect 1205 2825 1240 2925
rect 1260 2825 1295 2925
rect 1455 2825 1490 2925
rect 1510 2825 1545 2925
rect 1705 2825 1740 2925
rect 1760 2825 1795 2925
rect 1955 2825 1990 2925
rect 2010 2825 2045 2925
rect 2205 2825 2240 2925
rect 2260 2825 2295 2925
rect 2455 2825 2490 2925
rect 2510 2825 2545 2925
rect 2705 2825 2740 2925
rect 2760 2825 2795 2925
rect 2955 2825 2990 2925
rect 3010 2825 3045 2925
rect 3205 2825 3240 2925
rect 3260 2825 3295 2925
rect 3455 2825 3490 2925
rect 3510 2825 3545 2925
rect 3705 2825 3740 2925
rect 3760 2825 3795 2925
rect 3955 2825 3990 2925
rect 75 2760 175 2795
rect 325 2760 425 2795
rect 575 2760 675 2795
rect 825 2760 925 2795
rect 1075 2760 1175 2795
rect 1325 2760 1425 2795
rect 1575 2760 1675 2795
rect 1825 2760 1925 2795
rect 2075 2760 2175 2795
rect 2325 2760 2425 2795
rect 2575 2760 2675 2795
rect 2825 2760 2925 2795
rect 3075 2760 3175 2795
rect 3325 2760 3425 2795
rect 3575 2760 3675 2795
rect 3825 2760 3925 2795
rect 75 2705 175 2740
rect 325 2705 425 2740
rect 575 2705 675 2740
rect 825 2705 925 2740
rect 1075 2705 1175 2740
rect 1325 2705 1425 2740
rect 1575 2705 1675 2740
rect 1825 2705 1925 2740
rect 2075 2705 2175 2740
rect 2325 2705 2425 2740
rect 2575 2705 2675 2740
rect 2825 2705 2925 2740
rect 3075 2705 3175 2740
rect 3325 2705 3425 2740
rect 3575 2705 3675 2740
rect 3825 2705 3925 2740
rect 10 2575 45 2675
rect 205 2575 240 2675
rect 260 2575 295 2675
rect 455 2575 490 2675
rect 510 2575 545 2675
rect 705 2575 740 2675
rect 760 2575 795 2675
rect 955 2575 990 2675
rect 1010 2575 1045 2675
rect 1205 2575 1240 2675
rect 1260 2575 1295 2675
rect 1455 2575 1490 2675
rect 1510 2575 1545 2675
rect 1705 2575 1740 2675
rect 1760 2575 1795 2675
rect 1955 2575 1990 2675
rect 2010 2575 2045 2675
rect 2205 2575 2240 2675
rect 2260 2575 2295 2675
rect 2455 2575 2490 2675
rect 2510 2575 2545 2675
rect 2705 2575 2740 2675
rect 2760 2575 2795 2675
rect 2955 2575 2990 2675
rect 3010 2575 3045 2675
rect 3205 2575 3240 2675
rect 3260 2575 3295 2675
rect 3455 2575 3490 2675
rect 3510 2575 3545 2675
rect 3705 2575 3740 2675
rect 3760 2575 3795 2675
rect 3955 2575 3990 2675
rect 75 2510 175 2545
rect 325 2510 425 2545
rect 575 2510 675 2545
rect 825 2510 925 2545
rect 1075 2510 1175 2545
rect 1325 2510 1425 2545
rect 1575 2510 1675 2545
rect 1825 2510 1925 2545
rect 2075 2510 2175 2545
rect 2325 2510 2425 2545
rect 2575 2510 2675 2545
rect 2825 2510 2925 2545
rect 3075 2510 3175 2545
rect 3325 2510 3425 2545
rect 3575 2510 3675 2545
rect 3825 2510 3925 2545
rect 75 2455 175 2490
rect 325 2455 425 2490
rect 575 2455 675 2490
rect 825 2455 925 2490
rect 1075 2455 1175 2490
rect 1325 2455 1425 2490
rect 1575 2455 1675 2490
rect 1825 2455 1925 2490
rect 2075 2455 2175 2490
rect 2325 2455 2425 2490
rect 2575 2455 2675 2490
rect 2825 2455 2925 2490
rect 3075 2455 3175 2490
rect 3325 2455 3425 2490
rect 3575 2455 3675 2490
rect 3825 2455 3925 2490
rect 10 2325 45 2425
rect 205 2325 240 2425
rect 260 2325 295 2425
rect 455 2325 490 2425
rect 510 2325 545 2425
rect 705 2325 740 2425
rect 760 2325 795 2425
rect 955 2325 990 2425
rect 1010 2325 1045 2425
rect 1205 2325 1240 2425
rect 1260 2325 1295 2425
rect 1455 2325 1490 2425
rect 1510 2325 1545 2425
rect 1705 2325 1740 2425
rect 1760 2325 1795 2425
rect 1955 2325 1990 2425
rect 2010 2325 2045 2425
rect 2205 2325 2240 2425
rect 2260 2325 2295 2425
rect 2455 2325 2490 2425
rect 2510 2325 2545 2425
rect 2705 2325 2740 2425
rect 2760 2325 2795 2425
rect 2955 2325 2990 2425
rect 3010 2325 3045 2425
rect 3205 2325 3240 2425
rect 3260 2325 3295 2425
rect 3455 2325 3490 2425
rect 3510 2325 3545 2425
rect 3705 2325 3740 2425
rect 3760 2325 3795 2425
rect 3955 2325 3990 2425
rect 75 2260 175 2295
rect 325 2260 425 2295
rect 575 2260 675 2295
rect 825 2260 925 2295
rect 1075 2260 1175 2295
rect 1325 2260 1425 2295
rect 1575 2260 1675 2295
rect 1825 2260 1925 2295
rect 2075 2260 2175 2295
rect 2325 2260 2425 2295
rect 2575 2260 2675 2295
rect 2825 2260 2925 2295
rect 3075 2260 3175 2295
rect 3325 2260 3425 2295
rect 3575 2260 3675 2295
rect 3825 2260 3925 2295
rect 75 2205 175 2240
rect 325 2205 425 2240
rect 575 2205 675 2240
rect 825 2205 925 2240
rect 1075 2205 1175 2240
rect 1325 2205 1425 2240
rect 1575 2205 1675 2240
rect 1825 2205 1925 2240
rect 2075 2205 2175 2240
rect 2325 2205 2425 2240
rect 2575 2205 2675 2240
rect 2825 2205 2925 2240
rect 3075 2205 3175 2240
rect 3325 2205 3425 2240
rect 3575 2205 3675 2240
rect 3825 2205 3925 2240
rect 10 2075 45 2175
rect 205 2075 240 2175
rect 260 2075 295 2175
rect 455 2075 490 2175
rect 510 2075 545 2175
rect 705 2075 740 2175
rect 760 2075 795 2175
rect 955 2075 990 2175
rect 1010 2075 1045 2175
rect 1205 2075 1240 2175
rect 1260 2075 1295 2175
rect 1455 2075 1490 2175
rect 1510 2075 1545 2175
rect 1705 2075 1740 2175
rect 1760 2075 1795 2175
rect 1955 2075 1990 2175
rect 2010 2075 2045 2175
rect 2205 2075 2240 2175
rect 2260 2075 2295 2175
rect 2455 2075 2490 2175
rect 2510 2075 2545 2175
rect 2705 2075 2740 2175
rect 2760 2075 2795 2175
rect 2955 2075 2990 2175
rect 3010 2075 3045 2175
rect 3205 2075 3240 2175
rect 3260 2075 3295 2175
rect 3455 2075 3490 2175
rect 3510 2075 3545 2175
rect 3705 2075 3740 2175
rect 3760 2075 3795 2175
rect 3955 2075 3990 2175
rect 75 2010 175 2045
rect 325 2010 425 2045
rect 575 2010 675 2045
rect 825 2010 925 2045
rect 1075 2010 1175 2045
rect 1325 2010 1425 2045
rect 1575 2010 1675 2045
rect 1825 2010 1925 2045
rect 2075 2010 2175 2045
rect 2325 2010 2425 2045
rect 2575 2010 2675 2045
rect 2825 2010 2925 2045
rect 3075 2010 3175 2045
rect 3325 2010 3425 2045
rect 3575 2010 3675 2045
rect 3825 2010 3925 2045
rect 75 1955 175 1990
rect 325 1955 425 1990
rect 575 1955 675 1990
rect 825 1955 925 1990
rect 1075 1955 1175 1990
rect 1325 1955 1425 1990
rect 1575 1955 1675 1990
rect 1825 1955 1925 1990
rect 2075 1955 2175 1990
rect 2325 1955 2425 1990
rect 2575 1955 2675 1990
rect 2825 1955 2925 1990
rect 3075 1955 3175 1990
rect 3325 1955 3425 1990
rect 3575 1955 3675 1990
rect 3825 1955 3925 1990
rect 10 1825 45 1925
rect 205 1825 240 1925
rect 260 1825 295 1925
rect 455 1825 490 1925
rect 510 1825 545 1925
rect 705 1825 740 1925
rect 760 1825 795 1925
rect 955 1825 990 1925
rect 1010 1825 1045 1925
rect 1205 1825 1240 1925
rect 1260 1825 1295 1925
rect 1455 1825 1490 1925
rect 1510 1825 1545 1925
rect 1705 1825 1740 1925
rect 1760 1825 1795 1925
rect 1955 1825 1990 1925
rect 2010 1825 2045 1925
rect 2205 1825 2240 1925
rect 2260 1825 2295 1925
rect 2455 1825 2490 1925
rect 2510 1825 2545 1925
rect 2705 1825 2740 1925
rect 2760 1825 2795 1925
rect 2955 1825 2990 1925
rect 3010 1825 3045 1925
rect 3205 1825 3240 1925
rect 3260 1825 3295 1925
rect 3455 1825 3490 1925
rect 3510 1825 3545 1925
rect 3705 1825 3740 1925
rect 3760 1825 3795 1925
rect 3955 1825 3990 1925
rect 75 1760 175 1795
rect 325 1760 425 1795
rect 575 1760 675 1795
rect 825 1760 925 1795
rect 1075 1760 1175 1795
rect 1325 1760 1425 1795
rect 1575 1760 1675 1795
rect 1825 1760 1925 1795
rect 2075 1760 2175 1795
rect 2325 1760 2425 1795
rect 2575 1760 2675 1795
rect 2825 1760 2925 1795
rect 3075 1760 3175 1795
rect 3325 1760 3425 1795
rect 3575 1760 3675 1795
rect 3825 1760 3925 1795
rect 75 1705 175 1740
rect 325 1705 425 1740
rect 575 1705 675 1740
rect 825 1705 925 1740
rect 1075 1705 1175 1740
rect 1325 1705 1425 1740
rect 1575 1705 1675 1740
rect 1825 1705 1925 1740
rect 2075 1705 2175 1740
rect 2325 1705 2425 1740
rect 2575 1705 2675 1740
rect 2825 1705 2925 1740
rect 3075 1705 3175 1740
rect 3325 1705 3425 1740
rect 3575 1705 3675 1740
rect 3825 1705 3925 1740
rect 10 1575 45 1675
rect 205 1575 240 1675
rect 260 1575 295 1675
rect 455 1575 490 1675
rect 510 1575 545 1675
rect 705 1575 740 1675
rect 760 1575 795 1675
rect 955 1575 990 1675
rect 1010 1575 1045 1675
rect 1205 1575 1240 1675
rect 1260 1575 1295 1675
rect 1455 1575 1490 1675
rect 1510 1575 1545 1675
rect 1705 1575 1740 1675
rect 1760 1575 1795 1675
rect 1955 1575 1990 1675
rect 2010 1575 2045 1675
rect 2205 1575 2240 1675
rect 2260 1575 2295 1675
rect 2455 1575 2490 1675
rect 2510 1575 2545 1675
rect 2705 1575 2740 1675
rect 2760 1575 2795 1675
rect 2955 1575 2990 1675
rect 3010 1575 3045 1675
rect 3205 1575 3240 1675
rect 3260 1575 3295 1675
rect 3455 1575 3490 1675
rect 3510 1575 3545 1675
rect 3705 1575 3740 1675
rect 3760 1575 3795 1675
rect 3955 1575 3990 1675
rect 75 1510 175 1545
rect 325 1510 425 1545
rect 575 1510 675 1545
rect 825 1510 925 1545
rect 1075 1510 1175 1545
rect 1325 1510 1425 1545
rect 1575 1510 1675 1545
rect 1825 1510 1925 1545
rect 2075 1510 2175 1545
rect 2325 1510 2425 1545
rect 2575 1510 2675 1545
rect 2825 1510 2925 1545
rect 3075 1510 3175 1545
rect 3325 1510 3425 1545
rect 3575 1510 3675 1545
rect 3825 1510 3925 1545
rect 75 1455 175 1490
rect 325 1455 425 1490
rect 575 1455 675 1490
rect 825 1455 925 1490
rect 1075 1455 1175 1490
rect 1325 1455 1425 1490
rect 1575 1455 1675 1490
rect 1825 1455 1925 1490
rect 2075 1455 2175 1490
rect 2325 1455 2425 1490
rect 2575 1455 2675 1490
rect 2825 1455 2925 1490
rect 3075 1455 3175 1490
rect 3325 1455 3425 1490
rect 3575 1455 3675 1490
rect 3825 1455 3925 1490
rect 10 1325 45 1425
rect 205 1325 240 1425
rect 260 1325 295 1425
rect 455 1325 490 1425
rect 510 1325 545 1425
rect 705 1325 740 1425
rect 760 1325 795 1425
rect 955 1325 990 1425
rect 1010 1325 1045 1425
rect 1205 1325 1240 1425
rect 1260 1325 1295 1425
rect 1455 1325 1490 1425
rect 1510 1325 1545 1425
rect 1705 1325 1740 1425
rect 1760 1325 1795 1425
rect 1955 1325 1990 1425
rect 2010 1325 2045 1425
rect 2205 1325 2240 1425
rect 2260 1325 2295 1425
rect 2455 1325 2490 1425
rect 2510 1325 2545 1425
rect 2705 1325 2740 1425
rect 2760 1325 2795 1425
rect 2955 1325 2990 1425
rect 3010 1325 3045 1425
rect 3205 1325 3240 1425
rect 3260 1325 3295 1425
rect 3455 1325 3490 1425
rect 3510 1325 3545 1425
rect 3705 1325 3740 1425
rect 3760 1325 3795 1425
rect 3955 1325 3990 1425
rect 75 1260 175 1295
rect 325 1260 425 1295
rect 575 1260 675 1295
rect 825 1260 925 1295
rect 1075 1260 1175 1295
rect 1325 1260 1425 1295
rect 1575 1260 1675 1295
rect 1825 1260 1925 1295
rect 2075 1260 2175 1295
rect 2325 1260 2425 1295
rect 2575 1260 2675 1295
rect 2825 1260 2925 1295
rect 3075 1260 3175 1295
rect 3325 1260 3425 1295
rect 3575 1260 3675 1295
rect 3825 1260 3925 1295
rect 75 1205 175 1240
rect 325 1205 425 1240
rect 575 1205 675 1240
rect 825 1205 925 1240
rect 1075 1205 1175 1240
rect 1325 1205 1425 1240
rect 1575 1205 1675 1240
rect 1825 1205 1925 1240
rect 2075 1205 2175 1240
rect 2325 1205 2425 1240
rect 2575 1205 2675 1240
rect 2825 1205 2925 1240
rect 3075 1205 3175 1240
rect 3325 1205 3425 1240
rect 3575 1205 3675 1240
rect 3825 1205 3925 1240
rect 10 1075 45 1175
rect 205 1075 240 1175
rect 260 1075 295 1175
rect 455 1075 490 1175
rect 510 1075 545 1175
rect 705 1075 740 1175
rect 760 1075 795 1175
rect 955 1075 990 1175
rect 1010 1075 1045 1175
rect 1205 1075 1240 1175
rect 1260 1075 1295 1175
rect 1455 1075 1490 1175
rect 1510 1075 1545 1175
rect 1705 1075 1740 1175
rect 1760 1075 1795 1175
rect 1955 1075 1990 1175
rect 2010 1075 2045 1175
rect 2205 1075 2240 1175
rect 2260 1075 2295 1175
rect 2455 1075 2490 1175
rect 2510 1075 2545 1175
rect 2705 1075 2740 1175
rect 2760 1075 2795 1175
rect 2955 1075 2990 1175
rect 3010 1075 3045 1175
rect 3205 1075 3240 1175
rect 3260 1075 3295 1175
rect 3455 1075 3490 1175
rect 3510 1075 3545 1175
rect 3705 1075 3740 1175
rect 3760 1075 3795 1175
rect 3955 1075 3990 1175
rect 75 1010 175 1045
rect 325 1010 425 1045
rect 575 1010 675 1045
rect 825 1010 925 1045
rect 1075 1010 1175 1045
rect 1325 1010 1425 1045
rect 1575 1010 1675 1045
rect 1825 1010 1925 1045
rect 2075 1010 2175 1045
rect 2325 1010 2425 1045
rect 2575 1010 2675 1045
rect 2825 1010 2925 1045
rect 3075 1010 3175 1045
rect 3325 1010 3425 1045
rect 3575 1010 3675 1045
rect 3825 1010 3925 1045
rect 75 955 175 990
rect 325 955 425 990
rect 575 955 675 990
rect 825 955 925 990
rect 1075 955 1175 990
rect 1325 955 1425 990
rect 1575 955 1675 990
rect 1825 955 1925 990
rect 2075 955 2175 990
rect 2325 955 2425 990
rect 2575 955 2675 990
rect 2825 955 2925 990
rect 3075 955 3175 990
rect 3325 955 3425 990
rect 3575 955 3675 990
rect 3825 955 3925 990
rect 10 825 45 925
rect 205 825 240 925
rect 260 825 295 925
rect 455 825 490 925
rect 510 825 545 925
rect 705 825 740 925
rect 760 825 795 925
rect 955 825 990 925
rect 1010 825 1045 925
rect 1205 825 1240 925
rect 1260 825 1295 925
rect 1455 825 1490 925
rect 1510 825 1545 925
rect 1705 825 1740 925
rect 1760 825 1795 925
rect 1955 825 1990 925
rect 2010 825 2045 925
rect 2205 825 2240 925
rect 2260 825 2295 925
rect 2455 825 2490 925
rect 2510 825 2545 925
rect 2705 825 2740 925
rect 2760 825 2795 925
rect 2955 825 2990 925
rect 3010 825 3045 925
rect 3205 825 3240 925
rect 3260 825 3295 925
rect 3455 825 3490 925
rect 3510 825 3545 925
rect 3705 825 3740 925
rect 3760 825 3795 925
rect 3955 825 3990 925
rect 75 760 175 795
rect 325 760 425 795
rect 575 760 675 795
rect 825 760 925 795
rect 1075 760 1175 795
rect 1325 760 1425 795
rect 1575 760 1675 795
rect 1825 760 1925 795
rect 2075 760 2175 795
rect 2325 760 2425 795
rect 2575 760 2675 795
rect 2825 760 2925 795
rect 3075 760 3175 795
rect 3325 760 3425 795
rect 3575 760 3675 795
rect 3825 760 3925 795
rect 75 705 175 740
rect 325 705 425 740
rect 575 705 675 740
rect 825 705 925 740
rect 1075 705 1175 740
rect 1325 705 1425 740
rect 1575 705 1675 740
rect 1825 705 1925 740
rect 2075 705 2175 740
rect 2325 705 2425 740
rect 2575 705 2675 740
rect 2825 705 2925 740
rect 3075 705 3175 740
rect 3325 705 3425 740
rect 3575 705 3675 740
rect 3825 705 3925 740
rect 10 575 45 675
rect 205 575 240 675
rect 260 575 295 675
rect 455 575 490 675
rect 510 575 545 675
rect 705 575 740 675
rect 760 575 795 675
rect 955 575 990 675
rect 1010 575 1045 675
rect 1205 575 1240 675
rect 1260 575 1295 675
rect 1455 575 1490 675
rect 1510 575 1545 675
rect 1705 575 1740 675
rect 1760 575 1795 675
rect 1955 575 1990 675
rect 2010 575 2045 675
rect 2205 575 2240 675
rect 2260 575 2295 675
rect 2455 575 2490 675
rect 2510 575 2545 675
rect 2705 575 2740 675
rect 2760 575 2795 675
rect 2955 575 2990 675
rect 3010 575 3045 675
rect 3205 575 3240 675
rect 3260 575 3295 675
rect 3455 575 3490 675
rect 3510 575 3545 675
rect 3705 575 3740 675
rect 3760 575 3795 675
rect 3955 575 3990 675
rect 75 510 175 545
rect 325 510 425 545
rect 575 510 675 545
rect 825 510 925 545
rect 1075 510 1175 545
rect 1325 510 1425 545
rect 1575 510 1675 545
rect 1825 510 1925 545
rect 2075 510 2175 545
rect 2325 510 2425 545
rect 2575 510 2675 545
rect 2825 510 2925 545
rect 3075 510 3175 545
rect 3325 510 3425 545
rect 3575 510 3675 545
rect 3825 510 3925 545
rect 75 455 175 490
rect 325 455 425 490
rect 575 455 675 490
rect 825 455 925 490
rect 1075 455 1175 490
rect 1325 455 1425 490
rect 1575 455 1675 490
rect 1825 455 1925 490
rect 2075 455 2175 490
rect 2325 455 2425 490
rect 2575 455 2675 490
rect 2825 455 2925 490
rect 3075 455 3175 490
rect 3325 455 3425 490
rect 3575 455 3675 490
rect 3825 455 3925 490
rect 10 325 45 425
rect 205 325 240 425
rect 260 325 295 425
rect 455 325 490 425
rect 510 325 545 425
rect 705 325 740 425
rect 760 325 795 425
rect 955 325 990 425
rect 1010 325 1045 425
rect 1205 325 1240 425
rect 1260 325 1295 425
rect 1455 325 1490 425
rect 1510 325 1545 425
rect 1705 325 1740 425
rect 1760 325 1795 425
rect 1955 325 1990 425
rect 2010 325 2045 425
rect 2205 325 2240 425
rect 2260 325 2295 425
rect 2455 325 2490 425
rect 2510 325 2545 425
rect 2705 325 2740 425
rect 2760 325 2795 425
rect 2955 325 2990 425
rect 3010 325 3045 425
rect 3205 325 3240 425
rect 3260 325 3295 425
rect 3455 325 3490 425
rect 3510 325 3545 425
rect 3705 325 3740 425
rect 3760 325 3795 425
rect 3955 325 3990 425
rect 75 260 175 295
rect 325 260 425 295
rect 575 260 675 295
rect 825 260 925 295
rect 1075 260 1175 295
rect 1325 260 1425 295
rect 1575 260 1675 295
rect 1825 260 1925 295
rect 2075 260 2175 295
rect 2325 260 2425 295
rect 2575 260 2675 295
rect 2825 260 2925 295
rect 3075 260 3175 295
rect 3325 260 3425 295
rect 3575 260 3675 295
rect 3825 260 3925 295
rect 75 205 175 240
rect 325 205 425 240
rect 575 205 675 240
rect 825 205 925 240
rect 1075 205 1175 240
rect 1325 205 1425 240
rect 1575 205 1675 240
rect 1825 205 1925 240
rect 2075 205 2175 240
rect 2325 205 2425 240
rect 2575 205 2675 240
rect 2825 205 2925 240
rect 3075 205 3175 240
rect 3325 205 3425 240
rect 3575 205 3675 240
rect 3825 205 3925 240
rect 10 75 45 175
rect 205 75 240 175
rect 260 75 295 175
rect 455 75 490 175
rect 510 75 545 175
rect 705 75 740 175
rect 760 75 795 175
rect 955 75 990 175
rect 1010 75 1045 175
rect 1205 75 1240 175
rect 1260 75 1295 175
rect 1455 75 1490 175
rect 1510 75 1545 175
rect 1705 75 1740 175
rect 1760 75 1795 175
rect 1955 75 1990 175
rect 2010 75 2045 175
rect 2205 75 2240 175
rect 2260 75 2295 175
rect 2455 75 2490 175
rect 2510 75 2545 175
rect 2705 75 2740 175
rect 2760 75 2795 175
rect 2955 75 2990 175
rect 3010 75 3045 175
rect 3205 75 3240 175
rect 3260 75 3295 175
rect 3455 75 3490 175
rect 3510 75 3545 175
rect 3705 75 3740 175
rect 3760 75 3795 175
rect 3955 75 3990 175
rect 75 10 175 45
rect 325 10 425 45
rect 575 10 675 45
rect 825 10 925 45
rect 1075 10 1175 45
rect 1325 10 1425 45
rect 1575 10 1675 45
rect 1825 10 1925 45
rect 2075 10 2175 45
rect 2325 10 2425 45
rect 2575 10 2675 45
rect 2825 10 2925 45
rect 3075 10 3175 45
rect 3325 10 3425 45
rect 3575 10 3675 45
rect 3825 10 3925 45
<< metal2 >>
rect 70 3990 180 4000
rect 70 3955 75 3990
rect 175 3955 180 3990
rect 70 3930 180 3955
rect 320 3990 430 4000
rect 320 3955 325 3990
rect 425 3955 430 3990
rect 320 3930 430 3955
rect 570 3990 680 4000
rect 570 3955 575 3990
rect 675 3955 680 3990
rect 570 3930 680 3955
rect 820 3990 930 4000
rect 820 3955 825 3990
rect 925 3955 930 3990
rect 820 3930 930 3955
rect 1070 3990 1180 4000
rect 1070 3955 1075 3990
rect 1175 3955 1180 3990
rect 1070 3930 1180 3955
rect 1320 3990 1430 4000
rect 1320 3955 1325 3990
rect 1425 3955 1430 3990
rect 1320 3930 1430 3955
rect 1570 3990 1680 4000
rect 1570 3955 1575 3990
rect 1675 3955 1680 3990
rect 1570 3930 1680 3955
rect 1820 3990 1930 4000
rect 1820 3955 1825 3990
rect 1925 3955 1930 3990
rect 1820 3930 1930 3955
rect 2070 3990 2180 4000
rect 2070 3955 2075 3990
rect 2175 3955 2180 3990
rect 2070 3930 2180 3955
rect 2320 3990 2430 4000
rect 2320 3955 2325 3990
rect 2425 3955 2430 3990
rect 2320 3930 2430 3955
rect 2570 3990 2680 4000
rect 2570 3955 2575 3990
rect 2675 3955 2680 3990
rect 2570 3930 2680 3955
rect 2820 3990 2930 4000
rect 2820 3955 2825 3990
rect 2925 3955 2930 3990
rect 2820 3930 2930 3955
rect 3070 3990 3180 4000
rect 3070 3955 3075 3990
rect 3175 3955 3180 3990
rect 3070 3930 3180 3955
rect 3320 3990 3430 4000
rect 3320 3955 3325 3990
rect 3425 3955 3430 3990
rect 3320 3930 3430 3955
rect 3570 3990 3680 4000
rect 3570 3955 3575 3990
rect 3675 3955 3680 3990
rect 3570 3930 3680 3955
rect 3820 3990 3930 4000
rect 3820 3955 3825 3990
rect 3925 3955 3930 3990
rect 3820 3930 3930 3955
rect 0 3925 4000 3930
rect 0 3825 10 3925
rect 45 3825 205 3925
rect 240 3825 260 3925
rect 295 3825 455 3925
rect 490 3825 510 3925
rect 545 3825 705 3925
rect 740 3825 760 3925
rect 795 3825 955 3925
rect 990 3825 1010 3925
rect 1045 3825 1205 3925
rect 1240 3825 1260 3925
rect 1295 3825 1455 3925
rect 1490 3825 1510 3925
rect 1545 3825 1705 3925
rect 1740 3825 1760 3925
rect 1795 3825 1955 3925
rect 1990 3825 2010 3925
rect 2045 3825 2205 3925
rect 2240 3825 2260 3925
rect 2295 3825 2455 3925
rect 2490 3825 2510 3925
rect 2545 3825 2705 3925
rect 2740 3825 2760 3925
rect 2795 3825 2955 3925
rect 2990 3825 3010 3925
rect 3045 3825 3205 3925
rect 3240 3825 3260 3925
rect 3295 3825 3455 3925
rect 3490 3825 3510 3925
rect 3545 3825 3705 3925
rect 3740 3825 3760 3925
rect 3795 3825 3955 3925
rect 3990 3825 4000 3925
rect 0 3820 4000 3825
rect 70 3795 180 3820
rect 70 3760 75 3795
rect 175 3760 180 3795
rect 70 3740 180 3760
rect 70 3705 75 3740
rect 175 3705 180 3740
rect 70 3680 180 3705
rect 320 3795 430 3820
rect 320 3760 325 3795
rect 425 3760 430 3795
rect 320 3740 430 3760
rect 320 3705 325 3740
rect 425 3705 430 3740
rect 320 3680 430 3705
rect 570 3795 680 3820
rect 570 3760 575 3795
rect 675 3760 680 3795
rect 570 3740 680 3760
rect 570 3705 575 3740
rect 675 3705 680 3740
rect 570 3680 680 3705
rect 820 3795 930 3820
rect 820 3760 825 3795
rect 925 3760 930 3795
rect 820 3740 930 3760
rect 820 3705 825 3740
rect 925 3705 930 3740
rect 820 3680 930 3705
rect 1070 3795 1180 3820
rect 1070 3760 1075 3795
rect 1175 3760 1180 3795
rect 1070 3740 1180 3760
rect 1070 3705 1075 3740
rect 1175 3705 1180 3740
rect 1070 3680 1180 3705
rect 1320 3795 1430 3820
rect 1320 3760 1325 3795
rect 1425 3760 1430 3795
rect 1320 3740 1430 3760
rect 1320 3705 1325 3740
rect 1425 3705 1430 3740
rect 1320 3680 1430 3705
rect 1570 3795 1680 3820
rect 1570 3760 1575 3795
rect 1675 3760 1680 3795
rect 1570 3740 1680 3760
rect 1570 3705 1575 3740
rect 1675 3705 1680 3740
rect 1570 3680 1680 3705
rect 1820 3795 1930 3820
rect 1820 3760 1825 3795
rect 1925 3760 1930 3795
rect 1820 3740 1930 3760
rect 1820 3705 1825 3740
rect 1925 3705 1930 3740
rect 1820 3680 1930 3705
rect 2070 3795 2180 3820
rect 2070 3760 2075 3795
rect 2175 3760 2180 3795
rect 2070 3740 2180 3760
rect 2070 3705 2075 3740
rect 2175 3705 2180 3740
rect 2070 3680 2180 3705
rect 2320 3795 2430 3820
rect 2320 3760 2325 3795
rect 2425 3760 2430 3795
rect 2320 3740 2430 3760
rect 2320 3705 2325 3740
rect 2425 3705 2430 3740
rect 2320 3680 2430 3705
rect 2570 3795 2680 3820
rect 2570 3760 2575 3795
rect 2675 3760 2680 3795
rect 2570 3740 2680 3760
rect 2570 3705 2575 3740
rect 2675 3705 2680 3740
rect 2570 3680 2680 3705
rect 2820 3795 2930 3820
rect 2820 3760 2825 3795
rect 2925 3760 2930 3795
rect 2820 3740 2930 3760
rect 2820 3705 2825 3740
rect 2925 3705 2930 3740
rect 2820 3680 2930 3705
rect 3070 3795 3180 3820
rect 3070 3760 3075 3795
rect 3175 3760 3180 3795
rect 3070 3740 3180 3760
rect 3070 3705 3075 3740
rect 3175 3705 3180 3740
rect 3070 3680 3180 3705
rect 3320 3795 3430 3820
rect 3320 3760 3325 3795
rect 3425 3760 3430 3795
rect 3320 3740 3430 3760
rect 3320 3705 3325 3740
rect 3425 3705 3430 3740
rect 3320 3680 3430 3705
rect 3570 3795 3680 3820
rect 3570 3760 3575 3795
rect 3675 3760 3680 3795
rect 3570 3740 3680 3760
rect 3570 3705 3575 3740
rect 3675 3705 3680 3740
rect 3570 3680 3680 3705
rect 3820 3795 3930 3820
rect 3820 3760 3825 3795
rect 3925 3760 3930 3795
rect 3820 3740 3930 3760
rect 3820 3705 3825 3740
rect 3925 3705 3930 3740
rect 3820 3680 3930 3705
rect 0 3675 4000 3680
rect 0 3575 10 3675
rect 45 3575 205 3675
rect 240 3575 260 3675
rect 295 3575 455 3675
rect 490 3575 510 3675
rect 545 3575 705 3675
rect 740 3575 760 3675
rect 795 3575 955 3675
rect 990 3575 1010 3675
rect 1045 3575 1205 3675
rect 1240 3575 1260 3675
rect 1295 3575 1455 3675
rect 1490 3575 1510 3675
rect 1545 3575 1705 3675
rect 1740 3575 1760 3675
rect 1795 3575 1955 3675
rect 1990 3575 2010 3675
rect 2045 3575 2205 3675
rect 2240 3575 2260 3675
rect 2295 3575 2455 3675
rect 2490 3575 2510 3675
rect 2545 3575 2705 3675
rect 2740 3575 2760 3675
rect 2795 3575 2955 3675
rect 2990 3575 3010 3675
rect 3045 3575 3205 3675
rect 3240 3575 3260 3675
rect 3295 3575 3455 3675
rect 3490 3575 3510 3675
rect 3545 3575 3705 3675
rect 3740 3575 3760 3675
rect 3795 3575 3955 3675
rect 3990 3575 4000 3675
rect 0 3570 4000 3575
rect 70 3545 180 3570
rect 70 3510 75 3545
rect 175 3510 180 3545
rect 70 3490 180 3510
rect 70 3455 75 3490
rect 175 3455 180 3490
rect 70 3430 180 3455
rect 320 3545 430 3570
rect 320 3510 325 3545
rect 425 3510 430 3545
rect 320 3490 430 3510
rect 320 3455 325 3490
rect 425 3455 430 3490
rect 320 3430 430 3455
rect 570 3545 680 3570
rect 570 3510 575 3545
rect 675 3510 680 3545
rect 570 3490 680 3510
rect 570 3455 575 3490
rect 675 3455 680 3490
rect 570 3430 680 3455
rect 820 3545 930 3570
rect 820 3510 825 3545
rect 925 3510 930 3545
rect 820 3490 930 3510
rect 820 3455 825 3490
rect 925 3455 930 3490
rect 820 3430 930 3455
rect 1070 3545 1180 3570
rect 1070 3510 1075 3545
rect 1175 3510 1180 3545
rect 1070 3490 1180 3510
rect 1070 3455 1075 3490
rect 1175 3455 1180 3490
rect 1070 3430 1180 3455
rect 1320 3545 1430 3570
rect 1320 3510 1325 3545
rect 1425 3510 1430 3545
rect 1320 3490 1430 3510
rect 1320 3455 1325 3490
rect 1425 3455 1430 3490
rect 1320 3430 1430 3455
rect 1570 3545 1680 3570
rect 1570 3510 1575 3545
rect 1675 3510 1680 3545
rect 1570 3490 1680 3510
rect 1570 3455 1575 3490
rect 1675 3455 1680 3490
rect 1570 3430 1680 3455
rect 1820 3545 1930 3570
rect 1820 3510 1825 3545
rect 1925 3510 1930 3545
rect 1820 3490 1930 3510
rect 1820 3455 1825 3490
rect 1925 3455 1930 3490
rect 1820 3430 1930 3455
rect 2070 3545 2180 3570
rect 2070 3510 2075 3545
rect 2175 3510 2180 3545
rect 2070 3490 2180 3510
rect 2070 3455 2075 3490
rect 2175 3455 2180 3490
rect 2070 3430 2180 3455
rect 2320 3545 2430 3570
rect 2320 3510 2325 3545
rect 2425 3510 2430 3545
rect 2320 3490 2430 3510
rect 2320 3455 2325 3490
rect 2425 3455 2430 3490
rect 2320 3430 2430 3455
rect 2570 3545 2680 3570
rect 2570 3510 2575 3545
rect 2675 3510 2680 3545
rect 2570 3490 2680 3510
rect 2570 3455 2575 3490
rect 2675 3455 2680 3490
rect 2570 3430 2680 3455
rect 2820 3545 2930 3570
rect 2820 3510 2825 3545
rect 2925 3510 2930 3545
rect 2820 3490 2930 3510
rect 2820 3455 2825 3490
rect 2925 3455 2930 3490
rect 2820 3430 2930 3455
rect 3070 3545 3180 3570
rect 3070 3510 3075 3545
rect 3175 3510 3180 3545
rect 3070 3490 3180 3510
rect 3070 3455 3075 3490
rect 3175 3455 3180 3490
rect 3070 3430 3180 3455
rect 3320 3545 3430 3570
rect 3320 3510 3325 3545
rect 3425 3510 3430 3545
rect 3320 3490 3430 3510
rect 3320 3455 3325 3490
rect 3425 3455 3430 3490
rect 3320 3430 3430 3455
rect 3570 3545 3680 3570
rect 3570 3510 3575 3545
rect 3675 3510 3680 3545
rect 3570 3490 3680 3510
rect 3570 3455 3575 3490
rect 3675 3455 3680 3490
rect 3570 3430 3680 3455
rect 3820 3545 3930 3570
rect 3820 3510 3825 3545
rect 3925 3510 3930 3545
rect 3820 3490 3930 3510
rect 3820 3455 3825 3490
rect 3925 3455 3930 3490
rect 3820 3430 3930 3455
rect 0 3425 4000 3430
rect 0 3325 10 3425
rect 45 3325 205 3425
rect 240 3325 260 3425
rect 295 3325 455 3425
rect 490 3325 510 3425
rect 545 3325 705 3425
rect 740 3325 760 3425
rect 795 3325 955 3425
rect 990 3325 1010 3425
rect 1045 3325 1205 3425
rect 1240 3325 1260 3425
rect 1295 3325 1455 3425
rect 1490 3325 1510 3425
rect 1545 3325 1705 3425
rect 1740 3325 1760 3425
rect 1795 3325 1955 3425
rect 1990 3325 2010 3425
rect 2045 3325 2205 3425
rect 2240 3325 2260 3425
rect 2295 3325 2455 3425
rect 2490 3325 2510 3425
rect 2545 3325 2705 3425
rect 2740 3325 2760 3425
rect 2795 3325 2955 3425
rect 2990 3325 3010 3425
rect 3045 3325 3205 3425
rect 3240 3325 3260 3425
rect 3295 3325 3455 3425
rect 3490 3325 3510 3425
rect 3545 3325 3705 3425
rect 3740 3325 3760 3425
rect 3795 3325 3955 3425
rect 3990 3325 4000 3425
rect 0 3320 4000 3325
rect 70 3295 180 3320
rect 70 3260 75 3295
rect 175 3260 180 3295
rect 70 3240 180 3260
rect 70 3205 75 3240
rect 175 3205 180 3240
rect 70 3180 180 3205
rect 320 3295 430 3320
rect 320 3260 325 3295
rect 425 3260 430 3295
rect 320 3240 430 3260
rect 320 3205 325 3240
rect 425 3205 430 3240
rect 320 3180 430 3205
rect 570 3295 680 3320
rect 570 3260 575 3295
rect 675 3260 680 3295
rect 570 3240 680 3260
rect 570 3205 575 3240
rect 675 3205 680 3240
rect 570 3180 680 3205
rect 820 3295 930 3320
rect 820 3260 825 3295
rect 925 3260 930 3295
rect 820 3240 930 3260
rect 820 3205 825 3240
rect 925 3205 930 3240
rect 820 3180 930 3205
rect 1070 3295 1180 3320
rect 1070 3260 1075 3295
rect 1175 3260 1180 3295
rect 1070 3240 1180 3260
rect 1070 3205 1075 3240
rect 1175 3205 1180 3240
rect 1070 3180 1180 3205
rect 1320 3295 1430 3320
rect 1320 3260 1325 3295
rect 1425 3260 1430 3295
rect 1320 3240 1430 3260
rect 1320 3205 1325 3240
rect 1425 3205 1430 3240
rect 1320 3180 1430 3205
rect 1570 3295 1680 3320
rect 1570 3260 1575 3295
rect 1675 3260 1680 3295
rect 1570 3240 1680 3260
rect 1570 3205 1575 3240
rect 1675 3205 1680 3240
rect 1570 3180 1680 3205
rect 1820 3295 1930 3320
rect 1820 3260 1825 3295
rect 1925 3260 1930 3295
rect 1820 3240 1930 3260
rect 1820 3205 1825 3240
rect 1925 3205 1930 3240
rect 1820 3180 1930 3205
rect 2070 3295 2180 3320
rect 2070 3260 2075 3295
rect 2175 3260 2180 3295
rect 2070 3240 2180 3260
rect 2070 3205 2075 3240
rect 2175 3205 2180 3240
rect 2070 3180 2180 3205
rect 2320 3295 2430 3320
rect 2320 3260 2325 3295
rect 2425 3260 2430 3295
rect 2320 3240 2430 3260
rect 2320 3205 2325 3240
rect 2425 3205 2430 3240
rect 2320 3180 2430 3205
rect 2570 3295 2680 3320
rect 2570 3260 2575 3295
rect 2675 3260 2680 3295
rect 2570 3240 2680 3260
rect 2570 3205 2575 3240
rect 2675 3205 2680 3240
rect 2570 3180 2680 3205
rect 2820 3295 2930 3320
rect 2820 3260 2825 3295
rect 2925 3260 2930 3295
rect 2820 3240 2930 3260
rect 2820 3205 2825 3240
rect 2925 3205 2930 3240
rect 2820 3180 2930 3205
rect 3070 3295 3180 3320
rect 3070 3260 3075 3295
rect 3175 3260 3180 3295
rect 3070 3240 3180 3260
rect 3070 3205 3075 3240
rect 3175 3205 3180 3240
rect 3070 3180 3180 3205
rect 3320 3295 3430 3320
rect 3320 3260 3325 3295
rect 3425 3260 3430 3295
rect 3320 3240 3430 3260
rect 3320 3205 3325 3240
rect 3425 3205 3430 3240
rect 3320 3180 3430 3205
rect 3570 3295 3680 3320
rect 3570 3260 3575 3295
rect 3675 3260 3680 3295
rect 3570 3240 3680 3260
rect 3570 3205 3575 3240
rect 3675 3205 3680 3240
rect 3570 3180 3680 3205
rect 3820 3295 3930 3320
rect 3820 3260 3825 3295
rect 3925 3260 3930 3295
rect 3820 3240 3930 3260
rect 3820 3205 3825 3240
rect 3925 3205 3930 3240
rect 3820 3180 3930 3205
rect 0 3175 4000 3180
rect 0 3075 10 3175
rect 45 3075 205 3175
rect 240 3075 260 3175
rect 295 3075 455 3175
rect 490 3075 510 3175
rect 545 3075 705 3175
rect 740 3075 760 3175
rect 795 3075 955 3175
rect 990 3075 1010 3175
rect 1045 3075 1205 3175
rect 1240 3075 1260 3175
rect 1295 3075 1455 3175
rect 1490 3075 1510 3175
rect 1545 3075 1705 3175
rect 1740 3075 1760 3175
rect 1795 3075 1955 3175
rect 1990 3075 2010 3175
rect 2045 3075 2205 3175
rect 2240 3075 2260 3175
rect 2295 3075 2455 3175
rect 2490 3075 2510 3175
rect 2545 3075 2705 3175
rect 2740 3075 2760 3175
rect 2795 3075 2955 3175
rect 2990 3075 3010 3175
rect 3045 3075 3205 3175
rect 3240 3075 3260 3175
rect 3295 3075 3455 3175
rect 3490 3075 3510 3175
rect 3545 3075 3705 3175
rect 3740 3075 3760 3175
rect 3795 3075 3955 3175
rect 3990 3075 4000 3175
rect 0 3070 4000 3075
rect 70 3045 180 3070
rect 70 3010 75 3045
rect 175 3010 180 3045
rect 70 2990 180 3010
rect 70 2955 75 2990
rect 175 2955 180 2990
rect 70 2930 180 2955
rect 320 3045 430 3070
rect 320 3010 325 3045
rect 425 3010 430 3045
rect 320 2990 430 3010
rect 320 2955 325 2990
rect 425 2955 430 2990
rect 320 2930 430 2955
rect 570 3045 680 3070
rect 570 3010 575 3045
rect 675 3010 680 3045
rect 570 2990 680 3010
rect 570 2955 575 2990
rect 675 2955 680 2990
rect 570 2930 680 2955
rect 820 3045 930 3070
rect 820 3010 825 3045
rect 925 3010 930 3045
rect 820 2990 930 3010
rect 820 2955 825 2990
rect 925 2955 930 2990
rect 820 2930 930 2955
rect 1070 3045 1180 3070
rect 1070 3010 1075 3045
rect 1175 3010 1180 3045
rect 1070 2990 1180 3010
rect 1070 2955 1075 2990
rect 1175 2955 1180 2990
rect 1070 2930 1180 2955
rect 1320 3045 1430 3070
rect 1320 3010 1325 3045
rect 1425 3010 1430 3045
rect 1320 2990 1430 3010
rect 1320 2955 1325 2990
rect 1425 2955 1430 2990
rect 1320 2930 1430 2955
rect 1570 3045 1680 3070
rect 1570 3010 1575 3045
rect 1675 3010 1680 3045
rect 1570 2990 1680 3010
rect 1570 2955 1575 2990
rect 1675 2955 1680 2990
rect 1570 2930 1680 2955
rect 1820 3045 1930 3070
rect 1820 3010 1825 3045
rect 1925 3010 1930 3045
rect 1820 2990 1930 3010
rect 1820 2955 1825 2990
rect 1925 2955 1930 2990
rect 1820 2930 1930 2955
rect 2070 3045 2180 3070
rect 2070 3010 2075 3045
rect 2175 3010 2180 3045
rect 2070 2990 2180 3010
rect 2070 2955 2075 2990
rect 2175 2955 2180 2990
rect 2070 2930 2180 2955
rect 2320 3045 2430 3070
rect 2320 3010 2325 3045
rect 2425 3010 2430 3045
rect 2320 2990 2430 3010
rect 2320 2955 2325 2990
rect 2425 2955 2430 2990
rect 2320 2930 2430 2955
rect 2570 3045 2680 3070
rect 2570 3010 2575 3045
rect 2675 3010 2680 3045
rect 2570 2990 2680 3010
rect 2570 2955 2575 2990
rect 2675 2955 2680 2990
rect 2570 2930 2680 2955
rect 2820 3045 2930 3070
rect 2820 3010 2825 3045
rect 2925 3010 2930 3045
rect 2820 2990 2930 3010
rect 2820 2955 2825 2990
rect 2925 2955 2930 2990
rect 2820 2930 2930 2955
rect 3070 3045 3180 3070
rect 3070 3010 3075 3045
rect 3175 3010 3180 3045
rect 3070 2990 3180 3010
rect 3070 2955 3075 2990
rect 3175 2955 3180 2990
rect 3070 2930 3180 2955
rect 3320 3045 3430 3070
rect 3320 3010 3325 3045
rect 3425 3010 3430 3045
rect 3320 2990 3430 3010
rect 3320 2955 3325 2990
rect 3425 2955 3430 2990
rect 3320 2930 3430 2955
rect 3570 3045 3680 3070
rect 3570 3010 3575 3045
rect 3675 3010 3680 3045
rect 3570 2990 3680 3010
rect 3570 2955 3575 2990
rect 3675 2955 3680 2990
rect 3570 2930 3680 2955
rect 3820 3045 3930 3070
rect 3820 3010 3825 3045
rect 3925 3010 3930 3045
rect 3820 2990 3930 3010
rect 3820 2955 3825 2990
rect 3925 2955 3930 2990
rect 3820 2930 3930 2955
rect 0 2925 4000 2930
rect 0 2825 10 2925
rect 45 2825 205 2925
rect 240 2825 260 2925
rect 295 2825 455 2925
rect 490 2825 510 2925
rect 545 2825 705 2925
rect 740 2825 760 2925
rect 795 2825 955 2925
rect 990 2825 1010 2925
rect 1045 2825 1205 2925
rect 1240 2825 1260 2925
rect 1295 2825 1455 2925
rect 1490 2825 1510 2925
rect 1545 2825 1705 2925
rect 1740 2825 1760 2925
rect 1795 2825 1955 2925
rect 1990 2825 2010 2925
rect 2045 2825 2205 2925
rect 2240 2825 2260 2925
rect 2295 2825 2455 2925
rect 2490 2825 2510 2925
rect 2545 2825 2705 2925
rect 2740 2825 2760 2925
rect 2795 2825 2955 2925
rect 2990 2825 3010 2925
rect 3045 2825 3205 2925
rect 3240 2825 3260 2925
rect 3295 2825 3455 2925
rect 3490 2825 3510 2925
rect 3545 2825 3705 2925
rect 3740 2825 3760 2925
rect 3795 2825 3955 2925
rect 3990 2825 4000 2925
rect 0 2820 4000 2825
rect 70 2795 180 2820
rect 70 2760 75 2795
rect 175 2760 180 2795
rect 70 2740 180 2760
rect 70 2705 75 2740
rect 175 2705 180 2740
rect 70 2680 180 2705
rect 320 2795 430 2820
rect 320 2760 325 2795
rect 425 2760 430 2795
rect 320 2740 430 2760
rect 320 2705 325 2740
rect 425 2705 430 2740
rect 320 2680 430 2705
rect 570 2795 680 2820
rect 570 2760 575 2795
rect 675 2760 680 2795
rect 570 2740 680 2760
rect 570 2705 575 2740
rect 675 2705 680 2740
rect 570 2680 680 2705
rect 820 2795 930 2820
rect 820 2760 825 2795
rect 925 2760 930 2795
rect 820 2740 930 2760
rect 820 2705 825 2740
rect 925 2705 930 2740
rect 820 2680 930 2705
rect 1070 2795 1180 2820
rect 1070 2760 1075 2795
rect 1175 2760 1180 2795
rect 1070 2740 1180 2760
rect 1070 2705 1075 2740
rect 1175 2705 1180 2740
rect 1070 2680 1180 2705
rect 1320 2795 1430 2820
rect 1320 2760 1325 2795
rect 1425 2760 1430 2795
rect 1320 2740 1430 2760
rect 1320 2705 1325 2740
rect 1425 2705 1430 2740
rect 1320 2680 1430 2705
rect 1570 2795 1680 2820
rect 1570 2760 1575 2795
rect 1675 2760 1680 2795
rect 1570 2740 1680 2760
rect 1570 2705 1575 2740
rect 1675 2705 1680 2740
rect 1570 2680 1680 2705
rect 1820 2795 1930 2820
rect 1820 2760 1825 2795
rect 1925 2760 1930 2795
rect 1820 2740 1930 2760
rect 1820 2705 1825 2740
rect 1925 2705 1930 2740
rect 1820 2680 1930 2705
rect 2070 2795 2180 2820
rect 2070 2760 2075 2795
rect 2175 2760 2180 2795
rect 2070 2740 2180 2760
rect 2070 2705 2075 2740
rect 2175 2705 2180 2740
rect 2070 2680 2180 2705
rect 2320 2795 2430 2820
rect 2320 2760 2325 2795
rect 2425 2760 2430 2795
rect 2320 2740 2430 2760
rect 2320 2705 2325 2740
rect 2425 2705 2430 2740
rect 2320 2680 2430 2705
rect 2570 2795 2680 2820
rect 2570 2760 2575 2795
rect 2675 2760 2680 2795
rect 2570 2740 2680 2760
rect 2570 2705 2575 2740
rect 2675 2705 2680 2740
rect 2570 2680 2680 2705
rect 2820 2795 2930 2820
rect 2820 2760 2825 2795
rect 2925 2760 2930 2795
rect 2820 2740 2930 2760
rect 2820 2705 2825 2740
rect 2925 2705 2930 2740
rect 2820 2680 2930 2705
rect 3070 2795 3180 2820
rect 3070 2760 3075 2795
rect 3175 2760 3180 2795
rect 3070 2740 3180 2760
rect 3070 2705 3075 2740
rect 3175 2705 3180 2740
rect 3070 2680 3180 2705
rect 3320 2795 3430 2820
rect 3320 2760 3325 2795
rect 3425 2760 3430 2795
rect 3320 2740 3430 2760
rect 3320 2705 3325 2740
rect 3425 2705 3430 2740
rect 3320 2680 3430 2705
rect 3570 2795 3680 2820
rect 3570 2760 3575 2795
rect 3675 2760 3680 2795
rect 3570 2740 3680 2760
rect 3570 2705 3575 2740
rect 3675 2705 3680 2740
rect 3570 2680 3680 2705
rect 3820 2795 3930 2820
rect 3820 2760 3825 2795
rect 3925 2760 3930 2795
rect 3820 2740 3930 2760
rect 3820 2705 3825 2740
rect 3925 2705 3930 2740
rect 3820 2680 3930 2705
rect 0 2675 4000 2680
rect 0 2575 10 2675
rect 45 2575 205 2675
rect 240 2575 260 2675
rect 295 2575 455 2675
rect 490 2575 510 2675
rect 545 2575 705 2675
rect 740 2575 760 2675
rect 795 2575 955 2675
rect 990 2575 1010 2675
rect 1045 2575 1205 2675
rect 1240 2575 1260 2675
rect 1295 2575 1455 2675
rect 1490 2575 1510 2675
rect 1545 2575 1705 2675
rect 1740 2575 1760 2675
rect 1795 2575 1955 2675
rect 1990 2575 2010 2675
rect 2045 2575 2205 2675
rect 2240 2575 2260 2675
rect 2295 2575 2455 2675
rect 2490 2575 2510 2675
rect 2545 2575 2705 2675
rect 2740 2575 2760 2675
rect 2795 2575 2955 2675
rect 2990 2575 3010 2675
rect 3045 2575 3205 2675
rect 3240 2575 3260 2675
rect 3295 2575 3455 2675
rect 3490 2575 3510 2675
rect 3545 2575 3705 2675
rect 3740 2575 3760 2675
rect 3795 2575 3955 2675
rect 3990 2575 4000 2675
rect 0 2570 4000 2575
rect 70 2545 180 2570
rect 70 2510 75 2545
rect 175 2510 180 2545
rect 70 2490 180 2510
rect 70 2455 75 2490
rect 175 2455 180 2490
rect 70 2430 180 2455
rect 320 2545 430 2570
rect 320 2510 325 2545
rect 425 2510 430 2545
rect 320 2490 430 2510
rect 320 2455 325 2490
rect 425 2455 430 2490
rect 320 2430 430 2455
rect 570 2545 680 2570
rect 570 2510 575 2545
rect 675 2510 680 2545
rect 570 2490 680 2510
rect 570 2455 575 2490
rect 675 2455 680 2490
rect 570 2430 680 2455
rect 820 2545 930 2570
rect 820 2510 825 2545
rect 925 2510 930 2545
rect 820 2490 930 2510
rect 820 2455 825 2490
rect 925 2455 930 2490
rect 820 2430 930 2455
rect 1070 2545 1180 2570
rect 1070 2510 1075 2545
rect 1175 2510 1180 2545
rect 1070 2490 1180 2510
rect 1070 2455 1075 2490
rect 1175 2455 1180 2490
rect 1070 2430 1180 2455
rect 1320 2545 1430 2570
rect 1320 2510 1325 2545
rect 1425 2510 1430 2545
rect 1320 2490 1430 2510
rect 1320 2455 1325 2490
rect 1425 2455 1430 2490
rect 1320 2430 1430 2455
rect 1570 2545 1680 2570
rect 1570 2510 1575 2545
rect 1675 2510 1680 2545
rect 1570 2490 1680 2510
rect 1570 2455 1575 2490
rect 1675 2455 1680 2490
rect 1570 2430 1680 2455
rect 1820 2545 1930 2570
rect 1820 2510 1825 2545
rect 1925 2510 1930 2545
rect 1820 2490 1930 2510
rect 1820 2455 1825 2490
rect 1925 2455 1930 2490
rect 1820 2430 1930 2455
rect 2070 2545 2180 2570
rect 2070 2510 2075 2545
rect 2175 2510 2180 2545
rect 2070 2490 2180 2510
rect 2070 2455 2075 2490
rect 2175 2455 2180 2490
rect 2070 2430 2180 2455
rect 2320 2545 2430 2570
rect 2320 2510 2325 2545
rect 2425 2510 2430 2545
rect 2320 2490 2430 2510
rect 2320 2455 2325 2490
rect 2425 2455 2430 2490
rect 2320 2430 2430 2455
rect 2570 2545 2680 2570
rect 2570 2510 2575 2545
rect 2675 2510 2680 2545
rect 2570 2490 2680 2510
rect 2570 2455 2575 2490
rect 2675 2455 2680 2490
rect 2570 2430 2680 2455
rect 2820 2545 2930 2570
rect 2820 2510 2825 2545
rect 2925 2510 2930 2545
rect 2820 2490 2930 2510
rect 2820 2455 2825 2490
rect 2925 2455 2930 2490
rect 2820 2430 2930 2455
rect 3070 2545 3180 2570
rect 3070 2510 3075 2545
rect 3175 2510 3180 2545
rect 3070 2490 3180 2510
rect 3070 2455 3075 2490
rect 3175 2455 3180 2490
rect 3070 2430 3180 2455
rect 3320 2545 3430 2570
rect 3320 2510 3325 2545
rect 3425 2510 3430 2545
rect 3320 2490 3430 2510
rect 3320 2455 3325 2490
rect 3425 2455 3430 2490
rect 3320 2430 3430 2455
rect 3570 2545 3680 2570
rect 3570 2510 3575 2545
rect 3675 2510 3680 2545
rect 3570 2490 3680 2510
rect 3570 2455 3575 2490
rect 3675 2455 3680 2490
rect 3570 2430 3680 2455
rect 3820 2545 3930 2570
rect 3820 2510 3825 2545
rect 3925 2510 3930 2545
rect 3820 2490 3930 2510
rect 3820 2455 3825 2490
rect 3925 2455 3930 2490
rect 3820 2430 3930 2455
rect 0 2425 4000 2430
rect 0 2325 10 2425
rect 45 2325 205 2425
rect 240 2325 260 2425
rect 295 2325 455 2425
rect 490 2325 510 2425
rect 545 2325 705 2425
rect 740 2325 760 2425
rect 795 2325 955 2425
rect 990 2325 1010 2425
rect 1045 2325 1205 2425
rect 1240 2325 1260 2425
rect 1295 2325 1455 2425
rect 1490 2325 1510 2425
rect 1545 2325 1705 2425
rect 1740 2325 1760 2425
rect 1795 2325 1955 2425
rect 1990 2325 2010 2425
rect 2045 2325 2205 2425
rect 2240 2325 2260 2425
rect 2295 2325 2455 2425
rect 2490 2325 2510 2425
rect 2545 2325 2705 2425
rect 2740 2325 2760 2425
rect 2795 2325 2955 2425
rect 2990 2325 3010 2425
rect 3045 2325 3205 2425
rect 3240 2325 3260 2425
rect 3295 2325 3455 2425
rect 3490 2325 3510 2425
rect 3545 2325 3705 2425
rect 3740 2325 3760 2425
rect 3795 2325 3955 2425
rect 3990 2325 4000 2425
rect 0 2320 4000 2325
rect 70 2295 180 2320
rect 70 2260 75 2295
rect 175 2260 180 2295
rect 70 2240 180 2260
rect 70 2205 75 2240
rect 175 2205 180 2240
rect 70 2180 180 2205
rect 320 2295 430 2320
rect 320 2260 325 2295
rect 425 2260 430 2295
rect 320 2240 430 2260
rect 320 2205 325 2240
rect 425 2205 430 2240
rect 320 2180 430 2205
rect 570 2295 680 2320
rect 570 2260 575 2295
rect 675 2260 680 2295
rect 570 2240 680 2260
rect 570 2205 575 2240
rect 675 2205 680 2240
rect 570 2180 680 2205
rect 820 2295 930 2320
rect 820 2260 825 2295
rect 925 2260 930 2295
rect 820 2240 930 2260
rect 820 2205 825 2240
rect 925 2205 930 2240
rect 820 2180 930 2205
rect 1070 2295 1180 2320
rect 1070 2260 1075 2295
rect 1175 2260 1180 2295
rect 1070 2240 1180 2260
rect 1070 2205 1075 2240
rect 1175 2205 1180 2240
rect 1070 2180 1180 2205
rect 1320 2295 1430 2320
rect 1320 2260 1325 2295
rect 1425 2260 1430 2295
rect 1320 2240 1430 2260
rect 1320 2205 1325 2240
rect 1425 2205 1430 2240
rect 1320 2180 1430 2205
rect 1570 2295 1680 2320
rect 1570 2260 1575 2295
rect 1675 2260 1680 2295
rect 1570 2240 1680 2260
rect 1570 2205 1575 2240
rect 1675 2205 1680 2240
rect 1570 2180 1680 2205
rect 1820 2295 1930 2320
rect 1820 2260 1825 2295
rect 1925 2260 1930 2295
rect 1820 2240 1930 2260
rect 1820 2205 1825 2240
rect 1925 2205 1930 2240
rect 1820 2180 1930 2205
rect 2070 2295 2180 2320
rect 2070 2260 2075 2295
rect 2175 2260 2180 2295
rect 2070 2240 2180 2260
rect 2070 2205 2075 2240
rect 2175 2205 2180 2240
rect 2070 2180 2180 2205
rect 2320 2295 2430 2320
rect 2320 2260 2325 2295
rect 2425 2260 2430 2295
rect 2320 2240 2430 2260
rect 2320 2205 2325 2240
rect 2425 2205 2430 2240
rect 2320 2180 2430 2205
rect 2570 2295 2680 2320
rect 2570 2260 2575 2295
rect 2675 2260 2680 2295
rect 2570 2240 2680 2260
rect 2570 2205 2575 2240
rect 2675 2205 2680 2240
rect 2570 2180 2680 2205
rect 2820 2295 2930 2320
rect 2820 2260 2825 2295
rect 2925 2260 2930 2295
rect 2820 2240 2930 2260
rect 2820 2205 2825 2240
rect 2925 2205 2930 2240
rect 2820 2180 2930 2205
rect 3070 2295 3180 2320
rect 3070 2260 3075 2295
rect 3175 2260 3180 2295
rect 3070 2240 3180 2260
rect 3070 2205 3075 2240
rect 3175 2205 3180 2240
rect 3070 2180 3180 2205
rect 3320 2295 3430 2320
rect 3320 2260 3325 2295
rect 3425 2260 3430 2295
rect 3320 2240 3430 2260
rect 3320 2205 3325 2240
rect 3425 2205 3430 2240
rect 3320 2180 3430 2205
rect 3570 2295 3680 2320
rect 3570 2260 3575 2295
rect 3675 2260 3680 2295
rect 3570 2240 3680 2260
rect 3570 2205 3575 2240
rect 3675 2205 3680 2240
rect 3570 2180 3680 2205
rect 3820 2295 3930 2320
rect 3820 2260 3825 2295
rect 3925 2260 3930 2295
rect 3820 2240 3930 2260
rect 3820 2205 3825 2240
rect 3925 2205 3930 2240
rect 3820 2180 3930 2205
rect 0 2175 4000 2180
rect 0 2075 10 2175
rect 45 2075 205 2175
rect 240 2075 260 2175
rect 295 2075 455 2175
rect 490 2075 510 2175
rect 545 2075 705 2175
rect 740 2075 760 2175
rect 795 2075 955 2175
rect 990 2075 1010 2175
rect 1045 2075 1205 2175
rect 1240 2075 1260 2175
rect 1295 2075 1455 2175
rect 1490 2075 1510 2175
rect 1545 2075 1705 2175
rect 1740 2075 1760 2175
rect 1795 2075 1955 2175
rect 1990 2075 2010 2175
rect 2045 2075 2205 2175
rect 2240 2075 2260 2175
rect 2295 2075 2455 2175
rect 2490 2075 2510 2175
rect 2545 2075 2705 2175
rect 2740 2075 2760 2175
rect 2795 2075 2955 2175
rect 2990 2075 3010 2175
rect 3045 2075 3205 2175
rect 3240 2075 3260 2175
rect 3295 2075 3455 2175
rect 3490 2075 3510 2175
rect 3545 2075 3705 2175
rect 3740 2075 3760 2175
rect 3795 2075 3955 2175
rect 3990 2075 4000 2175
rect 0 2070 4000 2075
rect 70 2045 180 2070
rect 70 2010 75 2045
rect 175 2010 180 2045
rect 70 1990 180 2010
rect 70 1955 75 1990
rect 175 1955 180 1990
rect 70 1930 180 1955
rect 320 2045 430 2070
rect 320 2010 325 2045
rect 425 2010 430 2045
rect 320 1990 430 2010
rect 320 1955 325 1990
rect 425 1955 430 1990
rect 320 1930 430 1955
rect 570 2045 680 2070
rect 570 2010 575 2045
rect 675 2010 680 2045
rect 570 1990 680 2010
rect 570 1955 575 1990
rect 675 1955 680 1990
rect 570 1930 680 1955
rect 820 2045 930 2070
rect 820 2010 825 2045
rect 925 2010 930 2045
rect 820 1990 930 2010
rect 820 1955 825 1990
rect 925 1955 930 1990
rect 820 1930 930 1955
rect 1070 2045 1180 2070
rect 1070 2010 1075 2045
rect 1175 2010 1180 2045
rect 1070 1990 1180 2010
rect 1070 1955 1075 1990
rect 1175 1955 1180 1990
rect 1070 1930 1180 1955
rect 1320 2045 1430 2070
rect 1320 2010 1325 2045
rect 1425 2010 1430 2045
rect 1320 1990 1430 2010
rect 1320 1955 1325 1990
rect 1425 1955 1430 1990
rect 1320 1930 1430 1955
rect 1570 2045 1680 2070
rect 1570 2010 1575 2045
rect 1675 2010 1680 2045
rect 1570 1990 1680 2010
rect 1570 1955 1575 1990
rect 1675 1955 1680 1990
rect 1570 1930 1680 1955
rect 1820 2045 1930 2070
rect 1820 2010 1825 2045
rect 1925 2010 1930 2045
rect 1820 1990 1930 2010
rect 1820 1955 1825 1990
rect 1925 1955 1930 1990
rect 1820 1930 1930 1955
rect 2070 2045 2180 2070
rect 2070 2010 2075 2045
rect 2175 2010 2180 2045
rect 2070 1990 2180 2010
rect 2070 1955 2075 1990
rect 2175 1955 2180 1990
rect 2070 1930 2180 1955
rect 2320 2045 2430 2070
rect 2320 2010 2325 2045
rect 2425 2010 2430 2045
rect 2320 1990 2430 2010
rect 2320 1955 2325 1990
rect 2425 1955 2430 1990
rect 2320 1930 2430 1955
rect 2570 2045 2680 2070
rect 2570 2010 2575 2045
rect 2675 2010 2680 2045
rect 2570 1990 2680 2010
rect 2570 1955 2575 1990
rect 2675 1955 2680 1990
rect 2570 1930 2680 1955
rect 2820 2045 2930 2070
rect 2820 2010 2825 2045
rect 2925 2010 2930 2045
rect 2820 1990 2930 2010
rect 2820 1955 2825 1990
rect 2925 1955 2930 1990
rect 2820 1930 2930 1955
rect 3070 2045 3180 2070
rect 3070 2010 3075 2045
rect 3175 2010 3180 2045
rect 3070 1990 3180 2010
rect 3070 1955 3075 1990
rect 3175 1955 3180 1990
rect 3070 1930 3180 1955
rect 3320 2045 3430 2070
rect 3320 2010 3325 2045
rect 3425 2010 3430 2045
rect 3320 1990 3430 2010
rect 3320 1955 3325 1990
rect 3425 1955 3430 1990
rect 3320 1930 3430 1955
rect 3570 2045 3680 2070
rect 3570 2010 3575 2045
rect 3675 2010 3680 2045
rect 3570 1990 3680 2010
rect 3570 1955 3575 1990
rect 3675 1955 3680 1990
rect 3570 1930 3680 1955
rect 3820 2045 3930 2070
rect 3820 2010 3825 2045
rect 3925 2010 3930 2045
rect 3820 1990 3930 2010
rect 3820 1955 3825 1990
rect 3925 1955 3930 1990
rect 3820 1930 3930 1955
rect 0 1925 4000 1930
rect 0 1825 10 1925
rect 45 1825 205 1925
rect 240 1825 260 1925
rect 295 1825 455 1925
rect 490 1825 510 1925
rect 545 1825 705 1925
rect 740 1825 760 1925
rect 795 1825 955 1925
rect 990 1825 1010 1925
rect 1045 1825 1205 1925
rect 1240 1825 1260 1925
rect 1295 1825 1455 1925
rect 1490 1825 1510 1925
rect 1545 1825 1705 1925
rect 1740 1825 1760 1925
rect 1795 1825 1955 1925
rect 1990 1825 2010 1925
rect 2045 1825 2205 1925
rect 2240 1825 2260 1925
rect 2295 1825 2455 1925
rect 2490 1825 2510 1925
rect 2545 1825 2705 1925
rect 2740 1825 2760 1925
rect 2795 1825 2955 1925
rect 2990 1825 3010 1925
rect 3045 1825 3205 1925
rect 3240 1825 3260 1925
rect 3295 1825 3455 1925
rect 3490 1825 3510 1925
rect 3545 1825 3705 1925
rect 3740 1825 3760 1925
rect 3795 1825 3955 1925
rect 3990 1825 4000 1925
rect 0 1820 4000 1825
rect 70 1795 180 1820
rect 70 1760 75 1795
rect 175 1760 180 1795
rect 70 1740 180 1760
rect 70 1705 75 1740
rect 175 1705 180 1740
rect 70 1680 180 1705
rect 320 1795 430 1820
rect 320 1760 325 1795
rect 425 1760 430 1795
rect 320 1740 430 1760
rect 320 1705 325 1740
rect 425 1705 430 1740
rect 320 1680 430 1705
rect 570 1795 680 1820
rect 570 1760 575 1795
rect 675 1760 680 1795
rect 570 1740 680 1760
rect 570 1705 575 1740
rect 675 1705 680 1740
rect 570 1680 680 1705
rect 820 1795 930 1820
rect 820 1760 825 1795
rect 925 1760 930 1795
rect 820 1740 930 1760
rect 820 1705 825 1740
rect 925 1705 930 1740
rect 820 1680 930 1705
rect 1070 1795 1180 1820
rect 1070 1760 1075 1795
rect 1175 1760 1180 1795
rect 1070 1740 1180 1760
rect 1070 1705 1075 1740
rect 1175 1705 1180 1740
rect 1070 1680 1180 1705
rect 1320 1795 1430 1820
rect 1320 1760 1325 1795
rect 1425 1760 1430 1795
rect 1320 1740 1430 1760
rect 1320 1705 1325 1740
rect 1425 1705 1430 1740
rect 1320 1680 1430 1705
rect 1570 1795 1680 1820
rect 1570 1760 1575 1795
rect 1675 1760 1680 1795
rect 1570 1740 1680 1760
rect 1570 1705 1575 1740
rect 1675 1705 1680 1740
rect 1570 1680 1680 1705
rect 1820 1795 1930 1820
rect 1820 1760 1825 1795
rect 1925 1760 1930 1795
rect 1820 1740 1930 1760
rect 1820 1705 1825 1740
rect 1925 1705 1930 1740
rect 1820 1680 1930 1705
rect 2070 1795 2180 1820
rect 2070 1760 2075 1795
rect 2175 1760 2180 1795
rect 2070 1740 2180 1760
rect 2070 1705 2075 1740
rect 2175 1705 2180 1740
rect 2070 1680 2180 1705
rect 2320 1795 2430 1820
rect 2320 1760 2325 1795
rect 2425 1760 2430 1795
rect 2320 1740 2430 1760
rect 2320 1705 2325 1740
rect 2425 1705 2430 1740
rect 2320 1680 2430 1705
rect 2570 1795 2680 1820
rect 2570 1760 2575 1795
rect 2675 1760 2680 1795
rect 2570 1740 2680 1760
rect 2570 1705 2575 1740
rect 2675 1705 2680 1740
rect 2570 1680 2680 1705
rect 2820 1795 2930 1820
rect 2820 1760 2825 1795
rect 2925 1760 2930 1795
rect 2820 1740 2930 1760
rect 2820 1705 2825 1740
rect 2925 1705 2930 1740
rect 2820 1680 2930 1705
rect 3070 1795 3180 1820
rect 3070 1760 3075 1795
rect 3175 1760 3180 1795
rect 3070 1740 3180 1760
rect 3070 1705 3075 1740
rect 3175 1705 3180 1740
rect 3070 1680 3180 1705
rect 3320 1795 3430 1820
rect 3320 1760 3325 1795
rect 3425 1760 3430 1795
rect 3320 1740 3430 1760
rect 3320 1705 3325 1740
rect 3425 1705 3430 1740
rect 3320 1680 3430 1705
rect 3570 1795 3680 1820
rect 3570 1760 3575 1795
rect 3675 1760 3680 1795
rect 3570 1740 3680 1760
rect 3570 1705 3575 1740
rect 3675 1705 3680 1740
rect 3570 1680 3680 1705
rect 3820 1795 3930 1820
rect 3820 1760 3825 1795
rect 3925 1760 3930 1795
rect 3820 1740 3930 1760
rect 3820 1705 3825 1740
rect 3925 1705 3930 1740
rect 3820 1680 3930 1705
rect 0 1675 4000 1680
rect 0 1575 10 1675
rect 45 1575 205 1675
rect 240 1575 260 1675
rect 295 1575 455 1675
rect 490 1575 510 1675
rect 545 1575 705 1675
rect 740 1575 760 1675
rect 795 1575 955 1675
rect 990 1575 1010 1675
rect 1045 1575 1205 1675
rect 1240 1575 1260 1675
rect 1295 1575 1455 1675
rect 1490 1575 1510 1675
rect 1545 1575 1705 1675
rect 1740 1575 1760 1675
rect 1795 1575 1955 1675
rect 1990 1575 2010 1675
rect 2045 1575 2205 1675
rect 2240 1575 2260 1675
rect 2295 1575 2455 1675
rect 2490 1575 2510 1675
rect 2545 1575 2705 1675
rect 2740 1575 2760 1675
rect 2795 1575 2955 1675
rect 2990 1575 3010 1675
rect 3045 1575 3205 1675
rect 3240 1575 3260 1675
rect 3295 1575 3455 1675
rect 3490 1575 3510 1675
rect 3545 1575 3705 1675
rect 3740 1575 3760 1675
rect 3795 1575 3955 1675
rect 3990 1575 4000 1675
rect 0 1570 4000 1575
rect 70 1545 180 1570
rect 70 1510 75 1545
rect 175 1510 180 1545
rect 70 1490 180 1510
rect 70 1455 75 1490
rect 175 1455 180 1490
rect 70 1430 180 1455
rect 320 1545 430 1570
rect 320 1510 325 1545
rect 425 1510 430 1545
rect 320 1490 430 1510
rect 320 1455 325 1490
rect 425 1455 430 1490
rect 320 1430 430 1455
rect 570 1545 680 1570
rect 570 1510 575 1545
rect 675 1510 680 1545
rect 570 1490 680 1510
rect 570 1455 575 1490
rect 675 1455 680 1490
rect 570 1430 680 1455
rect 820 1545 930 1570
rect 820 1510 825 1545
rect 925 1510 930 1545
rect 820 1490 930 1510
rect 820 1455 825 1490
rect 925 1455 930 1490
rect 820 1430 930 1455
rect 1070 1545 1180 1570
rect 1070 1510 1075 1545
rect 1175 1510 1180 1545
rect 1070 1490 1180 1510
rect 1070 1455 1075 1490
rect 1175 1455 1180 1490
rect 1070 1430 1180 1455
rect 1320 1545 1430 1570
rect 1320 1510 1325 1545
rect 1425 1510 1430 1545
rect 1320 1490 1430 1510
rect 1320 1455 1325 1490
rect 1425 1455 1430 1490
rect 1320 1430 1430 1455
rect 1570 1545 1680 1570
rect 1570 1510 1575 1545
rect 1675 1510 1680 1545
rect 1570 1490 1680 1510
rect 1570 1455 1575 1490
rect 1675 1455 1680 1490
rect 1570 1430 1680 1455
rect 1820 1545 1930 1570
rect 1820 1510 1825 1545
rect 1925 1510 1930 1545
rect 1820 1490 1930 1510
rect 1820 1455 1825 1490
rect 1925 1455 1930 1490
rect 1820 1430 1930 1455
rect 2070 1545 2180 1570
rect 2070 1510 2075 1545
rect 2175 1510 2180 1545
rect 2070 1490 2180 1510
rect 2070 1455 2075 1490
rect 2175 1455 2180 1490
rect 2070 1430 2180 1455
rect 2320 1545 2430 1570
rect 2320 1510 2325 1545
rect 2425 1510 2430 1545
rect 2320 1490 2430 1510
rect 2320 1455 2325 1490
rect 2425 1455 2430 1490
rect 2320 1430 2430 1455
rect 2570 1545 2680 1570
rect 2570 1510 2575 1545
rect 2675 1510 2680 1545
rect 2570 1490 2680 1510
rect 2570 1455 2575 1490
rect 2675 1455 2680 1490
rect 2570 1430 2680 1455
rect 2820 1545 2930 1570
rect 2820 1510 2825 1545
rect 2925 1510 2930 1545
rect 2820 1490 2930 1510
rect 2820 1455 2825 1490
rect 2925 1455 2930 1490
rect 2820 1430 2930 1455
rect 3070 1545 3180 1570
rect 3070 1510 3075 1545
rect 3175 1510 3180 1545
rect 3070 1490 3180 1510
rect 3070 1455 3075 1490
rect 3175 1455 3180 1490
rect 3070 1430 3180 1455
rect 3320 1545 3430 1570
rect 3320 1510 3325 1545
rect 3425 1510 3430 1545
rect 3320 1490 3430 1510
rect 3320 1455 3325 1490
rect 3425 1455 3430 1490
rect 3320 1430 3430 1455
rect 3570 1545 3680 1570
rect 3570 1510 3575 1545
rect 3675 1510 3680 1545
rect 3570 1490 3680 1510
rect 3570 1455 3575 1490
rect 3675 1455 3680 1490
rect 3570 1430 3680 1455
rect 3820 1545 3930 1570
rect 3820 1510 3825 1545
rect 3925 1510 3930 1545
rect 3820 1490 3930 1510
rect 3820 1455 3825 1490
rect 3925 1455 3930 1490
rect 3820 1430 3930 1455
rect 0 1425 4000 1430
rect 0 1325 10 1425
rect 45 1325 205 1425
rect 240 1325 260 1425
rect 295 1325 455 1425
rect 490 1325 510 1425
rect 545 1325 705 1425
rect 740 1325 760 1425
rect 795 1325 955 1425
rect 990 1325 1010 1425
rect 1045 1325 1205 1425
rect 1240 1325 1260 1425
rect 1295 1325 1455 1425
rect 1490 1325 1510 1425
rect 1545 1325 1705 1425
rect 1740 1325 1760 1425
rect 1795 1325 1955 1425
rect 1990 1325 2010 1425
rect 2045 1325 2205 1425
rect 2240 1325 2260 1425
rect 2295 1325 2455 1425
rect 2490 1325 2510 1425
rect 2545 1325 2705 1425
rect 2740 1325 2760 1425
rect 2795 1325 2955 1425
rect 2990 1325 3010 1425
rect 3045 1325 3205 1425
rect 3240 1325 3260 1425
rect 3295 1325 3455 1425
rect 3490 1325 3510 1425
rect 3545 1325 3705 1425
rect 3740 1325 3760 1425
rect 3795 1325 3955 1425
rect 3990 1325 4000 1425
rect 0 1320 4000 1325
rect 70 1295 180 1320
rect 70 1260 75 1295
rect 175 1260 180 1295
rect 70 1240 180 1260
rect 70 1205 75 1240
rect 175 1205 180 1240
rect 70 1180 180 1205
rect 320 1295 430 1320
rect 320 1260 325 1295
rect 425 1260 430 1295
rect 320 1240 430 1260
rect 320 1205 325 1240
rect 425 1205 430 1240
rect 320 1180 430 1205
rect 570 1295 680 1320
rect 570 1260 575 1295
rect 675 1260 680 1295
rect 570 1240 680 1260
rect 570 1205 575 1240
rect 675 1205 680 1240
rect 570 1180 680 1205
rect 820 1295 930 1320
rect 820 1260 825 1295
rect 925 1260 930 1295
rect 820 1240 930 1260
rect 820 1205 825 1240
rect 925 1205 930 1240
rect 820 1180 930 1205
rect 1070 1295 1180 1320
rect 1070 1260 1075 1295
rect 1175 1260 1180 1295
rect 1070 1240 1180 1260
rect 1070 1205 1075 1240
rect 1175 1205 1180 1240
rect 1070 1180 1180 1205
rect 1320 1295 1430 1320
rect 1320 1260 1325 1295
rect 1425 1260 1430 1295
rect 1320 1240 1430 1260
rect 1320 1205 1325 1240
rect 1425 1205 1430 1240
rect 1320 1180 1430 1205
rect 1570 1295 1680 1320
rect 1570 1260 1575 1295
rect 1675 1260 1680 1295
rect 1570 1240 1680 1260
rect 1570 1205 1575 1240
rect 1675 1205 1680 1240
rect 1570 1180 1680 1205
rect 1820 1295 1930 1320
rect 1820 1260 1825 1295
rect 1925 1260 1930 1295
rect 1820 1240 1930 1260
rect 1820 1205 1825 1240
rect 1925 1205 1930 1240
rect 1820 1180 1930 1205
rect 2070 1295 2180 1320
rect 2070 1260 2075 1295
rect 2175 1260 2180 1295
rect 2070 1240 2180 1260
rect 2070 1205 2075 1240
rect 2175 1205 2180 1240
rect 2070 1180 2180 1205
rect 2320 1295 2430 1320
rect 2320 1260 2325 1295
rect 2425 1260 2430 1295
rect 2320 1240 2430 1260
rect 2320 1205 2325 1240
rect 2425 1205 2430 1240
rect 2320 1180 2430 1205
rect 2570 1295 2680 1320
rect 2570 1260 2575 1295
rect 2675 1260 2680 1295
rect 2570 1240 2680 1260
rect 2570 1205 2575 1240
rect 2675 1205 2680 1240
rect 2570 1180 2680 1205
rect 2820 1295 2930 1320
rect 2820 1260 2825 1295
rect 2925 1260 2930 1295
rect 2820 1240 2930 1260
rect 2820 1205 2825 1240
rect 2925 1205 2930 1240
rect 2820 1180 2930 1205
rect 3070 1295 3180 1320
rect 3070 1260 3075 1295
rect 3175 1260 3180 1295
rect 3070 1240 3180 1260
rect 3070 1205 3075 1240
rect 3175 1205 3180 1240
rect 3070 1180 3180 1205
rect 3320 1295 3430 1320
rect 3320 1260 3325 1295
rect 3425 1260 3430 1295
rect 3320 1240 3430 1260
rect 3320 1205 3325 1240
rect 3425 1205 3430 1240
rect 3320 1180 3430 1205
rect 3570 1295 3680 1320
rect 3570 1260 3575 1295
rect 3675 1260 3680 1295
rect 3570 1240 3680 1260
rect 3570 1205 3575 1240
rect 3675 1205 3680 1240
rect 3570 1180 3680 1205
rect 3820 1295 3930 1320
rect 3820 1260 3825 1295
rect 3925 1260 3930 1295
rect 3820 1240 3930 1260
rect 3820 1205 3825 1240
rect 3925 1205 3930 1240
rect 3820 1180 3930 1205
rect 0 1175 4000 1180
rect 0 1075 10 1175
rect 45 1075 205 1175
rect 240 1075 260 1175
rect 295 1075 455 1175
rect 490 1075 510 1175
rect 545 1075 705 1175
rect 740 1075 760 1175
rect 795 1075 955 1175
rect 990 1075 1010 1175
rect 1045 1075 1205 1175
rect 1240 1075 1260 1175
rect 1295 1075 1455 1175
rect 1490 1075 1510 1175
rect 1545 1075 1705 1175
rect 1740 1075 1760 1175
rect 1795 1075 1955 1175
rect 1990 1075 2010 1175
rect 2045 1075 2205 1175
rect 2240 1075 2260 1175
rect 2295 1075 2455 1175
rect 2490 1075 2510 1175
rect 2545 1075 2705 1175
rect 2740 1075 2760 1175
rect 2795 1075 2955 1175
rect 2990 1075 3010 1175
rect 3045 1075 3205 1175
rect 3240 1075 3260 1175
rect 3295 1075 3455 1175
rect 3490 1075 3510 1175
rect 3545 1075 3705 1175
rect 3740 1075 3760 1175
rect 3795 1075 3955 1175
rect 3990 1075 4000 1175
rect 0 1070 4000 1075
rect 70 1045 180 1070
rect 70 1010 75 1045
rect 175 1010 180 1045
rect 70 990 180 1010
rect 70 955 75 990
rect 175 955 180 990
rect 70 930 180 955
rect 320 1045 430 1070
rect 320 1010 325 1045
rect 425 1010 430 1045
rect 320 990 430 1010
rect 320 955 325 990
rect 425 955 430 990
rect 320 930 430 955
rect 570 1045 680 1070
rect 570 1010 575 1045
rect 675 1010 680 1045
rect 570 990 680 1010
rect 570 955 575 990
rect 675 955 680 990
rect 570 930 680 955
rect 820 1045 930 1070
rect 820 1010 825 1045
rect 925 1010 930 1045
rect 820 990 930 1010
rect 820 955 825 990
rect 925 955 930 990
rect 820 930 930 955
rect 1070 1045 1180 1070
rect 1070 1010 1075 1045
rect 1175 1010 1180 1045
rect 1070 990 1180 1010
rect 1070 955 1075 990
rect 1175 955 1180 990
rect 1070 930 1180 955
rect 1320 1045 1430 1070
rect 1320 1010 1325 1045
rect 1425 1010 1430 1045
rect 1320 990 1430 1010
rect 1320 955 1325 990
rect 1425 955 1430 990
rect 1320 930 1430 955
rect 1570 1045 1680 1070
rect 1570 1010 1575 1045
rect 1675 1010 1680 1045
rect 1570 990 1680 1010
rect 1570 955 1575 990
rect 1675 955 1680 990
rect 1570 930 1680 955
rect 1820 1045 1930 1070
rect 1820 1010 1825 1045
rect 1925 1010 1930 1045
rect 1820 990 1930 1010
rect 1820 955 1825 990
rect 1925 955 1930 990
rect 1820 930 1930 955
rect 2070 1045 2180 1070
rect 2070 1010 2075 1045
rect 2175 1010 2180 1045
rect 2070 990 2180 1010
rect 2070 955 2075 990
rect 2175 955 2180 990
rect 2070 930 2180 955
rect 2320 1045 2430 1070
rect 2320 1010 2325 1045
rect 2425 1010 2430 1045
rect 2320 990 2430 1010
rect 2320 955 2325 990
rect 2425 955 2430 990
rect 2320 930 2430 955
rect 2570 1045 2680 1070
rect 2570 1010 2575 1045
rect 2675 1010 2680 1045
rect 2570 990 2680 1010
rect 2570 955 2575 990
rect 2675 955 2680 990
rect 2570 930 2680 955
rect 2820 1045 2930 1070
rect 2820 1010 2825 1045
rect 2925 1010 2930 1045
rect 2820 990 2930 1010
rect 2820 955 2825 990
rect 2925 955 2930 990
rect 2820 930 2930 955
rect 3070 1045 3180 1070
rect 3070 1010 3075 1045
rect 3175 1010 3180 1045
rect 3070 990 3180 1010
rect 3070 955 3075 990
rect 3175 955 3180 990
rect 3070 930 3180 955
rect 3320 1045 3430 1070
rect 3320 1010 3325 1045
rect 3425 1010 3430 1045
rect 3320 990 3430 1010
rect 3320 955 3325 990
rect 3425 955 3430 990
rect 3320 930 3430 955
rect 3570 1045 3680 1070
rect 3570 1010 3575 1045
rect 3675 1010 3680 1045
rect 3570 990 3680 1010
rect 3570 955 3575 990
rect 3675 955 3680 990
rect 3570 930 3680 955
rect 3820 1045 3930 1070
rect 3820 1010 3825 1045
rect 3925 1010 3930 1045
rect 3820 990 3930 1010
rect 3820 955 3825 990
rect 3925 955 3930 990
rect 3820 930 3930 955
rect 0 925 4000 930
rect 0 825 10 925
rect 45 825 205 925
rect 240 825 260 925
rect 295 825 455 925
rect 490 825 510 925
rect 545 825 705 925
rect 740 825 760 925
rect 795 825 955 925
rect 990 825 1010 925
rect 1045 825 1205 925
rect 1240 825 1260 925
rect 1295 825 1455 925
rect 1490 825 1510 925
rect 1545 825 1705 925
rect 1740 825 1760 925
rect 1795 825 1955 925
rect 1990 825 2010 925
rect 2045 825 2205 925
rect 2240 825 2260 925
rect 2295 825 2455 925
rect 2490 825 2510 925
rect 2545 825 2705 925
rect 2740 825 2760 925
rect 2795 825 2955 925
rect 2990 825 3010 925
rect 3045 825 3205 925
rect 3240 825 3260 925
rect 3295 825 3455 925
rect 3490 825 3510 925
rect 3545 825 3705 925
rect 3740 825 3760 925
rect 3795 825 3955 925
rect 3990 825 4000 925
rect 0 820 4000 825
rect 70 795 180 820
rect 70 760 75 795
rect 175 760 180 795
rect 70 740 180 760
rect 70 705 75 740
rect 175 705 180 740
rect 70 680 180 705
rect 320 795 430 820
rect 320 760 325 795
rect 425 760 430 795
rect 320 740 430 760
rect 320 705 325 740
rect 425 705 430 740
rect 320 680 430 705
rect 570 795 680 820
rect 570 760 575 795
rect 675 760 680 795
rect 570 740 680 760
rect 570 705 575 740
rect 675 705 680 740
rect 570 680 680 705
rect 820 795 930 820
rect 820 760 825 795
rect 925 760 930 795
rect 820 740 930 760
rect 820 705 825 740
rect 925 705 930 740
rect 820 680 930 705
rect 1070 795 1180 820
rect 1070 760 1075 795
rect 1175 760 1180 795
rect 1070 740 1180 760
rect 1070 705 1075 740
rect 1175 705 1180 740
rect 1070 680 1180 705
rect 1320 795 1430 820
rect 1320 760 1325 795
rect 1425 760 1430 795
rect 1320 740 1430 760
rect 1320 705 1325 740
rect 1425 705 1430 740
rect 1320 680 1430 705
rect 1570 795 1680 820
rect 1570 760 1575 795
rect 1675 760 1680 795
rect 1570 740 1680 760
rect 1570 705 1575 740
rect 1675 705 1680 740
rect 1570 680 1680 705
rect 1820 795 1930 820
rect 1820 760 1825 795
rect 1925 760 1930 795
rect 1820 740 1930 760
rect 1820 705 1825 740
rect 1925 705 1930 740
rect 1820 680 1930 705
rect 2070 795 2180 820
rect 2070 760 2075 795
rect 2175 760 2180 795
rect 2070 740 2180 760
rect 2070 705 2075 740
rect 2175 705 2180 740
rect 2070 680 2180 705
rect 2320 795 2430 820
rect 2320 760 2325 795
rect 2425 760 2430 795
rect 2320 740 2430 760
rect 2320 705 2325 740
rect 2425 705 2430 740
rect 2320 680 2430 705
rect 2570 795 2680 820
rect 2570 760 2575 795
rect 2675 760 2680 795
rect 2570 740 2680 760
rect 2570 705 2575 740
rect 2675 705 2680 740
rect 2570 680 2680 705
rect 2820 795 2930 820
rect 2820 760 2825 795
rect 2925 760 2930 795
rect 2820 740 2930 760
rect 2820 705 2825 740
rect 2925 705 2930 740
rect 2820 680 2930 705
rect 3070 795 3180 820
rect 3070 760 3075 795
rect 3175 760 3180 795
rect 3070 740 3180 760
rect 3070 705 3075 740
rect 3175 705 3180 740
rect 3070 680 3180 705
rect 3320 795 3430 820
rect 3320 760 3325 795
rect 3425 760 3430 795
rect 3320 740 3430 760
rect 3320 705 3325 740
rect 3425 705 3430 740
rect 3320 680 3430 705
rect 3570 795 3680 820
rect 3570 760 3575 795
rect 3675 760 3680 795
rect 3570 740 3680 760
rect 3570 705 3575 740
rect 3675 705 3680 740
rect 3570 680 3680 705
rect 3820 795 3930 820
rect 3820 760 3825 795
rect 3925 760 3930 795
rect 3820 740 3930 760
rect 3820 705 3825 740
rect 3925 705 3930 740
rect 3820 680 3930 705
rect 0 675 4000 680
rect 0 575 10 675
rect 45 575 205 675
rect 240 575 260 675
rect 295 575 455 675
rect 490 575 510 675
rect 545 575 705 675
rect 740 575 760 675
rect 795 575 955 675
rect 990 575 1010 675
rect 1045 575 1205 675
rect 1240 575 1260 675
rect 1295 575 1455 675
rect 1490 575 1510 675
rect 1545 575 1705 675
rect 1740 575 1760 675
rect 1795 575 1955 675
rect 1990 575 2010 675
rect 2045 575 2205 675
rect 2240 575 2260 675
rect 2295 575 2455 675
rect 2490 575 2510 675
rect 2545 575 2705 675
rect 2740 575 2760 675
rect 2795 575 2955 675
rect 2990 575 3010 675
rect 3045 575 3205 675
rect 3240 575 3260 675
rect 3295 575 3455 675
rect 3490 575 3510 675
rect 3545 575 3705 675
rect 3740 575 3760 675
rect 3795 575 3955 675
rect 3990 575 4000 675
rect 0 570 4000 575
rect 70 545 180 570
rect 70 510 75 545
rect 175 510 180 545
rect 70 490 180 510
rect 70 455 75 490
rect 175 455 180 490
rect 70 430 180 455
rect 320 545 430 570
rect 320 510 325 545
rect 425 510 430 545
rect 320 490 430 510
rect 320 455 325 490
rect 425 455 430 490
rect 320 430 430 455
rect 570 545 680 570
rect 570 510 575 545
rect 675 510 680 545
rect 570 490 680 510
rect 570 455 575 490
rect 675 455 680 490
rect 570 430 680 455
rect 820 545 930 570
rect 820 510 825 545
rect 925 510 930 545
rect 820 490 930 510
rect 820 455 825 490
rect 925 455 930 490
rect 820 430 930 455
rect 1070 545 1180 570
rect 1070 510 1075 545
rect 1175 510 1180 545
rect 1070 490 1180 510
rect 1070 455 1075 490
rect 1175 455 1180 490
rect 1070 430 1180 455
rect 1320 545 1430 570
rect 1320 510 1325 545
rect 1425 510 1430 545
rect 1320 490 1430 510
rect 1320 455 1325 490
rect 1425 455 1430 490
rect 1320 430 1430 455
rect 1570 545 1680 570
rect 1570 510 1575 545
rect 1675 510 1680 545
rect 1570 490 1680 510
rect 1570 455 1575 490
rect 1675 455 1680 490
rect 1570 430 1680 455
rect 1820 545 1930 570
rect 1820 510 1825 545
rect 1925 510 1930 545
rect 1820 490 1930 510
rect 1820 455 1825 490
rect 1925 455 1930 490
rect 1820 430 1930 455
rect 2070 545 2180 570
rect 2070 510 2075 545
rect 2175 510 2180 545
rect 2070 490 2180 510
rect 2070 455 2075 490
rect 2175 455 2180 490
rect 2070 430 2180 455
rect 2320 545 2430 570
rect 2320 510 2325 545
rect 2425 510 2430 545
rect 2320 490 2430 510
rect 2320 455 2325 490
rect 2425 455 2430 490
rect 2320 430 2430 455
rect 2570 545 2680 570
rect 2570 510 2575 545
rect 2675 510 2680 545
rect 2570 490 2680 510
rect 2570 455 2575 490
rect 2675 455 2680 490
rect 2570 430 2680 455
rect 2820 545 2930 570
rect 2820 510 2825 545
rect 2925 510 2930 545
rect 2820 490 2930 510
rect 2820 455 2825 490
rect 2925 455 2930 490
rect 2820 430 2930 455
rect 3070 545 3180 570
rect 3070 510 3075 545
rect 3175 510 3180 545
rect 3070 490 3180 510
rect 3070 455 3075 490
rect 3175 455 3180 490
rect 3070 430 3180 455
rect 3320 545 3430 570
rect 3320 510 3325 545
rect 3425 510 3430 545
rect 3320 490 3430 510
rect 3320 455 3325 490
rect 3425 455 3430 490
rect 3320 430 3430 455
rect 3570 545 3680 570
rect 3570 510 3575 545
rect 3675 510 3680 545
rect 3570 490 3680 510
rect 3570 455 3575 490
rect 3675 455 3680 490
rect 3570 430 3680 455
rect 3820 545 3930 570
rect 3820 510 3825 545
rect 3925 510 3930 545
rect 3820 490 3930 510
rect 3820 455 3825 490
rect 3925 455 3930 490
rect 3820 430 3930 455
rect 0 425 4000 430
rect 0 325 10 425
rect 45 325 205 425
rect 240 325 260 425
rect 295 325 455 425
rect 490 325 510 425
rect 545 325 705 425
rect 740 325 760 425
rect 795 325 955 425
rect 990 325 1010 425
rect 1045 325 1205 425
rect 1240 325 1260 425
rect 1295 325 1455 425
rect 1490 325 1510 425
rect 1545 325 1705 425
rect 1740 325 1760 425
rect 1795 325 1955 425
rect 1990 325 2010 425
rect 2045 325 2205 425
rect 2240 325 2260 425
rect 2295 325 2455 425
rect 2490 325 2510 425
rect 2545 325 2705 425
rect 2740 325 2760 425
rect 2795 325 2955 425
rect 2990 325 3010 425
rect 3045 325 3205 425
rect 3240 325 3260 425
rect 3295 325 3455 425
rect 3490 325 3510 425
rect 3545 325 3705 425
rect 3740 325 3760 425
rect 3795 325 3955 425
rect 3990 325 4000 425
rect 0 320 4000 325
rect 70 295 180 320
rect 70 260 75 295
rect 175 260 180 295
rect 70 240 180 260
rect 70 205 75 240
rect 175 205 180 240
rect 70 180 180 205
rect 320 295 430 320
rect 320 260 325 295
rect 425 260 430 295
rect 320 240 430 260
rect 320 205 325 240
rect 425 205 430 240
rect 320 180 430 205
rect 570 295 680 320
rect 570 260 575 295
rect 675 260 680 295
rect 570 240 680 260
rect 570 205 575 240
rect 675 205 680 240
rect 570 180 680 205
rect 820 295 930 320
rect 820 260 825 295
rect 925 260 930 295
rect 820 240 930 260
rect 820 205 825 240
rect 925 205 930 240
rect 820 180 930 205
rect 1070 295 1180 320
rect 1070 260 1075 295
rect 1175 260 1180 295
rect 1070 240 1180 260
rect 1070 205 1075 240
rect 1175 205 1180 240
rect 1070 180 1180 205
rect 1320 295 1430 320
rect 1320 260 1325 295
rect 1425 260 1430 295
rect 1320 240 1430 260
rect 1320 205 1325 240
rect 1425 205 1430 240
rect 1320 180 1430 205
rect 1570 295 1680 320
rect 1570 260 1575 295
rect 1675 260 1680 295
rect 1570 240 1680 260
rect 1570 205 1575 240
rect 1675 205 1680 240
rect 1570 180 1680 205
rect 1820 295 1930 320
rect 1820 260 1825 295
rect 1925 260 1930 295
rect 1820 240 1930 260
rect 1820 205 1825 240
rect 1925 205 1930 240
rect 1820 180 1930 205
rect 2070 295 2180 320
rect 2070 260 2075 295
rect 2175 260 2180 295
rect 2070 240 2180 260
rect 2070 205 2075 240
rect 2175 205 2180 240
rect 2070 180 2180 205
rect 2320 295 2430 320
rect 2320 260 2325 295
rect 2425 260 2430 295
rect 2320 240 2430 260
rect 2320 205 2325 240
rect 2425 205 2430 240
rect 2320 180 2430 205
rect 2570 295 2680 320
rect 2570 260 2575 295
rect 2675 260 2680 295
rect 2570 240 2680 260
rect 2570 205 2575 240
rect 2675 205 2680 240
rect 2570 180 2680 205
rect 2820 295 2930 320
rect 2820 260 2825 295
rect 2925 260 2930 295
rect 2820 240 2930 260
rect 2820 205 2825 240
rect 2925 205 2930 240
rect 2820 180 2930 205
rect 3070 295 3180 320
rect 3070 260 3075 295
rect 3175 260 3180 295
rect 3070 240 3180 260
rect 3070 205 3075 240
rect 3175 205 3180 240
rect 3070 180 3180 205
rect 3320 295 3430 320
rect 3320 260 3325 295
rect 3425 260 3430 295
rect 3320 240 3430 260
rect 3320 205 3325 240
rect 3425 205 3430 240
rect 3320 180 3430 205
rect 3570 295 3680 320
rect 3570 260 3575 295
rect 3675 260 3680 295
rect 3570 240 3680 260
rect 3570 205 3575 240
rect 3675 205 3680 240
rect 3570 180 3680 205
rect 3820 295 3930 320
rect 3820 260 3825 295
rect 3925 260 3930 295
rect 3820 240 3930 260
rect 3820 205 3825 240
rect 3925 205 3930 240
rect 3820 180 3930 205
rect 0 175 4000 180
rect 0 75 10 175
rect 45 75 205 175
rect 240 75 260 175
rect 295 75 455 175
rect 490 75 510 175
rect 545 75 705 175
rect 740 75 760 175
rect 795 75 955 175
rect 990 75 1010 175
rect 1045 75 1205 175
rect 1240 75 1260 175
rect 1295 75 1455 175
rect 1490 75 1510 175
rect 1545 75 1705 175
rect 1740 75 1760 175
rect 1795 75 1955 175
rect 1990 75 2010 175
rect 2045 75 2205 175
rect 2240 75 2260 175
rect 2295 75 2455 175
rect 2490 75 2510 175
rect 2545 75 2705 175
rect 2740 75 2760 175
rect 2795 75 2955 175
rect 2990 75 3010 175
rect 3045 75 3205 175
rect 3240 75 3260 175
rect 3295 75 3455 175
rect 3490 75 3510 175
rect 3545 75 3705 175
rect 3740 75 3760 175
rect 3795 75 3955 175
rect 3990 75 4000 175
rect 0 70 4000 75
rect 70 45 180 70
rect 70 10 75 45
rect 175 10 180 45
rect 70 0 180 10
rect 320 45 430 70
rect 320 10 325 45
rect 425 10 430 45
rect 320 0 430 10
rect 570 45 680 70
rect 570 10 575 45
rect 675 10 680 45
rect 570 0 680 10
rect 820 45 930 70
rect 820 10 825 45
rect 925 10 930 45
rect 820 0 930 10
rect 1070 45 1180 70
rect 1070 10 1075 45
rect 1175 10 1180 45
rect 1070 0 1180 10
rect 1320 45 1430 70
rect 1320 10 1325 45
rect 1425 10 1430 45
rect 1320 0 1430 10
rect 1570 45 1680 70
rect 1570 10 1575 45
rect 1675 10 1680 45
rect 1570 0 1680 10
rect 1820 45 1930 70
rect 1820 10 1825 45
rect 1925 10 1930 45
rect 1820 0 1930 10
rect 2070 45 2180 70
rect 2070 10 2075 45
rect 2175 10 2180 45
rect 2070 0 2180 10
rect 2320 45 2430 70
rect 2320 10 2325 45
rect 2425 10 2430 45
rect 2320 0 2430 10
rect 2570 45 2680 70
rect 2570 10 2575 45
rect 2675 10 2680 45
rect 2570 0 2680 10
rect 2820 45 2930 70
rect 2820 10 2825 45
rect 2925 10 2930 45
rect 2820 0 2930 10
rect 3070 45 3180 70
rect 3070 10 3075 45
rect 3175 10 3180 45
rect 3070 0 3180 10
rect 3320 45 3430 70
rect 3320 10 3325 45
rect 3425 10 3430 45
rect 3320 0 3430 10
rect 3570 45 3680 70
rect 3570 10 3575 45
rect 3675 10 3680 45
rect 3570 0 3680 10
rect 3820 45 3930 70
rect 3820 10 3825 45
rect 3925 10 3930 45
rect 3820 0 3930 10
<< via2 >>
rect 75 3955 175 3990
rect 325 3955 425 3990
rect 575 3955 675 3990
rect 825 3955 925 3990
rect 1075 3955 1175 3990
rect 1325 3955 1425 3990
rect 1575 3955 1675 3990
rect 1825 3955 1925 3990
rect 2075 3955 2175 3990
rect 2325 3955 2425 3990
rect 2575 3955 2675 3990
rect 2825 3955 2925 3990
rect 3075 3955 3175 3990
rect 3325 3955 3425 3990
rect 3575 3955 3675 3990
rect 3825 3955 3925 3990
rect 10 3825 45 3925
rect 205 3825 240 3925
rect 260 3825 295 3925
rect 455 3825 490 3925
rect 510 3825 545 3925
rect 705 3825 740 3925
rect 760 3825 795 3925
rect 955 3825 990 3925
rect 1010 3825 1045 3925
rect 1205 3825 1240 3925
rect 1260 3825 1295 3925
rect 1455 3825 1490 3925
rect 1510 3825 1545 3925
rect 1705 3825 1740 3925
rect 1760 3825 1795 3925
rect 1955 3825 1990 3925
rect 2010 3825 2045 3925
rect 2205 3825 2240 3925
rect 2260 3825 2295 3925
rect 2455 3825 2490 3925
rect 2510 3825 2545 3925
rect 2705 3825 2740 3925
rect 2760 3825 2795 3925
rect 2955 3825 2990 3925
rect 3010 3825 3045 3925
rect 3205 3825 3240 3925
rect 3260 3825 3295 3925
rect 3455 3825 3490 3925
rect 3510 3825 3545 3925
rect 3705 3825 3740 3925
rect 3760 3825 3795 3925
rect 3955 3825 3990 3925
rect 75 3760 175 3795
rect 75 3705 175 3740
rect 325 3760 425 3795
rect 325 3705 425 3740
rect 575 3760 675 3795
rect 575 3705 675 3740
rect 825 3760 925 3795
rect 825 3705 925 3740
rect 1075 3760 1175 3795
rect 1075 3705 1175 3740
rect 1325 3760 1425 3795
rect 1325 3705 1425 3740
rect 1575 3760 1675 3795
rect 1575 3705 1675 3740
rect 1825 3760 1925 3795
rect 1825 3705 1925 3740
rect 2075 3760 2175 3795
rect 2075 3705 2175 3740
rect 2325 3760 2425 3795
rect 2325 3705 2425 3740
rect 2575 3760 2675 3795
rect 2575 3705 2675 3740
rect 2825 3760 2925 3795
rect 2825 3705 2925 3740
rect 3075 3760 3175 3795
rect 3075 3705 3175 3740
rect 3325 3760 3425 3795
rect 3325 3705 3425 3740
rect 3575 3760 3675 3795
rect 3575 3705 3675 3740
rect 3825 3760 3925 3795
rect 3825 3705 3925 3740
rect 10 3575 45 3675
rect 205 3575 240 3675
rect 260 3575 295 3675
rect 455 3575 490 3675
rect 510 3575 545 3675
rect 705 3575 740 3675
rect 760 3575 795 3675
rect 955 3575 990 3675
rect 1010 3575 1045 3675
rect 1205 3575 1240 3675
rect 1260 3575 1295 3675
rect 1455 3575 1490 3675
rect 1510 3575 1545 3675
rect 1705 3575 1740 3675
rect 1760 3575 1795 3675
rect 1955 3575 1990 3675
rect 2010 3575 2045 3675
rect 2205 3575 2240 3675
rect 2260 3575 2295 3675
rect 2455 3575 2490 3675
rect 2510 3575 2545 3675
rect 2705 3575 2740 3675
rect 2760 3575 2795 3675
rect 2955 3575 2990 3675
rect 3010 3575 3045 3675
rect 3205 3575 3240 3675
rect 3260 3575 3295 3675
rect 3455 3575 3490 3675
rect 3510 3575 3545 3675
rect 3705 3575 3740 3675
rect 3760 3575 3795 3675
rect 3955 3575 3990 3675
rect 75 3510 175 3545
rect 75 3455 175 3490
rect 325 3510 425 3545
rect 325 3455 425 3490
rect 575 3510 675 3545
rect 575 3455 675 3490
rect 825 3510 925 3545
rect 825 3455 925 3490
rect 1075 3510 1175 3545
rect 1075 3455 1175 3490
rect 1325 3510 1425 3545
rect 1325 3455 1425 3490
rect 1575 3510 1675 3545
rect 1575 3455 1675 3490
rect 1825 3510 1925 3545
rect 1825 3455 1925 3490
rect 2075 3510 2175 3545
rect 2075 3455 2175 3490
rect 2325 3510 2425 3545
rect 2325 3455 2425 3490
rect 2575 3510 2675 3545
rect 2575 3455 2675 3490
rect 2825 3510 2925 3545
rect 2825 3455 2925 3490
rect 3075 3510 3175 3545
rect 3075 3455 3175 3490
rect 3325 3510 3425 3545
rect 3325 3455 3425 3490
rect 3575 3510 3675 3545
rect 3575 3455 3675 3490
rect 3825 3510 3925 3545
rect 3825 3455 3925 3490
rect 10 3325 45 3425
rect 205 3325 240 3425
rect 260 3325 295 3425
rect 455 3325 490 3425
rect 510 3325 545 3425
rect 705 3325 740 3425
rect 760 3325 795 3425
rect 955 3325 990 3425
rect 1010 3325 1045 3425
rect 1205 3325 1240 3425
rect 1260 3325 1295 3425
rect 1455 3325 1490 3425
rect 1510 3325 1545 3425
rect 1705 3325 1740 3425
rect 1760 3325 1795 3425
rect 1955 3325 1990 3425
rect 2010 3325 2045 3425
rect 2205 3325 2240 3425
rect 2260 3325 2295 3425
rect 2455 3325 2490 3425
rect 2510 3325 2545 3425
rect 2705 3325 2740 3425
rect 2760 3325 2795 3425
rect 2955 3325 2990 3425
rect 3010 3325 3045 3425
rect 3205 3325 3240 3425
rect 3260 3325 3295 3425
rect 3455 3325 3490 3425
rect 3510 3325 3545 3425
rect 3705 3325 3740 3425
rect 3760 3325 3795 3425
rect 3955 3325 3990 3425
rect 75 3260 175 3295
rect 75 3205 175 3240
rect 325 3260 425 3295
rect 325 3205 425 3240
rect 575 3260 675 3295
rect 575 3205 675 3240
rect 825 3260 925 3295
rect 825 3205 925 3240
rect 1075 3260 1175 3295
rect 1075 3205 1175 3240
rect 1325 3260 1425 3295
rect 1325 3205 1425 3240
rect 1575 3260 1675 3295
rect 1575 3205 1675 3240
rect 1825 3260 1925 3295
rect 1825 3205 1925 3240
rect 2075 3260 2175 3295
rect 2075 3205 2175 3240
rect 2325 3260 2425 3295
rect 2325 3205 2425 3240
rect 2575 3260 2675 3295
rect 2575 3205 2675 3240
rect 2825 3260 2925 3295
rect 2825 3205 2925 3240
rect 3075 3260 3175 3295
rect 3075 3205 3175 3240
rect 3325 3260 3425 3295
rect 3325 3205 3425 3240
rect 3575 3260 3675 3295
rect 3575 3205 3675 3240
rect 3825 3260 3925 3295
rect 3825 3205 3925 3240
rect 10 3075 45 3175
rect 205 3075 240 3175
rect 260 3075 295 3175
rect 455 3075 490 3175
rect 510 3075 545 3175
rect 705 3075 740 3175
rect 760 3075 795 3175
rect 955 3075 990 3175
rect 1010 3075 1045 3175
rect 1205 3075 1240 3175
rect 1260 3075 1295 3175
rect 1455 3075 1490 3175
rect 1510 3075 1545 3175
rect 1705 3075 1740 3175
rect 1760 3075 1795 3175
rect 1955 3075 1990 3175
rect 2010 3075 2045 3175
rect 2205 3075 2240 3175
rect 2260 3075 2295 3175
rect 2455 3075 2490 3175
rect 2510 3075 2545 3175
rect 2705 3075 2740 3175
rect 2760 3075 2795 3175
rect 2955 3075 2990 3175
rect 3010 3075 3045 3175
rect 3205 3075 3240 3175
rect 3260 3075 3295 3175
rect 3455 3075 3490 3175
rect 3510 3075 3545 3175
rect 3705 3075 3740 3175
rect 3760 3075 3795 3175
rect 3955 3075 3990 3175
rect 75 3010 175 3045
rect 75 2955 175 2990
rect 325 3010 425 3045
rect 325 2955 425 2990
rect 575 3010 675 3045
rect 575 2955 675 2990
rect 825 3010 925 3045
rect 825 2955 925 2990
rect 1075 3010 1175 3045
rect 1075 2955 1175 2990
rect 1325 3010 1425 3045
rect 1325 2955 1425 2990
rect 1575 3010 1675 3045
rect 1575 2955 1675 2990
rect 1825 3010 1925 3045
rect 1825 2955 1925 2990
rect 2075 3010 2175 3045
rect 2075 2955 2175 2990
rect 2325 3010 2425 3045
rect 2325 2955 2425 2990
rect 2575 3010 2675 3045
rect 2575 2955 2675 2990
rect 2825 3010 2925 3045
rect 2825 2955 2925 2990
rect 3075 3010 3175 3045
rect 3075 2955 3175 2990
rect 3325 3010 3425 3045
rect 3325 2955 3425 2990
rect 3575 3010 3675 3045
rect 3575 2955 3675 2990
rect 3825 3010 3925 3045
rect 3825 2955 3925 2990
rect 10 2825 45 2925
rect 205 2825 240 2925
rect 260 2825 295 2925
rect 455 2825 490 2925
rect 510 2825 545 2925
rect 705 2825 740 2925
rect 760 2825 795 2925
rect 955 2825 990 2925
rect 1010 2825 1045 2925
rect 1205 2825 1240 2925
rect 1260 2825 1295 2925
rect 1455 2825 1490 2925
rect 1510 2825 1545 2925
rect 1705 2825 1740 2925
rect 1760 2825 1795 2925
rect 1955 2825 1990 2925
rect 2010 2825 2045 2925
rect 2205 2825 2240 2925
rect 2260 2825 2295 2925
rect 2455 2825 2490 2925
rect 2510 2825 2545 2925
rect 2705 2825 2740 2925
rect 2760 2825 2795 2925
rect 2955 2825 2990 2925
rect 3010 2825 3045 2925
rect 3205 2825 3240 2925
rect 3260 2825 3295 2925
rect 3455 2825 3490 2925
rect 3510 2825 3545 2925
rect 3705 2825 3740 2925
rect 3760 2825 3795 2925
rect 3955 2825 3990 2925
rect 75 2760 175 2795
rect 75 2705 175 2740
rect 325 2760 425 2795
rect 325 2705 425 2740
rect 575 2760 675 2795
rect 575 2705 675 2740
rect 825 2760 925 2795
rect 825 2705 925 2740
rect 1075 2760 1175 2795
rect 1075 2705 1175 2740
rect 1325 2760 1425 2795
rect 1325 2705 1425 2740
rect 1575 2760 1675 2795
rect 1575 2705 1675 2740
rect 1825 2760 1925 2795
rect 1825 2705 1925 2740
rect 2075 2760 2175 2795
rect 2075 2705 2175 2740
rect 2325 2760 2425 2795
rect 2325 2705 2425 2740
rect 2575 2760 2675 2795
rect 2575 2705 2675 2740
rect 2825 2760 2925 2795
rect 2825 2705 2925 2740
rect 3075 2760 3175 2795
rect 3075 2705 3175 2740
rect 3325 2760 3425 2795
rect 3325 2705 3425 2740
rect 3575 2760 3675 2795
rect 3575 2705 3675 2740
rect 3825 2760 3925 2795
rect 3825 2705 3925 2740
rect 10 2575 45 2675
rect 205 2575 240 2675
rect 260 2575 295 2675
rect 455 2575 490 2675
rect 510 2575 545 2675
rect 705 2575 740 2675
rect 760 2575 795 2675
rect 955 2575 990 2675
rect 1010 2575 1045 2675
rect 1205 2575 1240 2675
rect 1260 2575 1295 2675
rect 1455 2575 1490 2675
rect 1510 2575 1545 2675
rect 1705 2575 1740 2675
rect 1760 2575 1795 2675
rect 1955 2575 1990 2675
rect 2010 2575 2045 2675
rect 2205 2575 2240 2675
rect 2260 2575 2295 2675
rect 2455 2575 2490 2675
rect 2510 2575 2545 2675
rect 2705 2575 2740 2675
rect 2760 2575 2795 2675
rect 2955 2575 2990 2675
rect 3010 2575 3045 2675
rect 3205 2575 3240 2675
rect 3260 2575 3295 2675
rect 3455 2575 3490 2675
rect 3510 2575 3545 2675
rect 3705 2575 3740 2675
rect 3760 2575 3795 2675
rect 3955 2575 3990 2675
rect 75 2510 175 2545
rect 75 2455 175 2490
rect 325 2510 425 2545
rect 325 2455 425 2490
rect 575 2510 675 2545
rect 575 2455 675 2490
rect 825 2510 925 2545
rect 825 2455 925 2490
rect 1075 2510 1175 2545
rect 1075 2455 1175 2490
rect 1325 2510 1425 2545
rect 1325 2455 1425 2490
rect 1575 2510 1675 2545
rect 1575 2455 1675 2490
rect 1825 2510 1925 2545
rect 1825 2455 1925 2490
rect 2075 2510 2175 2545
rect 2075 2455 2175 2490
rect 2325 2510 2425 2545
rect 2325 2455 2425 2490
rect 2575 2510 2675 2545
rect 2575 2455 2675 2490
rect 2825 2510 2925 2545
rect 2825 2455 2925 2490
rect 3075 2510 3175 2545
rect 3075 2455 3175 2490
rect 3325 2510 3425 2545
rect 3325 2455 3425 2490
rect 3575 2510 3675 2545
rect 3575 2455 3675 2490
rect 3825 2510 3925 2545
rect 3825 2455 3925 2490
rect 10 2325 45 2425
rect 205 2325 240 2425
rect 260 2325 295 2425
rect 455 2325 490 2425
rect 510 2325 545 2425
rect 705 2325 740 2425
rect 760 2325 795 2425
rect 955 2325 990 2425
rect 1010 2325 1045 2425
rect 1205 2325 1240 2425
rect 1260 2325 1295 2425
rect 1455 2325 1490 2425
rect 1510 2325 1545 2425
rect 1705 2325 1740 2425
rect 1760 2325 1795 2425
rect 1955 2325 1990 2425
rect 2010 2325 2045 2425
rect 2205 2325 2240 2425
rect 2260 2325 2295 2425
rect 2455 2325 2490 2425
rect 2510 2325 2545 2425
rect 2705 2325 2740 2425
rect 2760 2325 2795 2425
rect 2955 2325 2990 2425
rect 3010 2325 3045 2425
rect 3205 2325 3240 2425
rect 3260 2325 3295 2425
rect 3455 2325 3490 2425
rect 3510 2325 3545 2425
rect 3705 2325 3740 2425
rect 3760 2325 3795 2425
rect 3955 2325 3990 2425
rect 75 2260 175 2295
rect 75 2205 175 2240
rect 325 2260 425 2295
rect 325 2205 425 2240
rect 575 2260 675 2295
rect 575 2205 675 2240
rect 825 2260 925 2295
rect 825 2205 925 2240
rect 1075 2260 1175 2295
rect 1075 2205 1175 2240
rect 1325 2260 1425 2295
rect 1325 2205 1425 2240
rect 1575 2260 1675 2295
rect 1575 2205 1675 2240
rect 1825 2260 1925 2295
rect 1825 2205 1925 2240
rect 2075 2260 2175 2295
rect 2075 2205 2175 2240
rect 2325 2260 2425 2295
rect 2325 2205 2425 2240
rect 2575 2260 2675 2295
rect 2575 2205 2675 2240
rect 2825 2260 2925 2295
rect 2825 2205 2925 2240
rect 3075 2260 3175 2295
rect 3075 2205 3175 2240
rect 3325 2260 3425 2295
rect 3325 2205 3425 2240
rect 3575 2260 3675 2295
rect 3575 2205 3675 2240
rect 3825 2260 3925 2295
rect 3825 2205 3925 2240
rect 10 2075 45 2175
rect 205 2075 240 2175
rect 260 2075 295 2175
rect 455 2075 490 2175
rect 510 2075 545 2175
rect 705 2075 740 2175
rect 760 2075 795 2175
rect 955 2075 990 2175
rect 1010 2075 1045 2175
rect 1205 2075 1240 2175
rect 1260 2075 1295 2175
rect 1455 2075 1490 2175
rect 1510 2075 1545 2175
rect 1705 2075 1740 2175
rect 1760 2075 1795 2175
rect 1955 2075 1990 2175
rect 2010 2075 2045 2175
rect 2205 2075 2240 2175
rect 2260 2075 2295 2175
rect 2455 2075 2490 2175
rect 2510 2075 2545 2175
rect 2705 2075 2740 2175
rect 2760 2075 2795 2175
rect 2955 2075 2990 2175
rect 3010 2075 3045 2175
rect 3205 2075 3240 2175
rect 3260 2075 3295 2175
rect 3455 2075 3490 2175
rect 3510 2075 3545 2175
rect 3705 2075 3740 2175
rect 3760 2075 3795 2175
rect 3955 2075 3990 2175
rect 75 2010 175 2045
rect 75 1955 175 1990
rect 325 2010 425 2045
rect 325 1955 425 1990
rect 575 2010 675 2045
rect 575 1955 675 1990
rect 825 2010 925 2045
rect 825 1955 925 1990
rect 1075 2010 1175 2045
rect 1075 1955 1175 1990
rect 1325 2010 1425 2045
rect 1325 1955 1425 1990
rect 1575 2010 1675 2045
rect 1575 1955 1675 1990
rect 1825 2010 1925 2045
rect 1825 1955 1925 1990
rect 2075 2010 2175 2045
rect 2075 1955 2175 1990
rect 2325 2010 2425 2045
rect 2325 1955 2425 1990
rect 2575 2010 2675 2045
rect 2575 1955 2675 1990
rect 2825 2010 2925 2045
rect 2825 1955 2925 1990
rect 3075 2010 3175 2045
rect 3075 1955 3175 1990
rect 3325 2010 3425 2045
rect 3325 1955 3425 1990
rect 3575 2010 3675 2045
rect 3575 1955 3675 1990
rect 3825 2010 3925 2045
rect 3825 1955 3925 1990
rect 10 1825 45 1925
rect 205 1825 240 1925
rect 260 1825 295 1925
rect 455 1825 490 1925
rect 510 1825 545 1925
rect 705 1825 740 1925
rect 760 1825 795 1925
rect 955 1825 990 1925
rect 1010 1825 1045 1925
rect 1205 1825 1240 1925
rect 1260 1825 1295 1925
rect 1455 1825 1490 1925
rect 1510 1825 1545 1925
rect 1705 1825 1740 1925
rect 1760 1825 1795 1925
rect 1955 1825 1990 1925
rect 2010 1825 2045 1925
rect 2205 1825 2240 1925
rect 2260 1825 2295 1925
rect 2455 1825 2490 1925
rect 2510 1825 2545 1925
rect 2705 1825 2740 1925
rect 2760 1825 2795 1925
rect 2955 1825 2990 1925
rect 3010 1825 3045 1925
rect 3205 1825 3240 1925
rect 3260 1825 3295 1925
rect 3455 1825 3490 1925
rect 3510 1825 3545 1925
rect 3705 1825 3740 1925
rect 3760 1825 3795 1925
rect 3955 1825 3990 1925
rect 75 1760 175 1795
rect 75 1705 175 1740
rect 325 1760 425 1795
rect 325 1705 425 1740
rect 575 1760 675 1795
rect 575 1705 675 1740
rect 825 1760 925 1795
rect 825 1705 925 1740
rect 1075 1760 1175 1795
rect 1075 1705 1175 1740
rect 1325 1760 1425 1795
rect 1325 1705 1425 1740
rect 1575 1760 1675 1795
rect 1575 1705 1675 1740
rect 1825 1760 1925 1795
rect 1825 1705 1925 1740
rect 2075 1760 2175 1795
rect 2075 1705 2175 1740
rect 2325 1760 2425 1795
rect 2325 1705 2425 1740
rect 2575 1760 2675 1795
rect 2575 1705 2675 1740
rect 2825 1760 2925 1795
rect 2825 1705 2925 1740
rect 3075 1760 3175 1795
rect 3075 1705 3175 1740
rect 3325 1760 3425 1795
rect 3325 1705 3425 1740
rect 3575 1760 3675 1795
rect 3575 1705 3675 1740
rect 3825 1760 3925 1795
rect 3825 1705 3925 1740
rect 10 1575 45 1675
rect 205 1575 240 1675
rect 260 1575 295 1675
rect 455 1575 490 1675
rect 510 1575 545 1675
rect 705 1575 740 1675
rect 760 1575 795 1675
rect 955 1575 990 1675
rect 1010 1575 1045 1675
rect 1205 1575 1240 1675
rect 1260 1575 1295 1675
rect 1455 1575 1490 1675
rect 1510 1575 1545 1675
rect 1705 1575 1740 1675
rect 1760 1575 1795 1675
rect 1955 1575 1990 1675
rect 2010 1575 2045 1675
rect 2205 1575 2240 1675
rect 2260 1575 2295 1675
rect 2455 1575 2490 1675
rect 2510 1575 2545 1675
rect 2705 1575 2740 1675
rect 2760 1575 2795 1675
rect 2955 1575 2990 1675
rect 3010 1575 3045 1675
rect 3205 1575 3240 1675
rect 3260 1575 3295 1675
rect 3455 1575 3490 1675
rect 3510 1575 3545 1675
rect 3705 1575 3740 1675
rect 3760 1575 3795 1675
rect 3955 1575 3990 1675
rect 75 1510 175 1545
rect 75 1455 175 1490
rect 325 1510 425 1545
rect 325 1455 425 1490
rect 575 1510 675 1545
rect 575 1455 675 1490
rect 825 1510 925 1545
rect 825 1455 925 1490
rect 1075 1510 1175 1545
rect 1075 1455 1175 1490
rect 1325 1510 1425 1545
rect 1325 1455 1425 1490
rect 1575 1510 1675 1545
rect 1575 1455 1675 1490
rect 1825 1510 1925 1545
rect 1825 1455 1925 1490
rect 2075 1510 2175 1545
rect 2075 1455 2175 1490
rect 2325 1510 2425 1545
rect 2325 1455 2425 1490
rect 2575 1510 2675 1545
rect 2575 1455 2675 1490
rect 2825 1510 2925 1545
rect 2825 1455 2925 1490
rect 3075 1510 3175 1545
rect 3075 1455 3175 1490
rect 3325 1510 3425 1545
rect 3325 1455 3425 1490
rect 3575 1510 3675 1545
rect 3575 1455 3675 1490
rect 3825 1510 3925 1545
rect 3825 1455 3925 1490
rect 10 1325 45 1425
rect 205 1325 240 1425
rect 260 1325 295 1425
rect 455 1325 490 1425
rect 510 1325 545 1425
rect 705 1325 740 1425
rect 760 1325 795 1425
rect 955 1325 990 1425
rect 1010 1325 1045 1425
rect 1205 1325 1240 1425
rect 1260 1325 1295 1425
rect 1455 1325 1490 1425
rect 1510 1325 1545 1425
rect 1705 1325 1740 1425
rect 1760 1325 1795 1425
rect 1955 1325 1990 1425
rect 2010 1325 2045 1425
rect 2205 1325 2240 1425
rect 2260 1325 2295 1425
rect 2455 1325 2490 1425
rect 2510 1325 2545 1425
rect 2705 1325 2740 1425
rect 2760 1325 2795 1425
rect 2955 1325 2990 1425
rect 3010 1325 3045 1425
rect 3205 1325 3240 1425
rect 3260 1325 3295 1425
rect 3455 1325 3490 1425
rect 3510 1325 3545 1425
rect 3705 1325 3740 1425
rect 3760 1325 3795 1425
rect 3955 1325 3990 1425
rect 75 1260 175 1295
rect 75 1205 175 1240
rect 325 1260 425 1295
rect 325 1205 425 1240
rect 575 1260 675 1295
rect 575 1205 675 1240
rect 825 1260 925 1295
rect 825 1205 925 1240
rect 1075 1260 1175 1295
rect 1075 1205 1175 1240
rect 1325 1260 1425 1295
rect 1325 1205 1425 1240
rect 1575 1260 1675 1295
rect 1575 1205 1675 1240
rect 1825 1260 1925 1295
rect 1825 1205 1925 1240
rect 2075 1260 2175 1295
rect 2075 1205 2175 1240
rect 2325 1260 2425 1295
rect 2325 1205 2425 1240
rect 2575 1260 2675 1295
rect 2575 1205 2675 1240
rect 2825 1260 2925 1295
rect 2825 1205 2925 1240
rect 3075 1260 3175 1295
rect 3075 1205 3175 1240
rect 3325 1260 3425 1295
rect 3325 1205 3425 1240
rect 3575 1260 3675 1295
rect 3575 1205 3675 1240
rect 3825 1260 3925 1295
rect 3825 1205 3925 1240
rect 10 1075 45 1175
rect 205 1075 240 1175
rect 260 1075 295 1175
rect 455 1075 490 1175
rect 510 1075 545 1175
rect 705 1075 740 1175
rect 760 1075 795 1175
rect 955 1075 990 1175
rect 1010 1075 1045 1175
rect 1205 1075 1240 1175
rect 1260 1075 1295 1175
rect 1455 1075 1490 1175
rect 1510 1075 1545 1175
rect 1705 1075 1740 1175
rect 1760 1075 1795 1175
rect 1955 1075 1990 1175
rect 2010 1075 2045 1175
rect 2205 1075 2240 1175
rect 2260 1075 2295 1175
rect 2455 1075 2490 1175
rect 2510 1075 2545 1175
rect 2705 1075 2740 1175
rect 2760 1075 2795 1175
rect 2955 1075 2990 1175
rect 3010 1075 3045 1175
rect 3205 1075 3240 1175
rect 3260 1075 3295 1175
rect 3455 1075 3490 1175
rect 3510 1075 3545 1175
rect 3705 1075 3740 1175
rect 3760 1075 3795 1175
rect 3955 1075 3990 1175
rect 75 1010 175 1045
rect 75 955 175 990
rect 325 1010 425 1045
rect 325 955 425 990
rect 575 1010 675 1045
rect 575 955 675 990
rect 825 1010 925 1045
rect 825 955 925 990
rect 1075 1010 1175 1045
rect 1075 955 1175 990
rect 1325 1010 1425 1045
rect 1325 955 1425 990
rect 1575 1010 1675 1045
rect 1575 955 1675 990
rect 1825 1010 1925 1045
rect 1825 955 1925 990
rect 2075 1010 2175 1045
rect 2075 955 2175 990
rect 2325 1010 2425 1045
rect 2325 955 2425 990
rect 2575 1010 2675 1045
rect 2575 955 2675 990
rect 2825 1010 2925 1045
rect 2825 955 2925 990
rect 3075 1010 3175 1045
rect 3075 955 3175 990
rect 3325 1010 3425 1045
rect 3325 955 3425 990
rect 3575 1010 3675 1045
rect 3575 955 3675 990
rect 3825 1010 3925 1045
rect 3825 955 3925 990
rect 10 825 45 925
rect 205 825 240 925
rect 260 825 295 925
rect 455 825 490 925
rect 510 825 545 925
rect 705 825 740 925
rect 760 825 795 925
rect 955 825 990 925
rect 1010 825 1045 925
rect 1205 825 1240 925
rect 1260 825 1295 925
rect 1455 825 1490 925
rect 1510 825 1545 925
rect 1705 825 1740 925
rect 1760 825 1795 925
rect 1955 825 1990 925
rect 2010 825 2045 925
rect 2205 825 2240 925
rect 2260 825 2295 925
rect 2455 825 2490 925
rect 2510 825 2545 925
rect 2705 825 2740 925
rect 2760 825 2795 925
rect 2955 825 2990 925
rect 3010 825 3045 925
rect 3205 825 3240 925
rect 3260 825 3295 925
rect 3455 825 3490 925
rect 3510 825 3545 925
rect 3705 825 3740 925
rect 3760 825 3795 925
rect 3955 825 3990 925
rect 75 760 175 795
rect 75 705 175 740
rect 325 760 425 795
rect 325 705 425 740
rect 575 760 675 795
rect 575 705 675 740
rect 825 760 925 795
rect 825 705 925 740
rect 1075 760 1175 795
rect 1075 705 1175 740
rect 1325 760 1425 795
rect 1325 705 1425 740
rect 1575 760 1675 795
rect 1575 705 1675 740
rect 1825 760 1925 795
rect 1825 705 1925 740
rect 2075 760 2175 795
rect 2075 705 2175 740
rect 2325 760 2425 795
rect 2325 705 2425 740
rect 2575 760 2675 795
rect 2575 705 2675 740
rect 2825 760 2925 795
rect 2825 705 2925 740
rect 3075 760 3175 795
rect 3075 705 3175 740
rect 3325 760 3425 795
rect 3325 705 3425 740
rect 3575 760 3675 795
rect 3575 705 3675 740
rect 3825 760 3925 795
rect 3825 705 3925 740
rect 10 575 45 675
rect 205 575 240 675
rect 260 575 295 675
rect 455 575 490 675
rect 510 575 545 675
rect 705 575 740 675
rect 760 575 795 675
rect 955 575 990 675
rect 1010 575 1045 675
rect 1205 575 1240 675
rect 1260 575 1295 675
rect 1455 575 1490 675
rect 1510 575 1545 675
rect 1705 575 1740 675
rect 1760 575 1795 675
rect 1955 575 1990 675
rect 2010 575 2045 675
rect 2205 575 2240 675
rect 2260 575 2295 675
rect 2455 575 2490 675
rect 2510 575 2545 675
rect 2705 575 2740 675
rect 2760 575 2795 675
rect 2955 575 2990 675
rect 3010 575 3045 675
rect 3205 575 3240 675
rect 3260 575 3295 675
rect 3455 575 3490 675
rect 3510 575 3545 675
rect 3705 575 3740 675
rect 3760 575 3795 675
rect 3955 575 3990 675
rect 75 510 175 545
rect 75 455 175 490
rect 325 510 425 545
rect 325 455 425 490
rect 575 510 675 545
rect 575 455 675 490
rect 825 510 925 545
rect 825 455 925 490
rect 1075 510 1175 545
rect 1075 455 1175 490
rect 1325 510 1425 545
rect 1325 455 1425 490
rect 1575 510 1675 545
rect 1575 455 1675 490
rect 1825 510 1925 545
rect 1825 455 1925 490
rect 2075 510 2175 545
rect 2075 455 2175 490
rect 2325 510 2425 545
rect 2325 455 2425 490
rect 2575 510 2675 545
rect 2575 455 2675 490
rect 2825 510 2925 545
rect 2825 455 2925 490
rect 3075 510 3175 545
rect 3075 455 3175 490
rect 3325 510 3425 545
rect 3325 455 3425 490
rect 3575 510 3675 545
rect 3575 455 3675 490
rect 3825 510 3925 545
rect 3825 455 3925 490
rect 10 325 45 425
rect 205 325 240 425
rect 260 325 295 425
rect 455 325 490 425
rect 510 325 545 425
rect 705 325 740 425
rect 760 325 795 425
rect 955 325 990 425
rect 1010 325 1045 425
rect 1205 325 1240 425
rect 1260 325 1295 425
rect 1455 325 1490 425
rect 1510 325 1545 425
rect 1705 325 1740 425
rect 1760 325 1795 425
rect 1955 325 1990 425
rect 2010 325 2045 425
rect 2205 325 2240 425
rect 2260 325 2295 425
rect 2455 325 2490 425
rect 2510 325 2545 425
rect 2705 325 2740 425
rect 2760 325 2795 425
rect 2955 325 2990 425
rect 3010 325 3045 425
rect 3205 325 3240 425
rect 3260 325 3295 425
rect 3455 325 3490 425
rect 3510 325 3545 425
rect 3705 325 3740 425
rect 3760 325 3795 425
rect 3955 325 3990 425
rect 75 260 175 295
rect 75 205 175 240
rect 325 260 425 295
rect 325 205 425 240
rect 575 260 675 295
rect 575 205 675 240
rect 825 260 925 295
rect 825 205 925 240
rect 1075 260 1175 295
rect 1075 205 1175 240
rect 1325 260 1425 295
rect 1325 205 1425 240
rect 1575 260 1675 295
rect 1575 205 1675 240
rect 1825 260 1925 295
rect 1825 205 1925 240
rect 2075 260 2175 295
rect 2075 205 2175 240
rect 2325 260 2425 295
rect 2325 205 2425 240
rect 2575 260 2675 295
rect 2575 205 2675 240
rect 2825 260 2925 295
rect 2825 205 2925 240
rect 3075 260 3175 295
rect 3075 205 3175 240
rect 3325 260 3425 295
rect 3325 205 3425 240
rect 3575 260 3675 295
rect 3575 205 3675 240
rect 3825 260 3925 295
rect 3825 205 3925 240
rect 10 75 45 175
rect 205 75 240 175
rect 260 75 295 175
rect 455 75 490 175
rect 510 75 545 175
rect 705 75 740 175
rect 760 75 795 175
rect 955 75 990 175
rect 1010 75 1045 175
rect 1205 75 1240 175
rect 1260 75 1295 175
rect 1455 75 1490 175
rect 1510 75 1545 175
rect 1705 75 1740 175
rect 1760 75 1795 175
rect 1955 75 1990 175
rect 2010 75 2045 175
rect 2205 75 2240 175
rect 2260 75 2295 175
rect 2455 75 2490 175
rect 2510 75 2545 175
rect 2705 75 2740 175
rect 2760 75 2795 175
rect 2955 75 2990 175
rect 3010 75 3045 175
rect 3205 75 3240 175
rect 3260 75 3295 175
rect 3455 75 3490 175
rect 3510 75 3545 175
rect 3705 75 3740 175
rect 3760 75 3795 175
rect 3955 75 3990 175
rect 75 10 175 45
rect 325 10 425 45
rect 575 10 675 45
rect 825 10 925 45
rect 1075 10 1175 45
rect 1325 10 1425 45
rect 1575 10 1675 45
rect 1825 10 1925 45
rect 2075 10 2175 45
rect 2325 10 2425 45
rect 2575 10 2675 45
rect 2825 10 2925 45
rect 3075 10 3175 45
rect 3325 10 3425 45
rect 3575 10 3675 45
rect 3825 10 3925 45
<< metal3 >>
rect 0 3990 4000 4000
rect 0 3955 75 3990
rect 175 3955 325 3990
rect 425 3955 575 3990
rect 675 3955 825 3990
rect 925 3955 1075 3990
rect 1175 3955 1325 3990
rect 1425 3955 1575 3990
rect 1675 3955 1825 3990
rect 1925 3955 2075 3990
rect 2175 3955 2325 3990
rect 2425 3955 2575 3990
rect 2675 3955 2825 3990
rect 2925 3955 3075 3990
rect 3175 3955 3325 3990
rect 3425 3955 3575 3990
rect 3675 3955 3825 3990
rect 3925 3955 4000 3990
rect 0 3950 4000 3955
rect 0 3940 60 3950
rect 190 3940 310 3950
rect 440 3940 560 3950
rect 690 3940 810 3950
rect 940 3940 1060 3950
rect 1190 3940 1310 3950
rect 1440 3940 1560 3950
rect 1690 3940 1810 3950
rect 1940 3940 2060 3950
rect 2190 3940 2310 3950
rect 2440 3940 2560 3950
rect 2690 3940 2810 3950
rect 2940 3940 3060 3950
rect 3190 3940 3310 3950
rect 3440 3940 3560 3950
rect 3690 3940 3810 3950
rect 3940 3940 4000 3950
rect 0 3925 50 3940
rect 0 3825 10 3925
rect 45 3825 50 3925
rect 0 3810 50 3825
rect 200 3925 300 3940
rect 200 3825 205 3925
rect 240 3825 260 3925
rect 295 3825 300 3925
rect 200 3810 300 3825
rect 450 3925 550 3940
rect 450 3825 455 3925
rect 490 3825 510 3925
rect 545 3825 550 3925
rect 450 3810 550 3825
rect 700 3925 800 3940
rect 700 3825 705 3925
rect 740 3825 760 3925
rect 795 3825 800 3925
rect 700 3810 800 3825
rect 950 3925 1050 3940
rect 950 3825 955 3925
rect 990 3825 1010 3925
rect 1045 3825 1050 3925
rect 950 3810 1050 3825
rect 1200 3925 1300 3940
rect 1200 3825 1205 3925
rect 1240 3825 1260 3925
rect 1295 3825 1300 3925
rect 1200 3810 1300 3825
rect 1450 3925 1550 3940
rect 1450 3825 1455 3925
rect 1490 3825 1510 3925
rect 1545 3825 1550 3925
rect 1450 3810 1550 3825
rect 1700 3925 1800 3940
rect 1700 3825 1705 3925
rect 1740 3825 1760 3925
rect 1795 3825 1800 3925
rect 1700 3810 1800 3825
rect 1950 3925 2050 3940
rect 1950 3825 1955 3925
rect 1990 3825 2010 3925
rect 2045 3825 2050 3925
rect 1950 3810 2050 3825
rect 2200 3925 2300 3940
rect 2200 3825 2205 3925
rect 2240 3825 2260 3925
rect 2295 3825 2300 3925
rect 2200 3810 2300 3825
rect 2450 3925 2550 3940
rect 2450 3825 2455 3925
rect 2490 3825 2510 3925
rect 2545 3825 2550 3925
rect 2450 3810 2550 3825
rect 2700 3925 2800 3940
rect 2700 3825 2705 3925
rect 2740 3825 2760 3925
rect 2795 3825 2800 3925
rect 2700 3810 2800 3825
rect 2950 3925 3050 3940
rect 2950 3825 2955 3925
rect 2990 3825 3010 3925
rect 3045 3825 3050 3925
rect 2950 3810 3050 3825
rect 3200 3925 3300 3940
rect 3200 3825 3205 3925
rect 3240 3825 3260 3925
rect 3295 3825 3300 3925
rect 3200 3810 3300 3825
rect 3450 3925 3550 3940
rect 3450 3825 3455 3925
rect 3490 3825 3510 3925
rect 3545 3825 3550 3925
rect 3450 3810 3550 3825
rect 3700 3925 3800 3940
rect 3700 3825 3705 3925
rect 3740 3825 3760 3925
rect 3795 3825 3800 3925
rect 3700 3810 3800 3825
rect 3950 3925 4000 3940
rect 3950 3825 3955 3925
rect 3990 3825 4000 3925
rect 3950 3810 4000 3825
rect 0 3800 60 3810
rect 190 3800 310 3810
rect 440 3800 560 3810
rect 690 3800 810 3810
rect 940 3800 1060 3810
rect 1190 3800 1310 3810
rect 1440 3800 1560 3810
rect 1690 3800 1810 3810
rect 1940 3800 2060 3810
rect 2190 3800 2310 3810
rect 2440 3800 2560 3810
rect 2690 3800 2810 3810
rect 2940 3800 3060 3810
rect 3190 3800 3310 3810
rect 3440 3800 3560 3810
rect 3690 3800 3810 3810
rect 3940 3800 4000 3810
rect 0 3795 200 3800
rect 0 3760 75 3795
rect 175 3760 200 3795
rect 0 3740 200 3760
rect 0 3705 75 3740
rect 175 3705 200 3740
rect 0 3700 200 3705
rect 300 3795 450 3800
rect 300 3760 325 3795
rect 425 3760 450 3795
rect 300 3740 450 3760
rect 300 3705 325 3740
rect 425 3705 450 3740
rect 300 3700 450 3705
rect 550 3795 700 3800
rect 550 3760 575 3795
rect 675 3760 700 3795
rect 550 3740 700 3760
rect 550 3705 575 3740
rect 675 3705 700 3740
rect 550 3700 700 3705
rect 800 3795 1200 3800
rect 800 3760 825 3795
rect 925 3760 1075 3795
rect 1175 3760 1200 3795
rect 800 3740 1200 3760
rect 800 3705 825 3740
rect 925 3705 1075 3740
rect 1175 3705 1200 3740
rect 800 3700 1200 3705
rect 1300 3795 1450 3800
rect 1300 3760 1325 3795
rect 1425 3760 1450 3795
rect 1300 3740 1450 3760
rect 1300 3705 1325 3740
rect 1425 3705 1450 3740
rect 1300 3700 1450 3705
rect 1550 3795 1700 3800
rect 1550 3760 1575 3795
rect 1675 3760 1700 3795
rect 1550 3740 1700 3760
rect 1550 3705 1575 3740
rect 1675 3705 1700 3740
rect 1550 3700 1700 3705
rect 1800 3795 2200 3800
rect 1800 3760 1825 3795
rect 1925 3760 2075 3795
rect 2175 3760 2200 3795
rect 1800 3740 2200 3760
rect 1800 3705 1825 3740
rect 1925 3705 2075 3740
rect 2175 3705 2200 3740
rect 1800 3700 2200 3705
rect 2300 3795 2450 3800
rect 2300 3760 2325 3795
rect 2425 3760 2450 3795
rect 2300 3740 2450 3760
rect 2300 3705 2325 3740
rect 2425 3705 2450 3740
rect 2300 3700 2450 3705
rect 2550 3795 2700 3800
rect 2550 3760 2575 3795
rect 2675 3760 2700 3795
rect 2550 3740 2700 3760
rect 2550 3705 2575 3740
rect 2675 3705 2700 3740
rect 2550 3700 2700 3705
rect 2800 3795 3200 3800
rect 2800 3760 2825 3795
rect 2925 3760 3075 3795
rect 3175 3760 3200 3795
rect 2800 3740 3200 3760
rect 2800 3705 2825 3740
rect 2925 3705 3075 3740
rect 3175 3705 3200 3740
rect 2800 3700 3200 3705
rect 3300 3795 3450 3800
rect 3300 3760 3325 3795
rect 3425 3760 3450 3795
rect 3300 3740 3450 3760
rect 3300 3705 3325 3740
rect 3425 3705 3450 3740
rect 3300 3700 3450 3705
rect 3550 3795 3700 3800
rect 3550 3760 3575 3795
rect 3675 3760 3700 3795
rect 3550 3740 3700 3760
rect 3550 3705 3575 3740
rect 3675 3705 3700 3740
rect 3550 3700 3700 3705
rect 3800 3795 4000 3800
rect 3800 3760 3825 3795
rect 3925 3760 4000 3795
rect 3800 3740 4000 3760
rect 3800 3705 3825 3740
rect 3925 3705 4000 3740
rect 3800 3700 4000 3705
rect 0 3690 60 3700
rect 190 3690 310 3700
rect 440 3690 560 3700
rect 690 3690 810 3700
rect 940 3690 1060 3700
rect 1190 3690 1310 3700
rect 1440 3690 1560 3700
rect 1690 3690 1810 3700
rect 1940 3690 2060 3700
rect 2190 3690 2310 3700
rect 2440 3690 2560 3700
rect 2690 3690 2810 3700
rect 2940 3690 3060 3700
rect 3190 3690 3310 3700
rect 3440 3690 3560 3700
rect 3690 3690 3810 3700
rect 3940 3690 4000 3700
rect 0 3675 50 3690
rect 0 3575 10 3675
rect 45 3575 50 3675
rect 0 3560 50 3575
rect 200 3675 300 3690
rect 200 3575 205 3675
rect 240 3575 260 3675
rect 295 3575 300 3675
rect 200 3560 300 3575
rect 450 3675 550 3690
rect 450 3575 455 3675
rect 490 3575 510 3675
rect 545 3575 550 3675
rect 450 3560 550 3575
rect 700 3675 800 3690
rect 700 3575 705 3675
rect 740 3575 760 3675
rect 795 3575 800 3675
rect 700 3560 800 3575
rect 950 3675 1050 3690
rect 950 3575 955 3675
rect 990 3575 1010 3675
rect 1045 3575 1050 3675
rect 950 3560 1050 3575
rect 1200 3675 1300 3690
rect 1200 3575 1205 3675
rect 1240 3575 1260 3675
rect 1295 3575 1300 3675
rect 1200 3560 1300 3575
rect 1450 3675 1550 3690
rect 1450 3575 1455 3675
rect 1490 3575 1510 3675
rect 1545 3575 1550 3675
rect 1450 3560 1550 3575
rect 1700 3675 1800 3690
rect 1700 3575 1705 3675
rect 1740 3575 1760 3675
rect 1795 3575 1800 3675
rect 1700 3560 1800 3575
rect 1950 3675 2050 3690
rect 1950 3575 1955 3675
rect 1990 3575 2010 3675
rect 2045 3575 2050 3675
rect 1950 3560 2050 3575
rect 2200 3675 2300 3690
rect 2200 3575 2205 3675
rect 2240 3575 2260 3675
rect 2295 3575 2300 3675
rect 2200 3560 2300 3575
rect 2450 3675 2550 3690
rect 2450 3575 2455 3675
rect 2490 3575 2510 3675
rect 2545 3575 2550 3675
rect 2450 3560 2550 3575
rect 2700 3675 2800 3690
rect 2700 3575 2705 3675
rect 2740 3575 2760 3675
rect 2795 3575 2800 3675
rect 2700 3560 2800 3575
rect 2950 3675 3050 3690
rect 2950 3575 2955 3675
rect 2990 3575 3010 3675
rect 3045 3575 3050 3675
rect 2950 3560 3050 3575
rect 3200 3675 3300 3690
rect 3200 3575 3205 3675
rect 3240 3575 3260 3675
rect 3295 3575 3300 3675
rect 3200 3560 3300 3575
rect 3450 3675 3550 3690
rect 3450 3575 3455 3675
rect 3490 3575 3510 3675
rect 3545 3575 3550 3675
rect 3450 3560 3550 3575
rect 3700 3675 3800 3690
rect 3700 3575 3705 3675
rect 3740 3575 3760 3675
rect 3795 3575 3800 3675
rect 3700 3560 3800 3575
rect 3950 3675 4000 3690
rect 3950 3575 3955 3675
rect 3990 3575 4000 3675
rect 3950 3560 4000 3575
rect 0 3550 60 3560
rect 190 3550 310 3560
rect 440 3550 560 3560
rect 690 3550 810 3560
rect 940 3550 1060 3560
rect 1190 3550 1310 3560
rect 1440 3550 1560 3560
rect 1690 3550 1810 3560
rect 1940 3550 2060 3560
rect 2190 3550 2310 3560
rect 2440 3550 2560 3560
rect 2690 3550 2810 3560
rect 2940 3550 3060 3560
rect 3190 3550 3310 3560
rect 3440 3550 3560 3560
rect 3690 3550 3810 3560
rect 3940 3550 4000 3560
rect 0 3545 200 3550
rect 0 3510 75 3545
rect 175 3510 200 3545
rect 0 3490 200 3510
rect 0 3455 75 3490
rect 175 3455 200 3490
rect 0 3450 200 3455
rect 300 3545 450 3550
rect 300 3510 325 3545
rect 425 3510 450 3545
rect 300 3490 450 3510
rect 300 3455 325 3490
rect 425 3455 450 3490
rect 300 3450 450 3455
rect 550 3545 700 3550
rect 550 3510 575 3545
rect 675 3510 700 3545
rect 550 3490 700 3510
rect 550 3455 575 3490
rect 675 3455 700 3490
rect 550 3450 700 3455
rect 800 3545 950 3550
rect 800 3510 825 3545
rect 925 3510 950 3545
rect 800 3490 950 3510
rect 800 3455 825 3490
rect 925 3455 950 3490
rect 800 3450 950 3455
rect 1050 3545 1200 3550
rect 1050 3510 1075 3545
rect 1175 3510 1200 3545
rect 1050 3490 1200 3510
rect 1050 3455 1075 3490
rect 1175 3455 1200 3490
rect 1050 3450 1200 3455
rect 1300 3545 1450 3550
rect 1300 3510 1325 3545
rect 1425 3510 1450 3545
rect 1300 3490 1450 3510
rect 1300 3455 1325 3490
rect 1425 3455 1450 3490
rect 1300 3450 1450 3455
rect 1550 3545 1700 3550
rect 1550 3510 1575 3545
rect 1675 3510 1700 3545
rect 1550 3490 1700 3510
rect 1550 3455 1575 3490
rect 1675 3455 1700 3490
rect 1550 3450 1700 3455
rect 1800 3545 2200 3550
rect 1800 3510 1825 3545
rect 1925 3510 2075 3545
rect 2175 3510 2200 3545
rect 1800 3490 2200 3510
rect 1800 3455 1825 3490
rect 1925 3455 2075 3490
rect 2175 3455 2200 3490
rect 1800 3450 2200 3455
rect 2300 3545 2450 3550
rect 2300 3510 2325 3545
rect 2425 3510 2450 3545
rect 2300 3490 2450 3510
rect 2300 3455 2325 3490
rect 2425 3455 2450 3490
rect 2300 3450 2450 3455
rect 2550 3545 2700 3550
rect 2550 3510 2575 3545
rect 2675 3510 2700 3545
rect 2550 3490 2700 3510
rect 2550 3455 2575 3490
rect 2675 3455 2700 3490
rect 2550 3450 2700 3455
rect 2800 3545 2950 3550
rect 2800 3510 2825 3545
rect 2925 3510 2950 3545
rect 2800 3490 2950 3510
rect 2800 3455 2825 3490
rect 2925 3455 2950 3490
rect 2800 3450 2950 3455
rect 3050 3545 3200 3550
rect 3050 3510 3075 3545
rect 3175 3510 3200 3545
rect 3050 3490 3200 3510
rect 3050 3455 3075 3490
rect 3175 3455 3200 3490
rect 3050 3450 3200 3455
rect 3300 3545 3450 3550
rect 3300 3510 3325 3545
rect 3425 3510 3450 3545
rect 3300 3490 3450 3510
rect 3300 3455 3325 3490
rect 3425 3455 3450 3490
rect 3300 3450 3450 3455
rect 3550 3545 3700 3550
rect 3550 3510 3575 3545
rect 3675 3510 3700 3545
rect 3550 3490 3700 3510
rect 3550 3455 3575 3490
rect 3675 3455 3700 3490
rect 3550 3450 3700 3455
rect 3800 3545 4000 3550
rect 3800 3510 3825 3545
rect 3925 3510 4000 3545
rect 3800 3490 4000 3510
rect 3800 3455 3825 3490
rect 3925 3455 4000 3490
rect 3800 3450 4000 3455
rect 0 3440 60 3450
rect 190 3440 310 3450
rect 440 3440 560 3450
rect 690 3440 810 3450
rect 940 3440 1060 3450
rect 1190 3440 1310 3450
rect 1440 3440 1560 3450
rect 1690 3440 1810 3450
rect 1940 3440 2060 3450
rect 2190 3440 2310 3450
rect 2440 3440 2560 3450
rect 2690 3440 2810 3450
rect 2940 3440 3060 3450
rect 3190 3440 3310 3450
rect 3440 3440 3560 3450
rect 3690 3440 3810 3450
rect 3940 3440 4000 3450
rect 0 3425 50 3440
rect 0 3325 10 3425
rect 45 3325 50 3425
rect 0 3310 50 3325
rect 200 3425 300 3440
rect 200 3325 205 3425
rect 240 3325 260 3425
rect 295 3325 300 3425
rect 200 3310 300 3325
rect 450 3425 550 3440
rect 450 3325 455 3425
rect 490 3325 510 3425
rect 545 3325 550 3425
rect 450 3310 550 3325
rect 700 3425 800 3440
rect 700 3325 705 3425
rect 740 3325 760 3425
rect 795 3325 800 3425
rect 700 3310 800 3325
rect 950 3425 1050 3440
rect 950 3325 955 3425
rect 990 3325 1010 3425
rect 1045 3325 1050 3425
rect 950 3310 1050 3325
rect 1200 3425 1300 3440
rect 1200 3325 1205 3425
rect 1240 3325 1260 3425
rect 1295 3325 1300 3425
rect 1200 3310 1300 3325
rect 1450 3425 1550 3440
rect 1450 3325 1455 3425
rect 1490 3325 1510 3425
rect 1545 3325 1550 3425
rect 1450 3310 1550 3325
rect 1700 3425 1800 3440
rect 1700 3325 1705 3425
rect 1740 3325 1760 3425
rect 1795 3325 1800 3425
rect 1700 3310 1800 3325
rect 1950 3425 2050 3440
rect 1950 3325 1955 3425
rect 1990 3325 2010 3425
rect 2045 3325 2050 3425
rect 1950 3310 2050 3325
rect 2200 3425 2300 3440
rect 2200 3325 2205 3425
rect 2240 3325 2260 3425
rect 2295 3325 2300 3425
rect 2200 3310 2300 3325
rect 2450 3425 2550 3440
rect 2450 3325 2455 3425
rect 2490 3325 2510 3425
rect 2545 3325 2550 3425
rect 2450 3310 2550 3325
rect 2700 3425 2800 3440
rect 2700 3325 2705 3425
rect 2740 3325 2760 3425
rect 2795 3325 2800 3425
rect 2700 3310 2800 3325
rect 2950 3425 3050 3440
rect 2950 3325 2955 3425
rect 2990 3325 3010 3425
rect 3045 3325 3050 3425
rect 2950 3310 3050 3325
rect 3200 3425 3300 3440
rect 3200 3325 3205 3425
rect 3240 3325 3260 3425
rect 3295 3325 3300 3425
rect 3200 3310 3300 3325
rect 3450 3425 3550 3440
rect 3450 3325 3455 3425
rect 3490 3325 3510 3425
rect 3545 3325 3550 3425
rect 3450 3310 3550 3325
rect 3700 3425 3800 3440
rect 3700 3325 3705 3425
rect 3740 3325 3760 3425
rect 3795 3325 3800 3425
rect 3700 3310 3800 3325
rect 3950 3425 4000 3440
rect 3950 3325 3955 3425
rect 3990 3325 4000 3425
rect 3950 3310 4000 3325
rect 0 3300 60 3310
rect 190 3300 310 3310
rect 440 3300 560 3310
rect 690 3300 810 3310
rect 940 3300 1060 3310
rect 1190 3300 1310 3310
rect 1440 3300 1560 3310
rect 1690 3300 1810 3310
rect 1940 3300 2060 3310
rect 2190 3300 2310 3310
rect 2440 3300 2560 3310
rect 2690 3300 2810 3310
rect 2940 3300 3060 3310
rect 3190 3300 3310 3310
rect 3440 3300 3560 3310
rect 3690 3300 3810 3310
rect 3940 3300 4000 3310
rect 0 3295 200 3300
rect 0 3260 75 3295
rect 175 3260 200 3295
rect 0 3240 200 3260
rect 0 3205 75 3240
rect 175 3205 200 3240
rect 0 3200 200 3205
rect 300 3295 450 3300
rect 300 3260 325 3295
rect 425 3260 450 3295
rect 300 3240 450 3260
rect 300 3205 325 3240
rect 425 3205 450 3240
rect 300 3200 450 3205
rect 550 3295 700 3300
rect 550 3260 575 3295
rect 675 3260 700 3295
rect 550 3240 700 3260
rect 550 3205 575 3240
rect 675 3205 700 3240
rect 550 3200 700 3205
rect 800 3295 1200 3300
rect 800 3260 825 3295
rect 925 3260 1075 3295
rect 1175 3260 1200 3295
rect 800 3240 1200 3260
rect 800 3205 825 3240
rect 925 3205 1075 3240
rect 1175 3205 1200 3240
rect 800 3200 1200 3205
rect 1300 3295 1450 3300
rect 1300 3260 1325 3295
rect 1425 3260 1450 3295
rect 1300 3240 1450 3260
rect 1300 3205 1325 3240
rect 1425 3205 1450 3240
rect 1300 3200 1450 3205
rect 1550 3295 1700 3300
rect 1550 3260 1575 3295
rect 1675 3260 1700 3295
rect 1550 3240 1700 3260
rect 1550 3205 1575 3240
rect 1675 3205 1700 3240
rect 1550 3200 1700 3205
rect 1800 3295 2200 3300
rect 1800 3260 1825 3295
rect 1925 3260 2075 3295
rect 2175 3260 2200 3295
rect 1800 3240 2200 3260
rect 1800 3205 1825 3240
rect 1925 3205 2075 3240
rect 2175 3205 2200 3240
rect 1800 3200 2200 3205
rect 2300 3295 2450 3300
rect 2300 3260 2325 3295
rect 2425 3260 2450 3295
rect 2300 3240 2450 3260
rect 2300 3205 2325 3240
rect 2425 3205 2450 3240
rect 2300 3200 2450 3205
rect 2550 3295 2700 3300
rect 2550 3260 2575 3295
rect 2675 3260 2700 3295
rect 2550 3240 2700 3260
rect 2550 3205 2575 3240
rect 2675 3205 2700 3240
rect 2550 3200 2700 3205
rect 2800 3295 3200 3300
rect 2800 3260 2825 3295
rect 2925 3260 3075 3295
rect 3175 3260 3200 3295
rect 2800 3240 3200 3260
rect 2800 3205 2825 3240
rect 2925 3205 3075 3240
rect 3175 3205 3200 3240
rect 2800 3200 3200 3205
rect 3300 3295 3450 3300
rect 3300 3260 3325 3295
rect 3425 3260 3450 3295
rect 3300 3240 3450 3260
rect 3300 3205 3325 3240
rect 3425 3205 3450 3240
rect 3300 3200 3450 3205
rect 3550 3295 3700 3300
rect 3550 3260 3575 3295
rect 3675 3260 3700 3295
rect 3550 3240 3700 3260
rect 3550 3205 3575 3240
rect 3675 3205 3700 3240
rect 3550 3200 3700 3205
rect 3800 3295 4000 3300
rect 3800 3260 3825 3295
rect 3925 3260 4000 3295
rect 3800 3240 4000 3260
rect 3800 3205 3825 3240
rect 3925 3205 4000 3240
rect 3800 3200 4000 3205
rect 0 3190 60 3200
rect 190 3190 310 3200
rect 440 3190 560 3200
rect 690 3190 810 3200
rect 940 3190 1060 3200
rect 1190 3190 1310 3200
rect 1440 3190 1560 3200
rect 1690 3190 1810 3200
rect 1940 3190 2060 3200
rect 2190 3190 2310 3200
rect 2440 3190 2560 3200
rect 2690 3190 2810 3200
rect 2940 3190 3060 3200
rect 3190 3190 3310 3200
rect 3440 3190 3560 3200
rect 3690 3190 3810 3200
rect 3940 3190 4000 3200
rect 0 3175 50 3190
rect 0 3075 10 3175
rect 45 3075 50 3175
rect 0 3060 50 3075
rect 200 3175 300 3190
rect 200 3075 205 3175
rect 240 3075 260 3175
rect 295 3075 300 3175
rect 200 3060 300 3075
rect 450 3175 550 3190
rect 450 3075 455 3175
rect 490 3075 510 3175
rect 545 3075 550 3175
rect 450 3060 550 3075
rect 700 3175 800 3190
rect 700 3075 705 3175
rect 740 3075 760 3175
rect 795 3075 800 3175
rect 700 3060 800 3075
rect 950 3175 1050 3190
rect 950 3075 955 3175
rect 990 3075 1010 3175
rect 1045 3075 1050 3175
rect 950 3060 1050 3075
rect 1200 3175 1300 3190
rect 1200 3075 1205 3175
rect 1240 3075 1260 3175
rect 1295 3075 1300 3175
rect 1200 3060 1300 3075
rect 1450 3175 1550 3190
rect 1450 3075 1455 3175
rect 1490 3075 1510 3175
rect 1545 3075 1550 3175
rect 1450 3060 1550 3075
rect 1700 3175 1800 3190
rect 1700 3075 1705 3175
rect 1740 3075 1760 3175
rect 1795 3075 1800 3175
rect 1700 3060 1800 3075
rect 1950 3175 2050 3190
rect 1950 3075 1955 3175
rect 1990 3075 2010 3175
rect 2045 3075 2050 3175
rect 1950 3060 2050 3075
rect 2200 3175 2300 3190
rect 2200 3075 2205 3175
rect 2240 3075 2260 3175
rect 2295 3075 2300 3175
rect 2200 3060 2300 3075
rect 2450 3175 2550 3190
rect 2450 3075 2455 3175
rect 2490 3075 2510 3175
rect 2545 3075 2550 3175
rect 2450 3060 2550 3075
rect 2700 3175 2800 3190
rect 2700 3075 2705 3175
rect 2740 3075 2760 3175
rect 2795 3075 2800 3175
rect 2700 3060 2800 3075
rect 2950 3175 3050 3190
rect 2950 3075 2955 3175
rect 2990 3075 3010 3175
rect 3045 3075 3050 3175
rect 2950 3060 3050 3075
rect 3200 3175 3300 3190
rect 3200 3075 3205 3175
rect 3240 3075 3260 3175
rect 3295 3075 3300 3175
rect 3200 3060 3300 3075
rect 3450 3175 3550 3190
rect 3450 3075 3455 3175
rect 3490 3075 3510 3175
rect 3545 3075 3550 3175
rect 3450 3060 3550 3075
rect 3700 3175 3800 3190
rect 3700 3075 3705 3175
rect 3740 3075 3760 3175
rect 3795 3075 3800 3175
rect 3700 3060 3800 3075
rect 3950 3175 4000 3190
rect 3950 3075 3955 3175
rect 3990 3075 4000 3175
rect 3950 3060 4000 3075
rect 0 3050 60 3060
rect 190 3050 310 3060
rect 440 3050 560 3060
rect 690 3050 810 3060
rect 940 3050 1060 3060
rect 1190 3050 1310 3060
rect 1440 3050 1560 3060
rect 1690 3050 1810 3060
rect 1940 3050 2060 3060
rect 2190 3050 2310 3060
rect 2440 3050 2560 3060
rect 2690 3050 2810 3060
rect 2940 3050 3060 3060
rect 3190 3050 3310 3060
rect 3440 3050 3560 3060
rect 3690 3050 3810 3060
rect 3940 3050 4000 3060
rect 0 3045 450 3050
rect 0 3010 75 3045
rect 175 3010 325 3045
rect 425 3010 450 3045
rect 0 2990 450 3010
rect 0 2955 75 2990
rect 175 2955 325 2990
rect 425 2955 450 2990
rect 0 2950 450 2955
rect 550 3045 1450 3050
rect 550 3010 575 3045
rect 675 3010 825 3045
rect 925 3010 1075 3045
rect 1175 3010 1325 3045
rect 1425 3010 1450 3045
rect 550 2990 1450 3010
rect 550 2955 575 2990
rect 675 2955 825 2990
rect 925 2955 1075 2990
rect 1175 2955 1325 2990
rect 1425 2955 1450 2990
rect 550 2950 1450 2955
rect 1550 3045 2450 3050
rect 1550 3010 1575 3045
rect 1675 3010 1825 3045
rect 1925 3010 2075 3045
rect 2175 3010 2325 3045
rect 2425 3010 2450 3045
rect 1550 2990 2450 3010
rect 1550 2955 1575 2990
rect 1675 2955 1825 2990
rect 1925 2955 2075 2990
rect 2175 2955 2325 2990
rect 2425 2955 2450 2990
rect 1550 2950 2450 2955
rect 2550 3045 3450 3050
rect 2550 3010 2575 3045
rect 2675 3010 2825 3045
rect 2925 3010 3075 3045
rect 3175 3010 3325 3045
rect 3425 3010 3450 3045
rect 2550 2990 3450 3010
rect 2550 2955 2575 2990
rect 2675 2955 2825 2990
rect 2925 2955 3075 2990
rect 3175 2955 3325 2990
rect 3425 2955 3450 2990
rect 2550 2950 3450 2955
rect 3550 3045 4000 3050
rect 3550 3010 3575 3045
rect 3675 3010 3825 3045
rect 3925 3010 4000 3045
rect 3550 2990 4000 3010
rect 3550 2955 3575 2990
rect 3675 2955 3825 2990
rect 3925 2955 4000 2990
rect 3550 2950 4000 2955
rect 0 2940 60 2950
rect 190 2940 310 2950
rect 440 2940 560 2950
rect 690 2940 810 2950
rect 940 2940 1060 2950
rect 1190 2940 1310 2950
rect 1440 2940 1560 2950
rect 1690 2940 1810 2950
rect 1940 2940 2060 2950
rect 2190 2940 2310 2950
rect 2440 2940 2560 2950
rect 2690 2940 2810 2950
rect 2940 2940 3060 2950
rect 3190 2940 3310 2950
rect 3440 2940 3560 2950
rect 3690 2940 3810 2950
rect 3940 2940 4000 2950
rect 0 2925 50 2940
rect 0 2825 10 2925
rect 45 2825 50 2925
rect 0 2810 50 2825
rect 200 2925 300 2940
rect 200 2825 205 2925
rect 240 2825 260 2925
rect 295 2825 300 2925
rect 200 2810 300 2825
rect 450 2925 550 2940
rect 450 2825 455 2925
rect 490 2825 510 2925
rect 545 2825 550 2925
rect 450 2810 550 2825
rect 700 2925 800 2940
rect 700 2825 705 2925
rect 740 2825 760 2925
rect 795 2825 800 2925
rect 700 2810 800 2825
rect 950 2925 1050 2940
rect 950 2825 955 2925
rect 990 2825 1010 2925
rect 1045 2825 1050 2925
rect 950 2810 1050 2825
rect 1200 2925 1300 2940
rect 1200 2825 1205 2925
rect 1240 2825 1260 2925
rect 1295 2825 1300 2925
rect 1200 2810 1300 2825
rect 1450 2925 1550 2940
rect 1450 2825 1455 2925
rect 1490 2825 1510 2925
rect 1545 2825 1550 2925
rect 1450 2810 1550 2825
rect 1700 2925 1800 2940
rect 1700 2825 1705 2925
rect 1740 2825 1760 2925
rect 1795 2825 1800 2925
rect 1700 2810 1800 2825
rect 1950 2925 2050 2940
rect 1950 2825 1955 2925
rect 1990 2825 2010 2925
rect 2045 2825 2050 2925
rect 1950 2810 2050 2825
rect 2200 2925 2300 2940
rect 2200 2825 2205 2925
rect 2240 2825 2260 2925
rect 2295 2825 2300 2925
rect 2200 2810 2300 2825
rect 2450 2925 2550 2940
rect 2450 2825 2455 2925
rect 2490 2825 2510 2925
rect 2545 2825 2550 2925
rect 2450 2810 2550 2825
rect 2700 2925 2800 2940
rect 2700 2825 2705 2925
rect 2740 2825 2760 2925
rect 2795 2825 2800 2925
rect 2700 2810 2800 2825
rect 2950 2925 3050 2940
rect 2950 2825 2955 2925
rect 2990 2825 3010 2925
rect 3045 2825 3050 2925
rect 2950 2810 3050 2825
rect 3200 2925 3300 2940
rect 3200 2825 3205 2925
rect 3240 2825 3260 2925
rect 3295 2825 3300 2925
rect 3200 2810 3300 2825
rect 3450 2925 3550 2940
rect 3450 2825 3455 2925
rect 3490 2825 3510 2925
rect 3545 2825 3550 2925
rect 3450 2810 3550 2825
rect 3700 2925 3800 2940
rect 3700 2825 3705 2925
rect 3740 2825 3760 2925
rect 3795 2825 3800 2925
rect 3700 2810 3800 2825
rect 3950 2925 4000 2940
rect 3950 2825 3955 2925
rect 3990 2825 4000 2925
rect 3950 2810 4000 2825
rect 0 2800 60 2810
rect 190 2800 310 2810
rect 440 2800 560 2810
rect 690 2800 810 2810
rect 940 2800 1060 2810
rect 1190 2800 1310 2810
rect 1440 2800 1560 2810
rect 1690 2800 1810 2810
rect 1940 2800 2060 2810
rect 2190 2800 2310 2810
rect 2440 2800 2560 2810
rect 2690 2800 2810 2810
rect 2940 2800 3060 2810
rect 3190 2800 3310 2810
rect 3440 2800 3560 2810
rect 3690 2800 3810 2810
rect 3940 2800 4000 2810
rect 0 2795 200 2800
rect 0 2760 75 2795
rect 175 2760 200 2795
rect 0 2740 200 2760
rect 0 2705 75 2740
rect 175 2705 200 2740
rect 0 2700 200 2705
rect 300 2795 450 2800
rect 300 2760 325 2795
rect 425 2760 450 2795
rect 300 2740 450 2760
rect 300 2705 325 2740
rect 425 2705 450 2740
rect 300 2700 450 2705
rect 550 2795 700 2800
rect 550 2760 575 2795
rect 675 2760 700 2795
rect 550 2740 700 2760
rect 550 2705 575 2740
rect 675 2705 700 2740
rect 550 2700 700 2705
rect 800 2795 1200 2800
rect 800 2760 825 2795
rect 925 2760 1075 2795
rect 1175 2760 1200 2795
rect 800 2740 1200 2760
rect 800 2705 825 2740
rect 925 2705 1075 2740
rect 1175 2705 1200 2740
rect 800 2700 1200 2705
rect 1300 2795 1450 2800
rect 1300 2760 1325 2795
rect 1425 2760 1450 2795
rect 1300 2740 1450 2760
rect 1300 2705 1325 2740
rect 1425 2705 1450 2740
rect 1300 2700 1450 2705
rect 1550 2795 1700 2800
rect 1550 2760 1575 2795
rect 1675 2760 1700 2795
rect 1550 2740 1700 2760
rect 1550 2705 1575 2740
rect 1675 2705 1700 2740
rect 1550 2700 1700 2705
rect 1800 2795 2200 2800
rect 1800 2760 1825 2795
rect 1925 2760 2075 2795
rect 2175 2760 2200 2795
rect 1800 2740 2200 2760
rect 1800 2705 1825 2740
rect 1925 2705 2075 2740
rect 2175 2705 2200 2740
rect 1800 2700 2200 2705
rect 2300 2795 2450 2800
rect 2300 2760 2325 2795
rect 2425 2760 2450 2795
rect 2300 2740 2450 2760
rect 2300 2705 2325 2740
rect 2425 2705 2450 2740
rect 2300 2700 2450 2705
rect 2550 2795 2700 2800
rect 2550 2760 2575 2795
rect 2675 2760 2700 2795
rect 2550 2740 2700 2760
rect 2550 2705 2575 2740
rect 2675 2705 2700 2740
rect 2550 2700 2700 2705
rect 2800 2795 3200 2800
rect 2800 2760 2825 2795
rect 2925 2760 3075 2795
rect 3175 2760 3200 2795
rect 2800 2740 3200 2760
rect 2800 2705 2825 2740
rect 2925 2705 3075 2740
rect 3175 2705 3200 2740
rect 2800 2700 3200 2705
rect 3300 2795 3450 2800
rect 3300 2760 3325 2795
rect 3425 2760 3450 2795
rect 3300 2740 3450 2760
rect 3300 2705 3325 2740
rect 3425 2705 3450 2740
rect 3300 2700 3450 2705
rect 3550 2795 3700 2800
rect 3550 2760 3575 2795
rect 3675 2760 3700 2795
rect 3550 2740 3700 2760
rect 3550 2705 3575 2740
rect 3675 2705 3700 2740
rect 3550 2700 3700 2705
rect 3800 2795 4000 2800
rect 3800 2760 3825 2795
rect 3925 2760 4000 2795
rect 3800 2740 4000 2760
rect 3800 2705 3825 2740
rect 3925 2705 4000 2740
rect 3800 2700 4000 2705
rect 0 2690 60 2700
rect 190 2690 310 2700
rect 440 2690 560 2700
rect 690 2690 810 2700
rect 940 2690 1060 2700
rect 1190 2690 1310 2700
rect 1440 2690 1560 2700
rect 1690 2690 1810 2700
rect 1940 2690 2060 2700
rect 2190 2690 2310 2700
rect 2440 2690 2560 2700
rect 2690 2690 2810 2700
rect 2940 2690 3060 2700
rect 3190 2690 3310 2700
rect 3440 2690 3560 2700
rect 3690 2690 3810 2700
rect 3940 2690 4000 2700
rect 0 2675 50 2690
rect 0 2575 10 2675
rect 45 2575 50 2675
rect 0 2560 50 2575
rect 200 2675 300 2690
rect 200 2575 205 2675
rect 240 2575 260 2675
rect 295 2575 300 2675
rect 200 2560 300 2575
rect 450 2675 550 2690
rect 450 2575 455 2675
rect 490 2575 510 2675
rect 545 2575 550 2675
rect 450 2560 550 2575
rect 700 2675 800 2690
rect 700 2575 705 2675
rect 740 2575 760 2675
rect 795 2575 800 2675
rect 700 2560 800 2575
rect 950 2675 1050 2690
rect 950 2575 955 2675
rect 990 2575 1010 2675
rect 1045 2575 1050 2675
rect 950 2560 1050 2575
rect 1200 2675 1300 2690
rect 1200 2575 1205 2675
rect 1240 2575 1260 2675
rect 1295 2575 1300 2675
rect 1200 2560 1300 2575
rect 1450 2675 1550 2690
rect 1450 2575 1455 2675
rect 1490 2575 1510 2675
rect 1545 2575 1550 2675
rect 1450 2560 1550 2575
rect 1700 2675 1800 2690
rect 1700 2575 1705 2675
rect 1740 2575 1760 2675
rect 1795 2575 1800 2675
rect 1700 2560 1800 2575
rect 1950 2675 2050 2690
rect 1950 2575 1955 2675
rect 1990 2575 2010 2675
rect 2045 2575 2050 2675
rect 1950 2560 2050 2575
rect 2200 2675 2300 2690
rect 2200 2575 2205 2675
rect 2240 2575 2260 2675
rect 2295 2575 2300 2675
rect 2200 2560 2300 2575
rect 2450 2675 2550 2690
rect 2450 2575 2455 2675
rect 2490 2575 2510 2675
rect 2545 2575 2550 2675
rect 2450 2560 2550 2575
rect 2700 2675 2800 2690
rect 2700 2575 2705 2675
rect 2740 2575 2760 2675
rect 2795 2575 2800 2675
rect 2700 2560 2800 2575
rect 2950 2675 3050 2690
rect 2950 2575 2955 2675
rect 2990 2575 3010 2675
rect 3045 2575 3050 2675
rect 2950 2560 3050 2575
rect 3200 2675 3300 2690
rect 3200 2575 3205 2675
rect 3240 2575 3260 2675
rect 3295 2575 3300 2675
rect 3200 2560 3300 2575
rect 3450 2675 3550 2690
rect 3450 2575 3455 2675
rect 3490 2575 3510 2675
rect 3545 2575 3550 2675
rect 3450 2560 3550 2575
rect 3700 2675 3800 2690
rect 3700 2575 3705 2675
rect 3740 2575 3760 2675
rect 3795 2575 3800 2675
rect 3700 2560 3800 2575
rect 3950 2675 4000 2690
rect 3950 2575 3955 2675
rect 3990 2575 4000 2675
rect 3950 2560 4000 2575
rect 0 2550 60 2560
rect 190 2550 310 2560
rect 440 2550 560 2560
rect 690 2550 810 2560
rect 940 2550 1060 2560
rect 1190 2550 1310 2560
rect 1440 2550 1560 2560
rect 1690 2550 1810 2560
rect 1940 2550 2060 2560
rect 2190 2550 2310 2560
rect 2440 2550 2560 2560
rect 2690 2550 2810 2560
rect 2940 2550 3060 2560
rect 3190 2550 3310 2560
rect 3440 2550 3560 2560
rect 3690 2550 3810 2560
rect 3940 2550 4000 2560
rect 0 2545 200 2550
rect 0 2510 75 2545
rect 175 2510 200 2545
rect 0 2490 200 2510
rect 0 2455 75 2490
rect 175 2455 200 2490
rect 0 2450 200 2455
rect 300 2545 450 2550
rect 300 2510 325 2545
rect 425 2510 450 2545
rect 300 2490 450 2510
rect 300 2455 325 2490
rect 425 2455 450 2490
rect 300 2450 450 2455
rect 550 2545 700 2550
rect 550 2510 575 2545
rect 675 2510 700 2545
rect 550 2490 700 2510
rect 550 2455 575 2490
rect 675 2455 700 2490
rect 550 2450 700 2455
rect 800 2545 950 2550
rect 800 2510 825 2545
rect 925 2510 950 2545
rect 800 2490 950 2510
rect 800 2455 825 2490
rect 925 2455 950 2490
rect 800 2450 950 2455
rect 1050 2545 1200 2550
rect 1050 2510 1075 2545
rect 1175 2510 1200 2545
rect 1050 2490 1200 2510
rect 1050 2455 1075 2490
rect 1175 2455 1200 2490
rect 1050 2450 1200 2455
rect 1300 2545 1450 2550
rect 1300 2510 1325 2545
rect 1425 2510 1450 2545
rect 1300 2490 1450 2510
rect 1300 2455 1325 2490
rect 1425 2455 1450 2490
rect 1300 2450 1450 2455
rect 1550 2545 1700 2550
rect 1550 2510 1575 2545
rect 1675 2510 1700 2545
rect 1550 2490 1700 2510
rect 1550 2455 1575 2490
rect 1675 2455 1700 2490
rect 1550 2450 1700 2455
rect 1800 2545 2200 2550
rect 1800 2510 1825 2545
rect 1925 2510 2075 2545
rect 2175 2510 2200 2545
rect 1800 2490 2200 2510
rect 1800 2455 1825 2490
rect 1925 2455 2075 2490
rect 2175 2455 2200 2490
rect 1800 2450 2200 2455
rect 2300 2545 2450 2550
rect 2300 2510 2325 2545
rect 2425 2510 2450 2545
rect 2300 2490 2450 2510
rect 2300 2455 2325 2490
rect 2425 2455 2450 2490
rect 2300 2450 2450 2455
rect 2550 2545 2700 2550
rect 2550 2510 2575 2545
rect 2675 2510 2700 2545
rect 2550 2490 2700 2510
rect 2550 2455 2575 2490
rect 2675 2455 2700 2490
rect 2550 2450 2700 2455
rect 2800 2545 2950 2550
rect 2800 2510 2825 2545
rect 2925 2510 2950 2545
rect 2800 2490 2950 2510
rect 2800 2455 2825 2490
rect 2925 2455 2950 2490
rect 2800 2450 2950 2455
rect 3050 2545 3200 2550
rect 3050 2510 3075 2545
rect 3175 2510 3200 2545
rect 3050 2490 3200 2510
rect 3050 2455 3075 2490
rect 3175 2455 3200 2490
rect 3050 2450 3200 2455
rect 3300 2545 3450 2550
rect 3300 2510 3325 2545
rect 3425 2510 3450 2545
rect 3300 2490 3450 2510
rect 3300 2455 3325 2490
rect 3425 2455 3450 2490
rect 3300 2450 3450 2455
rect 3550 2545 3700 2550
rect 3550 2510 3575 2545
rect 3675 2510 3700 2545
rect 3550 2490 3700 2510
rect 3550 2455 3575 2490
rect 3675 2455 3700 2490
rect 3550 2450 3700 2455
rect 3800 2545 4000 2550
rect 3800 2510 3825 2545
rect 3925 2510 4000 2545
rect 3800 2490 4000 2510
rect 3800 2455 3825 2490
rect 3925 2455 4000 2490
rect 3800 2450 4000 2455
rect 0 2440 60 2450
rect 190 2440 310 2450
rect 440 2440 560 2450
rect 690 2440 810 2450
rect 940 2440 1060 2450
rect 1190 2440 1310 2450
rect 1440 2440 1560 2450
rect 1690 2440 1810 2450
rect 1940 2440 2060 2450
rect 2190 2440 2310 2450
rect 2440 2440 2560 2450
rect 2690 2440 2810 2450
rect 2940 2440 3060 2450
rect 3190 2440 3310 2450
rect 3440 2440 3560 2450
rect 3690 2440 3810 2450
rect 3940 2440 4000 2450
rect 0 2425 50 2440
rect 0 2325 10 2425
rect 45 2325 50 2425
rect 0 2310 50 2325
rect 200 2425 300 2440
rect 200 2325 205 2425
rect 240 2325 260 2425
rect 295 2325 300 2425
rect 200 2310 300 2325
rect 450 2425 550 2440
rect 450 2325 455 2425
rect 490 2325 510 2425
rect 545 2325 550 2425
rect 450 2310 550 2325
rect 700 2425 800 2440
rect 700 2325 705 2425
rect 740 2325 760 2425
rect 795 2325 800 2425
rect 700 2310 800 2325
rect 950 2425 1050 2440
rect 950 2325 955 2425
rect 990 2325 1010 2425
rect 1045 2325 1050 2425
rect 950 2310 1050 2325
rect 1200 2425 1300 2440
rect 1200 2325 1205 2425
rect 1240 2325 1260 2425
rect 1295 2325 1300 2425
rect 1200 2310 1300 2325
rect 1450 2425 1550 2440
rect 1450 2325 1455 2425
rect 1490 2325 1510 2425
rect 1545 2325 1550 2425
rect 1450 2310 1550 2325
rect 1700 2425 1800 2440
rect 1700 2325 1705 2425
rect 1740 2325 1760 2425
rect 1795 2325 1800 2425
rect 1700 2310 1800 2325
rect 1950 2425 2050 2440
rect 1950 2325 1955 2425
rect 1990 2325 2010 2425
rect 2045 2325 2050 2425
rect 1950 2310 2050 2325
rect 2200 2425 2300 2440
rect 2200 2325 2205 2425
rect 2240 2325 2260 2425
rect 2295 2325 2300 2425
rect 2200 2310 2300 2325
rect 2450 2425 2550 2440
rect 2450 2325 2455 2425
rect 2490 2325 2510 2425
rect 2545 2325 2550 2425
rect 2450 2310 2550 2325
rect 2700 2425 2800 2440
rect 2700 2325 2705 2425
rect 2740 2325 2760 2425
rect 2795 2325 2800 2425
rect 2700 2310 2800 2325
rect 2950 2425 3050 2440
rect 2950 2325 2955 2425
rect 2990 2325 3010 2425
rect 3045 2325 3050 2425
rect 2950 2310 3050 2325
rect 3200 2425 3300 2440
rect 3200 2325 3205 2425
rect 3240 2325 3260 2425
rect 3295 2325 3300 2425
rect 3200 2310 3300 2325
rect 3450 2425 3550 2440
rect 3450 2325 3455 2425
rect 3490 2325 3510 2425
rect 3545 2325 3550 2425
rect 3450 2310 3550 2325
rect 3700 2425 3800 2440
rect 3700 2325 3705 2425
rect 3740 2325 3760 2425
rect 3795 2325 3800 2425
rect 3700 2310 3800 2325
rect 3950 2425 4000 2440
rect 3950 2325 3955 2425
rect 3990 2325 4000 2425
rect 3950 2310 4000 2325
rect 0 2300 60 2310
rect 190 2300 310 2310
rect 440 2300 560 2310
rect 690 2300 810 2310
rect 940 2300 1060 2310
rect 1190 2300 1310 2310
rect 1440 2300 1560 2310
rect 1690 2300 1810 2310
rect 1940 2300 2060 2310
rect 2190 2300 2310 2310
rect 2440 2300 2560 2310
rect 2690 2300 2810 2310
rect 2940 2300 3060 2310
rect 3190 2300 3310 2310
rect 3440 2300 3560 2310
rect 3690 2300 3810 2310
rect 3940 2300 4000 2310
rect 0 2295 200 2300
rect 0 2260 75 2295
rect 175 2260 200 2295
rect 0 2240 200 2260
rect 0 2205 75 2240
rect 175 2205 200 2240
rect 0 2200 200 2205
rect 300 2295 450 2300
rect 300 2260 325 2295
rect 425 2260 450 2295
rect 300 2240 450 2260
rect 300 2205 325 2240
rect 425 2205 450 2240
rect 300 2200 450 2205
rect 550 2295 700 2300
rect 550 2260 575 2295
rect 675 2260 700 2295
rect 550 2240 700 2260
rect 550 2205 575 2240
rect 675 2205 700 2240
rect 550 2200 700 2205
rect 800 2295 1200 2300
rect 800 2260 825 2295
rect 925 2260 1075 2295
rect 1175 2260 1200 2295
rect 800 2240 1200 2260
rect 800 2205 825 2240
rect 925 2205 1075 2240
rect 1175 2205 1200 2240
rect 800 2200 1200 2205
rect 1300 2295 1450 2300
rect 1300 2260 1325 2295
rect 1425 2260 1450 2295
rect 1300 2240 1450 2260
rect 1300 2205 1325 2240
rect 1425 2205 1450 2240
rect 1300 2200 1450 2205
rect 1550 2295 1700 2300
rect 1550 2260 1575 2295
rect 1675 2260 1700 2295
rect 1550 2240 1700 2260
rect 1550 2205 1575 2240
rect 1675 2205 1700 2240
rect 1550 2200 1700 2205
rect 1800 2295 2200 2300
rect 1800 2260 1825 2295
rect 1925 2260 2075 2295
rect 2175 2260 2200 2295
rect 1800 2240 2200 2260
rect 1800 2205 1825 2240
rect 1925 2205 2075 2240
rect 2175 2205 2200 2240
rect 1800 2200 2200 2205
rect 2300 2295 2450 2300
rect 2300 2260 2325 2295
rect 2425 2260 2450 2295
rect 2300 2240 2450 2260
rect 2300 2205 2325 2240
rect 2425 2205 2450 2240
rect 2300 2200 2450 2205
rect 2550 2295 2700 2300
rect 2550 2260 2575 2295
rect 2675 2260 2700 2295
rect 2550 2240 2700 2260
rect 2550 2205 2575 2240
rect 2675 2205 2700 2240
rect 2550 2200 2700 2205
rect 2800 2295 3200 2300
rect 2800 2260 2825 2295
rect 2925 2260 3075 2295
rect 3175 2260 3200 2295
rect 2800 2240 3200 2260
rect 2800 2205 2825 2240
rect 2925 2205 3075 2240
rect 3175 2205 3200 2240
rect 2800 2200 3200 2205
rect 3300 2295 3450 2300
rect 3300 2260 3325 2295
rect 3425 2260 3450 2295
rect 3300 2240 3450 2260
rect 3300 2205 3325 2240
rect 3425 2205 3450 2240
rect 3300 2200 3450 2205
rect 3550 2295 3700 2300
rect 3550 2260 3575 2295
rect 3675 2260 3700 2295
rect 3550 2240 3700 2260
rect 3550 2205 3575 2240
rect 3675 2205 3700 2240
rect 3550 2200 3700 2205
rect 3800 2295 4000 2300
rect 3800 2260 3825 2295
rect 3925 2260 4000 2295
rect 3800 2240 4000 2260
rect 3800 2205 3825 2240
rect 3925 2205 4000 2240
rect 3800 2200 4000 2205
rect 0 2190 60 2200
rect 190 2190 310 2200
rect 440 2190 560 2200
rect 690 2190 810 2200
rect 940 2190 1060 2200
rect 1190 2190 1310 2200
rect 1440 2190 1560 2200
rect 1690 2190 1810 2200
rect 1940 2190 2060 2200
rect 2190 2190 2310 2200
rect 2440 2190 2560 2200
rect 2690 2190 2810 2200
rect 2940 2190 3060 2200
rect 3190 2190 3310 2200
rect 3440 2190 3560 2200
rect 3690 2190 3810 2200
rect 3940 2190 4000 2200
rect 0 2175 50 2190
rect 0 2075 10 2175
rect 45 2075 50 2175
rect 0 2060 50 2075
rect 200 2175 300 2190
rect 200 2075 205 2175
rect 240 2075 260 2175
rect 295 2075 300 2175
rect 200 2060 300 2075
rect 450 2175 550 2190
rect 450 2075 455 2175
rect 490 2075 510 2175
rect 545 2075 550 2175
rect 450 2060 550 2075
rect 700 2175 800 2190
rect 700 2075 705 2175
rect 740 2075 760 2175
rect 795 2075 800 2175
rect 700 2060 800 2075
rect 950 2175 1050 2190
rect 950 2075 955 2175
rect 990 2075 1010 2175
rect 1045 2075 1050 2175
rect 950 2060 1050 2075
rect 1200 2175 1300 2190
rect 1200 2075 1205 2175
rect 1240 2075 1260 2175
rect 1295 2075 1300 2175
rect 1200 2060 1300 2075
rect 1450 2175 1550 2190
rect 1450 2075 1455 2175
rect 1490 2075 1510 2175
rect 1545 2075 1550 2175
rect 1450 2060 1550 2075
rect 1700 2175 1800 2190
rect 1700 2075 1705 2175
rect 1740 2075 1760 2175
rect 1795 2075 1800 2175
rect 1700 2060 1800 2075
rect 1950 2175 2050 2190
rect 1950 2075 1955 2175
rect 1990 2075 2010 2175
rect 2045 2075 2050 2175
rect 1950 2060 2050 2075
rect 2200 2175 2300 2190
rect 2200 2075 2205 2175
rect 2240 2075 2260 2175
rect 2295 2075 2300 2175
rect 2200 2060 2300 2075
rect 2450 2175 2550 2190
rect 2450 2075 2455 2175
rect 2490 2075 2510 2175
rect 2545 2075 2550 2175
rect 2450 2060 2550 2075
rect 2700 2175 2800 2190
rect 2700 2075 2705 2175
rect 2740 2075 2760 2175
rect 2795 2075 2800 2175
rect 2700 2060 2800 2075
rect 2950 2175 3050 2190
rect 2950 2075 2955 2175
rect 2990 2075 3010 2175
rect 3045 2075 3050 2175
rect 2950 2060 3050 2075
rect 3200 2175 3300 2190
rect 3200 2075 3205 2175
rect 3240 2075 3260 2175
rect 3295 2075 3300 2175
rect 3200 2060 3300 2075
rect 3450 2175 3550 2190
rect 3450 2075 3455 2175
rect 3490 2075 3510 2175
rect 3545 2075 3550 2175
rect 3450 2060 3550 2075
rect 3700 2175 3800 2190
rect 3700 2075 3705 2175
rect 3740 2075 3760 2175
rect 3795 2075 3800 2175
rect 3700 2060 3800 2075
rect 3950 2175 4000 2190
rect 3950 2075 3955 2175
rect 3990 2075 4000 2175
rect 3950 2060 4000 2075
rect 0 2050 60 2060
rect 190 2050 310 2060
rect 440 2050 560 2060
rect 690 2050 810 2060
rect 940 2050 1060 2060
rect 1190 2050 1310 2060
rect 1440 2050 1560 2060
rect 1690 2050 1810 2060
rect 1940 2050 2060 2060
rect 2190 2050 2310 2060
rect 2440 2050 2560 2060
rect 2690 2050 2810 2060
rect 2940 2050 3060 2060
rect 3190 2050 3310 2060
rect 3440 2050 3560 2060
rect 3690 2050 3810 2060
rect 3940 2050 4000 2060
rect 0 2045 4000 2050
rect 0 2010 75 2045
rect 175 2010 325 2045
rect 425 2010 575 2045
rect 675 2010 825 2045
rect 925 2010 1075 2045
rect 1175 2010 1325 2045
rect 1425 2010 1575 2045
rect 1675 2010 1825 2045
rect 1925 2010 2075 2045
rect 2175 2010 2325 2045
rect 2425 2010 2575 2045
rect 2675 2010 2825 2045
rect 2925 2010 3075 2045
rect 3175 2010 3325 2045
rect 3425 2010 3575 2045
rect 3675 2010 3825 2045
rect 3925 2010 4000 2045
rect 0 1990 4000 2010
rect 0 1955 75 1990
rect 175 1955 325 1990
rect 425 1955 575 1990
rect 675 1955 825 1990
rect 925 1955 1075 1990
rect 1175 1955 1325 1990
rect 1425 1955 1575 1990
rect 1675 1955 1825 1990
rect 1925 1955 2075 1990
rect 2175 1955 2325 1990
rect 2425 1955 2575 1990
rect 2675 1955 2825 1990
rect 2925 1955 3075 1990
rect 3175 1955 3325 1990
rect 3425 1955 3575 1990
rect 3675 1955 3825 1990
rect 3925 1955 4000 1990
rect 0 1950 4000 1955
rect 0 1940 60 1950
rect 190 1940 310 1950
rect 440 1940 560 1950
rect 690 1940 810 1950
rect 940 1940 1060 1950
rect 1190 1940 1310 1950
rect 1440 1940 1560 1950
rect 1690 1940 1810 1950
rect 1940 1940 2060 1950
rect 2190 1940 2310 1950
rect 2440 1940 2560 1950
rect 2690 1940 2810 1950
rect 2940 1940 3060 1950
rect 3190 1940 3310 1950
rect 3440 1940 3560 1950
rect 3690 1940 3810 1950
rect 3940 1940 4000 1950
rect 0 1925 50 1940
rect 0 1825 10 1925
rect 45 1825 50 1925
rect 0 1810 50 1825
rect 200 1925 300 1940
rect 200 1825 205 1925
rect 240 1825 260 1925
rect 295 1825 300 1925
rect 200 1810 300 1825
rect 450 1925 550 1940
rect 450 1825 455 1925
rect 490 1825 510 1925
rect 545 1825 550 1925
rect 450 1810 550 1825
rect 700 1925 800 1940
rect 700 1825 705 1925
rect 740 1825 760 1925
rect 795 1825 800 1925
rect 700 1810 800 1825
rect 950 1925 1050 1940
rect 950 1825 955 1925
rect 990 1825 1010 1925
rect 1045 1825 1050 1925
rect 950 1810 1050 1825
rect 1200 1925 1300 1940
rect 1200 1825 1205 1925
rect 1240 1825 1260 1925
rect 1295 1825 1300 1925
rect 1200 1810 1300 1825
rect 1450 1925 1550 1940
rect 1450 1825 1455 1925
rect 1490 1825 1510 1925
rect 1545 1825 1550 1925
rect 1450 1810 1550 1825
rect 1700 1925 1800 1940
rect 1700 1825 1705 1925
rect 1740 1825 1760 1925
rect 1795 1825 1800 1925
rect 1700 1810 1800 1825
rect 1950 1925 2050 1940
rect 1950 1825 1955 1925
rect 1990 1825 2010 1925
rect 2045 1825 2050 1925
rect 1950 1810 2050 1825
rect 2200 1925 2300 1940
rect 2200 1825 2205 1925
rect 2240 1825 2260 1925
rect 2295 1825 2300 1925
rect 2200 1810 2300 1825
rect 2450 1925 2550 1940
rect 2450 1825 2455 1925
rect 2490 1825 2510 1925
rect 2545 1825 2550 1925
rect 2450 1810 2550 1825
rect 2700 1925 2800 1940
rect 2700 1825 2705 1925
rect 2740 1825 2760 1925
rect 2795 1825 2800 1925
rect 2700 1810 2800 1825
rect 2950 1925 3050 1940
rect 2950 1825 2955 1925
rect 2990 1825 3010 1925
rect 3045 1825 3050 1925
rect 2950 1810 3050 1825
rect 3200 1925 3300 1940
rect 3200 1825 3205 1925
rect 3240 1825 3260 1925
rect 3295 1825 3300 1925
rect 3200 1810 3300 1825
rect 3450 1925 3550 1940
rect 3450 1825 3455 1925
rect 3490 1825 3510 1925
rect 3545 1825 3550 1925
rect 3450 1810 3550 1825
rect 3700 1925 3800 1940
rect 3700 1825 3705 1925
rect 3740 1825 3760 1925
rect 3795 1825 3800 1925
rect 3700 1810 3800 1825
rect 3950 1925 4000 1940
rect 3950 1825 3955 1925
rect 3990 1825 4000 1925
rect 3950 1810 4000 1825
rect 0 1800 60 1810
rect 190 1800 310 1810
rect 440 1800 560 1810
rect 690 1800 810 1810
rect 940 1800 1060 1810
rect 1190 1800 1310 1810
rect 1440 1800 1560 1810
rect 1690 1800 1810 1810
rect 1940 1800 2060 1810
rect 2190 1800 2310 1810
rect 2440 1800 2560 1810
rect 2690 1800 2810 1810
rect 2940 1800 3060 1810
rect 3190 1800 3310 1810
rect 3440 1800 3560 1810
rect 3690 1800 3810 1810
rect 3940 1800 4000 1810
rect 0 1795 200 1800
rect 0 1760 75 1795
rect 175 1760 200 1795
rect 0 1740 200 1760
rect 0 1705 75 1740
rect 175 1705 200 1740
rect 0 1700 200 1705
rect 300 1795 450 1800
rect 300 1760 325 1795
rect 425 1760 450 1795
rect 300 1740 450 1760
rect 300 1705 325 1740
rect 425 1705 450 1740
rect 300 1700 450 1705
rect 550 1795 700 1800
rect 550 1760 575 1795
rect 675 1760 700 1795
rect 550 1740 700 1760
rect 550 1705 575 1740
rect 675 1705 700 1740
rect 550 1700 700 1705
rect 800 1795 1200 1800
rect 800 1760 825 1795
rect 925 1760 1075 1795
rect 1175 1760 1200 1795
rect 800 1740 1200 1760
rect 800 1705 825 1740
rect 925 1705 1075 1740
rect 1175 1705 1200 1740
rect 800 1700 1200 1705
rect 1300 1795 1450 1800
rect 1300 1760 1325 1795
rect 1425 1760 1450 1795
rect 1300 1740 1450 1760
rect 1300 1705 1325 1740
rect 1425 1705 1450 1740
rect 1300 1700 1450 1705
rect 1550 1795 1700 1800
rect 1550 1760 1575 1795
rect 1675 1760 1700 1795
rect 1550 1740 1700 1760
rect 1550 1705 1575 1740
rect 1675 1705 1700 1740
rect 1550 1700 1700 1705
rect 1800 1795 2200 1800
rect 1800 1760 1825 1795
rect 1925 1760 2075 1795
rect 2175 1760 2200 1795
rect 1800 1740 2200 1760
rect 1800 1705 1825 1740
rect 1925 1705 2075 1740
rect 2175 1705 2200 1740
rect 1800 1700 2200 1705
rect 2300 1795 2450 1800
rect 2300 1760 2325 1795
rect 2425 1760 2450 1795
rect 2300 1740 2450 1760
rect 2300 1705 2325 1740
rect 2425 1705 2450 1740
rect 2300 1700 2450 1705
rect 2550 1795 2700 1800
rect 2550 1760 2575 1795
rect 2675 1760 2700 1795
rect 2550 1740 2700 1760
rect 2550 1705 2575 1740
rect 2675 1705 2700 1740
rect 2550 1700 2700 1705
rect 2800 1795 3200 1800
rect 2800 1760 2825 1795
rect 2925 1760 3075 1795
rect 3175 1760 3200 1795
rect 2800 1740 3200 1760
rect 2800 1705 2825 1740
rect 2925 1705 3075 1740
rect 3175 1705 3200 1740
rect 2800 1700 3200 1705
rect 3300 1795 3450 1800
rect 3300 1760 3325 1795
rect 3425 1760 3450 1795
rect 3300 1740 3450 1760
rect 3300 1705 3325 1740
rect 3425 1705 3450 1740
rect 3300 1700 3450 1705
rect 3550 1795 3700 1800
rect 3550 1760 3575 1795
rect 3675 1760 3700 1795
rect 3550 1740 3700 1760
rect 3550 1705 3575 1740
rect 3675 1705 3700 1740
rect 3550 1700 3700 1705
rect 3800 1795 4000 1800
rect 3800 1760 3825 1795
rect 3925 1760 4000 1795
rect 3800 1740 4000 1760
rect 3800 1705 3825 1740
rect 3925 1705 4000 1740
rect 3800 1700 4000 1705
rect 0 1690 60 1700
rect 190 1690 310 1700
rect 440 1690 560 1700
rect 690 1690 810 1700
rect 940 1690 1060 1700
rect 1190 1690 1310 1700
rect 1440 1690 1560 1700
rect 1690 1690 1810 1700
rect 1940 1690 2060 1700
rect 2190 1690 2310 1700
rect 2440 1690 2560 1700
rect 2690 1690 2810 1700
rect 2940 1690 3060 1700
rect 3190 1690 3310 1700
rect 3440 1690 3560 1700
rect 3690 1690 3810 1700
rect 3940 1690 4000 1700
rect 0 1675 50 1690
rect 0 1575 10 1675
rect 45 1575 50 1675
rect 0 1560 50 1575
rect 200 1675 300 1690
rect 200 1575 205 1675
rect 240 1575 260 1675
rect 295 1575 300 1675
rect 200 1560 300 1575
rect 450 1675 550 1690
rect 450 1575 455 1675
rect 490 1575 510 1675
rect 545 1575 550 1675
rect 450 1560 550 1575
rect 700 1675 800 1690
rect 700 1575 705 1675
rect 740 1575 760 1675
rect 795 1575 800 1675
rect 700 1560 800 1575
rect 950 1675 1050 1690
rect 950 1575 955 1675
rect 990 1575 1010 1675
rect 1045 1575 1050 1675
rect 950 1560 1050 1575
rect 1200 1675 1300 1690
rect 1200 1575 1205 1675
rect 1240 1575 1260 1675
rect 1295 1575 1300 1675
rect 1200 1560 1300 1575
rect 1450 1675 1550 1690
rect 1450 1575 1455 1675
rect 1490 1575 1510 1675
rect 1545 1575 1550 1675
rect 1450 1560 1550 1575
rect 1700 1675 1800 1690
rect 1700 1575 1705 1675
rect 1740 1575 1760 1675
rect 1795 1575 1800 1675
rect 1700 1560 1800 1575
rect 1950 1675 2050 1690
rect 1950 1575 1955 1675
rect 1990 1575 2010 1675
rect 2045 1575 2050 1675
rect 1950 1560 2050 1575
rect 2200 1675 2300 1690
rect 2200 1575 2205 1675
rect 2240 1575 2260 1675
rect 2295 1575 2300 1675
rect 2200 1560 2300 1575
rect 2450 1675 2550 1690
rect 2450 1575 2455 1675
rect 2490 1575 2510 1675
rect 2545 1575 2550 1675
rect 2450 1560 2550 1575
rect 2700 1675 2800 1690
rect 2700 1575 2705 1675
rect 2740 1575 2760 1675
rect 2795 1575 2800 1675
rect 2700 1560 2800 1575
rect 2950 1675 3050 1690
rect 2950 1575 2955 1675
rect 2990 1575 3010 1675
rect 3045 1575 3050 1675
rect 2950 1560 3050 1575
rect 3200 1675 3300 1690
rect 3200 1575 3205 1675
rect 3240 1575 3260 1675
rect 3295 1575 3300 1675
rect 3200 1560 3300 1575
rect 3450 1675 3550 1690
rect 3450 1575 3455 1675
rect 3490 1575 3510 1675
rect 3545 1575 3550 1675
rect 3450 1560 3550 1575
rect 3700 1675 3800 1690
rect 3700 1575 3705 1675
rect 3740 1575 3760 1675
rect 3795 1575 3800 1675
rect 3700 1560 3800 1575
rect 3950 1675 4000 1690
rect 3950 1575 3955 1675
rect 3990 1575 4000 1675
rect 3950 1560 4000 1575
rect 0 1550 60 1560
rect 190 1550 310 1560
rect 440 1550 560 1560
rect 690 1550 810 1560
rect 940 1550 1060 1560
rect 1190 1550 1310 1560
rect 1440 1550 1560 1560
rect 1690 1550 1810 1560
rect 1940 1550 2060 1560
rect 2190 1550 2310 1560
rect 2440 1550 2560 1560
rect 2690 1550 2810 1560
rect 2940 1550 3060 1560
rect 3190 1550 3310 1560
rect 3440 1550 3560 1560
rect 3690 1550 3810 1560
rect 3940 1550 4000 1560
rect 0 1545 200 1550
rect 0 1510 75 1545
rect 175 1510 200 1545
rect 0 1490 200 1510
rect 0 1455 75 1490
rect 175 1455 200 1490
rect 0 1450 200 1455
rect 300 1545 450 1550
rect 300 1510 325 1545
rect 425 1510 450 1545
rect 300 1490 450 1510
rect 300 1455 325 1490
rect 425 1455 450 1490
rect 300 1450 450 1455
rect 550 1545 700 1550
rect 550 1510 575 1545
rect 675 1510 700 1545
rect 550 1490 700 1510
rect 550 1455 575 1490
rect 675 1455 700 1490
rect 550 1450 700 1455
rect 800 1545 950 1550
rect 800 1510 825 1545
rect 925 1510 950 1545
rect 800 1490 950 1510
rect 800 1455 825 1490
rect 925 1455 950 1490
rect 800 1450 950 1455
rect 1050 1545 1200 1550
rect 1050 1510 1075 1545
rect 1175 1510 1200 1545
rect 1050 1490 1200 1510
rect 1050 1455 1075 1490
rect 1175 1455 1200 1490
rect 1050 1450 1200 1455
rect 1300 1545 1450 1550
rect 1300 1510 1325 1545
rect 1425 1510 1450 1545
rect 1300 1490 1450 1510
rect 1300 1455 1325 1490
rect 1425 1455 1450 1490
rect 1300 1450 1450 1455
rect 1550 1545 1700 1550
rect 1550 1510 1575 1545
rect 1675 1510 1700 1545
rect 1550 1490 1700 1510
rect 1550 1455 1575 1490
rect 1675 1455 1700 1490
rect 1550 1450 1700 1455
rect 1800 1545 2200 1550
rect 1800 1510 1825 1545
rect 1925 1510 2075 1545
rect 2175 1510 2200 1545
rect 1800 1490 2200 1510
rect 1800 1455 1825 1490
rect 1925 1455 2075 1490
rect 2175 1455 2200 1490
rect 1800 1450 2200 1455
rect 2300 1545 2450 1550
rect 2300 1510 2325 1545
rect 2425 1510 2450 1545
rect 2300 1490 2450 1510
rect 2300 1455 2325 1490
rect 2425 1455 2450 1490
rect 2300 1450 2450 1455
rect 2550 1545 2700 1550
rect 2550 1510 2575 1545
rect 2675 1510 2700 1545
rect 2550 1490 2700 1510
rect 2550 1455 2575 1490
rect 2675 1455 2700 1490
rect 2550 1450 2700 1455
rect 2800 1545 2950 1550
rect 2800 1510 2825 1545
rect 2925 1510 2950 1545
rect 2800 1490 2950 1510
rect 2800 1455 2825 1490
rect 2925 1455 2950 1490
rect 2800 1450 2950 1455
rect 3050 1545 3200 1550
rect 3050 1510 3075 1545
rect 3175 1510 3200 1545
rect 3050 1490 3200 1510
rect 3050 1455 3075 1490
rect 3175 1455 3200 1490
rect 3050 1450 3200 1455
rect 3300 1545 3450 1550
rect 3300 1510 3325 1545
rect 3425 1510 3450 1545
rect 3300 1490 3450 1510
rect 3300 1455 3325 1490
rect 3425 1455 3450 1490
rect 3300 1450 3450 1455
rect 3550 1545 3700 1550
rect 3550 1510 3575 1545
rect 3675 1510 3700 1545
rect 3550 1490 3700 1510
rect 3550 1455 3575 1490
rect 3675 1455 3700 1490
rect 3550 1450 3700 1455
rect 3800 1545 4000 1550
rect 3800 1510 3825 1545
rect 3925 1510 4000 1545
rect 3800 1490 4000 1510
rect 3800 1455 3825 1490
rect 3925 1455 4000 1490
rect 3800 1450 4000 1455
rect 0 1440 60 1450
rect 190 1440 310 1450
rect 440 1440 560 1450
rect 690 1440 810 1450
rect 940 1440 1060 1450
rect 1190 1440 1310 1450
rect 1440 1440 1560 1450
rect 1690 1440 1810 1450
rect 1940 1440 2060 1450
rect 2190 1440 2310 1450
rect 2440 1440 2560 1450
rect 2690 1440 2810 1450
rect 2940 1440 3060 1450
rect 3190 1440 3310 1450
rect 3440 1440 3560 1450
rect 3690 1440 3810 1450
rect 3940 1440 4000 1450
rect 0 1425 50 1440
rect 0 1325 10 1425
rect 45 1325 50 1425
rect 0 1310 50 1325
rect 200 1425 300 1440
rect 200 1325 205 1425
rect 240 1325 260 1425
rect 295 1325 300 1425
rect 200 1310 300 1325
rect 450 1425 550 1440
rect 450 1325 455 1425
rect 490 1325 510 1425
rect 545 1325 550 1425
rect 450 1310 550 1325
rect 700 1425 800 1440
rect 700 1325 705 1425
rect 740 1325 760 1425
rect 795 1325 800 1425
rect 700 1310 800 1325
rect 950 1425 1050 1440
rect 950 1325 955 1425
rect 990 1325 1010 1425
rect 1045 1325 1050 1425
rect 950 1310 1050 1325
rect 1200 1425 1300 1440
rect 1200 1325 1205 1425
rect 1240 1325 1260 1425
rect 1295 1325 1300 1425
rect 1200 1310 1300 1325
rect 1450 1425 1550 1440
rect 1450 1325 1455 1425
rect 1490 1325 1510 1425
rect 1545 1325 1550 1425
rect 1450 1310 1550 1325
rect 1700 1425 1800 1440
rect 1700 1325 1705 1425
rect 1740 1325 1760 1425
rect 1795 1325 1800 1425
rect 1700 1310 1800 1325
rect 1950 1425 2050 1440
rect 1950 1325 1955 1425
rect 1990 1325 2010 1425
rect 2045 1325 2050 1425
rect 1950 1310 2050 1325
rect 2200 1425 2300 1440
rect 2200 1325 2205 1425
rect 2240 1325 2260 1425
rect 2295 1325 2300 1425
rect 2200 1310 2300 1325
rect 2450 1425 2550 1440
rect 2450 1325 2455 1425
rect 2490 1325 2510 1425
rect 2545 1325 2550 1425
rect 2450 1310 2550 1325
rect 2700 1425 2800 1440
rect 2700 1325 2705 1425
rect 2740 1325 2760 1425
rect 2795 1325 2800 1425
rect 2700 1310 2800 1325
rect 2950 1425 3050 1440
rect 2950 1325 2955 1425
rect 2990 1325 3010 1425
rect 3045 1325 3050 1425
rect 2950 1310 3050 1325
rect 3200 1425 3300 1440
rect 3200 1325 3205 1425
rect 3240 1325 3260 1425
rect 3295 1325 3300 1425
rect 3200 1310 3300 1325
rect 3450 1425 3550 1440
rect 3450 1325 3455 1425
rect 3490 1325 3510 1425
rect 3545 1325 3550 1425
rect 3450 1310 3550 1325
rect 3700 1425 3800 1440
rect 3700 1325 3705 1425
rect 3740 1325 3760 1425
rect 3795 1325 3800 1425
rect 3700 1310 3800 1325
rect 3950 1425 4000 1440
rect 3950 1325 3955 1425
rect 3990 1325 4000 1425
rect 3950 1310 4000 1325
rect 0 1300 60 1310
rect 190 1300 310 1310
rect 440 1300 560 1310
rect 690 1300 810 1310
rect 940 1300 1060 1310
rect 1190 1300 1310 1310
rect 1440 1300 1560 1310
rect 1690 1300 1810 1310
rect 1940 1300 2060 1310
rect 2190 1300 2310 1310
rect 2440 1300 2560 1310
rect 2690 1300 2810 1310
rect 2940 1300 3060 1310
rect 3190 1300 3310 1310
rect 3440 1300 3560 1310
rect 3690 1300 3810 1310
rect 3940 1300 4000 1310
rect 0 1295 200 1300
rect 0 1260 75 1295
rect 175 1260 200 1295
rect 0 1240 200 1260
rect 0 1205 75 1240
rect 175 1205 200 1240
rect 0 1200 200 1205
rect 300 1295 450 1300
rect 300 1260 325 1295
rect 425 1260 450 1295
rect 300 1240 450 1260
rect 300 1205 325 1240
rect 425 1205 450 1240
rect 300 1200 450 1205
rect 550 1295 700 1300
rect 550 1260 575 1295
rect 675 1260 700 1295
rect 550 1240 700 1260
rect 550 1205 575 1240
rect 675 1205 700 1240
rect 550 1200 700 1205
rect 800 1295 1200 1300
rect 800 1260 825 1295
rect 925 1260 1075 1295
rect 1175 1260 1200 1295
rect 800 1240 1200 1260
rect 800 1205 825 1240
rect 925 1205 1075 1240
rect 1175 1205 1200 1240
rect 800 1200 1200 1205
rect 1300 1295 1450 1300
rect 1300 1260 1325 1295
rect 1425 1260 1450 1295
rect 1300 1240 1450 1260
rect 1300 1205 1325 1240
rect 1425 1205 1450 1240
rect 1300 1200 1450 1205
rect 1550 1295 1700 1300
rect 1550 1260 1575 1295
rect 1675 1260 1700 1295
rect 1550 1240 1700 1260
rect 1550 1205 1575 1240
rect 1675 1205 1700 1240
rect 1550 1200 1700 1205
rect 1800 1295 2200 1300
rect 1800 1260 1825 1295
rect 1925 1260 2075 1295
rect 2175 1260 2200 1295
rect 1800 1240 2200 1260
rect 1800 1205 1825 1240
rect 1925 1205 2075 1240
rect 2175 1205 2200 1240
rect 1800 1200 2200 1205
rect 2300 1295 2450 1300
rect 2300 1260 2325 1295
rect 2425 1260 2450 1295
rect 2300 1240 2450 1260
rect 2300 1205 2325 1240
rect 2425 1205 2450 1240
rect 2300 1200 2450 1205
rect 2550 1295 2700 1300
rect 2550 1260 2575 1295
rect 2675 1260 2700 1295
rect 2550 1240 2700 1260
rect 2550 1205 2575 1240
rect 2675 1205 2700 1240
rect 2550 1200 2700 1205
rect 2800 1295 3200 1300
rect 2800 1260 2825 1295
rect 2925 1260 3075 1295
rect 3175 1260 3200 1295
rect 2800 1240 3200 1260
rect 2800 1205 2825 1240
rect 2925 1205 3075 1240
rect 3175 1205 3200 1240
rect 2800 1200 3200 1205
rect 3300 1295 3450 1300
rect 3300 1260 3325 1295
rect 3425 1260 3450 1295
rect 3300 1240 3450 1260
rect 3300 1205 3325 1240
rect 3425 1205 3450 1240
rect 3300 1200 3450 1205
rect 3550 1295 3700 1300
rect 3550 1260 3575 1295
rect 3675 1260 3700 1295
rect 3550 1240 3700 1260
rect 3550 1205 3575 1240
rect 3675 1205 3700 1240
rect 3550 1200 3700 1205
rect 3800 1295 4000 1300
rect 3800 1260 3825 1295
rect 3925 1260 4000 1295
rect 3800 1240 4000 1260
rect 3800 1205 3825 1240
rect 3925 1205 4000 1240
rect 3800 1200 4000 1205
rect 0 1190 60 1200
rect 190 1190 310 1200
rect 440 1190 560 1200
rect 690 1190 810 1200
rect 940 1190 1060 1200
rect 1190 1190 1310 1200
rect 1440 1190 1560 1200
rect 1690 1190 1810 1200
rect 1940 1190 2060 1200
rect 2190 1190 2310 1200
rect 2440 1190 2560 1200
rect 2690 1190 2810 1200
rect 2940 1190 3060 1200
rect 3190 1190 3310 1200
rect 3440 1190 3560 1200
rect 3690 1190 3810 1200
rect 3940 1190 4000 1200
rect 0 1175 50 1190
rect 0 1075 10 1175
rect 45 1075 50 1175
rect 0 1060 50 1075
rect 200 1175 300 1190
rect 200 1075 205 1175
rect 240 1075 260 1175
rect 295 1075 300 1175
rect 200 1060 300 1075
rect 450 1175 550 1190
rect 450 1075 455 1175
rect 490 1075 510 1175
rect 545 1075 550 1175
rect 450 1060 550 1075
rect 700 1175 800 1190
rect 700 1075 705 1175
rect 740 1075 760 1175
rect 795 1075 800 1175
rect 700 1060 800 1075
rect 950 1175 1050 1190
rect 950 1075 955 1175
rect 990 1075 1010 1175
rect 1045 1075 1050 1175
rect 950 1060 1050 1075
rect 1200 1175 1300 1190
rect 1200 1075 1205 1175
rect 1240 1075 1260 1175
rect 1295 1075 1300 1175
rect 1200 1060 1300 1075
rect 1450 1175 1550 1190
rect 1450 1075 1455 1175
rect 1490 1075 1510 1175
rect 1545 1075 1550 1175
rect 1450 1060 1550 1075
rect 1700 1175 1800 1190
rect 1700 1075 1705 1175
rect 1740 1075 1760 1175
rect 1795 1075 1800 1175
rect 1700 1060 1800 1075
rect 1950 1175 2050 1190
rect 1950 1075 1955 1175
rect 1990 1075 2010 1175
rect 2045 1075 2050 1175
rect 1950 1060 2050 1075
rect 2200 1175 2300 1190
rect 2200 1075 2205 1175
rect 2240 1075 2260 1175
rect 2295 1075 2300 1175
rect 2200 1060 2300 1075
rect 2450 1175 2550 1190
rect 2450 1075 2455 1175
rect 2490 1075 2510 1175
rect 2545 1075 2550 1175
rect 2450 1060 2550 1075
rect 2700 1175 2800 1190
rect 2700 1075 2705 1175
rect 2740 1075 2760 1175
rect 2795 1075 2800 1175
rect 2700 1060 2800 1075
rect 2950 1175 3050 1190
rect 2950 1075 2955 1175
rect 2990 1075 3010 1175
rect 3045 1075 3050 1175
rect 2950 1060 3050 1075
rect 3200 1175 3300 1190
rect 3200 1075 3205 1175
rect 3240 1075 3260 1175
rect 3295 1075 3300 1175
rect 3200 1060 3300 1075
rect 3450 1175 3550 1190
rect 3450 1075 3455 1175
rect 3490 1075 3510 1175
rect 3545 1075 3550 1175
rect 3450 1060 3550 1075
rect 3700 1175 3800 1190
rect 3700 1075 3705 1175
rect 3740 1075 3760 1175
rect 3795 1075 3800 1175
rect 3700 1060 3800 1075
rect 3950 1175 4000 1190
rect 3950 1075 3955 1175
rect 3990 1075 4000 1175
rect 3950 1060 4000 1075
rect 0 1050 60 1060
rect 190 1050 310 1060
rect 440 1050 560 1060
rect 690 1050 810 1060
rect 940 1050 1060 1060
rect 1190 1050 1310 1060
rect 1440 1050 1560 1060
rect 1690 1050 1810 1060
rect 1940 1050 2060 1060
rect 2190 1050 2310 1060
rect 2440 1050 2560 1060
rect 2690 1050 2810 1060
rect 2940 1050 3060 1060
rect 3190 1050 3310 1060
rect 3440 1050 3560 1060
rect 3690 1050 3810 1060
rect 3940 1050 4000 1060
rect 0 1045 450 1050
rect 0 1010 75 1045
rect 175 1010 325 1045
rect 425 1010 450 1045
rect 0 990 450 1010
rect 0 955 75 990
rect 175 955 325 990
rect 425 955 450 990
rect 0 950 450 955
rect 550 1045 1450 1050
rect 550 1010 575 1045
rect 675 1010 825 1045
rect 925 1010 1075 1045
rect 1175 1010 1325 1045
rect 1425 1010 1450 1045
rect 550 990 1450 1010
rect 550 955 575 990
rect 675 955 825 990
rect 925 955 1075 990
rect 1175 955 1325 990
rect 1425 955 1450 990
rect 550 950 1450 955
rect 1550 1045 2450 1050
rect 1550 1010 1575 1045
rect 1675 1010 1825 1045
rect 1925 1010 2075 1045
rect 2175 1010 2325 1045
rect 2425 1010 2450 1045
rect 1550 990 2450 1010
rect 1550 955 1575 990
rect 1675 955 1825 990
rect 1925 955 2075 990
rect 2175 955 2325 990
rect 2425 955 2450 990
rect 1550 950 2450 955
rect 2550 1045 3450 1050
rect 2550 1010 2575 1045
rect 2675 1010 2825 1045
rect 2925 1010 3075 1045
rect 3175 1010 3325 1045
rect 3425 1010 3450 1045
rect 2550 990 3450 1010
rect 2550 955 2575 990
rect 2675 955 2825 990
rect 2925 955 3075 990
rect 3175 955 3325 990
rect 3425 955 3450 990
rect 2550 950 3450 955
rect 3550 1045 4000 1050
rect 3550 1010 3575 1045
rect 3675 1010 3825 1045
rect 3925 1010 4000 1045
rect 3550 990 4000 1010
rect 3550 955 3575 990
rect 3675 955 3825 990
rect 3925 955 4000 990
rect 3550 950 4000 955
rect 0 940 60 950
rect 190 940 310 950
rect 440 940 560 950
rect 690 940 810 950
rect 940 940 1060 950
rect 1190 940 1310 950
rect 1440 940 1560 950
rect 1690 940 1810 950
rect 1940 940 2060 950
rect 2190 940 2310 950
rect 2440 940 2560 950
rect 2690 940 2810 950
rect 2940 940 3060 950
rect 3190 940 3310 950
rect 3440 940 3560 950
rect 3690 940 3810 950
rect 3940 940 4000 950
rect 0 925 50 940
rect 0 825 10 925
rect 45 825 50 925
rect 0 810 50 825
rect 200 925 300 940
rect 200 825 205 925
rect 240 825 260 925
rect 295 825 300 925
rect 200 810 300 825
rect 450 925 550 940
rect 450 825 455 925
rect 490 825 510 925
rect 545 825 550 925
rect 450 810 550 825
rect 700 925 800 940
rect 700 825 705 925
rect 740 825 760 925
rect 795 825 800 925
rect 700 810 800 825
rect 950 925 1050 940
rect 950 825 955 925
rect 990 825 1010 925
rect 1045 825 1050 925
rect 950 810 1050 825
rect 1200 925 1300 940
rect 1200 825 1205 925
rect 1240 825 1260 925
rect 1295 825 1300 925
rect 1200 810 1300 825
rect 1450 925 1550 940
rect 1450 825 1455 925
rect 1490 825 1510 925
rect 1545 825 1550 925
rect 1450 810 1550 825
rect 1700 925 1800 940
rect 1700 825 1705 925
rect 1740 825 1760 925
rect 1795 825 1800 925
rect 1700 810 1800 825
rect 1950 925 2050 940
rect 1950 825 1955 925
rect 1990 825 2010 925
rect 2045 825 2050 925
rect 1950 810 2050 825
rect 2200 925 2300 940
rect 2200 825 2205 925
rect 2240 825 2260 925
rect 2295 825 2300 925
rect 2200 810 2300 825
rect 2450 925 2550 940
rect 2450 825 2455 925
rect 2490 825 2510 925
rect 2545 825 2550 925
rect 2450 810 2550 825
rect 2700 925 2800 940
rect 2700 825 2705 925
rect 2740 825 2760 925
rect 2795 825 2800 925
rect 2700 810 2800 825
rect 2950 925 3050 940
rect 2950 825 2955 925
rect 2990 825 3010 925
rect 3045 825 3050 925
rect 2950 810 3050 825
rect 3200 925 3300 940
rect 3200 825 3205 925
rect 3240 825 3260 925
rect 3295 825 3300 925
rect 3200 810 3300 825
rect 3450 925 3550 940
rect 3450 825 3455 925
rect 3490 825 3510 925
rect 3545 825 3550 925
rect 3450 810 3550 825
rect 3700 925 3800 940
rect 3700 825 3705 925
rect 3740 825 3760 925
rect 3795 825 3800 925
rect 3700 810 3800 825
rect 3950 925 4000 940
rect 3950 825 3955 925
rect 3990 825 4000 925
rect 3950 810 4000 825
rect 0 800 60 810
rect 190 800 310 810
rect 440 800 560 810
rect 690 800 810 810
rect 940 800 1060 810
rect 1190 800 1310 810
rect 1440 800 1560 810
rect 1690 800 1810 810
rect 1940 800 2060 810
rect 2190 800 2310 810
rect 2440 800 2560 810
rect 2690 800 2810 810
rect 2940 800 3060 810
rect 3190 800 3310 810
rect 3440 800 3560 810
rect 3690 800 3810 810
rect 3940 800 4000 810
rect 0 795 200 800
rect 0 760 75 795
rect 175 760 200 795
rect 0 740 200 760
rect 0 705 75 740
rect 175 705 200 740
rect 0 700 200 705
rect 300 795 450 800
rect 300 760 325 795
rect 425 760 450 795
rect 300 740 450 760
rect 300 705 325 740
rect 425 705 450 740
rect 300 700 450 705
rect 550 795 700 800
rect 550 760 575 795
rect 675 760 700 795
rect 550 740 700 760
rect 550 705 575 740
rect 675 705 700 740
rect 550 700 700 705
rect 800 795 1200 800
rect 800 760 825 795
rect 925 760 1075 795
rect 1175 760 1200 795
rect 800 740 1200 760
rect 800 705 825 740
rect 925 705 1075 740
rect 1175 705 1200 740
rect 800 700 1200 705
rect 1300 795 1450 800
rect 1300 760 1325 795
rect 1425 760 1450 795
rect 1300 740 1450 760
rect 1300 705 1325 740
rect 1425 705 1450 740
rect 1300 700 1450 705
rect 1550 795 1700 800
rect 1550 760 1575 795
rect 1675 760 1700 795
rect 1550 740 1700 760
rect 1550 705 1575 740
rect 1675 705 1700 740
rect 1550 700 1700 705
rect 1800 795 2200 800
rect 1800 760 1825 795
rect 1925 760 2075 795
rect 2175 760 2200 795
rect 1800 740 2200 760
rect 1800 705 1825 740
rect 1925 705 2075 740
rect 2175 705 2200 740
rect 1800 700 2200 705
rect 2300 795 2450 800
rect 2300 760 2325 795
rect 2425 760 2450 795
rect 2300 740 2450 760
rect 2300 705 2325 740
rect 2425 705 2450 740
rect 2300 700 2450 705
rect 2550 795 2700 800
rect 2550 760 2575 795
rect 2675 760 2700 795
rect 2550 740 2700 760
rect 2550 705 2575 740
rect 2675 705 2700 740
rect 2550 700 2700 705
rect 2800 795 3200 800
rect 2800 760 2825 795
rect 2925 760 3075 795
rect 3175 760 3200 795
rect 2800 740 3200 760
rect 2800 705 2825 740
rect 2925 705 3075 740
rect 3175 705 3200 740
rect 2800 700 3200 705
rect 3300 795 3450 800
rect 3300 760 3325 795
rect 3425 760 3450 795
rect 3300 740 3450 760
rect 3300 705 3325 740
rect 3425 705 3450 740
rect 3300 700 3450 705
rect 3550 795 3700 800
rect 3550 760 3575 795
rect 3675 760 3700 795
rect 3550 740 3700 760
rect 3550 705 3575 740
rect 3675 705 3700 740
rect 3550 700 3700 705
rect 3800 795 4000 800
rect 3800 760 3825 795
rect 3925 760 4000 795
rect 3800 740 4000 760
rect 3800 705 3825 740
rect 3925 705 4000 740
rect 3800 700 4000 705
rect 0 690 60 700
rect 190 690 310 700
rect 440 690 560 700
rect 690 690 810 700
rect 940 690 1060 700
rect 1190 690 1310 700
rect 1440 690 1560 700
rect 1690 690 1810 700
rect 1940 690 2060 700
rect 2190 690 2310 700
rect 2440 690 2560 700
rect 2690 690 2810 700
rect 2940 690 3060 700
rect 3190 690 3310 700
rect 3440 690 3560 700
rect 3690 690 3810 700
rect 3940 690 4000 700
rect 0 675 50 690
rect 0 575 10 675
rect 45 575 50 675
rect 0 560 50 575
rect 200 675 300 690
rect 200 575 205 675
rect 240 575 260 675
rect 295 575 300 675
rect 200 560 300 575
rect 450 675 550 690
rect 450 575 455 675
rect 490 575 510 675
rect 545 575 550 675
rect 450 560 550 575
rect 700 675 800 690
rect 700 575 705 675
rect 740 575 760 675
rect 795 575 800 675
rect 700 560 800 575
rect 950 675 1050 690
rect 950 575 955 675
rect 990 575 1010 675
rect 1045 575 1050 675
rect 950 560 1050 575
rect 1200 675 1300 690
rect 1200 575 1205 675
rect 1240 575 1260 675
rect 1295 575 1300 675
rect 1200 560 1300 575
rect 1450 675 1550 690
rect 1450 575 1455 675
rect 1490 575 1510 675
rect 1545 575 1550 675
rect 1450 560 1550 575
rect 1700 675 1800 690
rect 1700 575 1705 675
rect 1740 575 1760 675
rect 1795 575 1800 675
rect 1700 560 1800 575
rect 1950 675 2050 690
rect 1950 575 1955 675
rect 1990 575 2010 675
rect 2045 575 2050 675
rect 1950 560 2050 575
rect 2200 675 2300 690
rect 2200 575 2205 675
rect 2240 575 2260 675
rect 2295 575 2300 675
rect 2200 560 2300 575
rect 2450 675 2550 690
rect 2450 575 2455 675
rect 2490 575 2510 675
rect 2545 575 2550 675
rect 2450 560 2550 575
rect 2700 675 2800 690
rect 2700 575 2705 675
rect 2740 575 2760 675
rect 2795 575 2800 675
rect 2700 560 2800 575
rect 2950 675 3050 690
rect 2950 575 2955 675
rect 2990 575 3010 675
rect 3045 575 3050 675
rect 2950 560 3050 575
rect 3200 675 3300 690
rect 3200 575 3205 675
rect 3240 575 3260 675
rect 3295 575 3300 675
rect 3200 560 3300 575
rect 3450 675 3550 690
rect 3450 575 3455 675
rect 3490 575 3510 675
rect 3545 575 3550 675
rect 3450 560 3550 575
rect 3700 675 3800 690
rect 3700 575 3705 675
rect 3740 575 3760 675
rect 3795 575 3800 675
rect 3700 560 3800 575
rect 3950 675 4000 690
rect 3950 575 3955 675
rect 3990 575 4000 675
rect 3950 560 4000 575
rect 0 550 60 560
rect 190 550 310 560
rect 440 550 560 560
rect 690 550 810 560
rect 940 550 1060 560
rect 1190 550 1310 560
rect 1440 550 1560 560
rect 1690 550 1810 560
rect 1940 550 2060 560
rect 2190 550 2310 560
rect 2440 550 2560 560
rect 2690 550 2810 560
rect 2940 550 3060 560
rect 3190 550 3310 560
rect 3440 550 3560 560
rect 3690 550 3810 560
rect 3940 550 4000 560
rect 0 545 200 550
rect 0 510 75 545
rect 175 510 200 545
rect 0 490 200 510
rect 0 455 75 490
rect 175 455 200 490
rect 0 450 200 455
rect 300 545 450 550
rect 300 510 325 545
rect 425 510 450 545
rect 300 490 450 510
rect 300 455 325 490
rect 425 455 450 490
rect 300 450 450 455
rect 550 545 700 550
rect 550 510 575 545
rect 675 510 700 545
rect 550 490 700 510
rect 550 455 575 490
rect 675 455 700 490
rect 550 450 700 455
rect 800 545 950 550
rect 800 510 825 545
rect 925 510 950 545
rect 800 490 950 510
rect 800 455 825 490
rect 925 455 950 490
rect 800 450 950 455
rect 1050 545 1200 550
rect 1050 510 1075 545
rect 1175 510 1200 545
rect 1050 490 1200 510
rect 1050 455 1075 490
rect 1175 455 1200 490
rect 1050 450 1200 455
rect 1300 545 1450 550
rect 1300 510 1325 545
rect 1425 510 1450 545
rect 1300 490 1450 510
rect 1300 455 1325 490
rect 1425 455 1450 490
rect 1300 450 1450 455
rect 1550 545 1700 550
rect 1550 510 1575 545
rect 1675 510 1700 545
rect 1550 490 1700 510
rect 1550 455 1575 490
rect 1675 455 1700 490
rect 1550 450 1700 455
rect 1800 545 2200 550
rect 1800 510 1825 545
rect 1925 510 2075 545
rect 2175 510 2200 545
rect 1800 490 2200 510
rect 1800 455 1825 490
rect 1925 455 2075 490
rect 2175 455 2200 490
rect 1800 450 2200 455
rect 2300 545 2450 550
rect 2300 510 2325 545
rect 2425 510 2450 545
rect 2300 490 2450 510
rect 2300 455 2325 490
rect 2425 455 2450 490
rect 2300 450 2450 455
rect 2550 545 2700 550
rect 2550 510 2575 545
rect 2675 510 2700 545
rect 2550 490 2700 510
rect 2550 455 2575 490
rect 2675 455 2700 490
rect 2550 450 2700 455
rect 2800 545 2950 550
rect 2800 510 2825 545
rect 2925 510 2950 545
rect 2800 490 2950 510
rect 2800 455 2825 490
rect 2925 455 2950 490
rect 2800 450 2950 455
rect 3050 545 3200 550
rect 3050 510 3075 545
rect 3175 510 3200 545
rect 3050 490 3200 510
rect 3050 455 3075 490
rect 3175 455 3200 490
rect 3050 450 3200 455
rect 3300 545 3450 550
rect 3300 510 3325 545
rect 3425 510 3450 545
rect 3300 490 3450 510
rect 3300 455 3325 490
rect 3425 455 3450 490
rect 3300 450 3450 455
rect 3550 545 3700 550
rect 3550 510 3575 545
rect 3675 510 3700 545
rect 3550 490 3700 510
rect 3550 455 3575 490
rect 3675 455 3700 490
rect 3550 450 3700 455
rect 3800 545 4000 550
rect 3800 510 3825 545
rect 3925 510 4000 545
rect 3800 490 4000 510
rect 3800 455 3825 490
rect 3925 455 4000 490
rect 3800 450 4000 455
rect 0 440 60 450
rect 190 440 310 450
rect 440 440 560 450
rect 690 440 810 450
rect 940 440 1060 450
rect 1190 440 1310 450
rect 1440 440 1560 450
rect 1690 440 1810 450
rect 1940 440 2060 450
rect 2190 440 2310 450
rect 2440 440 2560 450
rect 2690 440 2810 450
rect 2940 440 3060 450
rect 3190 440 3310 450
rect 3440 440 3560 450
rect 3690 440 3810 450
rect 3940 440 4000 450
rect 0 425 50 440
rect 0 325 10 425
rect 45 325 50 425
rect 0 310 50 325
rect 200 425 300 440
rect 200 325 205 425
rect 240 325 260 425
rect 295 325 300 425
rect 200 310 300 325
rect 450 425 550 440
rect 450 325 455 425
rect 490 325 510 425
rect 545 325 550 425
rect 450 310 550 325
rect 700 425 800 440
rect 700 325 705 425
rect 740 325 760 425
rect 795 325 800 425
rect 700 310 800 325
rect 950 425 1050 440
rect 950 325 955 425
rect 990 325 1010 425
rect 1045 325 1050 425
rect 950 310 1050 325
rect 1200 425 1300 440
rect 1200 325 1205 425
rect 1240 325 1260 425
rect 1295 325 1300 425
rect 1200 310 1300 325
rect 1450 425 1550 440
rect 1450 325 1455 425
rect 1490 325 1510 425
rect 1545 325 1550 425
rect 1450 310 1550 325
rect 1700 425 1800 440
rect 1700 325 1705 425
rect 1740 325 1760 425
rect 1795 325 1800 425
rect 1700 310 1800 325
rect 1950 425 2050 440
rect 1950 325 1955 425
rect 1990 325 2010 425
rect 2045 325 2050 425
rect 1950 310 2050 325
rect 2200 425 2300 440
rect 2200 325 2205 425
rect 2240 325 2260 425
rect 2295 325 2300 425
rect 2200 310 2300 325
rect 2450 425 2550 440
rect 2450 325 2455 425
rect 2490 325 2510 425
rect 2545 325 2550 425
rect 2450 310 2550 325
rect 2700 425 2800 440
rect 2700 325 2705 425
rect 2740 325 2760 425
rect 2795 325 2800 425
rect 2700 310 2800 325
rect 2950 425 3050 440
rect 2950 325 2955 425
rect 2990 325 3010 425
rect 3045 325 3050 425
rect 2950 310 3050 325
rect 3200 425 3300 440
rect 3200 325 3205 425
rect 3240 325 3260 425
rect 3295 325 3300 425
rect 3200 310 3300 325
rect 3450 425 3550 440
rect 3450 325 3455 425
rect 3490 325 3510 425
rect 3545 325 3550 425
rect 3450 310 3550 325
rect 3700 425 3800 440
rect 3700 325 3705 425
rect 3740 325 3760 425
rect 3795 325 3800 425
rect 3700 310 3800 325
rect 3950 425 4000 440
rect 3950 325 3955 425
rect 3990 325 4000 425
rect 3950 310 4000 325
rect 0 300 60 310
rect 190 300 310 310
rect 440 300 560 310
rect 690 300 810 310
rect 940 300 1060 310
rect 1190 300 1310 310
rect 1440 300 1560 310
rect 1690 300 1810 310
rect 1940 300 2060 310
rect 2190 300 2310 310
rect 2440 300 2560 310
rect 2690 300 2810 310
rect 2940 300 3060 310
rect 3190 300 3310 310
rect 3440 300 3560 310
rect 3690 300 3810 310
rect 3940 300 4000 310
rect 0 295 200 300
rect 0 260 75 295
rect 175 260 200 295
rect 0 240 200 260
rect 0 205 75 240
rect 175 205 200 240
rect 0 200 200 205
rect 300 295 450 300
rect 300 260 325 295
rect 425 260 450 295
rect 300 240 450 260
rect 300 205 325 240
rect 425 205 450 240
rect 300 200 450 205
rect 550 295 700 300
rect 550 260 575 295
rect 675 260 700 295
rect 550 240 700 260
rect 550 205 575 240
rect 675 205 700 240
rect 550 200 700 205
rect 800 295 1200 300
rect 800 260 825 295
rect 925 260 1075 295
rect 1175 260 1200 295
rect 800 240 1200 260
rect 800 205 825 240
rect 925 205 1075 240
rect 1175 205 1200 240
rect 800 200 1200 205
rect 1300 295 1450 300
rect 1300 260 1325 295
rect 1425 260 1450 295
rect 1300 240 1450 260
rect 1300 205 1325 240
rect 1425 205 1450 240
rect 1300 200 1450 205
rect 1550 295 1700 300
rect 1550 260 1575 295
rect 1675 260 1700 295
rect 1550 240 1700 260
rect 1550 205 1575 240
rect 1675 205 1700 240
rect 1550 200 1700 205
rect 1800 295 2200 300
rect 1800 260 1825 295
rect 1925 260 2075 295
rect 2175 260 2200 295
rect 1800 240 2200 260
rect 1800 205 1825 240
rect 1925 205 2075 240
rect 2175 205 2200 240
rect 1800 200 2200 205
rect 2300 295 2450 300
rect 2300 260 2325 295
rect 2425 260 2450 295
rect 2300 240 2450 260
rect 2300 205 2325 240
rect 2425 205 2450 240
rect 2300 200 2450 205
rect 2550 295 2700 300
rect 2550 260 2575 295
rect 2675 260 2700 295
rect 2550 240 2700 260
rect 2550 205 2575 240
rect 2675 205 2700 240
rect 2550 200 2700 205
rect 2800 295 3200 300
rect 2800 260 2825 295
rect 2925 260 3075 295
rect 3175 260 3200 295
rect 2800 240 3200 260
rect 2800 205 2825 240
rect 2925 205 3075 240
rect 3175 205 3200 240
rect 2800 200 3200 205
rect 3300 295 3450 300
rect 3300 260 3325 295
rect 3425 260 3450 295
rect 3300 240 3450 260
rect 3300 205 3325 240
rect 3425 205 3450 240
rect 3300 200 3450 205
rect 3550 295 3700 300
rect 3550 260 3575 295
rect 3675 260 3700 295
rect 3550 240 3700 260
rect 3550 205 3575 240
rect 3675 205 3700 240
rect 3550 200 3700 205
rect 3800 295 4000 300
rect 3800 260 3825 295
rect 3925 260 4000 295
rect 3800 240 4000 260
rect 3800 205 3825 240
rect 3925 205 4000 240
rect 3800 200 4000 205
rect 0 190 60 200
rect 190 190 310 200
rect 440 190 560 200
rect 690 190 810 200
rect 940 190 1060 200
rect 1190 190 1310 200
rect 1440 190 1560 200
rect 1690 190 1810 200
rect 1940 190 2060 200
rect 2190 190 2310 200
rect 2440 190 2560 200
rect 2690 190 2810 200
rect 2940 190 3060 200
rect 3190 190 3310 200
rect 3440 190 3560 200
rect 3690 190 3810 200
rect 3940 190 4000 200
rect 0 175 50 190
rect 0 75 10 175
rect 45 75 50 175
rect 0 60 50 75
rect 200 175 300 190
rect 200 75 205 175
rect 240 75 260 175
rect 295 75 300 175
rect 200 60 300 75
rect 450 175 550 190
rect 450 75 455 175
rect 490 75 510 175
rect 545 75 550 175
rect 450 60 550 75
rect 700 175 800 190
rect 700 75 705 175
rect 740 75 760 175
rect 795 75 800 175
rect 700 60 800 75
rect 950 175 1050 190
rect 950 75 955 175
rect 990 75 1010 175
rect 1045 75 1050 175
rect 950 60 1050 75
rect 1200 175 1300 190
rect 1200 75 1205 175
rect 1240 75 1260 175
rect 1295 75 1300 175
rect 1200 60 1300 75
rect 1450 175 1550 190
rect 1450 75 1455 175
rect 1490 75 1510 175
rect 1545 75 1550 175
rect 1450 60 1550 75
rect 1700 175 1800 190
rect 1700 75 1705 175
rect 1740 75 1760 175
rect 1795 75 1800 175
rect 1700 60 1800 75
rect 1950 175 2050 190
rect 1950 75 1955 175
rect 1990 75 2010 175
rect 2045 75 2050 175
rect 1950 60 2050 75
rect 2200 175 2300 190
rect 2200 75 2205 175
rect 2240 75 2260 175
rect 2295 75 2300 175
rect 2200 60 2300 75
rect 2450 175 2550 190
rect 2450 75 2455 175
rect 2490 75 2510 175
rect 2545 75 2550 175
rect 2450 60 2550 75
rect 2700 175 2800 190
rect 2700 75 2705 175
rect 2740 75 2760 175
rect 2795 75 2800 175
rect 2700 60 2800 75
rect 2950 175 3050 190
rect 2950 75 2955 175
rect 2990 75 3010 175
rect 3045 75 3050 175
rect 2950 60 3050 75
rect 3200 175 3300 190
rect 3200 75 3205 175
rect 3240 75 3260 175
rect 3295 75 3300 175
rect 3200 60 3300 75
rect 3450 175 3550 190
rect 3450 75 3455 175
rect 3490 75 3510 175
rect 3545 75 3550 175
rect 3450 60 3550 75
rect 3700 175 3800 190
rect 3700 75 3705 175
rect 3740 75 3760 175
rect 3795 75 3800 175
rect 3700 60 3800 75
rect 3950 175 4000 190
rect 3950 75 3955 175
rect 3990 75 4000 175
rect 3950 60 4000 75
rect 0 50 60 60
rect 190 50 310 60
rect 440 50 560 60
rect 690 50 810 60
rect 940 50 1060 60
rect 1190 50 1310 60
rect 1440 50 1560 60
rect 1690 50 1810 60
rect 1940 50 2060 60
rect 2190 50 2310 60
rect 2440 50 2560 60
rect 2690 50 2810 60
rect 2940 50 3060 60
rect 3190 50 3310 60
rect 3440 50 3560 60
rect 3690 50 3810 60
rect 3940 50 4000 60
rect 0 45 4000 50
rect 0 10 75 45
rect 175 10 325 45
rect 425 10 575 45
rect 675 10 825 45
rect 925 10 1075 45
rect 1175 10 1325 45
rect 1425 10 1575 45
rect 1675 10 1825 45
rect 1925 10 2075 45
rect 2175 10 2325 45
rect 2425 10 2575 45
rect 2675 10 2825 45
rect 2925 10 3075 45
rect 3175 10 3325 45
rect 3425 10 3575 45
rect 3675 10 3825 45
rect 3925 10 4000 45
rect 0 0 4000 10
<< via3 >>
rect 200 3700 300 3800
rect 450 3700 550 3800
rect 700 3700 800 3800
rect 1200 3700 1300 3800
rect 1450 3700 1550 3800
rect 1700 3700 1800 3800
rect 2200 3700 2300 3800
rect 2450 3700 2550 3800
rect 2700 3700 2800 3800
rect 3200 3700 3300 3800
rect 3450 3700 3550 3800
rect 3700 3700 3800 3800
rect 200 3450 300 3550
rect 450 3450 550 3550
rect 700 3450 800 3550
rect 950 3450 1050 3550
rect 1200 3450 1300 3550
rect 1450 3450 1550 3550
rect 1700 3450 1800 3550
rect 2200 3450 2300 3550
rect 2450 3450 2550 3550
rect 2700 3450 2800 3550
rect 2950 3450 3050 3550
rect 3200 3450 3300 3550
rect 3450 3450 3550 3550
rect 3700 3450 3800 3550
rect 200 3200 300 3300
rect 450 3200 550 3300
rect 700 3200 800 3300
rect 1200 3200 1300 3300
rect 1450 3200 1550 3300
rect 1700 3200 1800 3300
rect 2200 3200 2300 3300
rect 2450 3200 2550 3300
rect 2700 3200 2800 3300
rect 3200 3200 3300 3300
rect 3450 3200 3550 3300
rect 3700 3200 3800 3300
rect 450 2950 550 3050
rect 1450 2950 1550 3050
rect 2450 2950 2550 3050
rect 3450 2950 3550 3050
rect 200 2700 300 2800
rect 450 2700 550 2800
rect 700 2700 800 2800
rect 1200 2700 1300 2800
rect 1450 2700 1550 2800
rect 1700 2700 1800 2800
rect 2200 2700 2300 2800
rect 2450 2700 2550 2800
rect 2700 2700 2800 2800
rect 3200 2700 3300 2800
rect 3450 2700 3550 2800
rect 3700 2700 3800 2800
rect 200 2450 300 2550
rect 450 2450 550 2550
rect 700 2450 800 2550
rect 950 2450 1050 2550
rect 1200 2450 1300 2550
rect 1450 2450 1550 2550
rect 1700 2450 1800 2550
rect 2200 2450 2300 2550
rect 2450 2450 2550 2550
rect 2700 2450 2800 2550
rect 2950 2450 3050 2550
rect 3200 2450 3300 2550
rect 3450 2450 3550 2550
rect 3700 2450 3800 2550
rect 200 2200 300 2300
rect 450 2200 550 2300
rect 700 2200 800 2300
rect 1200 2200 1300 2300
rect 1450 2200 1550 2300
rect 1700 2200 1800 2300
rect 2200 2200 2300 2300
rect 2450 2200 2550 2300
rect 2700 2200 2800 2300
rect 3200 2200 3300 2300
rect 3450 2200 3550 2300
rect 3700 2200 3800 2300
rect 200 1700 300 1800
rect 450 1700 550 1800
rect 700 1700 800 1800
rect 1200 1700 1300 1800
rect 1450 1700 1550 1800
rect 1700 1700 1800 1800
rect 2200 1700 2300 1800
rect 2450 1700 2550 1800
rect 2700 1700 2800 1800
rect 3200 1700 3300 1800
rect 3450 1700 3550 1800
rect 3700 1700 3800 1800
rect 200 1450 300 1550
rect 450 1450 550 1550
rect 700 1450 800 1550
rect 950 1450 1050 1550
rect 1200 1450 1300 1550
rect 1450 1450 1550 1550
rect 1700 1450 1800 1550
rect 2200 1450 2300 1550
rect 2450 1450 2550 1550
rect 2700 1450 2800 1550
rect 2950 1450 3050 1550
rect 3200 1450 3300 1550
rect 3450 1450 3550 1550
rect 3700 1450 3800 1550
rect 200 1200 300 1300
rect 450 1200 550 1300
rect 700 1200 800 1300
rect 1200 1200 1300 1300
rect 1450 1200 1550 1300
rect 1700 1200 1800 1300
rect 2200 1200 2300 1300
rect 2450 1200 2550 1300
rect 2700 1200 2800 1300
rect 3200 1200 3300 1300
rect 3450 1200 3550 1300
rect 3700 1200 3800 1300
rect 450 950 550 1050
rect 1450 950 1550 1050
rect 2450 950 2550 1050
rect 3450 950 3550 1050
rect 200 700 300 800
rect 450 700 550 800
rect 700 700 800 800
rect 1200 700 1300 800
rect 1450 700 1550 800
rect 1700 700 1800 800
rect 2200 700 2300 800
rect 2450 700 2550 800
rect 2700 700 2800 800
rect 3200 700 3300 800
rect 3450 700 3550 800
rect 3700 700 3800 800
rect 200 450 300 550
rect 450 450 550 550
rect 700 450 800 550
rect 950 450 1050 550
rect 1200 450 1300 550
rect 1450 450 1550 550
rect 1700 450 1800 550
rect 2200 450 2300 550
rect 2450 450 2550 550
rect 2700 450 2800 550
rect 2950 450 3050 550
rect 3200 450 3300 550
rect 3450 450 3550 550
rect 3700 450 3800 550
rect 200 200 300 300
rect 450 200 550 300
rect 700 200 800 300
rect 1200 200 1300 300
rect 1450 200 1550 300
rect 1700 200 1800 300
rect 2200 200 2300 300
rect 2450 200 2550 300
rect 2700 200 2800 300
rect 3200 200 3300 300
rect 3450 200 3550 300
rect 3700 200 3800 300
<< metal4 >>
rect 260 3820 740 4000
rect 1260 3820 1740 4000
rect 2260 3820 2740 4000
rect 3260 3820 3740 4000
rect 180 3800 820 3820
rect 180 3740 200 3800
rect 0 3700 200 3740
rect 300 3700 450 3800
rect 550 3700 700 3800
rect 800 3740 820 3800
rect 1180 3800 1820 3820
rect 1180 3740 1200 3800
rect 800 3700 1200 3740
rect 1300 3700 1450 3800
rect 1550 3700 1700 3800
rect 1800 3740 1820 3800
rect 2180 3800 2820 3820
rect 2180 3740 2200 3800
rect 1800 3700 2200 3740
rect 2300 3700 2450 3800
rect 2550 3700 2700 3800
rect 2800 3740 2820 3800
rect 3180 3800 3820 3820
rect 3180 3740 3200 3800
rect 2800 3700 3200 3740
rect 3300 3700 3450 3800
rect 3550 3700 3700 3800
rect 3800 3740 3820 3800
rect 3800 3700 4000 3740
rect 0 3550 4000 3700
rect 0 3450 200 3550
rect 300 3450 450 3550
rect 550 3450 700 3550
rect 800 3450 950 3550
rect 1050 3450 1200 3550
rect 1300 3450 1450 3550
rect 1550 3450 1700 3550
rect 1800 3450 2200 3550
rect 2300 3450 2450 3550
rect 2550 3450 2700 3550
rect 2800 3450 2950 3550
rect 3050 3450 3200 3550
rect 3300 3450 3450 3550
rect 3550 3450 3700 3550
rect 3800 3450 4000 3550
rect 0 3300 4000 3450
rect 0 3260 200 3300
rect 180 3200 200 3260
rect 300 3200 450 3300
rect 550 3200 700 3300
rect 800 3260 1200 3300
rect 800 3200 820 3260
rect 180 3180 820 3200
rect 1180 3200 1200 3260
rect 1300 3200 1450 3300
rect 1550 3200 1700 3300
rect 1800 3260 2200 3300
rect 1800 3200 1820 3260
rect 1180 3180 1820 3200
rect 2180 3200 2200 3260
rect 2300 3200 2450 3300
rect 2550 3200 2700 3300
rect 2800 3260 3200 3300
rect 2800 3200 2820 3260
rect 2180 3180 2820 3200
rect 3180 3200 3200 3260
rect 3300 3200 3450 3300
rect 3550 3200 3700 3300
rect 3800 3260 4000 3300
rect 3800 3200 3820 3260
rect 3180 3180 3820 3200
rect 260 3050 740 3180
rect 260 2950 450 3050
rect 550 2950 740 3050
rect 260 2820 740 2950
rect 1260 3050 1740 3180
rect 1260 2950 1450 3050
rect 1550 2950 1740 3050
rect 1260 2820 1740 2950
rect 2260 3050 2740 3180
rect 2260 2950 2450 3050
rect 2550 2950 2740 3050
rect 2260 2820 2740 2950
rect 3260 3050 3740 3180
rect 3260 2950 3450 3050
rect 3550 2950 3740 3050
rect 3260 2820 3740 2950
rect 180 2800 820 2820
rect 180 2740 200 2800
rect 0 2700 200 2740
rect 300 2700 450 2800
rect 550 2700 700 2800
rect 800 2740 820 2800
rect 1180 2800 1820 2820
rect 1180 2740 1200 2800
rect 800 2700 1200 2740
rect 1300 2700 1450 2800
rect 1550 2700 1700 2800
rect 1800 2740 1820 2800
rect 2180 2800 2820 2820
rect 2180 2740 2200 2800
rect 1800 2700 2200 2740
rect 2300 2700 2450 2800
rect 2550 2700 2700 2800
rect 2800 2740 2820 2800
rect 3180 2800 3820 2820
rect 3180 2740 3200 2800
rect 2800 2700 3200 2740
rect 3300 2700 3450 2800
rect 3550 2700 3700 2800
rect 3800 2740 3820 2800
rect 3800 2700 4000 2740
rect 0 2550 4000 2700
rect 0 2450 200 2550
rect 300 2450 450 2550
rect 550 2450 700 2550
rect 800 2450 950 2550
rect 1050 2450 1200 2550
rect 1300 2450 1450 2550
rect 1550 2450 1700 2550
rect 1800 2450 2200 2550
rect 2300 2450 2450 2550
rect 2550 2450 2700 2550
rect 2800 2450 2950 2550
rect 3050 2450 3200 2550
rect 3300 2450 3450 2550
rect 3550 2450 3700 2550
rect 3800 2450 4000 2550
rect 0 2300 4000 2450
rect 0 2260 200 2300
rect 180 2200 200 2260
rect 300 2200 450 2300
rect 550 2200 700 2300
rect 800 2260 1200 2300
rect 800 2200 820 2260
rect 180 2180 820 2200
rect 1180 2200 1200 2260
rect 1300 2200 1450 2300
rect 1550 2200 1700 2300
rect 1800 2260 2200 2300
rect 1800 2200 1820 2260
rect 1180 2180 1820 2200
rect 2180 2200 2200 2260
rect 2300 2200 2450 2300
rect 2550 2200 2700 2300
rect 2800 2260 3200 2300
rect 2800 2200 2820 2260
rect 2180 2180 2820 2200
rect 3180 2200 3200 2260
rect 3300 2200 3450 2300
rect 3550 2200 3700 2300
rect 3800 2260 4000 2300
rect 3800 2200 3820 2260
rect 3180 2180 3820 2200
rect 260 1820 740 2180
rect 1260 1820 1740 2180
rect 2260 1820 2740 2180
rect 3260 1820 3740 2180
rect 180 1800 820 1820
rect 180 1740 200 1800
rect 0 1700 200 1740
rect 300 1700 450 1800
rect 550 1700 700 1800
rect 800 1740 820 1800
rect 1180 1800 1820 1820
rect 1180 1740 1200 1800
rect 800 1700 1200 1740
rect 1300 1700 1450 1800
rect 1550 1700 1700 1800
rect 1800 1740 1820 1800
rect 2180 1800 2820 1820
rect 2180 1740 2200 1800
rect 1800 1700 2200 1740
rect 2300 1700 2450 1800
rect 2550 1700 2700 1800
rect 2800 1740 2820 1800
rect 3180 1800 3820 1820
rect 3180 1740 3200 1800
rect 2800 1700 3200 1740
rect 3300 1700 3450 1800
rect 3550 1700 3700 1800
rect 3800 1740 3820 1800
rect 3800 1700 4000 1740
rect 0 1550 4000 1700
rect 0 1450 200 1550
rect 300 1450 450 1550
rect 550 1450 700 1550
rect 800 1450 950 1550
rect 1050 1450 1200 1550
rect 1300 1450 1450 1550
rect 1550 1450 1700 1550
rect 1800 1450 2200 1550
rect 2300 1450 2450 1550
rect 2550 1450 2700 1550
rect 2800 1450 2950 1550
rect 3050 1450 3200 1550
rect 3300 1450 3450 1550
rect 3550 1450 3700 1550
rect 3800 1450 4000 1550
rect 0 1300 4000 1450
rect 0 1260 200 1300
rect 180 1200 200 1260
rect 300 1200 450 1300
rect 550 1200 700 1300
rect 800 1260 1200 1300
rect 800 1200 820 1260
rect 180 1180 820 1200
rect 1180 1200 1200 1260
rect 1300 1200 1450 1300
rect 1550 1200 1700 1300
rect 1800 1260 2200 1300
rect 1800 1200 1820 1260
rect 1180 1180 1820 1200
rect 2180 1200 2200 1260
rect 2300 1200 2450 1300
rect 2550 1200 2700 1300
rect 2800 1260 3200 1300
rect 2800 1200 2820 1260
rect 2180 1180 2820 1200
rect 3180 1200 3200 1260
rect 3300 1200 3450 1300
rect 3550 1200 3700 1300
rect 3800 1260 4000 1300
rect 3800 1200 3820 1260
rect 3180 1180 3820 1200
rect 260 1050 740 1180
rect 260 950 450 1050
rect 550 950 740 1050
rect 260 820 740 950
rect 1260 1050 1740 1180
rect 1260 950 1450 1050
rect 1550 950 1740 1050
rect 1260 820 1740 950
rect 2260 1050 2740 1180
rect 2260 950 2450 1050
rect 2550 950 2740 1050
rect 2260 820 2740 950
rect 3260 1050 3740 1180
rect 3260 950 3450 1050
rect 3550 950 3740 1050
rect 3260 820 3740 950
rect 180 800 820 820
rect 180 740 200 800
rect 0 700 200 740
rect 300 700 450 800
rect 550 700 700 800
rect 800 740 820 800
rect 1180 800 1820 820
rect 1180 740 1200 800
rect 800 700 1200 740
rect 1300 700 1450 800
rect 1550 700 1700 800
rect 1800 740 1820 800
rect 2180 800 2820 820
rect 2180 740 2200 800
rect 1800 700 2200 740
rect 2300 700 2450 800
rect 2550 700 2700 800
rect 2800 740 2820 800
rect 3180 800 3820 820
rect 3180 740 3200 800
rect 2800 700 3200 740
rect 3300 700 3450 800
rect 3550 700 3700 800
rect 3800 740 3820 800
rect 3800 700 4000 740
rect 0 550 4000 700
rect 0 450 200 550
rect 300 450 450 550
rect 550 450 700 550
rect 800 450 950 550
rect 1050 450 1200 550
rect 1300 450 1450 550
rect 1550 450 1700 550
rect 1800 450 2200 550
rect 2300 450 2450 550
rect 2550 450 2700 550
rect 2800 450 2950 550
rect 3050 450 3200 550
rect 3300 450 3450 550
rect 3550 450 3700 550
rect 3800 450 4000 550
rect 0 300 4000 450
rect 0 260 200 300
rect 180 200 200 260
rect 300 200 450 300
rect 550 200 700 300
rect 800 260 1200 300
rect 800 200 820 260
rect 180 180 820 200
rect 1180 200 1200 260
rect 1300 200 1450 300
rect 1550 200 1700 300
rect 1800 260 2200 300
rect 1800 200 1820 260
rect 1180 180 1820 200
rect 2180 200 2200 260
rect 2300 200 2450 300
rect 2550 200 2700 300
rect 2800 260 3200 300
rect 2800 200 2820 260
rect 2180 180 2820 200
rect 3180 200 3200 260
rect 3300 200 3450 300
rect 3550 200 3700 300
rect 3800 260 4000 300
rect 3800 200 3820 260
rect 3180 180 3820 200
rect 260 0 740 180
rect 1260 0 1740 180
rect 2260 0 2740 180
rect 3260 0 3740 180
<< end >>
