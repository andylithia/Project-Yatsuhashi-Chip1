magic
tech sky130B
magscale 1 2
timestamp 1661314321
<< metal4 >>
rect -35400 -22300 -26200 -22200
rect -35400 -27900 -30100 -22300
rect -26300 -27900 -26200 -22300
rect -35400 -28000 -26200 -27900
<< via4 >>
rect -30100 -27900 -26300 -22300
<< metal5 >>
tri -33442 -5000 -29442 -1000 se
rect -29442 -5000 -15358 -1000
tri -15358 -5000 -11358 -1000 sw
tri -35400 -6958 -33442 -5000 se
rect -33442 -5600 -28385 -5000
tri -28385 -5600 -27785 -5000 nw
tri -17015 -5600 -16415 -5000 ne
rect -16415 -5600 -11358 -5000
rect -33442 -6449 -29234 -5600
tri -29234 -6449 -28385 -5600 nw
tri -28385 -6449 -27536 -5600 se
rect -27536 -6449 -17264 -5600
tri -17264 -6449 -16415 -5600 sw
tri -16415 -6449 -15566 -5600 ne
rect -15566 -6449 -11358 -5600
rect -33442 -6958 -29951 -6449
tri -36457 -8015 -35400 -6958 se
rect -35400 -7166 -29951 -6958
tri -29951 -7166 -29234 -6449 nw
tri -29102 -7166 -28385 -6449 se
rect -28385 -7166 -16415 -6449
rect -35400 -8015 -30800 -7166
tri -30800 -8015 -29951 -7166 nw
tri -29951 -8015 -29102 -7166 se
rect -29102 -7298 -16415 -7166
tri -16415 -7298 -15566 -6449 sw
tri -15566 -7298 -14717 -6449 ne
rect -14717 -7298 -11358 -6449
rect -29102 -7902 -15566 -7298
tri -15566 -7902 -14962 -7298 sw
tri -14717 -7902 -14113 -7298 ne
rect -14113 -7902 -11358 -7298
rect -29102 -8015 -14962 -7902
tri -39400 -10958 -36457 -8015 se
rect -36457 -8864 -31649 -8015
tri -31649 -8864 -30800 -8015 nw
tri -30800 -8864 -29951 -8015 se
rect -29951 -8751 -14962 -8015
tri -14962 -8751 -14113 -7902 sw
tri -14113 -8751 -13264 -7902 ne
rect -13264 -8751 -11358 -7902
rect -29951 -8864 -14113 -8751
rect -36457 -9600 -32385 -8864
tri -32385 -9600 -31649 -8864 nw
tri -31536 -9600 -30800 -8864 se
rect -30800 -9600 -14113 -8864
tri -14113 -9600 -13264 -8751 sw
tri -13264 -9600 -12415 -8751 ne
rect -12415 -9600 -11358 -8751
tri -11358 -9600 -6758 -5000 sw
rect -36457 -10449 -33234 -9600
tri -33234 -10449 -32385 -9600 nw
tri -32385 -10449 -31536 -9600 se
rect -31536 -10449 -30800 -9600
rect -36457 -10958 -33936 -10449
rect -39400 -11151 -33936 -10958
tri -33936 -11151 -33234 -10449 nw
tri -33087 -11151 -32385 -10449 se
rect -32385 -11151 -30800 -10449
rect -39400 -12000 -34785 -11151
tri -34785 -12000 -33936 -11151 nw
tri -33936 -12000 -33087 -11151 se
rect -33087 -12000 -30800 -11151
rect -39400 -16000 -35400 -12000
tri -35400 -12615 -34785 -12000 nw
tri -34551 -12615 -33936 -12000 se
rect -33936 -12615 -30800 -12000
tri -34800 -12864 -34551 -12615 se
rect -34551 -12864 -30800 -12615
rect -34800 -29332 -30800 -12864
tri -30800 -14521 -25879 -9600 nw
tri -18921 -14521 -14000 -9600 ne
rect -14000 -10449 -13264 -9600
tri -13264 -10449 -12415 -9600 sw
tri -12415 -10449 -11566 -9600 ne
rect -11566 -10449 -6758 -9600
rect -14000 -11166 -12415 -10449
tri -12415 -11166 -11698 -10449 sw
tri -11566 -11166 -10849 -10449 ne
rect -10849 -10958 -6758 -10449
tri -6758 -10958 -5400 -9600 sw
rect -10849 -11166 -5400 -10958
rect -14000 -12015 -11698 -11166
tri -11698 -12015 -10849 -11166 sw
tri -10849 -12015 -10000 -11166 ne
rect -10000 -12015 -5400 -11166
rect -14000 -12864 -10849 -12015
tri -10849 -12864 -10000 -12015 sw
tri -10000 -12615 -9400 -12015 ne
rect -30200 -22300 -26200 -22200
rect -30200 -27900 -30100 -22300
rect -26300 -27900 -26200 -22300
rect -30200 -28484 -26200 -27900
tri -30800 -29332 -30200 -28732 sw
tri -30200 -29332 -29352 -28484 ne
rect -29352 -29332 -26200 -28484
rect -34800 -29552 -30200 -29332
tri -30200 -29552 -29980 -29332 sw
tri -29352 -29552 -29132 -29332 ne
rect -29132 -29552 -26200 -29332
rect -34800 -30389 -29980 -29552
tri -34800 -35000 -30189 -30389 ne
rect -30189 -30400 -29980 -30389
tri -29980 -30400 -29132 -29552 sw
tri -29132 -30400 -28284 -29552 ne
rect -28284 -30400 -26200 -29552
tri -26200 -30400 -22627 -26827 sw
tri -17573 -30400 -14000 -26827 se
rect -14000 -28484 -10000 -12864
rect -14000 -29332 -10848 -28484
tri -10848 -29332 -10000 -28484 nw
tri -10000 -29332 -9400 -28732 se
rect -9400 -29332 -5400 -12015
rect -14000 -29552 -11068 -29332
tri -11068 -29552 -10848 -29332 nw
tri -10220 -29552 -10000 -29332 se
rect -10000 -29552 -5400 -29332
rect -14000 -30400 -11916 -29552
tri -11916 -30400 -11068 -29552 nw
tri -11068 -30400 -10220 -29552 se
rect -10220 -30389 -5400 -29552
rect -10220 -30400 -10011 -30389
rect -30189 -31248 -29132 -30400
tri -29132 -31248 -28284 -30400 sw
tri -28284 -31248 -27436 -30400 ne
rect -27436 -31248 -12764 -30400
tri -12764 -31248 -11916 -30400 nw
tri -11916 -31248 -11068 -30400 se
rect -11068 -31248 -10011 -30400
rect -30189 -32096 -28284 -31248
tri -28284 -32096 -27436 -31248 sw
tri -27436 -32096 -26588 -31248 ne
rect -26588 -31636 -13152 -31248
tri -13152 -31636 -12764 -31248 nw
tri -12304 -31636 -11916 -31248 se
rect -11916 -31636 -10011 -31248
rect -26588 -32096 -14000 -31636
rect -30189 -32704 -27436 -32096
tri -27436 -32704 -26828 -32096 sw
tri -26588 -32704 -25980 -32096 ne
rect -25980 -32484 -14000 -32096
tri -14000 -32484 -13152 -31636 nw
tri -13152 -32484 -12304 -31636 se
rect -12304 -32484 -10011 -31636
rect -25980 -32704 -14848 -32484
rect -30189 -33552 -26828 -32704
tri -26828 -33552 -25980 -32704 sw
tri -25980 -33552 -25132 -32704 ne
rect -25132 -33332 -14848 -32704
tri -14848 -33332 -14000 -32484 nw
tri -14000 -33332 -13152 -32484 se
rect -13152 -33332 -10011 -32484
rect -25132 -33552 -15068 -33332
tri -15068 -33552 -14848 -33332 nw
tri -14220 -33552 -14000 -33332 se
rect -14000 -33552 -10011 -33332
rect -30189 -34400 -25980 -33552
tri -25980 -34400 -25132 -33552 sw
tri -25132 -34400 -24284 -33552 ne
rect -24284 -34400 -15916 -33552
tri -15916 -34400 -15068 -33552 nw
tri -15068 -34400 -14220 -33552 se
rect -14220 -34400 -10011 -33552
rect -30189 -35000 -25132 -34400
tri -25132 -35000 -24532 -34400 sw
tri -15668 -35000 -15068 -34400 se
rect -15068 -35000 -10011 -34400
tri -10011 -35000 -5400 -30389 nw
tri -30189 -39000 -26189 -35000 ne
rect -26189 -39000 -14011 -35000
tri -14011 -39000 -10011 -35000 nw
<< end >>
