magic
tech sky130A
timestamp 1659060853
<< metal1 >>
rect -1040 652 -1010 660
rect 870 652 900 660
rect -1040 552 -1003 652
rect -970 620 -780 630
rect -970 590 -960 620
rect -790 590 -780 620
rect -970 580 -780 590
rect -749 552 -720 652
rect -690 620 -490 630
rect -690 590 -680 620
rect -500 590 -490 620
rect -690 580 -490 590
rect -466 552 -437 652
rect -410 620 -210 630
rect -410 590 -400 620
rect -220 590 -210 620
rect -410 580 -210 590
rect -1040 55 -1010 552
rect -1040 -40 -1003 55
rect -980 20 -770 33
rect -980 -10 -970 20
rect -810 -10 -770 20
rect -980 -20 -770 -10
rect -749 -40 -720 55
rect -700 20 -490 30
rect -700 -10 -660 20
rect -520 -10 -490 20
rect -700 -20 -490 -10
rect -466 -40 -437 55
rect -410 20 -210 30
rect -410 -10 -380 20
rect -220 -10 -210 20
rect -410 -20 -210 -10
rect -183 -40 47 652
rect 70 620 270 630
rect 70 590 80 620
rect 260 590 270 620
rect 70 580 270 590
rect 301 552 330 652
rect 360 620 560 630
rect 360 590 370 620
rect 550 590 560 620
rect 360 580 560 590
rect 584 552 613 652
rect 640 620 840 630
rect 640 590 650 620
rect 830 590 840 620
rect 640 580 840 590
rect 867 552 900 652
rect 870 55 900 552
rect 70 20 270 30
rect 70 -10 80 20
rect 250 -10 270 20
rect 70 -20 270 -10
rect 301 -40 330 55
rect 360 20 560 30
rect 360 -10 380 20
rect 540 -10 560 20
rect 360 -20 560 -10
rect 584 -40 613 55
rect 640 20 840 30
rect 640 -10 660 20
rect 830 -10 840 20
rect 640 -20 840 -10
rect 867 -40 900 55
rect -1040 -60 900 -40
rect -1040 -120 -770 -60
rect -700 -120 -490 -60
rect -420 -120 280 -60
rect 350 -120 560 -60
rect 630 -120 900 -60
rect -1040 -130 900 -120
rect -130 -160 10 -130
<< via1 >>
rect -960 590 -790 620
rect -680 590 -500 620
rect -400 590 -220 620
rect -970 -10 -810 20
rect -660 -10 -520 20
rect -380 -10 -220 20
rect 80 590 260 620
rect 370 590 550 620
rect 650 590 830 620
rect 80 -10 250 20
rect 380 -10 540 20
rect 660 -10 830 20
rect -770 -120 -700 -60
rect -490 -120 -420 -60
rect 280 -120 350 -60
rect 560 -120 630 -60
<< metal2 >>
rect -970 620 -770 630
rect -970 590 -960 620
rect -780 590 -770 620
rect -970 580 -770 590
rect -690 620 -490 630
rect -690 590 -680 620
rect -500 590 -490 620
rect -690 580 -490 590
rect -410 620 -210 630
rect -410 590 -400 620
rect -220 590 -210 620
rect -410 580 -210 590
rect 70 620 270 630
rect 70 590 80 620
rect 260 590 270 620
rect 70 580 270 590
rect 360 620 560 630
rect 360 590 370 620
rect 550 590 560 620
rect 360 580 560 590
rect 640 620 840 630
rect 640 590 650 620
rect 830 590 840 620
rect 640 580 840 590
rect -780 40 -690 280
rect -500 40 -410 280
rect -196 55 16 291
rect 270 40 360 280
rect 550 50 640 280
rect 560 40 640 50
rect -980 20 -800 30
rect -980 -10 -970 20
rect -810 -10 -800 20
rect -980 -20 -800 -10
rect -770 -30 -700 40
rect -670 20 -510 30
rect -670 -10 -660 20
rect -520 -10 -510 20
rect -670 -20 -510 -10
rect -490 -30 -420 40
rect -390 20 -210 30
rect -390 -10 -380 20
rect -220 -10 -210 20
rect -390 -20 -210 -10
rect 70 20 260 30
rect 70 -10 80 20
rect 250 -10 260 20
rect 70 -20 260 -10
rect 280 -30 350 40
rect 370 20 550 30
rect 370 -10 380 20
rect 540 -10 550 20
rect 370 -20 550 -10
rect 570 -30 630 40
rect 650 20 840 30
rect 650 -10 660 20
rect 830 -10 840 20
rect 650 -20 840 -10
rect -780 -60 -690 -30
rect -780 -120 -770 -60
rect -700 -120 -690 -60
rect -780 -130 -690 -120
rect -500 -60 -410 -30
rect -500 -120 -490 -60
rect -420 -120 -410 -60
rect -500 -130 -410 -120
rect 270 -60 360 -30
rect 560 -40 630 -30
rect 270 -120 280 -60
rect 350 -120 360 -60
rect 270 -130 360 -120
rect 550 -60 640 -40
rect 550 -120 560 -60
rect 630 -120 640 -60
rect 550 -130 640 -120
<< via2 >>
rect -960 590 -790 620
rect -790 590 -780 620
rect -680 590 -500 620
rect -400 590 -220 620
rect 110 590 260 620
rect 370 590 550 620
rect 650 590 830 620
rect -240 330 -160 540
rect 20 330 100 540
rect -970 -10 -810 20
rect -660 -10 -520 20
rect -380 -10 -220 20
rect 80 -10 250 20
rect 380 -10 540 20
rect 660 -10 830 20
<< metal3 >>
rect -970 620 10 680
rect 100 670 840 680
rect 180 620 840 670
rect -970 590 -960 620
rect -780 590 -680 620
rect -500 590 -400 620
rect -220 590 10 620
rect 80 590 100 620
rect 260 590 370 620
rect 550 590 650 620
rect 830 590 840 620
rect -970 580 10 590
rect 100 580 840 590
rect -970 570 -290 580
rect -90 550 10 580
rect -250 540 -140 550
rect -250 330 -240 540
rect -160 330 -140 540
rect -250 320 -140 330
rect -90 540 110 550
rect -90 330 20 540
rect 100 330 110 540
rect -90 320 110 330
rect -980 30 -190 60
rect -90 30 10 320
rect -980 20 10 30
rect -980 -10 -970 20
rect -810 -10 -660 20
rect -520 -10 -380 20
rect -220 -10 10 20
rect -980 -50 10 -10
rect 70 20 860 50
rect 70 -10 80 20
rect 250 -10 380 20
rect 540 -10 660 20
rect 830 -10 860 20
rect 70 -40 100 -10
rect 180 -40 860 -10
rect 70 -50 860 -40
rect -280 -110 -180 -50
rect -280 -150 -270 -110
rect -190 -150 -180 -110
rect -280 -160 -180 -150
<< via3 >>
rect 100 620 180 670
rect 100 590 110 620
rect 110 590 180 620
rect -240 330 -160 540
rect 100 -10 180 20
rect 100 -40 180 -10
rect -270 -150 -190 -110
<< metal4 >>
rect -210 670 190 680
rect -210 590 100 670
rect 180 590 190 670
rect -210 580 190 590
rect -210 550 -90 580
rect -250 540 -90 550
rect -250 330 -240 540
rect -160 330 -90 540
rect -250 320 -90 330
rect -210 30 -90 320
rect -210 20 190 30
rect -210 -40 100 20
rect 180 -40 190 20
rect -210 -70 190 -40
rect -280 -110 -180 -100
rect -280 -150 -270 -110
rect -190 -150 -180 -110
rect -280 -160 -180 -150
rect 60 -160 160 -70
use sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_pr/mag
timestamp 1649977179
transform 1 0 0 0 1 0
box 0 0 348 607
use sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15_1
timestamp 1649977179
transform 1 0 283 0 1 0
box 0 0 348 607
use sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15_2
timestamp 1649977179
transform 1 0 566 0 1 0
box 0 0 348 607
use sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15_3
timestamp 1649977179
transform 1 0 -767 0 1 0
box 0 0 348 607
use sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15_4
timestamp 1649977179
transform 1 0 -1050 0 1 0
box 0 0 348 607
use sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aM04W5p00L0p15_5
timestamp 1649977179
transform 1 0 -484 0 1 0
box 0 0 348 607
<< labels >>
rlabel metal1 -130 -160 10 -130 1 SUB
rlabel metal4 60 -160 160 -130 1 G2
rlabel metal4 -280 -160 -180 -130 1 G1
<< end >>
