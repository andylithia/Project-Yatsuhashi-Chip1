** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/untitled-5.sch
**.subckt untitled-5
XM5 nop net5 GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=10
XM1 net1 net6 GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=10
Lload1 vsp net3 0.4n m=1
Lload2 net4 vsp 0.4n m=1
V1 net2 GND 0.9
I1 net2 net1 PULSE(0 10n 1n 10p 10p 1n 2)
R2 nop net6 3 m=1
R3 net5 net1 3 m=1
R1 net1 net3 1 m=1
I2 net2 vsp 10m
K1 Lload1 Lload2 0.9
R5 nop net1 200 m=1
R6 nop net4 1 m=1
C1 nop net1 100f m=1
C2 GND net1 10f m=1
C3 GND nop 10f m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice ff
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice



.subckt sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=2.828e+12p pd=2.132e+07u as=4.242e+12p
+ ps=3.198e+07u w=5.05e+06u l=150000u
X1 SOURCE SUBSTRATE SUBSTRATE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.03e+12p
+ ps=2.14e+07u w=5.05e+06u l=150000u
X2 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X5 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends
.options savecurrents
.tran 1ps 20ns
.control
run
display
plot v(nop)
plot v(nmid)
plot @I1[i]
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
