magic
tech sky130B
timestamp 1662232320
<< end >>
