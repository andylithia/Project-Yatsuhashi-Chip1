magic
tech sky130B
magscale 1 2
timestamp 1663446682
<< metal1 >>
rect 4270 40 4670 12480
rect 8870 40 9270 12480
rect 13470 40 13870 12480
<< metal2 >>
rect 0 12740 18000 13140
rect 0 12340 200 12740
rect 400 12340 600 12740
rect 800 12340 1000 12740
rect 1200 12340 1400 12740
rect 1600 12340 1800 12740
rect 2000 12340 2200 12740
rect 2400 12340 2600 12740
rect 2800 12340 3000 12740
rect 3200 12340 3400 12740
rect 3600 12340 3800 12740
rect 4000 12340 4200 12740
rect 4600 12340 4800 12740
rect 5000 12340 5200 12740
rect 5400 12340 5600 12740
rect 5800 12340 6000 12740
rect 6200 12340 6400 12740
rect 6600 12340 6800 12740
rect 7000 12340 7200 12740
rect 7400 12340 7600 12740
rect 7800 12340 8000 12740
rect 8200 12340 8400 12740
rect 8600 12340 8800 12740
rect 9200 12340 9400 12740
rect 9600 12340 9800 12740
rect 10000 12340 10200 12740
rect 10400 12340 10600 12740
rect 10800 12340 11000 12740
rect 11200 12340 11400 12740
rect 11600 12340 11800 12740
rect 12000 12340 12200 12740
rect 12400 12340 12600 12740
rect 12800 12340 13000 12740
rect 13200 12340 13400 12740
rect 13800 12340 14000 12740
rect 14200 12340 14400 12740
rect 14600 12340 14800 12740
rect 15000 12340 15200 12740
rect 15400 12340 15600 12740
rect 15800 12340 16000 12740
rect 16200 12340 16400 12740
rect 16600 12340 16800 12740
rect 17000 12340 17200 12740
rect 17400 12340 17600 12740
rect 17800 12340 18000 12740
rect 0 -200 200 200
rect 400 -200 600 200
rect 800 -200 1000 200
rect 1200 -200 1400 200
rect 1600 -200 1800 200
rect 2000 -200 2200 200
rect 2400 -200 2600 200
rect 2800 -200 3000 200
rect 3200 -200 3400 200
rect 3600 -200 3800 200
rect 4000 -200 4200 200
rect 4600 -200 4800 200
rect 5000 -200 5200 200
rect 5400 -200 5600 200
rect 5800 -200 6000 200
rect 6200 -200 6400 200
rect 6600 -200 6800 200
rect 7000 -200 7200 200
rect 7400 -200 7600 200
rect 7800 -200 8000 200
rect 8200 -200 8400 200
rect 8600 -200 8800 200
rect 9200 -200 9400 200
rect 9600 -200 9800 200
rect 10000 -200 10200 200
rect 10400 -200 10600 200
rect 10800 -200 11000 200
rect 11200 -200 11400 200
rect 11600 -200 11800 200
rect 12000 -200 12200 200
rect 12400 -200 12600 200
rect 12800 -200 13000 200
rect 13200 -200 13400 200
rect 13800 -200 14000 200
rect 14200 -200 14400 200
rect 14600 -200 14800 200
rect 15000 -200 15200 200
rect 15400 -200 15600 200
rect 15800 -200 16000 200
rect 16200 -200 16400 200
rect 16600 -200 16800 200
rect 17000 -200 17200 200
rect 17400 -200 17600 200
rect 17800 -200 18000 200
rect 0 -600 18000 -200
<< metal3 >>
rect 110 6470 150 12260
rect 4200 6600 4800 12000
rect 8800 6600 9400 12000
rect 13400 6600 14000 12000
rect 110 270 150 6060
rect 4200 400 4800 5800
rect 8800 400 9400 5800
rect 13400 400 14000 5800
use NMOS_50_0p5_25_1_alternative  NMOS_50_0p5_25_1_alternative_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/CLASSE
timestamp 1663444684
transform 1 0 65 0 1 65
box -65 -65 4283 12451
use NMOS_50_0p5_25_1_alternative  NMOS_50_0p5_25_1_alternative_1
timestamp 1663444684
transform 1 0 4665 0 1 65
box -65 -65 4283 12451
use NMOS_50_0p5_25_1_alternative  NMOS_50_0p5_25_1_alternative_2
timestamp 1663444684
transform 1 0 9265 0 1 65
box -65 -65 4283 12451
use NMOS_50_0p5_25_1_alternative  NMOS_50_0p5_25_1_alternative_3
timestamp 1663444684
transform 1 0 13865 0 1 65
box -65 -65 4283 12451
<< labels >>
rlabel metal2 0 12750 200 13140 1 G
rlabel metal3 110 6470 150 12260 1 SD1
rlabel metal3 110 270 150 6060 1 SD2
rlabel metal1 4420 60 4470 120 1 SUB
<< end >>
