magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< pwell >>
rect -26 -26 176 1026
<< scnmos >>
rect 60 0 90 1000
<< ndiff >>
rect 0 0 60 1000
rect 90 0 150 1000
<< poly >>
rect 60 1000 90 1026
rect 60 -26 90 0
<< locali >>
rect 8 467 42 533
rect 108 467 142 533
use sky130_sram_1r1w_24x128_8_contact_10  sky130_sram_1r1w_24x128_8_contact_10_0
timestamp 1661296025
transform 1 0 100 0 1 467
box -26 -22 76 88
use sky130_sram_1r1w_24x128_8_contact_10  sky130_sram_1r1w_24x128_8_contact_10_1
timestamp 1661296025
transform 1 0 0 0 1 467
box -26 -22 76 88
<< labels >>
rlabel poly s 75 500 75 500 4 G
port 1 nsew
rlabel locali s 25 500 25 500 4 S
port 2 nsew
rlabel locali s 125 500 125 500 4 D
port 3 nsew
<< properties >>
string FIXED_BBOX -25 -26 175 1026
<< end >>
