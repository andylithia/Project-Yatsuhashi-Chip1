** sch_path: /home/al/openmpw/Project-Yatsuhashi-Chip1/xschem/snh_clock_driver.sch
**.subckt snh_clock_driver vdd gnd CKIN CKN CKP CKOP CKON
*.iopin vdd
*.iopin gnd
*.ipin CKIN
*.opin CKN
*.opin CKP
*.opin CKOP
*.opin CKON
XC1 CKON CKN sky130_fd_pr__cap_mim_m3_1 W=10 L=5 MF=1 m=1
XC3 CKOP CKP sky130_fd_pr__cap_mim_m3_1 W=10 L=5 MF=1 m=1
x3 CKBUF gnd gnd vdd vdd CKP sky130_fd_sc_hd__clkinv_8
x2 CKBUF gnd gnd vdd vdd CKN sky130_fd_sc_hd__clkbuf_8
x1 net2 gnd gnd vdd vdd CKBUF sky130_fd_sc_hd__clkbuf_8
XM1 vdd CKON CKOP net1 sky130_fd_pr__nfet_03v3_nvt L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vdd CKOP CKON net1 sky130_fd_pr__nfet_03v3_nvt L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
x4 CKBUF gnd gnd vdd vdd CKP sky130_fd_sc_hd__clkinv_8
x5 CKBUF gnd gnd vdd vdd CKN sky130_fd_sc_hd__clkbuf_8
x6 CKIN gnd gnd vdd vdd net2 sky130_fd_sc_hd__clkbuf_2
**.ends
.end
