magic
tech sky130A
timestamp 1658607120
<< metal4 >>
rect 1700 -4400 2700 2000
rect 1700 -4600 1800 -4400
rect 2000 -4600 2100 -4400
rect 2300 -4600 2400 -4400
rect 2600 -4600 2700 -4400
rect 1700 -4700 2700 -4600
rect 1700 -4900 1800 -4700
rect 2000 -4900 2100 -4700
rect 2300 -4900 2400 -4700
rect 2600 -4900 2700 -4700
rect 1700 -5000 2700 -4900
rect 1700 -5200 1800 -5000
rect 2000 -5200 2100 -5000
rect 2300 -5200 2400 -5000
rect 2600 -5200 2700 -5000
rect 1700 -5300 2700 -5200
<< via4 >>
rect 1800 -4600 2000 -4400
rect 2100 -4600 2300 -4400
rect 2400 -4600 2600 -4400
rect 1800 -4900 2000 -4700
rect 2100 -4900 2300 -4700
rect 2400 -4900 2600 -4700
rect 1800 -5200 2000 -5000
rect 2100 -5200 2300 -5000
rect 2400 -5200 2600 -5000
<< metal5 >>
rect -2200 -100 13800 900
rect -2200 -1400 12500 -400
rect -2200 -14100 -1200 -1400
rect -900 -2700 11200 -1700
rect -900 -12800 100 -2700
rect 400 -4000 9900 -3000
rect 400 -11500 1400 -4000
rect 1700 -4400 2700 -4300
rect 1700 -4600 1800 -4400
rect 2000 -4600 2100 -4400
rect 2300 -4600 2400 -4400
rect 2600 -4600 2700 -4400
rect 1700 -4700 2700 -4600
rect 1700 -4900 1800 -4700
rect 2000 -4900 2100 -4700
rect 2300 -4900 2400 -4700
rect 2600 -4900 2700 -4700
rect 1700 -5000 2700 -4900
rect 1700 -5200 1800 -5000
rect 2000 -5200 2100 -5000
rect 2300 -5200 2400 -5000
rect 2600 -5200 2700 -5000
rect 1700 -10200 2700 -5200
rect 8900 -10200 9900 -4000
rect 1700 -11200 9900 -10200
rect 10200 -11500 11200 -2700
rect 400 -12500 11200 -11500
rect 11500 -12800 12500 -1400
rect -900 -13800 12500 -12800
rect 12800 -14100 13800 -100
rect -2200 -15100 13800 -14100
<< end >>
