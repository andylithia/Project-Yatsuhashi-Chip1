magic
tech sky130B
magscale 1 2
timestamp 1663980778
<< metal4 >>
rect -45500 -8112 -18500 -8000
rect -45500 -15888 -45388 -8112
rect -37612 -15888 -26388 -8112
rect -18612 -15888 -18500 -8112
rect -45500 -16000 -18500 -15888
<< via4 >>
rect -45388 -15888 -37612 -8112
rect -26388 -15888 -18612 -8112
<< metal5 >>
tri -25341 35728 -21069 40000 se
rect -21069 35728 12069 40000
tri 12069 35728 16341 40000 sw
tri -29069 32000 -25341 35728 se
rect -25341 32000 16341 35728
tri 16341 32000 20069 35728 sw
tri -36500 24569 -29069 32000 se
rect -29069 31000 -18755 32000
tri -18755 31000 -17755 32000 nw
tri 8755 31000 9755 32000 ne
rect 9755 31000 20069 32000
rect -29069 29586 -20169 31000
tri -20169 29586 -18755 31000 nw
tri -18755 29586 -17341 31000 se
rect -17341 29586 8341 31000
tri 8341 29586 9755 31000 sw
tri 9755 29586 11169 31000 ne
rect 11169 29586 20069 31000
rect -29069 28172 -21583 29586
tri -21583 28172 -20169 29586 nw
tri -20169 28172 -18755 29586 se
rect -18755 28172 9755 29586
tri 9755 28172 11169 29586 sw
tri 11169 28172 12583 29586 ne
rect 12583 28172 20069 29586
rect -29069 27242 -22513 28172
tri -22513 27242 -21583 28172 nw
tri -21099 27242 -20169 28172 se
rect -20169 27242 11169 28172
rect -29069 25828 -23927 27242
tri -23927 25828 -22513 27242 nw
tri -22513 25828 -21099 27242 se
rect -21099 26758 11169 27242
tri 11169 26758 12583 28172 sw
tri 12583 26758 13997 28172 ne
rect 13997 26758 20069 28172
rect -21099 25828 12583 26758
tri 12583 25828 13513 26758 sw
tri 13997 25828 14927 26758 ne
rect 14927 25828 20069 26758
rect -29069 24569 -25341 25828
tri -36655 24414 -36500 24569 se
rect -36500 24414 -25341 24569
tri -25341 24414 -23927 25828 nw
tri -23927 24414 -22513 25828 se
rect -22513 24414 13513 25828
tri 13513 24414 14927 25828 sw
tri 14927 24414 16341 25828 ne
rect 16341 24414 20069 25828
tri -44500 16569 -36655 24414 se
rect -36655 23000 -26755 24414
tri -26755 23000 -25341 24414 nw
tri -25341 23000 -23927 24414 se
rect -23927 23000 14927 24414
tri 14927 23000 16341 24414 sw
tri 16341 23000 17755 24414 ne
rect 17755 23000 20069 24414
rect -36655 21586 -28169 23000
tri -28169 21586 -26755 23000 nw
tri -26755 21586 -25341 23000 se
rect -25341 21586 -16186 23000
rect -36655 20172 -29583 21586
tri -29583 20172 -28169 21586 nw
tri -28169 20172 -26755 21586 se
rect -26755 20841 -16186 21586
tri -16186 20841 -14027 23000 nw
tri 5027 20841 7186 23000 ne
rect 7186 22255 16341 23000
tri 16341 22255 17086 23000 sw
tri 17755 22255 18500 23000 ne
rect 18500 22255 20069 23000
rect 7186 20841 17086 22255
tri 17086 20841 18500 22255 sw
tri 18500 20841 19914 22255 ne
rect 19914 20841 20069 22255
tri 20069 20841 31228 32000 sw
rect -26755 20172 -21027 20841
rect -36655 18828 -30927 20172
tri -30927 18828 -29583 20172 nw
tri -29513 18828 -28169 20172 se
rect -28169 18828 -21027 20172
rect -36655 17414 -32341 18828
tri -32341 17414 -30927 18828 nw
tri -30927 17414 -29513 18828 se
rect -29513 17414 -21027 18828
rect -36655 16569 -33755 17414
rect -44500 16000 -33755 16569
tri -33755 16000 -32341 17414 nw
tri -32341 16000 -30927 17414 se
rect -30927 16000 -21027 17414
tri -21027 16000 -16186 20841 nw
tri 7186 16000 12027 20841 ne
rect 12027 19427 18500 20841
tri 18500 19427 19914 20841 sw
tri 19914 19427 21328 20841 ne
rect 21328 19427 31228 20841
rect 12027 18013 19914 19427
tri 19914 18013 21328 19427 sw
tri 21328 18013 22742 19427 ne
rect 22742 18013 31228 19427
rect 12027 17083 21328 18013
tri 21328 17083 22258 18013 sw
tri 22742 17083 23672 18013 ne
rect 23672 17083 31228 18013
rect 12027 16000 22258 17083
rect -52500 14586 -35169 16000
tri -35169 14586 -33755 16000 nw
tri -33755 14586 -32341 16000 se
rect -32341 14586 -25341 16000
rect -52500 14255 -35500 14586
tri -35500 14255 -35169 14586 nw
tri -34086 14255 -33755 14586 se
rect -33755 14255 -25341 14586
rect -52500 8000 -36500 14255
tri -36500 13255 -35500 14255 nw
tri -35086 13255 -34086 14255 se
rect -34086 13255 -25341 14255
tri -35500 12841 -35086 13255 se
rect -35086 12841 -25341 13255
rect -35500 11686 -25341 12841
tri -25341 11686 -21027 16000 nw
tri 12027 11686 16341 16000 ne
rect 16341 15669 22258 16000
tri 22258 15669 23672 17083 sw
tri 23672 15669 25086 17083 ne
rect 25086 16569 31228 17083
tri 31228 16569 35500 20841 sw
rect 25086 15669 35500 16569
rect 16341 14255 23672 15669
tri 23672 14255 25086 15669 sw
tri 25086 14255 26500 15669 ne
rect 26500 14255 35500 15669
rect 16341 13255 25086 14255
tri 25086 13255 26086 14255 sw
tri 26500 13255 27500 14255 ne
rect 16341 12841 26086 13255
tri 26086 12841 26500 13255 sw
rect 16341 11686 26500 12841
rect -45500 -8112 -37500 -8000
rect -45500 -15888 -45388 -8112
rect -37612 -15888 -37500 -8112
rect -45500 -16000 -37500 -15888
rect -35500 -16891 -27500 11686
tri -27500 9527 -25341 11686 nw
tri 16341 9527 18500 11686 ne
rect -26500 -8112 -18500 -8000
rect -26500 -15888 -26388 -8112
rect -18612 -15888 -18500 -8112
tri -27500 -16891 -26500 -15891 sw
rect -26500 -16000 -18500 -15888
tri -25977 -16891 -25086 -16000 ne
rect -25086 -16891 -18500 -16000
rect -35500 -18305 -26500 -16891
tri -26500 -18305 -25086 -16891 sw
tri -25086 -18305 -23672 -16891 ne
rect -23672 -18305 -18500 -16891
rect -35500 -19205 -25086 -18305
tri -35500 -23000 -31705 -19205 ne
rect -31705 -19719 -25086 -19205
tri -25086 -19719 -23672 -18305 sw
tri -23672 -19719 -22258 -18305 ne
rect -22258 -19719 -18500 -18305
rect -31705 -20172 -23672 -19719
tri -23672 -20172 -23219 -19719 sw
tri -22258 -20172 -21805 -19719 ne
rect -21805 -20172 -18500 -19719
rect -31705 -21586 -23219 -20172
tri -23219 -21586 -21805 -20172 sw
tri -21805 -21586 -20391 -20172 ne
rect -20391 -21586 -18500 -20172
rect -31705 -23000 -21805 -21586
tri -21805 -23000 -20391 -21586 sw
tri -20391 -23000 -18977 -21586 ne
rect -18977 -23000 -18500 -21586
tri -18500 -23000 -7663 -12163 sw
tri 7663 -23000 18500 -12163 se
rect 18500 -15477 26500 11686
rect 18500 -15891 26086 -15477
tri 26086 -15891 26500 -15477 nw
rect 18500 -16891 25086 -15891
tri 25086 -16891 26086 -15891 nw
tri 26500 -16891 27500 -15891 se
rect 27500 -16891 35500 14255
rect 18500 -18305 23672 -16891
tri 23672 -18305 25086 -16891 nw
tri 25086 -18305 26500 -16891 se
rect 26500 -18305 35500 -16891
rect 18500 -19719 22258 -18305
tri 22258 -19719 23672 -18305 nw
tri 23672 -19719 25086 -18305 se
rect 25086 -19205 35500 -18305
rect 25086 -19719 29814 -19205
rect 18500 -20172 21805 -19719
tri 21805 -20172 22258 -19719 nw
tri 23219 -20172 23672 -19719 se
rect 23672 -20172 29814 -19719
rect 18500 -21586 20391 -20172
tri 20391 -21586 21805 -20172 nw
tri 21805 -21586 23219 -20172 se
rect 23219 -21586 29814 -20172
rect 18500 -23000 18977 -21586
tri 18977 -23000 20391 -21586 nw
tri 20391 -23000 21805 -21586 se
rect 21805 -23000 29814 -21586
tri -31705 -32000 -22705 -23000 ne
rect -22705 -24414 -20391 -23000
tri -20391 -24414 -18977 -23000 sw
tri -18977 -23477 -18500 -23000 ne
rect -18500 -23477 18500 -23000
tri 18500 -23477 18977 -23000 nw
tri 19914 -23477 20391 -23000 se
rect 20391 -23477 29814 -23000
tri -18500 -24414 -17563 -23477 ne
rect -17563 -24414 17086 -23477
rect -22705 -25828 -18977 -24414
tri -18977 -25828 -17563 -24414 sw
tri -17563 -25828 -16149 -24414 ne
rect -16149 -24891 17086 -24414
tri 17086 -24891 18500 -23477 nw
tri 18500 -24891 19914 -23477 se
rect 19914 -24891 29814 -23477
tri 29814 -24891 35500 -19205 nw
rect -16149 -25828 15672 -24891
rect -22705 -27242 -17563 -25828
tri -17563 -27242 -16149 -25828 sw
tri -16149 -27242 -14735 -25828 ne
rect -14735 -26305 15672 -25828
tri 15672 -26305 17086 -24891 nw
tri 17086 -26305 18500 -24891 se
rect 18500 -26305 27500 -24891
rect -14735 -27242 14258 -26305
rect -22705 -28172 -16149 -27242
tri -16149 -28172 -15219 -27242 sw
tri -14735 -28172 -13805 -27242 ne
rect -13805 -27719 14258 -27242
tri 14258 -27719 15672 -26305 nw
tri 15672 -27719 17086 -26305 se
rect 17086 -27205 27500 -26305
tri 27500 -27205 29814 -24891 nw
rect 17086 -27719 22705 -27205
rect -13805 -28172 13805 -27719
tri 13805 -28172 14258 -27719 nw
tri 15219 -28172 15672 -27719 se
rect 15672 -28172 22705 -27719
rect -22705 -29586 -15219 -28172
tri -15219 -29586 -13805 -28172 sw
tri -13805 -29586 -12391 -28172 ne
rect -12391 -29586 12391 -28172
tri 12391 -29586 13805 -28172 nw
tri 13805 -29586 15219 -28172 se
rect 15219 -29586 22705 -28172
rect -22705 -31000 -13805 -29586
tri -13805 -31000 -12391 -29586 sw
tri -12391 -31000 -10977 -29586 ne
rect -10977 -31000 10977 -29586
tri 10977 -31000 12391 -29586 nw
tri 12391 -31000 13805 -29586 se
rect 13805 -31000 22705 -29586
rect -22705 -32000 -12391 -31000
tri -12391 -32000 -11391 -31000 sw
tri 11391 -32000 12391 -31000 se
rect 12391 -32000 22705 -31000
tri 22705 -32000 27500 -27205 nw
tri -22705 -36205 -18500 -32000 ne
rect -18500 -36205 18500 -32000
tri 18500 -36205 22705 -32000 nw
tri -18500 -40000 -14705 -36205 ne
rect -14705 -40000 14705 -36205
tri 14705 -40000 18500 -36205 nw
<< end >>
