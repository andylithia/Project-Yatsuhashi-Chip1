magic
tech sky130A
timestamp 1658894606
use sky130_fd_pr__pfet_01v8_1um_10um_mult2  sky130_fd_pr__pfet_01v8_1um_10um_mult2_0
timestamp 1658894429
transform 1 0 0 0 1 0
box 0 0 539 1219
use sky130_fd_pr__pfet_01v8_1um_10um_mult2  sky130_fd_pr__pfet_01v8_1um_10um_mult2_1
timestamp 1658894429
transform 1 0 486 0 1 0
box 0 0 539 1219
use sky130_fd_pr__pfet_01v8_1um_10um_mult2  sky130_fd_pr__pfet_01v8_1um_10um_mult2_2
timestamp 1658894429
transform 1 0 972 0 1 0
box 0 0 539 1219
use sky130_fd_pr__pfet_01v8_1um_10um_mult2  sky130_fd_pr__pfet_01v8_1um_10um_mult2_3
timestamp 1658894429
transform 1 0 1458 0 1 0
box 0 0 539 1219
use sky130_fd_pr__pfet_01v8_1um_10um_mult2  sky130_fd_pr__pfet_01v8_1um_10um_mult2_4
timestamp 1658894429
transform 1 0 1944 0 1 0
box 0 0 539 1219
<< end >>
