magic
tech sky130B
magscale 1 2
timestamp 1659406861
<< metal4 >>
rect -39200 -16062 -36800 -15600
rect -39200 -17838 -38688 -16062
rect -36912 -17838 -36800 -16062
rect -39200 -18000 -36800 -17838
rect -39200 -22112 -31600 -21200
rect -39200 -23888 -33488 -22112
rect -31712 -23888 -31600 -22112
rect -39200 -24000 -31600 -23888
<< via4 >>
rect -38688 -17838 -36912 -16062
rect -33488 -23888 -31712 -22112
<< metal5 >>
tri -29472 -3423 -28549 -2500 se
rect -28549 -3423 -14051 -2500
tri -14051 -3423 -13128 -2500 sw
tri -30549 -4500 -29472 -3423 se
rect -29472 -4500 -13128 -3423
tri -13128 -4500 -12051 -3423 sw
tri -32301 -6252 -30549 -4500 se
rect -30549 -5100 -28320 -4500
tri -28320 -5100 -27720 -4500 nw
tri -14880 -5100 -14280 -4500 ne
rect -14280 -5100 -12051 -4500
rect -30549 -5948 -29168 -5100
tri -29168 -5948 -28320 -5100 nw
tri -28320 -5948 -27472 -5100 se
rect -27472 -5948 -15128 -5100
tri -15128 -5948 -14280 -5100 sw
tri -14280 -5948 -13432 -5100 ne
rect -13432 -5948 -12051 -5100
rect -30549 -6252 -29472 -5948
tri -29472 -6252 -29168 -5948 nw
tri -28624 -6252 -28320 -5948 se
rect -28320 -6252 -14280 -5948
tri -14280 -6252 -13976 -5948 sw
tri -13432 -6252 -13128 -5948 ne
rect -13128 -6252 -12051 -5948
tri -34200 -8151 -32301 -6252 se
rect -32301 -7100 -30320 -6252
tri -30320 -7100 -29472 -6252 nw
tri -29472 -7100 -28624 -6252 se
rect -28624 -7100 -13976 -6252
tri -13976 -7100 -13128 -6252 sw
tri -13128 -7100 -12280 -6252 ne
rect -12280 -7100 -12051 -6252
tri -12051 -7100 -9451 -4500 sw
rect -32301 -7948 -31168 -7100
tri -31168 -7948 -30320 -7100 nw
tri -30320 -7948 -29472 -7100 se
rect -29472 -7948 -28542 -7100
rect -32301 -8151 -31453 -7948
tri -35130 -9081 -34200 -8151 se
rect -34200 -8233 -31453 -8151
tri -31453 -8233 -31168 -7948 nw
tri -30605 -8233 -30320 -7948 se
rect -30320 -8233 -28542 -7948
rect -34200 -9081 -32301 -8233
tri -32301 -9081 -31453 -8233 nw
tri -31453 -9081 -30605 -8233 se
rect -30605 -8999 -28542 -8233
tri -28542 -8999 -26643 -7100 nw
tri -15957 -8999 -14058 -7100 ne
rect -14058 -7948 -13128 -7100
tri -13128 -7948 -12280 -7100 sw
tri -12280 -7948 -11432 -7100 ne
rect -11432 -7948 -9451 -7100
rect -14058 -8151 -12280 -7948
tri -12280 -8151 -12077 -7948 sw
tri -11432 -8151 -11229 -7948 ne
rect -11229 -8151 -9451 -7948
rect -14058 -8999 -12077 -8151
tri -12077 -8999 -11229 -8151 sw
tri -11229 -8999 -10381 -8151 ne
rect -10381 -8999 -9451 -8151
tri -9451 -8999 -7552 -7100 sw
rect -30605 -9081 -29472 -8999
tri -36800 -10751 -35130 -9081 se
rect -35130 -9929 -33149 -9081
tri -33149 -9929 -32301 -9081 nw
tri -32301 -9929 -31453 -9081 se
rect -31453 -9929 -29472 -9081
tri -29472 -9929 -28542 -8999 nw
tri -14058 -9929 -13128 -8999 ne
rect -13128 -9847 -11229 -8999
tri -11229 -9847 -10381 -8999 sw
tri -10381 -9847 -9533 -8999 ne
rect -9533 -9847 -7552 -8999
rect -13128 -9929 -10381 -9847
rect -35130 -10751 -33997 -9929
tri -37029 -10980 -36800 -10751 se
rect -36800 -10777 -33997 -10751
tri -33997 -10777 -33149 -9929 nw
tri -33149 -10777 -32301 -9929 se
rect -32301 -10777 -31371 -9929
rect -36800 -10980 -34200 -10777
tri -34200 -10980 -33997 -10777 nw
tri -33352 -10980 -33149 -10777 se
rect -33149 -10980 -31371 -10777
tri -38800 -12751 -37029 -10980 se
rect -37029 -11828 -35048 -10980
tri -35048 -11828 -34200 -10980 nw
tri -34200 -11828 -33352 -10980 se
rect -33352 -11828 -31371 -10980
tri -31371 -11828 -29472 -9929 nw
tri -13128 -11828 -11229 -9929 ne
rect -11229 -10132 -10381 -9929
tri -10381 -10132 -10096 -9847 sw
tri -9533 -10132 -9248 -9847 ne
rect -9248 -10132 -7552 -9847
rect -11229 -10980 -10096 -10132
tri -10096 -10980 -9248 -10132 sw
tri -9248 -10980 -8400 -10132 ne
rect -8400 -10980 -7552 -10132
rect -11229 -11828 -9248 -10980
tri -9248 -11828 -8400 -10980 sw
tri -8400 -11828 -7552 -10980 ne
tri -7552 -11828 -4723 -8999 sw
rect -37029 -12676 -35896 -11828
tri -35896 -12676 -35048 -11828 nw
tri -35048 -12676 -34200 -11828 se
rect -34200 -12676 -32301 -11828
rect -37029 -12751 -35978 -12676
rect -38800 -12758 -35978 -12751
tri -35978 -12758 -35896 -12676 nw
tri -35130 -12758 -35048 -12676 se
rect -35048 -12758 -32301 -12676
tri -32301 -12758 -31371 -11828 nw
tri -11229 -12758 -10299 -11828 ne
rect -10299 -12676 -8400 -11828
tri -8400 -12676 -7552 -11828 sw
tri -7552 -12676 -6704 -11828 ne
rect -6704 -12676 -4723 -11828
rect -10299 -12758 -7552 -12676
rect -38800 -12980 -36200 -12758
tri -36200 -12980 -35978 -12758 nw
tri -35352 -12980 -35130 -12758 se
rect -35130 -12980 -34200 -12758
rect -38800 -16062 -36800 -12980
tri -36800 -13580 -36200 -12980 nw
tri -35952 -13580 -35352 -12980 se
rect -35352 -13580 -34200 -12980
rect -38800 -17838 -38688 -16062
rect -36912 -17838 -36800 -16062
rect -38800 -17950 -36800 -17838
tri -36200 -13828 -35952 -13580 se
rect -35952 -13828 -34200 -13580
rect -36200 -27782 -34200 -13828
tri -34200 -14657 -32301 -12758 nw
tri -10299 -14657 -8400 -12758 ne
rect -8400 -12980 -7552 -12758
tri -7552 -12980 -7248 -12676 sw
tri -6704 -12980 -6400 -12676 ne
rect -6400 -12751 -4723 -12676
tri -4723 -12751 -3800 -11828 sw
rect -6400 -12980 -3800 -12751
rect -8400 -13580 -7248 -12980
tri -7248 -13580 -6648 -12980 sw
tri -6400 -13580 -5800 -12980 ne
rect -8400 -13828 -6648 -13580
tri -6648 -13828 -6400 -13580 sw
rect -33600 -22112 -31600 -22000
rect -33600 -23888 -33488 -22112
rect -31712 -23888 -31600 -22112
rect -33600 -26933 -31600 -23888
tri -33600 -27182 -33351 -26933 ne
rect -33351 -27182 -31600 -26933
tri -34200 -27782 -33600 -27182 sw
tri -33351 -27782 -32751 -27182 ne
rect -32751 -27782 -31600 -27182
rect -36200 -28010 -33600 -27782
tri -36200 -28933 -35277 -28010 ne
rect -35277 -28084 -33600 -28010
tri -33600 -28084 -33298 -27782 sw
tri -32751 -28084 -32449 -27782 ne
rect -32449 -28084 -31600 -27782
rect -35277 -28933 -33298 -28084
tri -33298 -28933 -32449 -28084 sw
tri -32449 -28933 -31600 -28084 ne
tri -31600 -28933 -28772 -26105 sw
tri -9539 -27244 -8400 -26105 se
rect -8400 -26933 -6400 -13828
rect -8400 -27182 -6649 -26933
tri -6649 -27182 -6400 -26933 nw
rect -8400 -27244 -6711 -27182
tri -6711 -27244 -6649 -27182 nw
tri -5862 -27244 -5800 -27182 se
rect -5800 -27244 -3800 -12980
tri -11228 -28933 -9539 -27244 se
rect -9539 -27782 -7249 -27244
tri -7249 -27782 -6711 -27244 nw
tri -6400 -27782 -5862 -27244 se
rect -5862 -27782 -3800 -27244
rect -9539 -28084 -7551 -27782
tri -7551 -28084 -7249 -27782 nw
tri -6702 -28084 -6400 -27782 se
rect -6400 -28010 -3800 -27782
rect -6400 -28084 -5572 -28010
rect -9539 -28933 -8400 -28084
tri -8400 -28933 -7551 -28084 nw
tri -7551 -28933 -6702 -28084 se
rect -6702 -28933 -5572 -28084
tri -35277 -31761 -32449 -28933 ne
tri -32449 -29782 -31600 -28933 sw
tri -31600 -29782 -30751 -28933 ne
rect -30751 -29782 -28772 -28933
rect -32449 -30631 -31600 -29782
tri -31600 -30631 -30751 -29782 sw
tri -30751 -30631 -29902 -29782 ne
rect -29902 -30631 -28772 -29782
rect -32449 -30912 -30751 -30631
tri -30751 -30912 -30470 -30631 sw
tri -29902 -30912 -29621 -30631 ne
rect -29621 -30912 -28772 -30631
rect -32449 -31761 -30470 -30912
tri -30470 -31761 -29621 -30912 sw
tri -29621 -31761 -28772 -30912 ne
tri -28772 -31761 -25944 -28933 sw
tri -12367 -30072 -11228 -28933 se
rect -11228 -29782 -9249 -28933
tri -9249 -29782 -8400 -28933 nw
tri -8400 -29782 -7551 -28933 se
rect -7551 -29782 -5572 -28933
tri -5572 -29782 -3800 -28010 nw
rect -11228 -30072 -9539 -29782
tri -9539 -30072 -9249 -29782 nw
tri -8690 -30072 -8400 -29782 se
rect -8400 -30010 -5800 -29782
tri -5800 -30010 -5572 -29782 nw
rect -8400 -30072 -6711 -30010
tri -14056 -31761 -12367 -30072 se
rect -12367 -30921 -10388 -30072
tri -10388 -30921 -9539 -30072 nw
tri -9539 -30921 -8690 -30072 se
rect -8690 -30921 -6711 -30072
tri -6711 -30921 -5800 -30010 nw
rect -12367 -31761 -11237 -30921
tri -32449 -32900 -31310 -31761 ne
rect -31310 -32610 -29621 -31761
tri -29621 -32610 -28772 -31761 sw
tri -28772 -32610 -27923 -31761 ne
rect -27923 -32610 -25944 -31761
rect -31310 -32900 -28772 -32610
tri -28772 -32900 -28482 -32610 sw
tri -27923 -32900 -27633 -32610 ne
rect -27633 -32900 -25944 -32610
tri -25944 -32900 -24805 -31761 sw
tri -15195 -32900 -14056 -31761 se
rect -14056 -31770 -11237 -31761
tri -11237 -31770 -10388 -30921 nw
tri -10388 -31770 -9539 -30921 se
rect -9539 -31770 -8400 -30921
rect -14056 -32051 -11518 -31770
tri -11518 -32051 -11237 -31770 nw
tri -10669 -32051 -10388 -31770 se
rect -10388 -32051 -8400 -31770
rect -14056 -32900 -12367 -32051
tri -12367 -32900 -11518 -32051 nw
tri -11518 -32900 -10669 -32051 se
rect -10669 -32610 -8400 -32051
tri -8400 -32610 -6711 -30921 nw
rect -10669 -32900 -9539 -32610
tri -31310 -35500 -28710 -32900 ne
rect -28710 -33749 -28482 -32900
tri -28482 -33749 -27633 -32900 sw
tri -27633 -33749 -26784 -32900 ne
rect -26784 -33749 -13216 -32900
tri -13216 -33749 -12367 -32900 nw
tri -12367 -33749 -11518 -32900 se
rect -11518 -33749 -9539 -32900
tri -9539 -33749 -8400 -32610 nw
rect -28710 -34051 -27633 -33749
tri -27633 -34051 -27331 -33749 sw
tri -26784 -34051 -26482 -33749 ne
rect -26482 -34051 -13518 -33749
tri -13518 -34051 -13216 -33749 nw
tri -12669 -34051 -12367 -33749 se
rect -12367 -34051 -11290 -33749
rect -28710 -34900 -27331 -34051
tri -27331 -34900 -26482 -34051 sw
tri -26482 -34900 -25633 -34051 ne
rect -25633 -34900 -14367 -34051
tri -14367 -34900 -13518 -34051 nw
tri -13518 -34900 -12669 -34051 se
rect -12669 -34900 -11290 -34051
rect -28710 -35500 -26482 -34900
tri -26482 -35500 -25882 -34900 sw
tri -14118 -35500 -13518 -34900 se
rect -13518 -35500 -11290 -34900
tri -11290 -35500 -9539 -33749 nw
tri -28710 -36577 -27633 -35500 ne
rect -27633 -36577 -12367 -35500
tri -12367 -36577 -11290 -35500 nw
tri -27633 -37500 -26710 -36577 ne
rect -26710 -37500 -13290 -36577
tri -13290 -37500 -12367 -36577 nw
<< end >>
