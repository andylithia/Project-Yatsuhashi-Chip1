** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/untitled.sch
**.subckt untitled
V1 vin GND dc 0 ac 1
R1 vmid vin 1k m=1
R2 vmid GND 1k m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.control
ac dec 10 1 10K
plot V(vmid) V(vin)

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
