magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< locali >>
rect 4021 25182 4967 25216
rect 6284 25143 6861 25177
rect 4341 25070 4857 25104
rect 4661 24980 4967 25014
rect 4661 24756 4967 24790
rect 4341 24666 4857 24700
rect 6284 24593 6861 24627
rect 3941 24554 4967 24588
rect 3861 24392 4967 24426
rect 6284 24353 6861 24387
rect 4341 24280 4857 24314
rect 4661 24190 4967 24224
rect 4661 23966 4967 24000
rect 4341 23876 4857 23910
rect 6284 23803 6861 23837
rect 3781 23764 4967 23798
rect 4021 23602 4967 23636
rect 6284 23563 6861 23597
rect 4261 23490 4857 23524
rect 4661 23400 4967 23434
rect 4661 23176 4967 23210
rect 4261 23086 4857 23120
rect 6284 23013 6861 23047
rect 3941 22974 4967 23008
rect 3861 22812 4967 22846
rect 6284 22773 6861 22807
rect 4261 22700 4857 22734
rect 4661 22610 4967 22644
rect 4661 22386 4967 22420
rect 4261 22296 4857 22330
rect 6284 22223 6861 22257
rect 3781 22184 4967 22218
rect 4021 22022 4967 22056
rect 6284 21983 6861 22017
rect 4181 21910 4857 21944
rect 4661 21820 4967 21854
rect 4661 21596 4967 21630
rect 4181 21506 4857 21540
rect 6284 21433 6861 21467
rect 3941 21394 4967 21428
rect 3861 21232 4967 21266
rect 6284 21193 6861 21227
rect 4181 21120 4857 21154
rect 4661 21030 4967 21064
rect 4661 20806 4967 20840
rect 4181 20716 4857 20750
rect 6284 20643 6861 20677
rect 3781 20604 4967 20638
rect 4021 20442 4967 20476
rect 6284 20403 6861 20437
rect 4101 20330 4857 20364
rect 4661 20240 4967 20274
rect 4661 20016 4967 20050
rect 4101 19926 4857 19960
rect 6284 19853 6861 19887
rect 3941 19814 4967 19848
rect 3861 19652 4967 19686
rect 6284 19613 6861 19647
rect 4101 19540 4857 19574
rect 4661 19450 4967 19484
rect 4661 19226 4967 19260
rect 4101 19136 4857 19170
rect 6284 19063 6861 19097
rect 3781 19024 4967 19058
rect 4021 18862 4967 18896
rect 6284 18823 6861 18857
rect 4341 18750 4857 18784
rect 4581 18660 4967 18694
rect 4581 18436 4967 18470
rect 4341 18346 4857 18380
rect 6284 18273 6861 18307
rect 3941 18234 4967 18268
rect 3861 18072 4967 18106
rect 6284 18033 6861 18067
rect 4341 17960 4857 17994
rect 4581 17870 4967 17904
rect 4581 17646 4967 17680
rect 4341 17556 4857 17590
rect 6284 17483 6861 17517
rect 3781 17444 4967 17478
rect 4021 17282 4967 17316
rect 6284 17243 6861 17277
rect 4261 17170 4857 17204
rect 4581 17080 4967 17114
rect 4581 16856 4967 16890
rect 4261 16766 4857 16800
rect 6284 16693 6861 16727
rect 3941 16654 4967 16688
rect 3861 16492 4967 16526
rect 6284 16453 6861 16487
rect 4261 16380 4857 16414
rect 4581 16290 4967 16324
rect 4581 16066 4967 16100
rect 4261 15976 4857 16010
rect 6284 15903 6861 15937
rect 3781 15864 4967 15898
rect 4021 15702 4967 15736
rect 6284 15663 6861 15697
rect 4181 15590 4857 15624
rect 4581 15500 4967 15534
rect 4581 15276 4967 15310
rect 4181 15186 4857 15220
rect 6284 15113 6861 15147
rect 3941 15074 4967 15108
rect 3861 14912 4967 14946
rect 6284 14873 6861 14907
rect 4181 14800 4857 14834
rect 4581 14710 4967 14744
rect 4581 14486 4967 14520
rect 4181 14396 4857 14430
rect 6284 14323 6861 14357
rect 3781 14284 4967 14318
rect 4021 14122 4967 14156
rect 6284 14083 6861 14117
rect 4101 14010 4857 14044
rect 4581 13920 4967 13954
rect 4581 13696 4967 13730
rect 4101 13606 4857 13640
rect 6284 13533 6861 13567
rect 3941 13494 4967 13528
rect 3861 13332 4967 13366
rect 6284 13293 6861 13327
rect 4101 13220 4857 13254
rect 4581 13130 4967 13164
rect 4581 12906 4967 12940
rect 4101 12816 4857 12850
rect 6284 12743 6861 12777
rect 3781 12704 4967 12738
rect 4021 12542 4967 12576
rect 6284 12503 6861 12537
rect 4341 12430 4857 12464
rect 4501 12340 4967 12374
rect 4501 12116 4967 12150
rect 4341 12026 4857 12060
rect 6284 11953 6861 11987
rect 3941 11914 4967 11948
rect 3861 11752 4967 11786
rect 6284 11713 6861 11747
rect 4341 11640 4857 11674
rect 4501 11550 4967 11584
rect 4501 11326 4967 11360
rect 4341 11236 4857 11270
rect 6284 11163 6861 11197
rect 3781 11124 4967 11158
rect 4021 10962 4967 10996
rect 6284 10923 6861 10957
rect 4261 10850 4857 10884
rect 4501 10760 4967 10794
rect 4501 10536 4967 10570
rect 4261 10446 4857 10480
rect 6284 10373 6861 10407
rect 3941 10334 4967 10368
rect 3861 10172 4967 10206
rect 6284 10133 6861 10167
rect 4261 10060 4857 10094
rect 4501 9970 4967 10004
rect 4501 9746 4967 9780
rect 4261 9656 4857 9690
rect 6284 9583 6861 9617
rect 3781 9544 4967 9578
rect 4021 9382 4967 9416
rect 6284 9343 6861 9377
rect 4181 9270 4857 9304
rect 4501 9180 4967 9214
rect 4501 8956 4967 8990
rect 4181 8866 4857 8900
rect 6284 8793 6861 8827
rect 3941 8754 4967 8788
rect 3861 8592 4967 8626
rect 6284 8553 6861 8587
rect 4181 8480 4857 8514
rect 4501 8390 4967 8424
rect 4501 8166 4967 8200
rect 4181 8076 4857 8110
rect 6284 8003 6861 8037
rect 3781 7964 4967 7998
rect 4021 7802 4967 7836
rect 6284 7763 6861 7797
rect 4101 7690 4857 7724
rect 4501 7600 4967 7634
rect 4501 7376 4967 7410
rect 4101 7286 4857 7320
rect 6284 7213 6861 7247
rect 3941 7174 4967 7208
rect 3861 7012 4967 7046
rect 6284 6973 6861 7007
rect 4101 6900 4857 6934
rect 4501 6810 4967 6844
rect 4501 6586 4967 6620
rect 4101 6496 4857 6530
rect 6284 6423 6861 6457
rect 3781 6384 4967 6418
rect 4021 6222 4967 6256
rect 6284 6183 6861 6217
rect 4341 6110 4857 6144
rect 4421 6020 4967 6054
rect 4421 5796 4967 5830
rect 4341 5706 4857 5740
rect 6284 5633 6861 5667
rect 3941 5594 4967 5628
rect 3861 5432 4967 5466
rect 6284 5393 6861 5427
rect 433 5343 701 5377
rect 4341 5320 4857 5354
rect 4421 5230 4967 5264
rect 4421 5006 4967 5040
rect 353 4893 621 4927
rect 4341 4916 4857 4950
rect 6284 4843 6861 4877
rect 3781 4804 4967 4838
rect 4021 4642 4967 4676
rect 6284 4603 6861 4637
rect 4261 4530 4857 4564
rect 4421 4440 4967 4474
rect 4421 4216 4967 4250
rect 4261 4126 4857 4160
rect 6284 4053 6861 4087
rect 3941 4014 4967 4048
rect 3861 3852 4967 3886
rect 6284 3813 6861 3847
rect 4261 3740 4857 3774
rect 4421 3650 4967 3684
rect 4421 3426 4967 3460
rect 4261 3336 4857 3370
rect 6284 3263 6861 3297
rect 3781 3224 4967 3258
rect 4021 3062 4967 3096
rect 6284 3023 6861 3057
rect 273 2973 701 3007
rect 4181 2950 4857 2984
rect 4421 2860 4967 2894
rect 4421 2636 4967 2670
rect 193 2523 621 2557
rect 4181 2546 4857 2580
rect 6284 2473 6861 2507
rect 3941 2434 4967 2468
rect 3861 2272 4967 2306
rect 6284 2233 6861 2267
rect 4181 2160 4857 2194
rect 4421 2070 4967 2104
rect 4421 1846 4967 1880
rect 4181 1756 4857 1790
rect 6284 1683 6861 1717
rect 3781 1644 4967 1678
rect 4021 1482 4967 1516
rect 6284 1443 6861 1477
rect 4101 1370 4857 1404
rect 4421 1280 4967 1314
rect 4421 1056 4967 1090
rect 4101 966 4857 1000
rect 6284 893 6861 927
rect 3941 854 4967 888
rect 3861 692 4967 726
rect 6284 653 6861 687
rect 113 603 701 637
rect 4101 580 4857 614
rect 4421 490 4967 524
rect 4421 266 4967 300
rect 33 153 621 187
rect 4101 176 4857 210
rect 6284 103 6861 137
rect 3781 64 4967 98
<< metal1 >>
rect 19 0 47 6320
rect 99 0 127 6320
rect 179 0 207 6320
rect 259 0 287 6320
rect 339 0 367 6320
rect 419 0 447 6320
rect 3655 6174 3719 6226
rect 3655 5624 3719 5676
rect 3655 5384 3719 5436
rect 3655 4834 3719 4886
rect 3655 3804 3719 3856
rect 3655 3254 3719 3306
rect 3655 3014 3719 3066
rect 3655 2464 3719 2516
rect 3655 1434 3719 1486
rect 3655 884 3719 936
rect 3655 644 3719 696
rect 3767 241 3795 25308
rect 3847 427 3875 25308
rect 3927 1031 3955 25308
rect 4007 1217 4035 25308
rect 4087 2402 4115 25308
rect 4167 2797 4195 25308
rect 4247 3192 4275 25308
rect 4327 3587 4355 25308
rect 4407 4772 4435 25308
rect 4487 5167 4515 25308
rect 4567 5562 4595 25308
rect 4647 5957 4675 25308
rect 5023 25045 5087 25097
rect 5495 25045 5559 25097
rect 5927 25045 5991 25097
rect 6271 25056 6335 25108
rect 6695 25056 6759 25108
rect 5023 24673 5087 24725
rect 5495 24673 5559 24725
rect 5927 24673 5991 24725
rect 6271 24662 6335 24714
rect 6695 24662 6759 24714
rect 5023 24255 5087 24307
rect 5495 24255 5559 24307
rect 5927 24255 5991 24307
rect 6271 24266 6335 24318
rect 6695 24266 6759 24318
rect 5023 23883 5087 23935
rect 5495 23883 5559 23935
rect 5927 23883 5991 23935
rect 6271 23872 6335 23924
rect 6695 23872 6759 23924
rect 5023 23465 5087 23517
rect 5495 23465 5559 23517
rect 5927 23465 5991 23517
rect 6271 23476 6335 23528
rect 6695 23476 6759 23528
rect 5023 23093 5087 23145
rect 5495 23093 5559 23145
rect 5927 23093 5991 23145
rect 6271 23082 6335 23134
rect 6695 23082 6759 23134
rect 5023 22675 5087 22727
rect 5495 22675 5559 22727
rect 5927 22675 5991 22727
rect 6271 22686 6335 22738
rect 6695 22686 6759 22738
rect 5023 22303 5087 22355
rect 5495 22303 5559 22355
rect 5927 22303 5991 22355
rect 6271 22292 6335 22344
rect 6695 22292 6759 22344
rect 5023 21885 5087 21937
rect 5495 21885 5559 21937
rect 5927 21885 5991 21937
rect 6271 21896 6335 21948
rect 6695 21896 6759 21948
rect 5023 21513 5087 21565
rect 5495 21513 5559 21565
rect 5927 21513 5991 21565
rect 6271 21502 6335 21554
rect 6695 21502 6759 21554
rect 5023 21095 5087 21147
rect 5495 21095 5559 21147
rect 5927 21095 5991 21147
rect 6271 21106 6335 21158
rect 6695 21106 6759 21158
rect 5023 20723 5087 20775
rect 5495 20723 5559 20775
rect 5927 20723 5991 20775
rect 6271 20712 6335 20764
rect 6695 20712 6759 20764
rect 5023 20305 5087 20357
rect 5495 20305 5559 20357
rect 5927 20305 5991 20357
rect 6271 20316 6335 20368
rect 6695 20316 6759 20368
rect 5023 19933 5087 19985
rect 5495 19933 5559 19985
rect 5927 19933 5991 19985
rect 6271 19922 6335 19974
rect 6695 19922 6759 19974
rect 5023 19515 5087 19567
rect 5495 19515 5559 19567
rect 5927 19515 5991 19567
rect 6271 19526 6335 19578
rect 6695 19526 6759 19578
rect 5023 19143 5087 19195
rect 5495 19143 5559 19195
rect 5927 19143 5991 19195
rect 6271 19132 6335 19184
rect 6695 19132 6759 19184
rect 5023 18725 5087 18777
rect 5495 18725 5559 18777
rect 5927 18725 5991 18777
rect 6271 18736 6335 18788
rect 6695 18736 6759 18788
rect 5023 18353 5087 18405
rect 5495 18353 5559 18405
rect 5927 18353 5991 18405
rect 6271 18342 6335 18394
rect 6695 18342 6759 18394
rect 5023 17935 5087 17987
rect 5495 17935 5559 17987
rect 5927 17935 5991 17987
rect 6271 17946 6335 17998
rect 6695 17946 6759 17998
rect 5023 17563 5087 17615
rect 5495 17563 5559 17615
rect 5927 17563 5991 17615
rect 6271 17552 6335 17604
rect 6695 17552 6759 17604
rect 5023 17145 5087 17197
rect 5495 17145 5559 17197
rect 5927 17145 5991 17197
rect 6271 17156 6335 17208
rect 6695 17156 6759 17208
rect 5023 16773 5087 16825
rect 5495 16773 5559 16825
rect 5927 16773 5991 16825
rect 6271 16762 6335 16814
rect 6695 16762 6759 16814
rect 5023 16355 5087 16407
rect 5495 16355 5559 16407
rect 5927 16355 5991 16407
rect 6271 16366 6335 16418
rect 6695 16366 6759 16418
rect 5023 15983 5087 16035
rect 5495 15983 5559 16035
rect 5927 15983 5991 16035
rect 6271 15972 6335 16024
rect 6695 15972 6759 16024
rect 5023 15565 5087 15617
rect 5495 15565 5559 15617
rect 5927 15565 5991 15617
rect 6271 15576 6335 15628
rect 6695 15576 6759 15628
rect 5023 15193 5087 15245
rect 5495 15193 5559 15245
rect 5927 15193 5991 15245
rect 6271 15182 6335 15234
rect 6695 15182 6759 15234
rect 5023 14775 5087 14827
rect 5495 14775 5559 14827
rect 5927 14775 5991 14827
rect 6271 14786 6335 14838
rect 6695 14786 6759 14838
rect 5023 14403 5087 14455
rect 5495 14403 5559 14455
rect 5927 14403 5991 14455
rect 6271 14392 6335 14444
rect 6695 14392 6759 14444
rect 5023 13985 5087 14037
rect 5495 13985 5559 14037
rect 5927 13985 5991 14037
rect 6271 13996 6335 14048
rect 6695 13996 6759 14048
rect 5023 13613 5087 13665
rect 5495 13613 5559 13665
rect 5927 13613 5991 13665
rect 6271 13602 6335 13654
rect 6695 13602 6759 13654
rect 5023 13195 5087 13247
rect 5495 13195 5559 13247
rect 5927 13195 5991 13247
rect 6271 13206 6335 13258
rect 6695 13206 6759 13258
rect 5023 12823 5087 12875
rect 5495 12823 5559 12875
rect 5927 12823 5991 12875
rect 6271 12812 6335 12864
rect 6695 12812 6759 12864
rect 5023 12405 5087 12457
rect 5495 12405 5559 12457
rect 5927 12405 5991 12457
rect 6271 12416 6335 12468
rect 6695 12416 6759 12468
rect 5023 12033 5087 12085
rect 5495 12033 5559 12085
rect 5927 12033 5991 12085
rect 6271 12022 6335 12074
rect 6695 12022 6759 12074
rect 5023 11615 5087 11667
rect 5495 11615 5559 11667
rect 5927 11615 5991 11667
rect 6271 11626 6335 11678
rect 6695 11626 6759 11678
rect 5023 11243 5087 11295
rect 5495 11243 5559 11295
rect 5927 11243 5991 11295
rect 6271 11232 6335 11284
rect 6695 11232 6759 11284
rect 5023 10825 5087 10877
rect 5495 10825 5559 10877
rect 5927 10825 5991 10877
rect 6271 10836 6335 10888
rect 6695 10836 6759 10888
rect 5023 10453 5087 10505
rect 5495 10453 5559 10505
rect 5927 10453 5991 10505
rect 6271 10442 6335 10494
rect 6695 10442 6759 10494
rect 5023 10035 5087 10087
rect 5495 10035 5559 10087
rect 5927 10035 5991 10087
rect 6271 10046 6335 10098
rect 6695 10046 6759 10098
rect 5023 9663 5087 9715
rect 5495 9663 5559 9715
rect 5927 9663 5991 9715
rect 6271 9652 6335 9704
rect 6695 9652 6759 9704
rect 5023 9245 5087 9297
rect 5495 9245 5559 9297
rect 5927 9245 5991 9297
rect 6271 9256 6335 9308
rect 6695 9256 6759 9308
rect 5023 8873 5087 8925
rect 5495 8873 5559 8925
rect 5927 8873 5991 8925
rect 6271 8862 6335 8914
rect 6695 8862 6759 8914
rect 5023 8455 5087 8507
rect 5495 8455 5559 8507
rect 5927 8455 5991 8507
rect 6271 8466 6335 8518
rect 6695 8466 6759 8518
rect 5023 8083 5087 8135
rect 5495 8083 5559 8135
rect 5927 8083 5991 8135
rect 6271 8072 6335 8124
rect 6695 8072 6759 8124
rect 5023 7665 5087 7717
rect 5495 7665 5559 7717
rect 5927 7665 5991 7717
rect 6271 7676 6335 7728
rect 6695 7676 6759 7728
rect 5023 7293 5087 7345
rect 5495 7293 5559 7345
rect 5927 7293 5991 7345
rect 6271 7282 6335 7334
rect 6695 7282 6759 7334
rect 5023 6875 5087 6927
rect 5495 6875 5559 6927
rect 5927 6875 5991 6927
rect 6271 6886 6335 6938
rect 6695 6886 6759 6938
rect 5023 6503 5087 6555
rect 5495 6503 5559 6555
rect 5927 6503 5991 6555
rect 6271 6492 6335 6544
rect 6695 6492 6759 6544
rect 5023 6085 5087 6137
rect 5495 6085 5559 6137
rect 5927 6085 5991 6137
rect 6271 6096 6335 6148
rect 6695 6096 6759 6148
rect 4635 5893 4687 5957
rect 4555 5498 4607 5562
rect 4475 5103 4527 5167
rect 4395 4708 4447 4772
rect 4315 3523 4367 3587
rect 4235 3128 4287 3192
rect 4155 2733 4207 2797
rect 4075 2338 4127 2402
rect 3995 1153 4047 1217
rect 3915 967 3967 1031
rect 3835 363 3887 427
rect 3755 177 3807 241
rect 3655 94 3719 146
rect 3767 0 3795 177
rect 3847 0 3875 363
rect 3927 0 3955 967
rect 4007 0 4035 1153
rect 4087 0 4115 2338
rect 4167 0 4195 2733
rect 4247 0 4275 3128
rect 4327 0 4355 3523
rect 4407 0 4435 4708
rect 4487 0 4515 5103
rect 4567 0 4595 5498
rect 4647 0 4675 5893
rect 5023 5713 5087 5765
rect 5495 5713 5559 5765
rect 5927 5713 5991 5765
rect 6271 5702 6335 5754
rect 6695 5702 6759 5754
rect 5023 5295 5087 5347
rect 5495 5295 5559 5347
rect 5927 5295 5991 5347
rect 6271 5306 6335 5358
rect 6695 5306 6759 5358
rect 5023 4923 5087 4975
rect 5495 4923 5559 4975
rect 5927 4923 5991 4975
rect 6271 4912 6335 4964
rect 6695 4912 6759 4964
rect 5023 4505 5087 4557
rect 5495 4505 5559 4557
rect 5927 4505 5991 4557
rect 6271 4516 6335 4568
rect 6695 4516 6759 4568
rect 5023 4133 5087 4185
rect 5495 4133 5559 4185
rect 5927 4133 5991 4185
rect 6271 4122 6335 4174
rect 6695 4122 6759 4174
rect 5023 3715 5087 3767
rect 5495 3715 5559 3767
rect 5927 3715 5991 3767
rect 6271 3726 6335 3778
rect 6695 3726 6759 3778
rect 5023 3343 5087 3395
rect 5495 3343 5559 3395
rect 5927 3343 5991 3395
rect 6271 3332 6335 3384
rect 6695 3332 6759 3384
rect 5023 2925 5087 2977
rect 5495 2925 5559 2977
rect 5927 2925 5991 2977
rect 6271 2936 6335 2988
rect 6695 2936 6759 2988
rect 5023 2553 5087 2605
rect 5495 2553 5559 2605
rect 5927 2553 5991 2605
rect 6271 2542 6335 2594
rect 6695 2542 6759 2594
rect 5023 2135 5087 2187
rect 5495 2135 5559 2187
rect 5927 2135 5991 2187
rect 6271 2146 6335 2198
rect 6695 2146 6759 2198
rect 5023 1763 5087 1815
rect 5495 1763 5559 1815
rect 5927 1763 5991 1815
rect 6271 1752 6335 1804
rect 6695 1752 6759 1804
rect 5023 1345 5087 1397
rect 5495 1345 5559 1397
rect 5927 1345 5991 1397
rect 6271 1356 6335 1408
rect 6695 1356 6759 1408
rect 5023 973 5087 1025
rect 5495 973 5559 1025
rect 5927 973 5991 1025
rect 6271 962 6335 1014
rect 6695 962 6759 1014
rect 5023 555 5087 607
rect 5495 555 5559 607
rect 5927 555 5991 607
rect 6271 566 6335 618
rect 6695 566 6759 618
rect 5023 183 5087 235
rect 5495 183 5559 235
rect 5927 183 5991 235
rect 6271 172 6335 224
rect 6695 172 6759 224
<< metal2 >>
rect 5027 25047 5083 25095
rect 5499 25047 5555 25095
rect 5931 25047 5987 25095
rect 6275 25058 6331 25106
rect 6699 25058 6755 25106
rect 5027 24675 5083 24723
rect 5499 24675 5555 24723
rect 5931 24675 5987 24723
rect 6275 24663 6331 24711
rect 6699 24663 6755 24711
rect 5027 24257 5083 24305
rect 5499 24257 5555 24305
rect 5931 24257 5987 24305
rect 6275 24268 6331 24316
rect 6699 24268 6755 24316
rect 5027 23885 5083 23933
rect 5499 23885 5555 23933
rect 5931 23885 5987 23933
rect 6275 23873 6331 23921
rect 6699 23873 6755 23921
rect 5027 23467 5083 23515
rect 5499 23467 5555 23515
rect 5931 23467 5987 23515
rect 6275 23478 6331 23526
rect 6699 23478 6755 23526
rect 5027 23095 5083 23143
rect 5499 23095 5555 23143
rect 5931 23095 5987 23143
rect 6275 23083 6331 23131
rect 6699 23083 6755 23131
rect 5027 22677 5083 22725
rect 5499 22677 5555 22725
rect 5931 22677 5987 22725
rect 6275 22688 6331 22736
rect 6699 22688 6755 22736
rect 5027 22305 5083 22353
rect 5499 22305 5555 22353
rect 5931 22305 5987 22353
rect 6275 22293 6331 22341
rect 6699 22293 6755 22341
rect 5027 21887 5083 21935
rect 5499 21887 5555 21935
rect 5931 21887 5987 21935
rect 6275 21898 6331 21946
rect 6699 21898 6755 21946
rect 5027 21515 5083 21563
rect 5499 21515 5555 21563
rect 5931 21515 5987 21563
rect 6275 21503 6331 21551
rect 6699 21503 6755 21551
rect 5027 21097 5083 21145
rect 5499 21097 5555 21145
rect 5931 21097 5987 21145
rect 6275 21108 6331 21156
rect 6699 21108 6755 21156
rect 5027 20725 5083 20773
rect 5499 20725 5555 20773
rect 5931 20725 5987 20773
rect 6275 20713 6331 20761
rect 6699 20713 6755 20761
rect 5027 20307 5083 20355
rect 5499 20307 5555 20355
rect 5931 20307 5987 20355
rect 6275 20318 6331 20366
rect 6699 20318 6755 20366
rect 5027 19935 5083 19983
rect 5499 19935 5555 19983
rect 5931 19935 5987 19983
rect 6275 19923 6331 19971
rect 6699 19923 6755 19971
rect 5027 19517 5083 19565
rect 5499 19517 5555 19565
rect 5931 19517 5987 19565
rect 6275 19528 6331 19576
rect 6699 19528 6755 19576
rect 5027 19145 5083 19193
rect 5499 19145 5555 19193
rect 5931 19145 5987 19193
rect 6275 19133 6331 19181
rect 6699 19133 6755 19181
rect 5027 18727 5083 18775
rect 5499 18727 5555 18775
rect 5931 18727 5987 18775
rect 6275 18738 6331 18786
rect 6699 18738 6755 18786
rect 5027 18355 5083 18403
rect 5499 18355 5555 18403
rect 5931 18355 5987 18403
rect 6275 18343 6331 18391
rect 6699 18343 6755 18391
rect 5027 17937 5083 17985
rect 5499 17937 5555 17985
rect 5931 17937 5987 17985
rect 6275 17948 6331 17996
rect 6699 17948 6755 17996
rect 5027 17565 5083 17613
rect 5499 17565 5555 17613
rect 5931 17565 5987 17613
rect 6275 17553 6331 17601
rect 6699 17553 6755 17601
rect 5027 17147 5083 17195
rect 5499 17147 5555 17195
rect 5931 17147 5987 17195
rect 6275 17158 6331 17206
rect 6699 17158 6755 17206
rect 5027 16775 5083 16823
rect 5499 16775 5555 16823
rect 5931 16775 5987 16823
rect 6275 16763 6331 16811
rect 6699 16763 6755 16811
rect 5027 16357 5083 16405
rect 5499 16357 5555 16405
rect 5931 16357 5987 16405
rect 6275 16368 6331 16416
rect 6699 16368 6755 16416
rect 5027 15985 5083 16033
rect 5499 15985 5555 16033
rect 5931 15985 5987 16033
rect 6275 15973 6331 16021
rect 6699 15973 6755 16021
rect 5027 15567 5083 15615
rect 5499 15567 5555 15615
rect 5931 15567 5987 15615
rect 6275 15578 6331 15626
rect 6699 15578 6755 15626
rect 5027 15195 5083 15243
rect 5499 15195 5555 15243
rect 5931 15195 5987 15243
rect 6275 15183 6331 15231
rect 6699 15183 6755 15231
rect 5027 14777 5083 14825
rect 5499 14777 5555 14825
rect 5931 14777 5987 14825
rect 6275 14788 6331 14836
rect 6699 14788 6755 14836
rect 5027 14405 5083 14453
rect 5499 14405 5555 14453
rect 5931 14405 5987 14453
rect 6275 14393 6331 14441
rect 6699 14393 6755 14441
rect 5027 13987 5083 14035
rect 5499 13987 5555 14035
rect 5931 13987 5987 14035
rect 6275 13998 6331 14046
rect 6699 13998 6755 14046
rect 5027 13615 5083 13663
rect 5499 13615 5555 13663
rect 5931 13615 5987 13663
rect 6275 13603 6331 13651
rect 6699 13603 6755 13651
rect 5027 13197 5083 13245
rect 5499 13197 5555 13245
rect 5931 13197 5987 13245
rect 6275 13208 6331 13256
rect 6699 13208 6755 13256
rect 5027 12825 5083 12873
rect 5499 12825 5555 12873
rect 5931 12825 5987 12873
rect 6275 12813 6331 12861
rect 6699 12813 6755 12861
rect 5027 12407 5083 12455
rect 5499 12407 5555 12455
rect 5931 12407 5987 12455
rect 6275 12418 6331 12466
rect 6699 12418 6755 12466
rect 5027 12035 5083 12083
rect 5499 12035 5555 12083
rect 5931 12035 5987 12083
rect 6275 12023 6331 12071
rect 6699 12023 6755 12071
rect 5027 11617 5083 11665
rect 5499 11617 5555 11665
rect 5931 11617 5987 11665
rect 6275 11628 6331 11676
rect 6699 11628 6755 11676
rect 5027 11245 5083 11293
rect 5499 11245 5555 11293
rect 5931 11245 5987 11293
rect 6275 11233 6331 11281
rect 6699 11233 6755 11281
rect 5027 10827 5083 10875
rect 5499 10827 5555 10875
rect 5931 10827 5987 10875
rect 6275 10838 6331 10886
rect 6699 10838 6755 10886
rect 5027 10455 5083 10503
rect 5499 10455 5555 10503
rect 5931 10455 5987 10503
rect 6275 10443 6331 10491
rect 6699 10443 6755 10491
rect 5027 10037 5083 10085
rect 5499 10037 5555 10085
rect 5931 10037 5987 10085
rect 6275 10048 6331 10096
rect 6699 10048 6755 10096
rect 5027 9665 5083 9713
rect 5499 9665 5555 9713
rect 5931 9665 5987 9713
rect 6275 9653 6331 9701
rect 6699 9653 6755 9701
rect 5027 9247 5083 9295
rect 5499 9247 5555 9295
rect 5931 9247 5987 9295
rect 6275 9258 6331 9306
rect 6699 9258 6755 9306
rect 5027 8875 5083 8923
rect 5499 8875 5555 8923
rect 5931 8875 5987 8923
rect 6275 8863 6331 8911
rect 6699 8863 6755 8911
rect 5027 8457 5083 8505
rect 5499 8457 5555 8505
rect 5931 8457 5987 8505
rect 6275 8468 6331 8516
rect 6699 8468 6755 8516
rect 5027 8085 5083 8133
rect 5499 8085 5555 8133
rect 5931 8085 5987 8133
rect 6275 8073 6331 8121
rect 6699 8073 6755 8121
rect 5027 7667 5083 7715
rect 5499 7667 5555 7715
rect 5931 7667 5987 7715
rect 6275 7678 6331 7726
rect 6699 7678 6755 7726
rect 5027 7295 5083 7343
rect 5499 7295 5555 7343
rect 5931 7295 5987 7343
rect 6275 7283 6331 7331
rect 6699 7283 6755 7331
rect 5027 6877 5083 6925
rect 5499 6877 5555 6925
rect 5931 6877 5987 6925
rect 6275 6888 6331 6936
rect 6699 6888 6755 6936
rect 5027 6505 5083 6553
rect 5499 6505 5555 6553
rect 5931 6505 5987 6553
rect 6275 6493 6331 6541
rect 6699 6493 6755 6541
rect 3673 5939 3701 6200
rect 5027 6087 5083 6135
rect 5499 6087 5555 6135
rect 5931 6087 5987 6135
rect 6275 6098 6331 6146
rect 6699 6098 6755 6146
rect 3673 5911 4661 5939
rect 5027 5715 5083 5763
rect 5499 5715 5555 5763
rect 5931 5715 5987 5763
rect 6275 5703 6331 5751
rect 6699 5703 6755 5751
rect 3673 5544 3701 5650
rect 3673 5516 4581 5544
rect 3673 5149 3701 5410
rect 5027 5297 5083 5345
rect 5499 5297 5555 5345
rect 5931 5297 5987 5345
rect 6275 5308 6331 5356
rect 6699 5308 6755 5356
rect 3673 5121 4501 5149
rect 5027 4925 5083 4973
rect 5499 4925 5555 4973
rect 5931 4925 5987 4973
rect 6275 4913 6331 4961
rect 6699 4913 6755 4961
rect 3673 4754 3701 4860
rect 3673 4726 4421 4754
rect 5027 4507 5083 4555
rect 5499 4507 5555 4555
rect 5931 4507 5987 4555
rect 6275 4518 6331 4566
rect 6699 4518 6755 4566
rect 5027 4135 5083 4183
rect 5499 4135 5555 4183
rect 5931 4135 5987 4183
rect 6275 4123 6331 4171
rect 6699 4123 6755 4171
rect 3673 3569 3701 3830
rect 5027 3717 5083 3765
rect 5499 3717 5555 3765
rect 5931 3717 5987 3765
rect 6275 3728 6331 3776
rect 6699 3728 6755 3776
rect 3673 3541 4341 3569
rect 5027 3345 5083 3393
rect 5499 3345 5555 3393
rect 5931 3345 5987 3393
rect 6275 3333 6331 3381
rect 6699 3333 6755 3381
rect 3673 3174 3701 3280
rect 3673 3146 4261 3174
rect 3673 2779 3701 3040
rect 5027 2927 5083 2975
rect 5499 2927 5555 2975
rect 5931 2927 5987 2975
rect 6275 2938 6331 2986
rect 6699 2938 6755 2986
rect 3673 2751 4181 2779
rect 5027 2555 5083 2603
rect 5499 2555 5555 2603
rect 5931 2555 5987 2603
rect 6275 2543 6331 2591
rect 6699 2543 6755 2591
rect 3673 2384 3701 2490
rect 3673 2356 4101 2384
rect 5027 2137 5083 2185
rect 5499 2137 5555 2185
rect 5931 2137 5987 2185
rect 6275 2148 6331 2196
rect 6699 2148 6755 2196
rect 5027 1765 5083 1813
rect 5499 1765 5555 1813
rect 5931 1765 5987 1813
rect 6275 1753 6331 1801
rect 6699 1753 6755 1801
rect 3673 1199 3701 1460
rect 5027 1347 5083 1395
rect 5499 1347 5555 1395
rect 5931 1347 5987 1395
rect 6275 1358 6331 1406
rect 6699 1358 6755 1406
rect 3673 1171 4021 1199
rect 3673 985 3941 1013
rect 3673 910 3701 985
rect 5027 975 5083 1023
rect 5499 975 5555 1023
rect 5931 975 5987 1023
rect 6275 963 6331 1011
rect 6699 963 6755 1011
rect 3673 409 3701 670
rect 5027 557 5083 605
rect 5499 557 5555 605
rect 5931 557 5987 605
rect 6275 568 6331 616
rect 6699 568 6755 616
rect 3673 381 3861 409
rect 3673 195 3781 223
rect 3673 120 3701 195
rect 5027 185 5083 233
rect 5499 185 5555 233
rect 5931 185 5987 233
rect 6275 173 6331 221
rect 6699 173 6755 221
<< metal3 >>
rect 4980 25039 5130 25103
rect 5452 25039 5602 25103
rect 5884 25039 6034 25103
rect 6228 25050 6378 25114
rect 6652 25050 6802 25114
rect 4980 24667 5130 24731
rect 5452 24667 5602 24731
rect 5884 24667 6034 24731
rect 6228 24656 6378 24720
rect 6652 24656 6802 24720
rect 4980 24249 5130 24313
rect 5452 24249 5602 24313
rect 5884 24249 6034 24313
rect 6228 24260 6378 24324
rect 6652 24260 6802 24324
rect 4980 23877 5130 23941
rect 5452 23877 5602 23941
rect 5884 23877 6034 23941
rect 6228 23866 6378 23930
rect 6652 23866 6802 23930
rect 4980 23459 5130 23523
rect 5452 23459 5602 23523
rect 5884 23459 6034 23523
rect 6228 23470 6378 23534
rect 6652 23470 6802 23534
rect 4980 23087 5130 23151
rect 5452 23087 5602 23151
rect 5884 23087 6034 23151
rect 6228 23076 6378 23140
rect 6652 23076 6802 23140
rect 4980 22669 5130 22733
rect 5452 22669 5602 22733
rect 5884 22669 6034 22733
rect 6228 22680 6378 22744
rect 6652 22680 6802 22744
rect 4980 22297 5130 22361
rect 5452 22297 5602 22361
rect 5884 22297 6034 22361
rect 6228 22286 6378 22350
rect 6652 22286 6802 22350
rect 4980 21879 5130 21943
rect 5452 21879 5602 21943
rect 5884 21879 6034 21943
rect 6228 21890 6378 21954
rect 6652 21890 6802 21954
rect 4980 21507 5130 21571
rect 5452 21507 5602 21571
rect 5884 21507 6034 21571
rect 6228 21496 6378 21560
rect 6652 21496 6802 21560
rect 4980 21089 5130 21153
rect 5452 21089 5602 21153
rect 5884 21089 6034 21153
rect 6228 21100 6378 21164
rect 6652 21100 6802 21164
rect 4980 20717 5130 20781
rect 5452 20717 5602 20781
rect 5884 20717 6034 20781
rect 6228 20706 6378 20770
rect 6652 20706 6802 20770
rect 4980 20299 5130 20363
rect 5452 20299 5602 20363
rect 5884 20299 6034 20363
rect 6228 20310 6378 20374
rect 6652 20310 6802 20374
rect 4980 19927 5130 19991
rect 5452 19927 5602 19991
rect 5884 19927 6034 19991
rect 6228 19916 6378 19980
rect 6652 19916 6802 19980
rect 4980 19509 5130 19573
rect 5452 19509 5602 19573
rect 5884 19509 6034 19573
rect 6228 19520 6378 19584
rect 6652 19520 6802 19584
rect 4980 19137 5130 19201
rect 5452 19137 5602 19201
rect 5884 19137 6034 19201
rect 6228 19126 6378 19190
rect 6652 19126 6802 19190
rect 4980 18719 5130 18783
rect 5452 18719 5602 18783
rect 5884 18719 6034 18783
rect 6228 18730 6378 18794
rect 6652 18730 6802 18794
rect 4980 18347 5130 18411
rect 5452 18347 5602 18411
rect 5884 18347 6034 18411
rect 6228 18336 6378 18400
rect 6652 18336 6802 18400
rect 4980 17929 5130 17993
rect 5452 17929 5602 17993
rect 5884 17929 6034 17993
rect 6228 17940 6378 18004
rect 6652 17940 6802 18004
rect 4980 17557 5130 17621
rect 5452 17557 5602 17621
rect 5884 17557 6034 17621
rect 6228 17546 6378 17610
rect 6652 17546 6802 17610
rect 4980 17139 5130 17203
rect 5452 17139 5602 17203
rect 5884 17139 6034 17203
rect 6228 17150 6378 17214
rect 6652 17150 6802 17214
rect 4980 16767 5130 16831
rect 5452 16767 5602 16831
rect 5884 16767 6034 16831
rect 6228 16756 6378 16820
rect 6652 16756 6802 16820
rect 4980 16349 5130 16413
rect 5452 16349 5602 16413
rect 5884 16349 6034 16413
rect 6228 16360 6378 16424
rect 6652 16360 6802 16424
rect 4980 15977 5130 16041
rect 5452 15977 5602 16041
rect 5884 15977 6034 16041
rect 6228 15966 6378 16030
rect 6652 15966 6802 16030
rect 4980 15559 5130 15623
rect 5452 15559 5602 15623
rect 5884 15559 6034 15623
rect 6228 15570 6378 15634
rect 6652 15570 6802 15634
rect 4980 15187 5130 15251
rect 5452 15187 5602 15251
rect 5884 15187 6034 15251
rect 6228 15176 6378 15240
rect 6652 15176 6802 15240
rect 4980 14769 5130 14833
rect 5452 14769 5602 14833
rect 5884 14769 6034 14833
rect 6228 14780 6378 14844
rect 6652 14780 6802 14844
rect 4980 14397 5130 14461
rect 5452 14397 5602 14461
rect 5884 14397 6034 14461
rect 6228 14386 6378 14450
rect 6652 14386 6802 14450
rect 4980 13979 5130 14043
rect 5452 13979 5602 14043
rect 5884 13979 6034 14043
rect 6228 13990 6378 14054
rect 6652 13990 6802 14054
rect 4980 13607 5130 13671
rect 5452 13607 5602 13671
rect 5884 13607 6034 13671
rect 6228 13596 6378 13660
rect 6652 13596 6802 13660
rect 4980 13189 5130 13253
rect 5452 13189 5602 13253
rect 5884 13189 6034 13253
rect 6228 13200 6378 13264
rect 6652 13200 6802 13264
rect 4980 12817 5130 12881
rect 5452 12817 5602 12881
rect 5884 12817 6034 12881
rect 6228 12806 6378 12870
rect 6652 12806 6802 12870
rect 4980 12399 5130 12463
rect 5452 12399 5602 12463
rect 5884 12399 6034 12463
rect 6228 12410 6378 12474
rect 6652 12410 6802 12474
rect 4980 12027 5130 12091
rect 5452 12027 5602 12091
rect 5884 12027 6034 12091
rect 6228 12016 6378 12080
rect 6652 12016 6802 12080
rect 4980 11609 5130 11673
rect 5452 11609 5602 11673
rect 5884 11609 6034 11673
rect 6228 11620 6378 11684
rect 6652 11620 6802 11684
rect 4980 11237 5130 11301
rect 5452 11237 5602 11301
rect 5884 11237 6034 11301
rect 6228 11226 6378 11290
rect 6652 11226 6802 11290
rect 4980 10819 5130 10883
rect 5452 10819 5602 10883
rect 5884 10819 6034 10883
rect 6228 10830 6378 10894
rect 6652 10830 6802 10894
rect 4980 10447 5130 10511
rect 5452 10447 5602 10511
rect 5884 10447 6034 10511
rect 6228 10436 6378 10500
rect 6652 10436 6802 10500
rect 4980 10029 5130 10093
rect 5452 10029 5602 10093
rect 5884 10029 6034 10093
rect 6228 10040 6378 10104
rect 6652 10040 6802 10104
rect 4980 9657 5130 9721
rect 5452 9657 5602 9721
rect 5884 9657 6034 9721
rect 6228 9646 6378 9710
rect 6652 9646 6802 9710
rect 4980 9239 5130 9303
rect 5452 9239 5602 9303
rect 5884 9239 6034 9303
rect 6228 9250 6378 9314
rect 6652 9250 6802 9314
rect 4980 8867 5130 8931
rect 5452 8867 5602 8931
rect 5884 8867 6034 8931
rect 6228 8856 6378 8920
rect 6652 8856 6802 8920
rect 4980 8449 5130 8513
rect 5452 8449 5602 8513
rect 5884 8449 6034 8513
rect 6228 8460 6378 8524
rect 6652 8460 6802 8524
rect 4980 8077 5130 8141
rect 5452 8077 5602 8141
rect 5884 8077 6034 8141
rect 6228 8066 6378 8130
rect 6652 8066 6802 8130
rect 4980 7659 5130 7723
rect 5452 7659 5602 7723
rect 5884 7659 6034 7723
rect 6228 7670 6378 7734
rect 6652 7670 6802 7734
rect 4980 7287 5130 7351
rect 5452 7287 5602 7351
rect 5884 7287 6034 7351
rect 6228 7276 6378 7340
rect 6652 7276 6802 7340
rect 4980 6869 5130 6933
rect 5452 6869 5602 6933
rect 5884 6869 6034 6933
rect 6228 6880 6378 6944
rect 6652 6880 6802 6944
rect 4980 6497 5130 6561
rect 5452 6497 5602 6561
rect 5884 6497 6034 6561
rect 6228 6486 6378 6550
rect 6652 6486 6802 6550
rect 4980 6079 5130 6143
rect 5452 6079 5602 6143
rect 5884 6079 6034 6143
rect 6228 6090 6378 6154
rect 6652 6090 6802 6154
rect 2290 5883 2388 5981
rect 2715 5883 2813 5981
rect 3094 5876 3192 5974
rect 3490 5876 3588 5974
rect 4980 5707 5130 5771
rect 5452 5707 5602 5771
rect 5884 5707 6034 5771
rect 6228 5696 6378 5760
rect 6652 5696 6802 5760
rect 4980 5289 5130 5353
rect 5452 5289 5602 5353
rect 5884 5289 6034 5353
rect 6228 5300 6378 5364
rect 6652 5300 6802 5364
rect 996 5086 1094 5184
rect 1392 5086 1490 5184
rect 2290 5093 2388 5191
rect 2715 5093 2813 5191
rect 3094 5086 3192 5184
rect 3490 5086 3588 5184
rect 4980 4917 5130 4981
rect 5452 4917 5602 4981
rect 5884 4917 6034 4981
rect 6228 4906 6378 4970
rect 6652 4906 6802 4970
rect 4980 4499 5130 4563
rect 5452 4499 5602 4563
rect 5884 4499 6034 4563
rect 6228 4510 6378 4574
rect 6652 4510 6802 4574
rect 4980 4127 5130 4191
rect 5452 4127 5602 4191
rect 5884 4127 6034 4191
rect 6228 4116 6378 4180
rect 6652 4116 6802 4180
rect 4980 3709 5130 3773
rect 5452 3709 5602 3773
rect 5884 3709 6034 3773
rect 6228 3720 6378 3784
rect 6652 3720 6802 3784
rect 2290 3513 2388 3611
rect 2715 3513 2813 3611
rect 3094 3506 3192 3604
rect 3490 3506 3588 3604
rect 4980 3337 5130 3401
rect 5452 3337 5602 3401
rect 5884 3337 6034 3401
rect 6228 3326 6378 3390
rect 6652 3326 6802 3390
rect 4980 2919 5130 2983
rect 5452 2919 5602 2983
rect 5884 2919 6034 2983
rect 6228 2930 6378 2994
rect 6652 2930 6802 2994
rect 996 2716 1094 2814
rect 1392 2716 1490 2814
rect 2290 2723 2388 2821
rect 2715 2723 2813 2821
rect 3094 2716 3192 2814
rect 3490 2716 3588 2814
rect 4980 2547 5130 2611
rect 5452 2547 5602 2611
rect 5884 2547 6034 2611
rect 6228 2536 6378 2600
rect 6652 2536 6802 2600
rect 4980 2129 5130 2193
rect 5452 2129 5602 2193
rect 5884 2129 6034 2193
rect 6228 2140 6378 2204
rect 6652 2140 6802 2204
rect 4980 1757 5130 1821
rect 5452 1757 5602 1821
rect 5884 1757 6034 1821
rect 6228 1746 6378 1810
rect 6652 1746 6802 1810
rect 4980 1339 5130 1403
rect 5452 1339 5602 1403
rect 5884 1339 6034 1403
rect 6228 1350 6378 1414
rect 6652 1350 6802 1414
rect 2290 1143 2388 1241
rect 2715 1143 2813 1241
rect 3094 1136 3192 1234
rect 3490 1136 3588 1234
rect 4980 967 5130 1031
rect 5452 967 5602 1031
rect 5884 967 6034 1031
rect 6228 956 6378 1020
rect 6652 956 6802 1020
rect 4980 549 5130 613
rect 5452 549 5602 613
rect 5884 549 6034 613
rect 6228 560 6378 624
rect 6652 560 6802 624
rect 996 346 1094 444
rect 1392 346 1490 444
rect 2290 353 2388 451
rect 2715 353 2813 451
rect 3094 346 3192 444
rect 3490 346 3588 444
rect 4980 177 5130 241
rect 5452 177 5602 241
rect 5884 177 6034 241
rect 6228 166 6378 230
rect 6652 166 6802 230
<< metal4 >>
rect 5022 -33 5088 25341
rect 5494 -33 5560 25341
rect 5926 -33 5992 25341
rect 6270 -33 6336 25341
rect 6694 -33 6760 25341
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_0
timestamp 1661296025
transform 1 0 4807 0 -1 25280
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_1
timestamp 1661296025
transform 1 0 4807 0 1 24490
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_2
timestamp 1661296025
transform 1 0 4807 0 -1 24490
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_3
timestamp 1661296025
transform 1 0 4807 0 1 23700
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_4
timestamp 1661296025
transform 1 0 4807 0 -1 23700
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_5
timestamp 1661296025
transform 1 0 4807 0 1 22910
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_6
timestamp 1661296025
transform 1 0 4807 0 -1 22910
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_7
timestamp 1661296025
transform 1 0 4807 0 1 22120
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_8
timestamp 1661296025
transform 1 0 4807 0 -1 22120
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_9
timestamp 1661296025
transform 1 0 4807 0 1 21330
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_10
timestamp 1661296025
transform 1 0 4807 0 -1 21330
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_11
timestamp 1661296025
transform 1 0 4807 0 1 20540
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_12
timestamp 1661296025
transform 1 0 4807 0 -1 20540
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_13
timestamp 1661296025
transform 1 0 4807 0 1 19750
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_14
timestamp 1661296025
transform 1 0 4807 0 -1 19750
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_15
timestamp 1661296025
transform 1 0 4807 0 1 18960
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_16
timestamp 1661296025
transform 1 0 4807 0 -1 18960
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_17
timestamp 1661296025
transform 1 0 4807 0 1 18170
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_18
timestamp 1661296025
transform 1 0 4807 0 -1 18170
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_19
timestamp 1661296025
transform 1 0 4807 0 1 17380
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_20
timestamp 1661296025
transform 1 0 4807 0 -1 17380
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_21
timestamp 1661296025
transform 1 0 4807 0 1 16590
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_22
timestamp 1661296025
transform 1 0 4807 0 -1 16590
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_23
timestamp 1661296025
transform 1 0 4807 0 1 15800
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_24
timestamp 1661296025
transform 1 0 4807 0 -1 15800
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_25
timestamp 1661296025
transform 1 0 4807 0 1 15010
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_26
timestamp 1661296025
transform 1 0 4807 0 -1 15010
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_27
timestamp 1661296025
transform 1 0 4807 0 1 14220
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_28
timestamp 1661296025
transform 1 0 4807 0 -1 14220
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_29
timestamp 1661296025
transform 1 0 4807 0 1 13430
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_30
timestamp 1661296025
transform 1 0 4807 0 -1 13430
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_31
timestamp 1661296025
transform 1 0 4807 0 1 12640
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_32
timestamp 1661296025
transform 1 0 4807 0 -1 12640
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_33
timestamp 1661296025
transform 1 0 4807 0 1 11850
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_34
timestamp 1661296025
transform 1 0 4807 0 -1 11850
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_35
timestamp 1661296025
transform 1 0 4807 0 1 11060
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_36
timestamp 1661296025
transform 1 0 4807 0 -1 11060
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_37
timestamp 1661296025
transform 1 0 4807 0 1 10270
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_38
timestamp 1661296025
transform 1 0 4807 0 -1 10270
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_39
timestamp 1661296025
transform 1 0 4807 0 1 9480
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_40
timestamp 1661296025
transform 1 0 4807 0 -1 9480
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_41
timestamp 1661296025
transform 1 0 4807 0 1 8690
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_42
timestamp 1661296025
transform 1 0 4807 0 -1 8690
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_43
timestamp 1661296025
transform 1 0 4807 0 1 7900
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_44
timestamp 1661296025
transform 1 0 4807 0 -1 7900
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_45
timestamp 1661296025
transform 1 0 4807 0 1 7110
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_46
timestamp 1661296025
transform 1 0 4807 0 -1 7110
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_47
timestamp 1661296025
transform 1 0 4807 0 1 6320
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_48
timestamp 1661296025
transform 1 0 4807 0 -1 6320
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_49
timestamp 1661296025
transform 1 0 4807 0 1 5530
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_50
timestamp 1661296025
transform 1 0 4807 0 -1 5530
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_51
timestamp 1661296025
transform 1 0 4807 0 1 4740
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_52
timestamp 1661296025
transform 1 0 4807 0 -1 4740
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_53
timestamp 1661296025
transform 1 0 4807 0 1 3950
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_54
timestamp 1661296025
transform 1 0 4807 0 -1 3950
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_55
timestamp 1661296025
transform 1 0 4807 0 1 3160
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_56
timestamp 1661296025
transform 1 0 4807 0 -1 3160
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_57
timestamp 1661296025
transform 1 0 4807 0 1 2370
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_58
timestamp 1661296025
transform 1 0 4807 0 -1 2370
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_59
timestamp 1661296025
transform 1 0 4807 0 1 1580
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_60
timestamp 1661296025
transform 1 0 4807 0 -1 1580
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_61
timestamp 1661296025
transform 1 0 4807 0 1 790
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_62
timestamp 1661296025
transform 1 0 4807 0 -1 790
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_and3_dec  sky130_sram_1r1w_24x128_8_and3_dec_63
timestamp 1661296025
transform 1 0 4807 0 1 0
box 0 -60 2072 490
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_0
timestamp 1661296025
transform 1 0 3658 0 1 6167
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_1
timestamp 1661296025
transform 1 0 3658 0 1 5617
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_2
timestamp 1661296025
transform 1 0 3658 0 1 5377
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_3
timestamp 1661296025
transform 1 0 3658 0 1 4827
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_4
timestamp 1661296025
transform 1 0 3658 0 1 3797
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_5
timestamp 1661296025
transform 1 0 3658 0 1 3247
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_6
timestamp 1661296025
transform 1 0 3658 0 1 3007
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_7
timestamp 1661296025
transform 1 0 3658 0 1 2457
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_8
timestamp 1661296025
transform 1 0 3658 0 1 1427
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_9
timestamp 1661296025
transform 1 0 3658 0 1 877
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_10
timestamp 1661296025
transform 1 0 3658 0 1 637
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_11
timestamp 1661296025
transform 1 0 3658 0 1 87
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_12
timestamp 1661296025
transform 1 0 672 0 1 5327
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_13
timestamp 1661296025
transform 1 0 592 0 1 4877
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_14
timestamp 1661296025
transform 1 0 672 0 1 2957
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_15
timestamp 1661296025
transform 1 0 592 0 1 2507
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_16
timestamp 1661296025
transform 1 0 672 0 1 587
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_17
timestamp 1661296025
transform 1 0 592 0 1 137
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_0
timestamp 1661296025
transform 1 0 4628 0 1 24968
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_1
timestamp 1661296025
transform 1 0 4308 0 1 25058
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_2
timestamp 1661296025
transform 1 0 3988 0 1 25170
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_3
timestamp 1661296025
transform 1 0 4628 0 1 24744
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_4
timestamp 1661296025
transform 1 0 4308 0 1 24654
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_5
timestamp 1661296025
transform 1 0 3908 0 1 24542
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_6
timestamp 1661296025
transform 1 0 4628 0 1 24178
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_7
timestamp 1661296025
transform 1 0 4308 0 1 24268
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_8
timestamp 1661296025
transform 1 0 3828 0 1 24380
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_9
timestamp 1661296025
transform 1 0 4628 0 1 23954
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_10
timestamp 1661296025
transform 1 0 4308 0 1 23864
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_11
timestamp 1661296025
transform 1 0 3748 0 1 23752
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_12
timestamp 1661296025
transform 1 0 4628 0 1 23388
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_13
timestamp 1661296025
transform 1 0 4228 0 1 23478
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_14
timestamp 1661296025
transform 1 0 3988 0 1 23590
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_15
timestamp 1661296025
transform 1 0 4628 0 1 23164
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_16
timestamp 1661296025
transform 1 0 4228 0 1 23074
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_17
timestamp 1661296025
transform 1 0 3908 0 1 22962
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_18
timestamp 1661296025
transform 1 0 4628 0 1 22598
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_19
timestamp 1661296025
transform 1 0 4228 0 1 22688
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_20
timestamp 1661296025
transform 1 0 3828 0 1 22800
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_21
timestamp 1661296025
transform 1 0 4628 0 1 22374
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_22
timestamp 1661296025
transform 1 0 4228 0 1 22284
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_23
timestamp 1661296025
transform 1 0 3748 0 1 22172
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_24
timestamp 1661296025
transform 1 0 4628 0 1 21808
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_25
timestamp 1661296025
transform 1 0 4148 0 1 21898
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_26
timestamp 1661296025
transform 1 0 3988 0 1 22010
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_27
timestamp 1661296025
transform 1 0 4628 0 1 21584
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_28
timestamp 1661296025
transform 1 0 4148 0 1 21494
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_29
timestamp 1661296025
transform 1 0 3908 0 1 21382
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_30
timestamp 1661296025
transform 1 0 4628 0 1 21018
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_31
timestamp 1661296025
transform 1 0 4148 0 1 21108
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_32
timestamp 1661296025
transform 1 0 3828 0 1 21220
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_33
timestamp 1661296025
transform 1 0 4628 0 1 20794
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_34
timestamp 1661296025
transform 1 0 4148 0 1 20704
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_35
timestamp 1661296025
transform 1 0 3748 0 1 20592
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_36
timestamp 1661296025
transform 1 0 4628 0 1 20228
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_37
timestamp 1661296025
transform 1 0 4068 0 1 20318
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_38
timestamp 1661296025
transform 1 0 3988 0 1 20430
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_39
timestamp 1661296025
transform 1 0 4628 0 1 20004
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_40
timestamp 1661296025
transform 1 0 4068 0 1 19914
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_41
timestamp 1661296025
transform 1 0 3908 0 1 19802
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_42
timestamp 1661296025
transform 1 0 4628 0 1 19438
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_43
timestamp 1661296025
transform 1 0 4068 0 1 19528
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_44
timestamp 1661296025
transform 1 0 3828 0 1 19640
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_45
timestamp 1661296025
transform 1 0 4628 0 1 19214
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_46
timestamp 1661296025
transform 1 0 4068 0 1 19124
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_47
timestamp 1661296025
transform 1 0 3748 0 1 19012
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_48
timestamp 1661296025
transform 1 0 4548 0 1 18648
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_49
timestamp 1661296025
transform 1 0 4308 0 1 18738
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_50
timestamp 1661296025
transform 1 0 3988 0 1 18850
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_51
timestamp 1661296025
transform 1 0 4548 0 1 18424
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_52
timestamp 1661296025
transform 1 0 4308 0 1 18334
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_53
timestamp 1661296025
transform 1 0 3908 0 1 18222
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_54
timestamp 1661296025
transform 1 0 4548 0 1 17858
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_55
timestamp 1661296025
transform 1 0 4308 0 1 17948
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_56
timestamp 1661296025
transform 1 0 3828 0 1 18060
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_57
timestamp 1661296025
transform 1 0 4548 0 1 17634
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_58
timestamp 1661296025
transform 1 0 4308 0 1 17544
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_59
timestamp 1661296025
transform 1 0 3748 0 1 17432
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_60
timestamp 1661296025
transform 1 0 4548 0 1 17068
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_61
timestamp 1661296025
transform 1 0 4228 0 1 17158
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_62
timestamp 1661296025
transform 1 0 3988 0 1 17270
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_63
timestamp 1661296025
transform 1 0 4548 0 1 16844
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_64
timestamp 1661296025
transform 1 0 4228 0 1 16754
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_65
timestamp 1661296025
transform 1 0 3908 0 1 16642
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_66
timestamp 1661296025
transform 1 0 4548 0 1 16278
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_67
timestamp 1661296025
transform 1 0 4228 0 1 16368
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_68
timestamp 1661296025
transform 1 0 3828 0 1 16480
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_69
timestamp 1661296025
transform 1 0 4548 0 1 16054
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_70
timestamp 1661296025
transform 1 0 4228 0 1 15964
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_71
timestamp 1661296025
transform 1 0 3748 0 1 15852
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_72
timestamp 1661296025
transform 1 0 4548 0 1 15488
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_73
timestamp 1661296025
transform 1 0 4148 0 1 15578
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_74
timestamp 1661296025
transform 1 0 3988 0 1 15690
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_75
timestamp 1661296025
transform 1 0 4548 0 1 15264
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_76
timestamp 1661296025
transform 1 0 4148 0 1 15174
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_77
timestamp 1661296025
transform 1 0 3908 0 1 15062
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_78
timestamp 1661296025
transform 1 0 4548 0 1 14698
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_79
timestamp 1661296025
transform 1 0 4148 0 1 14788
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_80
timestamp 1661296025
transform 1 0 3828 0 1 14900
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_81
timestamp 1661296025
transform 1 0 4548 0 1 14474
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_82
timestamp 1661296025
transform 1 0 4148 0 1 14384
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_83
timestamp 1661296025
transform 1 0 3748 0 1 14272
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_84
timestamp 1661296025
transform 1 0 4548 0 1 13908
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_85
timestamp 1661296025
transform 1 0 4068 0 1 13998
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_86
timestamp 1661296025
transform 1 0 3988 0 1 14110
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_87
timestamp 1661296025
transform 1 0 4548 0 1 13684
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_88
timestamp 1661296025
transform 1 0 4068 0 1 13594
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_89
timestamp 1661296025
transform 1 0 3908 0 1 13482
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_90
timestamp 1661296025
transform 1 0 4548 0 1 13118
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_91
timestamp 1661296025
transform 1 0 4068 0 1 13208
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_92
timestamp 1661296025
transform 1 0 3828 0 1 13320
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_93
timestamp 1661296025
transform 1 0 4548 0 1 12894
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_94
timestamp 1661296025
transform 1 0 4068 0 1 12804
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_95
timestamp 1661296025
transform 1 0 3748 0 1 12692
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_96
timestamp 1661296025
transform 1 0 4468 0 1 12328
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_97
timestamp 1661296025
transform 1 0 4308 0 1 12418
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_98
timestamp 1661296025
transform 1 0 3988 0 1 12530
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_99
timestamp 1661296025
transform 1 0 4468 0 1 12104
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_100
timestamp 1661296025
transform 1 0 4308 0 1 12014
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_101
timestamp 1661296025
transform 1 0 3908 0 1 11902
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_102
timestamp 1661296025
transform 1 0 4468 0 1 11538
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_103
timestamp 1661296025
transform 1 0 4308 0 1 11628
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_104
timestamp 1661296025
transform 1 0 3828 0 1 11740
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_105
timestamp 1661296025
transform 1 0 4468 0 1 11314
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_106
timestamp 1661296025
transform 1 0 4308 0 1 11224
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_107
timestamp 1661296025
transform 1 0 3748 0 1 11112
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_108
timestamp 1661296025
transform 1 0 4468 0 1 10748
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_109
timestamp 1661296025
transform 1 0 4228 0 1 10838
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_110
timestamp 1661296025
transform 1 0 3988 0 1 10950
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_111
timestamp 1661296025
transform 1 0 4468 0 1 10524
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_112
timestamp 1661296025
transform 1 0 4228 0 1 10434
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_113
timestamp 1661296025
transform 1 0 3908 0 1 10322
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_114
timestamp 1661296025
transform 1 0 4468 0 1 9958
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_115
timestamp 1661296025
transform 1 0 4228 0 1 10048
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_116
timestamp 1661296025
transform 1 0 3828 0 1 10160
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_117
timestamp 1661296025
transform 1 0 4468 0 1 9734
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_118
timestamp 1661296025
transform 1 0 4228 0 1 9644
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_119
timestamp 1661296025
transform 1 0 3748 0 1 9532
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_120
timestamp 1661296025
transform 1 0 4468 0 1 9168
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_121
timestamp 1661296025
transform 1 0 4148 0 1 9258
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_122
timestamp 1661296025
transform 1 0 3988 0 1 9370
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_123
timestamp 1661296025
transform 1 0 4468 0 1 8944
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_124
timestamp 1661296025
transform 1 0 4148 0 1 8854
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_125
timestamp 1661296025
transform 1 0 3908 0 1 8742
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_126
timestamp 1661296025
transform 1 0 4468 0 1 8378
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_127
timestamp 1661296025
transform 1 0 4148 0 1 8468
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_128
timestamp 1661296025
transform 1 0 3828 0 1 8580
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_129
timestamp 1661296025
transform 1 0 4468 0 1 8154
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_130
timestamp 1661296025
transform 1 0 4148 0 1 8064
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_131
timestamp 1661296025
transform 1 0 3748 0 1 7952
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_132
timestamp 1661296025
transform 1 0 4468 0 1 7588
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_133
timestamp 1661296025
transform 1 0 4068 0 1 7678
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_134
timestamp 1661296025
transform 1 0 3988 0 1 7790
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_135
timestamp 1661296025
transform 1 0 4468 0 1 7364
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_136
timestamp 1661296025
transform 1 0 4068 0 1 7274
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_137
timestamp 1661296025
transform 1 0 3908 0 1 7162
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_138
timestamp 1661296025
transform 1 0 4468 0 1 6798
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_139
timestamp 1661296025
transform 1 0 4068 0 1 6888
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_140
timestamp 1661296025
transform 1 0 3828 0 1 7000
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_141
timestamp 1661296025
transform 1 0 4468 0 1 6574
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_142
timestamp 1661296025
transform 1 0 4068 0 1 6484
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_143
timestamp 1661296025
transform 1 0 3748 0 1 6372
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_144
timestamp 1661296025
transform 1 0 4388 0 1 6008
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_145
timestamp 1661296025
transform 1 0 4308 0 1 6098
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_146
timestamp 1661296025
transform 1 0 3988 0 1 6210
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_147
timestamp 1661296025
transform 1 0 4388 0 1 5784
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_148
timestamp 1661296025
transform 1 0 4308 0 1 5694
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_149
timestamp 1661296025
transform 1 0 3908 0 1 5582
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_150
timestamp 1661296025
transform 1 0 4388 0 1 5218
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_151
timestamp 1661296025
transform 1 0 4308 0 1 5308
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_152
timestamp 1661296025
transform 1 0 3828 0 1 5420
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_153
timestamp 1661296025
transform 1 0 4388 0 1 4994
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_154
timestamp 1661296025
transform 1 0 4308 0 1 4904
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_155
timestamp 1661296025
transform 1 0 3748 0 1 4792
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_156
timestamp 1661296025
transform 1 0 4388 0 1 4428
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_157
timestamp 1661296025
transform 1 0 4228 0 1 4518
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_158
timestamp 1661296025
transform 1 0 3988 0 1 4630
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_159
timestamp 1661296025
transform 1 0 4388 0 1 4204
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_160
timestamp 1661296025
transform 1 0 4228 0 1 4114
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_161
timestamp 1661296025
transform 1 0 3908 0 1 4002
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_162
timestamp 1661296025
transform 1 0 4388 0 1 3638
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_163
timestamp 1661296025
transform 1 0 4228 0 1 3728
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_164
timestamp 1661296025
transform 1 0 3828 0 1 3840
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_165
timestamp 1661296025
transform 1 0 4388 0 1 3414
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_166
timestamp 1661296025
transform 1 0 4228 0 1 3324
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_167
timestamp 1661296025
transform 1 0 3748 0 1 3212
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_168
timestamp 1661296025
transform 1 0 4388 0 1 2848
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_169
timestamp 1661296025
transform 1 0 4148 0 1 2938
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_170
timestamp 1661296025
transform 1 0 3988 0 1 3050
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_171
timestamp 1661296025
transform 1 0 4388 0 1 2624
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_172
timestamp 1661296025
transform 1 0 4148 0 1 2534
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_173
timestamp 1661296025
transform 1 0 3908 0 1 2422
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_174
timestamp 1661296025
transform 1 0 4388 0 1 2058
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_175
timestamp 1661296025
transform 1 0 4148 0 1 2148
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_176
timestamp 1661296025
transform 1 0 3828 0 1 2260
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_177
timestamp 1661296025
transform 1 0 4388 0 1 1834
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_178
timestamp 1661296025
transform 1 0 4148 0 1 1744
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_179
timestamp 1661296025
transform 1 0 3748 0 1 1632
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_180
timestamp 1661296025
transform 1 0 4388 0 1 1268
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_181
timestamp 1661296025
transform 1 0 4068 0 1 1358
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_182
timestamp 1661296025
transform 1 0 3988 0 1 1470
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_183
timestamp 1661296025
transform 1 0 4388 0 1 1044
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_184
timestamp 1661296025
transform 1 0 4068 0 1 954
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_185
timestamp 1661296025
transform 1 0 3908 0 1 842
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_186
timestamp 1661296025
transform 1 0 4388 0 1 478
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_187
timestamp 1661296025
transform 1 0 4068 0 1 568
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_188
timestamp 1661296025
transform 1 0 3828 0 1 680
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_189
timestamp 1661296025
transform 1 0 4388 0 1 254
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_190
timestamp 1661296025
transform 1 0 4068 0 1 164
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_191
timestamp 1661296025
transform 1 0 3748 0 1 52
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_192
timestamp 1661296025
transform 1 0 400 0 1 5331
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_193
timestamp 1661296025
transform 1 0 320 0 1 4881
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_194
timestamp 1661296025
transform 1 0 240 0 1 2961
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_195
timestamp 1661296025
transform 1 0 160 0 1 2511
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_196
timestamp 1661296025
transform 1 0 80 0 1 591
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_197
timestamp 1661296025
transform 1 0 0 0 1 141
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_0
timestamp 1661296025
transform 1 0 5023 0 1 25039
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_1
timestamp 1661296025
transform 1 0 5023 0 1 24667
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_2
timestamp 1661296025
transform 1 0 5023 0 1 24249
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_3
timestamp 1661296025
transform 1 0 5023 0 1 23877
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_4
timestamp 1661296025
transform 1 0 5023 0 1 23459
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_5
timestamp 1661296025
transform 1 0 5023 0 1 23087
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_6
timestamp 1661296025
transform 1 0 5023 0 1 22669
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_7
timestamp 1661296025
transform 1 0 5023 0 1 22297
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_8
timestamp 1661296025
transform 1 0 5023 0 1 21879
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_9
timestamp 1661296025
transform 1 0 5023 0 1 21507
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_10
timestamp 1661296025
transform 1 0 5023 0 1 21089
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_11
timestamp 1661296025
transform 1 0 5023 0 1 20717
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_12
timestamp 1661296025
transform 1 0 5023 0 1 20299
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_13
timestamp 1661296025
transform 1 0 5023 0 1 19927
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_14
timestamp 1661296025
transform 1 0 5023 0 1 19509
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_15
timestamp 1661296025
transform 1 0 5023 0 1 19137
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_16
timestamp 1661296025
transform 1 0 5023 0 1 18719
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_17
timestamp 1661296025
transform 1 0 5023 0 1 18347
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_18
timestamp 1661296025
transform 1 0 5023 0 1 17929
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_19
timestamp 1661296025
transform 1 0 5023 0 1 17557
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_20
timestamp 1661296025
transform 1 0 5023 0 1 17139
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_21
timestamp 1661296025
transform 1 0 5023 0 1 16767
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_22
timestamp 1661296025
transform 1 0 5023 0 1 16349
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_23
timestamp 1661296025
transform 1 0 5023 0 1 15977
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_24
timestamp 1661296025
transform 1 0 5023 0 1 15559
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_25
timestamp 1661296025
transform 1 0 5023 0 1 15187
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_26
timestamp 1661296025
transform 1 0 5023 0 1 14769
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_27
timestamp 1661296025
transform 1 0 5023 0 1 14397
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_28
timestamp 1661296025
transform 1 0 5023 0 1 13979
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_29
timestamp 1661296025
transform 1 0 5023 0 1 13607
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_30
timestamp 1661296025
transform 1 0 5023 0 1 13189
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_31
timestamp 1661296025
transform 1 0 5023 0 1 12817
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_32
timestamp 1661296025
transform 1 0 5023 0 1 12399
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_33
timestamp 1661296025
transform 1 0 5023 0 1 12027
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_34
timestamp 1661296025
transform 1 0 5023 0 1 11609
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_35
timestamp 1661296025
transform 1 0 5023 0 1 11237
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_36
timestamp 1661296025
transform 1 0 5023 0 1 10819
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_37
timestamp 1661296025
transform 1 0 5023 0 1 10447
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_38
timestamp 1661296025
transform 1 0 5023 0 1 10029
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_39
timestamp 1661296025
transform 1 0 5023 0 1 9657
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_40
timestamp 1661296025
transform 1 0 5023 0 1 9239
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_41
timestamp 1661296025
transform 1 0 5023 0 1 8867
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_42
timestamp 1661296025
transform 1 0 5023 0 1 8449
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_43
timestamp 1661296025
transform 1 0 5023 0 1 8077
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_44
timestamp 1661296025
transform 1 0 5023 0 1 7659
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_45
timestamp 1661296025
transform 1 0 5023 0 1 7287
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_46
timestamp 1661296025
transform 1 0 5023 0 1 6869
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_47
timestamp 1661296025
transform 1 0 5023 0 1 6497
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_48
timestamp 1661296025
transform 1 0 5023 0 1 6079
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_49
timestamp 1661296025
transform 1 0 5023 0 1 5707
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_50
timestamp 1661296025
transform 1 0 5023 0 1 5289
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_51
timestamp 1661296025
transform 1 0 5023 0 1 4917
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_52
timestamp 1661296025
transform 1 0 5023 0 1 4499
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_53
timestamp 1661296025
transform 1 0 5023 0 1 4127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_54
timestamp 1661296025
transform 1 0 5023 0 1 3709
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_55
timestamp 1661296025
transform 1 0 5023 0 1 3337
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_56
timestamp 1661296025
transform 1 0 5023 0 1 2919
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_57
timestamp 1661296025
transform 1 0 5023 0 1 2547
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_58
timestamp 1661296025
transform 1 0 5023 0 1 2129
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_59
timestamp 1661296025
transform 1 0 5023 0 1 1757
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_60
timestamp 1661296025
transform 1 0 5023 0 1 1339
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_61
timestamp 1661296025
transform 1 0 5023 0 1 967
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_62
timestamp 1661296025
transform 1 0 5023 0 1 549
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_63
timestamp 1661296025
transform 1 0 5023 0 1 177
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_64
timestamp 1661296025
transform 1 0 6271 0 1 25050
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_65
timestamp 1661296025
transform 1 0 6271 0 1 24656
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_66
timestamp 1661296025
transform 1 0 6271 0 1 24260
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_67
timestamp 1661296025
transform 1 0 6271 0 1 23866
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_68
timestamp 1661296025
transform 1 0 6271 0 1 23470
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_69
timestamp 1661296025
transform 1 0 6271 0 1 23076
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_70
timestamp 1661296025
transform 1 0 6271 0 1 22680
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_71
timestamp 1661296025
transform 1 0 6271 0 1 22286
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_72
timestamp 1661296025
transform 1 0 6271 0 1 21890
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_73
timestamp 1661296025
transform 1 0 6271 0 1 21496
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_74
timestamp 1661296025
transform 1 0 6271 0 1 21100
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_75
timestamp 1661296025
transform 1 0 6271 0 1 20706
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_76
timestamp 1661296025
transform 1 0 6271 0 1 20310
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_77
timestamp 1661296025
transform 1 0 6271 0 1 19916
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_78
timestamp 1661296025
transform 1 0 6271 0 1 19520
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_79
timestamp 1661296025
transform 1 0 6271 0 1 19126
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_80
timestamp 1661296025
transform 1 0 6271 0 1 18730
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_81
timestamp 1661296025
transform 1 0 6271 0 1 18336
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_82
timestamp 1661296025
transform 1 0 6271 0 1 17940
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_83
timestamp 1661296025
transform 1 0 6271 0 1 17546
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_84
timestamp 1661296025
transform 1 0 6271 0 1 17150
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_85
timestamp 1661296025
transform 1 0 6271 0 1 16756
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_86
timestamp 1661296025
transform 1 0 6271 0 1 16360
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_87
timestamp 1661296025
transform 1 0 6271 0 1 15966
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_88
timestamp 1661296025
transform 1 0 6271 0 1 15570
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_89
timestamp 1661296025
transform 1 0 6271 0 1 15176
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_90
timestamp 1661296025
transform 1 0 6271 0 1 14780
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_91
timestamp 1661296025
transform 1 0 6271 0 1 14386
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_92
timestamp 1661296025
transform 1 0 6271 0 1 13990
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_93
timestamp 1661296025
transform 1 0 6271 0 1 13596
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_94
timestamp 1661296025
transform 1 0 6271 0 1 13200
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_95
timestamp 1661296025
transform 1 0 6271 0 1 12806
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_96
timestamp 1661296025
transform 1 0 6271 0 1 12410
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_97
timestamp 1661296025
transform 1 0 6271 0 1 12016
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_98
timestamp 1661296025
transform 1 0 6271 0 1 11620
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_99
timestamp 1661296025
transform 1 0 6271 0 1 11226
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_100
timestamp 1661296025
transform 1 0 6271 0 1 10830
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_101
timestamp 1661296025
transform 1 0 6271 0 1 10436
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_102
timestamp 1661296025
transform 1 0 6271 0 1 10040
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_103
timestamp 1661296025
transform 1 0 6271 0 1 9646
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_104
timestamp 1661296025
transform 1 0 6271 0 1 9250
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_105
timestamp 1661296025
transform 1 0 6271 0 1 8856
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_106
timestamp 1661296025
transform 1 0 6271 0 1 8460
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_107
timestamp 1661296025
transform 1 0 6271 0 1 8066
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_108
timestamp 1661296025
transform 1 0 6271 0 1 7670
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_109
timestamp 1661296025
transform 1 0 6271 0 1 7276
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_110
timestamp 1661296025
transform 1 0 6271 0 1 6880
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_111
timestamp 1661296025
transform 1 0 6271 0 1 6486
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_112
timestamp 1661296025
transform 1 0 6271 0 1 6090
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_113
timestamp 1661296025
transform 1 0 6271 0 1 5696
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_114
timestamp 1661296025
transform 1 0 6271 0 1 5300
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_115
timestamp 1661296025
transform 1 0 6271 0 1 4906
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_116
timestamp 1661296025
transform 1 0 6271 0 1 4510
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_117
timestamp 1661296025
transform 1 0 6271 0 1 4116
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_118
timestamp 1661296025
transform 1 0 6271 0 1 3720
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_119
timestamp 1661296025
transform 1 0 6271 0 1 3326
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_120
timestamp 1661296025
transform 1 0 6271 0 1 2930
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_121
timestamp 1661296025
transform 1 0 6271 0 1 2536
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_122
timestamp 1661296025
transform 1 0 6271 0 1 2140
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_123
timestamp 1661296025
transform 1 0 6271 0 1 1746
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_124
timestamp 1661296025
transform 1 0 6271 0 1 1350
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_125
timestamp 1661296025
transform 1 0 6271 0 1 956
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_126
timestamp 1661296025
transform 1 0 6271 0 1 560
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_127
timestamp 1661296025
transform 1 0 6271 0 1 166
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_128
timestamp 1661296025
transform 1 0 5927 0 1 25039
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_129
timestamp 1661296025
transform 1 0 5927 0 1 24667
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_130
timestamp 1661296025
transform 1 0 5927 0 1 24249
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_131
timestamp 1661296025
transform 1 0 5927 0 1 23877
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_132
timestamp 1661296025
transform 1 0 5927 0 1 23459
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_133
timestamp 1661296025
transform 1 0 5927 0 1 23087
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_134
timestamp 1661296025
transform 1 0 5927 0 1 22669
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_135
timestamp 1661296025
transform 1 0 5927 0 1 22297
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_136
timestamp 1661296025
transform 1 0 5927 0 1 21879
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_137
timestamp 1661296025
transform 1 0 5927 0 1 21507
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_138
timestamp 1661296025
transform 1 0 5927 0 1 21089
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_139
timestamp 1661296025
transform 1 0 5927 0 1 20717
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_140
timestamp 1661296025
transform 1 0 5927 0 1 20299
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_141
timestamp 1661296025
transform 1 0 5927 0 1 19927
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_142
timestamp 1661296025
transform 1 0 5927 0 1 19509
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_143
timestamp 1661296025
transform 1 0 5927 0 1 19137
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_144
timestamp 1661296025
transform 1 0 5927 0 1 18719
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_145
timestamp 1661296025
transform 1 0 5927 0 1 18347
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_146
timestamp 1661296025
transform 1 0 5927 0 1 17929
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_147
timestamp 1661296025
transform 1 0 5927 0 1 17557
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_148
timestamp 1661296025
transform 1 0 5927 0 1 17139
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_149
timestamp 1661296025
transform 1 0 5927 0 1 16767
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_150
timestamp 1661296025
transform 1 0 5927 0 1 16349
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_151
timestamp 1661296025
transform 1 0 5927 0 1 15977
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_152
timestamp 1661296025
transform 1 0 5927 0 1 15559
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_153
timestamp 1661296025
transform 1 0 5927 0 1 15187
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_154
timestamp 1661296025
transform 1 0 5927 0 1 14769
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_155
timestamp 1661296025
transform 1 0 5927 0 1 14397
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_156
timestamp 1661296025
transform 1 0 5927 0 1 13979
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_157
timestamp 1661296025
transform 1 0 5927 0 1 13607
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_158
timestamp 1661296025
transform 1 0 5927 0 1 13189
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_159
timestamp 1661296025
transform 1 0 5927 0 1 12817
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_160
timestamp 1661296025
transform 1 0 5927 0 1 12399
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_161
timestamp 1661296025
transform 1 0 5927 0 1 12027
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_162
timestamp 1661296025
transform 1 0 5927 0 1 11609
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_163
timestamp 1661296025
transform 1 0 5927 0 1 11237
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_164
timestamp 1661296025
transform 1 0 5927 0 1 10819
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_165
timestamp 1661296025
transform 1 0 5927 0 1 10447
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_166
timestamp 1661296025
transform 1 0 5927 0 1 10029
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_167
timestamp 1661296025
transform 1 0 5927 0 1 9657
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_168
timestamp 1661296025
transform 1 0 5927 0 1 9239
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_169
timestamp 1661296025
transform 1 0 5927 0 1 8867
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_170
timestamp 1661296025
transform 1 0 5927 0 1 8449
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_171
timestamp 1661296025
transform 1 0 5927 0 1 8077
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_172
timestamp 1661296025
transform 1 0 5927 0 1 7659
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_173
timestamp 1661296025
transform 1 0 5927 0 1 7287
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_174
timestamp 1661296025
transform 1 0 5927 0 1 6869
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_175
timestamp 1661296025
transform 1 0 5927 0 1 6497
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_176
timestamp 1661296025
transform 1 0 5927 0 1 6079
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_177
timestamp 1661296025
transform 1 0 5927 0 1 5707
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_178
timestamp 1661296025
transform 1 0 5927 0 1 5289
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_179
timestamp 1661296025
transform 1 0 5927 0 1 4917
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_180
timestamp 1661296025
transform 1 0 5927 0 1 4499
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_181
timestamp 1661296025
transform 1 0 5927 0 1 4127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_182
timestamp 1661296025
transform 1 0 5927 0 1 3709
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_183
timestamp 1661296025
transform 1 0 5927 0 1 3337
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_184
timestamp 1661296025
transform 1 0 5927 0 1 2919
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_185
timestamp 1661296025
transform 1 0 5927 0 1 2547
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_186
timestamp 1661296025
transform 1 0 5927 0 1 2129
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_187
timestamp 1661296025
transform 1 0 5927 0 1 1757
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_188
timestamp 1661296025
transform 1 0 5927 0 1 1339
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_189
timestamp 1661296025
transform 1 0 5927 0 1 967
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_190
timestamp 1661296025
transform 1 0 5927 0 1 549
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_191
timestamp 1661296025
transform 1 0 5927 0 1 177
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_192
timestamp 1661296025
transform 1 0 6695 0 1 25050
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_193
timestamp 1661296025
transform 1 0 6695 0 1 24656
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_194
timestamp 1661296025
transform 1 0 6695 0 1 24260
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_195
timestamp 1661296025
transform 1 0 6695 0 1 23866
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_196
timestamp 1661296025
transform 1 0 6695 0 1 23470
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_197
timestamp 1661296025
transform 1 0 6695 0 1 23076
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_198
timestamp 1661296025
transform 1 0 6695 0 1 22680
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_199
timestamp 1661296025
transform 1 0 6695 0 1 22286
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_200
timestamp 1661296025
transform 1 0 6695 0 1 21890
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_201
timestamp 1661296025
transform 1 0 6695 0 1 21496
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_202
timestamp 1661296025
transform 1 0 6695 0 1 21100
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_203
timestamp 1661296025
transform 1 0 6695 0 1 20706
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_204
timestamp 1661296025
transform 1 0 6695 0 1 20310
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_205
timestamp 1661296025
transform 1 0 6695 0 1 19916
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_206
timestamp 1661296025
transform 1 0 6695 0 1 19520
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_207
timestamp 1661296025
transform 1 0 6695 0 1 19126
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_208
timestamp 1661296025
transform 1 0 6695 0 1 18730
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_209
timestamp 1661296025
transform 1 0 6695 0 1 18336
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_210
timestamp 1661296025
transform 1 0 6695 0 1 17940
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_211
timestamp 1661296025
transform 1 0 6695 0 1 17546
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_212
timestamp 1661296025
transform 1 0 6695 0 1 17150
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_213
timestamp 1661296025
transform 1 0 6695 0 1 16756
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_214
timestamp 1661296025
transform 1 0 6695 0 1 16360
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_215
timestamp 1661296025
transform 1 0 6695 0 1 15966
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_216
timestamp 1661296025
transform 1 0 6695 0 1 15570
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_217
timestamp 1661296025
transform 1 0 6695 0 1 15176
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_218
timestamp 1661296025
transform 1 0 6695 0 1 14780
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_219
timestamp 1661296025
transform 1 0 6695 0 1 14386
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_220
timestamp 1661296025
transform 1 0 6695 0 1 13990
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_221
timestamp 1661296025
transform 1 0 6695 0 1 13596
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_222
timestamp 1661296025
transform 1 0 6695 0 1 13200
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_223
timestamp 1661296025
transform 1 0 6695 0 1 12806
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_224
timestamp 1661296025
transform 1 0 6695 0 1 12410
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_225
timestamp 1661296025
transform 1 0 6695 0 1 12016
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_226
timestamp 1661296025
transform 1 0 6695 0 1 11620
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_227
timestamp 1661296025
transform 1 0 6695 0 1 11226
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_228
timestamp 1661296025
transform 1 0 6695 0 1 10830
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_229
timestamp 1661296025
transform 1 0 6695 0 1 10436
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_230
timestamp 1661296025
transform 1 0 6695 0 1 10040
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_231
timestamp 1661296025
transform 1 0 6695 0 1 9646
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_232
timestamp 1661296025
transform 1 0 6695 0 1 9250
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_233
timestamp 1661296025
transform 1 0 6695 0 1 8856
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_234
timestamp 1661296025
transform 1 0 6695 0 1 8460
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_235
timestamp 1661296025
transform 1 0 6695 0 1 8066
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_236
timestamp 1661296025
transform 1 0 6695 0 1 7670
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_237
timestamp 1661296025
transform 1 0 6695 0 1 7276
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_238
timestamp 1661296025
transform 1 0 6695 0 1 6880
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_239
timestamp 1661296025
transform 1 0 6695 0 1 6486
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_240
timestamp 1661296025
transform 1 0 6695 0 1 6090
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_241
timestamp 1661296025
transform 1 0 6695 0 1 5696
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_242
timestamp 1661296025
transform 1 0 6695 0 1 5300
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_243
timestamp 1661296025
transform 1 0 6695 0 1 4906
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_244
timestamp 1661296025
transform 1 0 6695 0 1 4510
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_245
timestamp 1661296025
transform 1 0 6695 0 1 4116
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_246
timestamp 1661296025
transform 1 0 6695 0 1 3720
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_247
timestamp 1661296025
transform 1 0 6695 0 1 3326
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_248
timestamp 1661296025
transform 1 0 6695 0 1 2930
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_249
timestamp 1661296025
transform 1 0 6695 0 1 2536
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_250
timestamp 1661296025
transform 1 0 6695 0 1 2140
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_251
timestamp 1661296025
transform 1 0 6695 0 1 1746
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_252
timestamp 1661296025
transform 1 0 6695 0 1 1350
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_253
timestamp 1661296025
transform 1 0 6695 0 1 956
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_254
timestamp 1661296025
transform 1 0 6695 0 1 560
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_255
timestamp 1661296025
transform 1 0 6695 0 1 166
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_256
timestamp 1661296025
transform 1 0 5495 0 1 25039
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_257
timestamp 1661296025
transform 1 0 5495 0 1 24667
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_258
timestamp 1661296025
transform 1 0 5495 0 1 24249
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_259
timestamp 1661296025
transform 1 0 5495 0 1 23877
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_260
timestamp 1661296025
transform 1 0 5495 0 1 23459
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_261
timestamp 1661296025
transform 1 0 5495 0 1 23087
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_262
timestamp 1661296025
transform 1 0 5495 0 1 22669
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_263
timestamp 1661296025
transform 1 0 5495 0 1 22297
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_264
timestamp 1661296025
transform 1 0 5495 0 1 21879
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_265
timestamp 1661296025
transform 1 0 5495 0 1 21507
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_266
timestamp 1661296025
transform 1 0 5495 0 1 21089
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_267
timestamp 1661296025
transform 1 0 5495 0 1 20717
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_268
timestamp 1661296025
transform 1 0 5495 0 1 20299
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_269
timestamp 1661296025
transform 1 0 5495 0 1 19927
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_270
timestamp 1661296025
transform 1 0 5495 0 1 19509
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_271
timestamp 1661296025
transform 1 0 5495 0 1 19137
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_272
timestamp 1661296025
transform 1 0 5495 0 1 18719
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_273
timestamp 1661296025
transform 1 0 5495 0 1 18347
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_274
timestamp 1661296025
transform 1 0 5495 0 1 17929
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_275
timestamp 1661296025
transform 1 0 5495 0 1 17557
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_276
timestamp 1661296025
transform 1 0 5495 0 1 17139
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_277
timestamp 1661296025
transform 1 0 5495 0 1 16767
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_278
timestamp 1661296025
transform 1 0 5495 0 1 16349
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_279
timestamp 1661296025
transform 1 0 5495 0 1 15977
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_280
timestamp 1661296025
transform 1 0 5495 0 1 15559
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_281
timestamp 1661296025
transform 1 0 5495 0 1 15187
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_282
timestamp 1661296025
transform 1 0 5495 0 1 14769
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_283
timestamp 1661296025
transform 1 0 5495 0 1 14397
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_284
timestamp 1661296025
transform 1 0 5495 0 1 13979
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_285
timestamp 1661296025
transform 1 0 5495 0 1 13607
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_286
timestamp 1661296025
transform 1 0 5495 0 1 13189
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_287
timestamp 1661296025
transform 1 0 5495 0 1 12817
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_288
timestamp 1661296025
transform 1 0 5495 0 1 12399
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_289
timestamp 1661296025
transform 1 0 5495 0 1 12027
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_290
timestamp 1661296025
transform 1 0 5495 0 1 11609
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_291
timestamp 1661296025
transform 1 0 5495 0 1 11237
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_292
timestamp 1661296025
transform 1 0 5495 0 1 10819
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_293
timestamp 1661296025
transform 1 0 5495 0 1 10447
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_294
timestamp 1661296025
transform 1 0 5495 0 1 10029
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_295
timestamp 1661296025
transform 1 0 5495 0 1 9657
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_296
timestamp 1661296025
transform 1 0 5495 0 1 9239
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_297
timestamp 1661296025
transform 1 0 5495 0 1 8867
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_298
timestamp 1661296025
transform 1 0 5495 0 1 8449
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_299
timestamp 1661296025
transform 1 0 5495 0 1 8077
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_300
timestamp 1661296025
transform 1 0 5495 0 1 7659
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_301
timestamp 1661296025
transform 1 0 5495 0 1 7287
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_302
timestamp 1661296025
transform 1 0 5495 0 1 6869
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_303
timestamp 1661296025
transform 1 0 5495 0 1 6497
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_304
timestamp 1661296025
transform 1 0 5495 0 1 6079
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_305
timestamp 1661296025
transform 1 0 5495 0 1 5707
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_306
timestamp 1661296025
transform 1 0 5495 0 1 5289
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_307
timestamp 1661296025
transform 1 0 5495 0 1 4917
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_308
timestamp 1661296025
transform 1 0 5495 0 1 4499
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_309
timestamp 1661296025
transform 1 0 5495 0 1 4127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_310
timestamp 1661296025
transform 1 0 5495 0 1 3709
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_311
timestamp 1661296025
transform 1 0 5495 0 1 3337
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_312
timestamp 1661296025
transform 1 0 5495 0 1 2919
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_313
timestamp 1661296025
transform 1 0 5495 0 1 2547
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_314
timestamp 1661296025
transform 1 0 5495 0 1 2129
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_315
timestamp 1661296025
transform 1 0 5495 0 1 1757
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_316
timestamp 1661296025
transform 1 0 5495 0 1 1339
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_317
timestamp 1661296025
transform 1 0 5495 0 1 967
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_318
timestamp 1661296025
transform 1 0 5495 0 1 549
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_319
timestamp 1661296025
transform 1 0 5495 0 1 177
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_320
timestamp 1661296025
transform 1 0 3655 0 1 6168
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_321
timestamp 1661296025
transform 1 0 3655 0 1 5618
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_322
timestamp 1661296025
transform 1 0 3655 0 1 5378
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_323
timestamp 1661296025
transform 1 0 3655 0 1 4828
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_324
timestamp 1661296025
transform 1 0 3655 0 1 3798
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_325
timestamp 1661296025
transform 1 0 3655 0 1 3248
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_326
timestamp 1661296025
transform 1 0 3655 0 1 3008
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_327
timestamp 1661296025
transform 1 0 3655 0 1 2458
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_328
timestamp 1661296025
transform 1 0 3655 0 1 1428
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_329
timestamp 1661296025
transform 1 0 3655 0 1 878
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_330
timestamp 1661296025
transform 1 0 3655 0 1 638
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_331
timestamp 1661296025
transform 1 0 3655 0 1 88
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_0
timestamp 1661296025
transform 1 0 4629 0 1 5893
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_1
timestamp 1661296025
transform 1 0 4549 0 1 5498
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_2
timestamp 1661296025
transform 1 0 4469 0 1 5103
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_3
timestamp 1661296025
transform 1 0 4389 0 1 4708
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_4
timestamp 1661296025
transform 1 0 4309 0 1 3523
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_5
timestamp 1661296025
transform 1 0 4229 0 1 3128
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_6
timestamp 1661296025
transform 1 0 4149 0 1 2733
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_7
timestamp 1661296025
transform 1 0 4069 0 1 2338
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_8
timestamp 1661296025
transform 1 0 3989 0 1 1153
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_9
timestamp 1661296025
transform 1 0 3909 0 1 967
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_10
timestamp 1661296025
transform 1 0 3829 0 1 363
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_11
timestamp 1661296025
transform 1 0 3749 0 1 177
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_0
timestamp 1661296025
transform 1 0 5022 0 1 25034
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_1
timestamp 1661296025
transform 1 0 5022 0 1 24662
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_2
timestamp 1661296025
transform 1 0 5022 0 1 24244
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_3
timestamp 1661296025
transform 1 0 5022 0 1 23872
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_4
timestamp 1661296025
transform 1 0 5022 0 1 23454
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_5
timestamp 1661296025
transform 1 0 5022 0 1 23082
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_6
timestamp 1661296025
transform 1 0 5022 0 1 22664
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_7
timestamp 1661296025
transform 1 0 5022 0 1 22292
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_8
timestamp 1661296025
transform 1 0 5022 0 1 21874
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_9
timestamp 1661296025
transform 1 0 5022 0 1 21502
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_10
timestamp 1661296025
transform 1 0 5022 0 1 21084
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_11
timestamp 1661296025
transform 1 0 5022 0 1 20712
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_12
timestamp 1661296025
transform 1 0 5022 0 1 20294
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_13
timestamp 1661296025
transform 1 0 5022 0 1 19922
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_14
timestamp 1661296025
transform 1 0 5022 0 1 19504
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_15
timestamp 1661296025
transform 1 0 5022 0 1 19132
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_16
timestamp 1661296025
transform 1 0 5022 0 1 18714
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_17
timestamp 1661296025
transform 1 0 5022 0 1 18342
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_18
timestamp 1661296025
transform 1 0 5022 0 1 17924
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_19
timestamp 1661296025
transform 1 0 5022 0 1 17552
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_20
timestamp 1661296025
transform 1 0 5022 0 1 17134
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_21
timestamp 1661296025
transform 1 0 5022 0 1 16762
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_22
timestamp 1661296025
transform 1 0 5022 0 1 16344
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_23
timestamp 1661296025
transform 1 0 5022 0 1 15972
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_24
timestamp 1661296025
transform 1 0 5022 0 1 15554
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_25
timestamp 1661296025
transform 1 0 5022 0 1 15182
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_26
timestamp 1661296025
transform 1 0 5022 0 1 14764
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_27
timestamp 1661296025
transform 1 0 5022 0 1 14392
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_28
timestamp 1661296025
transform 1 0 5022 0 1 13974
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_29
timestamp 1661296025
transform 1 0 5022 0 1 13602
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_30
timestamp 1661296025
transform 1 0 5022 0 1 13184
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_31
timestamp 1661296025
transform 1 0 5022 0 1 12812
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_32
timestamp 1661296025
transform 1 0 5022 0 1 12394
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_33
timestamp 1661296025
transform 1 0 5022 0 1 12022
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_34
timestamp 1661296025
transform 1 0 5022 0 1 11604
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_35
timestamp 1661296025
transform 1 0 5022 0 1 11232
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_36
timestamp 1661296025
transform 1 0 5022 0 1 10814
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_37
timestamp 1661296025
transform 1 0 5022 0 1 10442
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_38
timestamp 1661296025
transform 1 0 5022 0 1 10024
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_39
timestamp 1661296025
transform 1 0 5022 0 1 9652
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_40
timestamp 1661296025
transform 1 0 5022 0 1 9234
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_41
timestamp 1661296025
transform 1 0 5022 0 1 8862
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_42
timestamp 1661296025
transform 1 0 5022 0 1 8444
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_43
timestamp 1661296025
transform 1 0 5022 0 1 8072
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_44
timestamp 1661296025
transform 1 0 5022 0 1 7654
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_45
timestamp 1661296025
transform 1 0 5022 0 1 7282
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_46
timestamp 1661296025
transform 1 0 5022 0 1 6864
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_47
timestamp 1661296025
transform 1 0 5022 0 1 6492
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_48
timestamp 1661296025
transform 1 0 5022 0 1 6074
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_49
timestamp 1661296025
transform 1 0 5022 0 1 5702
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_50
timestamp 1661296025
transform 1 0 5022 0 1 5284
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_51
timestamp 1661296025
transform 1 0 5022 0 1 4912
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_52
timestamp 1661296025
transform 1 0 5022 0 1 4494
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_53
timestamp 1661296025
transform 1 0 5022 0 1 4122
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_54
timestamp 1661296025
transform 1 0 5022 0 1 3704
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_55
timestamp 1661296025
transform 1 0 5022 0 1 3332
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_56
timestamp 1661296025
transform 1 0 5022 0 1 2914
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_57
timestamp 1661296025
transform 1 0 5022 0 1 2542
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_58
timestamp 1661296025
transform 1 0 5022 0 1 2124
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_59
timestamp 1661296025
transform 1 0 5022 0 1 1752
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_60
timestamp 1661296025
transform 1 0 5022 0 1 1334
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_61
timestamp 1661296025
transform 1 0 5022 0 1 962
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_62
timestamp 1661296025
transform 1 0 5022 0 1 544
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_63
timestamp 1661296025
transform 1 0 5022 0 1 172
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_64
timestamp 1661296025
transform 1 0 6270 0 1 25046
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_65
timestamp 1661296025
transform 1 0 6270 0 1 24650
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_66
timestamp 1661296025
transform 1 0 6270 0 1 24256
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_67
timestamp 1661296025
transform 1 0 6270 0 1 23860
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_68
timestamp 1661296025
transform 1 0 6270 0 1 23466
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_69
timestamp 1661296025
transform 1 0 6270 0 1 23070
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_70
timestamp 1661296025
transform 1 0 6270 0 1 22676
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_71
timestamp 1661296025
transform 1 0 6270 0 1 22280
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_72
timestamp 1661296025
transform 1 0 6270 0 1 21886
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_73
timestamp 1661296025
transform 1 0 6270 0 1 21490
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_74
timestamp 1661296025
transform 1 0 6270 0 1 21096
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_75
timestamp 1661296025
transform 1 0 6270 0 1 20700
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_76
timestamp 1661296025
transform 1 0 6270 0 1 20306
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_77
timestamp 1661296025
transform 1 0 6270 0 1 19910
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_78
timestamp 1661296025
transform 1 0 6270 0 1 19516
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_79
timestamp 1661296025
transform 1 0 6270 0 1 19120
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_80
timestamp 1661296025
transform 1 0 6270 0 1 18726
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_81
timestamp 1661296025
transform 1 0 6270 0 1 18330
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_82
timestamp 1661296025
transform 1 0 6270 0 1 17936
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_83
timestamp 1661296025
transform 1 0 6270 0 1 17540
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_84
timestamp 1661296025
transform 1 0 6270 0 1 17146
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_85
timestamp 1661296025
transform 1 0 6270 0 1 16750
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_86
timestamp 1661296025
transform 1 0 6270 0 1 16356
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_87
timestamp 1661296025
transform 1 0 6270 0 1 15960
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_88
timestamp 1661296025
transform 1 0 6270 0 1 15566
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_89
timestamp 1661296025
transform 1 0 6270 0 1 15170
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_90
timestamp 1661296025
transform 1 0 6270 0 1 14776
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_91
timestamp 1661296025
transform 1 0 6270 0 1 14380
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_92
timestamp 1661296025
transform 1 0 6270 0 1 13986
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_93
timestamp 1661296025
transform 1 0 6270 0 1 13590
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_94
timestamp 1661296025
transform 1 0 6270 0 1 13196
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_95
timestamp 1661296025
transform 1 0 6270 0 1 12800
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_96
timestamp 1661296025
transform 1 0 6270 0 1 12406
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_97
timestamp 1661296025
transform 1 0 6270 0 1 12010
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_98
timestamp 1661296025
transform 1 0 6270 0 1 11616
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_99
timestamp 1661296025
transform 1 0 6270 0 1 11220
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_100
timestamp 1661296025
transform 1 0 6270 0 1 10826
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_101
timestamp 1661296025
transform 1 0 6270 0 1 10430
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_102
timestamp 1661296025
transform 1 0 6270 0 1 10036
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_103
timestamp 1661296025
transform 1 0 6270 0 1 9640
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_104
timestamp 1661296025
transform 1 0 6270 0 1 9246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_105
timestamp 1661296025
transform 1 0 6270 0 1 8850
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_106
timestamp 1661296025
transform 1 0 6270 0 1 8456
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_107
timestamp 1661296025
transform 1 0 6270 0 1 8060
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_108
timestamp 1661296025
transform 1 0 6270 0 1 7666
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_109
timestamp 1661296025
transform 1 0 6270 0 1 7270
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_110
timestamp 1661296025
transform 1 0 6270 0 1 6876
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_111
timestamp 1661296025
transform 1 0 6270 0 1 6480
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_112
timestamp 1661296025
transform 1 0 6270 0 1 6086
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_113
timestamp 1661296025
transform 1 0 6270 0 1 5690
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_114
timestamp 1661296025
transform 1 0 6270 0 1 5296
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_115
timestamp 1661296025
transform 1 0 6270 0 1 4900
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_116
timestamp 1661296025
transform 1 0 6270 0 1 4506
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_117
timestamp 1661296025
transform 1 0 6270 0 1 4110
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_118
timestamp 1661296025
transform 1 0 6270 0 1 3716
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_119
timestamp 1661296025
transform 1 0 6270 0 1 3320
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_120
timestamp 1661296025
transform 1 0 6270 0 1 2926
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_121
timestamp 1661296025
transform 1 0 6270 0 1 2530
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_122
timestamp 1661296025
transform 1 0 6270 0 1 2136
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_123
timestamp 1661296025
transform 1 0 6270 0 1 1740
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_124
timestamp 1661296025
transform 1 0 6270 0 1 1346
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_125
timestamp 1661296025
transform 1 0 6270 0 1 950
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_126
timestamp 1661296025
transform 1 0 6270 0 1 556
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_127
timestamp 1661296025
transform 1 0 6270 0 1 160
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_128
timestamp 1661296025
transform 1 0 5926 0 1 25034
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_129
timestamp 1661296025
transform 1 0 5926 0 1 24662
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_130
timestamp 1661296025
transform 1 0 5926 0 1 24244
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_131
timestamp 1661296025
transform 1 0 5926 0 1 23872
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_132
timestamp 1661296025
transform 1 0 5926 0 1 23454
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_133
timestamp 1661296025
transform 1 0 5926 0 1 23082
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_134
timestamp 1661296025
transform 1 0 5926 0 1 22664
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_135
timestamp 1661296025
transform 1 0 5926 0 1 22292
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_136
timestamp 1661296025
transform 1 0 5926 0 1 21874
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_137
timestamp 1661296025
transform 1 0 5926 0 1 21502
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_138
timestamp 1661296025
transform 1 0 5926 0 1 21084
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_139
timestamp 1661296025
transform 1 0 5926 0 1 20712
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_140
timestamp 1661296025
transform 1 0 5926 0 1 20294
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_141
timestamp 1661296025
transform 1 0 5926 0 1 19922
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_142
timestamp 1661296025
transform 1 0 5926 0 1 19504
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_143
timestamp 1661296025
transform 1 0 5926 0 1 19132
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_144
timestamp 1661296025
transform 1 0 5926 0 1 18714
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_145
timestamp 1661296025
transform 1 0 5926 0 1 18342
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_146
timestamp 1661296025
transform 1 0 5926 0 1 17924
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_147
timestamp 1661296025
transform 1 0 5926 0 1 17552
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_148
timestamp 1661296025
transform 1 0 5926 0 1 17134
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_149
timestamp 1661296025
transform 1 0 5926 0 1 16762
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_150
timestamp 1661296025
transform 1 0 5926 0 1 16344
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_151
timestamp 1661296025
transform 1 0 5926 0 1 15972
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_152
timestamp 1661296025
transform 1 0 5926 0 1 15554
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_153
timestamp 1661296025
transform 1 0 5926 0 1 15182
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_154
timestamp 1661296025
transform 1 0 5926 0 1 14764
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_155
timestamp 1661296025
transform 1 0 5926 0 1 14392
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_156
timestamp 1661296025
transform 1 0 5926 0 1 13974
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_157
timestamp 1661296025
transform 1 0 5926 0 1 13602
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_158
timestamp 1661296025
transform 1 0 5926 0 1 13184
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_159
timestamp 1661296025
transform 1 0 5926 0 1 12812
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_160
timestamp 1661296025
transform 1 0 5926 0 1 12394
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_161
timestamp 1661296025
transform 1 0 5926 0 1 12022
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_162
timestamp 1661296025
transform 1 0 5926 0 1 11604
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_163
timestamp 1661296025
transform 1 0 5926 0 1 11232
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_164
timestamp 1661296025
transform 1 0 5926 0 1 10814
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_165
timestamp 1661296025
transform 1 0 5926 0 1 10442
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_166
timestamp 1661296025
transform 1 0 5926 0 1 10024
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_167
timestamp 1661296025
transform 1 0 5926 0 1 9652
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_168
timestamp 1661296025
transform 1 0 5926 0 1 9234
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_169
timestamp 1661296025
transform 1 0 5926 0 1 8862
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_170
timestamp 1661296025
transform 1 0 5926 0 1 8444
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_171
timestamp 1661296025
transform 1 0 5926 0 1 8072
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_172
timestamp 1661296025
transform 1 0 5926 0 1 7654
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_173
timestamp 1661296025
transform 1 0 5926 0 1 7282
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_174
timestamp 1661296025
transform 1 0 5926 0 1 6864
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_175
timestamp 1661296025
transform 1 0 5926 0 1 6492
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_176
timestamp 1661296025
transform 1 0 5926 0 1 6074
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_177
timestamp 1661296025
transform 1 0 5926 0 1 5702
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_178
timestamp 1661296025
transform 1 0 5926 0 1 5284
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_179
timestamp 1661296025
transform 1 0 5926 0 1 4912
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_180
timestamp 1661296025
transform 1 0 5926 0 1 4494
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_181
timestamp 1661296025
transform 1 0 5926 0 1 4122
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_182
timestamp 1661296025
transform 1 0 5926 0 1 3704
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_183
timestamp 1661296025
transform 1 0 5926 0 1 3332
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_184
timestamp 1661296025
transform 1 0 5926 0 1 2914
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_185
timestamp 1661296025
transform 1 0 5926 0 1 2542
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_186
timestamp 1661296025
transform 1 0 5926 0 1 2124
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_187
timestamp 1661296025
transform 1 0 5926 0 1 1752
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_188
timestamp 1661296025
transform 1 0 5926 0 1 1334
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_189
timestamp 1661296025
transform 1 0 5926 0 1 962
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_190
timestamp 1661296025
transform 1 0 5926 0 1 544
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_191
timestamp 1661296025
transform 1 0 5926 0 1 172
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_192
timestamp 1661296025
transform 1 0 6694 0 1 25046
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_193
timestamp 1661296025
transform 1 0 6694 0 1 24650
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_194
timestamp 1661296025
transform 1 0 6694 0 1 24256
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_195
timestamp 1661296025
transform 1 0 6694 0 1 23860
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_196
timestamp 1661296025
transform 1 0 6694 0 1 23466
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_197
timestamp 1661296025
transform 1 0 6694 0 1 23070
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_198
timestamp 1661296025
transform 1 0 6694 0 1 22676
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_199
timestamp 1661296025
transform 1 0 6694 0 1 22280
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_200
timestamp 1661296025
transform 1 0 6694 0 1 21886
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_201
timestamp 1661296025
transform 1 0 6694 0 1 21490
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_202
timestamp 1661296025
transform 1 0 6694 0 1 21096
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_203
timestamp 1661296025
transform 1 0 6694 0 1 20700
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_204
timestamp 1661296025
transform 1 0 6694 0 1 20306
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_205
timestamp 1661296025
transform 1 0 6694 0 1 19910
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_206
timestamp 1661296025
transform 1 0 6694 0 1 19516
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_207
timestamp 1661296025
transform 1 0 6694 0 1 19120
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_208
timestamp 1661296025
transform 1 0 6694 0 1 18726
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_209
timestamp 1661296025
transform 1 0 6694 0 1 18330
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_210
timestamp 1661296025
transform 1 0 6694 0 1 17936
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_211
timestamp 1661296025
transform 1 0 6694 0 1 17540
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_212
timestamp 1661296025
transform 1 0 6694 0 1 17146
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_213
timestamp 1661296025
transform 1 0 6694 0 1 16750
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_214
timestamp 1661296025
transform 1 0 6694 0 1 16356
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_215
timestamp 1661296025
transform 1 0 6694 0 1 15960
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_216
timestamp 1661296025
transform 1 0 6694 0 1 15566
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_217
timestamp 1661296025
transform 1 0 6694 0 1 15170
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_218
timestamp 1661296025
transform 1 0 6694 0 1 14776
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_219
timestamp 1661296025
transform 1 0 6694 0 1 14380
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_220
timestamp 1661296025
transform 1 0 6694 0 1 13986
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_221
timestamp 1661296025
transform 1 0 6694 0 1 13590
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_222
timestamp 1661296025
transform 1 0 6694 0 1 13196
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_223
timestamp 1661296025
transform 1 0 6694 0 1 12800
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_224
timestamp 1661296025
transform 1 0 6694 0 1 12406
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_225
timestamp 1661296025
transform 1 0 6694 0 1 12010
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_226
timestamp 1661296025
transform 1 0 6694 0 1 11616
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_227
timestamp 1661296025
transform 1 0 6694 0 1 11220
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_228
timestamp 1661296025
transform 1 0 6694 0 1 10826
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_229
timestamp 1661296025
transform 1 0 6694 0 1 10430
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_230
timestamp 1661296025
transform 1 0 6694 0 1 10036
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_231
timestamp 1661296025
transform 1 0 6694 0 1 9640
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_232
timestamp 1661296025
transform 1 0 6694 0 1 9246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_233
timestamp 1661296025
transform 1 0 6694 0 1 8850
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_234
timestamp 1661296025
transform 1 0 6694 0 1 8456
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_235
timestamp 1661296025
transform 1 0 6694 0 1 8060
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_236
timestamp 1661296025
transform 1 0 6694 0 1 7666
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_237
timestamp 1661296025
transform 1 0 6694 0 1 7270
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_238
timestamp 1661296025
transform 1 0 6694 0 1 6876
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_239
timestamp 1661296025
transform 1 0 6694 0 1 6480
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_240
timestamp 1661296025
transform 1 0 6694 0 1 6086
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_241
timestamp 1661296025
transform 1 0 6694 0 1 5690
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_242
timestamp 1661296025
transform 1 0 6694 0 1 5296
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_243
timestamp 1661296025
transform 1 0 6694 0 1 4900
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_244
timestamp 1661296025
transform 1 0 6694 0 1 4506
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_245
timestamp 1661296025
transform 1 0 6694 0 1 4110
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_246
timestamp 1661296025
transform 1 0 6694 0 1 3716
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_247
timestamp 1661296025
transform 1 0 6694 0 1 3320
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_248
timestamp 1661296025
transform 1 0 6694 0 1 2926
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_249
timestamp 1661296025
transform 1 0 6694 0 1 2530
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_250
timestamp 1661296025
transform 1 0 6694 0 1 2136
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_251
timestamp 1661296025
transform 1 0 6694 0 1 1740
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_252
timestamp 1661296025
transform 1 0 6694 0 1 1346
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_253
timestamp 1661296025
transform 1 0 6694 0 1 950
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_254
timestamp 1661296025
transform 1 0 6694 0 1 556
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_255
timestamp 1661296025
transform 1 0 6694 0 1 160
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_256
timestamp 1661296025
transform 1 0 5494 0 1 25034
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_257
timestamp 1661296025
transform 1 0 5494 0 1 24662
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_258
timestamp 1661296025
transform 1 0 5494 0 1 24244
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_259
timestamp 1661296025
transform 1 0 5494 0 1 23872
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_260
timestamp 1661296025
transform 1 0 5494 0 1 23454
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_261
timestamp 1661296025
transform 1 0 5494 0 1 23082
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_262
timestamp 1661296025
transform 1 0 5494 0 1 22664
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_263
timestamp 1661296025
transform 1 0 5494 0 1 22292
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_264
timestamp 1661296025
transform 1 0 5494 0 1 21874
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_265
timestamp 1661296025
transform 1 0 5494 0 1 21502
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_266
timestamp 1661296025
transform 1 0 5494 0 1 21084
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_267
timestamp 1661296025
transform 1 0 5494 0 1 20712
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_268
timestamp 1661296025
transform 1 0 5494 0 1 20294
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_269
timestamp 1661296025
transform 1 0 5494 0 1 19922
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_270
timestamp 1661296025
transform 1 0 5494 0 1 19504
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_271
timestamp 1661296025
transform 1 0 5494 0 1 19132
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_272
timestamp 1661296025
transform 1 0 5494 0 1 18714
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_273
timestamp 1661296025
transform 1 0 5494 0 1 18342
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_274
timestamp 1661296025
transform 1 0 5494 0 1 17924
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_275
timestamp 1661296025
transform 1 0 5494 0 1 17552
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_276
timestamp 1661296025
transform 1 0 5494 0 1 17134
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_277
timestamp 1661296025
transform 1 0 5494 0 1 16762
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_278
timestamp 1661296025
transform 1 0 5494 0 1 16344
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_279
timestamp 1661296025
transform 1 0 5494 0 1 15972
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_280
timestamp 1661296025
transform 1 0 5494 0 1 15554
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_281
timestamp 1661296025
transform 1 0 5494 0 1 15182
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_282
timestamp 1661296025
transform 1 0 5494 0 1 14764
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_283
timestamp 1661296025
transform 1 0 5494 0 1 14392
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_284
timestamp 1661296025
transform 1 0 5494 0 1 13974
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_285
timestamp 1661296025
transform 1 0 5494 0 1 13602
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_286
timestamp 1661296025
transform 1 0 5494 0 1 13184
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_287
timestamp 1661296025
transform 1 0 5494 0 1 12812
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_288
timestamp 1661296025
transform 1 0 5494 0 1 12394
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_289
timestamp 1661296025
transform 1 0 5494 0 1 12022
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_290
timestamp 1661296025
transform 1 0 5494 0 1 11604
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_291
timestamp 1661296025
transform 1 0 5494 0 1 11232
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_292
timestamp 1661296025
transform 1 0 5494 0 1 10814
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_293
timestamp 1661296025
transform 1 0 5494 0 1 10442
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_294
timestamp 1661296025
transform 1 0 5494 0 1 10024
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_295
timestamp 1661296025
transform 1 0 5494 0 1 9652
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_296
timestamp 1661296025
transform 1 0 5494 0 1 9234
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_297
timestamp 1661296025
transform 1 0 5494 0 1 8862
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_298
timestamp 1661296025
transform 1 0 5494 0 1 8444
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_299
timestamp 1661296025
transform 1 0 5494 0 1 8072
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_300
timestamp 1661296025
transform 1 0 5494 0 1 7654
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_301
timestamp 1661296025
transform 1 0 5494 0 1 7282
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_302
timestamp 1661296025
transform 1 0 5494 0 1 6864
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_303
timestamp 1661296025
transform 1 0 5494 0 1 6492
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_304
timestamp 1661296025
transform 1 0 5494 0 1 6074
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_305
timestamp 1661296025
transform 1 0 5494 0 1 5702
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_306
timestamp 1661296025
transform 1 0 5494 0 1 5284
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_307
timestamp 1661296025
transform 1 0 5494 0 1 4912
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_308
timestamp 1661296025
transform 1 0 5494 0 1 4494
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_309
timestamp 1661296025
transform 1 0 5494 0 1 4122
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_310
timestamp 1661296025
transform 1 0 5494 0 1 3704
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_311
timestamp 1661296025
transform 1 0 5494 0 1 3332
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_312
timestamp 1661296025
transform 1 0 5494 0 1 2914
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_313
timestamp 1661296025
transform 1 0 5494 0 1 2542
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_314
timestamp 1661296025
transform 1 0 5494 0 1 2124
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_315
timestamp 1661296025
transform 1 0 5494 0 1 1752
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_316
timestamp 1661296025
transform 1 0 5494 0 1 1334
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_317
timestamp 1661296025
transform 1 0 5494 0 1 962
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_318
timestamp 1661296025
transform 1 0 5494 0 1 544
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_319
timestamp 1661296025
transform 1 0 5494 0 1 172
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_0
timestamp 1661296025
transform 1 0 5017 0 1 25038
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_1
timestamp 1661296025
transform 1 0 5017 0 1 24666
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_2
timestamp 1661296025
transform 1 0 5017 0 1 24248
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_3
timestamp 1661296025
transform 1 0 5017 0 1 23876
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_4
timestamp 1661296025
transform 1 0 5017 0 1 23458
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_5
timestamp 1661296025
transform 1 0 5017 0 1 23086
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_6
timestamp 1661296025
transform 1 0 5017 0 1 22668
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_7
timestamp 1661296025
transform 1 0 5017 0 1 22296
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_8
timestamp 1661296025
transform 1 0 5017 0 1 21878
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_9
timestamp 1661296025
transform 1 0 5017 0 1 21506
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_10
timestamp 1661296025
transform 1 0 5017 0 1 21088
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_11
timestamp 1661296025
transform 1 0 5017 0 1 20716
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_12
timestamp 1661296025
transform 1 0 5017 0 1 20298
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_13
timestamp 1661296025
transform 1 0 5017 0 1 19926
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_14
timestamp 1661296025
transform 1 0 5017 0 1 19508
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_15
timestamp 1661296025
transform 1 0 5017 0 1 19136
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_16
timestamp 1661296025
transform 1 0 5017 0 1 18718
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_17
timestamp 1661296025
transform 1 0 5017 0 1 18346
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_18
timestamp 1661296025
transform 1 0 5017 0 1 17928
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_19
timestamp 1661296025
transform 1 0 5017 0 1 17556
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_20
timestamp 1661296025
transform 1 0 5017 0 1 17138
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_21
timestamp 1661296025
transform 1 0 5017 0 1 16766
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_22
timestamp 1661296025
transform 1 0 5017 0 1 16348
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_23
timestamp 1661296025
transform 1 0 5017 0 1 15976
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_24
timestamp 1661296025
transform 1 0 5017 0 1 15558
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_25
timestamp 1661296025
transform 1 0 5017 0 1 15186
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_26
timestamp 1661296025
transform 1 0 5017 0 1 14768
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_27
timestamp 1661296025
transform 1 0 5017 0 1 14396
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_28
timestamp 1661296025
transform 1 0 5017 0 1 13978
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_29
timestamp 1661296025
transform 1 0 5017 0 1 13606
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_30
timestamp 1661296025
transform 1 0 5017 0 1 13188
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_31
timestamp 1661296025
transform 1 0 5017 0 1 12816
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_32
timestamp 1661296025
transform 1 0 5017 0 1 12398
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_33
timestamp 1661296025
transform 1 0 5017 0 1 12026
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_34
timestamp 1661296025
transform 1 0 5017 0 1 11608
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_35
timestamp 1661296025
transform 1 0 5017 0 1 11236
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_36
timestamp 1661296025
transform 1 0 5017 0 1 10818
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_37
timestamp 1661296025
transform 1 0 5017 0 1 10446
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_38
timestamp 1661296025
transform 1 0 5017 0 1 10028
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_39
timestamp 1661296025
transform 1 0 5017 0 1 9656
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_40
timestamp 1661296025
transform 1 0 5017 0 1 9238
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_41
timestamp 1661296025
transform 1 0 5017 0 1 8866
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_42
timestamp 1661296025
transform 1 0 5017 0 1 8448
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_43
timestamp 1661296025
transform 1 0 5017 0 1 8076
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_44
timestamp 1661296025
transform 1 0 5017 0 1 7658
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_45
timestamp 1661296025
transform 1 0 5017 0 1 7286
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_46
timestamp 1661296025
transform 1 0 5017 0 1 6868
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_47
timestamp 1661296025
transform 1 0 5017 0 1 6496
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_48
timestamp 1661296025
transform 1 0 5017 0 1 6078
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_49
timestamp 1661296025
transform 1 0 5017 0 1 5706
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_50
timestamp 1661296025
transform 1 0 5017 0 1 5288
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_51
timestamp 1661296025
transform 1 0 5017 0 1 4916
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_52
timestamp 1661296025
transform 1 0 5017 0 1 4498
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_53
timestamp 1661296025
transform 1 0 5017 0 1 4126
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_54
timestamp 1661296025
transform 1 0 5017 0 1 3708
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_55
timestamp 1661296025
transform 1 0 5017 0 1 3336
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_56
timestamp 1661296025
transform 1 0 5017 0 1 2918
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_57
timestamp 1661296025
transform 1 0 5017 0 1 2546
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_58
timestamp 1661296025
transform 1 0 5017 0 1 2128
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_59
timestamp 1661296025
transform 1 0 5017 0 1 1756
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_60
timestamp 1661296025
transform 1 0 5017 0 1 1338
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_61
timestamp 1661296025
transform 1 0 5017 0 1 966
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_62
timestamp 1661296025
transform 1 0 5017 0 1 548
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_63
timestamp 1661296025
transform 1 0 5017 0 1 176
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_64
timestamp 1661296025
transform 1 0 6265 0 1 25050
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_65
timestamp 1661296025
transform 1 0 6265 0 1 24654
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_66
timestamp 1661296025
transform 1 0 6265 0 1 24260
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_67
timestamp 1661296025
transform 1 0 6265 0 1 23864
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_68
timestamp 1661296025
transform 1 0 6265 0 1 23470
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_69
timestamp 1661296025
transform 1 0 6265 0 1 23074
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_70
timestamp 1661296025
transform 1 0 6265 0 1 22680
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_71
timestamp 1661296025
transform 1 0 6265 0 1 22284
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_72
timestamp 1661296025
transform 1 0 6265 0 1 21890
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_73
timestamp 1661296025
transform 1 0 6265 0 1 21494
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_74
timestamp 1661296025
transform 1 0 6265 0 1 21100
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_75
timestamp 1661296025
transform 1 0 6265 0 1 20704
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_76
timestamp 1661296025
transform 1 0 6265 0 1 20310
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_77
timestamp 1661296025
transform 1 0 6265 0 1 19914
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_78
timestamp 1661296025
transform 1 0 6265 0 1 19520
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_79
timestamp 1661296025
transform 1 0 6265 0 1 19124
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_80
timestamp 1661296025
transform 1 0 6265 0 1 18730
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_81
timestamp 1661296025
transform 1 0 6265 0 1 18334
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_82
timestamp 1661296025
transform 1 0 6265 0 1 17940
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_83
timestamp 1661296025
transform 1 0 6265 0 1 17544
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_84
timestamp 1661296025
transform 1 0 6265 0 1 17150
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_85
timestamp 1661296025
transform 1 0 6265 0 1 16754
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_86
timestamp 1661296025
transform 1 0 6265 0 1 16360
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_87
timestamp 1661296025
transform 1 0 6265 0 1 15964
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_88
timestamp 1661296025
transform 1 0 6265 0 1 15570
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_89
timestamp 1661296025
transform 1 0 6265 0 1 15174
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_90
timestamp 1661296025
transform 1 0 6265 0 1 14780
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_91
timestamp 1661296025
transform 1 0 6265 0 1 14384
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_92
timestamp 1661296025
transform 1 0 6265 0 1 13990
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_93
timestamp 1661296025
transform 1 0 6265 0 1 13594
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_94
timestamp 1661296025
transform 1 0 6265 0 1 13200
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_95
timestamp 1661296025
transform 1 0 6265 0 1 12804
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_96
timestamp 1661296025
transform 1 0 6265 0 1 12410
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_97
timestamp 1661296025
transform 1 0 6265 0 1 12014
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_98
timestamp 1661296025
transform 1 0 6265 0 1 11620
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_99
timestamp 1661296025
transform 1 0 6265 0 1 11224
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_100
timestamp 1661296025
transform 1 0 6265 0 1 10830
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_101
timestamp 1661296025
transform 1 0 6265 0 1 10434
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_102
timestamp 1661296025
transform 1 0 6265 0 1 10040
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_103
timestamp 1661296025
transform 1 0 6265 0 1 9644
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_104
timestamp 1661296025
transform 1 0 6265 0 1 9250
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_105
timestamp 1661296025
transform 1 0 6265 0 1 8854
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_106
timestamp 1661296025
transform 1 0 6265 0 1 8460
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_107
timestamp 1661296025
transform 1 0 6265 0 1 8064
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_108
timestamp 1661296025
transform 1 0 6265 0 1 7670
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_109
timestamp 1661296025
transform 1 0 6265 0 1 7274
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_110
timestamp 1661296025
transform 1 0 6265 0 1 6880
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_111
timestamp 1661296025
transform 1 0 6265 0 1 6484
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_112
timestamp 1661296025
transform 1 0 6265 0 1 6090
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_113
timestamp 1661296025
transform 1 0 6265 0 1 5694
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_114
timestamp 1661296025
transform 1 0 6265 0 1 5300
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_115
timestamp 1661296025
transform 1 0 6265 0 1 4904
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_116
timestamp 1661296025
transform 1 0 6265 0 1 4510
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_117
timestamp 1661296025
transform 1 0 6265 0 1 4114
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_118
timestamp 1661296025
transform 1 0 6265 0 1 3720
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_119
timestamp 1661296025
transform 1 0 6265 0 1 3324
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_120
timestamp 1661296025
transform 1 0 6265 0 1 2930
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_121
timestamp 1661296025
transform 1 0 6265 0 1 2534
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_122
timestamp 1661296025
transform 1 0 6265 0 1 2140
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_123
timestamp 1661296025
transform 1 0 6265 0 1 1744
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_124
timestamp 1661296025
transform 1 0 6265 0 1 1350
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_125
timestamp 1661296025
transform 1 0 6265 0 1 954
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_126
timestamp 1661296025
transform 1 0 6265 0 1 560
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_127
timestamp 1661296025
transform 1 0 6265 0 1 164
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_128
timestamp 1661296025
transform 1 0 5921 0 1 25038
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_129
timestamp 1661296025
transform 1 0 5921 0 1 24666
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_130
timestamp 1661296025
transform 1 0 5921 0 1 24248
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_131
timestamp 1661296025
transform 1 0 5921 0 1 23876
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_132
timestamp 1661296025
transform 1 0 5921 0 1 23458
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_133
timestamp 1661296025
transform 1 0 5921 0 1 23086
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_134
timestamp 1661296025
transform 1 0 5921 0 1 22668
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_135
timestamp 1661296025
transform 1 0 5921 0 1 22296
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_136
timestamp 1661296025
transform 1 0 5921 0 1 21878
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_137
timestamp 1661296025
transform 1 0 5921 0 1 21506
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_138
timestamp 1661296025
transform 1 0 5921 0 1 21088
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_139
timestamp 1661296025
transform 1 0 5921 0 1 20716
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_140
timestamp 1661296025
transform 1 0 5921 0 1 20298
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_141
timestamp 1661296025
transform 1 0 5921 0 1 19926
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_142
timestamp 1661296025
transform 1 0 5921 0 1 19508
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_143
timestamp 1661296025
transform 1 0 5921 0 1 19136
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_144
timestamp 1661296025
transform 1 0 5921 0 1 18718
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_145
timestamp 1661296025
transform 1 0 5921 0 1 18346
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_146
timestamp 1661296025
transform 1 0 5921 0 1 17928
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_147
timestamp 1661296025
transform 1 0 5921 0 1 17556
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_148
timestamp 1661296025
transform 1 0 5921 0 1 17138
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_149
timestamp 1661296025
transform 1 0 5921 0 1 16766
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_150
timestamp 1661296025
transform 1 0 5921 0 1 16348
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_151
timestamp 1661296025
transform 1 0 5921 0 1 15976
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_152
timestamp 1661296025
transform 1 0 5921 0 1 15558
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_153
timestamp 1661296025
transform 1 0 5921 0 1 15186
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_154
timestamp 1661296025
transform 1 0 5921 0 1 14768
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_155
timestamp 1661296025
transform 1 0 5921 0 1 14396
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_156
timestamp 1661296025
transform 1 0 5921 0 1 13978
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_157
timestamp 1661296025
transform 1 0 5921 0 1 13606
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_158
timestamp 1661296025
transform 1 0 5921 0 1 13188
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_159
timestamp 1661296025
transform 1 0 5921 0 1 12816
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_160
timestamp 1661296025
transform 1 0 5921 0 1 12398
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_161
timestamp 1661296025
transform 1 0 5921 0 1 12026
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_162
timestamp 1661296025
transform 1 0 5921 0 1 11608
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_163
timestamp 1661296025
transform 1 0 5921 0 1 11236
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_164
timestamp 1661296025
transform 1 0 5921 0 1 10818
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_165
timestamp 1661296025
transform 1 0 5921 0 1 10446
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_166
timestamp 1661296025
transform 1 0 5921 0 1 10028
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_167
timestamp 1661296025
transform 1 0 5921 0 1 9656
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_168
timestamp 1661296025
transform 1 0 5921 0 1 9238
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_169
timestamp 1661296025
transform 1 0 5921 0 1 8866
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_170
timestamp 1661296025
transform 1 0 5921 0 1 8448
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_171
timestamp 1661296025
transform 1 0 5921 0 1 8076
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_172
timestamp 1661296025
transform 1 0 5921 0 1 7658
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_173
timestamp 1661296025
transform 1 0 5921 0 1 7286
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_174
timestamp 1661296025
transform 1 0 5921 0 1 6868
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_175
timestamp 1661296025
transform 1 0 5921 0 1 6496
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_176
timestamp 1661296025
transform 1 0 5921 0 1 6078
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_177
timestamp 1661296025
transform 1 0 5921 0 1 5706
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_178
timestamp 1661296025
transform 1 0 5921 0 1 5288
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_179
timestamp 1661296025
transform 1 0 5921 0 1 4916
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_180
timestamp 1661296025
transform 1 0 5921 0 1 4498
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_181
timestamp 1661296025
transform 1 0 5921 0 1 4126
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_182
timestamp 1661296025
transform 1 0 5921 0 1 3708
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_183
timestamp 1661296025
transform 1 0 5921 0 1 3336
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_184
timestamp 1661296025
transform 1 0 5921 0 1 2918
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_185
timestamp 1661296025
transform 1 0 5921 0 1 2546
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_186
timestamp 1661296025
transform 1 0 5921 0 1 2128
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_187
timestamp 1661296025
transform 1 0 5921 0 1 1756
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_188
timestamp 1661296025
transform 1 0 5921 0 1 1338
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_189
timestamp 1661296025
transform 1 0 5921 0 1 966
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_190
timestamp 1661296025
transform 1 0 5921 0 1 548
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_191
timestamp 1661296025
transform 1 0 5921 0 1 176
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_192
timestamp 1661296025
transform 1 0 6689 0 1 25050
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_193
timestamp 1661296025
transform 1 0 6689 0 1 24654
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_194
timestamp 1661296025
transform 1 0 6689 0 1 24260
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_195
timestamp 1661296025
transform 1 0 6689 0 1 23864
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_196
timestamp 1661296025
transform 1 0 6689 0 1 23470
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_197
timestamp 1661296025
transform 1 0 6689 0 1 23074
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_198
timestamp 1661296025
transform 1 0 6689 0 1 22680
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_199
timestamp 1661296025
transform 1 0 6689 0 1 22284
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_200
timestamp 1661296025
transform 1 0 6689 0 1 21890
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_201
timestamp 1661296025
transform 1 0 6689 0 1 21494
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_202
timestamp 1661296025
transform 1 0 6689 0 1 21100
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_203
timestamp 1661296025
transform 1 0 6689 0 1 20704
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_204
timestamp 1661296025
transform 1 0 6689 0 1 20310
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_205
timestamp 1661296025
transform 1 0 6689 0 1 19914
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_206
timestamp 1661296025
transform 1 0 6689 0 1 19520
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_207
timestamp 1661296025
transform 1 0 6689 0 1 19124
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_208
timestamp 1661296025
transform 1 0 6689 0 1 18730
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_209
timestamp 1661296025
transform 1 0 6689 0 1 18334
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_210
timestamp 1661296025
transform 1 0 6689 0 1 17940
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_211
timestamp 1661296025
transform 1 0 6689 0 1 17544
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_212
timestamp 1661296025
transform 1 0 6689 0 1 17150
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_213
timestamp 1661296025
transform 1 0 6689 0 1 16754
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_214
timestamp 1661296025
transform 1 0 6689 0 1 16360
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_215
timestamp 1661296025
transform 1 0 6689 0 1 15964
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_216
timestamp 1661296025
transform 1 0 6689 0 1 15570
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_217
timestamp 1661296025
transform 1 0 6689 0 1 15174
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_218
timestamp 1661296025
transform 1 0 6689 0 1 14780
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_219
timestamp 1661296025
transform 1 0 6689 0 1 14384
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_220
timestamp 1661296025
transform 1 0 6689 0 1 13990
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_221
timestamp 1661296025
transform 1 0 6689 0 1 13594
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_222
timestamp 1661296025
transform 1 0 6689 0 1 13200
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_223
timestamp 1661296025
transform 1 0 6689 0 1 12804
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_224
timestamp 1661296025
transform 1 0 6689 0 1 12410
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_225
timestamp 1661296025
transform 1 0 6689 0 1 12014
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_226
timestamp 1661296025
transform 1 0 6689 0 1 11620
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_227
timestamp 1661296025
transform 1 0 6689 0 1 11224
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_228
timestamp 1661296025
transform 1 0 6689 0 1 10830
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_229
timestamp 1661296025
transform 1 0 6689 0 1 10434
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_230
timestamp 1661296025
transform 1 0 6689 0 1 10040
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_231
timestamp 1661296025
transform 1 0 6689 0 1 9644
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_232
timestamp 1661296025
transform 1 0 6689 0 1 9250
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_233
timestamp 1661296025
transform 1 0 6689 0 1 8854
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_234
timestamp 1661296025
transform 1 0 6689 0 1 8460
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_235
timestamp 1661296025
transform 1 0 6689 0 1 8064
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_236
timestamp 1661296025
transform 1 0 6689 0 1 7670
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_237
timestamp 1661296025
transform 1 0 6689 0 1 7274
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_238
timestamp 1661296025
transform 1 0 6689 0 1 6880
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_239
timestamp 1661296025
transform 1 0 6689 0 1 6484
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_240
timestamp 1661296025
transform 1 0 6689 0 1 6090
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_241
timestamp 1661296025
transform 1 0 6689 0 1 5694
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_242
timestamp 1661296025
transform 1 0 6689 0 1 5300
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_243
timestamp 1661296025
transform 1 0 6689 0 1 4904
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_244
timestamp 1661296025
transform 1 0 6689 0 1 4510
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_245
timestamp 1661296025
transform 1 0 6689 0 1 4114
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_246
timestamp 1661296025
transform 1 0 6689 0 1 3720
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_247
timestamp 1661296025
transform 1 0 6689 0 1 3324
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_248
timestamp 1661296025
transform 1 0 6689 0 1 2930
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_249
timestamp 1661296025
transform 1 0 6689 0 1 2534
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_250
timestamp 1661296025
transform 1 0 6689 0 1 2140
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_251
timestamp 1661296025
transform 1 0 6689 0 1 1744
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_252
timestamp 1661296025
transform 1 0 6689 0 1 1350
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_253
timestamp 1661296025
transform 1 0 6689 0 1 954
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_254
timestamp 1661296025
transform 1 0 6689 0 1 560
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_255
timestamp 1661296025
transform 1 0 6689 0 1 164
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_256
timestamp 1661296025
transform 1 0 5489 0 1 25038
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_257
timestamp 1661296025
transform 1 0 5489 0 1 24666
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_258
timestamp 1661296025
transform 1 0 5489 0 1 24248
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_259
timestamp 1661296025
transform 1 0 5489 0 1 23876
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_260
timestamp 1661296025
transform 1 0 5489 0 1 23458
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_261
timestamp 1661296025
transform 1 0 5489 0 1 23086
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_262
timestamp 1661296025
transform 1 0 5489 0 1 22668
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_263
timestamp 1661296025
transform 1 0 5489 0 1 22296
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_264
timestamp 1661296025
transform 1 0 5489 0 1 21878
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_265
timestamp 1661296025
transform 1 0 5489 0 1 21506
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_266
timestamp 1661296025
transform 1 0 5489 0 1 21088
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_267
timestamp 1661296025
transform 1 0 5489 0 1 20716
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_268
timestamp 1661296025
transform 1 0 5489 0 1 20298
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_269
timestamp 1661296025
transform 1 0 5489 0 1 19926
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_270
timestamp 1661296025
transform 1 0 5489 0 1 19508
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_271
timestamp 1661296025
transform 1 0 5489 0 1 19136
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_272
timestamp 1661296025
transform 1 0 5489 0 1 18718
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_273
timestamp 1661296025
transform 1 0 5489 0 1 18346
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_274
timestamp 1661296025
transform 1 0 5489 0 1 17928
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_275
timestamp 1661296025
transform 1 0 5489 0 1 17556
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_276
timestamp 1661296025
transform 1 0 5489 0 1 17138
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_277
timestamp 1661296025
transform 1 0 5489 0 1 16766
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_278
timestamp 1661296025
transform 1 0 5489 0 1 16348
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_279
timestamp 1661296025
transform 1 0 5489 0 1 15976
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_280
timestamp 1661296025
transform 1 0 5489 0 1 15558
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_281
timestamp 1661296025
transform 1 0 5489 0 1 15186
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_282
timestamp 1661296025
transform 1 0 5489 0 1 14768
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_283
timestamp 1661296025
transform 1 0 5489 0 1 14396
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_284
timestamp 1661296025
transform 1 0 5489 0 1 13978
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_285
timestamp 1661296025
transform 1 0 5489 0 1 13606
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_286
timestamp 1661296025
transform 1 0 5489 0 1 13188
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_287
timestamp 1661296025
transform 1 0 5489 0 1 12816
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_288
timestamp 1661296025
transform 1 0 5489 0 1 12398
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_289
timestamp 1661296025
transform 1 0 5489 0 1 12026
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_290
timestamp 1661296025
transform 1 0 5489 0 1 11608
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_291
timestamp 1661296025
transform 1 0 5489 0 1 11236
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_292
timestamp 1661296025
transform 1 0 5489 0 1 10818
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_293
timestamp 1661296025
transform 1 0 5489 0 1 10446
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_294
timestamp 1661296025
transform 1 0 5489 0 1 10028
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_295
timestamp 1661296025
transform 1 0 5489 0 1 9656
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_296
timestamp 1661296025
transform 1 0 5489 0 1 9238
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_297
timestamp 1661296025
transform 1 0 5489 0 1 8866
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_298
timestamp 1661296025
transform 1 0 5489 0 1 8448
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_299
timestamp 1661296025
transform 1 0 5489 0 1 8076
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_300
timestamp 1661296025
transform 1 0 5489 0 1 7658
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_301
timestamp 1661296025
transform 1 0 5489 0 1 7286
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_302
timestamp 1661296025
transform 1 0 5489 0 1 6868
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_303
timestamp 1661296025
transform 1 0 5489 0 1 6496
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_304
timestamp 1661296025
transform 1 0 5489 0 1 6078
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_305
timestamp 1661296025
transform 1 0 5489 0 1 5706
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_306
timestamp 1661296025
transform 1 0 5489 0 1 5288
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_307
timestamp 1661296025
transform 1 0 5489 0 1 4916
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_308
timestamp 1661296025
transform 1 0 5489 0 1 4498
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_309
timestamp 1661296025
transform 1 0 5489 0 1 4126
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_310
timestamp 1661296025
transform 1 0 5489 0 1 3708
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_311
timestamp 1661296025
transform 1 0 5489 0 1 3336
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_312
timestamp 1661296025
transform 1 0 5489 0 1 2918
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_313
timestamp 1661296025
transform 1 0 5489 0 1 2546
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_314
timestamp 1661296025
transform 1 0 5489 0 1 2128
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_315
timestamp 1661296025
transform 1 0 5489 0 1 1756
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_316
timestamp 1661296025
transform 1 0 5489 0 1 1338
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_317
timestamp 1661296025
transform 1 0 5489 0 1 966
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_318
timestamp 1661296025
transform 1 0 5489 0 1 548
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_319
timestamp 1661296025
transform 1 0 5489 0 1 176
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_hierarchical_predecode2x4  sky130_sram_1r1w_24x128_8_hierarchical_predecode2x4_0
timestamp 1661296025
transform 1 0 527 0 1 4740
box 61 -56 3178 1636
use sky130_sram_1r1w_24x128_8_hierarchical_predecode2x4  sky130_sram_1r1w_24x128_8_hierarchical_predecode2x4_1
timestamp 1661296025
transform 1 0 527 0 1 2370
box 61 -56 3178 1636
use sky130_sram_1r1w_24x128_8_hierarchical_predecode2x4  sky130_sram_1r1w_24x128_8_hierarchical_predecode2x4_2
timestamp 1661296025
transform 1 0 527 0 1 0
box 61 -56 3178 1636
<< labels >>
rlabel metal1 s 19 0 47 6320 4 addr_0
port 1 nsew
rlabel metal1 s 99 0 127 6320 4 addr_1
port 2 nsew
rlabel metal1 s 179 0 207 6320 4 addr_2
port 3 nsew
rlabel metal1 s 259 0 287 6320 4 addr_3
port 4 nsew
rlabel metal1 s 339 0 367 6320 4 addr_4
port 5 nsew
rlabel metal1 s 419 0 447 6320 4 addr_5
port 6 nsew
rlabel locali s 6572 120 6572 120 4 decode_0
port 7 nsew
rlabel locali s 6572 670 6572 670 4 decode_1
port 8 nsew
rlabel locali s 6572 910 6572 910 4 decode_2
port 9 nsew
rlabel locali s 6572 1460 6572 1460 4 decode_3
port 10 nsew
rlabel locali s 6572 1700 6572 1700 4 decode_4
port 11 nsew
rlabel locali s 6572 2250 6572 2250 4 decode_5
port 12 nsew
rlabel locali s 6572 2490 6572 2490 4 decode_6
port 13 nsew
rlabel locali s 6572 3040 6572 3040 4 decode_7
port 14 nsew
rlabel locali s 6572 3280 6572 3280 4 decode_8
port 15 nsew
rlabel locali s 6572 3830 6572 3830 4 decode_9
port 16 nsew
rlabel locali s 6572 4070 6572 4070 4 decode_10
port 17 nsew
rlabel locali s 6572 4620 6572 4620 4 decode_11
port 18 nsew
rlabel locali s 6572 4860 6572 4860 4 decode_12
port 19 nsew
rlabel locali s 6572 5410 6572 5410 4 decode_13
port 20 nsew
rlabel locali s 6572 5650 6572 5650 4 decode_14
port 21 nsew
rlabel locali s 6572 6200 6572 6200 4 decode_15
port 22 nsew
rlabel locali s 6572 6440 6572 6440 4 decode_16
port 23 nsew
rlabel locali s 6572 6990 6572 6990 4 decode_17
port 24 nsew
rlabel locali s 6572 7230 6572 7230 4 decode_18
port 25 nsew
rlabel locali s 6572 7780 6572 7780 4 decode_19
port 26 nsew
rlabel locali s 6572 8020 6572 8020 4 decode_20
port 27 nsew
rlabel locali s 6572 8570 6572 8570 4 decode_21
port 28 nsew
rlabel locali s 6572 8810 6572 8810 4 decode_22
port 29 nsew
rlabel locali s 6572 9360 6572 9360 4 decode_23
port 30 nsew
rlabel locali s 6572 9600 6572 9600 4 decode_24
port 31 nsew
rlabel locali s 6572 10150 6572 10150 4 decode_25
port 32 nsew
rlabel locali s 6572 10390 6572 10390 4 decode_26
port 33 nsew
rlabel locali s 6572 10940 6572 10940 4 decode_27
port 34 nsew
rlabel locali s 6572 11180 6572 11180 4 decode_28
port 35 nsew
rlabel locali s 6572 11730 6572 11730 4 decode_29
port 36 nsew
rlabel locali s 6572 11970 6572 11970 4 decode_30
port 37 nsew
rlabel locali s 6572 12520 6572 12520 4 decode_31
port 38 nsew
rlabel locali s 6572 12760 6572 12760 4 decode_32
port 39 nsew
rlabel locali s 6572 13310 6572 13310 4 decode_33
port 40 nsew
rlabel locali s 6572 13550 6572 13550 4 decode_34
port 41 nsew
rlabel locali s 6572 14100 6572 14100 4 decode_35
port 42 nsew
rlabel locali s 6572 14340 6572 14340 4 decode_36
port 43 nsew
rlabel locali s 6572 14890 6572 14890 4 decode_37
port 44 nsew
rlabel locali s 6572 15130 6572 15130 4 decode_38
port 45 nsew
rlabel locali s 6572 15680 6572 15680 4 decode_39
port 46 nsew
rlabel locali s 6572 15920 6572 15920 4 decode_40
port 47 nsew
rlabel locali s 6572 16470 6572 16470 4 decode_41
port 48 nsew
rlabel locali s 6572 16710 6572 16710 4 decode_42
port 49 nsew
rlabel locali s 6572 17260 6572 17260 4 decode_43
port 50 nsew
rlabel locali s 6572 17500 6572 17500 4 decode_44
port 51 nsew
rlabel locali s 6572 18050 6572 18050 4 decode_45
port 52 nsew
rlabel locali s 6572 18290 6572 18290 4 decode_46
port 53 nsew
rlabel locali s 6572 18840 6572 18840 4 decode_47
port 54 nsew
rlabel locali s 6572 19080 6572 19080 4 decode_48
port 55 nsew
rlabel locali s 6572 19630 6572 19630 4 decode_49
port 56 nsew
rlabel locali s 6572 19870 6572 19870 4 decode_50
port 57 nsew
rlabel locali s 6572 20420 6572 20420 4 decode_51
port 58 nsew
rlabel locali s 6572 20660 6572 20660 4 decode_52
port 59 nsew
rlabel locali s 6572 21210 6572 21210 4 decode_53
port 60 nsew
rlabel locali s 6572 21450 6572 21450 4 decode_54
port 61 nsew
rlabel locali s 6572 22000 6572 22000 4 decode_55
port 62 nsew
rlabel locali s 6572 22240 6572 22240 4 decode_56
port 63 nsew
rlabel locali s 6572 22790 6572 22790 4 decode_57
port 64 nsew
rlabel locali s 6572 23030 6572 23030 4 decode_58
port 65 nsew
rlabel locali s 6572 23580 6572 23580 4 decode_59
port 66 nsew
rlabel locali s 6572 23820 6572 23820 4 decode_60
port 67 nsew
rlabel locali s 6572 24370 6572 24370 4 decode_61
port 68 nsew
rlabel locali s 6572 24610 6572 24610 4 decode_62
port 69 nsew
rlabel locali s 6572 25160 6572 25160 4 decode_63
port 70 nsew
rlabel metal4 s 6694 -33 6760 25341 4 vdd
port 71 nsew
rlabel metal3 s 1392 5086 1490 5184 4 vdd
port 71 nsew
rlabel metal3 s 2715 2723 2813 2821 4 vdd
port 71 nsew
rlabel metal3 s 1392 2716 1490 2814 4 vdd
port 71 nsew
rlabel metal3 s 1392 346 1490 444 4 vdd
port 71 nsew
rlabel metal3 s 3490 1136 3588 1234 4 vdd
port 71 nsew
rlabel metal3 s 2715 3513 2813 3611 4 vdd
port 71 nsew
rlabel metal3 s 3490 5876 3588 5974 4 vdd
port 71 nsew
rlabel metal3 s 3490 3506 3588 3604 4 vdd
port 71 nsew
rlabel metal3 s 2715 1143 2813 1241 4 vdd
port 71 nsew
rlabel metal4 s 5494 -33 5560 25341 4 vdd
port 71 nsew
rlabel metal4 s 5926 -33 5992 25341 4 vdd
port 71 nsew
rlabel metal3 s 3490 346 3588 444 4 vdd
port 71 nsew
rlabel metal3 s 3490 5086 3588 5184 4 vdd
port 71 nsew
rlabel metal3 s 2715 353 2813 451 4 vdd
port 71 nsew
rlabel metal3 s 3490 2716 3588 2814 4 vdd
port 71 nsew
rlabel metal3 s 2715 5093 2813 5191 4 vdd
port 71 nsew
rlabel metal3 s 2715 5883 2813 5981 4 vdd
port 71 nsew
rlabel metal3 s 3094 3506 3192 3604 4 gnd
port 72 nsew
rlabel metal3 s 2290 2723 2388 2821 4 gnd
port 72 nsew
rlabel metal4 s 6270 -33 6336 25341 4 gnd
port 72 nsew
rlabel metal3 s 2290 353 2388 451 4 gnd
port 72 nsew
rlabel metal3 s 3094 346 3192 444 4 gnd
port 72 nsew
rlabel metal3 s 3094 5086 3192 5184 4 gnd
port 72 nsew
rlabel metal3 s 996 5086 1094 5184 4 gnd
port 72 nsew
rlabel metal3 s 2290 5093 2388 5191 4 gnd
port 72 nsew
rlabel metal3 s 3094 5876 3192 5974 4 gnd
port 72 nsew
rlabel metal3 s 3094 2716 3192 2814 4 gnd
port 72 nsew
rlabel metal3 s 2290 1143 2388 1241 4 gnd
port 72 nsew
rlabel metal3 s 996 346 1094 444 4 gnd
port 72 nsew
rlabel metal3 s 2290 3513 2388 3611 4 gnd
port 72 nsew
rlabel metal3 s 3094 1136 3192 1234 4 gnd
port 72 nsew
rlabel metal3 s 2290 5883 2388 5981 4 gnd
port 72 nsew
rlabel metal3 s 996 2716 1094 2814 4 gnd
port 72 nsew
rlabel metal4 s 5022 -33 5088 25341 4 gnd
port 72 nsew
<< properties >>
string FIXED_BBOX 0 0 6861 25308
<< end >>
