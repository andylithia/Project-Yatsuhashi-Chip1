magic
tech sky130B
magscale 1 2
timestamp 1660526289
<< metal4 >>
rect -28400 -4112 -14600 -4000
rect -28400 -7888 -28288 -4112
rect -24512 -7888 -18488 -4112
rect -14712 -7888 -14600 -4112
rect -28400 -8000 -14600 -7888
<< via4 >>
rect -28288 -7888 -24512 -4112
rect -18488 -7888 -14712 -4112
<< metal5 >>
tri -15074 20906 -12980 23000 se
rect -12980 20906 8380 23000
tri 8380 20906 10474 23000 sw
tri -16980 19000 -15074 20906 se
rect -15074 19000 10474 20906
tri 10474 19000 12380 20906 sw
tri -19200 16780 -16980 19000 se
rect -16980 18400 -11923 19000
tri -11923 18400 -11323 19000 nw
tri 6723 18400 7323 19000 ne
rect 7323 18400 12380 19000
rect -16980 17551 -12772 18400
tri -12772 17551 -11923 18400 nw
tri -11923 17551 -11074 18400 se
rect -11074 17551 6474 18400
tri 6474 17551 7323 18400 sw
tri 7323 17551 8172 18400 ne
rect 8172 17551 12380 18400
rect -16980 16780 -13621 17551
tri -20731 15249 -19200 16780 se
rect -19200 16702 -13621 16780
tri -13621 16702 -12772 17551 nw
tri -12772 16702 -11923 17551 se
rect -11923 16702 7323 17551
tri 7323 16702 8172 17551 sw
tri 8172 16702 9021 17551 ne
rect 9021 16702 12380 17551
rect -19200 16098 -14225 16702
tri -14225 16098 -13621 16702 nw
tri -13376 16098 -12772 16702 se
rect -12772 16098 8172 16702
tri 8172 16098 8776 16702 sw
tri 9021 16098 9625 16702 ne
rect 9625 16098 12380 16702
rect -19200 15249 -15074 16098
tri -15074 15249 -14225 16098 nw
tri -14225 15249 -13376 16098 se
rect -13376 15249 8776 16098
tri 8776 15249 9625 16098 sw
tri 9625 15249 10474 16098 ne
rect 10474 15249 12380 16098
tri -23800 12180 -20731 15249 se
rect -20731 14400 -15923 15249
tri -15923 14400 -15074 15249 nw
tri -15074 14400 -14225 15249 se
rect -14225 14400 9625 15249
tri 9625 14400 10474 15249 sw
tri 10474 14400 11323 15249 ne
rect 11323 14400 12380 15249
tri 12380 14400 16980 19000 sw
rect -20731 13551 -16772 14400
tri -16772 13551 -15923 14400 nw
tri -15923 13551 -15074 14400 se
rect -15074 13551 -13543 14400
rect -20731 12702 -17621 13551
tri -17621 12702 -16772 13551 nw
tri -16772 12702 -15923 13551 se
rect -15923 12702 -13543 13551
rect -20731 12180 -18351 12702
tri -24857 11123 -23800 12180 se
rect -23800 11972 -18351 12180
tri -18351 11972 -17621 12702 nw
tri -17502 11972 -16772 12702 se
rect -16772 11972 -13543 12702
rect -23800 11123 -19200 11972
tri -19200 11123 -18351 11972 nw
tri -18351 11123 -17502 11972 se
rect -17502 11123 -13543 11972
tri -27800 8180 -24857 11123 se
rect -24857 10274 -20049 11123
tri -20049 10274 -19200 11123 nw
tri -19200 10274 -18351 11123 se
rect -18351 10274 -13543 11123
tri -13543 10274 -9417 14400 nw
tri 4817 10274 8943 14400 ne
rect 8943 13551 10474 14400
tri 10474 13551 11323 14400 sw
tri 11323 13551 12172 14400 ne
rect 12172 13551 16980 14400
rect 8943 12702 11323 13551
tri 11323 12702 12172 13551 sw
tri 12172 12702 13021 13551 ne
rect 13021 12702 16980 13551
rect 8943 11972 12172 12702
tri 12172 11972 12902 12702 sw
tri 13021 11972 13751 12702 ne
rect 13751 11972 16980 12702
rect 8943 11123 12902 11972
tri 12902 11123 13751 11972 sw
tri 13751 11123 14600 11972 ne
rect 14600 11123 16980 11972
rect 8943 10274 13751 11123
tri 13751 10274 14600 11123 sw
tri 14600 10274 15449 11123 ne
rect 15449 10274 16980 11123
tri 16980 10274 21106 14400 sw
rect -24857 9425 -20898 10274
tri -20898 9425 -20049 10274 nw
tri -20049 9425 -19200 10274 se
rect -19200 9425 -15074 10274
rect -24857 8743 -21580 9425
tri -21580 8743 -20898 9425 nw
tri -20731 8743 -20049 9425 se
rect -20049 8743 -15074 9425
tri -15074 8743 -13543 10274 nw
tri 8943 8743 10474 10274 ne
rect 10474 9425 14600 10274
tri 14600 9425 15449 10274 sw
tri 15449 9425 16298 10274 ne
rect 16298 9425 21106 10274
rect 10474 8743 15449 9425
rect -24857 8180 -22323 8743
rect -27800 8000 -22323 8180
tri -22323 8000 -21580 8743 nw
tri -21474 8000 -20731 8743 se
rect -20731 8000 -15817 8743
tri -15817 8000 -15074 8743 nw
tri 10474 8000 11217 8743 ne
rect 11217 8576 15449 8743
tri 15449 8576 16298 9425 sw
tri 16298 8576 17147 9425 ne
rect 17147 8576 21106 9425
rect 11217 8000 16298 8576
rect -31800 7151 -23172 8000
tri -23172 7151 -22323 8000 nw
tri -22323 7151 -21474 8000 se
rect -21474 7151 -19200 8000
rect -31800 7123 -23200 7151
tri -23200 7123 -23172 7151 nw
tri -22351 7123 -22323 7151 se
rect -22323 7123 -19200 7151
rect -31800 4000 -23800 7123
tri -23800 6523 -23200 7123 nw
tri -22951 6523 -22351 7123 se
rect -22351 6523 -19200 7123
tri -23200 6274 -22951 6523 se
rect -22951 6274 -19200 6523
rect -28400 -4112 -24400 -4000
rect -28400 -7888 -28288 -4112
rect -24512 -7888 -24400 -4112
rect -28400 -8000 -24400 -7888
rect -23200 -8470 -19200 6274
tri -19200 4617 -15817 8000 nw
tri 11217 4617 14600 8000 ne
rect 14600 7972 16298 8000
tri 16298 7972 16902 8576 sw
tri 17147 7972 17751 8576 ne
rect 17751 8180 21106 8576
tri 21106 8180 23200 10274 sw
rect 17751 7972 23200 8180
rect 14600 7123 16902 7972
tri 16902 7123 17751 7972 sw
tri 17751 7123 18600 7972 ne
rect 18600 7123 23200 7972
rect 14600 6523 17751 7123
tri 17751 6523 18351 7123 sw
tri 18600 6523 19200 7123 ne
rect 14600 6274 18351 6523
tri 18351 6274 18600 6523 sw
rect -18600 -4112 -14600 -4000
tri -19200 -8470 -18600 -7870 sw
rect -18600 -7888 -18488 -4112
rect -14712 -7888 -14600 -4112
rect -18600 -8000 -14600 -7888
tri -18222 -8470 -17752 -8000 ne
rect -17752 -8470 -14600 -8000
rect -23200 -9318 -18600 -8470
tri -18600 -9318 -17752 -8470 sw
tri -17752 -9318 -16904 -8470 ne
rect -16904 -9318 -14600 -8470
rect -23200 -9527 -17752 -9318
tri -23200 -11622 -21105 -9527 ne
rect -21105 -9926 -17752 -9527
tri -17752 -9926 -17144 -9318 sw
tri -16904 -9926 -16296 -9318 ne
rect -16296 -9926 -14600 -9318
rect -21105 -10774 -17144 -9926
tri -17144 -10774 -16296 -9926 sw
tri -16296 -10774 -15448 -9926 ne
rect -15448 -10774 -14600 -9926
rect -21105 -11622 -16296 -10774
tri -16296 -11622 -15448 -10774 sw
tri -15448 -11622 -14600 -10774 ne
tri -14600 -11622 -8943 -5965 sw
tri 11822 -8743 14600 -5965 se
rect 14600 -7622 18600 6274
rect 14600 -7870 18352 -7622
tri 18352 -7870 18600 -7622 nw
rect 14600 -8470 17752 -7870
tri 17752 -8470 18352 -7870 nw
tri 18600 -8470 19200 -7870 se
rect 19200 -8470 23200 7123
rect 14600 -8743 17479 -8470
tri 17479 -8743 17752 -8470 nw
tri 18327 -8743 18600 -8470 se
rect 18600 -8743 23200 -8470
tri 8943 -11622 11822 -8743 se
rect 11822 -9591 16631 -8743
tri 16631 -9591 17479 -8743 nw
tri 17479 -9591 18327 -8743 se
rect 18327 -9527 23200 -8743
rect 18327 -9591 20257 -9527
rect 11822 -9926 16296 -9591
tri 16296 -9926 16631 -9591 nw
tri 17144 -9926 17479 -9591 se
rect 17479 -9926 20257 -9591
rect 11822 -10774 15448 -9926
tri 15448 -10774 16296 -9926 nw
tri 16296 -10774 17144 -9926 se
rect 17144 -10774 20257 -9926
rect 11822 -11622 14600 -10774
tri 14600 -11622 15448 -10774 nw
tri 15448 -11622 16296 -10774 se
rect 16296 -11622 20257 -10774
tri -21105 -14400 -18327 -11622 ne
rect -18327 -12470 -15448 -11622
tri -15448 -12470 -14600 -11622 sw
tri -14600 -12470 -13752 -11622 ne
rect -13752 -12470 -8943 -11622
rect -18327 -13318 -14600 -12470
tri -14600 -13318 -13752 -12470 sw
tri -13752 -13318 -12904 -12470 ne
rect -12904 -13318 -8943 -12470
rect -18327 -13552 -13752 -13318
tri -13752 -13552 -13518 -13318 sw
tri -12904 -13552 -12670 -13318 ne
rect -12670 -13552 -8943 -13318
rect -18327 -14400 -13518 -13552
tri -13518 -14400 -12670 -13552 sw
tri -12670 -14400 -11822 -13552 ne
rect -11822 -14400 -8943 -13552
tri -8943 -14400 -6165 -11622 sw
tri 6165 -14400 8943 -11622 se
rect 8943 -12470 13752 -11622
tri 13752 -12470 14600 -11622 nw
tri 14600 -12470 15448 -11622 se
rect 15448 -12470 20257 -11622
tri 20257 -12470 23200 -9527 nw
rect 8943 -13318 12904 -12470
tri 12904 -13318 13752 -12470 nw
tri 13752 -13318 14600 -12470 se
rect 14600 -13318 19200 -12470
rect 8943 -13552 12670 -13318
tri 12670 -13552 12904 -13318 nw
tri 13518 -13552 13752 -13318 se
rect 13752 -13527 19200 -13318
tri 19200 -13527 20257 -12470 nw
rect 13752 -13552 17479 -13527
rect 8943 -14400 11822 -13552
tri 11822 -14400 12670 -13552 nw
tri 12670 -14400 13518 -13552 se
rect 13518 -14400 17479 -13552
tri -18327 -19000 -13727 -14400 ne
rect -13727 -15248 -12670 -14400
tri -12670 -15248 -11822 -14400 sw
tri -11822 -15248 -10974 -14400 ne
rect -10974 -15248 10974 -14400
tri 10974 -15248 11822 -14400 nw
tri 11822 -15248 12670 -14400 se
rect 12670 -15248 17479 -14400
tri 17479 -15248 19200 -13527 nw
rect -13727 -16096 -11822 -15248
tri -11822 -16096 -10974 -15248 sw
tri -10974 -16096 -10126 -15248 ne
rect -10126 -16096 10126 -15248
tri 10126 -16096 10974 -15248 nw
tri 10974 -16096 11822 -15248 se
rect 11822 -16096 14600 -15248
rect -13727 -16704 -10974 -16096
tri -10974 -16704 -10366 -16096 sw
tri -10126 -16704 -9518 -16096 ne
rect -9518 -16704 9518 -16096
tri 9518 -16704 10126 -16096 nw
tri 10366 -16704 10974 -16096 se
rect 10974 -16704 14600 -16096
rect -13727 -17552 -10366 -16704
tri -10366 -17552 -9518 -16704 sw
tri -9518 -17552 -8670 -16704 ne
rect -8670 -17552 8670 -16704
tri 8670 -17552 9518 -16704 nw
tri 9518 -17552 10366 -16704 se
rect 10366 -17552 14600 -16704
rect -13727 -18400 -9518 -17552
tri -9518 -18400 -8670 -17552 sw
tri -8670 -18400 -7822 -17552 ne
rect -7822 -18400 7822 -17552
tri 7822 -18400 8670 -17552 nw
tri 8670 -18400 9518 -17552 se
rect 9518 -18127 14600 -17552
tri 14600 -18127 17479 -15248 nw
rect 9518 -18400 13727 -18127
rect -13727 -19000 -8670 -18400
tri -8670 -19000 -8070 -18400 sw
tri 8070 -19000 8670 -18400 se
rect 8670 -19000 13727 -18400
tri 13727 -19000 14600 -18127 nw
tri -13727 -20905 -11822 -19000 ne
rect -11822 -20905 11822 -19000
tri 11822 -20905 13727 -19000 nw
tri -11822 -23000 -9727 -20905 ne
rect -9727 -23000 9727 -20905
tri 9727 -23000 11822 -20905 nw
<< end >>
