magic
tech sky130A
magscale 1 2
timestamp 1658894429
<< nwell >>
rect 486 0 1078 2438
<< pmos >>
rect 682 219 882 2219
<< pdiff >>
rect 624 2207 682 2219
rect 624 231 636 2207
rect 670 231 682 2207
rect 624 219 682 231
rect 882 2207 940 2219
rect 882 231 894 2207
rect 928 231 940 2207
rect 882 219 940 231
<< pdiffc >>
rect 636 231 670 2207
rect 894 231 928 2207
<< nsubdiff >>
rect 522 2368 618 2402
rect 946 2368 1042 2402
rect 522 2306 556 2368
rect 1008 2306 1042 2368
rect 522 70 556 132
rect 1008 70 1042 132
rect 522 36 618 70
rect 946 36 1042 70
<< nsubdiffcont >>
rect 618 2368 946 2402
rect 522 132 556 2306
rect 1008 132 1042 2306
rect 618 36 946 70
<< poly >>
rect 682 2300 882 2316
rect 682 2266 698 2300
rect 866 2266 882 2300
rect 682 2219 882 2266
rect 682 172 882 219
rect 682 138 698 172
rect 866 138 882 172
rect 682 122 882 138
<< polycont >>
rect 698 2266 866 2300
rect 698 138 866 172
<< locali >>
rect 522 2368 618 2402
rect 946 2368 1042 2402
rect 522 2306 556 2368
rect 1008 2306 1042 2368
rect 682 2266 698 2300
rect 866 2266 882 2300
rect 636 2207 670 2223
rect 636 215 670 231
rect 894 2207 928 2223
rect 894 215 928 231
rect 682 138 698 172
rect 866 138 882 172
rect 522 70 556 132
rect 1008 70 1042 132
rect 522 36 618 70
rect 946 36 1042 70
<< viali >>
rect 698 2266 866 2300
rect 636 231 670 2207
rect 894 231 928 2207
rect 698 138 866 172
<< metal1 >>
rect 686 2300 878 2306
rect 686 2266 698 2300
rect 866 2266 878 2300
rect 686 2260 878 2266
rect 630 2207 676 2219
rect 630 231 636 2207
rect 670 231 676 2207
rect 630 219 676 231
rect 888 2207 934 2219
rect 888 231 894 2207
rect 928 231 934 2207
rect 888 219 934 231
rect 686 172 878 178
rect 686 138 698 172
rect 866 138 878 172
rect 686 132 878 138
use sky130_fd_pr__pfet_01v8_1um_10um  sky130_fd_pr__pfet_01v8_1um_10um_0
timestamp 1658894378
transform 1 0 53 0 1 53
box -53 -53 539 2385
<< end >>
