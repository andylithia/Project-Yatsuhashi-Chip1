magic
tech sky130B
magscale 1 2
timestamp 1606063140
<< nwell >>
rect -338 -497 338 497
<< mvpmos >>
rect -80 -200 80 200
<< mvpdiff >>
rect -138 188 -80 200
rect -138 -188 -126 188
rect -92 -188 -80 188
rect -138 -200 -80 -188
rect 80 188 138 200
rect 80 -188 92 188
rect 126 -188 138 188
rect 80 -200 138 -188
<< mvpdiffc >>
rect -126 -188 -92 188
rect 92 -188 126 188
<< mvnsubdiff >>
rect -272 419 272 431
rect -272 385 -164 419
rect 164 385 272 419
rect -272 373 272 385
rect -272 323 -214 373
rect -272 -323 -260 323
rect -226 -323 -214 323
rect 214 323 272 373
rect -272 -373 -214 -323
rect 214 -323 226 323
rect 260 -323 272 323
rect 214 -373 272 -323
rect -272 -385 272 -373
rect -272 -419 -164 -385
rect 164 -419 272 -385
rect -272 -431 272 -419
<< mvnsubdiffcont >>
rect -164 385 164 419
rect -260 -323 -226 323
rect 226 -323 260 323
rect -164 -419 164 -385
<< poly >>
rect -80 281 80 297
rect -80 247 -64 281
rect 64 247 80 281
rect -80 200 80 247
rect -80 -247 80 -200
rect -80 -281 -64 -247
rect 64 -281 80 -247
rect -80 -297 80 -281
<< polycont >>
rect -64 247 64 281
rect -64 -281 64 -247
<< locali >>
rect -260 385 -181 419
rect 181 385 260 419
rect -260 323 -226 385
rect 226 323 260 385
rect -80 247 -64 281
rect 64 247 80 281
rect -126 188 -92 204
rect -126 -204 -92 -188
rect 92 188 126 204
rect 92 -204 126 -188
rect -80 -281 -64 -247
rect 64 -281 80 -247
rect -260 -385 -226 -323
rect 226 -385 260 -323
rect -260 -419 -164 -385
rect 164 -419 260 -385
<< viali >>
rect -181 385 -164 419
rect -164 385 164 419
rect 164 385 181 419
rect -64 247 64 281
rect -126 -188 -92 188
rect 92 -188 126 188
rect -64 -281 64 -247
<< metal1 >>
rect -193 419 193 425
rect -193 385 -181 419
rect 181 385 193 419
rect -193 379 193 385
rect -76 281 76 287
rect -76 247 -64 281
rect 64 247 76 281
rect -76 241 76 247
rect -132 188 -86 200
rect -132 -188 -126 188
rect -92 -188 -86 188
rect -132 -200 -86 -188
rect 86 188 132 200
rect 86 -188 92 188
rect 126 -188 132 188
rect 86 -200 132 -188
rect -76 -247 76 -241
rect -76 -281 -64 -247
rect 64 -281 76 -247
rect -76 -287 76 -281
<< properties >>
string FIXED_BBOX -243 -402 243 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.00 l 0.80 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 80 viagb 0 viagate 100 viadrn 100 viasrc 100
<< end >>
