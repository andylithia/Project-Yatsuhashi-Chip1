magic
tech sky130B
timestamp 1659320289
<< metal1 >>
rect -1200 7650 7700 7700
rect -1200 -1950 -1150 7650
rect -650 7100 7150 7150
rect -650 6900 -600 7100
rect -400 6950 -100 7100
rect -350 6900 -100 6950
rect -650 6850 -450 6900
rect -300 6850 -100 6900
rect -650 6800 -400 6850
rect -250 6800 -100 6850
rect -650 6750 -350 6800
rect -200 6750 -100 6800
rect -650 6700 -300 6750
rect -150 6700 -100 6750
rect -650 6650 -250 6700
rect -650 6600 -200 6650
rect -650 6400 -600 6600
rect 100 6450 400 7100
rect 150 6400 400 6450
rect -650 6350 50 6400
rect 200 6350 400 6400
rect -650 6300 100 6350
rect 250 6300 400 6350
rect -650 6250 150 6300
rect 300 6250 400 6300
rect -650 6200 200 6250
rect 350 6200 400 6250
rect -650 6150 250 6200
rect -650 6100 300 6150
rect -650 5900 -600 6100
rect 600 5950 900 7100
rect 650 5900 900 5950
rect -650 5850 550 5900
rect 700 5850 900 5900
rect -650 5800 600 5850
rect 750 5800 900 5850
rect -650 5750 650 5800
rect 800 5750 900 5800
rect -650 5700 700 5750
rect 850 5700 900 5750
rect -650 5650 750 5700
rect -650 5600 800 5650
rect -650 5400 -600 5600
rect 1100 5450 1400 7100
rect 1150 5400 1400 5450
rect -650 5350 1050 5400
rect 1200 5350 1400 5400
rect -650 5300 1100 5350
rect 1250 5300 1400 5350
rect -650 5250 1150 5300
rect 1300 5250 1400 5300
rect -650 5200 1200 5250
rect 1350 5200 1400 5250
rect -650 5150 1250 5200
rect -650 5100 1300 5150
rect -650 4900 -600 5100
rect 1600 4950 1900 7100
rect 1650 4900 1900 4950
rect -650 4850 1550 4900
rect 1700 4850 1900 4900
rect -650 4800 1600 4850
rect 1750 4800 1900 4850
rect -650 4750 1650 4800
rect 1800 4750 1900 4800
rect -650 4700 1700 4750
rect 1850 4700 1900 4750
rect -650 4650 1750 4700
rect -650 4600 1800 4650
rect -650 4400 -600 4600
rect 2100 4450 2400 7100
rect 2150 4400 2400 4450
rect -650 4350 2050 4400
rect 2200 4350 2400 4400
rect -650 4300 2100 4350
rect 2250 4300 2400 4350
rect -650 4250 2150 4300
rect 2300 4250 2400 4300
rect -650 4200 2200 4250
rect 2350 4200 2400 4250
rect -650 4150 2250 4200
rect -650 4100 2300 4150
rect -650 3900 -600 4100
rect 2600 3950 2900 7100
rect 2650 3900 2900 3950
rect -650 3850 2550 3900
rect 2700 3850 2900 3900
rect -650 3800 2600 3850
rect 2750 3800 2900 3850
rect -650 3750 2650 3800
rect 2800 3750 2900 3800
rect -650 3700 2700 3750
rect 2850 3700 2900 3750
rect 3100 3700 3400 7100
rect 3600 3950 3900 7100
rect 4100 4450 4400 7100
rect 4600 4950 4900 7100
rect 5100 5450 5400 7100
rect 5600 5950 5900 7100
rect 6100 6450 6400 7100
rect 6600 6950 6900 7100
rect 6600 6900 6850 6950
rect 7100 6900 7150 7100
rect 6600 6850 6800 6900
rect 6950 6850 7150 6900
rect 6600 6800 6750 6850
rect 6900 6800 7150 6850
rect 6600 6750 6700 6800
rect 6850 6750 7150 6800
rect 6600 6700 6650 6750
rect 6800 6700 7150 6750
rect 6750 6650 7150 6700
rect 6700 6600 7150 6650
rect 6100 6400 6350 6450
rect 7100 6400 7150 6600
rect 6100 6350 6300 6400
rect 6450 6350 7150 6400
rect 6100 6300 6250 6350
rect 6400 6300 7150 6350
rect 6100 6250 6200 6300
rect 6350 6250 7150 6300
rect 6100 6200 6150 6250
rect 6300 6200 7150 6250
rect 6250 6150 7150 6200
rect 6200 6100 7150 6150
rect 5600 5900 5850 5950
rect 7100 5900 7150 6100
rect 5600 5850 5800 5900
rect 5950 5850 7150 5900
rect 5600 5800 5750 5850
rect 5900 5800 7150 5850
rect 5600 5750 5700 5800
rect 5850 5750 7150 5800
rect 5600 5700 5650 5750
rect 5800 5700 7150 5750
rect 5750 5650 7150 5700
rect 5700 5600 7150 5650
rect 5100 5400 5350 5450
rect 7100 5400 7150 5600
rect 5100 5350 5300 5400
rect 5450 5350 7150 5400
rect 5100 5300 5250 5350
rect 5400 5300 7150 5350
rect 5100 5250 5200 5300
rect 5350 5250 7150 5300
rect 5100 5200 5150 5250
rect 5300 5200 7150 5250
rect 5250 5150 7150 5200
rect 5200 5100 7150 5150
rect 4600 4900 4850 4950
rect 7100 4900 7150 5100
rect 4600 4850 4800 4900
rect 4950 4850 7150 4900
rect 4600 4800 4750 4850
rect 4900 4800 7150 4850
rect 4600 4750 4700 4800
rect 4850 4750 7150 4800
rect 4600 4700 4650 4750
rect 4800 4700 7150 4750
rect 4750 4650 7150 4700
rect 4700 4600 7150 4650
rect 4100 4400 4350 4450
rect 7100 4400 7150 4600
rect 4100 4350 4300 4400
rect 4450 4350 7150 4400
rect 4100 4300 4250 4350
rect 4400 4300 7150 4350
rect 4100 4250 4200 4300
rect 4350 4250 7150 4300
rect 4100 4200 4150 4250
rect 4300 4200 7150 4250
rect 4250 4150 7150 4200
rect 4200 4100 7150 4150
rect 3600 3900 3850 3950
rect 7100 3900 7150 4100
rect 3600 3850 3800 3900
rect 3950 3850 7150 3900
rect 3600 3800 3750 3850
rect 3900 3800 7150 3850
rect 3600 3750 3700 3800
rect 3850 3750 7150 3800
rect 3600 3700 3650 3750
rect 3800 3700 7150 3750
rect -650 3650 2750 3700
rect 3750 3650 7150 3700
rect -650 3600 2800 3650
rect 3700 3600 7150 3650
rect -650 3400 -600 3600
rect 7100 3400 7150 3600
rect -650 3100 2800 3400
rect 3700 3100 7150 3400
rect -650 2900 -600 3100
rect 7100 2900 7150 3100
rect -650 2850 2800 2900
rect 3700 2850 7150 2900
rect -650 2800 2750 2850
rect 3750 2800 7150 2850
rect -650 2750 2700 2800
rect 2850 2750 2900 2800
rect -650 2700 2650 2750
rect 2800 2700 2900 2750
rect -650 2650 2600 2700
rect 2750 2650 2900 2700
rect -650 2600 2550 2650
rect 2700 2600 2900 2650
rect -650 2400 -600 2600
rect 2650 2550 2900 2600
rect -650 2350 2300 2400
rect -650 2300 2250 2350
rect -650 2250 2200 2300
rect 2350 2250 2400 2300
rect -650 2200 2150 2250
rect 2300 2200 2400 2250
rect -650 2150 2100 2200
rect 2250 2150 2400 2200
rect -650 2100 2050 2150
rect 2200 2100 2400 2150
rect -650 1900 -600 2100
rect 2150 2050 2400 2100
rect -650 1850 1800 1900
rect -650 1800 1750 1850
rect -650 1750 1700 1800
rect 1850 1750 1900 1800
rect -650 1700 1650 1750
rect 1800 1700 1900 1750
rect -650 1650 1600 1700
rect 1750 1650 1900 1700
rect -650 1600 1550 1650
rect 1700 1600 1900 1650
rect -650 1400 -600 1600
rect 1650 1550 1900 1600
rect -650 1350 1300 1400
rect -650 1300 1250 1350
rect -650 1250 1200 1300
rect 1350 1250 1400 1300
rect -650 1200 1150 1250
rect 1300 1200 1400 1250
rect -650 1150 1100 1200
rect 1250 1150 1400 1200
rect -650 1100 1050 1150
rect 1200 1100 1400 1150
rect -650 900 -600 1100
rect 1150 1050 1400 1100
rect -650 850 800 900
rect -650 800 750 850
rect -650 750 700 800
rect 850 750 900 800
rect -650 700 650 750
rect 800 700 900 750
rect -650 650 600 700
rect 750 650 900 700
rect -650 600 550 650
rect 700 600 900 650
rect -650 400 -600 600
rect 650 550 900 600
rect -650 350 300 400
rect -650 300 250 350
rect -650 250 200 300
rect 350 250 400 300
rect -650 200 150 250
rect 300 200 400 250
rect -650 150 100 200
rect 250 150 400 200
rect -650 100 50 150
rect 200 100 400 150
rect -650 -100 -600 100
rect 150 50 400 100
rect -650 -150 -200 -100
rect -650 -200 -250 -150
rect -650 -250 -300 -200
rect -150 -250 -100 -200
rect -650 -300 -350 -250
rect -200 -300 -100 -250
rect -650 -350 -400 -300
rect -250 -350 -100 -300
rect -650 -400 -450 -350
rect -300 -400 -100 -350
rect -650 -1400 -600 -400
rect -350 -450 -100 -400
rect -400 -1400 -100 -450
rect 100 -1400 400 50
rect 600 -1400 900 550
rect 1100 -1400 1400 1050
rect 1600 -1400 1900 1550
rect 2100 -1400 2400 2050
rect 2600 -1400 2900 2550
rect 3100 -1400 3400 2800
rect 3600 2750 3650 2800
rect 3800 2750 7150 2800
rect 3600 2700 3700 2750
rect 3850 2700 7150 2750
rect 3600 2650 3750 2700
rect 3900 2650 7150 2700
rect 3600 2600 3800 2650
rect 3950 2600 7150 2650
rect 3600 2550 3850 2600
rect 3600 -1400 3900 2550
rect 7100 2400 7150 2600
rect 4200 2350 7150 2400
rect 4250 2300 7150 2350
rect 4100 2250 4150 2300
rect 4300 2250 7150 2300
rect 4100 2200 4200 2250
rect 4350 2200 7150 2250
rect 4100 2150 4250 2200
rect 4400 2150 7150 2200
rect 4100 2100 4300 2150
rect 4450 2100 7150 2150
rect 4100 2050 4350 2100
rect 4100 -1400 4400 2050
rect 7100 1900 7150 2100
rect 4700 1850 7150 1900
rect 4750 1800 7150 1850
rect 4600 1750 4650 1800
rect 4800 1750 7150 1800
rect 4600 1700 4700 1750
rect 4850 1700 7150 1750
rect 4600 1650 4750 1700
rect 4900 1650 7150 1700
rect 4600 1600 4800 1650
rect 4950 1600 7150 1650
rect 4600 1550 4850 1600
rect 4600 -1400 4900 1550
rect 7100 1400 7150 1600
rect 5200 1350 7150 1400
rect 5250 1300 7150 1350
rect 5100 1250 5150 1300
rect 5300 1250 7150 1300
rect 5100 1200 5200 1250
rect 5350 1200 7150 1250
rect 5100 1150 5250 1200
rect 5400 1150 7150 1200
rect 5100 1100 5300 1150
rect 5450 1100 7150 1150
rect 5100 1050 5350 1100
rect 5100 -1400 5400 1050
rect 7100 900 7150 1100
rect 5700 850 7150 900
rect 5750 800 7150 850
rect 5600 750 5650 800
rect 5800 750 7150 800
rect 5600 700 5700 750
rect 5850 700 7150 750
rect 5600 650 5750 700
rect 5900 650 7150 700
rect 5600 600 5800 650
rect 5950 600 7150 650
rect 5600 550 5850 600
rect 5600 -1400 5900 550
rect 7100 400 7150 600
rect 6200 350 7150 400
rect 6250 300 7150 350
rect 6100 250 6150 300
rect 6300 250 7150 300
rect 6100 200 6200 250
rect 6350 200 7150 250
rect 6100 150 6250 200
rect 6400 150 7150 200
rect 6100 100 6300 150
rect 6450 100 7150 150
rect 6100 50 6350 100
rect 6100 -1400 6400 50
rect 7100 -100 7150 100
rect 6700 -150 7150 -100
rect 6750 -200 7150 -150
rect 6600 -250 6650 -200
rect 6800 -250 7150 -200
rect 6600 -300 6700 -250
rect 6850 -300 7150 -250
rect 6600 -350 6750 -300
rect 6900 -350 7150 -300
rect 6600 -400 6800 -350
rect 6950 -400 7150 -350
rect 6600 -450 6850 -400
rect 6600 -1400 6900 -450
rect 7100 -1400 7150 -400
rect -650 -1450 7150 -1400
rect 7650 -1950 7700 7650
rect -1200 -2000 7700 -1950
<< via1 >>
rect -1150 7150 7650 7650
rect -1150 -1450 -650 7150
rect 7150 -1450 7650 7150
rect -1150 -1950 7650 -1450
<< metal2 >>
rect -1200 7650 7700 7700
rect -1200 -1950 -1150 7650
rect -650 7100 7150 7150
rect -650 6900 -600 7100
rect -400 6950 -100 7100
rect -350 6900 -100 6950
rect -650 6850 -450 6900
rect -300 6850 -100 6900
rect -650 6800 -400 6850
rect -250 6800 -100 6850
rect -650 6750 -350 6800
rect -200 6750 -100 6800
rect -650 6700 -300 6750
rect -150 6700 -100 6750
rect -650 6650 -250 6700
rect -650 6600 -200 6650
rect -650 6400 -600 6600
rect 100 6450 400 7100
rect 150 6400 400 6450
rect -650 6350 50 6400
rect 200 6350 400 6400
rect -650 6300 100 6350
rect 250 6300 400 6350
rect -650 6250 150 6300
rect 300 6250 400 6300
rect -650 6200 200 6250
rect 350 6200 400 6250
rect -650 6150 250 6200
rect -650 6100 300 6150
rect -650 5900 -600 6100
rect 600 5950 900 7100
rect 650 5900 900 5950
rect -650 5850 550 5900
rect 700 5850 900 5900
rect -650 5800 600 5850
rect 750 5800 900 5850
rect -650 5750 650 5800
rect 800 5750 900 5800
rect -650 5700 700 5750
rect 850 5700 900 5750
rect -650 5650 750 5700
rect -650 5600 800 5650
rect -650 5400 -600 5600
rect 1100 5450 1400 7100
rect 1150 5400 1400 5450
rect -650 5350 1050 5400
rect 1200 5350 1400 5400
rect -650 5300 1100 5350
rect 1250 5300 1400 5350
rect -650 5250 1150 5300
rect 1300 5250 1400 5300
rect -650 5200 1200 5250
rect 1350 5200 1400 5250
rect -650 5150 1250 5200
rect -650 5100 1300 5150
rect -650 4900 -600 5100
rect 1600 4950 1900 7100
rect 1650 4900 1900 4950
rect -650 4850 1550 4900
rect 1700 4850 1900 4900
rect -650 4800 1600 4850
rect 1750 4800 1900 4850
rect -650 4750 1650 4800
rect 1800 4750 1900 4800
rect -650 4700 1700 4750
rect 1850 4700 1900 4750
rect -650 4650 1750 4700
rect -650 4600 1800 4650
rect -650 4400 -600 4600
rect 2100 4450 2400 7100
rect 2150 4400 2400 4450
rect -650 4350 2050 4400
rect 2200 4350 2400 4400
rect -650 4300 2100 4350
rect 2250 4300 2400 4350
rect -650 4250 2150 4300
rect 2300 4250 2400 4300
rect -650 4200 2200 4250
rect 2350 4200 2400 4250
rect -650 4150 2250 4200
rect -650 4100 2300 4150
rect -650 3900 -600 4100
rect 2600 3950 2900 7100
rect 2650 3900 2900 3950
rect -650 3850 2550 3900
rect 2700 3850 2900 3900
rect -650 3800 2600 3850
rect 2750 3800 2900 3850
rect -650 3750 2650 3800
rect 2800 3750 2900 3800
rect -650 3700 2700 3750
rect 2850 3700 2900 3750
rect 3100 3700 3400 7100
rect 3600 3950 3900 7100
rect 4100 4450 4400 7100
rect 4600 4950 4900 7100
rect 5100 5450 5400 7100
rect 5600 5950 5900 7100
rect 6100 6450 6400 7100
rect 6600 6950 6900 7100
rect 6600 6900 6850 6950
rect 7100 6900 7150 7100
rect 6600 6850 6800 6900
rect 6950 6850 7150 6900
rect 6600 6800 6750 6850
rect 6900 6800 7150 6850
rect 6600 6750 6700 6800
rect 6850 6750 7150 6800
rect 6600 6700 6650 6750
rect 6800 6700 7150 6750
rect 6750 6650 7150 6700
rect 6700 6600 7150 6650
rect 6100 6400 6350 6450
rect 7100 6400 7150 6600
rect 6100 6350 6300 6400
rect 6450 6350 7150 6400
rect 6100 6300 6250 6350
rect 6400 6300 7150 6350
rect 6100 6250 6200 6300
rect 6350 6250 7150 6300
rect 6100 6200 6150 6250
rect 6300 6200 7150 6250
rect 6250 6150 7150 6200
rect 6200 6100 7150 6150
rect 5600 5900 5850 5950
rect 7100 5900 7150 6100
rect 5600 5850 5800 5900
rect 5950 5850 7150 5900
rect 5600 5800 5750 5850
rect 5900 5800 7150 5850
rect 5600 5750 5700 5800
rect 5850 5750 7150 5800
rect 5600 5700 5650 5750
rect 5800 5700 7150 5750
rect 5750 5650 7150 5700
rect 5700 5600 7150 5650
rect 5100 5400 5350 5450
rect 7100 5400 7150 5600
rect 5100 5350 5300 5400
rect 5450 5350 7150 5400
rect 5100 5300 5250 5350
rect 5400 5300 7150 5350
rect 5100 5250 5200 5300
rect 5350 5250 7150 5300
rect 5100 5200 5150 5250
rect 5300 5200 7150 5250
rect 5250 5150 7150 5200
rect 5200 5100 7150 5150
rect 4600 4900 4850 4950
rect 7100 4900 7150 5100
rect 4600 4850 4800 4900
rect 4950 4850 7150 4900
rect 4600 4800 4750 4850
rect 4900 4800 7150 4850
rect 4600 4750 4700 4800
rect 4850 4750 7150 4800
rect 4600 4700 4650 4750
rect 4800 4700 7150 4750
rect 4750 4650 7150 4700
rect 4700 4600 7150 4650
rect 4100 4400 4350 4450
rect 7100 4400 7150 4600
rect 4100 4350 4300 4400
rect 4450 4350 7150 4400
rect 4100 4300 4250 4350
rect 4400 4300 7150 4350
rect 4100 4250 4200 4300
rect 4350 4250 7150 4300
rect 4100 4200 4150 4250
rect 4300 4200 7150 4250
rect 4250 4150 7150 4200
rect 4200 4100 7150 4150
rect 3600 3900 3850 3950
rect 7100 3900 7150 4100
rect 3600 3850 3800 3900
rect 3950 3850 7150 3900
rect 3600 3800 3750 3850
rect 3900 3800 7150 3850
rect 3600 3750 3700 3800
rect 3850 3750 7150 3800
rect 3600 3700 3650 3750
rect 3800 3700 7150 3750
rect -650 3650 2750 3700
rect 3750 3650 7150 3700
rect -650 3600 2800 3650
rect 3700 3600 7150 3650
rect -650 3400 -600 3600
rect 7100 3400 7150 3600
rect -650 3100 2800 3400
rect 3700 3100 7150 3400
rect -650 2900 -600 3100
rect 7100 2900 7150 3100
rect -650 2850 2800 2900
rect 3700 2850 7150 2900
rect -650 2800 2750 2850
rect 3750 2800 7150 2850
rect -650 2750 2700 2800
rect 2850 2750 2900 2800
rect -650 2700 2650 2750
rect 2800 2700 2900 2750
rect -650 2650 2600 2700
rect 2750 2650 2900 2700
rect -650 2600 2550 2650
rect 2700 2600 2900 2650
rect -650 2400 -600 2600
rect 2650 2550 2900 2600
rect -650 2350 2300 2400
rect -650 2300 2250 2350
rect -650 2250 2200 2300
rect 2350 2250 2400 2300
rect -650 2200 2150 2250
rect 2300 2200 2400 2250
rect -650 2150 2100 2200
rect 2250 2150 2400 2200
rect -650 2100 2050 2150
rect 2200 2100 2400 2150
rect -650 1900 -600 2100
rect 2150 2050 2400 2100
rect -650 1850 1800 1900
rect -650 1800 1750 1850
rect -650 1750 1700 1800
rect 1850 1750 1900 1800
rect -650 1700 1650 1750
rect 1800 1700 1900 1750
rect -650 1650 1600 1700
rect 1750 1650 1900 1700
rect -650 1600 1550 1650
rect 1700 1600 1900 1650
rect -650 1400 -600 1600
rect 1650 1550 1900 1600
rect -650 1350 1300 1400
rect -650 1300 1250 1350
rect -650 1250 1200 1300
rect 1350 1250 1400 1300
rect -650 1200 1150 1250
rect 1300 1200 1400 1250
rect -650 1150 1100 1200
rect 1250 1150 1400 1200
rect -650 1100 1050 1150
rect 1200 1100 1400 1150
rect -650 900 -600 1100
rect 1150 1050 1400 1100
rect -650 850 800 900
rect -650 800 750 850
rect -650 750 700 800
rect 850 750 900 800
rect -650 700 650 750
rect 800 700 900 750
rect -650 650 600 700
rect 750 650 900 700
rect -650 600 550 650
rect 700 600 900 650
rect -650 400 -600 600
rect 650 550 900 600
rect -650 350 300 400
rect -650 300 250 350
rect -650 250 200 300
rect 350 250 400 300
rect -650 200 150 250
rect 300 200 400 250
rect -650 150 100 200
rect 250 150 400 200
rect -650 100 50 150
rect 200 100 400 150
rect -650 -100 -600 100
rect 150 50 400 100
rect -650 -150 -200 -100
rect -650 -200 -250 -150
rect -650 -250 -300 -200
rect -150 -250 -100 -200
rect -650 -300 -350 -250
rect -200 -300 -100 -250
rect -650 -350 -400 -300
rect -250 -350 -100 -300
rect -650 -400 -450 -350
rect -300 -400 -100 -350
rect -650 -1400 -600 -400
rect -350 -450 -100 -400
rect -400 -1400 -100 -450
rect 100 -1400 400 50
rect 600 -1400 900 550
rect 1100 -1400 1400 1050
rect 1600 -1400 1900 1550
rect 2100 -1400 2400 2050
rect 2600 -1400 2900 2550
rect 3100 -1400 3400 2800
rect 3600 2750 3650 2800
rect 3800 2750 7150 2800
rect 3600 2700 3700 2750
rect 3850 2700 7150 2750
rect 3600 2650 3750 2700
rect 3900 2650 7150 2700
rect 3600 2600 3800 2650
rect 3950 2600 7150 2650
rect 3600 2550 3850 2600
rect 3600 -1400 3900 2550
rect 7100 2400 7150 2600
rect 4200 2350 7150 2400
rect 4250 2300 7150 2350
rect 4100 2250 4150 2300
rect 4300 2250 7150 2300
rect 4100 2200 4200 2250
rect 4350 2200 7150 2250
rect 4100 2150 4250 2200
rect 4400 2150 7150 2200
rect 4100 2100 4300 2150
rect 4450 2100 7150 2150
rect 4100 2050 4350 2100
rect 4100 -1400 4400 2050
rect 7100 1900 7150 2100
rect 4700 1850 7150 1900
rect 4750 1800 7150 1850
rect 4600 1750 4650 1800
rect 4800 1750 7150 1800
rect 4600 1700 4700 1750
rect 4850 1700 7150 1750
rect 4600 1650 4750 1700
rect 4900 1650 7150 1700
rect 4600 1600 4800 1650
rect 4950 1600 7150 1650
rect 4600 1550 4850 1600
rect 4600 -1400 4900 1550
rect 7100 1400 7150 1600
rect 5200 1350 7150 1400
rect 5250 1300 7150 1350
rect 5100 1250 5150 1300
rect 5300 1250 7150 1300
rect 5100 1200 5200 1250
rect 5350 1200 7150 1250
rect 5100 1150 5250 1200
rect 5400 1150 7150 1200
rect 5100 1100 5300 1150
rect 5450 1100 7150 1150
rect 5100 1050 5350 1100
rect 5100 -1400 5400 1050
rect 7100 900 7150 1100
rect 5700 850 7150 900
rect 5750 800 7150 850
rect 5600 750 5650 800
rect 5800 750 7150 800
rect 5600 700 5700 750
rect 5850 700 7150 750
rect 5600 650 5750 700
rect 5900 650 7150 700
rect 5600 600 5800 650
rect 5950 600 7150 650
rect 5600 550 5850 600
rect 5600 -1400 5900 550
rect 7100 400 7150 600
rect 6200 350 7150 400
rect 6250 300 7150 350
rect 6100 250 6150 300
rect 6300 250 7150 300
rect 6100 200 6200 250
rect 6350 200 7150 250
rect 6100 150 6250 200
rect 6400 150 7150 200
rect 6100 100 6300 150
rect 6450 100 7150 150
rect 6100 50 6350 100
rect 6100 -1400 6400 50
rect 7100 -100 7150 100
rect 6700 -150 7150 -100
rect 6750 -200 7150 -150
rect 6600 -250 6650 -200
rect 6800 -250 7150 -200
rect 6600 -300 6700 -250
rect 6850 -300 7150 -250
rect 6600 -350 6750 -300
rect 6900 -350 7150 -300
rect 6600 -400 6800 -350
rect 6950 -400 7150 -350
rect 6600 -450 6850 -400
rect 6600 -1400 6900 -450
rect 7100 -1400 7150 -400
rect -650 -1450 7150 -1400
rect 7650 -1950 7700 7650
rect -1200 -2000 7700 -1950
<< via2 >>
rect -1150 7150 7650 7650
rect -1150 -1450 -650 7150
rect 7150 -1450 7650 7150
rect -1150 -1950 7650 -1450
<< metal3 >>
rect -1200 7650 7700 7700
rect -1200 -1950 -1150 7650
rect -650 7100 7150 7150
rect -650 6900 -600 7100
rect -400 6950 -100 7100
rect -350 6900 -100 6950
rect -650 6850 -450 6900
rect -300 6850 -100 6900
rect -650 6800 -400 6850
rect -250 6800 -100 6850
rect -650 6750 -350 6800
rect -200 6750 -100 6800
rect -650 6700 -300 6750
rect -150 6700 -100 6750
rect -650 6650 -250 6700
rect -650 6600 -200 6650
rect -650 6400 -600 6600
rect 100 6450 400 7100
rect 150 6400 400 6450
rect -650 6350 50 6400
rect 200 6350 400 6400
rect -650 6300 100 6350
rect 250 6300 400 6350
rect -650 6250 150 6300
rect 300 6250 400 6300
rect -650 6200 200 6250
rect 350 6200 400 6250
rect -650 6150 250 6200
rect -650 6100 300 6150
rect -650 5900 -600 6100
rect 600 5950 900 7100
rect 650 5900 900 5950
rect -650 5850 550 5900
rect 700 5850 900 5900
rect -650 5800 600 5850
rect 750 5800 900 5850
rect -650 5750 650 5800
rect 800 5750 900 5800
rect -650 5700 700 5750
rect 850 5700 900 5750
rect -650 5650 750 5700
rect -650 5600 800 5650
rect -650 5400 -600 5600
rect 1100 5450 1400 7100
rect 1150 5400 1400 5450
rect -650 5350 1050 5400
rect 1200 5350 1400 5400
rect -650 5300 1100 5350
rect 1250 5300 1400 5350
rect -650 5250 1150 5300
rect 1300 5250 1400 5300
rect -650 5200 1200 5250
rect 1350 5200 1400 5250
rect -650 5150 1250 5200
rect -650 5100 1300 5150
rect -650 4900 -600 5100
rect 1600 4950 1900 7100
rect 1650 4900 1900 4950
rect -650 4850 1550 4900
rect 1700 4850 1900 4900
rect -650 4800 1600 4850
rect 1750 4800 1900 4850
rect -650 4750 1650 4800
rect 1800 4750 1900 4800
rect -650 4700 1700 4750
rect 1850 4700 1900 4750
rect -650 4650 1750 4700
rect -650 4600 1800 4650
rect -650 4400 -600 4600
rect 2100 4450 2400 7100
rect 2150 4400 2400 4450
rect -650 4350 2050 4400
rect 2200 4350 2400 4400
rect -650 4300 2100 4350
rect 2250 4300 2400 4350
rect -650 4250 2150 4300
rect 2300 4250 2400 4300
rect -650 4200 2200 4250
rect 2350 4200 2400 4250
rect -650 4150 2250 4200
rect -650 4100 2300 4150
rect -650 3900 -600 4100
rect 2600 3950 2900 7100
rect 2650 3900 2900 3950
rect -650 3850 2550 3900
rect 2700 3850 2900 3900
rect -650 3800 2600 3850
rect 2750 3800 2900 3850
rect -650 3750 2650 3800
rect 2800 3750 2900 3800
rect -650 3700 2700 3750
rect 2850 3700 2900 3750
rect 3100 3700 3400 7100
rect 3600 3950 3900 7100
rect 4100 4450 4400 7100
rect 4600 4950 4900 7100
rect 5100 5450 5400 7100
rect 5600 5950 5900 7100
rect 6100 6450 6400 7100
rect 6600 6950 6900 7100
rect 6600 6900 6850 6950
rect 7100 6900 7150 7100
rect 6600 6850 6800 6900
rect 6950 6850 7150 6900
rect 6600 6800 6750 6850
rect 6900 6800 7150 6850
rect 6600 6750 6700 6800
rect 6850 6750 7150 6800
rect 6600 6700 6650 6750
rect 6800 6700 7150 6750
rect 6750 6650 7150 6700
rect 6700 6600 7150 6650
rect 6100 6400 6350 6450
rect 7100 6400 7150 6600
rect 6100 6350 6300 6400
rect 6450 6350 7150 6400
rect 6100 6300 6250 6350
rect 6400 6300 7150 6350
rect 6100 6250 6200 6300
rect 6350 6250 7150 6300
rect 6100 6200 6150 6250
rect 6300 6200 7150 6250
rect 6250 6150 7150 6200
rect 6200 6100 7150 6150
rect 5600 5900 5850 5950
rect 7100 5900 7150 6100
rect 5600 5850 5800 5900
rect 5950 5850 7150 5900
rect 5600 5800 5750 5850
rect 5900 5800 7150 5850
rect 5600 5750 5700 5800
rect 5850 5750 7150 5800
rect 5600 5700 5650 5750
rect 5800 5700 7150 5750
rect 5750 5650 7150 5700
rect 5700 5600 7150 5650
rect 5100 5400 5350 5450
rect 7100 5400 7150 5600
rect 5100 5350 5300 5400
rect 5450 5350 7150 5400
rect 5100 5300 5250 5350
rect 5400 5300 7150 5350
rect 5100 5250 5200 5300
rect 5350 5250 7150 5300
rect 5100 5200 5150 5250
rect 5300 5200 7150 5250
rect 5250 5150 7150 5200
rect 5200 5100 7150 5150
rect 4600 4900 4850 4950
rect 7100 4900 7150 5100
rect 4600 4850 4800 4900
rect 4950 4850 7150 4900
rect 4600 4800 4750 4850
rect 4900 4800 7150 4850
rect 4600 4750 4700 4800
rect 4850 4750 7150 4800
rect 4600 4700 4650 4750
rect 4800 4700 7150 4750
rect 4750 4650 7150 4700
rect 4700 4600 7150 4650
rect 4100 4400 4350 4450
rect 7100 4400 7150 4600
rect 4100 4350 4300 4400
rect 4450 4350 7150 4400
rect 4100 4300 4250 4350
rect 4400 4300 7150 4350
rect 4100 4250 4200 4300
rect 4350 4250 7150 4300
rect 4100 4200 4150 4250
rect 4300 4200 7150 4250
rect 4250 4150 7150 4200
rect 4200 4100 7150 4150
rect 3600 3900 3850 3950
rect 7100 3900 7150 4100
rect 3600 3850 3800 3900
rect 3950 3850 7150 3900
rect 3600 3800 3750 3850
rect 3900 3800 7150 3850
rect 3600 3750 3700 3800
rect 3850 3750 7150 3800
rect 3600 3700 3650 3750
rect 3800 3700 7150 3750
rect -650 3650 2750 3700
rect 3750 3650 7150 3700
rect -650 3600 2800 3650
rect 3700 3600 7150 3650
rect -650 3400 -600 3600
rect 7100 3400 7150 3600
rect -650 3100 2800 3400
rect 3700 3100 7150 3400
rect -650 2900 -600 3100
rect 7100 2900 7150 3100
rect -650 2850 2800 2900
rect 3700 2850 7150 2900
rect -650 2800 2750 2850
rect 3750 2800 7150 2850
rect -650 2750 2700 2800
rect 2850 2750 2900 2800
rect -650 2700 2650 2750
rect 2800 2700 2900 2750
rect -650 2650 2600 2700
rect 2750 2650 2900 2700
rect -650 2600 2550 2650
rect 2700 2600 2900 2650
rect -650 2400 -600 2600
rect 2650 2550 2900 2600
rect -650 2350 2300 2400
rect -650 2300 2250 2350
rect -650 2250 2200 2300
rect 2350 2250 2400 2300
rect -650 2200 2150 2250
rect 2300 2200 2400 2250
rect -650 2150 2100 2200
rect 2250 2150 2400 2200
rect -650 2100 2050 2150
rect 2200 2100 2400 2150
rect -650 1900 -600 2100
rect 2150 2050 2400 2100
rect -650 1850 1800 1900
rect -650 1800 1750 1850
rect -650 1750 1700 1800
rect 1850 1750 1900 1800
rect -650 1700 1650 1750
rect 1800 1700 1900 1750
rect -650 1650 1600 1700
rect 1750 1650 1900 1700
rect -650 1600 1550 1650
rect 1700 1600 1900 1650
rect -650 1400 -600 1600
rect 1650 1550 1900 1600
rect -650 1350 1300 1400
rect -650 1300 1250 1350
rect -650 1250 1200 1300
rect 1350 1250 1400 1300
rect -650 1200 1150 1250
rect 1300 1200 1400 1250
rect -650 1150 1100 1200
rect 1250 1150 1400 1200
rect -650 1100 1050 1150
rect 1200 1100 1400 1150
rect -650 900 -600 1100
rect 1150 1050 1400 1100
rect -650 850 800 900
rect -650 800 750 850
rect -650 750 700 800
rect 850 750 900 800
rect -650 700 650 750
rect 800 700 900 750
rect -650 650 600 700
rect 750 650 900 700
rect -650 600 550 650
rect 700 600 900 650
rect -650 400 -600 600
rect 650 550 900 600
rect -650 350 300 400
rect -650 300 250 350
rect -650 250 200 300
rect 350 250 400 300
rect -650 200 150 250
rect 300 200 400 250
rect -650 150 100 200
rect 250 150 400 200
rect -650 100 50 150
rect 200 100 400 150
rect -650 -100 -600 100
rect 150 50 400 100
rect -650 -150 -200 -100
rect -650 -200 -250 -150
rect -650 -250 -300 -200
rect -150 -250 -100 -200
rect -650 -300 -350 -250
rect -200 -300 -100 -250
rect -650 -350 -400 -300
rect -250 -350 -100 -300
rect -650 -400 -450 -350
rect -300 -400 -100 -350
rect -650 -1400 -600 -400
rect -350 -450 -100 -400
rect -400 -1400 -100 -450
rect 100 -1400 400 50
rect 600 -1400 900 550
rect 1100 -1400 1400 1050
rect 1600 -1400 1900 1550
rect 2100 -1400 2400 2050
rect 2600 -1400 2900 2550
rect 3100 -1400 3400 2800
rect 3600 2750 3650 2800
rect 3800 2750 7150 2800
rect 3600 2700 3700 2750
rect 3850 2700 7150 2750
rect 3600 2650 3750 2700
rect 3900 2650 7150 2700
rect 3600 2600 3800 2650
rect 3950 2600 7150 2650
rect 3600 2550 3850 2600
rect 3600 -1400 3900 2550
rect 7100 2400 7150 2600
rect 4200 2350 7150 2400
rect 4250 2300 7150 2350
rect 4100 2250 4150 2300
rect 4300 2250 7150 2300
rect 4100 2200 4200 2250
rect 4350 2200 7150 2250
rect 4100 2150 4250 2200
rect 4400 2150 7150 2200
rect 4100 2100 4300 2150
rect 4450 2100 7150 2150
rect 4100 2050 4350 2100
rect 4100 -1400 4400 2050
rect 7100 1900 7150 2100
rect 4700 1850 7150 1900
rect 4750 1800 7150 1850
rect 4600 1750 4650 1800
rect 4800 1750 7150 1800
rect 4600 1700 4700 1750
rect 4850 1700 7150 1750
rect 4600 1650 4750 1700
rect 4900 1650 7150 1700
rect 4600 1600 4800 1650
rect 4950 1600 7150 1650
rect 4600 1550 4850 1600
rect 4600 -1400 4900 1550
rect 7100 1400 7150 1600
rect 5200 1350 7150 1400
rect 5250 1300 7150 1350
rect 5100 1250 5150 1300
rect 5300 1250 7150 1300
rect 5100 1200 5200 1250
rect 5350 1200 7150 1250
rect 5100 1150 5250 1200
rect 5400 1150 7150 1200
rect 5100 1100 5300 1150
rect 5450 1100 7150 1150
rect 5100 1050 5350 1100
rect 5100 -1400 5400 1050
rect 7100 900 7150 1100
rect 5700 850 7150 900
rect 5750 800 7150 850
rect 5600 750 5650 800
rect 5800 750 7150 800
rect 5600 700 5700 750
rect 5850 700 7150 750
rect 5600 650 5750 700
rect 5900 650 7150 700
rect 5600 600 5800 650
rect 5950 600 7150 650
rect 5600 550 5850 600
rect 5600 -1400 5900 550
rect 7100 400 7150 600
rect 6200 350 7150 400
rect 6250 300 7150 350
rect 6100 250 6150 300
rect 6300 250 7150 300
rect 6100 200 6200 250
rect 6350 200 7150 250
rect 6100 150 6250 200
rect 6400 150 7150 200
rect 6100 100 6300 150
rect 6450 100 7150 150
rect 6100 50 6350 100
rect 6100 -1400 6400 50
rect 7100 -100 7150 100
rect 6700 -150 7150 -100
rect 6750 -200 7150 -150
rect 6600 -250 6650 -200
rect 6800 -250 7150 -200
rect 6600 -300 6700 -250
rect 6850 -300 7150 -250
rect 6600 -350 6750 -300
rect 6900 -350 7150 -300
rect 6600 -400 6800 -350
rect 6950 -400 7150 -350
rect 6600 -450 6850 -400
rect 6600 -1400 6900 -450
rect 7100 -1400 7150 -400
rect -650 -1450 7150 -1400
rect 7650 -1950 7700 7650
rect -1200 -2000 7700 -1950
<< via3 >>
rect -1150 7150 7650 7650
rect -1150 -1950 -650 7150
rect 7150 4300 7650 7150
rect 7150 2500 7650 3800
rect 7150 -1450 7650 2300
rect 1150 -1950 7650 -1450
<< metal4 >>
rect -1200 7650 7700 7700
rect -1200 -1950 -1150 7650
rect -650 7100 7150 7150
rect -650 3600 -600 7100
rect 7100 4300 7150 7100
rect 7650 4300 7700 7650
rect 7100 3800 7700 4300
rect -650 3400 3600 3600
rect -650 2900 3000 3400
rect -650 -1950 -600 2900
rect 7100 2500 7150 3800
rect 7650 2500 7700 3800
rect 7100 2300 7700 2500
rect 7100 -1400 7150 2300
rect -1200 -2000 -600 -1950
rect 1100 -1450 7150 -1400
rect 1100 -1950 1150 -1450
rect 7650 -1950 7700 2300
rect 1100 -2000 7700 -1950
<< via4 >>
rect 3000 2900 3600 3400
<< metal5 >>
rect 0 6000 6500 6500
rect 0 -300 500 6000
rect 800 5200 5700 5700
rect 800 500 1300 5200
rect 1600 4400 4900 4900
rect 1600 1300 2100 4400
rect 2400 3400 3700 3500
rect 2400 2900 3000 3400
rect 3600 2900 3700 3400
rect 2400 2800 3700 2900
rect 2400 2100 2900 2800
rect 4400 2100 4900 4400
rect 2400 1600 4900 2100
rect 5200 1300 5700 5200
rect 1600 800 5700 1300
rect 6000 500 6500 6000
rect 800 0 6500 500
rect 0 -400 600 -300
rect 0 -500 700 -400
rect 0 -2200 800 -500
<< end >>
