magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< locali >>
rect 5634 9881 10346 9915
rect 3386 8467 5634 8501
rect 3754 7053 10346 7087
rect 3733 6790 3952 6824
rect 3918 6308 3952 6790
rect 3386 5639 6514 5673
rect 4780 4225 10346 4259
rect 3386 2811 5148 2845
rect 3715 2541 3900 2575
rect 3715 2176 3749 2541
rect 3582 2142 3749 2176
rect 5148 1397 10346 1431
rect 3386 -17 10346 17
<< metal1 >>
rect 10314 9872 10378 9924
rect 2980 9140 3467 9168
rect 4786 9165 4850 9217
rect 3354 8458 3418 8510
rect 2896 7801 3467 7829
rect 3550 7789 3614 7841
rect 10314 7044 10378 7096
rect 5880 6337 5944 6389
rect 2896 6160 3615 6188
rect 3064 5912 3515 5940
rect 3354 5630 3418 5682
rect 3232 5372 3482 5400
rect 2812 5248 3615 5276
rect 2980 5124 3748 5152
rect 4896 4923 4960 4975
rect 1553 4308 2896 4336
rect 10314 4216 10378 4268
rect 383 4148 3148 4176
rect 4254 3493 4318 3545
rect 3232 3332 3615 3360
rect 3148 3084 3515 3112
rect 3354 2802 3418 2854
rect 3951 2284 4015 2336
rect 3148 2145 3467 2173
rect 4622 2111 4686 2163
rect 10314 1388 10378 1440
rect 3435 643 3499 695
rect 8524 681 8588 733
rect 3354 -26 3418 26
<< metal2 >>
rect -57 17699 -29 17727
rect 1539 4322 1567 6401
rect 369 1414 397 4162
rect 1844 861 1900 909
rect 137 538 203 590
rect 2798 0 2826 9938
rect 2882 0 2910 9938
rect 2966 0 2994 9938
rect 3050 0 3078 9938
rect 3134 0 3162 9938
rect 3218 0 3246 9938
rect 10318 9874 10374 9922
rect 4818 9177 10430 9205
rect 3358 8460 3414 8508
rect 3568 7391 3596 7815
rect 10318 7046 10374 7094
rect 5912 6349 10430 6377
rect 3358 5632 3414 5680
rect 4928 4935 10430 4963
rect 10318 4218 10374 4266
rect 4258 3495 4314 3543
rect 3358 2804 3414 2852
rect 3955 2286 4011 2334
rect 4640 1713 4668 2137
rect 10318 1390 10374 1438
rect 8556 707 10430 721
rect 8542 693 10430 707
rect 3453 655 3481 683
rect 8542 283 8570 693
rect 3358 -24 3414 24
<< metal3 >>
rect 10271 9866 10421 9930
rect 3311 8452 3461 8516
rect 2812 7361 3582 7421
rect 10271 7038 10421 7102
rect 3311 5624 3461 5688
rect 10271 4210 10421 4274
rect 3064 3489 4286 3549
rect 3311 2796 3461 2860
rect 3232 2280 3983 2340
rect 2980 1683 4654 1743
rect 1228 1365 1326 1463
rect 10271 1382 10421 1446
rect 1872 855 3232 915
rect 3148 253 8556 313
rect 1228 -49 1326 49
rect 3311 -32 3461 32
<< metal4 >>
rect 335 5606 401 18415
rect 1439 5623 1505 18432
rect 3353 -33 3419 8517
rect 10313 1381 10379 9931
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_0
timestamp 1661296025
transform 1 0 3357 0 1 8451
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_1
timestamp 1661296025
transform 1 0 10317 0 1 9865
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_2
timestamp 1661296025
transform 1 0 3357 0 1 8451
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_3
timestamp 1661296025
transform 1 0 10317 0 1 7037
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_4
timestamp 1661296025
transform 1 0 3357 0 1 5623
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_5
timestamp 1661296025
transform 1 0 10317 0 1 7037
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_6
timestamp 1661296025
transform 1 0 3357 0 1 5623
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_7
timestamp 1661296025
transform 1 0 10317 0 1 4209
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_8
timestamp 1661296025
transform 1 0 3357 0 1 2795
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_9
timestamp 1661296025
transform 1 0 10317 0 1 4209
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_10
timestamp 1661296025
transform 1 0 3357 0 1 2795
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_11
timestamp 1661296025
transform 1 0 10317 0 1 1381
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_12
timestamp 1661296025
transform 1 0 3357 0 1 -33
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_13
timestamp 1661296025
transform 1 0 10317 0 1 1381
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_14
timestamp 1661296025
transform 1 0 4257 0 1 3486
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_15
timestamp 1661296025
transform 1 0 4257 0 1 3486
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_16
timestamp 1661296025
transform 1 0 3586 0 1 3313
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_17
timestamp 1661296025
transform 1 0 3486 0 1 3065
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_18
timestamp 1661296025
transform 1 0 4625 0 1 2104
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_19
timestamp 1661296025
transform 1 0 3954 0 1 2277
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_20
timestamp 1661296025
transform 1 0 3954 0 1 2277
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_21
timestamp 1661296025
transform 1 0 3438 0 1 2126
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_22
timestamp 1661296025
transform 1 0 8527 0 1 674
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_23
timestamp 1661296025
transform 1 0 8527 0 1 674
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_24
timestamp 1661296025
transform 1 0 3438 0 1 636
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_25
timestamp 1661296025
transform 1 0 5883 0 1 6330
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_26
timestamp 1661296025
transform 1 0 3586 0 1 6141
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_27
timestamp 1661296025
transform 1 0 3486 0 1 5893
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_28
timestamp 1661296025
transform 1 0 4899 0 1 4916
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_29
timestamp 1661296025
transform 1 0 3719 0 1 5105
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_30
timestamp 1661296025
transform 1 0 3586 0 1 5229
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_31
timestamp 1661296025
transform 1 0 3453 0 1 5353
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_32
timestamp 1661296025
transform 1 0 3438 0 1 7782
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_33
timestamp 1661296025
transform 1 0 3553 0 1 7782
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_34
timestamp 1661296025
transform 1 0 4789 0 1 9158
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_35
timestamp 1661296025
transform 1 0 3438 0 1 9121
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_0
timestamp 1661296025
transform 1 0 3354 0 1 8452
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_1
timestamp 1661296025
transform 1 0 10314 0 1 9866
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_2
timestamp 1661296025
transform 1 0 3354 0 1 8452
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_3
timestamp 1661296025
transform 1 0 10314 0 1 7038
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_4
timestamp 1661296025
transform 1 0 3354 0 1 5624
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_5
timestamp 1661296025
transform 1 0 10314 0 1 7038
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_6
timestamp 1661296025
transform 1 0 3354 0 1 5624
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_7
timestamp 1661296025
transform 1 0 10314 0 1 4210
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_8
timestamp 1661296025
transform 1 0 3354 0 1 2796
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_9
timestamp 1661296025
transform 1 0 10314 0 1 4210
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_10
timestamp 1661296025
transform 1 0 3354 0 1 2796
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_11
timestamp 1661296025
transform 1 0 10314 0 1 1382
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_12
timestamp 1661296025
transform 1 0 3354 0 1 -32
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_13
timestamp 1661296025
transform 1 0 10314 0 1 1382
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_14
timestamp 1661296025
transform 1 0 4254 0 1 3487
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_15
timestamp 1661296025
transform 1 0 4254 0 1 3487
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_16
timestamp 1661296025
transform 1 0 3200 0 1 3314
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_17
timestamp 1661296025
transform 1 0 3116 0 1 3066
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_18
timestamp 1661296025
transform 1 0 4622 0 1 2105
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_19
timestamp 1661296025
transform 1 0 3951 0 1 2278
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_20
timestamp 1661296025
transform 1 0 3951 0 1 2278
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_21
timestamp 1661296025
transform 1 0 3116 0 1 2127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_22
timestamp 1661296025
transform 1 0 8524 0 1 675
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_23
timestamp 1661296025
transform 1 0 8524 0 1 675
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_24
timestamp 1661296025
transform 1 0 3435 0 1 637
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_25
timestamp 1661296025
transform 1 0 5880 0 1 6331
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_26
timestamp 1661296025
transform 1 0 2864 0 1 6142
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_27
timestamp 1661296025
transform 1 0 3032 0 1 5894
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_28
timestamp 1661296025
transform 1 0 2864 0 1 4290
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_29
timestamp 1661296025
transform 1 0 1521 0 1 4290
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_30
timestamp 1661296025
transform 1 0 4896 0 1 4917
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_31
timestamp 1661296025
transform 1 0 2948 0 1 5106
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_32
timestamp 1661296025
transform 1 0 2780 0 1 5230
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_33
timestamp 1661296025
transform 1 0 3200 0 1 5354
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_34
timestamp 1661296025
transform 1 0 2864 0 1 7783
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_35
timestamp 1661296025
transform 1 0 3550 0 1 7783
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_36
timestamp 1661296025
transform 1 0 4786 0 1 9159
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_37
timestamp 1661296025
transform 1 0 2948 0 1 9122
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_38
timestamp 1661296025
transform 1 0 3116 0 1 4130
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_39
timestamp 1661296025
transform 1 0 351 0 1 4130
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_0
timestamp 1661296025
transform 1 0 3353 0 1 8447
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_1
timestamp 1661296025
transform 1 0 10313 0 1 9861
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_2
timestamp 1661296025
transform 1 0 3353 0 1 8447
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_3
timestamp 1661296025
transform 1 0 10313 0 1 7033
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_4
timestamp 1661296025
transform 1 0 3353 0 1 5619
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_5
timestamp 1661296025
transform 1 0 10313 0 1 7033
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_6
timestamp 1661296025
transform 1 0 3353 0 1 5619
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_7
timestamp 1661296025
transform 1 0 10313 0 1 4205
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_8
timestamp 1661296025
transform 1 0 3353 0 1 2791
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_9
timestamp 1661296025
transform 1 0 10313 0 1 4205
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_10
timestamp 1661296025
transform 1 0 3353 0 1 2791
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_11
timestamp 1661296025
transform 1 0 10313 0 1 1377
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_12
timestamp 1661296025
transform 1 0 3353 0 1 -37
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_13
timestamp 1661296025
transform 1 0 10313 0 1 1377
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_14
timestamp 1661296025
transform 1 0 4253 0 1 3482
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_15
timestamp 1661296025
transform 1 0 3950 0 1 2273
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_16
timestamp 1661296025
transform 1 0 3950 0 1 2273
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_17
timestamp 1661296025
transform 1 0 1839 0 1 848
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_0
timestamp 1661296025
transform 1 0 3348 0 1 8451
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_1
timestamp 1661296025
transform 1 0 10308 0 1 9865
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_2
timestamp 1661296025
transform 1 0 3348 0 1 8451
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_3
timestamp 1661296025
transform 1 0 10308 0 1 7037
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_4
timestamp 1661296025
transform 1 0 3348 0 1 5623
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_5
timestamp 1661296025
transform 1 0 10308 0 1 7037
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_6
timestamp 1661296025
transform 1 0 3348 0 1 5623
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_7
timestamp 1661296025
transform 1 0 10308 0 1 4209
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_8
timestamp 1661296025
transform 1 0 3348 0 1 2795
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_9
timestamp 1661296025
transform 1 0 10308 0 1 4209
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_10
timestamp 1661296025
transform 1 0 3348 0 1 2795
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_11
timestamp 1661296025
transform 1 0 10308 0 1 1381
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_12
timestamp 1661296025
transform 1 0 3348 0 1 -33
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_13
timestamp 1661296025
transform 1 0 10308 0 1 1381
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_0
timestamp 1661296025
transform 1 0 3031 0 1 3482
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_1
timestamp 1661296025
transform 1 0 2947 0 1 1676
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_2
timestamp 1661296025
transform 1 0 4621 0 1 1676
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_3
timestamp 1661296025
transform 1 0 3199 0 1 2273
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_4
timestamp 1661296025
transform 1 0 3115 0 1 246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_5
timestamp 1661296025
transform 1 0 8523 0 1 246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_6
timestamp 1661296025
transform 1 0 2779 0 1 7354
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_7
timestamp 1661296025
transform 1 0 3549 0 1 7354
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_8
timestamp 1661296025
transform 1 0 3199 0 1 848
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_delay_chain  sky130_sram_1r1w_24x128_8_delay_chain_0
timestamp 1661296025
transform 1 0 0 0 -1 18382
box -75 -50 1876 12783
use sky130_sram_1r1w_24x128_8_dff_buf_array  sky130_sram_1r1w_24x128_8_dff_buf_array_0
timestamp 1661296025
transform 1 0 0 0 1 0
box -36 -49 2590 1471
use sky130_sram_1r1w_24x128_8_pand2  sky130_sram_1r1w_24x128_8_pand2_0
timestamp 1661296025
transform 1 0 3386 0 1 2828
box -36 -17 1430 1471
use sky130_sram_1r1w_24x128_8_pand2  sky130_sram_1r1w_24x128_8_pand2_1
timestamp 1661296025
transform 1 0 3754 0 -1 2828
box -36 -17 1430 1471
use sky130_sram_1r1w_24x128_8_pand3  sky130_sram_1r1w_24x128_8_pand3_0
timestamp 1661296025
transform 1 0 3386 0 -1 5656
box -36 -17 2718 1471
use sky130_sram_1r1w_24x128_8_pdriver_0  sky130_sram_1r1w_24x128_8_pdriver_0_0
timestamp 1661296025
transform 1 0 3386 0 1 0
box -36 -17 6996 1471
use sky130_sram_1r1w_24x128_8_pdriver_1  sky130_sram_1r1w_24x128_8_pdriver_1_0
timestamp 1661296025
transform 1 0 3386 0 1 8484
box -36 -17 2284 1471
use sky130_sram_1r1w_24x128_8_pdriver_4  sky130_sram_1r1w_24x128_8_pdriver_4_0
timestamp 1661296025
transform 1 0 3854 0 1 5656
box -36 -17 2696 1471
use sky130_sram_1r1w_24x128_8_pinv  sky130_sram_1r1w_24x128_8_pinv_0
timestamp 1661296025
transform 1 0 3386 0 -1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv  sky130_sram_1r1w_24x128_8_pinv_1
timestamp 1661296025
transform 1 0 3386 0 -1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pnand2_0  sky130_sram_1r1w_24x128_8_pnand2_0_0
timestamp 1661296025
transform 1 0 3386 0 1 5656
box -36 -17 504 1471
<< labels >>
rlabel metal2 s 137 538 203 590 4 csb
port 1 nsew
rlabel metal2 s 4818 9177 10430 9205 4 wl_en
port 2 nsew
rlabel metal2 s 4928 4935 10430 4963 4 w_en
port 3 nsew
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
port 4 nsew
rlabel metal2 s 5912 6349 10430 6377 4 p_en_bar
port 5 nsew
rlabel metal2 s 3453 655 3481 683 4 clk
port 6 nsew
rlabel metal2 s 8556 693 10430 721 4 clk_buf
port 7 nsew
rlabel metal4 s 10313 1381 10379 9931 4 vdd
port 8 nsew
rlabel metal4 s 335 5606 401 18415 4 vdd
port 8 nsew
rlabel metal3 s 1228 1365 1326 1463 4 vdd
port 8 nsew
rlabel metal4 s 1439 5623 1505 18432 4 gnd
port 9 nsew
rlabel metal4 s 3353 -33 3419 8517 4 gnd
port 9 nsew
rlabel metal3 s 1228 -49 1326 49 4 gnd
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 10430 18542
<< end >>
