magic
tech sky130B
magscale 1 2
timestamp 1659664599
<< error_p >>
rect -1421 481 -1363 487
rect -1229 481 -1171 487
rect -1037 481 -979 487
rect -845 481 -787 487
rect -653 481 -595 487
rect -461 481 -403 487
rect -269 481 -211 487
rect -77 481 -19 487
rect 115 481 173 487
rect 307 481 365 487
rect 499 481 557 487
rect 691 481 749 487
rect 883 481 941 487
rect 1075 481 1133 487
rect 1267 481 1325 487
rect 1459 481 1517 487
rect -1421 447 -1409 481
rect -1229 447 -1217 481
rect -1037 447 -1025 481
rect -845 447 -833 481
rect -653 447 -641 481
rect -461 447 -449 481
rect -269 447 -257 481
rect -77 447 -65 481
rect 115 447 127 481
rect 307 447 319 481
rect 499 447 511 481
rect 691 447 703 481
rect 883 447 895 481
rect 1075 447 1087 481
rect 1267 447 1279 481
rect 1459 447 1471 481
rect -1421 441 -1363 447
rect -1229 441 -1171 447
rect -1037 441 -979 447
rect -845 441 -787 447
rect -653 441 -595 447
rect -461 441 -403 447
rect -269 441 -211 447
rect -77 441 -19 447
rect 115 441 173 447
rect 307 441 365 447
rect 499 441 557 447
rect 691 441 749 447
rect 883 441 941 447
rect 1075 441 1133 447
rect 1267 441 1325 447
rect 1459 441 1517 447
rect -1517 -447 -1459 -441
rect -1325 -447 -1267 -441
rect -1133 -447 -1075 -441
rect -941 -447 -883 -441
rect -749 -447 -691 -441
rect -557 -447 -499 -441
rect -365 -447 -307 -441
rect -173 -447 -115 -441
rect 19 -447 77 -441
rect 211 -447 269 -441
rect 403 -447 461 -441
rect 595 -447 653 -441
rect 787 -447 845 -441
rect 979 -447 1037 -441
rect 1171 -447 1229 -441
rect 1363 -447 1421 -441
rect -1517 -481 -1505 -447
rect -1325 -481 -1313 -447
rect -1133 -481 -1121 -447
rect -941 -481 -929 -447
rect -749 -481 -737 -447
rect -557 -481 -545 -447
rect -365 -481 -353 -447
rect -173 -481 -161 -447
rect 19 -481 31 -447
rect 211 -481 223 -447
rect 403 -481 415 -447
rect 595 -481 607 -447
rect 787 -481 799 -447
rect 979 -481 991 -447
rect 1171 -481 1183 -447
rect 1363 -481 1375 -447
rect -1517 -487 -1459 -481
rect -1325 -487 -1267 -481
rect -1133 -487 -1075 -481
rect -941 -487 -883 -481
rect -749 -487 -691 -481
rect -557 -487 -499 -481
rect -365 -487 -307 -481
rect -173 -487 -115 -481
rect 19 -487 77 -481
rect 211 -487 269 -481
rect 403 -487 461 -481
rect 595 -487 653 -481
rect 787 -487 845 -481
rect 979 -487 1037 -481
rect 1171 -487 1229 -481
rect 1363 -487 1421 -481
<< nwell >>
rect -1703 -619 1703 619
<< pmos >>
rect -1503 -400 -1473 400
rect -1407 -400 -1377 400
rect -1311 -400 -1281 400
rect -1215 -400 -1185 400
rect -1119 -400 -1089 400
rect -1023 -400 -993 400
rect -927 -400 -897 400
rect -831 -400 -801 400
rect -735 -400 -705 400
rect -639 -400 -609 400
rect -543 -400 -513 400
rect -447 -400 -417 400
rect -351 -400 -321 400
rect -255 -400 -225 400
rect -159 -400 -129 400
rect -63 -400 -33 400
rect 33 -400 63 400
rect 129 -400 159 400
rect 225 -400 255 400
rect 321 -400 351 400
rect 417 -400 447 400
rect 513 -400 543 400
rect 609 -400 639 400
rect 705 -400 735 400
rect 801 -400 831 400
rect 897 -400 927 400
rect 993 -400 1023 400
rect 1089 -400 1119 400
rect 1185 -400 1215 400
rect 1281 -400 1311 400
rect 1377 -400 1407 400
rect 1473 -400 1503 400
<< pdiff >>
rect -1565 388 -1503 400
rect -1565 -388 -1553 388
rect -1519 -388 -1503 388
rect -1565 -400 -1503 -388
rect -1473 388 -1407 400
rect -1473 -388 -1457 388
rect -1423 -388 -1407 388
rect -1473 -400 -1407 -388
rect -1377 388 -1311 400
rect -1377 -388 -1361 388
rect -1327 -388 -1311 388
rect -1377 -400 -1311 -388
rect -1281 388 -1215 400
rect -1281 -388 -1265 388
rect -1231 -388 -1215 388
rect -1281 -400 -1215 -388
rect -1185 388 -1119 400
rect -1185 -388 -1169 388
rect -1135 -388 -1119 388
rect -1185 -400 -1119 -388
rect -1089 388 -1023 400
rect -1089 -388 -1073 388
rect -1039 -388 -1023 388
rect -1089 -400 -1023 -388
rect -993 388 -927 400
rect -993 -388 -977 388
rect -943 -388 -927 388
rect -993 -400 -927 -388
rect -897 388 -831 400
rect -897 -388 -881 388
rect -847 -388 -831 388
rect -897 -400 -831 -388
rect -801 388 -735 400
rect -801 -388 -785 388
rect -751 -388 -735 388
rect -801 -400 -735 -388
rect -705 388 -639 400
rect -705 -388 -689 388
rect -655 -388 -639 388
rect -705 -400 -639 -388
rect -609 388 -543 400
rect -609 -388 -593 388
rect -559 -388 -543 388
rect -609 -400 -543 -388
rect -513 388 -447 400
rect -513 -388 -497 388
rect -463 -388 -447 388
rect -513 -400 -447 -388
rect -417 388 -351 400
rect -417 -388 -401 388
rect -367 -388 -351 388
rect -417 -400 -351 -388
rect -321 388 -255 400
rect -321 -388 -305 388
rect -271 -388 -255 388
rect -321 -400 -255 -388
rect -225 388 -159 400
rect -225 -388 -209 388
rect -175 -388 -159 388
rect -225 -400 -159 -388
rect -129 388 -63 400
rect -129 -388 -113 388
rect -79 -388 -63 388
rect -129 -400 -63 -388
rect -33 388 33 400
rect -33 -388 -17 388
rect 17 -388 33 388
rect -33 -400 33 -388
rect 63 388 129 400
rect 63 -388 79 388
rect 113 -388 129 388
rect 63 -400 129 -388
rect 159 388 225 400
rect 159 -388 175 388
rect 209 -388 225 388
rect 159 -400 225 -388
rect 255 388 321 400
rect 255 -388 271 388
rect 305 -388 321 388
rect 255 -400 321 -388
rect 351 388 417 400
rect 351 -388 367 388
rect 401 -388 417 388
rect 351 -400 417 -388
rect 447 388 513 400
rect 447 -388 463 388
rect 497 -388 513 388
rect 447 -400 513 -388
rect 543 388 609 400
rect 543 -388 559 388
rect 593 -388 609 388
rect 543 -400 609 -388
rect 639 388 705 400
rect 639 -388 655 388
rect 689 -388 705 388
rect 639 -400 705 -388
rect 735 388 801 400
rect 735 -388 751 388
rect 785 -388 801 388
rect 735 -400 801 -388
rect 831 388 897 400
rect 831 -388 847 388
rect 881 -388 897 388
rect 831 -400 897 -388
rect 927 388 993 400
rect 927 -388 943 388
rect 977 -388 993 388
rect 927 -400 993 -388
rect 1023 388 1089 400
rect 1023 -388 1039 388
rect 1073 -388 1089 388
rect 1023 -400 1089 -388
rect 1119 388 1185 400
rect 1119 -388 1135 388
rect 1169 -388 1185 388
rect 1119 -400 1185 -388
rect 1215 388 1281 400
rect 1215 -388 1231 388
rect 1265 -388 1281 388
rect 1215 -400 1281 -388
rect 1311 388 1377 400
rect 1311 -388 1327 388
rect 1361 -388 1377 388
rect 1311 -400 1377 -388
rect 1407 388 1473 400
rect 1407 -388 1423 388
rect 1457 -388 1473 388
rect 1407 -400 1473 -388
rect 1503 388 1565 400
rect 1503 -388 1519 388
rect 1553 -388 1565 388
rect 1503 -400 1565 -388
<< pdiffc >>
rect -1553 -388 -1519 388
rect -1457 -388 -1423 388
rect -1361 -388 -1327 388
rect -1265 -388 -1231 388
rect -1169 -388 -1135 388
rect -1073 -388 -1039 388
rect -977 -388 -943 388
rect -881 -388 -847 388
rect -785 -388 -751 388
rect -689 -388 -655 388
rect -593 -388 -559 388
rect -497 -388 -463 388
rect -401 -388 -367 388
rect -305 -388 -271 388
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect 271 -388 305 388
rect 367 -388 401 388
rect 463 -388 497 388
rect 559 -388 593 388
rect 655 -388 689 388
rect 751 -388 785 388
rect 847 -388 881 388
rect 943 -388 977 388
rect 1039 -388 1073 388
rect 1135 -388 1169 388
rect 1231 -388 1265 388
rect 1327 -388 1361 388
rect 1423 -388 1457 388
rect 1519 -388 1553 388
<< nsubdiff >>
rect -1667 549 -1571 583
rect 1571 549 1667 583
rect -1667 487 -1633 549
rect 1633 487 1667 549
rect -1667 -549 -1633 -487
rect 1633 -549 1667 -487
rect -1667 -583 -1571 -549
rect 1571 -583 1667 -549
<< nsubdiffcont >>
rect -1571 549 1571 583
rect -1667 -487 -1633 487
rect 1633 -487 1667 487
rect -1571 -583 1571 -549
<< poly >>
rect -1425 481 -1359 497
rect -1425 447 -1409 481
rect -1375 447 -1359 481
rect -1425 431 -1359 447
rect -1233 481 -1167 497
rect -1233 447 -1217 481
rect -1183 447 -1167 481
rect -1233 431 -1167 447
rect -1041 481 -975 497
rect -1041 447 -1025 481
rect -991 447 -975 481
rect -1041 431 -975 447
rect -849 481 -783 497
rect -849 447 -833 481
rect -799 447 -783 481
rect -849 431 -783 447
rect -657 481 -591 497
rect -657 447 -641 481
rect -607 447 -591 481
rect -657 431 -591 447
rect -465 481 -399 497
rect -465 447 -449 481
rect -415 447 -399 481
rect -465 431 -399 447
rect -273 481 -207 497
rect -273 447 -257 481
rect -223 447 -207 481
rect -273 431 -207 447
rect -81 481 -15 497
rect -81 447 -65 481
rect -31 447 -15 481
rect -81 431 -15 447
rect 111 481 177 497
rect 111 447 127 481
rect 161 447 177 481
rect 111 431 177 447
rect 303 481 369 497
rect 303 447 319 481
rect 353 447 369 481
rect 303 431 369 447
rect 495 481 561 497
rect 495 447 511 481
rect 545 447 561 481
rect 495 431 561 447
rect 687 481 753 497
rect 687 447 703 481
rect 737 447 753 481
rect 687 431 753 447
rect 879 481 945 497
rect 879 447 895 481
rect 929 447 945 481
rect 879 431 945 447
rect 1071 481 1137 497
rect 1071 447 1087 481
rect 1121 447 1137 481
rect 1071 431 1137 447
rect 1263 481 1329 497
rect 1263 447 1279 481
rect 1313 447 1329 481
rect 1263 431 1329 447
rect 1455 481 1521 497
rect 1455 447 1471 481
rect 1505 447 1521 481
rect 1455 431 1521 447
rect -1503 400 -1473 426
rect -1407 400 -1377 431
rect -1311 400 -1281 426
rect -1215 400 -1185 431
rect -1119 400 -1089 426
rect -1023 400 -993 431
rect -927 400 -897 426
rect -831 400 -801 431
rect -735 400 -705 426
rect -639 400 -609 431
rect -543 400 -513 426
rect -447 400 -417 431
rect -351 400 -321 426
rect -255 400 -225 431
rect -159 400 -129 426
rect -63 400 -33 431
rect 33 400 63 426
rect 129 400 159 431
rect 225 400 255 426
rect 321 400 351 431
rect 417 400 447 426
rect 513 400 543 431
rect 609 400 639 426
rect 705 400 735 431
rect 801 400 831 426
rect 897 400 927 431
rect 993 400 1023 426
rect 1089 400 1119 431
rect 1185 400 1215 426
rect 1281 400 1311 431
rect 1377 400 1407 426
rect 1473 400 1503 431
rect -1503 -431 -1473 -400
rect -1407 -426 -1377 -400
rect -1311 -431 -1281 -400
rect -1215 -426 -1185 -400
rect -1119 -431 -1089 -400
rect -1023 -426 -993 -400
rect -927 -431 -897 -400
rect -831 -426 -801 -400
rect -735 -431 -705 -400
rect -639 -426 -609 -400
rect -543 -431 -513 -400
rect -447 -426 -417 -400
rect -351 -431 -321 -400
rect -255 -426 -225 -400
rect -159 -431 -129 -400
rect -63 -426 -33 -400
rect 33 -431 63 -400
rect 129 -426 159 -400
rect 225 -431 255 -400
rect 321 -426 351 -400
rect 417 -431 447 -400
rect 513 -426 543 -400
rect 609 -431 639 -400
rect 705 -426 735 -400
rect 801 -431 831 -400
rect 897 -426 927 -400
rect 993 -431 1023 -400
rect 1089 -426 1119 -400
rect 1185 -431 1215 -400
rect 1281 -426 1311 -400
rect 1377 -431 1407 -400
rect 1473 -426 1503 -400
rect -1521 -447 -1455 -431
rect -1521 -481 -1505 -447
rect -1471 -481 -1455 -447
rect -1521 -497 -1455 -481
rect -1329 -447 -1263 -431
rect -1329 -481 -1313 -447
rect -1279 -481 -1263 -447
rect -1329 -497 -1263 -481
rect -1137 -447 -1071 -431
rect -1137 -481 -1121 -447
rect -1087 -481 -1071 -447
rect -1137 -497 -1071 -481
rect -945 -447 -879 -431
rect -945 -481 -929 -447
rect -895 -481 -879 -447
rect -945 -497 -879 -481
rect -753 -447 -687 -431
rect -753 -481 -737 -447
rect -703 -481 -687 -447
rect -753 -497 -687 -481
rect -561 -447 -495 -431
rect -561 -481 -545 -447
rect -511 -481 -495 -447
rect -561 -497 -495 -481
rect -369 -447 -303 -431
rect -369 -481 -353 -447
rect -319 -481 -303 -447
rect -369 -497 -303 -481
rect -177 -447 -111 -431
rect -177 -481 -161 -447
rect -127 -481 -111 -447
rect -177 -497 -111 -481
rect 15 -447 81 -431
rect 15 -481 31 -447
rect 65 -481 81 -447
rect 15 -497 81 -481
rect 207 -447 273 -431
rect 207 -481 223 -447
rect 257 -481 273 -447
rect 207 -497 273 -481
rect 399 -447 465 -431
rect 399 -481 415 -447
rect 449 -481 465 -447
rect 399 -497 465 -481
rect 591 -447 657 -431
rect 591 -481 607 -447
rect 641 -481 657 -447
rect 591 -497 657 -481
rect 783 -447 849 -431
rect 783 -481 799 -447
rect 833 -481 849 -447
rect 783 -497 849 -481
rect 975 -447 1041 -431
rect 975 -481 991 -447
rect 1025 -481 1041 -447
rect 975 -497 1041 -481
rect 1167 -447 1233 -431
rect 1167 -481 1183 -447
rect 1217 -481 1233 -447
rect 1167 -497 1233 -481
rect 1359 -447 1425 -431
rect 1359 -481 1375 -447
rect 1409 -481 1425 -447
rect 1359 -497 1425 -481
<< polycont >>
rect -1409 447 -1375 481
rect -1217 447 -1183 481
rect -1025 447 -991 481
rect -833 447 -799 481
rect -641 447 -607 481
rect -449 447 -415 481
rect -257 447 -223 481
rect -65 447 -31 481
rect 127 447 161 481
rect 319 447 353 481
rect 511 447 545 481
rect 703 447 737 481
rect 895 447 929 481
rect 1087 447 1121 481
rect 1279 447 1313 481
rect 1471 447 1505 481
rect -1505 -481 -1471 -447
rect -1313 -481 -1279 -447
rect -1121 -481 -1087 -447
rect -929 -481 -895 -447
rect -737 -481 -703 -447
rect -545 -481 -511 -447
rect -353 -481 -319 -447
rect -161 -481 -127 -447
rect 31 -481 65 -447
rect 223 -481 257 -447
rect 415 -481 449 -447
rect 607 -481 641 -447
rect 799 -481 833 -447
rect 991 -481 1025 -447
rect 1183 -481 1217 -447
rect 1375 -481 1409 -447
<< locali >>
rect -1667 549 -1571 583
rect 1571 549 1667 583
rect -1667 487 -1633 549
rect 1633 487 1667 549
rect -1425 447 -1409 481
rect -1375 447 -1359 481
rect -1233 447 -1217 481
rect -1183 447 -1167 481
rect -1041 447 -1025 481
rect -991 447 -975 481
rect -849 447 -833 481
rect -799 447 -783 481
rect -657 447 -641 481
rect -607 447 -591 481
rect -465 447 -449 481
rect -415 447 -399 481
rect -273 447 -257 481
rect -223 447 -207 481
rect -81 447 -65 481
rect -31 447 -15 481
rect 111 447 127 481
rect 161 447 177 481
rect 303 447 319 481
rect 353 447 369 481
rect 495 447 511 481
rect 545 447 561 481
rect 687 447 703 481
rect 737 447 753 481
rect 879 447 895 481
rect 929 447 945 481
rect 1071 447 1087 481
rect 1121 447 1137 481
rect 1263 447 1279 481
rect 1313 447 1329 481
rect 1455 447 1471 481
rect 1505 447 1521 481
rect -1553 388 -1519 404
rect -1553 -404 -1519 -388
rect -1457 388 -1423 404
rect -1457 -404 -1423 -388
rect -1361 388 -1327 404
rect -1361 -404 -1327 -388
rect -1265 388 -1231 404
rect -1265 -404 -1231 -388
rect -1169 388 -1135 404
rect -1169 -404 -1135 -388
rect -1073 388 -1039 404
rect -1073 -404 -1039 -388
rect -977 388 -943 404
rect -977 -404 -943 -388
rect -881 388 -847 404
rect -881 -404 -847 -388
rect -785 388 -751 404
rect -785 -404 -751 -388
rect -689 388 -655 404
rect -689 -404 -655 -388
rect -593 388 -559 404
rect -593 -404 -559 -388
rect -497 388 -463 404
rect -497 -404 -463 -388
rect -401 388 -367 404
rect -401 -404 -367 -388
rect -305 388 -271 404
rect -305 -404 -271 -388
rect -209 388 -175 404
rect -209 -404 -175 -388
rect -113 388 -79 404
rect -113 -404 -79 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 79 388 113 404
rect 79 -404 113 -388
rect 175 388 209 404
rect 175 -404 209 -388
rect 271 388 305 404
rect 271 -404 305 -388
rect 367 388 401 404
rect 367 -404 401 -388
rect 463 388 497 404
rect 463 -404 497 -388
rect 559 388 593 404
rect 559 -404 593 -388
rect 655 388 689 404
rect 655 -404 689 -388
rect 751 388 785 404
rect 751 -404 785 -388
rect 847 388 881 404
rect 847 -404 881 -388
rect 943 388 977 404
rect 943 -404 977 -388
rect 1039 388 1073 404
rect 1039 -404 1073 -388
rect 1135 388 1169 404
rect 1135 -404 1169 -388
rect 1231 388 1265 404
rect 1231 -404 1265 -388
rect 1327 388 1361 404
rect 1327 -404 1361 -388
rect 1423 388 1457 404
rect 1423 -404 1457 -388
rect 1519 388 1553 404
rect 1519 -404 1553 -388
rect -1521 -481 -1505 -447
rect -1471 -481 -1455 -447
rect -1329 -481 -1313 -447
rect -1279 -481 -1263 -447
rect -1137 -481 -1121 -447
rect -1087 -481 -1071 -447
rect -945 -481 -929 -447
rect -895 -481 -879 -447
rect -753 -481 -737 -447
rect -703 -481 -687 -447
rect -561 -481 -545 -447
rect -511 -481 -495 -447
rect -369 -481 -353 -447
rect -319 -481 -303 -447
rect -177 -481 -161 -447
rect -127 -481 -111 -447
rect 15 -481 31 -447
rect 65 -481 81 -447
rect 207 -481 223 -447
rect 257 -481 273 -447
rect 399 -481 415 -447
rect 449 -481 465 -447
rect 591 -481 607 -447
rect 641 -481 657 -447
rect 783 -481 799 -447
rect 833 -481 849 -447
rect 975 -481 991 -447
rect 1025 -481 1041 -447
rect 1167 -481 1183 -447
rect 1217 -481 1233 -447
rect 1359 -481 1375 -447
rect 1409 -481 1425 -447
rect -1667 -549 -1633 -487
rect 1633 -549 1667 -487
rect -1667 -583 -1571 -549
rect 1571 -583 1667 -549
<< viali >>
rect -1409 447 -1375 481
rect -1217 447 -1183 481
rect -1025 447 -991 481
rect -833 447 -799 481
rect -641 447 -607 481
rect -449 447 -415 481
rect -257 447 -223 481
rect -65 447 -31 481
rect 127 447 161 481
rect 319 447 353 481
rect 511 447 545 481
rect 703 447 737 481
rect 895 447 929 481
rect 1087 447 1121 481
rect 1279 447 1313 481
rect 1471 447 1505 481
rect -1553 -388 -1519 388
rect -1457 -388 -1423 388
rect -1361 -388 -1327 388
rect -1265 -388 -1231 388
rect -1169 -388 -1135 388
rect -1073 -388 -1039 388
rect -977 -388 -943 388
rect -881 -388 -847 388
rect -785 -388 -751 388
rect -689 -388 -655 388
rect -593 -388 -559 388
rect -497 -388 -463 388
rect -401 -388 -367 388
rect -305 -388 -271 388
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect 271 -388 305 388
rect 367 -388 401 388
rect 463 -388 497 388
rect 559 -388 593 388
rect 655 -388 689 388
rect 751 -388 785 388
rect 847 -388 881 388
rect 943 -388 977 388
rect 1039 -388 1073 388
rect 1135 -388 1169 388
rect 1231 -388 1265 388
rect 1327 -388 1361 388
rect 1423 -388 1457 388
rect 1519 -388 1553 388
rect -1505 -481 -1471 -447
rect -1313 -481 -1279 -447
rect -1121 -481 -1087 -447
rect -929 -481 -895 -447
rect -737 -481 -703 -447
rect -545 -481 -511 -447
rect -353 -481 -319 -447
rect -161 -481 -127 -447
rect 31 -481 65 -447
rect 223 -481 257 -447
rect 415 -481 449 -447
rect 607 -481 641 -447
rect 799 -481 833 -447
rect 991 -481 1025 -447
rect 1183 -481 1217 -447
rect 1375 -481 1409 -447
<< metal1 >>
rect -1421 481 -1363 487
rect -1421 447 -1409 481
rect -1375 447 -1363 481
rect -1421 441 -1363 447
rect -1229 481 -1171 487
rect -1229 447 -1217 481
rect -1183 447 -1171 481
rect -1229 441 -1171 447
rect -1037 481 -979 487
rect -1037 447 -1025 481
rect -991 447 -979 481
rect -1037 441 -979 447
rect -845 481 -787 487
rect -845 447 -833 481
rect -799 447 -787 481
rect -845 441 -787 447
rect -653 481 -595 487
rect -653 447 -641 481
rect -607 447 -595 481
rect -653 441 -595 447
rect -461 481 -403 487
rect -461 447 -449 481
rect -415 447 -403 481
rect -461 441 -403 447
rect -269 481 -211 487
rect -269 447 -257 481
rect -223 447 -211 481
rect -269 441 -211 447
rect -77 481 -19 487
rect -77 447 -65 481
rect -31 447 -19 481
rect -77 441 -19 447
rect 115 481 173 487
rect 115 447 127 481
rect 161 447 173 481
rect 115 441 173 447
rect 307 481 365 487
rect 307 447 319 481
rect 353 447 365 481
rect 307 441 365 447
rect 499 481 557 487
rect 499 447 511 481
rect 545 447 557 481
rect 499 441 557 447
rect 691 481 749 487
rect 691 447 703 481
rect 737 447 749 481
rect 691 441 749 447
rect 883 481 941 487
rect 883 447 895 481
rect 929 447 941 481
rect 883 441 941 447
rect 1075 481 1133 487
rect 1075 447 1087 481
rect 1121 447 1133 481
rect 1075 441 1133 447
rect 1267 481 1325 487
rect 1267 447 1279 481
rect 1313 447 1325 481
rect 1267 441 1325 447
rect 1459 481 1517 487
rect 1459 447 1471 481
rect 1505 447 1517 481
rect 1459 441 1517 447
rect -1559 388 -1513 400
rect -1559 -388 -1553 388
rect -1519 -388 -1513 388
rect -1559 -400 -1513 -388
rect -1463 388 -1417 400
rect -1463 -388 -1457 388
rect -1423 -388 -1417 388
rect -1463 -400 -1417 -388
rect -1367 388 -1321 400
rect -1367 -388 -1361 388
rect -1327 -388 -1321 388
rect -1367 -400 -1321 -388
rect -1271 388 -1225 400
rect -1271 -388 -1265 388
rect -1231 -388 -1225 388
rect -1271 -400 -1225 -388
rect -1175 388 -1129 400
rect -1175 -388 -1169 388
rect -1135 -388 -1129 388
rect -1175 -400 -1129 -388
rect -1079 388 -1033 400
rect -1079 -388 -1073 388
rect -1039 -388 -1033 388
rect -1079 -400 -1033 -388
rect -983 388 -937 400
rect -983 -388 -977 388
rect -943 -388 -937 388
rect -983 -400 -937 -388
rect -887 388 -841 400
rect -887 -388 -881 388
rect -847 -388 -841 388
rect -887 -400 -841 -388
rect -791 388 -745 400
rect -791 -388 -785 388
rect -751 -388 -745 388
rect -791 -400 -745 -388
rect -695 388 -649 400
rect -695 -388 -689 388
rect -655 -388 -649 388
rect -695 -400 -649 -388
rect -599 388 -553 400
rect -599 -388 -593 388
rect -559 -388 -553 388
rect -599 -400 -553 -388
rect -503 388 -457 400
rect -503 -388 -497 388
rect -463 -388 -457 388
rect -503 -400 -457 -388
rect -407 388 -361 400
rect -407 -388 -401 388
rect -367 -388 -361 388
rect -407 -400 -361 -388
rect -311 388 -265 400
rect -311 -388 -305 388
rect -271 -388 -265 388
rect -311 -400 -265 -388
rect -215 388 -169 400
rect -215 -388 -209 388
rect -175 -388 -169 388
rect -215 -400 -169 -388
rect -119 388 -73 400
rect -119 -388 -113 388
rect -79 -388 -73 388
rect -119 -400 -73 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 73 388 119 400
rect 73 -388 79 388
rect 113 -388 119 388
rect 73 -400 119 -388
rect 169 388 215 400
rect 169 -388 175 388
rect 209 -388 215 388
rect 169 -400 215 -388
rect 265 388 311 400
rect 265 -388 271 388
rect 305 -388 311 388
rect 265 -400 311 -388
rect 361 388 407 400
rect 361 -388 367 388
rect 401 -388 407 388
rect 361 -400 407 -388
rect 457 388 503 400
rect 457 -388 463 388
rect 497 -388 503 388
rect 457 -400 503 -388
rect 553 388 599 400
rect 553 -388 559 388
rect 593 -388 599 388
rect 553 -400 599 -388
rect 649 388 695 400
rect 649 -388 655 388
rect 689 -388 695 388
rect 649 -400 695 -388
rect 745 388 791 400
rect 745 -388 751 388
rect 785 -388 791 388
rect 745 -400 791 -388
rect 841 388 887 400
rect 841 -388 847 388
rect 881 -388 887 388
rect 841 -400 887 -388
rect 937 388 983 400
rect 937 -388 943 388
rect 977 -388 983 388
rect 937 -400 983 -388
rect 1033 388 1079 400
rect 1033 -388 1039 388
rect 1073 -388 1079 388
rect 1033 -400 1079 -388
rect 1129 388 1175 400
rect 1129 -388 1135 388
rect 1169 -388 1175 388
rect 1129 -400 1175 -388
rect 1225 388 1271 400
rect 1225 -388 1231 388
rect 1265 -388 1271 388
rect 1225 -400 1271 -388
rect 1321 388 1367 400
rect 1321 -388 1327 388
rect 1361 -388 1367 388
rect 1321 -400 1367 -388
rect 1417 388 1463 400
rect 1417 -388 1423 388
rect 1457 -388 1463 388
rect 1417 -400 1463 -388
rect 1513 388 1559 400
rect 1513 -388 1519 388
rect 1553 -388 1559 388
rect 1513 -400 1559 -388
rect -1517 -447 -1459 -441
rect -1517 -481 -1505 -447
rect -1471 -481 -1459 -447
rect -1517 -487 -1459 -481
rect -1325 -447 -1267 -441
rect -1325 -481 -1313 -447
rect -1279 -481 -1267 -447
rect -1325 -487 -1267 -481
rect -1133 -447 -1075 -441
rect -1133 -481 -1121 -447
rect -1087 -481 -1075 -447
rect -1133 -487 -1075 -481
rect -941 -447 -883 -441
rect -941 -481 -929 -447
rect -895 -481 -883 -447
rect -941 -487 -883 -481
rect -749 -447 -691 -441
rect -749 -481 -737 -447
rect -703 -481 -691 -447
rect -749 -487 -691 -481
rect -557 -447 -499 -441
rect -557 -481 -545 -447
rect -511 -481 -499 -447
rect -557 -487 -499 -481
rect -365 -447 -307 -441
rect -365 -481 -353 -447
rect -319 -481 -307 -447
rect -365 -487 -307 -481
rect -173 -447 -115 -441
rect -173 -481 -161 -447
rect -127 -481 -115 -447
rect -173 -487 -115 -481
rect 19 -447 77 -441
rect 19 -481 31 -447
rect 65 -481 77 -447
rect 19 -487 77 -481
rect 211 -447 269 -441
rect 211 -481 223 -447
rect 257 -481 269 -447
rect 211 -487 269 -481
rect 403 -447 461 -441
rect 403 -481 415 -447
rect 449 -481 461 -447
rect 403 -487 461 -481
rect 595 -447 653 -441
rect 595 -481 607 -447
rect 641 -481 653 -447
rect 595 -487 653 -481
rect 787 -447 845 -441
rect 787 -481 799 -447
rect 833 -481 845 -447
rect 787 -487 845 -481
rect 979 -447 1037 -441
rect 979 -481 991 -447
rect 1025 -481 1037 -447
rect 979 -487 1037 -481
rect 1171 -447 1229 -441
rect 1171 -481 1183 -447
rect 1217 -481 1229 -447
rect 1171 -487 1229 -481
rect 1363 -447 1421 -441
rect 1363 -481 1375 -447
rect 1409 -481 1421 -447
rect 1363 -487 1421 -481
<< properties >>
string FIXED_BBOX -1650 -566 1650 566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 0.15 m 1 nf 32 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
