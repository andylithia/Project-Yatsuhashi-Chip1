** sch_path: /home/al/openmpw/Project-Yatsuhashi-Chip1/xschem/LNA5_with_output_buf_4_SP_captune.sch
**.subckt LNA5_with_output_buf_4_SP_captune
V1 VDD GND 1.8
V2 net3 GND dc 0.9 ac 1 portnum 1 z0 50
I0 VDDI Vref 1m
XM1 Vref Vref GNDI GNDI sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=2.5u l=0.15u m=1
XC7 Vref GNDI sky130_fd_pr__cap_mim_m3_1 W=20 L=30 MF=1 m=1
Ldeg5 net1 VDDI 2n m=1
R3 net1 VDD 3 m=1
Ldeg6 net2 GND 2n m=1
R4 net2 GNDI 3 m=1
C17 net7 net4 0.3p m=1
L2 VDDI net4 2.5n m=1
XC3 net12 GNDI sky130_fd_pr__cap_mim_m3_1 W=40 L=60 MF=8 m=8
C8 GNDI GND 1 m=1
C19 VDD VDDI 1 m=1
R2 net12 VDDI 5 m=1
C1 net5 net3 1n m=1
Ldeg1 net6 net5 2n m=1
L1 net10 vmid 0.7n m=1
Ldeg2 net9 net6 0.5n m=1
XC4 net13 GNDI sky130_fd_pr__cap_mim_m3_1 W=40 L=60 MF=8 m=8
R8 net13 VDDI 5 m=1
L4 net8 GNDI 1n m=1
V3 net7 GNDI dc 0.9 ac 1 portnum 2 z0 50
R7 g_top_ref VDDI 5k m=1
C5 GNDI g_top_ref 50f m=1
x3 VDDI net4 GNDI VDDI GNDI GNDI __UNCONNECTED_PIN__0 net11 net11 net10 vmid net8 Vref net9 GNDI
+ LNA_complete_2_wo_ind_PEX
**** begin user architecture code


.subckt sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=2.828e+12p pd=2.132e+07u as=4.242e+12p
+ ps=3.198e+07u w=5.05e+06u l=150000u
X1 SOURCE SUBSTRATE SUBSTRATE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.03e+12p
+ ps=2.14e+07u w=5.05e+06u l=150000u
X2 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X5 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends
.sp dec 1000 1e9 10e9 1
* .ac dec 1000 0.01e9 100e9
.control
run
display
let z11=50*(1+s_1_1)/(1-s_1_1)
let z22=50*(1+s_2_2)/(1-s_2_2)
let S11 = S_1_1
let S21 = S_2_1
let S12 = S_1_2
let S22 = S_2_2

* Stability
let delta=S11*S22-S12*S21
let K    = (1-mag(S11)^2-mag(S22)^2+mag(delta)^2)/(2*mag(S12*S21))
let mu   = (1-mag(S11)^2)/(mag(S22-conj(S11)*delta)+mag(S21*S12))
* plot real(z11) real(z22)
* plot imag(z11) imag(z22)
plot db(S_1_1) db(S_2_2) db(S_2_1)

plot db(K)
plot mag(delta)
plot db(mu)
plot NF NFmin
.endc


.lib /home/al/openmpw/pdk_1/sky130B/libs.tech/ngspice/sky130.lib.spice tt
* .include /home/al/openmpw/pdk_1/sky130B/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

**** end user architecture code
**.ends

* expanding   symbol:  LNA_complete_2_wo_ind_PEX.sym # of pins=15
** sym_path: /home/al/openmpw/Project-Yatsuhashi-Chip1/xschem/LNA_complete_2_wo_ind_PEX.sym
** sch_path: /home/al/openmpw/Project-Yatsuhashi-Chip1/xschem/LNA_complete_2_wo_ind_PEX.sch
.subckt LNA_complete_2_wo_ind_PEX VHI VOUT G4 G8 G2 G1 RFB_MID G_TOP BIAS_TOP S1 D1 SS BIAS_BOT VIN
+ VLO
*.iopin VHI
*.iopin VLO
*.iopin VOUT
*.iopin VIN
*.iopin SS
*.iopin D1
*.iopin S1
*.iopin BIAS_BOT
*.iopin BIAS_TOP
*.iopin G_TOP
*.iopin G2
*.iopin G8
*.iopin G4
*.iopin G1
*.iopin RFB_MID
**** begin user architecture code


* NGSPICE file created from flat3.ext - technology: sky130B
* lna_complete_2_wo_ind_flat_220831_2340
X0 S1.t23 G_TOP VOUT.t17 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X1 SS.t15 VIN D1.t11 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X2 VHI VLO sky130_fd_pr__cap_mim_m3_2 l=4.4e+07u w=5e+07u
X3 VOUT.t16 G_TOP S1.t22 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 SS.t14 VIN D1.t5 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X5 D1.t14 VIN SS.t13 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X6 VHI a_n6328_16092.t0 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2.5e+06u
X7 D1.t13 VIN SS.t12 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X8 S1.t21 G_TOP VOUT.t29 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X9 SS.t11 VIN D1.t4 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X10 D1.t8 VIN SS.t10 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X11 VLO VHI sky130_fd_pr__cap_mim_m3_1 l=4.4e+07u w=5e+07u
X12 BIAS_TOP VLO sky130_fd_pr__cap_mim_m3_2 l=7.5e+06u w=4.5e+06u
X13 SS.t9 VIN D1.t10 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X14 SS.t8 VIN D1.t0 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X15 BIAS_BOT VLO sky130_fd_pr__cap_mim_m3_2 l=1.15e+07u w=9.5e+06u
X16 S1.t20 G_TOP VOUT.t28 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X17 VOUT.t31 G_TOP S1.t19 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X18 D1.t12 VIN SS.t7 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X19 D1.t6 VIN SS.t6 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X20 VOUT.t30 G_TOP S1.t18 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X21 SS.t5 VIN D1.t15 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X22 VLO BIAS_TOP sky130_fd_pr__cap_mim_m3_1 l=7.5e+06u w=4.5e+06u
X23 a_n6328_16092.t2 G1 VOUT.t0 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X24 a_n5540_16092.t2 G4 VOUT.t6 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X25 S1.t17 G_TOP VOUT.t15 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
R0 RFB_MID VOUT sky130_fd_pr__res_generic_po w=330000u l=1.28e+07u
X26 D1.t3 VIN SS.t4 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X27 VOUT.t4 G2 a_n6722_16092.t2 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X28 VOUT.t2 G8 a_n5934_16092.t2 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X29 VOUT.t14 G_TOP S1.t16 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X30 VLO BIAS_BOT sky130_fd_pr__cap_mim_m3_1 l=1.15e+07u w=9.5e+06u
X31 S1.t15 G_TOP VOUT.t27 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X32 SS.t3 VIN D1.t7 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X33 D1.t2 VIN SS.t2 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X34 VOUT.t26 G_TOP S1.t14 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X35 VOUT.t11 G_TOP S1.t13 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X36 VOUT.t10 G_TOP S1.t12 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X37 S1.t11 G_TOP VOUT.t13 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X38 D1.t9 VIN SS.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X39 VHI a_n5934_16092.t0 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=8e+06u
X40 S1.t10 G_TOP VOUT.t12 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X41 VIN RFB_MID sky130_fd_pr__cap_mim_m3_2 l=2.05e+07u w=1.15e+07u
X42 VOUT.t1 G1 a_n6328_16092.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X43 VOUT.t7 G4 a_n5540_16092.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X44 VOUT.t21 G_TOP S1.t9 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X45 a_n5934_16092.t1 G8 VOUT.t3 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
R1 VHI BIAS_TOP sky130_fd_pr__res_generic_po w=330000u l=1.28e+07u
X46 S1.t8 G_TOP VOUT.t20 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
R2 BIAS_BOT VIN sky130_fd_pr__res_generic_po w=330000u l=2.068e+07u
X47 VOUT.t19 G_TOP S1.t7 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X48 RFB_MID VIN sky130_fd_pr__cap_mim_m3_1 l=2.05e+07u w=1.15e+07u
X49 VOUT.t18 G_TOP S1.t6 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X50 S1.t5 G_TOP VOUT.t25 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X51 VHI a_n5540_16092.t0 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=4e+06u
X52 S1.t4 G_TOP VOUT.t24 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X53 S1.t3 G_TOP VOUT.t23 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X54 VOUT.t22 G_TOP S1.t2 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X55 VOUT.t9 G_TOP S1.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X56 VHI a_n6722_16092.t0 sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=2.5e+06u
X57 S1.t0 G_TOP VOUT.t8 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X58 a_n6722_16092.t1 G2 VOUT.t5 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X59 SS.t0 VIN D1.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
C0 m5_n800_n3000# SS 3.92fF
C1 BIAS_BOT VIN 2.13fF
C2 RFB_MID VIN 40.06fF
C3 VIN D1 3.39fF
C4 VIN SS 14.77fF
C5 VOUT VHI 2.58fF
C6 D1 SS 26.96fF
C7 G_TOP VOUT 5.37fF
C8 m5_n800_n3000# VIN 1.17fF
C9 G_TOP S1 3.12fF
C10 S1 VOUT 41.75fF
R3 VOUT.n237 VOUT.n1279 9.305
R4 VOUT.n238 VOUT.n1159 9.305
R5 VOUT.n239 VOUT.n1259 9.305
R6 VOUT.n1281 VOUT.n1282 9.3
R7 VOUT.n155 VOUT.n1294 9.3
R8 VOUT.n27 VOUT.n1305 9.3
R9 VOUT.n141 VOUT.n1285 9.3
R10 VOUT.n1288 VOUT.n1287 9.3
R11 VOUT.n154 VOUT.n1291 9.3
R12 VOUT.n155 VOUT.n1293 9.3
R13 VOUT.n215 VOUT.n1297 9.3
R14 VOUT.n216 VOUT.n1300 9.3
R15 VOUT.n216 VOUT.n1299 9.3
R16 VOUT.n240 VOUT.n1303 9.3
R17 VOUT.n156 VOUT.n1278 9.3
R18 VOUT.n27 VOUT.n1306 9.3
R19 VOUT.n158 VOUT.n1174 9.3
R20 VOUT.n157 VOUT.n1171 9.3
R21 VOUT.n217 VOUT.n1177 9.3
R22 VOUT.n1168 VOUT.n1167 9.3
R23 VOUT.n138 VOUT.n1165 9.3
R24 VOUT.n1161 VOUT.n1162 9.3
R25 VOUT.n218 VOUT.n1180 9.3
R26 VOUT.n26 VOUT.n1186 9.3
R27 VOUT.n26 VOUT.n1185 9.3
R28 VOUT.n159 VOUT.n1158 9.3
R29 VOUT.n241 VOUT.n1183 9.3
R30 VOUT.n218 VOUT.n1179 9.3
R31 VOUT.n158 VOUT.n1173 9.3
R32 VOUT.n1261 VOUT.n1262 9.3
R33 VOUT.n1268 VOUT.n1267 9.3
R34 VOUT.n163 VOUT.n1255 9.3
R35 VOUT.n24 VOUT.n1244 9.3
R36 VOUT.n164 VOUT.n1258 9.3
R37 VOUT.n163 VOUT.n1256 9.3
R38 VOUT.n221 VOUT.n1253 9.3
R39 VOUT.n1239 VOUT.n1238 9.3
R40 VOUT.n1251 VOUT.n1250 9.3
R41 VOUT.n243 VOUT.n1242 9.3
R42 VOUT.n165 VOUT.n1232 9.3
R43 VOUT.n24 VOUT.n1245 9.3
R44 VOUT.n140 VOUT.n1265 9.3
R45 VOUT.n191 VOUT.n699 9.3
R46 VOUT.n115 VOUT.n687 9.3
R47 VOUT.n192 VOUT.n676 9.3
R48 VOUT.n222 VOUT.n680 9.3
R49 VOUT.n222 VOUT.n681 9.3
R50 VOUT.n684 VOUT.n683 9.3
R51 VOUT.n114 VOUT.n686 9.3
R52 VOUT.n115 VOUT.n689 9.3
R53 VOUT.n245 VOUT.n690 9.3
R54 VOUT.n244 VOUT.n691 9.3
R55 VOUT.n244 VOUT.n693 9.3
R56 VOUT.n23 VOUT.n695 9.3
R57 VOUT.n191 VOUT.n697 9.3
R58 VOUT.n64 VOUT.n701 9.3
R59 VOUT.n0 VOUT.n703 9.3
R60 VOUT.n52 VOUT.n704 9.3
R61 VOUT.n147 VOUT.n636 9.3
R62 VOUT.n50 VOUT.n658 9.3
R63 VOUT.n167 VOUT.n671 9.3
R64 VOUT.n166 VOUT.n670 9.3
R65 VOUT.n166 VOUT.n669 9.3
R66 VOUT.n66 VOUT.n650 9.3
R67 VOUT.n67 VOUT.n651 9.3
R68 VOUT.n65 VOUT.n654 9.3
R69 VOUT.n645 VOUT.n655 9.3
R70 VOUT.n50 VOUT.n659 9.3
R71 VOUT.n51 VOUT.n660 9.3
R72 VOUT.n675 VOUT.n674 9.3
R73 VOUT.n192 VOUT.n677 9.3
R74 VOUT.n193 VOUT.n626 9.3
R75 VOUT.n117 VOUT.n614 9.3
R76 VOUT.n194 VOUT.n603 9.3
R77 VOUT.n223 VOUT.n607 9.3
R78 VOUT.n223 VOUT.n608 9.3
R79 VOUT.n611 VOUT.n610 9.3
R80 VOUT.n116 VOUT.n613 9.3
R81 VOUT.n117 VOUT.n616 9.3
R82 VOUT.n247 VOUT.n617 9.3
R83 VOUT.n246 VOUT.n618 9.3
R84 VOUT.n246 VOUT.n620 9.3
R85 VOUT.n22 VOUT.n622 9.3
R86 VOUT.n193 VOUT.n624 9.3
R87 VOUT.n68 VOUT.n628 9.3
R88 VOUT.n1 VOUT.n630 9.3
R89 VOUT.n53 VOUT.n631 9.3
R90 VOUT.n146 VOUT.n563 9.3
R91 VOUT.n48 VOUT.n585 9.3
R92 VOUT.n169 VOUT.n598 9.3
R93 VOUT.n168 VOUT.n597 9.3
R94 VOUT.n168 VOUT.n596 9.3
R95 VOUT.n70 VOUT.n577 9.3
R96 VOUT.n71 VOUT.n578 9.3
R97 VOUT.n69 VOUT.n581 9.3
R98 VOUT.n572 VOUT.n582 9.3
R99 VOUT.n48 VOUT.n586 9.3
R100 VOUT.n49 VOUT.n587 9.3
R101 VOUT.n602 VOUT.n601 9.3
R102 VOUT.n194 VOUT.n604 9.3
R103 VOUT.n195 VOUT.n553 9.3
R104 VOUT.n119 VOUT.n541 9.3
R105 VOUT.n196 VOUT.n530 9.3
R106 VOUT.n224 VOUT.n534 9.3
R107 VOUT.n224 VOUT.n535 9.3
R108 VOUT.n538 VOUT.n537 9.3
R109 VOUT.n118 VOUT.n540 9.3
R110 VOUT.n119 VOUT.n543 9.3
R111 VOUT.n249 VOUT.n544 9.3
R112 VOUT.n248 VOUT.n545 9.3
R113 VOUT.n248 VOUT.n547 9.3
R114 VOUT.n21 VOUT.n549 9.3
R115 VOUT.n195 VOUT.n551 9.3
R116 VOUT.n72 VOUT.n555 9.3
R117 VOUT.n2 VOUT.n557 9.3
R118 VOUT.n54 VOUT.n558 9.3
R119 VOUT.n145 VOUT.n490 9.3
R120 VOUT.n46 VOUT.n512 9.3
R121 VOUT.n171 VOUT.n525 9.3
R122 VOUT.n170 VOUT.n524 9.3
R123 VOUT.n170 VOUT.n523 9.3
R124 VOUT.n74 VOUT.n504 9.3
R125 VOUT.n75 VOUT.n505 9.3
R126 VOUT.n73 VOUT.n508 9.3
R127 VOUT.n499 VOUT.n509 9.3
R128 VOUT.n46 VOUT.n513 9.3
R129 VOUT.n47 VOUT.n514 9.3
R130 VOUT.n529 VOUT.n528 9.3
R131 VOUT.n196 VOUT.n531 9.3
R132 VOUT.n197 VOUT.n480 9.3
R133 VOUT.n121 VOUT.n468 9.3
R134 VOUT.n198 VOUT.n457 9.3
R135 VOUT.n225 VOUT.n461 9.3
R136 VOUT.n225 VOUT.n462 9.3
R137 VOUT.n465 VOUT.n464 9.3
R138 VOUT.n120 VOUT.n467 9.3
R139 VOUT.n121 VOUT.n470 9.3
R140 VOUT.n251 VOUT.n471 9.3
R141 VOUT.n250 VOUT.n472 9.3
R142 VOUT.n250 VOUT.n474 9.3
R143 VOUT.n20 VOUT.n476 9.3
R144 VOUT.n197 VOUT.n478 9.3
R145 VOUT.n76 VOUT.n482 9.3
R146 VOUT.n3 VOUT.n484 9.3
R147 VOUT.n55 VOUT.n485 9.3
R148 VOUT.n144 VOUT.n417 9.3
R149 VOUT.n44 VOUT.n439 9.3
R150 VOUT.n173 VOUT.n452 9.3
R151 VOUT.n172 VOUT.n451 9.3
R152 VOUT.n172 VOUT.n450 9.3
R153 VOUT.n78 VOUT.n431 9.3
R154 VOUT.n79 VOUT.n432 9.3
R155 VOUT.n77 VOUT.n435 9.3
R156 VOUT.n426 VOUT.n436 9.3
R157 VOUT.n44 VOUT.n440 9.3
R158 VOUT.n45 VOUT.n441 9.3
R159 VOUT.n456 VOUT.n455 9.3
R160 VOUT.n198 VOUT.n458 9.3
R161 VOUT.n199 VOUT.n407 9.3
R162 VOUT.n123 VOUT.n395 9.3
R163 VOUT.n200 VOUT.n384 9.3
R164 VOUT.n226 VOUT.n388 9.3
R165 VOUT.n226 VOUT.n389 9.3
R166 VOUT.n392 VOUT.n391 9.3
R167 VOUT.n122 VOUT.n394 9.3
R168 VOUT.n123 VOUT.n397 9.3
R169 VOUT.n253 VOUT.n398 9.3
R170 VOUT.n252 VOUT.n399 9.3
R171 VOUT.n252 VOUT.n401 9.3
R172 VOUT.n19 VOUT.n403 9.3
R173 VOUT.n199 VOUT.n405 9.3
R174 VOUT.n80 VOUT.n409 9.3
R175 VOUT.n4 VOUT.n411 9.3
R176 VOUT.n56 VOUT.n412 9.3
R177 VOUT.n143 VOUT.n344 9.3
R178 VOUT.n42 VOUT.n366 9.3
R179 VOUT.n175 VOUT.n379 9.3
R180 VOUT.n174 VOUT.n378 9.3
R181 VOUT.n174 VOUT.n377 9.3
R182 VOUT.n82 VOUT.n358 9.3
R183 VOUT.n83 VOUT.n359 9.3
R184 VOUT.n81 VOUT.n362 9.3
R185 VOUT.n353 VOUT.n363 9.3
R186 VOUT.n42 VOUT.n367 9.3
R187 VOUT.n43 VOUT.n368 9.3
R188 VOUT.n383 VOUT.n382 9.3
R189 VOUT.n200 VOUT.n385 9.3
R190 VOUT.n201 VOUT.n334 9.3
R191 VOUT.n125 VOUT.n322 9.3
R192 VOUT.n202 VOUT.n311 9.3
R193 VOUT.n227 VOUT.n315 9.3
R194 VOUT.n227 VOUT.n316 9.3
R195 VOUT.n319 VOUT.n318 9.3
R196 VOUT.n124 VOUT.n321 9.3
R197 VOUT.n125 VOUT.n324 9.3
R198 VOUT.n255 VOUT.n325 9.3
R199 VOUT.n254 VOUT.n326 9.3
R200 VOUT.n254 VOUT.n328 9.3
R201 VOUT.n18 VOUT.n330 9.3
R202 VOUT.n201 VOUT.n332 9.3
R203 VOUT.n84 VOUT.n336 9.3
R204 VOUT.n5 VOUT.n338 9.3
R205 VOUT.n57 VOUT.n339 9.3
R206 VOUT.n142 VOUT.n271 9.3
R207 VOUT.n40 VOUT.n293 9.3
R208 VOUT.n177 VOUT.n306 9.3
R209 VOUT.n176 VOUT.n305 9.3
R210 VOUT.n176 VOUT.n304 9.3
R211 VOUT.n86 VOUT.n285 9.3
R212 VOUT.n87 VOUT.n286 9.3
R213 VOUT.n85 VOUT.n289 9.3
R214 VOUT.n280 VOUT.n290 9.3
R215 VOUT.n40 VOUT.n294 9.3
R216 VOUT.n41 VOUT.n295 9.3
R217 VOUT.n310 VOUT.n309 9.3
R218 VOUT.n202 VOUT.n312 9.3
R219 VOUT.n203 VOUT.n1142 9.3
R220 VOUT.n127 VOUT.n1130 9.3
R221 VOUT.n204 VOUT.n1119 9.3
R222 VOUT.n228 VOUT.n1123 9.3
R223 VOUT.n228 VOUT.n1124 9.3
R224 VOUT.n1127 VOUT.n1126 9.3
R225 VOUT.n126 VOUT.n1129 9.3
R226 VOUT.n127 VOUT.n1132 9.3
R227 VOUT.n257 VOUT.n1133 9.3
R228 VOUT.n256 VOUT.n1134 9.3
R229 VOUT.n256 VOUT.n1136 9.3
R230 VOUT.n17 VOUT.n1138 9.3
R231 VOUT.n203 VOUT.n1140 9.3
R232 VOUT.n88 VOUT.n1144 9.3
R233 VOUT.n6 VOUT.n1146 9.3
R234 VOUT.n58 VOUT.n1147 9.3
R235 VOUT.n153 VOUT.n1079 9.3
R236 VOUT.n38 VOUT.n1101 9.3
R237 VOUT.n179 VOUT.n1114 9.3
R238 VOUT.n178 VOUT.n1113 9.3
R239 VOUT.n178 VOUT.n1112 9.3
R240 VOUT.n90 VOUT.n1093 9.3
R241 VOUT.n91 VOUT.n1094 9.3
R242 VOUT.n89 VOUT.n1097 9.3
R243 VOUT.n1088 VOUT.n1098 9.3
R244 VOUT.n38 VOUT.n1102 9.3
R245 VOUT.n39 VOUT.n1103 9.3
R246 VOUT.n1118 VOUT.n1117 9.3
R247 VOUT.n204 VOUT.n1120 9.3
R248 VOUT.n205 VOUT.n1069 9.3
R249 VOUT.n129 VOUT.n1057 9.3
R250 VOUT.n206 VOUT.n1046 9.3
R251 VOUT.n229 VOUT.n1050 9.3
R252 VOUT.n229 VOUT.n1051 9.3
R253 VOUT.n1054 VOUT.n1053 9.3
R254 VOUT.n128 VOUT.n1056 9.3
R255 VOUT.n129 VOUT.n1059 9.3
R256 VOUT.n259 VOUT.n1060 9.3
R257 VOUT.n258 VOUT.n1061 9.3
R258 VOUT.n258 VOUT.n1063 9.3
R259 VOUT.n16 VOUT.n1065 9.3
R260 VOUT.n205 VOUT.n1067 9.3
R261 VOUT.n92 VOUT.n1071 9.3
R262 VOUT.n7 VOUT.n1073 9.3
R263 VOUT.n59 VOUT.n1074 9.3
R264 VOUT.n152 VOUT.n1006 9.3
R265 VOUT.n36 VOUT.n1028 9.3
R266 VOUT.n181 VOUT.n1041 9.3
R267 VOUT.n180 VOUT.n1040 9.3
R268 VOUT.n180 VOUT.n1039 9.3
R269 VOUT.n94 VOUT.n1020 9.3
R270 VOUT.n95 VOUT.n1021 9.3
R271 VOUT.n93 VOUT.n1024 9.3
R272 VOUT.n1015 VOUT.n1025 9.3
R273 VOUT.n36 VOUT.n1029 9.3
R274 VOUT.n37 VOUT.n1030 9.3
R275 VOUT.n1045 VOUT.n1044 9.3
R276 VOUT.n206 VOUT.n1047 9.3
R277 VOUT.n207 VOUT.n996 9.3
R278 VOUT.n131 VOUT.n984 9.3
R279 VOUT.n208 VOUT.n973 9.3
R280 VOUT.n230 VOUT.n977 9.3
R281 VOUT.n230 VOUT.n978 9.3
R282 VOUT.n981 VOUT.n980 9.3
R283 VOUT.n130 VOUT.n983 9.3
R284 VOUT.n131 VOUT.n986 9.3
R285 VOUT.n261 VOUT.n987 9.3
R286 VOUT.n260 VOUT.n988 9.3
R287 VOUT.n260 VOUT.n990 9.3
R288 VOUT.n15 VOUT.n992 9.3
R289 VOUT.n207 VOUT.n994 9.3
R290 VOUT.n96 VOUT.n998 9.3
R291 VOUT.n8 VOUT.n1000 9.3
R292 VOUT.n60 VOUT.n1001 9.3
R293 VOUT.n151 VOUT.n933 9.3
R294 VOUT.n34 VOUT.n955 9.3
R295 VOUT.n183 VOUT.n968 9.3
R296 VOUT.n182 VOUT.n967 9.3
R297 VOUT.n182 VOUT.n966 9.3
R298 VOUT.n98 VOUT.n947 9.3
R299 VOUT.n99 VOUT.n948 9.3
R300 VOUT.n97 VOUT.n951 9.3
R301 VOUT.n942 VOUT.n952 9.3
R302 VOUT.n34 VOUT.n956 9.3
R303 VOUT.n35 VOUT.n957 9.3
R304 VOUT.n972 VOUT.n971 9.3
R305 VOUT.n208 VOUT.n974 9.3
R306 VOUT.n209 VOUT.n774 9.3
R307 VOUT.n133 VOUT.n762 9.3
R308 VOUT.n210 VOUT.n751 9.3
R309 VOUT.n231 VOUT.n755 9.3
R310 VOUT.n231 VOUT.n756 9.3
R311 VOUT.n759 VOUT.n758 9.3
R312 VOUT.n132 VOUT.n761 9.3
R313 VOUT.n133 VOUT.n764 9.3
R314 VOUT.n263 VOUT.n765 9.3
R315 VOUT.n262 VOUT.n766 9.3
R316 VOUT.n262 VOUT.n768 9.3
R317 VOUT.n14 VOUT.n770 9.3
R318 VOUT.n209 VOUT.n772 9.3
R319 VOUT.n100 VOUT.n776 9.3
R320 VOUT.n9 VOUT.n778 9.3
R321 VOUT.n61 VOUT.n779 9.3
R322 VOUT.n148 VOUT.n711 9.3
R323 VOUT.n32 VOUT.n733 9.3
R324 VOUT.n185 VOUT.n746 9.3
R325 VOUT.n184 VOUT.n745 9.3
R326 VOUT.n184 VOUT.n744 9.3
R327 VOUT.n102 VOUT.n725 9.3
R328 VOUT.n103 VOUT.n726 9.3
R329 VOUT.n101 VOUT.n729 9.3
R330 VOUT.n720 VOUT.n730 9.3
R331 VOUT.n32 VOUT.n734 9.3
R332 VOUT.n33 VOUT.n735 9.3
R333 VOUT.n750 VOUT.n749 9.3
R334 VOUT.n210 VOUT.n752 9.3
R335 VOUT.n211 VOUT.n847 9.3
R336 VOUT.n135 VOUT.n835 9.3
R337 VOUT.n212 VOUT.n824 9.3
R338 VOUT.n232 VOUT.n828 9.3
R339 VOUT.n232 VOUT.n829 9.3
R340 VOUT.n832 VOUT.n831 9.3
R341 VOUT.n134 VOUT.n834 9.3
R342 VOUT.n135 VOUT.n837 9.3
R343 VOUT.n265 VOUT.n838 9.3
R344 VOUT.n264 VOUT.n839 9.3
R345 VOUT.n264 VOUT.n841 9.3
R346 VOUT.n13 VOUT.n843 9.3
R347 VOUT.n211 VOUT.n845 9.3
R348 VOUT.n104 VOUT.n849 9.3
R349 VOUT.n10 VOUT.n851 9.3
R350 VOUT.n62 VOUT.n852 9.3
R351 VOUT.n149 VOUT.n784 9.3
R352 VOUT.n30 VOUT.n806 9.3
R353 VOUT.n187 VOUT.n819 9.3
R354 VOUT.n186 VOUT.n818 9.3
R355 VOUT.n186 VOUT.n817 9.3
R356 VOUT.n106 VOUT.n798 9.3
R357 VOUT.n107 VOUT.n799 9.3
R358 VOUT.n105 VOUT.n802 9.3
R359 VOUT.n793 VOUT.n803 9.3
R360 VOUT.n30 VOUT.n807 9.3
R361 VOUT.n31 VOUT.n808 9.3
R362 VOUT.n823 VOUT.n822 9.3
R363 VOUT.n212 VOUT.n825 9.3
R364 VOUT.n213 VOUT.n920 9.3
R365 VOUT.n137 VOUT.n908 9.3
R366 VOUT.n214 VOUT.n897 9.3
R367 VOUT.n233 VOUT.n901 9.3
R368 VOUT.n233 VOUT.n902 9.3
R369 VOUT.n905 VOUT.n904 9.3
R370 VOUT.n136 VOUT.n907 9.3
R371 VOUT.n137 VOUT.n910 9.3
R372 VOUT.n267 VOUT.n911 9.3
R373 VOUT.n266 VOUT.n912 9.3
R374 VOUT.n266 VOUT.n914 9.3
R375 VOUT.n12 VOUT.n916 9.3
R376 VOUT.n213 VOUT.n918 9.3
R377 VOUT.n108 VOUT.n922 9.3
R378 VOUT.n11 VOUT.n924 9.3
R379 VOUT.n63 VOUT.n925 9.3
R380 VOUT.n150 VOUT.n857 9.3
R381 VOUT.n28 VOUT.n879 9.3
R382 VOUT.n189 VOUT.n892 9.3
R383 VOUT.n188 VOUT.n891 9.3
R384 VOUT.n188 VOUT.n890 9.3
R385 VOUT.n110 VOUT.n871 9.3
R386 VOUT.n111 VOUT.n872 9.3
R387 VOUT.n109 VOUT.n875 9.3
R388 VOUT.n866 VOUT.n876 9.3
R389 VOUT.n28 VOUT.n880 9.3
R390 VOUT.n29 VOUT.n881 9.3
R391 VOUT.n896 VOUT.n895 9.3
R392 VOUT.n214 VOUT.n898 9.3
R393 VOUT.n162 VOUT.n1226 9.3
R394 VOUT.n1193 VOUT.n1192 9.3
R395 VOUT.n25 VOUT.n1199 9.3
R396 VOUT.n25 VOUT.n1198 9.3
R397 VOUT.n160 VOUT.n1208 9.3
R398 VOUT.n160 VOUT.n1209 9.3
R399 VOUT.n1222 VOUT.n1221 9.3
R400 VOUT.n1215 VOUT.n1216 9.3
R401 VOUT.n1203 VOUT.n1202 9.3
R402 VOUT.n220 VOUT.n1206 9.3
R403 VOUT.n242 VOUT.n1196 9.3
R404 VOUT.n161 VOUT.n1212 9.3
R405 VOUT.n139 VOUT.n1219 9.3
R406 VOUT.n219 VOUT.n1213 9.3
R407 VOUT.n142 VOUT.n272 9
R408 VOUT.n5 VOUT.n273 9
R409 VOUT.n18 VOUT.n331 9
R410 VOUT.n255 VOUT.n274 9
R411 VOUT.n124 VOUT.n320 9
R412 VOUT.n314 VOUT.n276 9
R413 VOUT.n86 VOUT.n282 9
R414 VOUT.n85 VOUT.n281 9
R415 VOUT.n41 VOUT.n279 9
R416 VOUT.n177 VOUT.n307 9
R417 VOUT.n313 VOUT.n277 9
R418 VOUT.n143 VOUT.n345 9
R419 VOUT.n4 VOUT.n346 9
R420 VOUT.n19 VOUT.n404 9
R421 VOUT.n253 VOUT.n347 9
R422 VOUT.n122 VOUT.n393 9
R423 VOUT.n387 VOUT.n349 9
R424 VOUT.n82 VOUT.n355 9
R425 VOUT.n81 VOUT.n354 9
R426 VOUT.n43 VOUT.n352 9
R427 VOUT.n175 VOUT.n380 9
R428 VOUT.n386 VOUT.n350 9
R429 VOUT.n144 VOUT.n418 9
R430 VOUT.n3 VOUT.n419 9
R431 VOUT.n20 VOUT.n477 9
R432 VOUT.n251 VOUT.n420 9
R433 VOUT.n120 VOUT.n466 9
R434 VOUT.n460 VOUT.n422 9
R435 VOUT.n78 VOUT.n428 9
R436 VOUT.n77 VOUT.n427 9
R437 VOUT.n45 VOUT.n425 9
R438 VOUT.n173 VOUT.n453 9
R439 VOUT.n459 VOUT.n423 9
R440 VOUT.n145 VOUT.n491 9
R441 VOUT.n2 VOUT.n492 9
R442 VOUT.n21 VOUT.n550 9
R443 VOUT.n249 VOUT.n493 9
R444 VOUT.n118 VOUT.n539 9
R445 VOUT.n533 VOUT.n495 9
R446 VOUT.n74 VOUT.n501 9
R447 VOUT.n73 VOUT.n500 9
R448 VOUT.n47 VOUT.n498 9
R449 VOUT.n171 VOUT.n526 9
R450 VOUT.n532 VOUT.n496 9
R451 VOUT.n146 VOUT.n564 9
R452 VOUT.n1 VOUT.n565 9
R453 VOUT.n22 VOUT.n623 9
R454 VOUT.n247 VOUT.n566 9
R455 VOUT.n116 VOUT.n612 9
R456 VOUT.n606 VOUT.n568 9
R457 VOUT.n70 VOUT.n574 9
R458 VOUT.n69 VOUT.n573 9
R459 VOUT.n49 VOUT.n571 9
R460 VOUT.n169 VOUT.n599 9
R461 VOUT.n605 VOUT.n569 9
R462 VOUT.n147 VOUT.n637 9
R463 VOUT.n0 VOUT.n638 9
R464 VOUT.n23 VOUT.n696 9
R465 VOUT.n245 VOUT.n639 9
R466 VOUT.n114 VOUT.n685 9
R467 VOUT.n679 VOUT.n641 9
R468 VOUT.n66 VOUT.n647 9
R469 VOUT.n65 VOUT.n646 9
R470 VOUT.n51 VOUT.n644 9
R471 VOUT.n167 VOUT.n672 9
R472 VOUT.n678 VOUT.n642 9
R473 VOUT.n153 VOUT.n1080 9
R474 VOUT.n6 VOUT.n1081 9
R475 VOUT.n17 VOUT.n1139 9
R476 VOUT.n257 VOUT.n1082 9
R477 VOUT.n126 VOUT.n1128 9
R478 VOUT.n1122 VOUT.n1084 9
R479 VOUT.n90 VOUT.n1090 9
R480 VOUT.n89 VOUT.n1089 9
R481 VOUT.n39 VOUT.n1087 9
R482 VOUT.n179 VOUT.n1115 9
R483 VOUT.n1121 VOUT.n1085 9
R484 VOUT.n152 VOUT.n1007 9
R485 VOUT.n7 VOUT.n1008 9
R486 VOUT.n16 VOUT.n1066 9
R487 VOUT.n259 VOUT.n1009 9
R488 VOUT.n128 VOUT.n1055 9
R489 VOUT.n1049 VOUT.n1011 9
R490 VOUT.n94 VOUT.n1017 9
R491 VOUT.n93 VOUT.n1016 9
R492 VOUT.n37 VOUT.n1014 9
R493 VOUT.n181 VOUT.n1042 9
R494 VOUT.n1048 VOUT.n1012 9
R495 VOUT.n151 VOUT.n934 9
R496 VOUT.n8 VOUT.n935 9
R497 VOUT.n15 VOUT.n993 9
R498 VOUT.n261 VOUT.n936 9
R499 VOUT.n130 VOUT.n982 9
R500 VOUT.n976 VOUT.n938 9
R501 VOUT.n98 VOUT.n944 9
R502 VOUT.n97 VOUT.n943 9
R503 VOUT.n35 VOUT.n941 9
R504 VOUT.n183 VOUT.n969 9
R505 VOUT.n975 VOUT.n939 9
R506 VOUT.n148 VOUT.n712 9
R507 VOUT.n9 VOUT.n713 9
R508 VOUT.n14 VOUT.n771 9
R509 VOUT.n263 VOUT.n714 9
R510 VOUT.n132 VOUT.n760 9
R511 VOUT.n754 VOUT.n716 9
R512 VOUT.n102 VOUT.n722 9
R513 VOUT.n101 VOUT.n721 9
R514 VOUT.n33 VOUT.n719 9
R515 VOUT.n185 VOUT.n747 9
R516 VOUT.n753 VOUT.n717 9
R517 VOUT.n149 VOUT.n785 9
R518 VOUT.n10 VOUT.n786 9
R519 VOUT.n13 VOUT.n844 9
R520 VOUT.n265 VOUT.n787 9
R521 VOUT.n134 VOUT.n833 9
R522 VOUT.n827 VOUT.n789 9
R523 VOUT.n106 VOUT.n795 9
R524 VOUT.n105 VOUT.n794 9
R525 VOUT.n31 VOUT.n792 9
R526 VOUT.n187 VOUT.n820 9
R527 VOUT.n826 VOUT.n790 9
R528 VOUT.n150 VOUT.n858 9
R529 VOUT.n11 VOUT.n859 9
R530 VOUT.n12 VOUT.n917 9
R531 VOUT.n267 VOUT.n860 9
R532 VOUT.n136 VOUT.n906 9
R533 VOUT.n900 VOUT.n862 9
R534 VOUT.n110 VOUT.n868 9
R535 VOUT.n109 VOUT.n867 9
R536 VOUT.n29 VOUT.n865 9
R537 VOUT.n189 VOUT.n893 9
R538 VOUT.n899 VOUT.n863 9
R539 VOUT.n159 VOUT.n1154 9
R540 VOUT.n156 VOUT.n1274 9
R541 VOUT.n138 VOUT.n1166 9
R542 VOUT.n238 VOUT.n1160 9
R543 VOUT.n141 VOUT.n1286 9
R544 VOUT.n154 VOUT.n1292 9
R545 VOUT.n215 VOUT.n1298 9
R546 VOUT.n165 VOUT.n1233 9
R547 VOUT.n164 VOUT.n1248 9
R548 VOUT.n221 VOUT.n1249 9
R549 VOUT.n24 VOUT.n1246 9
R550 VOUT.n243 VOUT.n1243 9
R551 VOUT.n140 VOUT.n1266 9
R552 VOUT.n26 VOUT.n1187 9
R553 VOUT.n27 VOUT.n1307 9
R554 VOUT.n240 VOUT.n1304 9
R555 VOUT.n241 VOUT.n1184 9
R556 VOUT.n217 VOUT.n1178 9
R557 VOUT.n237 VOUT.n1280 9
R558 VOUT.n157 VOUT.n1172 9
R559 VOUT.n239 VOUT.n1260 9
R560 VOUT.n219 VOUT.n1214 9
R561 VOUT.n139 VOUT.n1220 9
R562 VOUT.n161 VOUT.n1210 9
R563 VOUT.n162 VOUT.n1227 9
R564 VOUT.n25 VOUT.n1200 9
R565 VOUT.n242 VOUT.n1197 9
R566 VOUT.n220 VOUT.n1204 9
R567 VOUT.n641 VOUT.n640 8.282
R568 VOUT.n568 VOUT.n567 8.282
R569 VOUT.n495 VOUT.n494 8.282
R570 VOUT.n422 VOUT.n421 8.282
R571 VOUT.n349 VOUT.n348 8.282
R572 VOUT.n276 VOUT.n275 8.282
R573 VOUT.n1084 VOUT.n1083 8.282
R574 VOUT.n1011 VOUT.n1010 8.282
R575 VOUT.n938 VOUT.n937 8.282
R576 VOUT.n716 VOUT.n715 8.282
R577 VOUT.n789 VOUT.n788 8.282
R578 VOUT.n862 VOUT.n861 8.282
R579 VOUT.n635 VOUT.n634 7.853
R580 VOUT.n562 VOUT.n561 7.853
R581 VOUT.n489 VOUT.n488 7.853
R582 VOUT.n416 VOUT.n415 7.853
R583 VOUT.n343 VOUT.n342 7.853
R584 VOUT.n270 VOUT.n269 7.853
R585 VOUT.n1078 VOUT.n1077 7.853
R586 VOUT.n1005 VOUT.n1004 7.853
R587 VOUT.n932 VOUT.n931 7.853
R588 VOUT.n710 VOUT.n709 7.853
R589 VOUT.n783 VOUT.n782 7.853
R590 VOUT.n856 VOUT.n855 7.853
R591 VOUT.n649 VOUT.n648 7.851
R592 VOUT.n576 VOUT.n575 7.851
R593 VOUT.n503 VOUT.n502 7.851
R594 VOUT.n430 VOUT.n429 7.851
R595 VOUT.n357 VOUT.n356 7.851
R596 VOUT.n284 VOUT.n283 7.851
R597 VOUT.n1092 VOUT.n1091 7.851
R598 VOUT.n1019 VOUT.n1018 7.851
R599 VOUT.n946 VOUT.n945 7.851
R600 VOUT.n724 VOUT.n723 7.851
R601 VOUT.n797 VOUT.n796 7.851
R602 VOUT.n870 VOUT.n869 7.851
R603 VOUT.n664 VOUT.n663 4.65
R604 VOUT.n591 VOUT.n590 4.65
R605 VOUT.n518 VOUT.n517 4.65
R606 VOUT.n445 VOUT.n444 4.65
R607 VOUT.n372 VOUT.n371 4.65
R608 VOUT.n299 VOUT.n298 4.65
R609 VOUT.n1107 VOUT.n1106 4.65
R610 VOUT.n1034 VOUT.n1033 4.65
R611 VOUT.n961 VOUT.n960 4.65
R612 VOUT.n739 VOUT.n738 4.65
R613 VOUT.n812 VOUT.n811 4.65
R614 VOUT.n885 VOUT.n884 4.65
R615 VOUT.n1201 VOUT.n1191 4.61
R616 VOUT.n1247 VOUT.n1237 4.61
R617 VOUT.n300 VOUT.n278 4.574
R618 VOUT.n373 VOUT.n351 4.574
R619 VOUT.n446 VOUT.n424 4.574
R620 VOUT.n519 VOUT.n497 4.574
R621 VOUT.n592 VOUT.n570 4.574
R622 VOUT.n665 VOUT.n643 4.574
R623 VOUT.n1108 VOUT.n1086 4.574
R624 VOUT.n1035 VOUT.n1013 4.574
R625 VOUT.n962 VOUT.n940 4.574
R626 VOUT.n740 VOUT.n718 4.574
R627 VOUT.n813 VOUT.n791 4.574
R628 VOUT.n886 VOUT.n864 4.574
R629 VOUT.n1153 VOUT.n1152 4.574
R630 VOUT.n1273 VOUT.n1272 4.574
R631 VOUT.n1272 VOUT.n1271 3.388
R632 VOUT.n1152 VOUT.n1151 3.388
R633 VOUT.n1237 VOUT.n1236 3.388
R634 VOUT.n1191 VOUT.n1190 3.388
R635 VOUT.n1275 VOUT.t6 3.326
R636 VOUT.n1275 VOUT.t7 3.326
R637 VOUT.n1155 VOUT.t3 3.326
R638 VOUT.n1155 VOUT.t2 3.326
R639 VOUT.n1230 VOUT.t5 3.326
R640 VOUT.n1230 VOUT.t4 3.326
R641 VOUT.n633 VOUT.t20 3.326
R642 VOUT.n633 VOUT.t9 3.326
R643 VOUT.n560 VOUT.t25 3.326
R644 VOUT.n560 VOUT.t21 3.326
R645 VOUT.n487 VOUT.t23 3.326
R646 VOUT.n487 VOUT.t19 3.326
R647 VOUT.n414 VOUT.t8 3.326
R648 VOUT.n414 VOUT.t22 3.326
R649 VOUT.n341 VOUT.t12 3.326
R650 VOUT.n341 VOUT.t18 3.326
R651 VOUT.n268 VOUT.t24 3.326
R652 VOUT.n268 VOUT.t11 3.326
R653 VOUT.n1076 VOUT.t17 3.326
R654 VOUT.n1076 VOUT.t16 3.326
R655 VOUT.n1003 VOUT.t28 3.326
R656 VOUT.n1003 VOUT.t10 3.326
R657 VOUT.n930 VOUT.t29 3.326
R658 VOUT.n930 VOUT.t14 3.326
R659 VOUT.n708 VOUT.t15 3.326
R660 VOUT.n708 VOUT.t31 3.326
R661 VOUT.n781 VOUT.t13 3.326
R662 VOUT.n781 VOUT.t26 3.326
R663 VOUT.n854 VOUT.t27 3.326
R664 VOUT.n854 VOUT.t30 3.326
R665 VOUT.n1224 VOUT.t0 3.326
R666 VOUT.n1224 VOUT.t1 3.326
R667 VOUT.n699 VOUT.n698 3.191
R668 VOUT.n626 VOUT.n625 3.191
R669 VOUT.n553 VOUT.n552 3.191
R670 VOUT.n480 VOUT.n479 3.191
R671 VOUT.n407 VOUT.n406 3.191
R672 VOUT.n334 VOUT.n333 3.191
R673 VOUT.n1142 VOUT.n1141 3.191
R674 VOUT.n1069 VOUT.n1068 3.191
R675 VOUT.n996 VOUT.n995 3.191
R676 VOUT.n774 VOUT.n773 3.191
R677 VOUT.n847 VOUT.n846 3.191
R678 VOUT.n920 VOUT.n919 3.191
R679 VOUT.n340 VOUT.n142 3.055
R680 VOUT.n413 VOUT.n143 3.055
R681 VOUT.n486 VOUT.n144 3.055
R682 VOUT.n559 VOUT.n145 3.055
R683 VOUT.n632 VOUT.n146 3.055
R684 VOUT.n705 VOUT.n147 3.055
R685 VOUT.n1148 VOUT.n153 3.055
R686 VOUT.n1075 VOUT.n152 3.055
R687 VOUT.n1002 VOUT.n151 3.055
R688 VOUT.n780 VOUT.n148 3.055
R689 VOUT.n853 VOUT.n149 3.055
R690 VOUT.n926 VOUT.n150 3.055
R691 VOUT.n1229 VOUT.n1247 2.989
R692 VOUT.n234 VOUT.n1201 2.989
R693 VOUT.n1229 VOUT.n1234 2.987
R694 VOUT.n234 VOUT.n1228 2.987
R695 VOUT.n1229 VOUT.n1269 2.979
R696 VOUT.n234 VOUT.n1223 2.979
R697 VOUT.n658 VOUT.n657 2.814
R698 VOUT.n585 VOUT.n584 2.814
R699 VOUT.n512 VOUT.n511 2.814
R700 VOUT.n439 VOUT.n438 2.814
R701 VOUT.n366 VOUT.n365 2.814
R702 VOUT.n293 VOUT.n292 2.814
R703 VOUT.n1101 VOUT.n1100 2.814
R704 VOUT.n1028 VOUT.n1027 2.814
R705 VOUT.n955 VOUT.n954 2.814
R706 VOUT.n733 VOUT.n732 2.814
R707 VOUT.n806 VOUT.n805 2.814
R708 VOUT.n879 VOUT.n878 2.814
R709 VOUT.n236 VOUT.n1308 2.231
R710 VOUT.n235 VOUT.n1188 2.231
R711 VOUT.n634 VOUT.n633 2.082
R712 VOUT.n561 VOUT.n560 2.082
R713 VOUT.n488 VOUT.n487 2.082
R714 VOUT.n415 VOUT.n414 2.082
R715 VOUT.n342 VOUT.n341 2.082
R716 VOUT.n269 VOUT.n268 2.082
R717 VOUT.n1077 VOUT.n1076 2.082
R718 VOUT.n1004 VOUT.n1003 2.082
R719 VOUT.n931 VOUT.n930 2.082
R720 VOUT.n709 VOUT.n708 2.082
R721 VOUT.n782 VOUT.n781 2.082
R722 VOUT.n855 VOUT.n854 2.082
R723 VOUT.n1231 VOUT.n1230 1.155
R724 VOUT.n1225 VOUT.n1224 1.155
R725 VOUT.n1276 VOUT.n1275 1.155
R726 VOUT.n1156 VOUT.n1155 1.155
R727 VOUT.n928 VOUT.n927 0.926
R728 VOUT.n1234 VOUT.n1231 0.921
R729 VOUT.n1157 VOUT.n1156 0.921
R730 VOUT.n1228 VOUT.n1225 0.921
R731 VOUT.n1277 VOUT.n1276 0.903
R732 VOUT.n683 VOUT.n682 0.536
R733 VOUT.n674 VOUT.n673 0.536
R734 VOUT.n610 VOUT.n609 0.536
R735 VOUT.n601 VOUT.n600 0.536
R736 VOUT.n537 VOUT.n536 0.536
R737 VOUT.n528 VOUT.n527 0.536
R738 VOUT.n464 VOUT.n463 0.536
R739 VOUT.n455 VOUT.n454 0.536
R740 VOUT.n391 VOUT.n390 0.536
R741 VOUT.n382 VOUT.n381 0.536
R742 VOUT.n318 VOUT.n317 0.536
R743 VOUT.n309 VOUT.n308 0.536
R744 VOUT.n1126 VOUT.n1125 0.536
R745 VOUT.n1117 VOUT.n1116 0.536
R746 VOUT.n1053 VOUT.n1052 0.536
R747 VOUT.n1044 VOUT.n1043 0.536
R748 VOUT.n980 VOUT.n979 0.536
R749 VOUT.n971 VOUT.n970 0.536
R750 VOUT.n758 VOUT.n757 0.536
R751 VOUT.n749 VOUT.n748 0.536
R752 VOUT.n831 VOUT.n830 0.536
R753 VOUT.n822 VOUT.n821 0.536
R754 VOUT.n904 VOUT.n903 0.536
R755 VOUT.n895 VOUT.n894 0.536
R756 VOUT.n1272 VOUT.n1270 0.506
R757 VOUT.n1152 VOUT.n1150 0.506
R758 VOUT.n1237 VOUT.n1235 0.506
R759 VOUT.n689 VOUT.n688 0.506
R760 VOUT.n669 VOUT.n668 0.506
R761 VOUT.n616 VOUT.n615 0.506
R762 VOUT.n596 VOUT.n595 0.506
R763 VOUT.n543 VOUT.n542 0.506
R764 VOUT.n523 VOUT.n522 0.506
R765 VOUT.n470 VOUT.n469 0.506
R766 VOUT.n450 VOUT.n449 0.506
R767 VOUT.n397 VOUT.n396 0.506
R768 VOUT.n377 VOUT.n376 0.506
R769 VOUT.n324 VOUT.n323 0.506
R770 VOUT.n304 VOUT.n303 0.506
R771 VOUT.n1132 VOUT.n1131 0.506
R772 VOUT.n1112 VOUT.n1111 0.506
R773 VOUT.n1059 VOUT.n1058 0.506
R774 VOUT.n1039 VOUT.n1038 0.506
R775 VOUT.n986 VOUT.n985 0.506
R776 VOUT.n966 VOUT.n965 0.506
R777 VOUT.n764 VOUT.n763 0.506
R778 VOUT.n744 VOUT.n743 0.506
R779 VOUT.n837 VOUT.n836 0.506
R780 VOUT.n817 VOUT.n816 0.506
R781 VOUT.n910 VOUT.n909 0.506
R782 VOUT.n890 VOUT.n889 0.506
R783 VOUT.n1191 VOUT.n1189 0.506
R784 VOUT.n1303 VOUT.n1302 0.476
R785 VOUT.n1183 VOUT.n1182 0.476
R786 VOUT.n1242 VOUT.n1241 0.476
R787 VOUT.n693 VOUT.n692 0.476
R788 VOUT.n663 VOUT.n662 0.476
R789 VOUT.n620 VOUT.n619 0.476
R790 VOUT.n590 VOUT.n589 0.476
R791 VOUT.n547 VOUT.n546 0.476
R792 VOUT.n517 VOUT.n516 0.476
R793 VOUT.n474 VOUT.n473 0.476
R794 VOUT.n444 VOUT.n443 0.476
R795 VOUT.n401 VOUT.n400 0.476
R796 VOUT.n371 VOUT.n370 0.476
R797 VOUT.n328 VOUT.n327 0.476
R798 VOUT.n298 VOUT.n297 0.476
R799 VOUT.n1136 VOUT.n1135 0.476
R800 VOUT.n1106 VOUT.n1105 0.476
R801 VOUT.n1063 VOUT.n1062 0.476
R802 VOUT.n1033 VOUT.n1032 0.476
R803 VOUT.n990 VOUT.n989 0.476
R804 VOUT.n960 VOUT.n959 0.476
R805 VOUT.n768 VOUT.n767 0.476
R806 VOUT.n738 VOUT.n737 0.476
R807 VOUT.n841 VOUT.n840 0.476
R808 VOUT.n811 VOUT.n810 0.476
R809 VOUT.n914 VOUT.n913 0.476
R810 VOUT.n884 VOUT.n883 0.476
R811 VOUT.n1196 VOUT.n1195 0.476
R812 VOUT.n1297 VOUT.n1296 0.445
R813 VOUT.n1177 VOUT.n1176 0.445
R814 VOUT.n1253 VOUT.n1252 0.445
R815 VOUT.n1206 VOUT.n1205 0.445
R816 VOUT.n1291 VOUT.n1290 0.414
R817 VOUT.n1171 VOUT.n1170 0.414
R818 VOUT.n1258 VOUT.n1257 0.414
R819 VOUT.n703 VOUT.n702 0.414
R820 VOUT.n654 VOUT.n653 0.414
R821 VOUT.n630 VOUT.n629 0.414
R822 VOUT.n581 VOUT.n580 0.414
R823 VOUT.n557 VOUT.n556 0.414
R824 VOUT.n508 VOUT.n507 0.414
R825 VOUT.n484 VOUT.n483 0.414
R826 VOUT.n435 VOUT.n434 0.414
R827 VOUT.n411 VOUT.n410 0.414
R828 VOUT.n362 VOUT.n361 0.414
R829 VOUT.n338 VOUT.n337 0.414
R830 VOUT.n289 VOUT.n288 0.414
R831 VOUT.n1146 VOUT.n1145 0.414
R832 VOUT.n1097 VOUT.n1096 0.414
R833 VOUT.n1073 VOUT.n1072 0.414
R834 VOUT.n1024 VOUT.n1023 0.414
R835 VOUT.n1000 VOUT.n999 0.414
R836 VOUT.n951 VOUT.n950 0.414
R837 VOUT.n778 VOUT.n777 0.414
R838 VOUT.n729 VOUT.n728 0.414
R839 VOUT.n851 VOUT.n850 0.414
R840 VOUT.n802 VOUT.n801 0.414
R841 VOUT.n924 VOUT.n923 0.414
R842 VOUT.n875 VOUT.n874 0.414
R843 VOUT.n1212 VOUT.n1211 0.413
R844 VOUT.n1285 VOUT.n1284 0.382
R845 VOUT.n1165 VOUT.n1164 0.382
R846 VOUT.n1265 VOUT.n1264 0.382
R847 VOUT.n1219 VOUT.n1218 0.382
R848 VOUT.n1149 VOUT.n1148 0.271
R849 VOUT.n1309 VOUT.n236 0.244
R850 VOUT.n706 VOUT.n340 0.228
R851 VOUT.n706 VOUT.n413 0.228
R852 VOUT.n706 VOUT.n486 0.228
R853 VOUT.n706 VOUT.n559 0.228
R854 VOUT.n706 VOUT.n632 0.228
R855 VOUT.n706 VOUT.n705 0.228
R856 VOUT.n1149 VOUT.n1075 0.228
R857 VOUT.n113 VOUT.n1002 0.228
R858 VOUT.n112 VOUT.n780 0.228
R859 VOUT.n929 VOUT.n853 0.228
R860 VOUT.n928 VOUT.n926 0.228
R861 VOUT.n190 VOUT.n707 0.169
R862 VOUT.n234 VOUT.n1229 0.103
R863 VOUT.n52 VOUT.n0 0.079
R864 VOUT.n700 VOUT.n191 0.079
R865 VOUT.n664 VOUT.n661 0.079
R866 VOUT.n50 VOUT.n656 0.079
R867 VOUT.n652 VOUT.n67 0.079
R868 VOUT.n53 VOUT.n1 0.079
R869 VOUT.n627 VOUT.n193 0.079
R870 VOUT.n591 VOUT.n588 0.079
R871 VOUT.n48 VOUT.n583 0.079
R872 VOUT.n579 VOUT.n71 0.079
R873 VOUT.n54 VOUT.n2 0.079
R874 VOUT.n554 VOUT.n195 0.079
R875 VOUT.n518 VOUT.n515 0.079
R876 VOUT.n46 VOUT.n510 0.079
R877 VOUT.n506 VOUT.n75 0.079
R878 VOUT.n55 VOUT.n3 0.079
R879 VOUT.n481 VOUT.n197 0.079
R880 VOUT.n445 VOUT.n442 0.079
R881 VOUT.n44 VOUT.n437 0.079
R882 VOUT.n433 VOUT.n79 0.079
R883 VOUT.n56 VOUT.n4 0.079
R884 VOUT.n408 VOUT.n199 0.079
R885 VOUT.n372 VOUT.n369 0.079
R886 VOUT.n42 VOUT.n364 0.079
R887 VOUT.n360 VOUT.n83 0.079
R888 VOUT.n57 VOUT.n5 0.079
R889 VOUT.n335 VOUT.n201 0.079
R890 VOUT.n299 VOUT.n296 0.079
R891 VOUT.n40 VOUT.n291 0.079
R892 VOUT.n287 VOUT.n87 0.079
R893 VOUT.n58 VOUT.n6 0.079
R894 VOUT.n1143 VOUT.n203 0.079
R895 VOUT.n1107 VOUT.n1104 0.079
R896 VOUT.n38 VOUT.n1099 0.079
R897 VOUT.n1095 VOUT.n91 0.079
R898 VOUT.n59 VOUT.n7 0.079
R899 VOUT.n1070 VOUT.n205 0.079
R900 VOUT.n1034 VOUT.n1031 0.079
R901 VOUT.n36 VOUT.n1026 0.079
R902 VOUT.n1022 VOUT.n95 0.079
R903 VOUT.n60 VOUT.n8 0.079
R904 VOUT.n997 VOUT.n207 0.079
R905 VOUT.n961 VOUT.n958 0.079
R906 VOUT.n34 VOUT.n953 0.079
R907 VOUT.n949 VOUT.n99 0.079
R908 VOUT.n61 VOUT.n9 0.079
R909 VOUT.n775 VOUT.n209 0.079
R910 VOUT.n739 VOUT.n736 0.079
R911 VOUT.n32 VOUT.n731 0.079
R912 VOUT.n727 VOUT.n103 0.079
R913 VOUT.n62 VOUT.n10 0.079
R914 VOUT.n848 VOUT.n211 0.079
R915 VOUT.n812 VOUT.n809 0.079
R916 VOUT.n30 VOUT.n804 0.079
R917 VOUT.n800 VOUT.n107 0.079
R918 VOUT.n63 VOUT.n11 0.079
R919 VOUT.n921 VOUT.n213 0.079
R920 VOUT.n885 VOUT.n882 0.079
R921 VOUT.n28 VOUT.n877 0.079
R922 VOUT.n873 VOUT.n111 0.079
R923 VOUT.n694 VOUT.n244 0.076
R924 VOUT.n621 VOUT.n246 0.076
R925 VOUT.n548 VOUT.n248 0.076
R926 VOUT.n475 VOUT.n250 0.076
R927 VOUT.n402 VOUT.n252 0.076
R928 VOUT.n329 VOUT.n254 0.076
R929 VOUT.n1137 VOUT.n256 0.076
R930 VOUT.n1064 VOUT.n258 0.076
R931 VOUT.n991 VOUT.n260 0.076
R932 VOUT.n769 VOUT.n262 0.076
R933 VOUT.n842 VOUT.n264 0.076
R934 VOUT.n915 VOUT.n266 0.076
R935 VOUT.n1295 VOUT.n155 0.073
R936 VOUT.n1175 VOUT.n158 0.073
R937 VOUT.n160 VOUT.n1207 0.073
R938 VOUT.n163 VOUT.n1254 0.073
R939 VOUT.n1309 VOUT.n190 0.073
R940 VOUT.n141 VOUT.n1283 0.073
R941 VOUT.n138 VOUT.n1163 0.073
R942 VOUT.n139 VOUT.n1217 0.073
R943 VOUT.n140 VOUT.n1263 0.073
R944 VOUT.n1169 VOUT.n1168 0.072
R945 VOUT.n1201 VOUT.n25 0.072
R946 VOUT.n1247 VOUT.n24 0.072
R947 VOUT.n1289 VOUT.n1288 0.072
R948 VOUT.n1223 VOUT.n1222 0.072
R949 VOUT.n1269 VOUT.n1268 0.072
R950 VOUT.n1301 VOUT.n216 0.068
R951 VOUT.n1181 VOUT.n218 0.068
R952 VOUT.n1194 VOUT.n1193 0.068
R953 VOUT.n1240 VOUT.n1239 0.068
R954 VOUT.n166 VOUT.n667 0.064
R955 VOUT.n168 VOUT.n594 0.064
R956 VOUT.n170 VOUT.n521 0.064
R957 VOUT.n172 VOUT.n448 0.064
R958 VOUT.n174 VOUT.n375 0.064
R959 VOUT.n176 VOUT.n302 0.064
R960 VOUT.n178 VOUT.n1110 0.064
R961 VOUT.n180 VOUT.n1037 0.064
R962 VOUT.n182 VOUT.n964 0.064
R963 VOUT.n184 VOUT.n742 0.064
R964 VOUT.n186 VOUT.n815 0.064
R965 VOUT.n188 VOUT.n888 0.064
R966 VOUT.n245 VOUT.n115 0.126
R967 VOUT.n247 VOUT.n117 0.126
R968 VOUT.n249 VOUT.n119 0.126
R969 VOUT.n251 VOUT.n121 0.126
R970 VOUT.n253 VOUT.n123 0.126
R971 VOUT.n255 VOUT.n125 0.126
R972 VOUT.n257 VOUT.n127 0.126
R973 VOUT.n259 VOUT.n129 0.126
R974 VOUT.n261 VOUT.n131 0.126
R975 VOUT.n263 VOUT.n133 0.126
R976 VOUT.n265 VOUT.n135 0.126
R977 VOUT.n267 VOUT.n137 0.126
R978 VOUT.n1269 VOUT.n164 0.057
R979 VOUT.n154 VOUT.n1289 0.057
R980 VOUT.n1223 VOUT.n161 0.057
R981 VOUT.n157 VOUT.n1169 0.057
R982 VOUT.n1283 VOUT.n1281 0.054
R983 VOUT.n1163 VOUT.n1161 0.054
R984 VOUT.n1217 VOUT.n1215 0.054
R985 VOUT.n1263 VOUT.n1261 0.054
R986 VOUT.n1308 VOUT.n1273 0.054
R987 VOUT.n1188 VOUT.n1153 0.054
R988 VOUT.n1188 VOUT.n26 0.054
R989 VOUT.n1308 VOUT.n27 0.054
R990 VOUT.n156 VOUT.n1277 0.053
R991 VOUT.n679 VOUT.n678 0.106
R992 VOUT.n606 VOUT.n605 0.106
R993 VOUT.n533 VOUT.n532 0.106
R994 VOUT.n460 VOUT.n459 0.106
R995 VOUT.n387 VOUT.n386 0.106
R996 VOUT.n314 VOUT.n313 0.106
R997 VOUT.n1122 VOUT.n1121 0.106
R998 VOUT.n1049 VOUT.n1048 0.106
R999 VOUT.n976 VOUT.n975 0.106
R1000 VOUT.n754 VOUT.n753 0.106
R1001 VOUT.n827 VOUT.n826 0.106
R1002 VOUT.n900 VOUT.n899 0.106
R1003 VOUT VOUT.n1309 0.052
R1004 VOUT.n675 VOUT.n167 0.112
R1005 VOUT.n602 VOUT.n169 0.112
R1006 VOUT.n529 VOUT.n171 0.112
R1007 VOUT.n456 VOUT.n173 0.112
R1008 VOUT.n383 VOUT.n175 0.112
R1009 VOUT.n310 VOUT.n177 0.112
R1010 VOUT.n1118 VOUT.n179 0.112
R1011 VOUT.n1045 VOUT.n181 0.112
R1012 VOUT.n972 VOUT.n183 0.112
R1013 VOUT.n750 VOUT.n185 0.112
R1014 VOUT.n823 VOUT.n187 0.112
R1015 VOUT.n896 VOUT.n189 0.112
R1016 VOUT.n240 VOUT.n1301 0.048
R1017 VOUT.n241 VOUT.n1181 0.048
R1018 VOUT.n242 VOUT.n1194 0.048
R1019 VOUT.n243 VOUT.n1240 0.048
R1020 VOUT.n114 VOUT.n684 0.109
R1021 VOUT.n116 VOUT.n611 0.109
R1022 VOUT.n118 VOUT.n538 0.109
R1023 VOUT.n120 VOUT.n465 0.109
R1024 VOUT.n122 VOUT.n392 0.109
R1025 VOUT.n124 VOUT.n319 0.109
R1026 VOUT.n126 VOUT.n1127 0.109
R1027 VOUT.n128 VOUT.n1054 0.109
R1028 VOUT.n130 VOUT.n981 0.109
R1029 VOUT.n132 VOUT.n759 0.109
R1030 VOUT.n134 VOUT.n832 0.109
R1031 VOUT.n136 VOUT.n905 0.109
R1032 VOUT.n235 VOUT.n234 0.109
R1033 VOUT.n236 VOUT.n235 0.103
R1034 VOUT.n11 VOUT.n108 0.066
R1035 VOUT.n10 VOUT.n104 0.066
R1036 VOUT.n9 VOUT.n100 0.066
R1037 VOUT.n8 VOUT.n96 0.066
R1038 VOUT.n7 VOUT.n92 0.066
R1039 VOUT.n6 VOUT.n88 0.066
R1040 VOUT.n5 VOUT.n84 0.066
R1041 VOUT.n4 VOUT.n80 0.066
R1042 VOUT.n3 VOUT.n76 0.066
R1043 VOUT.n2 VOUT.n72 0.066
R1044 VOUT.n1 VOUT.n68 0.066
R1045 VOUT.n0 VOUT.n64 0.066
R1046 VOUT.n23 VOUT.n694 0.062
R1047 VOUT.n22 VOUT.n621 0.062
R1048 VOUT.n21 VOUT.n548 0.062
R1049 VOUT.n20 VOUT.n475 0.062
R1050 VOUT.n19 VOUT.n402 0.062
R1051 VOUT.n18 VOUT.n329 0.062
R1052 VOUT.n17 VOUT.n1137 0.062
R1053 VOUT.n16 VOUT.n1064 0.062
R1054 VOUT.n15 VOUT.n991 0.062
R1055 VOUT.n14 VOUT.n769 0.062
R1056 VOUT.n13 VOUT.n842 0.062
R1057 VOUT.n12 VOUT.n915 0.062
R1058 VOUT.n150 VOUT.n63 0.061
R1059 VOUT.n149 VOUT.n62 0.061
R1060 VOUT.n148 VOUT.n61 0.061
R1061 VOUT.n151 VOUT.n60 0.061
R1062 VOUT.n152 VOUT.n59 0.061
R1063 VOUT.n153 VOUT.n58 0.061
R1064 VOUT.n142 VOUT.n57 0.061
R1065 VOUT.n143 VOUT.n56 0.061
R1066 VOUT.n144 VOUT.n55 0.061
R1067 VOUT.n145 VOUT.n54 0.061
R1068 VOUT.n146 VOUT.n53 0.061
R1069 VOUT.n147 VOUT.n52 0.061
R1070 VOUT.n661 VOUT.n51 0.061
R1071 VOUT.n588 VOUT.n49 0.061
R1072 VOUT.n515 VOUT.n47 0.061
R1073 VOUT.n442 VOUT.n45 0.061
R1074 VOUT.n369 VOUT.n43 0.061
R1075 VOUT.n296 VOUT.n41 0.061
R1076 VOUT.n1104 VOUT.n39 0.061
R1077 VOUT.n1031 VOUT.n37 0.061
R1078 VOUT.n958 VOUT.n35 0.061
R1079 VOUT.n736 VOUT.n33 0.061
R1080 VOUT.n809 VOUT.n31 0.061
R1081 VOUT.n882 VOUT.n29 0.061
R1082 VOUT.n111 VOUT.n110 0.059
R1083 VOUT.n107 VOUT.n106 0.059
R1084 VOUT.n103 VOUT.n102 0.059
R1085 VOUT.n99 VOUT.n98 0.059
R1086 VOUT.n95 VOUT.n94 0.059
R1087 VOUT.n91 VOUT.n90 0.059
R1088 VOUT.n87 VOUT.n86 0.059
R1089 VOUT.n83 VOUT.n82 0.059
R1090 VOUT.n79 VOUT.n78 0.059
R1091 VOUT.n75 VOUT.n74 0.059
R1092 VOUT.n71 VOUT.n70 0.059
R1093 VOUT.n67 VOUT.n66 0.059
R1094 VOUT.n27 VOUT.n240 0.058
R1095 VOUT.n26 VOUT.n241 0.058
R1096 VOUT.n25 VOUT.n242 0.058
R1097 VOUT.n24 VOUT.n243 0.058
R1098 VOUT.n137 VOUT.n136 0.056
R1099 VOUT.n135 VOUT.n134 0.056
R1100 VOUT.n133 VOUT.n132 0.056
R1101 VOUT.n131 VOUT.n130 0.056
R1102 VOUT.n129 VOUT.n128 0.056
R1103 VOUT.n127 VOUT.n126 0.056
R1104 VOUT.n125 VOUT.n124 0.056
R1105 VOUT.n123 VOUT.n122 0.056
R1106 VOUT.n121 VOUT.n120 0.056
R1107 VOUT.n119 VOUT.n118 0.056
R1108 VOUT.n117 VOUT.n116 0.056
R1109 VOUT.n115 VOUT.n114 0.056
R1110 VOUT.n189 VOUT.n188 0.054
R1111 VOUT.n187 VOUT.n186 0.054
R1112 VOUT.n185 VOUT.n184 0.054
R1113 VOUT.n183 VOUT.n182 0.054
R1114 VOUT.n181 VOUT.n180 0.054
R1115 VOUT.n179 VOUT.n178 0.054
R1116 VOUT.n177 VOUT.n176 0.054
R1117 VOUT.n175 VOUT.n174 0.054
R1118 VOUT.n173 VOUT.n172 0.054
R1119 VOUT.n171 VOUT.n170 0.054
R1120 VOUT.n169 VOUT.n168 0.054
R1121 VOUT.n167 VOUT.n166 0.054
R1122 VOUT.n164 VOUT.n163 0.054
R1123 VOUT.n161 VOUT.n160 0.054
R1124 VOUT.n158 VOUT.n157 0.054
R1125 VOUT.n1273 VOUT.n156 0.054
R1126 VOUT.n155 VOUT.n154 0.054
R1127 VOUT.n1234 VOUT.n165 0.05
R1128 VOUT.n1228 VOUT.n162 0.05
R1129 VOUT.n159 VOUT.n1157 0.05
R1130 VOUT.n217 VOUT.n1175 0.048
R1131 VOUT.n215 VOUT.n1295 0.048
R1132 VOUT.n190 VOUT.n113 0.048
R1133 VOUT.n66 VOUT.n649 0.043
R1134 VOUT.n70 VOUT.n576 0.043
R1135 VOUT.n74 VOUT.n503 0.043
R1136 VOUT.n78 VOUT.n430 0.043
R1137 VOUT.n82 VOUT.n357 0.043
R1138 VOUT.n86 VOUT.n284 0.043
R1139 VOUT.n707 VOUT.n706 0.043
R1140 VOUT.n90 VOUT.n1092 0.043
R1141 VOUT.n94 VOUT.n1019 0.043
R1142 VOUT.n98 VOUT.n946 0.043
R1143 VOUT.n102 VOUT.n724 0.043
R1144 VOUT.n106 VOUT.n797 0.043
R1145 VOUT.n110 VOUT.n870 0.043
R1146 VOUT.n929 VOUT.n928 0.043
R1147 VOUT.n112 VOUT.n929 0.043
R1148 VOUT.n113 VOUT.n1149 0.043
R1149 VOUT.n113 VOUT.n112 0.042
R1150 VOUT.n1288 VOUT.n141 0.041
R1151 VOUT.n1268 VOUT.n140 0.041
R1152 VOUT.n1222 VOUT.n139 0.041
R1153 VOUT.n1168 VOUT.n138 0.041
R1154 VOUT.n1153 VOUT.n159 0.04
R1155 VOUT.n147 VOUT.n635 0.04
R1156 VOUT.n665 VOUT.n664 0.04
R1157 VOUT.n146 VOUT.n562 0.04
R1158 VOUT.n592 VOUT.n591 0.04
R1159 VOUT.n145 VOUT.n489 0.04
R1160 VOUT.n519 VOUT.n518 0.04
R1161 VOUT.n144 VOUT.n416 0.04
R1162 VOUT.n446 VOUT.n445 0.04
R1163 VOUT.n143 VOUT.n343 0.04
R1164 VOUT.n373 VOUT.n372 0.04
R1165 VOUT.n142 VOUT.n270 0.04
R1166 VOUT.n300 VOUT.n299 0.04
R1167 VOUT.n153 VOUT.n1078 0.04
R1168 VOUT.n1108 VOUT.n1107 0.04
R1169 VOUT.n152 VOUT.n1005 0.04
R1170 VOUT.n1035 VOUT.n1034 0.04
R1171 VOUT.n151 VOUT.n932 0.04
R1172 VOUT.n962 VOUT.n961 0.04
R1173 VOUT.n148 VOUT.n710 0.04
R1174 VOUT.n740 VOUT.n739 0.04
R1175 VOUT.n149 VOUT.n783 0.04
R1176 VOUT.n813 VOUT.n812 0.04
R1177 VOUT.n150 VOUT.n856 0.04
R1178 VOUT.n886 VOUT.n885 0.04
R1179 VOUT.n266 VOUT.n267 0.04
R1180 VOUT.n264 VOUT.n265 0.04
R1181 VOUT.n262 VOUT.n263 0.04
R1182 VOUT.n260 VOUT.n261 0.04
R1183 VOUT.n258 VOUT.n259 0.04
R1184 VOUT.n256 VOUT.n257 0.04
R1185 VOUT.n254 VOUT.n255 0.04
R1186 VOUT.n252 VOUT.n253 0.04
R1187 VOUT.n250 VOUT.n251 0.04
R1188 VOUT.n248 VOUT.n249 0.04
R1189 VOUT.n246 VOUT.n247 0.04
R1190 VOUT.n244 VOUT.n245 0.04
R1191 VOUT.n905 VOUT.n233 0.04
R1192 VOUT.n832 VOUT.n232 0.04
R1193 VOUT.n759 VOUT.n231 0.04
R1194 VOUT.n981 VOUT.n230 0.04
R1195 VOUT.n1054 VOUT.n229 0.04
R1196 VOUT.n1127 VOUT.n228 0.04
R1197 VOUT.n319 VOUT.n227 0.04
R1198 VOUT.n392 VOUT.n226 0.04
R1199 VOUT.n465 VOUT.n225 0.04
R1200 VOUT.n538 VOUT.n224 0.04
R1201 VOUT.n611 VOUT.n223 0.04
R1202 VOUT.n684 VOUT.n222 0.04
R1203 VOUT.n221 VOUT.n1251 0.04
R1204 VOUT.n220 VOUT.n1203 0.04
R1205 VOUT.n1215 VOUT.n219 0.04
R1206 VOUT.n218 VOUT.n217 0.04
R1207 VOUT.n216 VOUT.n215 0.04
R1208 VOUT.n899 VOUT.n214 0.04
R1209 VOUT.n213 VOUT.n12 0.04
R1210 VOUT.n826 VOUT.n212 0.04
R1211 VOUT.n211 VOUT.n13 0.04
R1212 VOUT.n753 VOUT.n210 0.04
R1213 VOUT.n209 VOUT.n14 0.04
R1214 VOUT.n975 VOUT.n208 0.04
R1215 VOUT.n207 VOUT.n15 0.04
R1216 VOUT.n1048 VOUT.n206 0.04
R1217 VOUT.n205 VOUT.n16 0.04
R1218 VOUT.n1121 VOUT.n204 0.04
R1219 VOUT.n203 VOUT.n17 0.04
R1220 VOUT.n313 VOUT.n202 0.04
R1221 VOUT.n201 VOUT.n18 0.04
R1222 VOUT.n386 VOUT.n200 0.04
R1223 VOUT.n199 VOUT.n19 0.04
R1224 VOUT.n459 VOUT.n198 0.04
R1225 VOUT.n197 VOUT.n20 0.04
R1226 VOUT.n532 VOUT.n196 0.04
R1227 VOUT.n195 VOUT.n21 0.04
R1228 VOUT.n605 VOUT.n194 0.04
R1229 VOUT.n193 VOUT.n22 0.04
R1230 VOUT.n678 VOUT.n192 0.04
R1231 VOUT.n191 VOUT.n23 0.04
R1232 VOUT.n29 VOUT.n28 0.04
R1233 VOUT.n31 VOUT.n30 0.04
R1234 VOUT.n33 VOUT.n32 0.04
R1235 VOUT.n35 VOUT.n34 0.04
R1236 VOUT.n37 VOUT.n36 0.04
R1237 VOUT.n39 VOUT.n38 0.04
R1238 VOUT.n41 VOUT.n40 0.04
R1239 VOUT.n43 VOUT.n42 0.04
R1240 VOUT.n45 VOUT.n44 0.04
R1241 VOUT.n47 VOUT.n46 0.04
R1242 VOUT.n49 VOUT.n48 0.04
R1243 VOUT.n51 VOUT.n50 0.04
R1244 VOUT.n866 VOUT.n109 0.04
R1245 VOUT.n793 VOUT.n105 0.04
R1246 VOUT.n720 VOUT.n101 0.04
R1247 VOUT.n942 VOUT.n97 0.04
R1248 VOUT.n1015 VOUT.n93 0.04
R1249 VOUT.n1088 VOUT.n89 0.04
R1250 VOUT.n280 VOUT.n85 0.04
R1251 VOUT.n353 VOUT.n81 0.04
R1252 VOUT.n426 VOUT.n77 0.04
R1253 VOUT.n499 VOUT.n73 0.04
R1254 VOUT.n572 VOUT.n69 0.04
R1255 VOUT.n645 VOUT.n65 0.04
R1256 VOUT.n1207 VOUT.n220 0.039
R1257 VOUT.n1254 VOUT.n221 0.039
R1258 VOUT.n64 VOUT.n700 0.036
R1259 VOUT.n68 VOUT.n627 0.036
R1260 VOUT.n72 VOUT.n554 0.036
R1261 VOUT.n76 VOUT.n481 0.036
R1262 VOUT.n80 VOUT.n408 0.036
R1263 VOUT.n84 VOUT.n335 0.036
R1264 VOUT.n88 VOUT.n1143 0.036
R1265 VOUT.n92 VOUT.n1070 0.036
R1266 VOUT.n96 VOUT.n997 0.036
R1267 VOUT.n100 VOUT.n775 0.036
R1268 VOUT.n104 VOUT.n848 0.036
R1269 VOUT.n108 VOUT.n921 0.036
R1270 VOUT.n1261 VOUT.n239 0.036
R1271 VOUT.n1161 VOUT.n238 0.036
R1272 VOUT.n1281 VOUT.n237 0.036
R1273 VOUT.n666 VOUT.n665 0.033
R1274 VOUT.n656 VOUT.n645 0.033
R1275 VOUT.n593 VOUT.n592 0.033
R1276 VOUT.n583 VOUT.n572 0.033
R1277 VOUT.n520 VOUT.n519 0.033
R1278 VOUT.n510 VOUT.n499 0.033
R1279 VOUT.n447 VOUT.n446 0.033
R1280 VOUT.n437 VOUT.n426 0.033
R1281 VOUT.n374 VOUT.n373 0.033
R1282 VOUT.n364 VOUT.n353 0.033
R1283 VOUT.n301 VOUT.n300 0.033
R1284 VOUT.n291 VOUT.n280 0.033
R1285 VOUT.n1109 VOUT.n1108 0.033
R1286 VOUT.n1099 VOUT.n1088 0.033
R1287 VOUT.n1036 VOUT.n1035 0.033
R1288 VOUT.n1026 VOUT.n1015 0.033
R1289 VOUT.n963 VOUT.n962 0.033
R1290 VOUT.n953 VOUT.n942 0.033
R1291 VOUT.n741 VOUT.n740 0.033
R1292 VOUT.n731 VOUT.n720 0.033
R1293 VOUT.n814 VOUT.n813 0.033
R1294 VOUT.n804 VOUT.n793 0.033
R1295 VOUT.n887 VOUT.n886 0.033
R1296 VOUT.n877 VOUT.n866 0.033
R1297 VOUT.n222 VOUT.n679 0.031
R1298 VOUT.n223 VOUT.n606 0.031
R1299 VOUT.n224 VOUT.n533 0.031
R1300 VOUT.n225 VOUT.n460 0.031
R1301 VOUT.n226 VOUT.n387 0.031
R1302 VOUT.n227 VOUT.n314 0.031
R1303 VOUT.n228 VOUT.n1122 0.031
R1304 VOUT.n229 VOUT.n1049 0.031
R1305 VOUT.n230 VOUT.n976 0.031
R1306 VOUT.n231 VOUT.n754 0.031
R1307 VOUT.n232 VOUT.n827 0.031
R1308 VOUT.n233 VOUT.n900 0.031
R1309 VOUT.n192 VOUT.n675 0.028
R1310 VOUT.n667 VOUT.n666 0.028
R1311 VOUT.n65 VOUT.n652 0.028
R1312 VOUT.n194 VOUT.n602 0.028
R1313 VOUT.n594 VOUT.n593 0.028
R1314 VOUT.n69 VOUT.n579 0.028
R1315 VOUT.n196 VOUT.n529 0.028
R1316 VOUT.n521 VOUT.n520 0.028
R1317 VOUT.n73 VOUT.n506 0.028
R1318 VOUT.n198 VOUT.n456 0.028
R1319 VOUT.n448 VOUT.n447 0.028
R1320 VOUT.n77 VOUT.n433 0.028
R1321 VOUT.n200 VOUT.n383 0.028
R1322 VOUT.n375 VOUT.n374 0.028
R1323 VOUT.n81 VOUT.n360 0.028
R1324 VOUT.n202 VOUT.n310 0.028
R1325 VOUT.n302 VOUT.n301 0.028
R1326 VOUT.n85 VOUT.n287 0.028
R1327 VOUT.n204 VOUT.n1118 0.028
R1328 VOUT.n1110 VOUT.n1109 0.028
R1329 VOUT.n89 VOUT.n1095 0.028
R1330 VOUT.n206 VOUT.n1045 0.028
R1331 VOUT.n1037 VOUT.n1036 0.028
R1332 VOUT.n93 VOUT.n1022 0.028
R1333 VOUT.n208 VOUT.n972 0.028
R1334 VOUT.n964 VOUT.n963 0.028
R1335 VOUT.n97 VOUT.n949 0.028
R1336 VOUT.n210 VOUT.n750 0.028
R1337 VOUT.n742 VOUT.n741 0.028
R1338 VOUT.n101 VOUT.n727 0.028
R1339 VOUT.n212 VOUT.n823 0.028
R1340 VOUT.n815 VOUT.n814 0.028
R1341 VOUT.n105 VOUT.n800 0.028
R1342 VOUT.n214 VOUT.n896 0.028
R1343 VOUT.n888 VOUT.n887 0.028
R1344 VOUT.n109 VOUT.n873 0.028
R1345 S1.n18 S1.t22 5.393
R1346 S1.n8 S1.t3 5.393
R1347 S1.n3 S1.t13 5.393
R1348 S1.n13 S1.t15 5.393
R1349 S1.n7 S1.t7 3.326
R1350 S1.n7 S1.t0 3.326
R1351 S1.n6 S1.t2 3.326
R1352 S1.n6 S1.t5 3.326
R1353 S1.n0 S1.t9 3.326
R1354 S1.n0 S1.t10 3.326
R1355 S1.n1 S1.t6 3.326
R1356 S1.n1 S1.t8 3.326
R1357 S1.n2 S1.t1 3.326
R1358 S1.n2 S1.t4 3.326
R1359 S1.n12 S1.t18 3.326
R1360 S1.n12 S1.t11 3.326
R1361 S1.n11 S1.t14 3.326
R1362 S1.n11 S1.t17 3.326
R1363 S1.n15 S1.t19 3.326
R1364 S1.n15 S1.t21 3.326
R1365 S1.n16 S1.t16 3.326
R1366 S1.n16 S1.t20 3.326
R1367 S1.n17 S1.t12 3.326
R1368 S1.n17 S1.t23 3.326
R1369 S1.n8 S1.n7 1.79
R1370 S1.n9 S1.n6 1.79
R1371 S1.n5 S1.n0 1.79
R1372 S1.n4 S1.n1 1.79
R1373 S1.n3 S1.n2 1.79
R1374 S1.n13 S1.n12 1.79
R1375 S1.n14 S1.n11 1.79
R1376 S1.n20 S1.n15 1.79
R1377 S1.n19 S1.n16 1.79
R1378 S1.n18 S1.n17 1.79
R1379 S1.n9 S1.n8 0.307
R1380 S1.n5 S1.n4 0.307
R1381 S1.n4 S1.n3 0.307
R1382 S1.n14 S1.n13 0.307
R1383 S1.n20 S1.n19 0.307
R1384 S1.n19 S1.n18 0.307
R1385 S1.n10 S1.n9 0.3
R1386 S1.n21 S1.n14 0.3
R1387 S1.n22 S1.n21 0.049
R1388 S1.n23 S1 0.03
R1389 S1.n23 S1.n22 0.028
R1390 S1 S1.n23 0.024
R1391 S1.n10 S1.n5 0.007
R1392 S1.n21 S1.n20 0.007
R1393 S1.n22 S1.n10 0.001
R1394 D1.n6 D1.t14 5.416
R1395 D1.n8 D1.t6 5.416
R1396 D1.n11 D1.t0 5.414
R1397 D1.n4 D1.t11 5.414
R1398 D1.n3 D1.t4 3.326
R1399 D1.n3 D1.t13 3.326
R1400 D1.n2 D1.t5 3.326
R1401 D1.n2 D1.t12 3.326
R1402 D1.n5 D1.t1 3.326
R1403 D1.n5 D1.t8 3.326
R1404 D1.n10 D1.t7 3.326
R1405 D1.n10 D1.t3 3.326
R1406 D1.n9 D1.t15 3.326
R1407 D1.n9 D1.t9 3.326
R1408 D1.n7 D1.t10 3.326
R1409 D1.n7 D1.t2 3.326
R1410 D1.n4 D1.n3 1.766
R1411 D1.n0 D1.n2 1.766
R1412 D1.n6 D1.n5 1.766
R1413 D1.n11 D1.n10 1.766
R1414 D1.n1 D1.n9 1.766
R1415 D1.n8 D1.n7 1.766
R1416 D1.n0 D1.n4 0.352
R1417 D1.n1 D1.n11 0.352
R1418 D1.n0 D1.n6 0.35
R1419 D1.n1 D1.n8 0.35
R1420 D1.n12 D1.n0 0.106
R1421 D1 D1.n12 0.098
R1422 D1.n12 D1.n1 0.056
R1423 SS.n539 SS.n538 9.3
R1424 SS.n559 SS.n558 9.3
R1425 SS.n583 SS.n582 9.3
R1426 SS.n520 SS.n519 9.3
R1427 SS.n525 SS.n524 9.3
R1428 SS.n530 SS.n529 9.3
R1429 SS.n535 SS.n534 9.3
R1430 SS.n541 SS.n540 9.3
R1431 SS.n545 SS.n544 9.3
R1432 SS.n557 SS.n556 9.3
R1433 SS.n561 SS.n560 9.3
R1434 SS.n568 SS.n567 9.3
R1435 SS.n570 SS.n569 9.3
R1436 SS.n572 SS.n571 9.3
R1437 SS.n597 SS.n596 9.3
R1438 SS.n605 SS.n604 9.3
R1439 SS.n616 SS.n615 9.3
R1440 SS.n619 SS.n618 9.3
R1441 SS.n622 SS.n621 9.3
R1442 SS.n638 SS.n637 9.3
R1443 SS.n632 SS.n631 9.3
R1444 SS.n628 SS.n627 9.3
R1445 SS.n612 SS.n611 9.3
R1446 SS.n608 SS.n607 9.3
R1447 SS.n603 SS.n602 9.3
R1448 SS.n594 SS.n593 9.3
R1449 SS.n592 SS.n591 9.3
R1450 SS.n586 SS.n585 9.3
R1451 SS.n581 SS.n580 9.3
R1452 SS.n378 SS.n377 9.3
R1453 SS.n398 SS.n397 9.3
R1454 SS.n422 SS.n421 9.3
R1455 SS.n359 SS.n358 9.3
R1456 SS.n364 SS.n363 9.3
R1457 SS.n369 SS.n368 9.3
R1458 SS.n374 SS.n373 9.3
R1459 SS.n380 SS.n379 9.3
R1460 SS.n384 SS.n383 9.3
R1461 SS.n396 SS.n395 9.3
R1462 SS.n400 SS.n399 9.3
R1463 SS.n407 SS.n406 9.3
R1464 SS.n409 SS.n408 9.3
R1465 SS.n411 SS.n410 9.3
R1466 SS.n436 SS.n435 9.3
R1467 SS.n444 SS.n443 9.3
R1468 SS.n455 SS.n454 9.3
R1469 SS.n458 SS.n457 9.3
R1470 SS.n461 SS.n460 9.3
R1471 SS.n477 SS.n476 9.3
R1472 SS.n471 SS.n470 9.3
R1473 SS.n467 SS.n466 9.3
R1474 SS.n451 SS.n450 9.3
R1475 SS.n447 SS.n446 9.3
R1476 SS.n442 SS.n441 9.3
R1477 SS.n433 SS.n432 9.3
R1478 SS.n431 SS.n430 9.3
R1479 SS.n425 SS.n424 9.3
R1480 SS.n420 SS.n419 9.3
R1481 SS.n217 SS.n216 9.3
R1482 SS.n237 SS.n236 9.3
R1483 SS.n261 SS.n260 9.3
R1484 SS.n198 SS.n197 9.3
R1485 SS.n203 SS.n202 9.3
R1486 SS.n208 SS.n207 9.3
R1487 SS.n213 SS.n212 9.3
R1488 SS.n219 SS.n218 9.3
R1489 SS.n223 SS.n222 9.3
R1490 SS.n235 SS.n234 9.3
R1491 SS.n239 SS.n238 9.3
R1492 SS.n246 SS.n245 9.3
R1493 SS.n248 SS.n247 9.3
R1494 SS.n250 SS.n249 9.3
R1495 SS.n275 SS.n274 9.3
R1496 SS.n283 SS.n282 9.3
R1497 SS.n294 SS.n293 9.3
R1498 SS.n297 SS.n296 9.3
R1499 SS.n300 SS.n299 9.3
R1500 SS.n316 SS.n315 9.3
R1501 SS.n310 SS.n309 9.3
R1502 SS.n306 SS.n305 9.3
R1503 SS.n290 SS.n289 9.3
R1504 SS.n286 SS.n285 9.3
R1505 SS.n281 SS.n280 9.3
R1506 SS.n272 SS.n271 9.3
R1507 SS.n270 SS.n269 9.3
R1508 SS.n264 SS.n263 9.3
R1509 SS.n259 SS.n258 9.3
R1510 SS.n56 SS.n55 9.3
R1511 SS.n76 SS.n75 9.3
R1512 SS.n100 SS.n99 9.3
R1513 SS.n37 SS.n36 9.3
R1514 SS.n42 SS.n41 9.3
R1515 SS.n47 SS.n46 9.3
R1516 SS.n52 SS.n51 9.3
R1517 SS.n58 SS.n57 9.3
R1518 SS.n62 SS.n61 9.3
R1519 SS.n74 SS.n73 9.3
R1520 SS.n78 SS.n77 9.3
R1521 SS.n85 SS.n84 9.3
R1522 SS.n87 SS.n86 9.3
R1523 SS.n89 SS.n88 9.3
R1524 SS.n114 SS.n113 9.3
R1525 SS.n122 SS.n121 9.3
R1526 SS.n133 SS.n132 9.3
R1527 SS.n136 SS.n135 9.3
R1528 SS.n139 SS.n138 9.3
R1529 SS.n155 SS.n154 9.3
R1530 SS.n149 SS.n148 9.3
R1531 SS.n145 SS.n144 9.3
R1532 SS.n129 SS.n128 9.3
R1533 SS.n125 SS.n124 9.3
R1534 SS.n120 SS.n119 9.3
R1535 SS.n111 SS.n110 9.3
R1536 SS.n109 SS.n108 9.3
R1537 SS.n103 SS.n102 9.3
R1538 SS.n98 SS.n97 9.3
R1539 SS.n704 SS.n703 9.3
R1540 SS.n724 SS.n723 9.3
R1541 SS.n748 SS.n747 9.3
R1542 SS.n685 SS.n684 9.3
R1543 SS.n690 SS.n689 9.3
R1544 SS.n695 SS.n694 9.3
R1545 SS.n700 SS.n699 9.3
R1546 SS.n706 SS.n705 9.3
R1547 SS.n710 SS.n709 9.3
R1548 SS.n722 SS.n721 9.3
R1549 SS.n726 SS.n725 9.3
R1550 SS.n733 SS.n732 9.3
R1551 SS.n735 SS.n734 9.3
R1552 SS.n737 SS.n736 9.3
R1553 SS.n762 SS.n761 9.3
R1554 SS.n770 SS.n769 9.3
R1555 SS.n781 SS.n780 9.3
R1556 SS.n784 SS.n783 9.3
R1557 SS.n787 SS.n786 9.3
R1558 SS.n803 SS.n802 9.3
R1559 SS.n797 SS.n796 9.3
R1560 SS.n793 SS.n792 9.3
R1561 SS.n777 SS.n776 9.3
R1562 SS.n773 SS.n772 9.3
R1563 SS.n768 SS.n767 9.3
R1564 SS.n759 SS.n758 9.3
R1565 SS.n757 SS.n756 9.3
R1566 SS.n751 SS.n750 9.3
R1567 SS.n746 SS.n745 9.3
R1568 SS.n865 SS.n864 9.3
R1569 SS.n885 SS.n884 9.3
R1570 SS.n909 SS.n908 9.3
R1571 SS.n846 SS.n845 9.3
R1572 SS.n851 SS.n850 9.3
R1573 SS.n856 SS.n855 9.3
R1574 SS.n861 SS.n860 9.3
R1575 SS.n867 SS.n866 9.3
R1576 SS.n871 SS.n870 9.3
R1577 SS.n883 SS.n882 9.3
R1578 SS.n887 SS.n886 9.3
R1579 SS.n894 SS.n893 9.3
R1580 SS.n896 SS.n895 9.3
R1581 SS.n898 SS.n897 9.3
R1582 SS.n923 SS.n922 9.3
R1583 SS.n931 SS.n930 9.3
R1584 SS.n942 SS.n941 9.3
R1585 SS.n945 SS.n944 9.3
R1586 SS.n948 SS.n947 9.3
R1587 SS.n964 SS.n963 9.3
R1588 SS.n958 SS.n957 9.3
R1589 SS.n954 SS.n953 9.3
R1590 SS.n938 SS.n937 9.3
R1591 SS.n934 SS.n933 9.3
R1592 SS.n929 SS.n928 9.3
R1593 SS.n920 SS.n919 9.3
R1594 SS.n918 SS.n917 9.3
R1595 SS.n912 SS.n911 9.3
R1596 SS.n907 SS.n906 9.3
R1597 SS.n1192 SS.n1191 9.3
R1598 SS.n1212 SS.n1211 9.3
R1599 SS.n1236 SS.n1235 9.3
R1600 SS.n1225 SS.n1224 9.3
R1601 SS.n1223 SS.n1222 9.3
R1602 SS.n1221 SS.n1220 9.3
R1603 SS.n1214 SS.n1213 9.3
R1604 SS.n1210 SS.n1209 9.3
R1605 SS.n1198 SS.n1197 9.3
R1606 SS.n1194 SS.n1193 9.3
R1607 SS.n1188 SS.n1187 9.3
R1608 SS.n1183 SS.n1182 9.3
R1609 SS.n1178 SS.n1177 9.3
R1610 SS.n1173 SS.n1172 9.3
R1611 SS.n1272 SS.n1271 9.3
R1612 SS.n1258 SS.n1257 9.3
R1613 SS.n1245 SS.n1244 9.3
R1614 SS.n1247 SS.n1246 9.3
R1615 SS.n1250 SS.n1249 9.3
R1616 SS.n1291 SS.n1290 9.3
R1617 SS.n1285 SS.n1284 9.3
R1618 SS.n1281 SS.n1280 9.3
R1619 SS.n1275 SS.n1274 9.3
R1620 SS.n1269 SS.n1268 9.3
R1621 SS.n1265 SS.n1264 9.3
R1622 SS.n1261 SS.n1260 9.3
R1623 SS.n1256 SS.n1255 9.3
R1624 SS.n1239 SS.n1238 9.3
R1625 SS.n1234 SS.n1233 9.3
R1626 SS.n1027 SS.n1026 9.3
R1627 SS.n1047 SS.n1046 9.3
R1628 SS.n1071 SS.n1070 9.3
R1629 SS.n1013 SS.n1012 9.3
R1630 SS.n1023 SS.n1022 9.3
R1631 SS.n1033 SS.n1032 9.3
R1632 SS.n1049 SS.n1048 9.3
R1633 SS.n1058 SS.n1057 9.3
R1634 SS.n1060 SS.n1059 9.3
R1635 SS.n1093 SS.n1092 9.3
R1636 SS.n1107 SS.n1106 9.3
R1637 SS.n1110 SS.n1109 9.3
R1638 SS.n1120 SS.n1119 9.3
R1639 SS.n1100 SS.n1099 9.3
R1640 SS.n1091 SS.n1090 9.3
R1641 SS.n1082 SS.n1081 9.3
R1642 SS.n1080 SS.n1079 9.3
R1643 SS.n1069 SS.n1068 9.3
R1644 SS.n1008 SS.n1007 9.3
R1645 SS.n1018 SS.n1017 9.3
R1646 SS.n1029 SS.n1028 9.3
R1647 SS.n1045 SS.n1044 9.3
R1648 SS.n1056 SS.n1055 9.3
R1649 SS.n1085 SS.n1084 9.3
R1650 SS.n1104 SS.n1103 9.3
R1651 SS.n1126 SS.n1125 9.3
R1652 SS.n1116 SS.n1115 9.3
R1653 SS.n1096 SS.n1095 9.3
R1654 SS.n1074 SS.n1073 9.3
R1655 SS.n640 SS.n633 9
R1656 SS.n523 SS.n522 9
R1657 SS.n532 SS.n531 9
R1658 SS.n543 SS.n542 9
R1659 SS.n563 SS.n562 9
R1660 SS.n574 SS.n573 9
R1661 SS.n590 SS.n589 9
R1662 SS.n625 SS.n624 9
R1663 SS.n614 SS.n613 9
R1664 SS.n601 SS.n600 9
R1665 SS.n579 SS.n578 9
R1666 SS.n479 SS.n472 9
R1667 SS.n362 SS.n361 9
R1668 SS.n371 SS.n370 9
R1669 SS.n382 SS.n381 9
R1670 SS.n402 SS.n401 9
R1671 SS.n413 SS.n412 9
R1672 SS.n429 SS.n428 9
R1673 SS.n464 SS.n463 9
R1674 SS.n453 SS.n452 9
R1675 SS.n440 SS.n439 9
R1676 SS.n418 SS.n417 9
R1677 SS.n318 SS.n311 9
R1678 SS.n201 SS.n200 9
R1679 SS.n210 SS.n209 9
R1680 SS.n221 SS.n220 9
R1681 SS.n241 SS.n240 9
R1682 SS.n252 SS.n251 9
R1683 SS.n268 SS.n267 9
R1684 SS.n303 SS.n302 9
R1685 SS.n292 SS.n291 9
R1686 SS.n279 SS.n278 9
R1687 SS.n257 SS.n256 9
R1688 SS.n157 SS.n150 9
R1689 SS.n40 SS.n39 9
R1690 SS.n49 SS.n48 9
R1691 SS.n60 SS.n59 9
R1692 SS.n80 SS.n79 9
R1693 SS.n91 SS.n90 9
R1694 SS.n107 SS.n106 9
R1695 SS.n142 SS.n141 9
R1696 SS.n131 SS.n130 9
R1697 SS.n118 SS.n117 9
R1698 SS.n96 SS.n95 9
R1699 SS.n805 SS.n798 9
R1700 SS.n688 SS.n687 9
R1701 SS.n697 SS.n696 9
R1702 SS.n708 SS.n707 9
R1703 SS.n728 SS.n727 9
R1704 SS.n739 SS.n738 9
R1705 SS.n755 SS.n754 9
R1706 SS.n790 SS.n789 9
R1707 SS.n779 SS.n778 9
R1708 SS.n766 SS.n765 9
R1709 SS.n744 SS.n743 9
R1710 SS.n966 SS.n959 9
R1711 SS.n849 SS.n848 9
R1712 SS.n858 SS.n857 9
R1713 SS.n869 SS.n868 9
R1714 SS.n889 SS.n888 9
R1715 SS.n900 SS.n899 9
R1716 SS.n916 SS.n915 9
R1717 SS.n951 SS.n950 9
R1718 SS.n940 SS.n939 9
R1719 SS.n927 SS.n926 9
R1720 SS.n905 SS.n904 9
R1721 SS.n1176 SS.n1175 9
R1722 SS.n1185 SS.n1184 9
R1723 SS.n1196 SS.n1195 9
R1724 SS.n1216 SS.n1215 9
R1725 SS.n1227 SS.n1226 9
R1726 SS.n1293 SS.n1286 9
R1727 SS.n1278 SS.n1277 9
R1728 SS.n1267 SS.n1266 9
R1729 SS.n1243 SS.n1242 9
R1730 SS.n1254 SS.n1253 9
R1731 SS.n1232 SS.n1231 9
R1732 SS.n1128 SS.n1121 9
R1733 SS.n1011 SS.n1010 9
R1734 SS.n1020 SS.n1019 9
R1735 SS.n1031 SS.n1030 9
R1736 SS.n1051 SS.n1050 9
R1737 SS.n1062 SS.n1061 9
R1738 SS.n1078 SS.n1077 9
R1739 SS.n1113 SS.n1112 9
R1740 SS.n1102 SS.n1101 9
R1741 SS.n1089 SS.n1088 9
R1742 SS.n1067 SS.n1066 9
R1743 SS.n578 SS.n577 8.282
R1744 SS.n417 SS.n416 8.282
R1745 SS.n256 SS.n255 8.282
R1746 SS.n95 SS.n94 8.282
R1747 SS.n743 SS.n742 8.282
R1748 SS.n904 SS.n903 8.282
R1749 SS.n1231 SS.n1230 8.282
R1750 SS.n1066 SS.n1065 8.282
R1751 SS.n636 SS.n635 7.853
R1752 SS.n475 SS.n474 7.853
R1753 SS.n314 SS.n313 7.853
R1754 SS.n153 SS.n152 7.853
R1755 SS.n801 SS.n800 7.853
R1756 SS.n962 SS.n961 7.853
R1757 SS.n1289 SS.n1288 7.853
R1758 SS.n1124 SS.n1123 7.853
R1759 SS.n1006 SS.n1005 7.852
R1760 SS.n518 SS.n517 7.851
R1761 SS.n357 SS.n356 7.851
R1762 SS.n196 SS.n195 7.851
R1763 SS.n35 SS.n34 7.851
R1764 SS.n683 SS.n682 7.851
R1765 SS.n844 SS.n843 7.851
R1766 SS.n1171 SS.n1170 7.851
R1767 SS.n550 SS.n549 4.65
R1768 SS.n389 SS.n388 4.65
R1769 SS.n228 SS.n227 4.65
R1770 SS.n67 SS.n66 4.65
R1771 SS.n715 SS.n714 4.65
R1772 SS.n876 SS.n875 4.65
R1773 SS.n1203 SS.n1202 4.65
R1774 SS.n1038 SS.n1037 4.65
R1775 SS.n552 SS.n551 4.574
R1776 SS.n391 SS.n390 4.574
R1777 SS.n230 SS.n229 4.574
R1778 SS.n69 SS.n68 4.574
R1779 SS.n717 SS.n716 4.574
R1780 SS.n878 SS.n877 4.574
R1781 SS.n1205 SS.n1204 4.574
R1782 SS.n1040 SS.n1039 4.574
R1783 SS.n634 SS.t6 3.326
R1784 SS.n634 SS.t9 3.326
R1785 SS.n473 SS.t2 3.326
R1786 SS.n473 SS.t5 3.326
R1787 SS.n312 SS.t1 3.326
R1788 SS.n312 SS.t3 3.326
R1789 SS.n151 SS.t4 3.326
R1790 SS.n151 SS.t8 3.326
R1791 SS.n799 SS.t13 3.326
R1792 SS.n799 SS.t0 3.326
R1793 SS.n960 SS.t7 3.326
R1794 SS.n960 SS.t11 3.326
R1795 SS.n1287 SS.t12 3.326
R1796 SS.n1287 SS.t15 3.326
R1797 SS.n1122 SS.t10 3.326
R1798 SS.n1122 SS.t14 3.326
R1799 SS.n618 SS.n617 3.191
R1800 SS.n457 SS.n456 3.191
R1801 SS.n296 SS.n295 3.191
R1802 SS.n135 SS.n134 3.191
R1803 SS.n783 SS.n782 3.191
R1804 SS.n944 SS.n943 3.191
R1805 SS.n1271 SS.n1270 3.191
R1806 SS.n1106 SS.n1105 3.191
R1807 SS.n641 SS.n640 3
R1808 SS.n480 SS.n479 3
R1809 SS.n319 SS.n318 3
R1810 SS.n158 SS.n157 3
R1811 SS.n806 SS.n805 3
R1812 SS.n967 SS.n966 3
R1813 SS.n1294 SS.n1293 3
R1814 SS.n1129 SS.n1128 3
R1815 SS.n538 SS.n537 2.814
R1816 SS.n377 SS.n376 2.814
R1817 SS.n216 SS.n215 2.814
R1818 SS.n55 SS.n54 2.814
R1819 SS.n703 SS.n702 2.814
R1820 SS.n864 SS.n863 2.814
R1821 SS.n1191 SS.n1190 2.814
R1822 SS.n1026 SS.n1025 2.814
R1823 SS.n635 SS.n634 2.082
R1824 SS.n474 SS.n473 2.082
R1825 SS.n313 SS.n312 2.082
R1826 SS.n152 SS.n151 2.082
R1827 SS.n800 SS.n799 2.082
R1828 SS.n961 SS.n960 2.082
R1829 SS.n1288 SS.n1287 2.082
R1830 SS.n1123 SS.n1122 2.082
R1831 SS.n1298 SS.n1297 0.704
R1832 SS.n567 SS.n566 0.536
R1833 SS.n585 SS.n584 0.536
R1834 SS.n406 SS.n405 0.536
R1835 SS.n424 SS.n423 0.536
R1836 SS.n245 SS.n244 0.536
R1837 SS.n263 SS.n262 0.536
R1838 SS.n84 SS.n83 0.536
R1839 SS.n102 SS.n101 0.536
R1840 SS.n732 SS.n731 0.536
R1841 SS.n750 SS.n749 0.536
R1842 SS.n893 SS.n892 0.536
R1843 SS.n911 SS.n910 0.536
R1844 SS.n1220 SS.n1219 0.536
R1845 SS.n1238 SS.n1237 0.536
R1846 SS.n1073 SS.n1072 0.536
R1847 SS.n1055 SS.n1054 0.536
R1848 SS.n556 SS.n555 0.506
R1849 SS.n596 SS.n595 0.506
R1850 SS.n395 SS.n394 0.506
R1851 SS.n435 SS.n434 0.506
R1852 SS.n234 SS.n233 0.506
R1853 SS.n274 SS.n273 0.506
R1854 SS.n73 SS.n72 0.506
R1855 SS.n113 SS.n112 0.506
R1856 SS.n721 SS.n720 0.506
R1857 SS.n761 SS.n760 0.506
R1858 SS.n882 SS.n881 0.506
R1859 SS.n922 SS.n921 0.506
R1860 SS.n1209 SS.n1208 0.506
R1861 SS.n1249 SS.n1248 0.506
R1862 SS.n1084 SS.n1083 0.506
R1863 SS.n1044 SS.n1043 0.506
R1864 SS.n549 SS.n548 0.476
R1865 SS.n607 SS.n606 0.476
R1866 SS.n388 SS.n387 0.476
R1867 SS.n446 SS.n445 0.476
R1868 SS.n227 SS.n226 0.476
R1869 SS.n285 SS.n284 0.476
R1870 SS.n66 SS.n65 0.476
R1871 SS.n124 SS.n123 0.476
R1872 SS.n714 SS.n713 0.476
R1873 SS.n772 SS.n771 0.476
R1874 SS.n875 SS.n874 0.476
R1875 SS.n933 SS.n932 0.476
R1876 SS.n1202 SS.n1201 0.476
R1877 SS.n1260 SS.n1259 0.476
R1878 SS.n1095 SS.n1094 0.476
R1879 SS.n1037 SS.n1036 0.475
R1880 SS.n529 SS.n528 0.414
R1881 SS.n627 SS.n626 0.414
R1882 SS.n368 SS.n367 0.414
R1883 SS.n466 SS.n465 0.414
R1884 SS.n207 SS.n206 0.414
R1885 SS.n305 SS.n304 0.414
R1886 SS.n46 SS.n45 0.414
R1887 SS.n144 SS.n143 0.414
R1888 SS.n694 SS.n693 0.414
R1889 SS.n792 SS.n791 0.414
R1890 SS.n855 SS.n854 0.414
R1891 SS.n953 SS.n952 0.414
R1892 SS.n1182 SS.n1181 0.414
R1893 SS.n1280 SS.n1279 0.414
R1894 SS.n1115 SS.n1114 0.414
R1895 SS.n1017 SS.n1016 0.413
R1896 SS.n1135 SS.n1134 0.312
R1897 SS SS.n1298 0.264
R1898 SS.n1134 SS.n1133 0.217
R1899 SS.n1134 SS.n647 0.192
R1900 SS.n644 SS.n643 0.18
R1901 SS.n645 SS.n482 0.18
R1902 SS.n646 SS.n321 0.18
R1903 SS.n647 SS.n160 0.18
R1904 SS.n1133 SS.n808 0.18
R1905 SS.n970 SS.n969 0.18
R1906 SS.n1297 SS.n1296 0.18
R1907 SS.n1132 SS.n1131 0.18
R1908 SS.n490 SS.n489 0.12
R1909 SS.n493 SS.n492 0.12
R1910 SS.n496 SS.n495 0.12
R1911 SS.n499 SS.n498 0.12
R1912 SS.n503 SS.n502 0.12
R1913 SS.n506 SS.n505 0.12
R1914 SS.n509 SS.n508 0.12
R1915 SS.n512 SS.n511 0.12
R1916 SS.n329 SS.n328 0.12
R1917 SS.n332 SS.n331 0.12
R1918 SS.n335 SS.n334 0.12
R1919 SS.n338 SS.n337 0.12
R1920 SS.n342 SS.n341 0.12
R1921 SS.n345 SS.n344 0.12
R1922 SS.n348 SS.n347 0.12
R1923 SS.n351 SS.n350 0.12
R1924 SS.n168 SS.n167 0.12
R1925 SS.n171 SS.n170 0.12
R1926 SS.n174 SS.n173 0.12
R1927 SS.n177 SS.n176 0.12
R1928 SS.n181 SS.n180 0.12
R1929 SS.n184 SS.n183 0.12
R1930 SS.n187 SS.n186 0.12
R1931 SS.n190 SS.n189 0.12
R1932 SS.n7 SS.n6 0.12
R1933 SS.n10 SS.n9 0.12
R1934 SS.n13 SS.n12 0.12
R1935 SS.n16 SS.n15 0.12
R1936 SS.n20 SS.n19 0.12
R1937 SS.n23 SS.n22 0.12
R1938 SS.n26 SS.n25 0.12
R1939 SS.n29 SS.n28 0.12
R1940 SS.n655 SS.n654 0.12
R1941 SS.n658 SS.n657 0.12
R1942 SS.n661 SS.n660 0.12
R1943 SS.n664 SS.n663 0.12
R1944 SS.n668 SS.n667 0.12
R1945 SS.n671 SS.n670 0.12
R1946 SS.n674 SS.n673 0.12
R1947 SS.n677 SS.n676 0.12
R1948 SS.n816 SS.n815 0.12
R1949 SS.n819 SS.n818 0.12
R1950 SS.n822 SS.n821 0.12
R1951 SS.n825 SS.n824 0.12
R1952 SS.n829 SS.n828 0.12
R1953 SS.n832 SS.n831 0.12
R1954 SS.n835 SS.n834 0.12
R1955 SS.n838 SS.n837 0.12
R1956 SS.n1143 SS.n1142 0.12
R1957 SS.n1146 SS.n1145 0.12
R1958 SS.n1149 SS.n1148 0.12
R1959 SS.n1152 SS.n1151 0.12
R1960 SS.n1156 SS.n1155 0.12
R1961 SS.n1159 SS.n1158 0.12
R1962 SS.n1162 SS.n1161 0.12
R1963 SS.n1165 SS.n1164 0.12
R1964 SS.n978 SS.n977 0.12
R1965 SS.n981 SS.n980 0.12
R1966 SS.n984 SS.n983 0.12
R1967 SS.n987 SS.n986 0.12
R1968 SS.n991 SS.n990 0.12
R1969 SS.n994 SS.n993 0.12
R1970 SS.n997 SS.n996 0.12
R1971 SS.n1000 SS.n999 0.12
R1972 SS.n1015 SS.n1014 0.079
R1973 SS.n1027 SS.n1024 0.079
R1974 SS.n1038 SS.n1035 0.079
R1975 SS.n1108 SS.n1107 0.079
R1976 SS.n1118 SS.n1117 0.079
R1977 SS.n527 SS.n526 0.079
R1978 SS.n539 SS.n536 0.079
R1979 SS.n550 SS.n547 0.079
R1980 SS.n620 SS.n619 0.079
R1981 SS.n630 SS.n629 0.079
R1982 SS.n486 SS.n485 0.079
R1983 SS.n516 SS.n515 0.079
R1984 SS.n366 SS.n365 0.079
R1985 SS.n378 SS.n375 0.079
R1986 SS.n389 SS.n386 0.079
R1987 SS.n459 SS.n458 0.079
R1988 SS.n469 SS.n468 0.079
R1989 SS.n325 SS.n324 0.079
R1990 SS.n355 SS.n354 0.079
R1991 SS.n205 SS.n204 0.079
R1992 SS.n217 SS.n214 0.079
R1993 SS.n228 SS.n225 0.079
R1994 SS.n298 SS.n297 0.079
R1995 SS.n308 SS.n307 0.079
R1996 SS.n164 SS.n163 0.079
R1997 SS.n194 SS.n193 0.079
R1998 SS.n44 SS.n43 0.079
R1999 SS.n56 SS.n53 0.079
R2000 SS.n67 SS.n64 0.079
R2001 SS.n137 SS.n136 0.079
R2002 SS.n147 SS.n146 0.079
R2003 SS.n3 SS.n2 0.079
R2004 SS.n33 SS.n32 0.079
R2005 SS.n692 SS.n691 0.079
R2006 SS.n704 SS.n701 0.079
R2007 SS.n715 SS.n712 0.079
R2008 SS.n785 SS.n784 0.079
R2009 SS.n795 SS.n794 0.079
R2010 SS.n651 SS.n650 0.079
R2011 SS.n681 SS.n680 0.079
R2012 SS.n853 SS.n852 0.079
R2013 SS.n865 SS.n862 0.079
R2014 SS.n876 SS.n873 0.079
R2015 SS.n946 SS.n945 0.079
R2016 SS.n956 SS.n955 0.079
R2017 SS.n812 SS.n811 0.079
R2018 SS.n842 SS.n841 0.079
R2019 SS.n1180 SS.n1179 0.079
R2020 SS.n1192 SS.n1189 0.079
R2021 SS.n1203 SS.n1200 0.079
R2022 SS.n1273 SS.n1272 0.079
R2023 SS.n1283 SS.n1282 0.079
R2024 SS.n1139 SS.n1138 0.079
R2025 SS.n1169 SS.n1168 0.079
R2026 SS.n974 SS.n973 0.079
R2027 SS.n1004 SS.n1003 0.079
R2028 SS.n1097 SS.n1096 0.076
R2029 SS.n609 SS.n608 0.076
R2030 SS.n448 SS.n447 0.076
R2031 SS.n287 SS.n286 0.076
R2032 SS.n126 SS.n125 0.076
R2033 SS.n774 SS.n773 0.076
R2034 SS.n935 SS.n934 0.076
R2035 SS.n1262 SS.n1261 0.076
R2036 SS.n645 SS.n644 0.071
R2037 SS.n646 SS.n645 0.071
R2038 SS.n647 SS.n646 0.071
R2039 SS.n1133 SS.n1132 0.071
R2040 SS.n1132 SS.n970 0.071
R2041 SS.n1045 SS.n1042 0.064
R2042 SS.n557 SS.n554 0.064
R2043 SS.n396 SS.n393 0.064
R2044 SS.n235 SS.n232 0.064
R2045 SS.n74 SS.n71 0.064
R2046 SS.n722 SS.n719 0.064
R2047 SS.n883 SS.n880 0.064
R2048 SS.n1210 SS.n1207 0.064
R2049 SS.n1086 SS.n1085 0.062
R2050 SS.n598 SS.n597 0.062
R2051 SS.n437 SS.n436 0.062
R2052 SS.n276 SS.n275 0.062
R2053 SS.n115 SS.n114 0.062
R2054 SS.n763 SS.n762 0.062
R2055 SS.n924 SS.n923 0.062
R2056 SS.n1251 SS.n1250 0.062
R2057 SS.n1063 SS.n1062 0.052
R2058 SS.n1067 SS.n1064 0.052
R2059 SS.n575 SS.n574 0.052
R2060 SS.n579 SS.n576 0.052
R2061 SS.n500 SS.n499 0.052
R2062 SS.n502 SS.n501 0.052
R2063 SS.n414 SS.n413 0.052
R2064 SS.n418 SS.n415 0.052
R2065 SS.n339 SS.n338 0.052
R2066 SS.n341 SS.n340 0.052
R2067 SS.n253 SS.n252 0.052
R2068 SS.n257 SS.n254 0.052
R2069 SS.n178 SS.n177 0.052
R2070 SS.n180 SS.n179 0.052
R2071 SS.n92 SS.n91 0.052
R2072 SS.n96 SS.n93 0.052
R2073 SS.n17 SS.n16 0.052
R2074 SS.n19 SS.n18 0.052
R2075 SS.n740 SS.n739 0.052
R2076 SS.n744 SS.n741 0.052
R2077 SS.n665 SS.n664 0.052
R2078 SS.n667 SS.n666 0.052
R2079 SS.n901 SS.n900 0.052
R2080 SS.n905 SS.n902 0.052
R2081 SS.n826 SS.n825 0.052
R2082 SS.n828 SS.n827 0.052
R2083 SS.n1228 SS.n1227 0.052
R2084 SS.n1232 SS.n1229 0.052
R2085 SS.n1153 SS.n1152 0.052
R2086 SS.n1155 SS.n1154 0.052
R2087 SS.n988 SS.n987 0.052
R2088 SS.n990 SS.n989 0.052
R2089 SS.n1056 SS.n1053 0.05
R2090 SS.n568 SS.n565 0.05
R2091 SS.n407 SS.n404 0.05
R2092 SS.n246 SS.n243 0.05
R2093 SS.n85 SS.n82 0.05
R2094 SS.n733 SS.n730 0.05
R2095 SS.n894 SS.n891 0.05
R2096 SS.n1221 SS.n1218 0.05
R2097 SS.n1075 SS.n1074 0.048
R2098 SS.n587 SS.n586 0.048
R2099 SS.n487 SS.n486 0.048
R2100 SS.n489 SS.n488 0.048
R2101 SS.n641 SS.n516 0.048
R2102 SS.n643 SS.n642 0.048
R2103 SS.n426 SS.n425 0.048
R2104 SS.n326 SS.n325 0.048
R2105 SS.n328 SS.n327 0.048
R2106 SS.n480 SS.n355 0.048
R2107 SS.n482 SS.n481 0.048
R2108 SS.n265 SS.n264 0.048
R2109 SS.n165 SS.n164 0.048
R2110 SS.n167 SS.n166 0.048
R2111 SS.n319 SS.n194 0.048
R2112 SS.n321 SS.n320 0.048
R2113 SS.n104 SS.n103 0.048
R2114 SS.n4 SS.n3 0.048
R2115 SS.n6 SS.n5 0.048
R2116 SS.n158 SS.n33 0.048
R2117 SS.n160 SS.n159 0.048
R2118 SS.n1298 SS.n1135 0.048
R2119 SS.n752 SS.n751 0.048
R2120 SS.n652 SS.n651 0.048
R2121 SS.n654 SS.n653 0.048
R2122 SS.n806 SS.n681 0.048
R2123 SS.n808 SS.n807 0.048
R2124 SS.n913 SS.n912 0.048
R2125 SS.n813 SS.n812 0.048
R2126 SS.n815 SS.n814 0.048
R2127 SS.n967 SS.n842 0.048
R2128 SS.n969 SS.n968 0.048
R2129 SS.n1240 SS.n1239 0.048
R2130 SS.n1140 SS.n1139 0.048
R2131 SS.n1142 SS.n1141 0.048
R2132 SS.n1294 SS.n1169 0.048
R2133 SS.n1296 SS.n1295 0.048
R2134 SS.n975 SS.n974 0.048
R2135 SS.n977 SS.n976 0.048
R2136 SS.n1129 SS.n1004 0.048
R2137 SS.n1131 SS.n1130 0.048
R2138 SS.n1078 SS.n1076 0.045
R2139 SS.n590 SS.n588 0.045
R2140 SS.n485 SS.n484 0.045
R2141 SS.n505 SS.n504 0.045
R2142 SS.n513 SS.n512 0.045
R2143 SS.n515 SS.n514 0.045
R2144 SS.n429 SS.n427 0.045
R2145 SS.n324 SS.n323 0.045
R2146 SS.n344 SS.n343 0.045
R2147 SS.n352 SS.n351 0.045
R2148 SS.n354 SS.n353 0.045
R2149 SS.n268 SS.n266 0.045
R2150 SS.n163 SS.n162 0.045
R2151 SS.n183 SS.n182 0.045
R2152 SS.n191 SS.n190 0.045
R2153 SS.n193 SS.n192 0.045
R2154 SS.n107 SS.n105 0.045
R2155 SS.n2 SS.n1 0.045
R2156 SS.n22 SS.n21 0.045
R2157 SS.n30 SS.n29 0.045
R2158 SS.n32 SS.n31 0.045
R2159 SS.n755 SS.n753 0.045
R2160 SS.n650 SS.n649 0.045
R2161 SS.n670 SS.n669 0.045
R2162 SS.n678 SS.n677 0.045
R2163 SS.n680 SS.n679 0.045
R2164 SS.n916 SS.n914 0.045
R2165 SS.n811 SS.n810 0.045
R2166 SS.n831 SS.n830 0.045
R2167 SS.n839 SS.n838 0.045
R2168 SS.n841 SS.n840 0.045
R2169 SS.n1243 SS.n1241 0.045
R2170 SS.n1138 SS.n1137 0.045
R2171 SS.n1158 SS.n1157 0.045
R2172 SS.n1166 SS.n1165 0.045
R2173 SS.n1168 SS.n1167 0.045
R2174 SS.n973 SS.n972 0.045
R2175 SS.n993 SS.n992 0.045
R2176 SS.n1001 SS.n1000 0.045
R2177 SS.n1003 SS.n1002 0.045
R2178 SS.n1008 SS.n1006 0.043
R2179 SS.n1052 SS.n1051 0.043
R2180 SS.n520 SS.n518 0.043
R2181 SS.n564 SS.n563 0.043
R2182 SS.n497 SS.n496 0.043
R2183 SS.n359 SS.n357 0.043
R2184 SS.n403 SS.n402 0.043
R2185 SS.n336 SS.n335 0.043
R2186 SS.n198 SS.n196 0.043
R2187 SS.n242 SS.n241 0.043
R2188 SS.n175 SS.n174 0.043
R2189 SS.n37 SS.n35 0.043
R2190 SS.n81 SS.n80 0.043
R2191 SS.n14 SS.n13 0.043
R2192 SS.n685 SS.n683 0.043
R2193 SS.n729 SS.n728 0.043
R2194 SS.n662 SS.n661 0.043
R2195 SS.n846 SS.n844 0.043
R2196 SS.n890 SS.n889 0.043
R2197 SS.n823 SS.n822 0.043
R2198 SS.n1173 SS.n1171 0.043
R2199 SS.n1217 SS.n1216 0.043
R2200 SS.n1150 SS.n1149 0.043
R2201 SS.n985 SS.n984 0.043
R2202 SS.n1040 SS.n1038 0.04
R2203 SS.n1126 SS.n1124 0.04
R2204 SS.n552 SS.n550 0.04
R2205 SS.n638 SS.n636 0.04
R2206 SS.n391 SS.n389 0.04
R2207 SS.n477 SS.n475 0.04
R2208 SS.n230 SS.n228 0.04
R2209 SS.n316 SS.n314 0.04
R2210 SS.n69 SS.n67 0.04
R2211 SS.n155 SS.n153 0.04
R2212 SS.n717 SS.n715 0.04
R2213 SS.n803 SS.n801 0.04
R2214 SS.n878 SS.n876 0.04
R2215 SS.n964 SS.n962 0.04
R2216 SS.n1205 SS.n1203 0.04
R2217 SS.n1291 SS.n1289 0.04
R2218 SS.n1035 SS.n1034 0.038
R2219 SS.n1093 SS.n1091 0.038
R2220 SS.n547 SS.n546 0.038
R2221 SS.n605 SS.n603 0.038
R2222 SS.n492 SS.n491 0.038
R2223 SS.n386 SS.n385 0.038
R2224 SS.n444 SS.n442 0.038
R2225 SS.n331 SS.n330 0.038
R2226 SS.n225 SS.n224 0.038
R2227 SS.n283 SS.n281 0.038
R2228 SS.n170 SS.n169 0.038
R2229 SS.n64 SS.n63 0.038
R2230 SS.n122 SS.n120 0.038
R2231 SS.n9 SS.n8 0.038
R2232 SS.n712 SS.n711 0.038
R2233 SS.n770 SS.n768 0.038
R2234 SS.n657 SS.n656 0.038
R2235 SS.n873 SS.n872 0.038
R2236 SS.n931 SS.n929 0.038
R2237 SS.n818 SS.n817 0.038
R2238 SS.n1200 SS.n1199 0.038
R2239 SS.n1258 SS.n1256 0.038
R2240 SS.n1145 SS.n1144 0.038
R2241 SS.n980 SS.n979 0.038
R2242 SS.n1089 SS.n1087 0.036
R2243 SS.n1098 SS.n1097 0.036
R2244 SS.n1110 SS.n1108 0.036
R2245 SS.n601 SS.n599 0.036
R2246 SS.n610 SS.n609 0.036
R2247 SS.n622 SS.n620 0.036
R2248 SS.n508 SS.n507 0.036
R2249 SS.n510 SS.n509 0.036
R2250 SS.n440 SS.n438 0.036
R2251 SS.n449 SS.n448 0.036
R2252 SS.n461 SS.n459 0.036
R2253 SS.n347 SS.n346 0.036
R2254 SS.n349 SS.n348 0.036
R2255 SS.n279 SS.n277 0.036
R2256 SS.n288 SS.n287 0.036
R2257 SS.n300 SS.n298 0.036
R2258 SS.n186 SS.n185 0.036
R2259 SS.n188 SS.n187 0.036
R2260 SS.n118 SS.n116 0.036
R2261 SS.n127 SS.n126 0.036
R2262 SS.n139 SS.n137 0.036
R2263 SS.n25 SS.n24 0.036
R2264 SS.n27 SS.n26 0.036
R2265 SS.n766 SS.n764 0.036
R2266 SS.n775 SS.n774 0.036
R2267 SS.n787 SS.n785 0.036
R2268 SS.n673 SS.n672 0.036
R2269 SS.n675 SS.n674 0.036
R2270 SS.n927 SS.n925 0.036
R2271 SS.n936 SS.n935 0.036
R2272 SS.n948 SS.n946 0.036
R2273 SS.n834 SS.n833 0.036
R2274 SS.n836 SS.n835 0.036
R2275 SS.n1254 SS.n1252 0.036
R2276 SS.n1263 SS.n1262 0.036
R2277 SS.n1275 SS.n1273 0.036
R2278 SS.n1161 SS.n1160 0.036
R2279 SS.n1163 SS.n1162 0.036
R2280 SS.n996 SS.n995 0.036
R2281 SS.n998 SS.n997 0.036
R2282 SS.n1024 SS.n1023 0.033
R2283 SS.n1041 SS.n1040 0.033
R2284 SS.n536 SS.n535 0.033
R2285 SS.n553 SS.n552 0.033
R2286 SS.n494 SS.n493 0.033
R2287 SS.n375 SS.n374 0.033
R2288 SS.n392 SS.n391 0.033
R2289 SS.n333 SS.n332 0.033
R2290 SS.n214 SS.n213 0.033
R2291 SS.n231 SS.n230 0.033
R2292 SS.n172 SS.n171 0.033
R2293 SS.n53 SS.n52 0.033
R2294 SS.n70 SS.n69 0.033
R2295 SS.n11 SS.n10 0.033
R2296 SS.n701 SS.n700 0.033
R2297 SS.n718 SS.n717 0.033
R2298 SS.n659 SS.n658 0.033
R2299 SS.n862 SS.n861 0.033
R2300 SS.n879 SS.n878 0.033
R2301 SS.n820 SS.n819 0.033
R2302 SS.n1189 SS.n1188 0.033
R2303 SS.n1206 SS.n1205 0.033
R2304 SS.n1147 SS.n1146 0.033
R2305 SS.n982 SS.n981 0.033
R2306 SS.n1069 SS.n1067 0.031
R2307 SS.n1074 SS.n1071 0.031
R2308 SS.n581 SS.n579 0.031
R2309 SS.n586 SS.n583 0.031
R2310 SS.n420 SS.n418 0.031
R2311 SS.n425 SS.n422 0.031
R2312 SS.n259 SS.n257 0.031
R2313 SS.n264 SS.n261 0.031
R2314 SS.n98 SS.n96 0.031
R2315 SS.n103 SS.n100 0.031
R2316 SS.n746 SS.n744 0.031
R2317 SS.n751 SS.n748 0.031
R2318 SS.n907 SS.n905 0.031
R2319 SS.n912 SS.n909 0.031
R2320 SS.n1234 SS.n1232 0.031
R2321 SS.n1239 SS.n1236 0.031
R2322 SS.n1018 SS.n1015 0.028
R2323 SS.n1042 SS.n1041 0.028
R2324 SS.n1058 SS.n1056 0.028
R2325 SS.n1062 SS.n1060 0.028
R2326 SS.n1104 SS.n1102 0.028
R2327 SS.n530 SS.n527 0.028
R2328 SS.n554 SS.n553 0.028
R2329 SS.n570 SS.n568 0.028
R2330 SS.n574 SS.n572 0.028
R2331 SS.n616 SS.n614 0.028
R2332 SS.n495 SS.n494 0.028
R2333 SS.n369 SS.n366 0.028
R2334 SS.n393 SS.n392 0.028
R2335 SS.n409 SS.n407 0.028
R2336 SS.n413 SS.n411 0.028
R2337 SS.n455 SS.n453 0.028
R2338 SS.n334 SS.n333 0.028
R2339 SS.n208 SS.n205 0.028
R2340 SS.n232 SS.n231 0.028
R2341 SS.n248 SS.n246 0.028
R2342 SS.n252 SS.n250 0.028
R2343 SS.n294 SS.n292 0.028
R2344 SS.n173 SS.n172 0.028
R2345 SS.n47 SS.n44 0.028
R2346 SS.n71 SS.n70 0.028
R2347 SS.n87 SS.n85 0.028
R2348 SS.n91 SS.n89 0.028
R2349 SS.n133 SS.n131 0.028
R2350 SS.n12 SS.n11 0.028
R2351 SS.n695 SS.n692 0.028
R2352 SS.n719 SS.n718 0.028
R2353 SS.n735 SS.n733 0.028
R2354 SS.n739 SS.n737 0.028
R2355 SS.n781 SS.n779 0.028
R2356 SS.n660 SS.n659 0.028
R2357 SS.n856 SS.n853 0.028
R2358 SS.n880 SS.n879 0.028
R2359 SS.n896 SS.n894 0.028
R2360 SS.n900 SS.n898 0.028
R2361 SS.n942 SS.n940 0.028
R2362 SS.n821 SS.n820 0.028
R2363 SS.n1183 SS.n1180 0.028
R2364 SS.n1207 SS.n1206 0.028
R2365 SS.n1223 SS.n1221 0.028
R2366 SS.n1227 SS.n1225 0.028
R2367 SS.n1269 SS.n1267 0.028
R2368 SS.n1148 SS.n1147 0.028
R2369 SS.n983 SS.n982 0.028
R2370 SS.n1013 SS.n1011 0.026
R2371 SS.n1031 SS.n1029 0.026
R2372 SS.n1049 SS.n1047 0.026
R2373 SS.n1087 SS.n1086 0.026
R2374 SS.n1117 SS.n1116 0.026
R2375 SS.n1128 SS.n1120 0.026
R2376 SS.n525 SS.n523 0.026
R2377 SS.n543 SS.n541 0.026
R2378 SS.n561 SS.n559 0.026
R2379 SS.n599 SS.n598 0.026
R2380 SS.n629 SS.n628 0.026
R2381 SS.n640 SS.n632 0.026
R2382 SS.n507 SS.n506 0.026
R2383 SS.n511 SS.n510 0.026
R2384 SS.n364 SS.n362 0.026
R2385 SS.n382 SS.n380 0.026
R2386 SS.n400 SS.n398 0.026
R2387 SS.n438 SS.n437 0.026
R2388 SS.n468 SS.n467 0.026
R2389 SS.n479 SS.n471 0.026
R2390 SS.n346 SS.n345 0.026
R2391 SS.n350 SS.n349 0.026
R2392 SS.n203 SS.n201 0.026
R2393 SS.n221 SS.n219 0.026
R2394 SS.n239 SS.n237 0.026
R2395 SS.n277 SS.n276 0.026
R2396 SS.n307 SS.n306 0.026
R2397 SS.n318 SS.n310 0.026
R2398 SS.n185 SS.n184 0.026
R2399 SS.n189 SS.n188 0.026
R2400 SS.n42 SS.n40 0.026
R2401 SS.n60 SS.n58 0.026
R2402 SS.n78 SS.n76 0.026
R2403 SS.n116 SS.n115 0.026
R2404 SS.n146 SS.n145 0.026
R2405 SS.n157 SS.n149 0.026
R2406 SS.n24 SS.n23 0.026
R2407 SS.n28 SS.n27 0.026
R2408 SS.n690 SS.n688 0.026
R2409 SS.n708 SS.n706 0.026
R2410 SS.n726 SS.n724 0.026
R2411 SS.n764 SS.n763 0.026
R2412 SS.n794 SS.n793 0.026
R2413 SS.n805 SS.n797 0.026
R2414 SS.n672 SS.n671 0.026
R2415 SS.n676 SS.n675 0.026
R2416 SS.n851 SS.n849 0.026
R2417 SS.n869 SS.n867 0.026
R2418 SS.n887 SS.n885 0.026
R2419 SS.n925 SS.n924 0.026
R2420 SS.n955 SS.n954 0.026
R2421 SS.n966 SS.n958 0.026
R2422 SS.n833 SS.n832 0.026
R2423 SS.n837 SS.n836 0.026
R2424 SS.n1178 SS.n1176 0.026
R2425 SS.n1196 SS.n1194 0.026
R2426 SS.n1214 SS.n1212 0.026
R2427 SS.n1252 SS.n1251 0.026
R2428 SS.n1282 SS.n1281 0.026
R2429 SS.n1293 SS.n1285 0.026
R2430 SS.n1160 SS.n1159 0.026
R2431 SS.n1164 SS.n1163 0.026
R2432 SS.n995 SS.n994 0.026
R2433 SS.n999 SS.n998 0.026
R2434 SS.n1082 SS.n1080 0.024
R2435 SS.n594 SS.n592 0.024
R2436 SS.n491 SS.n490 0.024
R2437 SS.n433 SS.n431 0.024
R2438 SS.n330 SS.n329 0.024
R2439 SS.n272 SS.n270 0.024
R2440 SS.n169 SS.n168 0.024
R2441 SS.n111 SS.n109 0.024
R2442 SS.n8 SS.n7 0.024
R2443 SS.n759 SS.n757 0.024
R2444 SS.n656 SS.n655 0.024
R2445 SS.n920 SS.n918 0.024
R2446 SS.n817 SS.n816 0.024
R2447 SS.n1247 SS.n1245 0.024
R2448 SS.n1144 SS.n1143 0.024
R2449 SS.n979 SS.n978 0.024
R2450 SS.n1120 SS.n1118 0.021
R2451 SS.n632 SS.n630 0.021
R2452 SS.n471 SS.n469 0.021
R2453 SS.n310 SS.n308 0.021
R2454 SS.n149 SS.n147 0.021
R2455 SS.n797 SS.n795 0.021
R2456 SS.n958 SS.n956 0.021
R2457 SS.n1285 SS.n1283 0.021
R2458 SS.n1014 SS.n1013 0.019
R2459 SS.n1020 SS.n1018 0.019
R2460 SS.n1053 SS.n1052 0.019
R2461 SS.n1116 SS.n1113 0.019
R2462 SS.n526 SS.n525 0.019
R2463 SS.n532 SS.n530 0.019
R2464 SS.n565 SS.n564 0.019
R2465 SS.n628 SS.n625 0.019
R2466 SS.n498 SS.n497 0.019
R2467 SS.n365 SS.n364 0.019
R2468 SS.n371 SS.n369 0.019
R2469 SS.n404 SS.n403 0.019
R2470 SS.n467 SS.n464 0.019
R2471 SS.n337 SS.n336 0.019
R2472 SS.n204 SS.n203 0.019
R2473 SS.n210 SS.n208 0.019
R2474 SS.n243 SS.n242 0.019
R2475 SS.n306 SS.n303 0.019
R2476 SS.n176 SS.n175 0.019
R2477 SS.n43 SS.n42 0.019
R2478 SS.n49 SS.n47 0.019
R2479 SS.n82 SS.n81 0.019
R2480 SS.n145 SS.n142 0.019
R2481 SS.n15 SS.n14 0.019
R2482 SS.n691 SS.n690 0.019
R2483 SS.n697 SS.n695 0.019
R2484 SS.n730 SS.n729 0.019
R2485 SS.n793 SS.n790 0.019
R2486 SS.n663 SS.n662 0.019
R2487 SS.n852 SS.n851 0.019
R2488 SS.n858 SS.n856 0.019
R2489 SS.n891 SS.n890 0.019
R2490 SS.n954 SS.n951 0.019
R2491 SS.n824 SS.n823 0.019
R2492 SS.n1179 SS.n1178 0.019
R2493 SS.n1185 SS.n1183 0.019
R2494 SS.n1218 SS.n1217 0.019
R2495 SS.n1281 SS.n1278 0.019
R2496 SS.n1151 SS.n1150 0.019
R2497 SS.n986 SS.n985 0.019
R2498 SS.n1076 SS.n1075 0.016
R2499 SS.n1080 SS.n1078 0.016
R2500 SS.n1085 SS.n1082 0.016
R2501 SS.n588 SS.n587 0.016
R2502 SS.n592 SS.n590 0.016
R2503 SS.n597 SS.n594 0.016
R2504 SS.n504 SS.n503 0.016
R2505 SS.n427 SS.n426 0.016
R2506 SS.n431 SS.n429 0.016
R2507 SS.n436 SS.n433 0.016
R2508 SS.n343 SS.n342 0.016
R2509 SS.n266 SS.n265 0.016
R2510 SS.n270 SS.n268 0.016
R2511 SS.n275 SS.n272 0.016
R2512 SS.n182 SS.n181 0.016
R2513 SS.n105 SS.n104 0.016
R2514 SS.n109 SS.n107 0.016
R2515 SS.n114 SS.n111 0.016
R2516 SS.n21 SS.n20 0.016
R2517 SS.n753 SS.n752 0.016
R2518 SS.n757 SS.n755 0.016
R2519 SS.n762 SS.n759 0.016
R2520 SS.n669 SS.n668 0.016
R2521 SS.n914 SS.n913 0.016
R2522 SS.n918 SS.n916 0.016
R2523 SS.n923 SS.n920 0.016
R2524 SS.n830 SS.n829 0.016
R2525 SS.n1241 SS.n1240 0.016
R2526 SS.n1245 SS.n1243 0.016
R2527 SS.n1250 SS.n1247 0.016
R2528 SS.n1157 SS.n1156 0.016
R2529 SS.n992 SS.n991 0.016
R2530 SS.n1023 SS.n1021 0.014
R2531 SS.n1029 SS.n1027 0.014
R2532 SS.n1033 SS.n1031 0.014
R2533 SS.n1047 SS.n1045 0.014
R2534 SS.n1051 SS.n1049 0.014
R2535 SS.n1100 SS.n1098 0.014
R2536 SS.n535 SS.n533 0.014
R2537 SS.n541 SS.n539 0.014
R2538 SS.n545 SS.n543 0.014
R2539 SS.n559 SS.n557 0.014
R2540 SS.n563 SS.n561 0.014
R2541 SS.n612 SS.n610 0.014
R2542 SS.n374 SS.n372 0.014
R2543 SS.n380 SS.n378 0.014
R2544 SS.n384 SS.n382 0.014
R2545 SS.n398 SS.n396 0.014
R2546 SS.n402 SS.n400 0.014
R2547 SS.n451 SS.n449 0.014
R2548 SS.n213 SS.n211 0.014
R2549 SS.n219 SS.n217 0.014
R2550 SS.n223 SS.n221 0.014
R2551 SS.n237 SS.n235 0.014
R2552 SS.n241 SS.n239 0.014
R2553 SS.n290 SS.n288 0.014
R2554 SS.n52 SS.n50 0.014
R2555 SS.n58 SS.n56 0.014
R2556 SS.n62 SS.n60 0.014
R2557 SS.n76 SS.n74 0.014
R2558 SS.n80 SS.n78 0.014
R2559 SS.n129 SS.n127 0.014
R2560 SS.n700 SS.n698 0.014
R2561 SS.n706 SS.n704 0.014
R2562 SS.n710 SS.n708 0.014
R2563 SS.n724 SS.n722 0.014
R2564 SS.n728 SS.n726 0.014
R2565 SS.n777 SS.n775 0.014
R2566 SS.n861 SS.n859 0.014
R2567 SS.n867 SS.n865 0.014
R2568 SS.n871 SS.n869 0.014
R2569 SS.n885 SS.n883 0.014
R2570 SS.n889 SS.n887 0.014
R2571 SS.n938 SS.n936 0.014
R2572 SS.n1188 SS.n1186 0.014
R2573 SS.n1194 SS.n1192 0.014
R2574 SS.n1198 SS.n1196 0.014
R2575 SS.n1212 SS.n1210 0.014
R2576 SS.n1216 SS.n1214 0.014
R2577 SS.n1265 SS.n1263 0.014
R2578 SS.n1011 SS.n1009 0.012
R2579 SS.n1060 SS.n1058 0.012
R2580 SS.n1102 SS.n1100 0.012
R2581 SS.n1107 SS.n1104 0.012
R2582 SS.n1113 SS.n1111 0.012
R2583 SS.n523 SS.n521 0.012
R2584 SS.n572 SS.n570 0.012
R2585 SS.n614 SS.n612 0.012
R2586 SS.n619 SS.n616 0.012
R2587 SS.n625 SS.n623 0.012
R2588 SS.n484 SS.n483 0.012
R2589 SS.n514 SS.n513 0.012
R2590 SS.n362 SS.n360 0.012
R2591 SS.n411 SS.n409 0.012
R2592 SS.n453 SS.n451 0.012
R2593 SS.n458 SS.n455 0.012
R2594 SS.n464 SS.n462 0.012
R2595 SS.n323 SS.n322 0.012
R2596 SS.n353 SS.n352 0.012
R2597 SS.n201 SS.n199 0.012
R2598 SS.n250 SS.n248 0.012
R2599 SS.n292 SS.n290 0.012
R2600 SS.n297 SS.n294 0.012
R2601 SS.n303 SS.n301 0.012
R2602 SS.n162 SS.n161 0.012
R2603 SS.n192 SS.n191 0.012
R2604 SS.n40 SS.n38 0.012
R2605 SS.n89 SS.n87 0.012
R2606 SS.n131 SS.n129 0.012
R2607 SS.n136 SS.n133 0.012
R2608 SS.n142 SS.n140 0.012
R2609 SS.n1 SS.n0 0.012
R2610 SS.n31 SS.n30 0.012
R2611 SS.n688 SS.n686 0.012
R2612 SS.n737 SS.n735 0.012
R2613 SS.n779 SS.n777 0.012
R2614 SS.n784 SS.n781 0.012
R2615 SS.n790 SS.n788 0.012
R2616 SS.n649 SS.n648 0.012
R2617 SS.n679 SS.n678 0.012
R2618 SS.n849 SS.n847 0.012
R2619 SS.n898 SS.n896 0.012
R2620 SS.n940 SS.n938 0.012
R2621 SS.n945 SS.n942 0.012
R2622 SS.n951 SS.n949 0.012
R2623 SS.n810 SS.n809 0.012
R2624 SS.n840 SS.n839 0.012
R2625 SS.n1176 SS.n1174 0.012
R2626 SS.n1225 SS.n1223 0.012
R2627 SS.n1267 SS.n1265 0.012
R2628 SS.n1272 SS.n1269 0.012
R2629 SS.n1278 SS.n1276 0.012
R2630 SS.n1137 SS.n1136 0.012
R2631 SS.n1167 SS.n1166 0.012
R2632 SS.n972 SS.n971 0.012
R2633 SS.n1002 SS.n1001 0.012
R2634 SS.n1034 SS.n1033 0.009
R2635 SS.n1071 SS.n1069 0.009
R2636 SS.n1111 SS.n1110 0.009
R2637 SS.n546 SS.n545 0.009
R2638 SS.n583 SS.n581 0.009
R2639 SS.n623 SS.n622 0.009
R2640 SS.n385 SS.n384 0.009
R2641 SS.n422 SS.n420 0.009
R2642 SS.n462 SS.n461 0.009
R2643 SS.n224 SS.n223 0.009
R2644 SS.n261 SS.n259 0.009
R2645 SS.n301 SS.n300 0.009
R2646 SS.n63 SS.n62 0.009
R2647 SS.n100 SS.n98 0.009
R2648 SS.n140 SS.n139 0.009
R2649 SS.n711 SS.n710 0.009
R2650 SS.n748 SS.n746 0.009
R2651 SS.n788 SS.n787 0.009
R2652 SS.n872 SS.n871 0.009
R2653 SS.n909 SS.n907 0.009
R2654 SS.n949 SS.n948 0.009
R2655 SS.n1199 SS.n1198 0.009
R2656 SS.n1236 SS.n1234 0.009
R2657 SS.n1276 SS.n1275 0.009
R2658 SS.n1021 SS.n1020 0.007
R2659 SS.n1128 SS.n1127 0.007
R2660 SS.n1127 SS.n1126 0.007
R2661 SS.n533 SS.n532 0.007
R2662 SS.n640 SS.n639 0.007
R2663 SS.n639 SS.n638 0.007
R2664 SS.n488 SS.n487 0.007
R2665 SS.n642 SS.n641 0.007
R2666 SS.n372 SS.n371 0.007
R2667 SS.n479 SS.n478 0.007
R2668 SS.n478 SS.n477 0.007
R2669 SS.n327 SS.n326 0.007
R2670 SS.n481 SS.n480 0.007
R2671 SS.n211 SS.n210 0.007
R2672 SS.n318 SS.n317 0.007
R2673 SS.n317 SS.n316 0.007
R2674 SS.n166 SS.n165 0.007
R2675 SS.n320 SS.n319 0.007
R2676 SS.n50 SS.n49 0.007
R2677 SS.n157 SS.n156 0.007
R2678 SS.n156 SS.n155 0.007
R2679 SS.n5 SS.n4 0.007
R2680 SS.n159 SS.n158 0.007
R2681 SS.n698 SS.n697 0.007
R2682 SS.n805 SS.n804 0.007
R2683 SS.n804 SS.n803 0.007
R2684 SS.n653 SS.n652 0.007
R2685 SS.n807 SS.n806 0.007
R2686 SS.n859 SS.n858 0.007
R2687 SS.n966 SS.n965 0.007
R2688 SS.n965 SS.n964 0.007
R2689 SS.n814 SS.n813 0.007
R2690 SS.n968 SS.n967 0.007
R2691 SS.n1186 SS.n1185 0.007
R2692 SS.n1293 SS.n1292 0.007
R2693 SS.n1292 SS.n1291 0.007
R2694 SS.n1141 SS.n1140 0.007
R2695 SS.n1295 SS.n1294 0.007
R2696 SS.n976 SS.n975 0.007
R2697 SS.n1130 SS.n1129 0.007
R2698 SS.n1009 SS.n1008 0.002
R2699 SS.n1064 SS.n1063 0.002
R2700 SS.n1091 SS.n1089 0.002
R2701 SS.n1096 SS.n1093 0.002
R2702 SS.n521 SS.n520 0.002
R2703 SS.n576 SS.n575 0.002
R2704 SS.n603 SS.n601 0.002
R2705 SS.n608 SS.n605 0.002
R2706 SS.n501 SS.n500 0.002
R2707 SS.n360 SS.n359 0.002
R2708 SS.n415 SS.n414 0.002
R2709 SS.n442 SS.n440 0.002
R2710 SS.n447 SS.n444 0.002
R2711 SS.n340 SS.n339 0.002
R2712 SS.n199 SS.n198 0.002
R2713 SS.n254 SS.n253 0.002
R2714 SS.n281 SS.n279 0.002
R2715 SS.n286 SS.n283 0.002
R2716 SS.n179 SS.n178 0.002
R2717 SS.n38 SS.n37 0.002
R2718 SS.n93 SS.n92 0.002
R2719 SS.n120 SS.n118 0.002
R2720 SS.n125 SS.n122 0.002
R2721 SS.n18 SS.n17 0.002
R2722 SS.n686 SS.n685 0.002
R2723 SS.n741 SS.n740 0.002
R2724 SS.n768 SS.n766 0.002
R2725 SS.n773 SS.n770 0.002
R2726 SS.n666 SS.n665 0.002
R2727 SS.n847 SS.n846 0.002
R2728 SS.n902 SS.n901 0.002
R2729 SS.n929 SS.n927 0.002
R2730 SS.n934 SS.n931 0.002
R2731 SS.n827 SS.n826 0.002
R2732 SS.n1174 SS.n1173 0.002
R2733 SS.n1229 SS.n1228 0.002
R2734 SS.n1256 SS.n1254 0.002
R2735 SS.n1261 SS.n1258 0.002
R2736 SS.n1154 SS.n1153 0.002
R2737 SS.n989 SS.n988 0.002
R2738 a_n6328_16092.n12 a_n6328_16092.n74 9.3
R2739 a_n6328_16092.n13 a_n6328_16092.n80 9.3
R2740 a_n6328_16092.n6 a_n6328_16092.n87 9.3
R2741 a_n6328_16092.n5 a_n6328_16092.n82 9.3
R2742 a_n6328_16092.n5 a_n6328_16092.n83 9.3
R2743 a_n6328_16092.n101 a_n6328_16092.n100 9.3
R2744 a_n6328_16092.n103 a_n6328_16092.n107 9.3
R2745 a_n6328_16092.n110 a_n6328_16092.n109 9.3
R2746 a_n6328_16092.n10 a_n6328_16092.n112 9.3
R2747 a_n6328_16092.n1 a_n6328_16092.n96 9.3
R2748 a_n6328_16092.n92 a_n6328_16092.n91 9.3
R2749 a_n6328_16092.n90 a_n6328_16092.n89 9.3
R2750 a_n6328_16092.n12 a_n6328_16092.n75 9.3
R2751 a_n6328_16092.n65 a_n6328_16092.n64 9.3
R2752 a_n6328_16092.n14 a_n6328_16092.n47 9.3
R2753 a_n6328_16092.n9 a_n6328_16092.n45 9.3
R2754 a_n6328_16092.n9 a_n6328_16092.n44 9.3
R2755 a_n6328_16092.n14 a_n6328_16092.n48 9.3
R2756 a_n6328_16092.n58 a_n6328_16092.n57 9.3
R2757 a_n6328_16092.n36 a_n6328_16092.n35 9.3
R2758 a_n6328_16092.n31 a_n6328_16092.n30 9.3
R2759 a_n6328_16092.n39 a_n6328_16092.n38 9.3
R2760 a_n6328_16092.n41 a_n6328_16092.n40 9.3
R2761 a_n6328_16092.n11 a_n6328_16092.n111 9
R2762 a_n6328_16092.n104 a_n6328_16092.n102 9
R2763 a_n6328_16092.n97 a_n6328_16092.n93 9
R2764 a_n6328_16092.n6 a_n6328_16092.n88 9
R2765 a_n6328_16092.n13 a_n6328_16092.n81 9
R2766 a_n6328_16092.n76 a_n6328_16092.n73 9
R2767 a_n6328_16092.n66 a_n6328_16092.n63 9
R2768 a_n6328_16092.n114 a_n6328_16092.n113 9
R2769 a_n6328_16092.n50 a_n6328_16092.n49 9
R2770 a_n6328_16092.n118 a_n6328_16092.n25 8.473
R2771 a_n6328_16092.n118 a_n6328_16092.n28 8.096
R2772 a_n6328_16092.n118 a_n6328_16092.n23 8.069
R2773 a_n6328_16092.n118 a_n6328_16092.n20 8.042
R2774 a_n6328_16092.n118 a_n6328_16092.n17 8.016
R2775 a_n6328_16092.n72 a_n6328_16092.n71 4.574
R2776 a_n6328_16092.n55 a_n6328_16092.n54 4.574
R2777 a_n6328_16092.n71 a_n6328_16092.n69 3.388
R2778 a_n6328_16092.n54 a_n6328_16092.n52 3.388
R2779 a_n6328_16092.n59 a_n6328_16092.t2 3.326
R2780 a_n6328_16092.t1 a_n6328_16092.n118 3.326
R2781 a_n6328_16092.n0 a_n6328_16092.n6 3
R2782 a_n6328_16092.n98 a_n6328_16092.n97 3
R2783 a_n6328_16092.n7 a_n6328_16092.n104 3
R2784 a_n6328_16092.n8 a_n6328_16092.n11 3
R2785 a_n6328_16092.n4 a_n6328_16092.n13 3
R2786 a_n6328_16092.n4 a_n6328_16092.n76 3
R2787 a_n6328_16092.n2 a_n6328_16092.n72 3
R2788 a_n6328_16092.n2 a_n6328_16092.n66 3
R2789 a_n6328_16092.n114 a_n6328_16092.n2 3
R2790 a_n6328_16092.n22 a_n6328_16092.n21 2.258
R2791 a_n6328_16092.n27 a_n6328_16092.n26 2.258
R2792 a_n6328_16092.n19 a_n6328_16092.n18 1.505
R2793 a_n6328_16092.n25 a_n6328_16092.n24 1.505
R2794 a_n6328_16092.n118 a_n6328_16092.n117 1.155
R2795 a_n6328_16092.n60 a_n6328_16092.n59 1.155
R2796 a_n6328_16092.n117 a_n6328_16092.n116 0.893
R2797 a_n6328_16092.n61 a_n6328_16092.n60 0.893
R2798 a_n6328_16092.n16 a_n6328_16092.n15 0.752
R2799 a_n6328_16092.n71 a_n6328_16092.n70 0.506
R2800 a_n6328_16092.n54 a_n6328_16092.n53 0.506
R2801 a_n6328_16092.n80 a_n6328_16092.n79 0.476
R2802 a_n6328_16092.n17 a_n6328_16092.n16 0.476
R2803 a_n6328_16092.n87 a_n6328_16092.n86 0.445
R2804 a_n6328_16092.n20 a_n6328_16092.n19 0.445
R2805 a_n6328_16092.n96 a_n6328_16092.n95 0.414
R2806 a_n6328_16092.n23 a_n6328_16092.n22 0.414
R2807 a_n6328_16092.n107 a_n6328_16092.n106 0.382
R2808 a_n6328_16092.n28 a_n6328_16092.n27 0.382
R2809 a_n6328_16092.n8 a_n6328_16092.t0 0.224
R2810 a_n6328_16092.n42 a_n6328_16092.n41 0.06
R2811 a_n6328_16092.n33 a_n6328_16092.n32 0.06
R2812 a_n6328_16092.n72 a_n6328_16092.n68 0.053
R2813 a_n6328_16092.n55 a_n6328_16092.n51 0.053
R2814 a_n6328_16092.n51 a_n6328_16092.n50 0.053
R2815 a_n6328_16092.n66 a_n6328_16092.n62 0.043
R2816 a_n6328_16092.n103 a_n6328_16092.n105 0.043
R2817 a_n6328_16092.n115 a_n6328_16092.n114 0.043
R2818 a_n6328_16092.n34 a_n6328_16092.n33 0.043
R2819 a_n6328_16092.n14 a_n6328_16092.n46 0.091
R2820 a_n6328_16092.n46 a_n6328_16092.n9 0.069
R2821 a_n6328_16092.n13 a_n6328_16092.n78 0.044
R2822 a_n6328_16092.n36 a_n6328_16092.n34 0.04
R2823 a_n6328_16092.n31 a_n6328_16092.n29 0.04
R2824 a_n6328_16092.n1 a_n6328_16092.n94 0.036
R2825 a_n6328_16092.n9 a_n6328_16092.n43 0.066
R2826 a_n6328_16092.n7 a_n6328_16092.n8 0.042
R2827 a_n6328_16092.n6 a_n6328_16092.n5 0.04
R2828 a_n6328_16092.n6 a_n6328_16092.n85 0.035
R2829 a_n6328_16092.n98 a_n6328_16092.n7 0.033
R2830 a_n6328_16092.n2 a_n6328_16092.n4 0.031
R2831 a_n6328_16092.n85 a_n6328_16092.n84 0.026
R2832 a_n6328_16092.n97 a_n6328_16092.n92 0.026
R2833 a_n6328_16092.n104 a_n6328_16092.n101 0.026
R2834 a_n6328_16092.n43 a_n6328_16092.n42 0.026
R2835 a_n6328_16092.n39 a_n6328_16092.n37 0.148
R2836 a_n6328_16092.n3 a_n6328_16092.n0 0.032
R2837 a_n6328_16092.n97 a_n6328_16092.n1 0.026
R2838 a_n6328_16092.n110 a_n6328_16092.n108 0.024
R2839 a_n6328_16092.n11 a_n6328_16092.n110 0.024
R2840 a_n6328_16092.n32 a_n6328_16092.n31 0.024
R2841 a_n6328_16092.n50 a_n6328_16092.n14 0.023
R2842 a_n6328_16092.n76 a_n6328_16092.n12 0.023
R2843 a_n6328_16092.n4 a_n6328_16092.n3 0.023
R2844 a_n6328_16092.n72 a_n6328_16092.n67 0.021
R2845 a_n6328_16092.n56 a_n6328_16092.n55 0.021
R2846 a_n6328_16092.n0 a_n6328_16092.n98 0.02
R2847 a_n6328_16092.n62 a_n6328_16092.n61 0.019
R2848 a_n6328_16092.n101 a_n6328_16092.n99 0.019
R2849 a_n6328_16092.n116 a_n6328_16092.n115 0.019
R2850 a_n6328_16092.n58 a_n6328_16092.n56 0.019
R2851 a_n6328_16092.n37 a_n6328_16092.n36 0.019
R2852 a_n6328_16092.n78 a_n6328_16092.n77 0.016
R2853 a_n6328_16092.n11 a_n6328_16092.n10 0.016
R2854 a_n6328_16092.n104 a_n6328_16092.n103 0.014
R2855 a_n6328_16092.n66 a_n6328_16092.n65 0.014
R2856 a_n6328_16092.n92 a_n6328_16092.n90 0.014
R2857 a_n6328_16092.n114 a_n6328_16092.n58 0.014
R2858 a_n6328_16092.n41 a_n6328_16092.n39 0.014
R2859 a_n5540_16092.n80 a_n5540_16092.n78 9.469
R2860 a_n5540_16092.n6 a_n5540_16092.n67 9.3
R2861 a_n5540_16092.n7 a_n5540_16092.n65 9.3
R2862 a_n5540_16092.n31 a_n5540_16092.n30 9.3
R2863 a_n5540_16092.n2 a_n5540_16092.n41 9.3
R2864 a_n5540_16092.n1 a_n5540_16092.n37 9.3
R2865 a_n5540_16092.n26 a_n5540_16092.n34 9.3
R2866 a_n5540_16092.n36 a_n5540_16092.n35 9.3
R2867 a_n5540_16092.n51 a_n5540_16092.n50 9.3
R2868 a_n5540_16092.n46 a_n5540_16092.n45 9.3
R2869 a_n5540_16092.n44 a_n5540_16092.n43 9.3
R2870 a_n5540_16092.n1 a_n5540_16092.n38 9.3
R2871 a_n5540_16092.n0 a_n5540_16092.n29 9.3
R2872 a_n5540_16092.n6 a_n5540_16092.n68 9.3
R2873 a_n5540_16092.n59 a_n5540_16092.n58 9.3
R2874 a_n5540_16092.n8 a_n5540_16092.n90 9.3
R2875 a_n5540_16092.n3 a_n5540_16092.n89 9.3
R2876 a_n5540_16092.n3 a_n5540_16092.n88 9.3
R2877 a_n5540_16092.n80 a_n5540_16092.n79 9.3
R2878 a_n5540_16092.n85 a_n5540_16092.n84 9.3
R2879 a_n5540_16092.n87 a_n5540_16092.n86 9.3
R2880 a_n5540_16092.n8 a_n5540_16092.n91 9.3
R2881 a_n5540_16092.n101 a_n5540_16092.n100 9.3
R2882 a_n5540_16092.n48 a_n5540_16092.n47 9
R2883 a_n5540_16092.n27 a_n5540_16092.n25 9
R2884 a_n5540_16092.n2 a_n5540_16092.n39 9
R2885 a_n5540_16092.n0 a_n5540_16092.n28 9
R2886 a_n5540_16092.n7 a_n5540_16092.n66 9
R2887 a_n5540_16092.n69 a_n5540_16092.n62 9
R2888 a_n5540_16092.n60 a_n5540_16092.n57 9
R2889 a_n5540_16092.n103 a_n5540_16092.n102 9
R2890 a_n5540_16092.n93 a_n5540_16092.n92 9
R2891 a_n5540_16092.n106 a_n5540_16092.n22 8.474
R2892 a_n5540_16092.n106 a_n5540_16092.n20 8.096
R2893 a_n5540_16092.n106 a_n5540_16092.n17 8.069
R2894 a_n5540_16092.n106 a_n5540_16092.n14 8.042
R2895 a_n5540_16092.n106 a_n5540_16092.n11 8.016
R2896 a_n5540_16092.n74 a_n5540_16092.n73 4.574
R2897 a_n5540_16092.n98 a_n5540_16092.n97 4.574
R2898 a_n5540_16092.n73 a_n5540_16092.n71 3.388
R2899 a_n5540_16092.n97 a_n5540_16092.n95 3.388
R2900 a_n5540_16092.n55 a_n5540_16092.t2 3.326
R2901 a_n5540_16092.t1 a_n5540_16092.n106 3.326
R2902 a_n5540_16092.n54 a_n5540_16092.n75 2.989
R2903 a_n5540_16092.n54 a_n5540_16092.n61 2.987
R2904 a_n5540_16092.n104 a_n5540_16092.n24 2.987
R2905 a_n5540_16092.n5 a_n5540_16092.n52 2.979
R2906 a_n5540_16092.n16 a_n5540_16092.n15 2.258
R2907 a_n5540_16092.n19 a_n5540_16092.n18 2.258
R2908 a_n5540_16092.n13 a_n5540_16092.n12 1.505
R2909 a_n5540_16092.n22 a_n5540_16092.n21 1.505
R2910 a_n5540_16092.n106 a_n5540_16092.n105 1.155
R2911 a_n5540_16092.n56 a_n5540_16092.n55 1.155
R2912 a_n5540_16092.n105 a_n5540_16092.n104 0.921
R2913 a_n5540_16092.n61 a_n5540_16092.n56 0.921
R2914 a_n5540_16092.n10 a_n5540_16092.n9 0.752
R2915 a_n5540_16092.n73 a_n5540_16092.n72 0.506
R2916 a_n5540_16092.n97 a_n5540_16092.n96 0.506
R2917 a_n5540_16092.n65 a_n5540_16092.n64 0.476
R2918 a_n5540_16092.n11 a_n5540_16092.n10 0.476
R2919 a_n5540_16092.n41 a_n5540_16092.n40 0.445
R2920 a_n5540_16092.n14 a_n5540_16092.n13 0.445
R2921 a_n5540_16092.n50 a_n5540_16092.n49 0.414
R2922 a_n5540_16092.n17 a_n5540_16092.n16 0.414
R2923 a_n5540_16092.n34 a_n5540_16092.n33 0.382
R2924 a_n5540_16092.n20 a_n5540_16092.n19 0.382
R2925 a_n5540_16092.n8 a_n5540_16092.n3 0.161
R2926 a_n5540_16092.n4 a_n5540_16092.t0 0.119
R2927 a_n5540_16092.n44 a_n5540_16092.n42 0.073
R2928 a_n5540_16092.n3 a_n5540_16092.n87 0.153
R2929 a_n5540_16092.n26 a_n5540_16092.n32 0.073
R2930 a_n5540_16092.n52 a_n5540_16092.n36 0.072
R2931 a_n5540_16092.n81 a_n5540_16092.n80 0.072
R2932 a_n5540_16092.n75 a_n5540_16092.n69 0.071
R2933 a_n5540_16092.n94 a_n5540_16092.n93 0.071
R2934 a_n5540_16092.n52 a_n5540_16092.n51 0.057
R2935 a_n5540_16092.n82 a_n5540_16092.n81 0.057
R2936 a_n5540_16092.n76 a_n5540_16092.n54 0.056
R2937 a_n5540_16092.n32 a_n5540_16092.n31 0.054
R2938 a_n5540_16092.n2 a_n5540_16092.n1 0.049
R2939 a_n5540_16092.n7 a_n5540_16092.n63 0.048
R2940 a_n5540_16092.n31 a_n5540_16092.n0 0.041
R2941 a_n5540_16092.n42 a_n5540_16092.n2 0.039
R2942 a_n5540_16092.n23 a_n5540_16092.n76 0.038
R2943 a_n5540_16092.n76 a_n5540_16092.n107 0.037
R2944 a_n5540_16092.n75 a_n5540_16092.n74 0.036
R2945 a_n5540_16092.n98 a_n5540_16092.n94 0.036
R2946 a_n5540_16092.n61 a_n5540_16092.n60 0.036
R2947 a_n5540_16092.n104 a_n5540_16092.n103 0.036
R2948 a_n5540_16092.n6 a_n5540_16092.n7 0.035
R2949 a_n5540_16092.n48 a_n5540_16092.n46 0.026
R2950 a_n5540_16092.n36 a_n5540_16092.n27 0.026
R2951 a_n5540_16092.n85 a_n5540_16092.n83 0.026
R2952 a_n5540_16092.n76 a_n5540_16092.n5 0.023
R2953 a_n5540_16092.n93 a_n5540_16092.n8 0.023
R2954 a_n5540_16092.n69 a_n5540_16092.n6 0.023
R2955 a_n5540_16092.n74 a_n5540_16092.n70 0.021
R2956 a_n5540_16092.n99 a_n5540_16092.n98 0.021
R2957 a_n5540_16092.n101 a_n5540_16092.n99 0.019
R2958 a_n5540_16092.n5 a_n5540_16092.n4 0.016
R2959 a_n5540_16092.n27 a_n5540_16092.n26 0.015
R2960 a_n5540_16092.n60 a_n5540_16092.n59 0.014
R2961 a_n5540_16092.n46 a_n5540_16092.n44 0.014
R2962 a_n5540_16092.n51 a_n5540_16092.n48 0.014
R2963 a_n5540_16092.n103 a_n5540_16092.n101 0.014
R2964 a_n5540_16092.n87 a_n5540_16092.n85 0.014
R2965 a_n5540_16092.n83 a_n5540_16092.n82 0.014
R2966 a_n5540_16092.n54 a_n5540_16092.n53 0.014
R2967 a_n5540_16092.n24 a_n5540_16092.n23 0.014
R2968 a_n5540_16092.n24 a_n5540_16092.n77 0.014
R2969 a_n6722_16092.n24 a_n6722_16092.n22 9.468
R2970 a_n6722_16092.n5 a_n6722_16092.n75 9.3
R2971 a_n6722_16092.n6 a_n6722_16092.n73 9.3
R2972 a_n6722_16092.n1 a_n6722_16092.n33 9.3
R2973 a_n6722_16092.n1 a_n6722_16092.n34 9.3
R2974 a_n6722_16092.n2 a_n6722_16092.n37 9.3
R2975 a_n6722_16092.n5 a_n6722_16092.n76 9.3
R2976 a_n6722_16092.n65 a_n6722_16092.n64 9.3
R2977 a_n6722_16092.n59 a_n6722_16092.n58 9.3
R2978 a_n6722_16092.n49 a_n6722_16092.n57 9.3
R2979 a_n6722_16092.n54 a_n6722_16092.n53 9.3
R2980 a_n6722_16092.n0 a_n6722_16092.n52 9.3
R2981 a_n6722_16092.n47 a_n6722_16092.n46 9.3
R2982 a_n6722_16092.n42 a_n6722_16092.n41 9.3
R2983 a_n6722_16092.n40 a_n6722_16092.n39 9.3
R2984 a_n6722_16092.n7 a_n6722_16092.n29 9.3
R2985 a_n6722_16092.n3 a_n6722_16092.n28 9.3
R2986 a_n6722_16092.n3 a_n6722_16092.n27 9.3
R2987 a_n6722_16092.n24 a_n6722_16092.n23 9.3
R2988 a_n6722_16092.n26 a_n6722_16092.n25 9.3
R2989 a_n6722_16092.n7 a_n6722_16092.n30 9.3
R2990 a_n6722_16092.n92 a_n6722_16092.n91 9.3
R2991 a_n6722_16092.n0 a_n6722_16092.n51 9
R2992 a_n6722_16092.n50 a_n6722_16092.n48 9
R2993 a_n6722_16092.n44 a_n6722_16092.n43 9
R2994 a_n6722_16092.n2 a_n6722_16092.n35 9
R2995 a_n6722_16092.n66 a_n6722_16092.n63 9
R2996 a_n6722_16092.n6 a_n6722_16092.n74 9
R2997 a_n6722_16092.n77 a_n6722_16092.n70 9
R2998 a_n6722_16092.n32 a_n6722_16092.n31 9
R2999 a_n6722_16092.n94 a_n6722_16092.n93 9
R3000 a_n6722_16092.n97 a_n6722_16092.n15 8.473
R3001 a_n6722_16092.n97 a_n6722_16092.n18 8.096
R3002 a_n6722_16092.n97 a_n6722_16092.n13 8.069
R3003 a_n6722_16092.n97 a_n6722_16092.n21 8.043
R3004 a_n6722_16092.n97 a_n6722_16092.n10 8.016
R3005 a_n6722_16092.n82 a_n6722_16092.n81 4.574
R3006 a_n6722_16092.n89 a_n6722_16092.n88 4.574
R3007 a_n6722_16092.n81 a_n6722_16092.n79 3.388
R3008 a_n6722_16092.n88 a_n6722_16092.n86 3.388
R3009 a_n6722_16092.n67 a_n6722_16092.t2 3.326
R3010 a_n6722_16092.t1 a_n6722_16092.n97 3.326
R3011 a_n6722_16092.n62 a_n6722_16092.n83 2.989
R3012 a_n6722_16092.n62 a_n6722_16092.n69 2.987
R3013 a_n6722_16092.n4 a_n6722_16092.n60 2.979
R3014 a_n6722_16092.n85 a_n6722_16092.n84 2.286
R3015 a_n6722_16092.n12 a_n6722_16092.n11 2.258
R3016 a_n6722_16092.n17 a_n6722_16092.n16 2.258
R3017 a_n6722_16092.n20 a_n6722_16092.n19 1.505
R3018 a_n6722_16092.n15 a_n6722_16092.n14 1.505
R3019 a_n6722_16092.n68 a_n6722_16092.n67 1.155
R3020 a_n6722_16092.n97 a_n6722_16092.n96 1.155
R3021 a_n6722_16092.n69 a_n6722_16092.n68 0.921
R3022 a_n6722_16092.n96 a_n6722_16092.n95 0.903
R3023 a_n6722_16092.n9 a_n6722_16092.n8 0.752
R3024 a_n6722_16092.n81 a_n6722_16092.n80 0.506
R3025 a_n6722_16092.n88 a_n6722_16092.n87 0.506
R3026 a_n6722_16092.n73 a_n6722_16092.n72 0.476
R3027 a_n6722_16092.n10 a_n6722_16092.n9 0.476
R3028 a_n6722_16092.n21 a_n6722_16092.n20 0.445
R3029 a_n6722_16092.n37 a_n6722_16092.n36 0.445
R3030 a_n6722_16092.n46 a_n6722_16092.n45 0.414
R3031 a_n6722_16092.n13 a_n6722_16092.n12 0.413
R3032 a_n6722_16092.n57 a_n6722_16092.n56 0.382
R3033 a_n6722_16092.n18 a_n6722_16092.n17 0.382
R3034 a_n6722_16092.n7 a_n6722_16092.n3 0.161
R3035 a_n6722_16092.n4 a_n6722_16092.t0 0.135
R3036 a_n6722_16092.n40 a_n6722_16092.n38 0.073
R3037 a_n6722_16092.n3 a_n6722_16092.n26 0.153
R3038 a_n6722_16092.n49 a_n6722_16092.n55 0.073
R3039 a_n6722_16092.n60 a_n6722_16092.n59 0.072
R3040 a_n6722_16092.n83 a_n6722_16092.n77 0.071
R3041 a_n6722_16092.n60 a_n6722_16092.n47 0.057
R3042 a_n6722_16092.n55 a_n6722_16092.n54 0.054
R3043 a_n6722_16092.n89 a_n6722_16092.n85 0.054
R3044 a_n6722_16092.n85 a_n6722_16092.n32 0.054
R3045 a_n6722_16092.n84 a_n6722_16092.n62 0.053
R3046 a_n6722_16092.n95 a_n6722_16092.n94 0.053
R3047 a_n6722_16092.n2 a_n6722_16092.n1 0.049
R3048 a_n6722_16092.n6 a_n6722_16092.n71 0.048
R3049 a_n6722_16092.n54 a_n6722_16092.n0 0.041
R3050 a_n6722_16092.n38 a_n6722_16092.n2 0.039
R3051 a_n6722_16092.n83 a_n6722_16092.n82 0.036
R3052 a_n6722_16092.n69 a_n6722_16092.n66 0.036
R3053 a_n6722_16092.n5 a_n6722_16092.n6 0.035
R3054 a_n6722_16092.n84 a_n6722_16092.n4 0.029
R3055 a_n6722_16092.n44 a_n6722_16092.n42 0.026
R3056 a_n6722_16092.n59 a_n6722_16092.n50 0.026
R3057 a_n6722_16092.n32 a_n6722_16092.n7 0.023
R3058 a_n6722_16092.n77 a_n6722_16092.n5 0.023
R3059 a_n6722_16092.n82 a_n6722_16092.n78 0.021
R3060 a_n6722_16092.n90 a_n6722_16092.n89 0.021
R3061 a_n6722_16092.n92 a_n6722_16092.n90 0.019
R3062 a_n6722_16092.n50 a_n6722_16092.n49 0.015
R3063 a_n6722_16092.n66 a_n6722_16092.n65 0.014
R3064 a_n6722_16092.n42 a_n6722_16092.n40 0.014
R3065 a_n6722_16092.n47 a_n6722_16092.n44 0.014
R3066 a_n6722_16092.n94 a_n6722_16092.n92 0.014
R3067 a_n6722_16092.n26 a_n6722_16092.n24 0.014
R3068 a_n6722_16092.n62 a_n6722_16092.n61 0.014
R3069 a_n5934_16092.n5 a_n5934_16092.n93 9.3
R3070 a_n5934_16092.n7 a_n5934_16092.n85 9.3
R3071 a_n5934_16092.n8 a_n5934_16092.n83 9.3
R3072 a_n5934_16092.n2 a_n5934_16092.n79 9.3
R3073 a_n5934_16092.n73 a_n5934_16092.n72 9.3
R3074 a_n5934_16092.n2 a_n5934_16092.n78 9.3
R3075 a_n5934_16092.n3 a_n5934_16092.n77 9.3
R3076 a_n5934_16092.n71 a_n5934_16092.n70 9.3
R3077 a_n5934_16092.n0 a_n5934_16092.n67 9.3
R3078 a_n5934_16092.n63 a_n5934_16092.n62 9.3
R3079 a_n5934_16092.n57 a_n5934_16092.n61 9.3
R3080 a_n5934_16092.n7 a_n5934_16092.n86 9.3
R3081 a_n5934_16092.n49 a_n5934_16092.n48 9.3
R3082 a_n5934_16092.n4 a_n5934_16092.n94 9.3
R3083 a_n5934_16092.n1 a_n5934_16092.n35 9.3
R3084 a_n5934_16092.n31 a_n5934_16092.n30 9.3
R3085 a_n5934_16092.n6 a_n5934_16092.n37 9.3
R3086 a_n5934_16092.n103 a_n5934_16092.n102 9.3
R3087 a_n5934_16092.n26 a_n5934_16092.n25 9.3
R3088 a_n5934_16092.n29 a_n5934_16092.n28 9.3
R3089 a_n5934_16092.n1 a_n5934_16092.n34 9.3
R3090 a_n5934_16092.n6 a_n5934_16092.n38 9.3
R3091 a_n5934_16092.n47 a_n5934_16092.n46 9
R3092 a_n5934_16092.n3 a_n5934_16092.n55 9
R3093 a_n5934_16092.n69 a_n5934_16092.n68 9
R3094 a_n5934_16092.n58 a_n5934_16092.n56 9
R3095 a_n5934_16092.n8 a_n5934_16092.n84 9
R3096 a_n5934_16092.n88 a_n5934_16092.n87 9
R3097 a_n5934_16092.n4 a_n5934_16092.n95 9
R3098 a_n5934_16092.n105 a_n5934_16092.n104 9
R3099 a_n5934_16092.n40 a_n5934_16092.n39 9
R3100 a_n5934_16092.n110 a_n5934_16092.n17 8.473
R3101 a_n5934_16092.n110 a_n5934_16092.n20 8.097
R3102 a_n5934_16092.n110 a_n5934_16092.n15 8.069
R3103 a_n5934_16092.n110 a_n5934_16092.n23 8.043
R3104 a_n5934_16092.n110 a_n5934_16092.n12 8.016
R3105 a_n5934_16092.n54 a_n5934_16092.n53 4.574
R3106 a_n5934_16092.n100 a_n5934_16092.n99 4.574
R3107 a_n5934_16092.n53 a_n5934_16092.n51 3.388
R3108 a_n5934_16092.n99 a_n5934_16092.n97 3.388
R3109 a_n5934_16092.n41 a_n5934_16092.t2 3.326
R3110 a_n5934_16092.t1 a_n5934_16092.n110 3.326
R3111 a_n5934_16092.n9 a_n5934_16092.n5 2.561
R3112 a_n5934_16092.n96 a_n5934_16092.n90 2.473
R3113 a_n5934_16092.n14 a_n5934_16092.n13 2.258
R3114 a_n5934_16092.n19 a_n5934_16092.n18 2.258
R3115 a_n5934_16092.n90 a_n5934_16092.n89 1.94
R3116 a_n5934_16092.n22 a_n5934_16092.n21 1.505
R3117 a_n5934_16092.n17 a_n5934_16092.n16 1.505
R3118 a_n5934_16092.n42 a_n5934_16092.n41 1.155
R3119 a_n5934_16092.n110 a_n5934_16092.n109 1.155
R3120 a_n5934_16092.n43 a_n5934_16092.n42 0.852
R3121 a_n5934_16092.n109 a_n5934_16092.n108 0.852
R3122 a_n5934_16092.n11 a_n5934_16092.n10 0.752
R3123 a_n5934_16092.n99 a_n5934_16092.n98 0.506
R3124 a_n5934_16092.n53 a_n5934_16092.n52 0.506
R3125 a_n5934_16092.n83 a_n5934_16092.n82 0.476
R3126 a_n5934_16092.n12 a_n5934_16092.n11 0.476
R3127 a_n5934_16092.n23 a_n5934_16092.n22 0.445
R3128 a_n5934_16092.n77 a_n5934_16092.n76 0.445
R3129 a_n5934_16092.n67 a_n5934_16092.n66 0.414
R3130 a_n5934_16092.n15 a_n5934_16092.n14 0.414
R3131 a_n5934_16092.n20 a_n5934_16092.n19 0.382
R3132 a_n5934_16092.n61 a_n5934_16092.n60 0.382
R3133 a_n5934_16092.n9 a_n5934_16092.t0 0.179
R3134 a_n5934_16092.n32 a_n5934_16092.n31 0.06
R3135 a_n5934_16092.n80 a_n5934_16092.n2 0.06
R3136 a_n5934_16092.n74 a_n5934_16092.n73 0.06
R3137 a_n5934_16092.n65 a_n5934_16092.n64 0.06
R3138 a_n5934_16092.n90 a_n5934_16092.n9 0.056
R3139 a_n5934_16092.n89 a_n5934_16092.n54 0.054
R3140 a_n5934_16092.n100 a_n5934_16092.n96 0.054
R3141 a_n5934_16092.n96 a_n5934_16092.n40 0.053
R3142 a_n5934_16092.n89 a_n5934_16092.n88 0.053
R3143 a_n5934_16092.n57 a_n5934_16092.n59 0.043
R3144 a_n5934_16092.n108 a_n5934_16092.n107 0.04
R3145 a_n5934_16092.n106 a_n5934_16092.n105 0.04
R3146 a_n5934_16092.n6 a_n5934_16092.n36 0.091
R3147 a_n5934_16092.n26 a_n5934_16092.n24 9.474
R3148 a_n5934_16092.n36 a_n5934_16092.n1 0.069
R3149 a_n5934_16092.n44 a_n5934_16092.n43 0.04
R3150 a_n5934_16092.n47 a_n5934_16092.n45 0.04
R3151 a_n5934_16092.n8 a_n5934_16092.n81 0.04
R3152 a_n5934_16092.n5 a_n5934_16092.n4 0.04
R3153 a_n5934_16092.n2 a_n5934_16092.n3 0.04
R3154 a_n5934_16092.n0 a_n5934_16092.n65 0.036
R3155 a_n5934_16092.n7 a_n5934_16092.n8 0.035
R3156 a_n5934_16092.n3 a_n5934_16092.n75 0.035
R3157 a_n5934_16092.n1 a_n5934_16092.n33 0.066
R3158 a_n5934_16092.n9 a_n5934_16092.n91 0.027
R3159 a_n5934_16092.n33 a_n5934_16092.n32 0.026
R3160 a_n5934_16092.n29 a_n5934_16092.n27 0.148
R3161 a_n5934_16092.n75 a_n5934_16092.n74 0.026
R3162 a_n5934_16092.n71 a_n5934_16092.n69 0.026
R3163 a_n5934_16092.n63 a_n5934_16092.n58 0.026
R3164 a_n5934_16092.n69 a_n5934_16092.n0 0.026
R3165 a_n5934_16092.n5 a_n5934_16092.n92 0.024
R3166 a_n5934_16092.n88 a_n5934_16092.n7 0.023
R3167 a_n5934_16092.n40 a_n5934_16092.n6 0.023
R3168 a_n5934_16092.n107 a_n5934_16092.n106 0.021
R3169 a_n5934_16092.n101 a_n5934_16092.n100 0.021
R3170 a_n5934_16092.n45 a_n5934_16092.n44 0.021
R3171 a_n5934_16092.n54 a_n5934_16092.n50 0.021
R3172 a_n5934_16092.n103 a_n5934_16092.n101 0.019
R3173 a_n5934_16092.n27 a_n5934_16092.n26 0.019
R3174 a_n5934_16092.n50 a_n5934_16092.n49 0.019
R3175 a_n5934_16092.n64 a_n5934_16092.n63 0.019
R3176 a_n5934_16092.n81 a_n5934_16092.n80 0.016
R3177 a_n5934_16092.n58 a_n5934_16092.n57 0.014
R3178 a_n5934_16092.n105 a_n5934_16092.n103 0.014
R3179 a_n5934_16092.n31 a_n5934_16092.n29 0.014
R3180 a_n5934_16092.n49 a_n5934_16092.n47 0.014
R3181 a_n5934_16092.n73 a_n5934_16092.n71 0.014
C11 BIAS_BOT VLO 28.25fF $ **FLOATING
C12 SS VLO 11.81fF
C13 D1 VLO 37.75fF
C14 VIN VLO 23.70fF $ **FLOATING
C15 RFB_MID VLO 5.66fF $ **FLOATING
C16 S1 VLO 52.77fF
C17 G_TOP VLO 6.51fF $ **FLOATING
C18 BIAS_TOP VLO 14.02fF $ **FLOATING
C19 VHI VLO 432.32fF $ **FLOATING
C20 VOUT VLO 75.58fF $ **FLOATING
C21 G4 VLO 1.28fF $ **FLOATING
C22 G8 VLO 1.10fF $ **FLOATING
C23 G1 VLO 1.06fF $ **FLOATING
C24 G2 VLO 1.29fF $ **FLOATING
C25 a_n5934_16092.n9 VLO 1.46fF
C26 a_n5934_16092.t0 VLO 9.51fF $ **FLOATING
C27 a_n6722_16092.t0 VLO 3.28fF $ **FLOATING
C28 a_n5540_16092.n4 VLO 1.02fF
C29 a_n5540_16092.t0 VLO 6.31fF $ **FLOATING
C30 a_n6328_16092.t0 VLO 2.94fF $ **FLOATING
C31 SS.n644 VLO 2.06fF
C32 SS.n1134 VLO 1.69fF
C33 SS.n1135 VLO 7.88fF
C34 SS.n1297 VLO 1.19fF
C35 SS.n1298 VLO 38.42fF
C36 D1.n0 VLO 3.62fF
C37 D1.n12 VLO 19.83fF
C38 S1.n21 VLO 5.21fF
C39 S1.n22 VLO 5.35fF
C40 S1.n23 VLO 14.34fF
C41 VOUT.n190 VLO 20.71fF
C42 VOUT.n236 VLO 1.35fF
C43 VOUT.n707 VLO 2.07fF
C44 VOUT.n1309 VLO 67.82fF


**** end user architecture code
.ends

.GLOBAL GND
.GLOBAL GNDI
.end
