magic
tech sky130A
timestamp 1665276793
<< metal3 >>
rect -30800 4300 -25200 4400
rect -30800 -1400 -30700 4300
rect -30000 -1400 -25200 4300
rect -30800 -1500 -25200 -1400
rect -24800 4300 -19200 4400
rect -24800 -1400 -20000 4300
rect -19300 -1400 -19200 4300
rect -24800 -1500 -19200 -1400
rect -40500 -3600 -27500 -3500
rect -40500 -7900 -28800 -3600
rect -27600 -7900 -27500 -3600
rect -40500 -8000 -27500 -7900
rect -22500 -3600 -9500 -3500
rect -22500 -7900 -22400 -3600
rect -21200 -7900 -9500 -3600
rect -22500 -8000 -9500 -7900
rect -36500 -27900 -31195 -27885
rect -36500 -28175 -31375 -27900
rect -31210 -28175 -31195 -27900
rect -36500 -28190 -31195 -28175
rect -36500 -28245 -31380 -28190
rect -18805 -28210 -18610 -28195
rect -36500 -48600 -36000 -28245
rect -18805 -28590 -18790 -28210
rect -18625 -28245 -18610 -28210
rect -18625 -28590 -13500 -28245
rect -18805 -28605 -13500 -28590
rect -35500 -46600 -14500 -32500
rect -35500 -48400 -35400 -46600
rect -14600 -48400 -14500 -46600
rect -35500 -48500 -14500 -48400
rect -14000 -48500 -13500 -28605
<< via3 >>
rect -30700 -1400 -30000 4300
rect -20000 -1400 -19300 4300
rect -28800 -7900 -27600 -3600
rect -22400 -7900 -21200 -3600
rect -31375 -28175 -31210 -27900
rect -18790 -28590 -18625 -28210
rect -35400 -48400 -14600 -46600
<< mimcap >>
rect -29500 4200 -25300 4300
rect -29500 -1300 -29400 4200
rect -25400 -1300 -25300 4200
rect -29500 -1400 -25300 -1300
rect -24700 4200 -20500 4300
rect -24700 -1300 -24600 4200
rect -20600 -1300 -20500 4200
rect -24700 -1400 -20500 -1300
rect -40400 -3700 -29300 -3600
rect -40400 -7800 -40300 -3700
rect -29400 -7800 -29300 -3700
rect -40400 -7900 -29300 -7800
rect -20700 -3700 -9600 -3600
rect -20700 -7800 -20600 -3700
rect -9700 -7800 -9600 -3700
rect -20700 -7900 -9600 -7800
rect -35400 -32700 -14600 -32600
rect -35400 -45300 -35300 -32700
rect -14700 -45300 -14600 -32700
rect -35400 -45400 -14600 -45300
<< mimcapcontact >>
rect -29400 -1300 -25400 4200
rect -24600 -1300 -20600 4200
rect -40300 -7800 -29400 -3700
rect -20600 -7800 -9700 -3700
rect -35300 -45300 -14700 -32700
<< metal4 >>
rect -30800 4300 -29900 4400
rect -30800 -1400 -30700 4300
rect -30000 -1400 -29900 4300
rect -30800 -1500 -29900 -1400
rect -29600 4200 -20400 4400
rect -29600 -1300 -29400 4200
rect -25400 -1300 -24600 4200
rect -20600 -1300 -20400 4200
rect -29600 -1500 -20400 -1300
rect -20100 4300 -19200 4400
rect -20100 -1400 -20000 4300
rect -19300 -1400 -19200 4300
rect -20100 -1500 -19200 -1400
rect -40500 -3700 -29200 -3500
rect -40500 -7800 -40300 -3700
rect -29400 -7800 -29200 -3700
rect -40500 -8000 -29200 -7800
rect -28900 -3600 -27500 -3500
rect -28900 -7900 -28800 -3600
rect -27600 -7900 -27500 -3600
rect -28900 -8000 -27500 -7900
rect -22500 -3600 -21100 -3500
rect -22500 -7900 -22400 -3600
rect -21200 -7900 -21100 -3600
rect -22500 -8000 -21100 -7900
rect -20800 -3700 -9500 -3500
rect -20800 -7800 -20600 -3700
rect -9700 -7800 -9500 -3700
rect -20800 -8000 -9500 -7800
rect -40500 -10300 -34900 -8000
rect -15100 -10300 -9500 -8000
rect -31390 -27900 -31195 -27885
rect -31390 -28175 -31375 -27900
rect -31210 -28175 -31195 -27900
rect -31390 -28190 -31195 -28175
rect -18805 -28210 -18610 -28195
rect -18805 -28590 -18790 -28210
rect -18625 -28590 -18610 -28210
rect -18805 -28605 -18610 -28590
rect -48500 -32700 -1500 -32500
rect -48500 -33000 -35300 -32700
rect -48500 -45000 -48000 -33000
rect -37500 -45000 -35300 -33000
rect -48500 -45300 -35300 -45000
rect -14700 -33000 -1500 -32700
rect -14700 -45000 -12500 -33000
rect -2000 -45000 -1500 -33000
rect -14700 -45300 -1500 -45000
rect -48500 -45500 -1500 -45300
rect -35500 -46600 -14500 -46500
rect -35500 -48400 -35400 -46600
rect -14600 -48400 -14500 -46600
rect -35500 -48500 -14500 -48400
<< via4 >>
rect -30700 -1400 -30000 4300
rect -20000 -1400 -19300 4300
rect -28800 -7900 -27600 -3600
rect -22400 -7900 -21200 -3600
rect -31375 -28175 -31210 -27900
rect -18790 -28590 -18625 -28210
rect -48000 -45000 -37500 -33000
rect -12500 -45000 -2000 -33000
rect -35400 -48400 -14600 -46600
<< mimcap2 >>
rect -29500 4200 -25300 4300
rect -29500 -1300 -29400 4200
rect -25400 -1300 -25300 4200
rect -29500 -1400 -25300 -1300
rect -24700 4200 -20500 4300
rect -24700 -1300 -24600 4200
rect -20600 -1300 -20500 4200
rect -24700 -1400 -20500 -1300
rect -35400 -32700 -14600 -32600
rect -35400 -45300 -35300 -32700
rect -14700 -45300 -14600 -32700
rect -35400 -45400 -14600 -45300
<< mimcap2contact >>
rect -29400 -1300 -25400 4200
rect -24600 -1300 -20600 4200
rect -35300 -45300 -14700 -32700
<< metal5 >>
rect -29500 10200 -27500 11600
rect -30700 8900 -27500 10200
rect -22500 10200 -20500 11600
rect -22500 8900 -19300 10200
rect -30700 8200 -29500 8900
rect -32300 6400 -29500 8200
rect -35900 5900 -29500 6400
rect -36500 4400 -29500 5900
rect -20500 8200 -19300 8900
rect -20500 6400 -17700 8200
rect -20500 5900 -14100 6400
rect -20500 4400 -13500 5900
rect -36500 4300 -25200 4400
rect -36500 -1400 -30700 4300
rect -30000 4200 -25200 4300
rect -30000 -1300 -29400 4200
rect -25400 -1300 -25200 4200
rect -30000 -1400 -25200 -1300
rect -36500 -1500 -25200 -1400
rect -24800 4300 -13500 4400
rect -24800 4200 -20000 4300
rect -24800 -1300 -24600 4200
rect -20600 -1300 -20000 4200
rect -24800 -1400 -20000 -1300
rect -19300 -1400 -13500 4300
rect -24800 -1500 -13500 -1400
rect -36500 -3500 -29500 -1500
rect -20500 -3500 -13500 -1500
rect -40500 -3600 -27500 -3500
rect -40500 -7900 -28800 -3600
rect -27600 -7900 -27500 -3600
rect -40500 -8000 -27500 -7900
rect -22500 -3600 -9500 -3500
rect -22500 -7900 -22400 -3600
rect -21200 -7900 -9500 -3600
rect -22500 -8000 -9500 -7900
rect -31100 -8400 -28900 -8000
rect -21100 -8400 -18900 -8000
rect -31100 -8500 -30300 -8400
rect -19700 -8500 -18900 -8400
rect -40900 -26000 -37300 -23300
rect -43600 -28700 -37300 -26000
rect -12700 -26000 -9100 -23300
rect -31390 -27900 -31195 -27885
rect -31390 -28175 -31375 -27900
rect -31210 -28175 -31195 -27900
rect -31390 -28190 -31195 -28175
rect -18805 -28210 -18610 -28195
rect -18805 -28590 -18790 -28210
rect -18625 -28590 -18610 -28210
rect -18805 -28605 -18610 -28590
rect -45700 -31500 -37300 -28700
rect -48500 -32500 -37300 -31500
rect -12700 -28700 -6400 -26000
rect -12700 -31500 -4300 -28700
rect -35400 -32500 -14600 -32100
rect -12700 -32500 -1500 -31500
rect -48500 -33000 -37000 -32500
rect -48500 -33500 -48000 -33000
rect -50800 -36300 -48000 -33500
rect -52900 -38400 -48000 -36300
rect -57500 -40000 -48000 -38400
rect -48500 -45000 -48000 -40000
rect -37500 -45000 -37000 -33000
rect -48500 -45500 -37000 -45000
rect -35500 -32700 -14500 -32500
rect -35500 -45300 -35300 -32700
rect -14700 -45300 -14500 -32700
rect -35500 -46600 -14500 -45300
rect -13000 -33000 -1500 -32500
rect -13000 -45000 -12500 -33000
rect -2000 -33500 -1500 -33000
rect -2000 -36300 800 -33500
rect -2000 -38400 2900 -36300
rect -2000 -40000 7500 -38400
rect -2000 -45000 -1500 -40000
rect -13000 -45500 -1500 -45000
rect -35500 -48400 -35400 -46600
rect -14600 -48400 -14500 -46600
rect -35500 -48500 -14500 -48400
<< comment >>
rect -31390 -27875 -31385 -27870
use cascode_complete_3  cascode_complete_3_0
timestamp 1665275542
transform 1 0 -31700 0 1 -32700
box -3600 0 17000 24250
use octa_ind_1p5n_highQ  octa_ind_1p5n_highQ_0
timestamp 1665275929
transform 0 -1 -21000 1 0 33600
box -30500 -21500 10500 1500
use octa_ind_1p5n_highQ  octa_ind_1p5n_highQ_1
timestamp 1665275929
transform 0 1 -29000 1 0 33600
box -30500 -21500 10500 1500
use octa_ind_3p5n_highQ  octa_ind_3p5n_highQ_0
timestamp 1665269856
transform 1 0 29300 0 -1 -23800
box -42000 -36250 18000 16250
use octa_ind_3p5n_highQ  octa_ind_3p5n_highQ_1
timestamp 1665269856
transform -1 0 -79300 0 -1 -23800
box -42000 -36250 18000 16250
<< end >>
