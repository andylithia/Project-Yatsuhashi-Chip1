magic
tech sky130B
magscale 1 2
timestamp 1662258694
<< error_p >>
rect -293 757 -247 769
rect -185 757 -139 769
rect -77 757 -31 769
rect 31 757 77 769
rect 139 757 185 769
rect 247 757 293 769
rect -293 717 -287 757
rect -185 717 -179 757
rect -77 717 -71 757
rect 31 717 37 757
rect 139 717 145 757
rect 247 717 253 757
rect -293 705 -247 717
rect -185 705 -139 717
rect -77 705 -31 717
rect 31 705 77 717
rect 139 705 185 717
rect 247 705 293 717
rect -293 -717 -247 -705
rect -185 -717 -139 -705
rect -77 -717 -31 -705
rect 31 -717 77 -705
rect 139 -717 185 -705
rect 247 -717 293 -705
rect -293 -757 -287 -717
rect -185 -757 -179 -717
rect -77 -757 -71 -717
rect 31 -757 37 -717
rect 139 -757 145 -717
rect 247 -757 253 -717
rect -293 -769 -247 -757
rect -185 -769 -139 -757
rect -77 -769 -31 -757
rect 31 -769 77 -757
rect 139 -769 185 -757
rect 247 -769 293 -757
<< pwell >>
rect -469 -939 469 939
<< psubdiff >>
rect -433 869 -337 903
rect 337 869 433 903
rect -433 807 -399 869
rect 399 807 433 869
rect -433 -869 -399 -807
rect 399 -869 433 -807
rect -433 -903 -337 -869
rect 337 -903 433 -869
<< psubdiffcont >>
rect -337 869 337 903
rect -433 -807 -399 807
rect 399 -807 433 807
rect -337 -903 337 -869
<< poly >>
rect -303 757 -237 773
rect -303 723 -287 757
rect -253 723 -237 757
rect -303 700 -237 723
rect -303 -723 -237 -700
rect -303 -757 -287 -723
rect -253 -757 -237 -723
rect -303 -773 -237 -757
rect -195 757 -129 773
rect -195 723 -179 757
rect -145 723 -129 757
rect -195 700 -129 723
rect -195 -723 -129 -700
rect -195 -757 -179 -723
rect -145 -757 -129 -723
rect -195 -773 -129 -757
rect -87 757 -21 773
rect -87 723 -71 757
rect -37 723 -21 757
rect -87 700 -21 723
rect -87 -723 -21 -700
rect -87 -757 -71 -723
rect -37 -757 -21 -723
rect -87 -773 -21 -757
rect 21 757 87 773
rect 21 723 37 757
rect 71 723 87 757
rect 21 700 87 723
rect 21 -723 87 -700
rect 21 -757 37 -723
rect 71 -757 87 -723
rect 21 -773 87 -757
rect 129 757 195 773
rect 129 723 145 757
rect 179 723 195 757
rect 129 700 195 723
rect 129 -723 195 -700
rect 129 -757 145 -723
rect 179 -757 195 -723
rect 129 -773 195 -757
rect 237 757 303 773
rect 237 723 253 757
rect 287 723 303 757
rect 237 700 303 723
rect 237 -723 303 -700
rect 237 -757 253 -723
rect 287 -757 303 -723
rect 237 -773 303 -757
<< polycont >>
rect -287 723 -253 757
rect -287 -757 -253 -723
rect -179 723 -145 757
rect -179 -757 -145 -723
rect -71 723 -37 757
rect -71 -757 -37 -723
rect 37 723 71 757
rect 37 -757 71 -723
rect 145 723 179 757
rect 145 -757 179 -723
rect 253 723 287 757
rect 253 -757 287 -723
<< npolyres >>
rect -303 -700 -237 700
rect -195 -700 -129 700
rect -87 -700 -21 700
rect 21 -700 87 700
rect 129 -700 195 700
rect 237 -700 303 700
<< locali >>
rect -433 869 -337 903
rect 337 869 433 903
rect -433 807 -399 869
rect 399 807 433 869
rect -303 723 -287 757
rect -253 723 -237 757
rect -195 723 -179 757
rect -145 723 -129 757
rect -87 723 -71 757
rect -37 723 -21 757
rect 21 723 37 757
rect 71 723 87 757
rect 129 723 145 757
rect 179 723 195 757
rect 237 723 253 757
rect 287 723 303 757
rect -303 -757 -287 -723
rect -253 -757 -237 -723
rect -195 -757 -179 -723
rect -145 -757 -129 -723
rect -87 -757 -71 -723
rect -37 -757 -21 -723
rect 21 -757 37 -723
rect 71 -757 87 -723
rect 129 -757 145 -723
rect 179 -757 195 -723
rect 237 -757 253 -723
rect 287 -757 303 -723
rect -433 -869 -399 -807
rect 399 -869 433 -807
rect -433 -903 -337 -869
rect 337 -903 433 -869
<< viali >>
rect -287 723 -253 757
rect -179 723 -145 757
rect -71 723 -37 757
rect 37 723 71 757
rect 145 723 179 757
rect 253 723 287 757
rect -287 717 -253 723
rect -179 717 -145 723
rect -71 717 -37 723
rect 37 717 71 723
rect 145 717 179 723
rect 253 717 287 723
rect -287 -723 -253 -717
rect -179 -723 -145 -717
rect -71 -723 -37 -717
rect 37 -723 71 -717
rect 145 -723 179 -717
rect 253 -723 287 -717
rect -287 -757 -253 -723
rect -179 -757 -145 -723
rect -71 -757 -37 -723
rect 37 -757 71 -723
rect 145 -757 179 -723
rect 253 -757 287 -723
<< metal1 >>
rect -293 757 -247 769
rect -293 717 -287 757
rect -253 717 -247 757
rect -293 705 -247 717
rect -185 757 -139 769
rect -185 717 -179 757
rect -145 717 -139 757
rect -185 705 -139 717
rect -77 757 -31 769
rect -77 717 -71 757
rect -37 717 -31 757
rect -77 705 -31 717
rect 31 757 77 769
rect 31 717 37 757
rect 71 717 77 757
rect 31 705 77 717
rect 139 757 185 769
rect 139 717 145 757
rect 179 717 185 757
rect 139 705 185 717
rect 247 757 293 769
rect 247 717 253 757
rect 287 717 293 757
rect 247 705 293 717
rect -293 -717 -247 -705
rect -293 -757 -287 -717
rect -253 -757 -247 -717
rect -293 -769 -247 -757
rect -185 -717 -139 -705
rect -185 -757 -179 -717
rect -145 -757 -139 -717
rect -185 -769 -139 -757
rect -77 -717 -31 -705
rect -77 -757 -71 -717
rect -37 -757 -31 -717
rect -77 -769 -31 -757
rect 31 -717 77 -705
rect 31 -757 37 -717
rect 71 -757 77 -717
rect 31 -769 77 -757
rect 139 -717 185 -705
rect 139 -757 145 -717
rect 179 -757 185 -717
rect 139 -769 185 -757
rect 247 -717 293 -705
rect 247 -757 253 -717
rect 287 -757 293 -717
rect 247 -769 293 -757
<< properties >>
string FIXED_BBOX -416 -886 416 886
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 7 m 1 nx 6 wmin 0.330 lmin 1.650 rho 48.2 val 1.022k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
