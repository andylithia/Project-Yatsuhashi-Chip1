* NGSPICE file created from pex_test.ext - technology: sky130B

C0 B VSUBS 109.26fF $ **FLOATING
