magic
tech sky130A
timestamp 1664804552
<< metal4 >>
rect -300 23750 400 23800
rect -300 23250 -250 23750
rect 350 23250 400 23750
rect -300 23200 400 23250
rect -500 23000 400 23200
rect -1700 20400 400 23000
rect -500 19550 400 20400
rect -1700 19300 -800 19350
rect -1700 18800 -1450 19300
rect -850 18800 -800 19300
rect -1700 12450 -800 18800
rect -3050 7150 -800 12450
rect -1700 6900 -800 7150
rect -1700 6400 -1650 6900
rect -850 6400 -800 6900
rect -1700 6350 -800 6400
rect -500 12750 -300 19550
rect 350 12750 400 19550
rect -500 11600 400 12750
rect -500 7350 -300 11600
rect 350 7350 400 11600
rect -500 1800 400 7350
rect 13000 23750 13700 23800
rect 13000 23250 13050 23750
rect 13650 23250 13700 23750
rect 13000 23200 13700 23250
rect 13000 23000 13900 23200
rect 13000 20400 15100 23000
rect 13000 19100 13900 20400
rect 13000 12300 13050 19100
rect 13700 12300 13900 19100
rect 13000 11150 13900 12300
rect 13000 7350 13050 11150
rect 13700 7800 13900 11150
rect 13850 7350 13900 7800
rect 13000 1800 13900 7350
rect 14100 19300 15000 19350
rect 14100 18800 14150 19300
rect 14750 18800 15000 19300
rect 14100 12450 15000 18800
rect 14100 7150 16350 12450
rect 14100 6900 15000 7150
rect 14100 6400 14150 6900
rect 14950 6400 15000 6900
rect 14100 6350 15000 6400
<< via4 >>
rect -250 23250 350 23750
rect -1450 18800 -850 19300
rect -1650 6400 -850 6900
rect -300 12750 350 19550
rect -300 7350 350 11600
rect 13050 23250 13650 23750
rect 13050 12300 13700 19100
rect 13050 7800 13700 11150
rect 13050 7350 13850 7800
rect 14150 18800 14750 19300
rect 14150 6400 14950 6900
<< mimcap2 >>
rect -1650 22900 350 22950
rect -1650 20500 -1600 22900
rect 300 20500 350 22900
rect -1650 20450 350 20500
rect 13050 22900 15050 22950
rect 13050 20500 13100 22900
rect 15000 20500 15050 22900
rect 13050 20450 15050 20500
rect -1650 18450 -850 18500
rect -1650 13350 -1600 18450
rect -900 13350 -850 18450
rect -1650 13300 -850 13350
rect 14150 18450 14950 18500
rect 14150 13350 14200 18450
rect 14900 13350 14950 18450
rect 14150 13300 14950 13350
rect -3000 7200 -850 12400
rect 14150 7200 16300 12400
rect -450 7000 350 7050
rect -450 1900 -400 7000
rect 300 1900 350 7000
rect -450 1850 350 1900
rect 13050 7000 13850 7050
rect 13050 1900 13100 7000
rect 13800 1900 13850 7000
rect 13050 1850 13850 1900
<< mimcap2contact >>
rect -1600 20500 300 22900
rect 13100 20500 15000 22900
rect -1600 13350 -900 18450
rect 14200 13350 14900 18450
rect -400 1900 300 7000
rect 13100 1900 13800 7000
<< metal5 >>
rect -300 23750 650 23800
rect -300 23250 -250 23750
rect 350 23350 650 23750
rect 12750 23750 13700 23800
rect 12750 23350 13050 23750
rect 350 23250 400 23350
rect -300 23200 400 23250
rect 13000 23250 13050 23350
rect 13650 23250 13700 23750
rect 13000 23200 13700 23250
rect -1700 22900 400 23000
rect -1700 20500 -1600 22900
rect 300 20500 400 22900
rect -1700 20400 400 20500
rect 13000 22900 15100 23000
rect 13000 20500 13100 22900
rect 15000 20500 15100 22900
rect 13000 20400 15100 20500
rect -1500 19850 600 20100
rect -1500 19300 -800 19850
rect -1500 18800 -1450 19300
rect -850 18800 -800 19300
rect -1500 18750 -800 18800
rect -350 19550 400 19600
rect -1700 18450 -800 18550
rect -1700 13350 -1600 18450
rect -900 13350 -800 18450
rect -1700 13250 -800 13350
rect -350 12750 -300 19550
rect 350 12750 400 19550
rect 12700 19400 14800 19650
rect 14100 19300 14800 19400
rect -350 12700 400 12750
rect 13000 19100 13750 19150
rect -3050 12200 600 12450
rect 13000 12300 13050 19100
rect 13700 12300 13750 19100
rect 14100 18800 14150 19300
rect 14750 18800 14800 19300
rect 14100 18750 14800 18800
rect 14100 18450 15000 18550
rect 14100 13350 14200 18450
rect 14900 13350 15000 18450
rect 14100 13250 15000 13350
rect 13000 12250 13750 12300
rect -3050 11900 150 12200
rect 14100 12000 16350 12450
rect -3050 7150 -800 11900
rect 12700 11750 16350 12000
rect -350 11600 400 11650
rect -350 7350 -300 11600
rect 350 8950 400 11600
rect 13150 11450 16350 11750
rect 13000 11150 13750 11200
rect 350 8250 650 8950
rect 350 7350 400 8250
rect 13000 7850 13050 11150
rect -350 7300 400 7350
rect 12750 7350 13050 7850
rect 13700 7850 13750 11150
rect 13700 7800 13900 7850
rect 13850 7350 13900 7800
rect 12750 7300 13900 7350
rect 14100 7150 16350 11450
rect -500 7000 400 7100
rect -1700 6900 -800 6950
rect -1700 6400 -1650 6900
rect -850 6400 -800 6900
rect -1700 1800 -800 6400
rect -500 1900 -400 7000
rect 300 1900 400 7000
rect -500 1800 400 1900
rect 13000 7000 13900 7100
rect 13000 1900 13100 7000
rect 13800 1900 13900 7000
rect 13000 1800 13900 1900
rect 14100 6900 15000 6950
rect 14100 6400 14150 6900
rect 14950 6400 15000 6900
rect 14100 1800 15000 6400
rect -1700 1100 700 1800
rect 12000 1100 15000 1800
rect 12000 850 12750 1100
use cascode_1  cascode_1_0
timestamp 1664506494
transform 1 0 7350 0 1 -1850
box -7350 1850 5400 26100
<< end >>
