magic
tech sky130B
magscale 1 2
timestamp 1661915753
<< pwell >>
rect 0 66 1686 1128
<< nmos >>
rect 194 92 224 1102
rect 280 92 310 1102
rect 588 92 618 1102
rect 674 92 704 1102
rect 982 92 1012 1102
rect 1068 92 1098 1102
rect 1376 92 1406 1102
rect 1462 92 1492 1102
<< ndiff >>
rect 138 1090 194 1102
rect 138 1056 149 1090
rect 183 1056 194 1090
rect 138 1022 194 1056
rect 138 988 149 1022
rect 183 988 194 1022
rect 138 954 194 988
rect 138 920 149 954
rect 183 920 194 954
rect 138 886 194 920
rect 138 852 149 886
rect 183 852 194 886
rect 138 818 194 852
rect 138 784 149 818
rect 183 784 194 818
rect 138 750 194 784
rect 138 716 149 750
rect 183 716 194 750
rect 138 682 194 716
rect 138 648 149 682
rect 183 648 194 682
rect 138 614 194 648
rect 138 580 149 614
rect 183 580 194 614
rect 138 546 194 580
rect 138 512 149 546
rect 183 512 194 546
rect 138 478 194 512
rect 138 444 149 478
rect 183 444 194 478
rect 138 410 194 444
rect 138 376 149 410
rect 183 376 194 410
rect 138 342 194 376
rect 138 308 149 342
rect 183 308 194 342
rect 138 274 194 308
rect 138 240 149 274
rect 183 240 194 274
rect 138 206 194 240
rect 138 172 149 206
rect 183 172 194 206
rect 138 138 194 172
rect 138 104 149 138
rect 183 104 194 138
rect 138 92 194 104
rect 224 1090 280 1102
rect 224 1056 235 1090
rect 269 1056 280 1090
rect 224 1022 280 1056
rect 224 988 235 1022
rect 269 988 280 1022
rect 224 954 280 988
rect 224 920 235 954
rect 269 920 280 954
rect 224 886 280 920
rect 224 852 235 886
rect 269 852 280 886
rect 224 818 280 852
rect 224 784 235 818
rect 269 784 280 818
rect 224 750 280 784
rect 224 716 235 750
rect 269 716 280 750
rect 224 682 280 716
rect 224 648 235 682
rect 269 648 280 682
rect 224 614 280 648
rect 224 580 235 614
rect 269 580 280 614
rect 224 546 280 580
rect 224 512 235 546
rect 269 512 280 546
rect 224 478 280 512
rect 224 444 235 478
rect 269 444 280 478
rect 224 410 280 444
rect 224 376 235 410
rect 269 376 280 410
rect 224 342 280 376
rect 224 308 235 342
rect 269 308 280 342
rect 224 274 280 308
rect 224 240 235 274
rect 269 240 280 274
rect 224 206 280 240
rect 224 172 235 206
rect 269 172 280 206
rect 224 138 280 172
rect 224 104 235 138
rect 269 104 280 138
rect 224 92 280 104
rect 310 1090 366 1102
rect 310 1056 321 1090
rect 355 1056 366 1090
rect 310 1022 366 1056
rect 310 988 321 1022
rect 355 988 366 1022
rect 310 954 366 988
rect 310 920 321 954
rect 355 920 366 954
rect 310 886 366 920
rect 310 852 321 886
rect 355 852 366 886
rect 310 818 366 852
rect 310 784 321 818
rect 355 784 366 818
rect 310 750 366 784
rect 310 716 321 750
rect 355 716 366 750
rect 310 682 366 716
rect 310 648 321 682
rect 355 648 366 682
rect 310 614 366 648
rect 310 580 321 614
rect 355 580 366 614
rect 310 546 366 580
rect 310 512 321 546
rect 355 512 366 546
rect 310 478 366 512
rect 310 444 321 478
rect 355 444 366 478
rect 310 410 366 444
rect 310 376 321 410
rect 355 376 366 410
rect 310 342 366 376
rect 310 308 321 342
rect 355 308 366 342
rect 310 274 366 308
rect 310 240 321 274
rect 355 240 366 274
rect 310 206 366 240
rect 310 172 321 206
rect 355 172 366 206
rect 310 138 366 172
rect 310 104 321 138
rect 355 104 366 138
rect 310 92 366 104
rect 532 1090 588 1102
rect 532 1056 543 1090
rect 577 1056 588 1090
rect 532 1022 588 1056
rect 532 988 543 1022
rect 577 988 588 1022
rect 532 954 588 988
rect 532 920 543 954
rect 577 920 588 954
rect 532 886 588 920
rect 532 852 543 886
rect 577 852 588 886
rect 532 818 588 852
rect 532 784 543 818
rect 577 784 588 818
rect 532 750 588 784
rect 532 716 543 750
rect 577 716 588 750
rect 532 682 588 716
rect 532 648 543 682
rect 577 648 588 682
rect 532 614 588 648
rect 532 580 543 614
rect 577 580 588 614
rect 532 546 588 580
rect 532 512 543 546
rect 577 512 588 546
rect 532 478 588 512
rect 532 444 543 478
rect 577 444 588 478
rect 532 410 588 444
rect 532 376 543 410
rect 577 376 588 410
rect 532 342 588 376
rect 532 308 543 342
rect 577 308 588 342
rect 532 274 588 308
rect 532 240 543 274
rect 577 240 588 274
rect 532 206 588 240
rect 532 172 543 206
rect 577 172 588 206
rect 532 138 588 172
rect 532 104 543 138
rect 577 104 588 138
rect 532 92 588 104
rect 618 1090 674 1102
rect 618 1056 629 1090
rect 663 1056 674 1090
rect 618 1022 674 1056
rect 618 988 629 1022
rect 663 988 674 1022
rect 618 954 674 988
rect 618 920 629 954
rect 663 920 674 954
rect 618 886 674 920
rect 618 852 629 886
rect 663 852 674 886
rect 618 818 674 852
rect 618 784 629 818
rect 663 784 674 818
rect 618 750 674 784
rect 618 716 629 750
rect 663 716 674 750
rect 618 682 674 716
rect 618 648 629 682
rect 663 648 674 682
rect 618 614 674 648
rect 618 580 629 614
rect 663 580 674 614
rect 618 546 674 580
rect 618 512 629 546
rect 663 512 674 546
rect 618 478 674 512
rect 618 444 629 478
rect 663 444 674 478
rect 618 410 674 444
rect 618 376 629 410
rect 663 376 674 410
rect 618 342 674 376
rect 618 308 629 342
rect 663 308 674 342
rect 618 274 674 308
rect 618 240 629 274
rect 663 240 674 274
rect 618 206 674 240
rect 618 172 629 206
rect 663 172 674 206
rect 618 138 674 172
rect 618 104 629 138
rect 663 104 674 138
rect 618 92 674 104
rect 704 1090 760 1102
rect 704 1056 715 1090
rect 749 1056 760 1090
rect 704 1022 760 1056
rect 704 988 715 1022
rect 749 988 760 1022
rect 704 954 760 988
rect 704 920 715 954
rect 749 920 760 954
rect 704 886 760 920
rect 704 852 715 886
rect 749 852 760 886
rect 704 818 760 852
rect 704 784 715 818
rect 749 784 760 818
rect 704 750 760 784
rect 704 716 715 750
rect 749 716 760 750
rect 704 682 760 716
rect 704 648 715 682
rect 749 648 760 682
rect 704 614 760 648
rect 704 580 715 614
rect 749 580 760 614
rect 704 546 760 580
rect 704 512 715 546
rect 749 512 760 546
rect 704 478 760 512
rect 704 444 715 478
rect 749 444 760 478
rect 704 410 760 444
rect 704 376 715 410
rect 749 376 760 410
rect 704 342 760 376
rect 704 308 715 342
rect 749 308 760 342
rect 704 274 760 308
rect 704 240 715 274
rect 749 240 760 274
rect 704 206 760 240
rect 704 172 715 206
rect 749 172 760 206
rect 704 138 760 172
rect 704 104 715 138
rect 749 104 760 138
rect 704 92 760 104
rect 926 1090 982 1102
rect 926 1056 937 1090
rect 971 1056 982 1090
rect 926 1022 982 1056
rect 926 988 937 1022
rect 971 988 982 1022
rect 926 954 982 988
rect 926 920 937 954
rect 971 920 982 954
rect 926 886 982 920
rect 926 852 937 886
rect 971 852 982 886
rect 926 818 982 852
rect 926 784 937 818
rect 971 784 982 818
rect 926 750 982 784
rect 926 716 937 750
rect 971 716 982 750
rect 926 682 982 716
rect 926 648 937 682
rect 971 648 982 682
rect 926 614 982 648
rect 926 580 937 614
rect 971 580 982 614
rect 926 546 982 580
rect 926 512 937 546
rect 971 512 982 546
rect 926 478 982 512
rect 926 444 937 478
rect 971 444 982 478
rect 926 410 982 444
rect 926 376 937 410
rect 971 376 982 410
rect 926 342 982 376
rect 926 308 937 342
rect 971 308 982 342
rect 926 274 982 308
rect 926 240 937 274
rect 971 240 982 274
rect 926 206 982 240
rect 926 172 937 206
rect 971 172 982 206
rect 926 138 982 172
rect 926 104 937 138
rect 971 104 982 138
rect 926 92 982 104
rect 1012 1090 1068 1102
rect 1012 1056 1023 1090
rect 1057 1056 1068 1090
rect 1012 1022 1068 1056
rect 1012 988 1023 1022
rect 1057 988 1068 1022
rect 1012 954 1068 988
rect 1012 920 1023 954
rect 1057 920 1068 954
rect 1012 886 1068 920
rect 1012 852 1023 886
rect 1057 852 1068 886
rect 1012 818 1068 852
rect 1012 784 1023 818
rect 1057 784 1068 818
rect 1012 750 1068 784
rect 1012 716 1023 750
rect 1057 716 1068 750
rect 1012 682 1068 716
rect 1012 648 1023 682
rect 1057 648 1068 682
rect 1012 614 1068 648
rect 1012 580 1023 614
rect 1057 580 1068 614
rect 1012 546 1068 580
rect 1012 512 1023 546
rect 1057 512 1068 546
rect 1012 478 1068 512
rect 1012 444 1023 478
rect 1057 444 1068 478
rect 1012 410 1068 444
rect 1012 376 1023 410
rect 1057 376 1068 410
rect 1012 342 1068 376
rect 1012 308 1023 342
rect 1057 308 1068 342
rect 1012 274 1068 308
rect 1012 240 1023 274
rect 1057 240 1068 274
rect 1012 206 1068 240
rect 1012 172 1023 206
rect 1057 172 1068 206
rect 1012 138 1068 172
rect 1012 104 1023 138
rect 1057 104 1068 138
rect 1012 92 1068 104
rect 1098 1090 1154 1102
rect 1098 1056 1109 1090
rect 1143 1056 1154 1090
rect 1098 1022 1154 1056
rect 1098 988 1109 1022
rect 1143 988 1154 1022
rect 1098 954 1154 988
rect 1098 920 1109 954
rect 1143 920 1154 954
rect 1098 886 1154 920
rect 1098 852 1109 886
rect 1143 852 1154 886
rect 1098 818 1154 852
rect 1098 784 1109 818
rect 1143 784 1154 818
rect 1098 750 1154 784
rect 1098 716 1109 750
rect 1143 716 1154 750
rect 1098 682 1154 716
rect 1098 648 1109 682
rect 1143 648 1154 682
rect 1098 614 1154 648
rect 1098 580 1109 614
rect 1143 580 1154 614
rect 1098 546 1154 580
rect 1098 512 1109 546
rect 1143 512 1154 546
rect 1098 478 1154 512
rect 1098 444 1109 478
rect 1143 444 1154 478
rect 1098 410 1154 444
rect 1098 376 1109 410
rect 1143 376 1154 410
rect 1098 342 1154 376
rect 1098 308 1109 342
rect 1143 308 1154 342
rect 1098 274 1154 308
rect 1098 240 1109 274
rect 1143 240 1154 274
rect 1098 206 1154 240
rect 1098 172 1109 206
rect 1143 172 1154 206
rect 1098 138 1154 172
rect 1098 104 1109 138
rect 1143 104 1154 138
rect 1098 92 1154 104
rect 1320 1090 1376 1102
rect 1320 1056 1331 1090
rect 1365 1056 1376 1090
rect 1320 1022 1376 1056
rect 1320 988 1331 1022
rect 1365 988 1376 1022
rect 1320 954 1376 988
rect 1320 920 1331 954
rect 1365 920 1376 954
rect 1320 886 1376 920
rect 1320 852 1331 886
rect 1365 852 1376 886
rect 1320 818 1376 852
rect 1320 784 1331 818
rect 1365 784 1376 818
rect 1320 750 1376 784
rect 1320 716 1331 750
rect 1365 716 1376 750
rect 1320 682 1376 716
rect 1320 648 1331 682
rect 1365 648 1376 682
rect 1320 614 1376 648
rect 1320 580 1331 614
rect 1365 580 1376 614
rect 1320 546 1376 580
rect 1320 512 1331 546
rect 1365 512 1376 546
rect 1320 478 1376 512
rect 1320 444 1331 478
rect 1365 444 1376 478
rect 1320 410 1376 444
rect 1320 376 1331 410
rect 1365 376 1376 410
rect 1320 342 1376 376
rect 1320 308 1331 342
rect 1365 308 1376 342
rect 1320 274 1376 308
rect 1320 240 1331 274
rect 1365 240 1376 274
rect 1320 206 1376 240
rect 1320 172 1331 206
rect 1365 172 1376 206
rect 1320 138 1376 172
rect 1320 104 1331 138
rect 1365 104 1376 138
rect 1320 92 1376 104
rect 1406 1090 1462 1102
rect 1406 1056 1417 1090
rect 1451 1056 1462 1090
rect 1406 1022 1462 1056
rect 1406 988 1417 1022
rect 1451 988 1462 1022
rect 1406 954 1462 988
rect 1406 920 1417 954
rect 1451 920 1462 954
rect 1406 886 1462 920
rect 1406 852 1417 886
rect 1451 852 1462 886
rect 1406 818 1462 852
rect 1406 784 1417 818
rect 1451 784 1462 818
rect 1406 750 1462 784
rect 1406 716 1417 750
rect 1451 716 1462 750
rect 1406 682 1462 716
rect 1406 648 1417 682
rect 1451 648 1462 682
rect 1406 614 1462 648
rect 1406 580 1417 614
rect 1451 580 1462 614
rect 1406 546 1462 580
rect 1406 512 1417 546
rect 1451 512 1462 546
rect 1406 478 1462 512
rect 1406 444 1417 478
rect 1451 444 1462 478
rect 1406 410 1462 444
rect 1406 376 1417 410
rect 1451 376 1462 410
rect 1406 342 1462 376
rect 1406 308 1417 342
rect 1451 308 1462 342
rect 1406 274 1462 308
rect 1406 240 1417 274
rect 1451 240 1462 274
rect 1406 206 1462 240
rect 1406 172 1417 206
rect 1451 172 1462 206
rect 1406 138 1462 172
rect 1406 104 1417 138
rect 1451 104 1462 138
rect 1406 92 1462 104
rect 1492 1090 1548 1102
rect 1492 1056 1503 1090
rect 1537 1056 1548 1090
rect 1492 1022 1548 1056
rect 1492 988 1503 1022
rect 1537 988 1548 1022
rect 1492 954 1548 988
rect 1492 920 1503 954
rect 1537 920 1548 954
rect 1492 886 1548 920
rect 1492 852 1503 886
rect 1537 852 1548 886
rect 1492 818 1548 852
rect 1492 784 1503 818
rect 1537 784 1548 818
rect 1492 750 1548 784
rect 1492 716 1503 750
rect 1537 716 1548 750
rect 1492 682 1548 716
rect 1492 648 1503 682
rect 1537 648 1548 682
rect 1492 614 1548 648
rect 1492 580 1503 614
rect 1537 580 1548 614
rect 1492 546 1548 580
rect 1492 512 1503 546
rect 1537 512 1548 546
rect 1492 478 1548 512
rect 1492 444 1503 478
rect 1537 444 1548 478
rect 1492 410 1548 444
rect 1492 376 1503 410
rect 1537 376 1548 410
rect 1492 342 1548 376
rect 1492 308 1503 342
rect 1537 308 1548 342
rect 1492 274 1548 308
rect 1492 240 1503 274
rect 1537 240 1548 274
rect 1492 206 1548 240
rect 1492 172 1503 206
rect 1537 172 1548 206
rect 1492 138 1548 172
rect 1492 104 1503 138
rect 1537 104 1548 138
rect 1492 92 1548 104
<< ndiffc >>
rect 149 1056 183 1090
rect 149 988 183 1022
rect 149 920 183 954
rect 149 852 183 886
rect 149 784 183 818
rect 149 716 183 750
rect 149 648 183 682
rect 149 580 183 614
rect 149 512 183 546
rect 149 444 183 478
rect 149 376 183 410
rect 149 308 183 342
rect 149 240 183 274
rect 149 172 183 206
rect 149 104 183 138
rect 235 1056 269 1090
rect 235 988 269 1022
rect 235 920 269 954
rect 235 852 269 886
rect 235 784 269 818
rect 235 716 269 750
rect 235 648 269 682
rect 235 580 269 614
rect 235 512 269 546
rect 235 444 269 478
rect 235 376 269 410
rect 235 308 269 342
rect 235 240 269 274
rect 235 172 269 206
rect 235 104 269 138
rect 321 1056 355 1090
rect 321 988 355 1022
rect 321 920 355 954
rect 321 852 355 886
rect 321 784 355 818
rect 321 716 355 750
rect 321 648 355 682
rect 321 580 355 614
rect 321 512 355 546
rect 321 444 355 478
rect 321 376 355 410
rect 321 308 355 342
rect 321 240 355 274
rect 321 172 355 206
rect 321 104 355 138
rect 543 1056 577 1090
rect 543 988 577 1022
rect 543 920 577 954
rect 543 852 577 886
rect 543 784 577 818
rect 543 716 577 750
rect 543 648 577 682
rect 543 580 577 614
rect 543 512 577 546
rect 543 444 577 478
rect 543 376 577 410
rect 543 308 577 342
rect 543 240 577 274
rect 543 172 577 206
rect 543 104 577 138
rect 629 1056 663 1090
rect 629 988 663 1022
rect 629 920 663 954
rect 629 852 663 886
rect 629 784 663 818
rect 629 716 663 750
rect 629 648 663 682
rect 629 580 663 614
rect 629 512 663 546
rect 629 444 663 478
rect 629 376 663 410
rect 629 308 663 342
rect 629 240 663 274
rect 629 172 663 206
rect 629 104 663 138
rect 715 1056 749 1090
rect 715 988 749 1022
rect 715 920 749 954
rect 715 852 749 886
rect 715 784 749 818
rect 715 716 749 750
rect 715 648 749 682
rect 715 580 749 614
rect 715 512 749 546
rect 715 444 749 478
rect 715 376 749 410
rect 715 308 749 342
rect 715 240 749 274
rect 715 172 749 206
rect 715 104 749 138
rect 937 1056 971 1090
rect 937 988 971 1022
rect 937 920 971 954
rect 937 852 971 886
rect 937 784 971 818
rect 937 716 971 750
rect 937 648 971 682
rect 937 580 971 614
rect 937 512 971 546
rect 937 444 971 478
rect 937 376 971 410
rect 937 308 971 342
rect 937 240 971 274
rect 937 172 971 206
rect 937 104 971 138
rect 1023 1056 1057 1090
rect 1023 988 1057 1022
rect 1023 920 1057 954
rect 1023 852 1057 886
rect 1023 784 1057 818
rect 1023 716 1057 750
rect 1023 648 1057 682
rect 1023 580 1057 614
rect 1023 512 1057 546
rect 1023 444 1057 478
rect 1023 376 1057 410
rect 1023 308 1057 342
rect 1023 240 1057 274
rect 1023 172 1057 206
rect 1023 104 1057 138
rect 1109 1056 1143 1090
rect 1109 988 1143 1022
rect 1109 920 1143 954
rect 1109 852 1143 886
rect 1109 784 1143 818
rect 1109 716 1143 750
rect 1109 648 1143 682
rect 1109 580 1143 614
rect 1109 512 1143 546
rect 1109 444 1143 478
rect 1109 376 1143 410
rect 1109 308 1143 342
rect 1109 240 1143 274
rect 1109 172 1143 206
rect 1109 104 1143 138
rect 1331 1056 1365 1090
rect 1331 988 1365 1022
rect 1331 920 1365 954
rect 1331 852 1365 886
rect 1331 784 1365 818
rect 1331 716 1365 750
rect 1331 648 1365 682
rect 1331 580 1365 614
rect 1331 512 1365 546
rect 1331 444 1365 478
rect 1331 376 1365 410
rect 1331 308 1365 342
rect 1331 240 1365 274
rect 1331 172 1365 206
rect 1331 104 1365 138
rect 1417 1056 1451 1090
rect 1417 988 1451 1022
rect 1417 920 1451 954
rect 1417 852 1451 886
rect 1417 784 1451 818
rect 1417 716 1451 750
rect 1417 648 1451 682
rect 1417 580 1451 614
rect 1417 512 1451 546
rect 1417 444 1451 478
rect 1417 376 1451 410
rect 1417 308 1451 342
rect 1417 240 1451 274
rect 1417 172 1451 206
rect 1417 104 1451 138
rect 1503 1056 1537 1090
rect 1503 988 1537 1022
rect 1503 920 1537 954
rect 1503 852 1537 886
rect 1503 784 1537 818
rect 1503 716 1537 750
rect 1503 648 1537 682
rect 1503 580 1537 614
rect 1503 512 1537 546
rect 1503 444 1537 478
rect 1503 376 1537 410
rect 1503 308 1537 342
rect 1503 240 1537 274
rect 1503 172 1537 206
rect 1503 104 1537 138
<< psubdiff >>
rect 26 1056 84 1102
rect 26 1022 38 1056
rect 72 1022 84 1056
rect 26 988 84 1022
rect 26 954 38 988
rect 72 954 84 988
rect 26 920 84 954
rect 26 886 38 920
rect 72 886 84 920
rect 26 852 84 886
rect 26 818 38 852
rect 72 818 84 852
rect 26 784 84 818
rect 26 750 38 784
rect 72 750 84 784
rect 26 716 84 750
rect 26 682 38 716
rect 72 682 84 716
rect 26 648 84 682
rect 26 614 38 648
rect 72 614 84 648
rect 26 580 84 614
rect 26 546 38 580
rect 72 546 84 580
rect 26 512 84 546
rect 26 478 38 512
rect 72 478 84 512
rect 26 444 84 478
rect 26 410 38 444
rect 72 410 84 444
rect 26 376 84 410
rect 26 342 38 376
rect 72 342 84 376
rect 26 308 84 342
rect 26 274 38 308
rect 72 274 84 308
rect 26 240 84 274
rect 26 206 38 240
rect 72 206 84 240
rect 26 172 84 206
rect 26 138 38 172
rect 72 138 84 172
rect 26 92 84 138
rect 420 1056 478 1102
rect 420 1022 432 1056
rect 466 1022 478 1056
rect 420 988 478 1022
rect 420 954 432 988
rect 466 954 478 988
rect 420 920 478 954
rect 420 886 432 920
rect 466 886 478 920
rect 420 852 478 886
rect 420 818 432 852
rect 466 818 478 852
rect 420 784 478 818
rect 420 750 432 784
rect 466 750 478 784
rect 420 716 478 750
rect 420 682 432 716
rect 466 682 478 716
rect 420 648 478 682
rect 420 614 432 648
rect 466 614 478 648
rect 420 580 478 614
rect 420 546 432 580
rect 466 546 478 580
rect 420 512 478 546
rect 420 478 432 512
rect 466 478 478 512
rect 420 444 478 478
rect 420 410 432 444
rect 466 410 478 444
rect 420 376 478 410
rect 420 342 432 376
rect 466 342 478 376
rect 420 308 478 342
rect 420 274 432 308
rect 466 274 478 308
rect 420 240 478 274
rect 420 206 432 240
rect 466 206 478 240
rect 420 172 478 206
rect 420 138 432 172
rect 466 138 478 172
rect 420 92 478 138
rect 814 1056 872 1102
rect 814 1022 826 1056
rect 860 1022 872 1056
rect 814 988 872 1022
rect 814 954 826 988
rect 860 954 872 988
rect 814 920 872 954
rect 814 886 826 920
rect 860 886 872 920
rect 814 852 872 886
rect 814 818 826 852
rect 860 818 872 852
rect 814 784 872 818
rect 814 750 826 784
rect 860 750 872 784
rect 814 716 872 750
rect 814 682 826 716
rect 860 682 872 716
rect 814 648 872 682
rect 814 614 826 648
rect 860 614 872 648
rect 814 580 872 614
rect 814 546 826 580
rect 860 546 872 580
rect 814 512 872 546
rect 814 478 826 512
rect 860 478 872 512
rect 814 444 872 478
rect 814 410 826 444
rect 860 410 872 444
rect 814 376 872 410
rect 814 342 826 376
rect 860 342 872 376
rect 814 308 872 342
rect 814 274 826 308
rect 860 274 872 308
rect 814 240 872 274
rect 814 206 826 240
rect 860 206 872 240
rect 814 172 872 206
rect 814 138 826 172
rect 860 138 872 172
rect 814 92 872 138
rect 1208 1056 1266 1102
rect 1208 1022 1220 1056
rect 1254 1022 1266 1056
rect 1208 988 1266 1022
rect 1208 954 1220 988
rect 1254 954 1266 988
rect 1208 920 1266 954
rect 1208 886 1220 920
rect 1254 886 1266 920
rect 1208 852 1266 886
rect 1208 818 1220 852
rect 1254 818 1266 852
rect 1208 784 1266 818
rect 1208 750 1220 784
rect 1254 750 1266 784
rect 1208 716 1266 750
rect 1208 682 1220 716
rect 1254 682 1266 716
rect 1208 648 1266 682
rect 1208 614 1220 648
rect 1254 614 1266 648
rect 1208 580 1266 614
rect 1208 546 1220 580
rect 1254 546 1266 580
rect 1208 512 1266 546
rect 1208 478 1220 512
rect 1254 478 1266 512
rect 1208 444 1266 478
rect 1208 410 1220 444
rect 1254 410 1266 444
rect 1208 376 1266 410
rect 1208 342 1220 376
rect 1254 342 1266 376
rect 1208 308 1266 342
rect 1208 274 1220 308
rect 1254 274 1266 308
rect 1208 240 1266 274
rect 1208 206 1220 240
rect 1254 206 1266 240
rect 1208 172 1266 206
rect 1208 138 1220 172
rect 1254 138 1266 172
rect 1208 92 1266 138
rect 1602 1056 1660 1102
rect 1602 1022 1614 1056
rect 1648 1022 1660 1056
rect 1602 988 1660 1022
rect 1602 954 1614 988
rect 1648 954 1660 988
rect 1602 920 1660 954
rect 1602 886 1614 920
rect 1648 886 1660 920
rect 1602 852 1660 886
rect 1602 818 1614 852
rect 1648 818 1660 852
rect 1602 784 1660 818
rect 1602 750 1614 784
rect 1648 750 1660 784
rect 1602 716 1660 750
rect 1602 682 1614 716
rect 1648 682 1660 716
rect 1602 648 1660 682
rect 1602 614 1614 648
rect 1648 614 1660 648
rect 1602 580 1660 614
rect 1602 546 1614 580
rect 1648 546 1660 580
rect 1602 512 1660 546
rect 1602 478 1614 512
rect 1648 478 1660 512
rect 1602 444 1660 478
rect 1602 410 1614 444
rect 1648 410 1660 444
rect 1602 376 1660 410
rect 1602 342 1614 376
rect 1648 342 1660 376
rect 1602 308 1660 342
rect 1602 274 1614 308
rect 1648 274 1660 308
rect 1602 240 1660 274
rect 1602 206 1614 240
rect 1648 206 1660 240
rect 1602 172 1660 206
rect 1602 138 1614 172
rect 1648 138 1660 172
rect 1602 92 1660 138
<< psubdiffcont >>
rect 38 1022 72 1056
rect 38 954 72 988
rect 38 886 72 920
rect 38 818 72 852
rect 38 750 72 784
rect 38 682 72 716
rect 38 614 72 648
rect 38 546 72 580
rect 38 478 72 512
rect 38 410 72 444
rect 38 342 72 376
rect 38 274 72 308
rect 38 206 72 240
rect 38 138 72 172
rect 432 1022 466 1056
rect 432 954 466 988
rect 432 886 466 920
rect 432 818 466 852
rect 432 750 466 784
rect 432 682 466 716
rect 432 614 466 648
rect 432 546 466 580
rect 432 478 466 512
rect 432 410 466 444
rect 432 342 466 376
rect 432 274 466 308
rect 432 206 466 240
rect 432 138 466 172
rect 826 1022 860 1056
rect 826 954 860 988
rect 826 886 860 920
rect 826 818 860 852
rect 826 750 860 784
rect 826 682 860 716
rect 826 614 860 648
rect 826 546 860 580
rect 826 478 860 512
rect 826 410 860 444
rect 826 342 860 376
rect 826 274 860 308
rect 826 206 860 240
rect 826 138 860 172
rect 1220 1022 1254 1056
rect 1220 954 1254 988
rect 1220 886 1254 920
rect 1220 818 1254 852
rect 1220 750 1254 784
rect 1220 682 1254 716
rect 1220 614 1254 648
rect 1220 546 1254 580
rect 1220 478 1254 512
rect 1220 410 1254 444
rect 1220 342 1254 376
rect 1220 274 1254 308
rect 1220 206 1254 240
rect 1220 138 1254 172
rect 1614 1022 1648 1056
rect 1614 954 1648 988
rect 1614 886 1648 920
rect 1614 818 1648 852
rect 1614 750 1648 784
rect 1614 682 1648 716
rect 1614 614 1648 648
rect 1614 546 1648 580
rect 1614 478 1648 512
rect 1614 410 1648 444
rect 1614 342 1648 376
rect 1614 274 1648 308
rect 1614 206 1648 240
rect 1614 138 1648 172
<< poly >>
rect 151 1174 353 1194
rect 151 1140 167 1174
rect 201 1140 235 1174
rect 269 1140 303 1174
rect 337 1140 353 1174
rect 151 1124 353 1140
rect 545 1174 747 1194
rect 545 1140 561 1174
rect 595 1140 629 1174
rect 663 1140 697 1174
rect 731 1140 747 1174
rect 545 1124 747 1140
rect 939 1174 1141 1194
rect 939 1140 955 1174
rect 989 1140 1023 1174
rect 1057 1140 1091 1174
rect 1125 1140 1141 1174
rect 939 1124 1141 1140
rect 1333 1174 1535 1194
rect 1333 1140 1349 1174
rect 1383 1140 1417 1174
rect 1451 1140 1485 1174
rect 1519 1140 1535 1174
rect 1333 1124 1535 1140
rect 194 1102 224 1124
rect 280 1102 310 1124
rect 588 1102 618 1124
rect 674 1102 704 1124
rect 982 1102 1012 1124
rect 1068 1102 1098 1124
rect 1376 1102 1406 1124
rect 1462 1102 1492 1124
rect 194 70 224 92
rect 280 70 310 92
rect 588 70 618 92
rect 674 70 704 92
rect 982 70 1012 92
rect 1068 70 1098 92
rect 1376 70 1406 92
rect 1462 70 1492 92
rect 151 54 353 70
rect 151 20 167 54
rect 201 20 235 54
rect 269 20 303 54
rect 337 20 353 54
rect 151 0 353 20
rect 545 54 747 70
rect 545 20 561 54
rect 595 20 629 54
rect 663 20 697 54
rect 731 20 747 54
rect 545 0 747 20
rect 939 54 1141 70
rect 939 20 955 54
rect 989 20 1023 54
rect 1057 20 1091 54
rect 1125 20 1141 54
rect 939 0 1141 20
rect 1333 54 1535 70
rect 1333 20 1349 54
rect 1383 20 1417 54
rect 1451 20 1485 54
rect 1519 20 1535 54
rect 1333 0 1535 20
<< polycont >>
rect 167 1140 201 1174
rect 235 1140 269 1174
rect 303 1140 337 1174
rect 561 1140 595 1174
rect 629 1140 663 1174
rect 697 1140 731 1174
rect 955 1140 989 1174
rect 1023 1140 1057 1174
rect 1091 1140 1125 1174
rect 1349 1140 1383 1174
rect 1417 1140 1451 1174
rect 1485 1140 1519 1174
rect 167 20 201 54
rect 235 20 269 54
rect 303 20 337 54
rect 561 20 595 54
rect 629 20 663 54
rect 697 20 731 54
rect 955 20 989 54
rect 1023 20 1057 54
rect 1091 20 1125 54
rect 1349 20 1383 54
rect 1417 20 1451 54
rect 1485 20 1519 54
<< locali >>
rect 151 1140 163 1174
rect 201 1140 235 1174
rect 269 1140 303 1174
rect 341 1140 353 1174
rect 545 1140 557 1174
rect 595 1140 629 1174
rect 663 1140 697 1174
rect 735 1140 747 1174
rect 939 1140 951 1174
rect 989 1140 1023 1174
rect 1057 1140 1091 1174
rect 1129 1140 1141 1174
rect 1333 1140 1345 1174
rect 1383 1140 1417 1174
rect 1451 1140 1485 1174
rect 1523 1140 1535 1174
rect 149 1090 183 1106
rect 38 1010 72 1022
rect 38 938 72 954
rect 38 866 72 886
rect 38 794 72 818
rect 38 722 72 750
rect 38 650 72 682
rect 38 580 72 614
rect 38 512 72 544
rect 38 444 72 472
rect 38 376 72 400
rect 38 308 72 328
rect 38 240 72 256
rect 38 172 72 184
rect 149 1022 183 1048
rect 149 954 183 976
rect 149 886 183 904
rect 149 818 183 832
rect 149 750 183 760
rect 149 682 183 688
rect 149 614 183 616
rect 149 578 183 580
rect 149 506 183 512
rect 149 434 183 444
rect 149 362 183 376
rect 149 290 183 308
rect 149 218 183 240
rect 149 146 183 172
rect 149 88 183 104
rect 235 1090 269 1106
rect 235 1022 269 1048
rect 235 954 269 976
rect 235 886 269 904
rect 235 818 269 832
rect 235 750 269 760
rect 235 682 269 688
rect 235 614 269 616
rect 235 578 269 580
rect 235 506 269 512
rect 235 434 269 444
rect 235 362 269 376
rect 235 290 269 308
rect 235 218 269 240
rect 235 146 269 172
rect 235 88 269 104
rect 321 1090 355 1106
rect 543 1090 577 1106
rect 321 1022 355 1048
rect 321 954 355 976
rect 321 886 355 904
rect 321 818 355 832
rect 321 750 355 760
rect 321 682 355 688
rect 321 614 355 616
rect 321 578 355 580
rect 321 506 355 512
rect 321 434 355 444
rect 321 362 355 376
rect 321 290 355 308
rect 321 218 355 240
rect 321 146 355 172
rect 432 1010 466 1022
rect 432 938 466 954
rect 432 866 466 886
rect 432 794 466 818
rect 432 722 466 750
rect 432 650 466 682
rect 432 580 466 614
rect 432 512 466 544
rect 432 444 466 472
rect 432 376 466 400
rect 432 308 466 328
rect 432 240 466 256
rect 432 172 466 184
rect 543 1022 577 1048
rect 543 954 577 976
rect 543 886 577 904
rect 543 818 577 832
rect 543 750 577 760
rect 543 682 577 688
rect 543 614 577 616
rect 543 578 577 580
rect 543 506 577 512
rect 543 434 577 444
rect 543 362 577 376
rect 543 290 577 308
rect 543 218 577 240
rect 543 146 577 172
rect 321 88 355 104
rect 543 88 577 104
rect 629 1090 663 1106
rect 629 1022 663 1048
rect 629 954 663 976
rect 629 886 663 904
rect 629 818 663 832
rect 629 750 663 760
rect 629 682 663 688
rect 629 614 663 616
rect 629 578 663 580
rect 629 506 663 512
rect 629 434 663 444
rect 629 362 663 376
rect 629 290 663 308
rect 629 218 663 240
rect 629 146 663 172
rect 629 88 663 104
rect 715 1090 749 1106
rect 937 1090 971 1106
rect 715 1022 749 1048
rect 715 954 749 976
rect 715 886 749 904
rect 715 818 749 832
rect 715 750 749 760
rect 715 682 749 688
rect 715 614 749 616
rect 715 578 749 580
rect 715 506 749 512
rect 715 434 749 444
rect 715 362 749 376
rect 715 290 749 308
rect 715 218 749 240
rect 715 146 749 172
rect 826 1010 860 1022
rect 826 938 860 954
rect 826 866 860 886
rect 826 794 860 818
rect 826 722 860 750
rect 826 650 860 682
rect 826 580 860 614
rect 826 512 860 544
rect 826 444 860 472
rect 826 376 860 400
rect 826 308 860 328
rect 826 240 860 256
rect 826 172 860 184
rect 937 1022 971 1048
rect 937 954 971 976
rect 937 886 971 904
rect 937 818 971 832
rect 937 750 971 760
rect 937 682 971 688
rect 937 614 971 616
rect 937 578 971 580
rect 937 506 971 512
rect 937 434 971 444
rect 937 362 971 376
rect 937 290 971 308
rect 937 218 971 240
rect 937 146 971 172
rect 715 88 749 104
rect 937 88 971 104
rect 1023 1090 1057 1106
rect 1023 1022 1057 1048
rect 1023 954 1057 976
rect 1023 886 1057 904
rect 1023 818 1057 832
rect 1023 750 1057 760
rect 1023 682 1057 688
rect 1023 614 1057 616
rect 1023 578 1057 580
rect 1023 506 1057 512
rect 1023 434 1057 444
rect 1023 362 1057 376
rect 1023 290 1057 308
rect 1023 218 1057 240
rect 1023 146 1057 172
rect 1023 88 1057 104
rect 1109 1090 1143 1106
rect 1331 1090 1365 1106
rect 1109 1022 1143 1048
rect 1109 954 1143 976
rect 1109 886 1143 904
rect 1109 818 1143 832
rect 1109 750 1143 760
rect 1109 682 1143 688
rect 1109 614 1143 616
rect 1109 578 1143 580
rect 1109 506 1143 512
rect 1109 434 1143 444
rect 1109 362 1143 376
rect 1109 290 1143 308
rect 1109 218 1143 240
rect 1109 146 1143 172
rect 1220 1010 1254 1022
rect 1220 938 1254 954
rect 1220 866 1254 886
rect 1220 794 1254 818
rect 1220 722 1254 750
rect 1220 650 1254 682
rect 1220 580 1254 614
rect 1220 512 1254 544
rect 1220 444 1254 472
rect 1220 376 1254 400
rect 1220 308 1254 328
rect 1220 240 1254 256
rect 1220 172 1254 184
rect 1331 1022 1365 1048
rect 1331 954 1365 976
rect 1331 886 1365 904
rect 1331 818 1365 832
rect 1331 750 1365 760
rect 1331 682 1365 688
rect 1331 614 1365 616
rect 1331 578 1365 580
rect 1331 506 1365 512
rect 1331 434 1365 444
rect 1331 362 1365 376
rect 1331 290 1365 308
rect 1331 218 1365 240
rect 1331 146 1365 172
rect 1109 88 1143 104
rect 1331 88 1365 104
rect 1417 1090 1451 1106
rect 1417 1022 1451 1048
rect 1417 954 1451 976
rect 1417 886 1451 904
rect 1417 818 1451 832
rect 1417 750 1451 760
rect 1417 682 1451 688
rect 1417 614 1451 616
rect 1417 578 1451 580
rect 1417 506 1451 512
rect 1417 434 1451 444
rect 1417 362 1451 376
rect 1417 290 1451 308
rect 1417 218 1451 240
rect 1417 146 1451 172
rect 1417 88 1451 104
rect 1503 1090 1537 1106
rect 1503 1022 1537 1048
rect 1503 954 1537 976
rect 1503 886 1537 904
rect 1503 818 1537 832
rect 1503 750 1537 760
rect 1503 682 1537 688
rect 1503 614 1537 616
rect 1503 578 1537 580
rect 1503 506 1537 512
rect 1503 434 1537 444
rect 1503 362 1537 376
rect 1503 290 1537 308
rect 1503 218 1537 240
rect 1503 146 1537 172
rect 1614 1010 1648 1022
rect 1614 938 1648 954
rect 1614 866 1648 886
rect 1614 794 1648 818
rect 1614 722 1648 750
rect 1614 650 1648 682
rect 1614 580 1648 614
rect 1614 512 1648 544
rect 1614 444 1648 472
rect 1614 376 1648 400
rect 1614 308 1648 328
rect 1614 240 1648 256
rect 1614 172 1648 184
rect 1503 88 1537 104
rect 151 20 163 54
rect 201 20 235 54
rect 269 20 303 54
rect 341 20 353 54
rect 545 20 557 54
rect 595 20 629 54
rect 663 20 697 54
rect 735 20 747 54
rect 939 20 951 54
rect 989 20 1023 54
rect 1057 20 1091 54
rect 1129 20 1141 54
rect 1333 20 1345 54
rect 1383 20 1417 54
rect 1451 20 1485 54
rect 1523 20 1535 54
<< viali >>
rect 163 1140 167 1174
rect 167 1140 197 1174
rect 235 1140 269 1174
rect 307 1140 337 1174
rect 337 1140 341 1174
rect 557 1140 561 1174
rect 561 1140 591 1174
rect 629 1140 663 1174
rect 701 1140 731 1174
rect 731 1140 735 1174
rect 951 1140 955 1174
rect 955 1140 985 1174
rect 1023 1140 1057 1174
rect 1095 1140 1125 1174
rect 1125 1140 1129 1174
rect 1345 1140 1349 1174
rect 1349 1140 1379 1174
rect 1417 1140 1451 1174
rect 1489 1140 1519 1174
rect 1519 1140 1523 1174
rect 38 1056 72 1082
rect 38 1048 72 1056
rect 38 988 72 1010
rect 38 976 72 988
rect 38 920 72 938
rect 38 904 72 920
rect 38 852 72 866
rect 38 832 72 852
rect 38 784 72 794
rect 38 760 72 784
rect 38 716 72 722
rect 38 688 72 716
rect 38 648 72 650
rect 38 616 72 648
rect 38 546 72 578
rect 38 544 72 546
rect 38 478 72 506
rect 38 472 72 478
rect 38 410 72 434
rect 38 400 72 410
rect 38 342 72 362
rect 38 328 72 342
rect 38 274 72 290
rect 38 256 72 274
rect 38 206 72 218
rect 38 184 72 206
rect 38 138 72 146
rect 38 112 72 138
rect 149 1056 183 1082
rect 149 1048 183 1056
rect 149 988 183 1010
rect 149 976 183 988
rect 149 920 183 938
rect 149 904 183 920
rect 149 852 183 866
rect 149 832 183 852
rect 149 784 183 794
rect 149 760 183 784
rect 149 716 183 722
rect 149 688 183 716
rect 149 648 183 650
rect 149 616 183 648
rect 149 546 183 578
rect 149 544 183 546
rect 149 478 183 506
rect 149 472 183 478
rect 149 410 183 434
rect 149 400 183 410
rect 149 342 183 362
rect 149 328 183 342
rect 149 274 183 290
rect 149 256 183 274
rect 149 206 183 218
rect 149 184 183 206
rect 149 138 183 146
rect 149 112 183 138
rect 235 1056 269 1082
rect 235 1048 269 1056
rect 235 988 269 1010
rect 235 976 269 988
rect 235 920 269 938
rect 235 904 269 920
rect 235 852 269 866
rect 235 832 269 852
rect 235 784 269 794
rect 235 760 269 784
rect 235 716 269 722
rect 235 688 269 716
rect 235 648 269 650
rect 235 616 269 648
rect 235 546 269 578
rect 235 544 269 546
rect 235 478 269 506
rect 235 472 269 478
rect 235 410 269 434
rect 235 400 269 410
rect 235 342 269 362
rect 235 328 269 342
rect 235 274 269 290
rect 235 256 269 274
rect 235 206 269 218
rect 235 184 269 206
rect 235 138 269 146
rect 235 112 269 138
rect 321 1056 355 1082
rect 321 1048 355 1056
rect 321 988 355 1010
rect 321 976 355 988
rect 321 920 355 938
rect 321 904 355 920
rect 321 852 355 866
rect 321 832 355 852
rect 321 784 355 794
rect 321 760 355 784
rect 321 716 355 722
rect 321 688 355 716
rect 321 648 355 650
rect 321 616 355 648
rect 321 546 355 578
rect 321 544 355 546
rect 321 478 355 506
rect 321 472 355 478
rect 321 410 355 434
rect 321 400 355 410
rect 321 342 355 362
rect 321 328 355 342
rect 321 274 355 290
rect 321 256 355 274
rect 321 206 355 218
rect 321 184 355 206
rect 321 138 355 146
rect 321 112 355 138
rect 432 1056 466 1082
rect 432 1048 466 1056
rect 432 988 466 1010
rect 432 976 466 988
rect 432 920 466 938
rect 432 904 466 920
rect 432 852 466 866
rect 432 832 466 852
rect 432 784 466 794
rect 432 760 466 784
rect 432 716 466 722
rect 432 688 466 716
rect 432 648 466 650
rect 432 616 466 648
rect 432 546 466 578
rect 432 544 466 546
rect 432 478 466 506
rect 432 472 466 478
rect 432 410 466 434
rect 432 400 466 410
rect 432 342 466 362
rect 432 328 466 342
rect 432 274 466 290
rect 432 256 466 274
rect 432 206 466 218
rect 432 184 466 206
rect 432 138 466 146
rect 432 112 466 138
rect 543 1056 577 1082
rect 543 1048 577 1056
rect 543 988 577 1010
rect 543 976 577 988
rect 543 920 577 938
rect 543 904 577 920
rect 543 852 577 866
rect 543 832 577 852
rect 543 784 577 794
rect 543 760 577 784
rect 543 716 577 722
rect 543 688 577 716
rect 543 648 577 650
rect 543 616 577 648
rect 543 546 577 578
rect 543 544 577 546
rect 543 478 577 506
rect 543 472 577 478
rect 543 410 577 434
rect 543 400 577 410
rect 543 342 577 362
rect 543 328 577 342
rect 543 274 577 290
rect 543 256 577 274
rect 543 206 577 218
rect 543 184 577 206
rect 543 138 577 146
rect 543 112 577 138
rect 629 1056 663 1082
rect 629 1048 663 1056
rect 629 988 663 1010
rect 629 976 663 988
rect 629 920 663 938
rect 629 904 663 920
rect 629 852 663 866
rect 629 832 663 852
rect 629 784 663 794
rect 629 760 663 784
rect 629 716 663 722
rect 629 688 663 716
rect 629 648 663 650
rect 629 616 663 648
rect 629 546 663 578
rect 629 544 663 546
rect 629 478 663 506
rect 629 472 663 478
rect 629 410 663 434
rect 629 400 663 410
rect 629 342 663 362
rect 629 328 663 342
rect 629 274 663 290
rect 629 256 663 274
rect 629 206 663 218
rect 629 184 663 206
rect 629 138 663 146
rect 629 112 663 138
rect 715 1056 749 1082
rect 715 1048 749 1056
rect 715 988 749 1010
rect 715 976 749 988
rect 715 920 749 938
rect 715 904 749 920
rect 715 852 749 866
rect 715 832 749 852
rect 715 784 749 794
rect 715 760 749 784
rect 715 716 749 722
rect 715 688 749 716
rect 715 648 749 650
rect 715 616 749 648
rect 715 546 749 578
rect 715 544 749 546
rect 715 478 749 506
rect 715 472 749 478
rect 715 410 749 434
rect 715 400 749 410
rect 715 342 749 362
rect 715 328 749 342
rect 715 274 749 290
rect 715 256 749 274
rect 715 206 749 218
rect 715 184 749 206
rect 715 138 749 146
rect 715 112 749 138
rect 826 1056 860 1082
rect 826 1048 860 1056
rect 826 988 860 1010
rect 826 976 860 988
rect 826 920 860 938
rect 826 904 860 920
rect 826 852 860 866
rect 826 832 860 852
rect 826 784 860 794
rect 826 760 860 784
rect 826 716 860 722
rect 826 688 860 716
rect 826 648 860 650
rect 826 616 860 648
rect 826 546 860 578
rect 826 544 860 546
rect 826 478 860 506
rect 826 472 860 478
rect 826 410 860 434
rect 826 400 860 410
rect 826 342 860 362
rect 826 328 860 342
rect 826 274 860 290
rect 826 256 860 274
rect 826 206 860 218
rect 826 184 860 206
rect 826 138 860 146
rect 826 112 860 138
rect 937 1056 971 1082
rect 937 1048 971 1056
rect 937 988 971 1010
rect 937 976 971 988
rect 937 920 971 938
rect 937 904 971 920
rect 937 852 971 866
rect 937 832 971 852
rect 937 784 971 794
rect 937 760 971 784
rect 937 716 971 722
rect 937 688 971 716
rect 937 648 971 650
rect 937 616 971 648
rect 937 546 971 578
rect 937 544 971 546
rect 937 478 971 506
rect 937 472 971 478
rect 937 410 971 434
rect 937 400 971 410
rect 937 342 971 362
rect 937 328 971 342
rect 937 274 971 290
rect 937 256 971 274
rect 937 206 971 218
rect 937 184 971 206
rect 937 138 971 146
rect 937 112 971 138
rect 1023 1056 1057 1082
rect 1023 1048 1057 1056
rect 1023 988 1057 1010
rect 1023 976 1057 988
rect 1023 920 1057 938
rect 1023 904 1057 920
rect 1023 852 1057 866
rect 1023 832 1057 852
rect 1023 784 1057 794
rect 1023 760 1057 784
rect 1023 716 1057 722
rect 1023 688 1057 716
rect 1023 648 1057 650
rect 1023 616 1057 648
rect 1023 546 1057 578
rect 1023 544 1057 546
rect 1023 478 1057 506
rect 1023 472 1057 478
rect 1023 410 1057 434
rect 1023 400 1057 410
rect 1023 342 1057 362
rect 1023 328 1057 342
rect 1023 274 1057 290
rect 1023 256 1057 274
rect 1023 206 1057 218
rect 1023 184 1057 206
rect 1023 138 1057 146
rect 1023 112 1057 138
rect 1109 1056 1143 1082
rect 1109 1048 1143 1056
rect 1109 988 1143 1010
rect 1109 976 1143 988
rect 1109 920 1143 938
rect 1109 904 1143 920
rect 1109 852 1143 866
rect 1109 832 1143 852
rect 1109 784 1143 794
rect 1109 760 1143 784
rect 1109 716 1143 722
rect 1109 688 1143 716
rect 1109 648 1143 650
rect 1109 616 1143 648
rect 1109 546 1143 578
rect 1109 544 1143 546
rect 1109 478 1143 506
rect 1109 472 1143 478
rect 1109 410 1143 434
rect 1109 400 1143 410
rect 1109 342 1143 362
rect 1109 328 1143 342
rect 1109 274 1143 290
rect 1109 256 1143 274
rect 1109 206 1143 218
rect 1109 184 1143 206
rect 1109 138 1143 146
rect 1109 112 1143 138
rect 1220 1056 1254 1082
rect 1220 1048 1254 1056
rect 1220 988 1254 1010
rect 1220 976 1254 988
rect 1220 920 1254 938
rect 1220 904 1254 920
rect 1220 852 1254 866
rect 1220 832 1254 852
rect 1220 784 1254 794
rect 1220 760 1254 784
rect 1220 716 1254 722
rect 1220 688 1254 716
rect 1220 648 1254 650
rect 1220 616 1254 648
rect 1220 546 1254 578
rect 1220 544 1254 546
rect 1220 478 1254 506
rect 1220 472 1254 478
rect 1220 410 1254 434
rect 1220 400 1254 410
rect 1220 342 1254 362
rect 1220 328 1254 342
rect 1220 274 1254 290
rect 1220 256 1254 274
rect 1220 206 1254 218
rect 1220 184 1254 206
rect 1220 138 1254 146
rect 1220 112 1254 138
rect 1331 1056 1365 1082
rect 1331 1048 1365 1056
rect 1331 988 1365 1010
rect 1331 976 1365 988
rect 1331 920 1365 938
rect 1331 904 1365 920
rect 1331 852 1365 866
rect 1331 832 1365 852
rect 1331 784 1365 794
rect 1331 760 1365 784
rect 1331 716 1365 722
rect 1331 688 1365 716
rect 1331 648 1365 650
rect 1331 616 1365 648
rect 1331 546 1365 578
rect 1331 544 1365 546
rect 1331 478 1365 506
rect 1331 472 1365 478
rect 1331 410 1365 434
rect 1331 400 1365 410
rect 1331 342 1365 362
rect 1331 328 1365 342
rect 1331 274 1365 290
rect 1331 256 1365 274
rect 1331 206 1365 218
rect 1331 184 1365 206
rect 1331 138 1365 146
rect 1331 112 1365 138
rect 1417 1056 1451 1082
rect 1417 1048 1451 1056
rect 1417 988 1451 1010
rect 1417 976 1451 988
rect 1417 920 1451 938
rect 1417 904 1451 920
rect 1417 852 1451 866
rect 1417 832 1451 852
rect 1417 784 1451 794
rect 1417 760 1451 784
rect 1417 716 1451 722
rect 1417 688 1451 716
rect 1417 648 1451 650
rect 1417 616 1451 648
rect 1417 546 1451 578
rect 1417 544 1451 546
rect 1417 478 1451 506
rect 1417 472 1451 478
rect 1417 410 1451 434
rect 1417 400 1451 410
rect 1417 342 1451 362
rect 1417 328 1451 342
rect 1417 274 1451 290
rect 1417 256 1451 274
rect 1417 206 1451 218
rect 1417 184 1451 206
rect 1417 138 1451 146
rect 1417 112 1451 138
rect 1503 1056 1537 1082
rect 1503 1048 1537 1056
rect 1503 988 1537 1010
rect 1503 976 1537 988
rect 1503 920 1537 938
rect 1503 904 1537 920
rect 1503 852 1537 866
rect 1503 832 1537 852
rect 1503 784 1537 794
rect 1503 760 1537 784
rect 1503 716 1537 722
rect 1503 688 1537 716
rect 1503 648 1537 650
rect 1503 616 1537 648
rect 1503 546 1537 578
rect 1503 544 1537 546
rect 1503 478 1537 506
rect 1503 472 1537 478
rect 1503 410 1537 434
rect 1503 400 1537 410
rect 1503 342 1537 362
rect 1503 328 1537 342
rect 1503 274 1537 290
rect 1503 256 1537 274
rect 1503 206 1537 218
rect 1503 184 1537 206
rect 1503 138 1537 146
rect 1503 112 1537 138
rect 1614 1056 1648 1082
rect 1614 1048 1648 1056
rect 1614 988 1648 1010
rect 1614 976 1648 988
rect 1614 920 1648 938
rect 1614 904 1648 920
rect 1614 852 1648 866
rect 1614 832 1648 852
rect 1614 784 1648 794
rect 1614 760 1648 784
rect 1614 716 1648 722
rect 1614 688 1648 716
rect 1614 648 1648 650
rect 1614 616 1648 648
rect 1614 546 1648 578
rect 1614 544 1648 546
rect 1614 478 1648 506
rect 1614 472 1648 478
rect 1614 410 1648 434
rect 1614 400 1648 410
rect 1614 342 1648 362
rect 1614 328 1648 342
rect 1614 274 1648 290
rect 1614 256 1648 274
rect 1614 206 1648 218
rect 1614 184 1648 206
rect 1614 138 1648 146
rect 1614 112 1648 138
rect 163 20 167 54
rect 167 20 197 54
rect 235 20 269 54
rect 307 20 337 54
rect 337 20 341 54
rect 557 20 561 54
rect 561 20 591 54
rect 629 20 663 54
rect 701 20 731 54
rect 731 20 735 54
rect 951 20 955 54
rect 955 20 985 54
rect 1023 20 1057 54
rect 1095 20 1125 54
rect 1125 20 1129 54
rect 1345 20 1349 54
rect 1349 20 1379 54
rect 1417 20 1451 54
rect 1489 20 1519 54
rect 1519 20 1523 54
<< metal1 >>
rect 20 1094 80 1280
rect 140 1240 360 1260
rect 140 1160 160 1240
rect 340 1174 360 1240
rect 140 1140 163 1160
rect 197 1140 235 1160
rect 269 1140 307 1160
rect 341 1140 360 1174
rect 151 1128 353 1140
rect 20 1082 84 1094
rect 20 1048 38 1082
rect 72 1048 84 1082
rect 20 1010 84 1048
rect 20 976 38 1010
rect 72 976 84 1010
rect 20 938 84 976
rect 20 904 38 938
rect 72 904 84 938
rect 20 866 84 904
rect 20 832 38 866
rect 72 832 84 866
rect 20 794 84 832
rect 20 760 38 794
rect 72 760 84 794
rect 20 722 84 760
rect 20 688 38 722
rect 72 688 84 722
rect 20 650 84 688
rect 20 616 38 650
rect 72 616 84 650
rect 20 578 84 616
rect 20 544 38 578
rect 72 544 84 578
rect 20 506 84 544
rect 20 472 38 506
rect 72 472 84 506
rect 20 434 84 472
rect 20 400 38 434
rect 72 400 84 434
rect 20 362 84 400
rect 20 328 38 362
rect 72 328 84 362
rect 20 290 84 328
rect 20 256 38 290
rect 72 256 84 290
rect 20 218 84 256
rect 20 184 38 218
rect 72 184 84 218
rect 20 146 84 184
rect 20 112 38 146
rect 72 112 84 146
rect 20 100 84 112
rect 140 1082 192 1094
rect 140 1048 149 1082
rect 183 1048 192 1082
rect 140 1010 192 1048
rect 140 976 149 1010
rect 183 976 192 1010
rect 140 938 192 976
rect 140 904 149 938
rect 183 904 192 938
rect 140 866 192 904
rect 140 832 149 866
rect 183 832 192 866
rect 140 794 192 832
rect 140 760 149 794
rect 183 760 192 794
rect 140 722 192 760
rect 140 688 149 722
rect 183 688 192 722
rect 140 650 192 688
rect 140 616 149 650
rect 183 616 192 650
rect 140 578 192 616
rect 140 544 149 578
rect 183 544 192 578
rect 140 542 192 544
rect 140 478 149 490
rect 183 478 192 490
rect 140 414 149 426
rect 183 414 192 426
rect 140 350 149 362
rect 183 350 192 362
rect 140 290 192 298
rect 140 286 149 290
rect 183 286 192 290
rect 140 222 192 234
rect 140 158 192 170
rect 140 100 192 106
rect 226 1088 278 1094
rect 226 1024 278 1036
rect 226 960 278 972
rect 226 904 235 908
rect 269 904 278 908
rect 226 896 278 904
rect 226 832 235 844
rect 269 832 278 844
rect 226 768 235 780
rect 269 768 278 780
rect 226 704 235 716
rect 269 704 278 716
rect 226 650 278 652
rect 226 616 235 650
rect 269 616 278 650
rect 226 578 278 616
rect 226 544 235 578
rect 269 544 278 578
rect 226 506 278 544
rect 226 472 235 506
rect 269 472 278 506
rect 226 434 278 472
rect 226 400 235 434
rect 269 400 278 434
rect 226 362 278 400
rect 226 328 235 362
rect 269 328 278 362
rect 226 290 278 328
rect 226 256 235 290
rect 269 256 278 290
rect 226 218 278 256
rect 226 184 235 218
rect 269 184 278 218
rect 226 146 278 184
rect 226 112 235 146
rect 269 112 278 146
rect 226 100 278 112
rect 312 1082 364 1094
rect 312 1048 321 1082
rect 355 1048 364 1082
rect 312 1010 364 1048
rect 312 976 321 1010
rect 355 976 364 1010
rect 312 938 364 976
rect 312 904 321 938
rect 355 904 364 938
rect 312 866 364 904
rect 312 832 321 866
rect 355 832 364 866
rect 312 794 364 832
rect 312 760 321 794
rect 355 760 364 794
rect 312 722 364 760
rect 312 688 321 722
rect 355 688 364 722
rect 312 650 364 688
rect 312 616 321 650
rect 355 616 364 650
rect 312 578 364 616
rect 312 544 321 578
rect 355 544 364 578
rect 312 542 364 544
rect 312 478 321 490
rect 355 478 364 490
rect 312 414 321 426
rect 355 414 364 426
rect 312 350 321 362
rect 355 350 364 362
rect 312 290 364 298
rect 312 286 321 290
rect 355 286 364 290
rect 312 222 364 234
rect 312 158 364 170
rect 312 100 364 106
rect 420 1082 480 1280
rect 540 1240 760 1260
rect 540 1174 560 1240
rect 540 1140 557 1174
rect 740 1160 760 1240
rect 591 1140 629 1160
rect 663 1140 701 1160
rect 735 1140 760 1160
rect 545 1128 747 1140
rect 820 1094 880 1280
rect 940 1240 1160 1260
rect 940 1194 960 1240
rect 939 1174 960 1194
rect 939 1140 951 1174
rect 1140 1160 1160 1240
rect 985 1140 1023 1160
rect 1057 1140 1095 1160
rect 1129 1140 1160 1160
rect 939 1128 1141 1140
rect 1200 1094 1260 1280
rect 1320 1240 1540 1260
rect 1320 1160 1340 1240
rect 1520 1174 1540 1240
rect 1320 1140 1345 1160
rect 1379 1140 1417 1160
rect 1451 1140 1489 1160
rect 1523 1140 1540 1174
rect 1333 1128 1535 1140
rect 420 1048 432 1082
rect 466 1048 480 1082
rect 420 1010 480 1048
rect 420 976 432 1010
rect 466 976 480 1010
rect 420 938 480 976
rect 420 904 432 938
rect 466 904 480 938
rect 420 866 480 904
rect 420 832 432 866
rect 466 832 480 866
rect 420 794 480 832
rect 420 760 432 794
rect 466 760 480 794
rect 420 722 480 760
rect 420 688 432 722
rect 466 688 480 722
rect 420 650 480 688
rect 420 616 432 650
rect 466 616 480 650
rect 420 578 480 616
rect 420 544 432 578
rect 466 544 480 578
rect 420 506 480 544
rect 420 472 432 506
rect 466 472 480 506
rect 420 434 480 472
rect 420 400 432 434
rect 466 400 480 434
rect 420 362 480 400
rect 420 328 432 362
rect 466 328 480 362
rect 420 290 480 328
rect 420 256 432 290
rect 466 256 480 290
rect 420 218 480 256
rect 420 184 432 218
rect 466 184 480 218
rect 420 146 480 184
rect 420 112 432 146
rect 466 112 480 146
rect 20 -80 80 100
rect 151 54 353 66
rect 151 20 163 54
rect 197 20 235 54
rect 269 20 307 54
rect 341 20 353 54
rect 151 0 353 20
rect 420 -80 480 112
rect 534 1082 586 1094
rect 534 1048 543 1082
rect 577 1048 586 1082
rect 534 1010 586 1048
rect 534 976 543 1010
rect 577 976 586 1010
rect 534 938 586 976
rect 534 904 543 938
rect 577 904 586 938
rect 534 866 586 904
rect 534 832 543 866
rect 577 832 586 866
rect 534 794 586 832
rect 534 760 543 794
rect 577 760 586 794
rect 534 722 586 760
rect 534 688 543 722
rect 577 688 586 722
rect 534 650 586 688
rect 534 616 543 650
rect 577 616 586 650
rect 534 578 586 616
rect 534 544 543 578
rect 577 544 586 578
rect 534 542 586 544
rect 534 478 543 490
rect 577 478 586 490
rect 534 414 543 426
rect 577 414 586 426
rect 534 350 543 362
rect 577 350 586 362
rect 534 290 586 298
rect 534 286 543 290
rect 577 286 586 290
rect 534 222 586 234
rect 534 158 586 170
rect 534 100 586 106
rect 620 1088 672 1094
rect 620 1024 672 1036
rect 620 960 672 972
rect 620 904 629 908
rect 663 904 672 908
rect 620 896 672 904
rect 620 832 629 844
rect 663 832 672 844
rect 620 768 629 780
rect 663 768 672 780
rect 620 704 629 716
rect 663 704 672 716
rect 620 650 672 652
rect 620 616 629 650
rect 663 616 672 650
rect 620 578 672 616
rect 620 544 629 578
rect 663 544 672 578
rect 620 506 672 544
rect 620 472 629 506
rect 663 472 672 506
rect 620 434 672 472
rect 620 400 629 434
rect 663 400 672 434
rect 620 362 672 400
rect 620 328 629 362
rect 663 328 672 362
rect 620 290 672 328
rect 620 256 629 290
rect 663 256 672 290
rect 620 218 672 256
rect 620 184 629 218
rect 663 184 672 218
rect 620 146 672 184
rect 620 112 629 146
rect 663 112 672 146
rect 620 100 672 112
rect 706 1082 758 1094
rect 706 1048 715 1082
rect 749 1048 758 1082
rect 706 1010 758 1048
rect 706 976 715 1010
rect 749 976 758 1010
rect 706 938 758 976
rect 706 904 715 938
rect 749 904 758 938
rect 706 866 758 904
rect 706 832 715 866
rect 749 832 758 866
rect 706 794 758 832
rect 706 760 715 794
rect 749 760 758 794
rect 706 722 758 760
rect 706 688 715 722
rect 749 688 758 722
rect 706 650 758 688
rect 706 616 715 650
rect 749 616 758 650
rect 706 578 758 616
rect 706 544 715 578
rect 749 544 758 578
rect 706 542 758 544
rect 706 478 715 490
rect 749 478 758 490
rect 706 414 715 426
rect 749 414 758 426
rect 706 350 715 362
rect 749 350 758 362
rect 706 290 758 298
rect 706 286 715 290
rect 749 286 758 290
rect 706 222 758 234
rect 706 158 758 170
rect 706 100 758 106
rect 814 1082 880 1094
rect 814 1048 826 1082
rect 860 1048 880 1082
rect 814 1010 880 1048
rect 814 976 826 1010
rect 860 976 880 1010
rect 814 938 880 976
rect 814 904 826 938
rect 860 904 880 938
rect 814 866 880 904
rect 814 832 826 866
rect 860 832 880 866
rect 814 794 880 832
rect 814 760 826 794
rect 860 760 880 794
rect 814 722 880 760
rect 814 688 826 722
rect 860 688 880 722
rect 814 650 880 688
rect 814 616 826 650
rect 860 616 880 650
rect 814 578 880 616
rect 814 544 826 578
rect 860 544 880 578
rect 814 506 880 544
rect 814 472 826 506
rect 860 472 880 506
rect 814 434 880 472
rect 814 400 826 434
rect 860 400 880 434
rect 814 362 880 400
rect 814 328 826 362
rect 860 328 880 362
rect 814 290 880 328
rect 814 256 826 290
rect 860 256 880 290
rect 814 218 880 256
rect 814 184 826 218
rect 860 184 880 218
rect 814 146 880 184
rect 814 112 826 146
rect 860 112 880 146
rect 814 100 880 112
rect 928 1082 980 1094
rect 928 1048 937 1082
rect 971 1048 980 1082
rect 928 1010 980 1048
rect 928 976 937 1010
rect 971 976 980 1010
rect 928 938 980 976
rect 928 904 937 938
rect 971 904 980 938
rect 928 866 980 904
rect 928 832 937 866
rect 971 832 980 866
rect 928 794 980 832
rect 928 760 937 794
rect 971 760 980 794
rect 928 722 980 760
rect 928 688 937 722
rect 971 688 980 722
rect 928 650 980 688
rect 928 616 937 650
rect 971 616 980 650
rect 928 578 980 616
rect 928 544 937 578
rect 971 544 980 578
rect 928 542 980 544
rect 928 478 937 490
rect 971 478 980 490
rect 928 414 937 426
rect 971 414 980 426
rect 928 350 937 362
rect 971 350 980 362
rect 928 290 980 298
rect 928 286 937 290
rect 971 286 980 290
rect 928 222 980 234
rect 928 158 980 170
rect 928 100 980 106
rect 1014 1088 1066 1094
rect 1014 1024 1066 1036
rect 1014 960 1066 972
rect 1014 904 1023 908
rect 1057 904 1066 908
rect 1014 896 1066 904
rect 1014 832 1023 844
rect 1057 832 1066 844
rect 1014 768 1023 780
rect 1057 768 1066 780
rect 1014 704 1023 716
rect 1057 704 1066 716
rect 1014 650 1066 652
rect 1014 616 1023 650
rect 1057 616 1066 650
rect 1014 578 1066 616
rect 1014 544 1023 578
rect 1057 544 1066 578
rect 1014 506 1066 544
rect 1014 472 1023 506
rect 1057 472 1066 506
rect 1014 434 1066 472
rect 1014 400 1023 434
rect 1057 400 1066 434
rect 1014 362 1066 400
rect 1014 328 1023 362
rect 1057 328 1066 362
rect 1014 290 1066 328
rect 1014 256 1023 290
rect 1057 256 1066 290
rect 1014 218 1066 256
rect 1014 184 1023 218
rect 1057 184 1066 218
rect 1014 146 1066 184
rect 1014 112 1023 146
rect 1057 112 1066 146
rect 1014 100 1066 112
rect 1100 1082 1152 1094
rect 1100 1048 1109 1082
rect 1143 1048 1152 1082
rect 1100 1010 1152 1048
rect 1100 976 1109 1010
rect 1143 976 1152 1010
rect 1100 938 1152 976
rect 1100 904 1109 938
rect 1143 904 1152 938
rect 1100 866 1152 904
rect 1100 832 1109 866
rect 1143 832 1152 866
rect 1100 794 1152 832
rect 1100 760 1109 794
rect 1143 760 1152 794
rect 1100 722 1152 760
rect 1100 688 1109 722
rect 1143 688 1152 722
rect 1100 650 1152 688
rect 1100 616 1109 650
rect 1143 616 1152 650
rect 1100 578 1152 616
rect 1100 544 1109 578
rect 1143 544 1152 578
rect 1100 542 1152 544
rect 1100 478 1109 490
rect 1143 478 1152 490
rect 1100 414 1109 426
rect 1143 414 1152 426
rect 1100 350 1109 362
rect 1143 350 1152 362
rect 1100 290 1152 298
rect 1100 286 1109 290
rect 1143 286 1152 290
rect 1100 222 1152 234
rect 1100 158 1152 170
rect 1100 100 1152 106
rect 1200 1082 1266 1094
rect 1200 1048 1220 1082
rect 1254 1048 1266 1082
rect 1200 1010 1266 1048
rect 1200 976 1220 1010
rect 1254 976 1266 1010
rect 1200 938 1266 976
rect 1200 904 1220 938
rect 1254 904 1266 938
rect 1200 866 1266 904
rect 1200 832 1220 866
rect 1254 832 1266 866
rect 1200 794 1266 832
rect 1200 760 1220 794
rect 1254 760 1266 794
rect 1200 722 1266 760
rect 1200 688 1220 722
rect 1254 688 1266 722
rect 1200 650 1266 688
rect 1200 616 1220 650
rect 1254 616 1266 650
rect 1200 578 1266 616
rect 1200 544 1220 578
rect 1254 544 1266 578
rect 1200 506 1266 544
rect 1200 472 1220 506
rect 1254 472 1266 506
rect 1200 434 1266 472
rect 1200 400 1220 434
rect 1254 400 1266 434
rect 1200 362 1266 400
rect 1200 328 1220 362
rect 1254 328 1266 362
rect 1200 290 1266 328
rect 1200 256 1220 290
rect 1254 256 1266 290
rect 1200 218 1266 256
rect 1200 184 1220 218
rect 1254 184 1266 218
rect 1200 146 1266 184
rect 1200 112 1220 146
rect 1254 112 1266 146
rect 1200 100 1266 112
rect 1322 1082 1374 1094
rect 1322 1048 1331 1082
rect 1365 1048 1374 1082
rect 1322 1010 1374 1048
rect 1322 976 1331 1010
rect 1365 976 1374 1010
rect 1322 938 1374 976
rect 1322 904 1331 938
rect 1365 904 1374 938
rect 1322 866 1374 904
rect 1322 832 1331 866
rect 1365 832 1374 866
rect 1322 794 1374 832
rect 1322 760 1331 794
rect 1365 760 1374 794
rect 1322 722 1374 760
rect 1322 688 1331 722
rect 1365 688 1374 722
rect 1322 650 1374 688
rect 1322 616 1331 650
rect 1365 616 1374 650
rect 1322 578 1374 616
rect 1322 544 1331 578
rect 1365 544 1374 578
rect 1322 542 1374 544
rect 1322 478 1331 490
rect 1365 478 1374 490
rect 1322 414 1331 426
rect 1365 414 1374 426
rect 1322 350 1331 362
rect 1365 350 1374 362
rect 1322 290 1374 298
rect 1322 286 1331 290
rect 1365 286 1374 290
rect 1322 222 1374 234
rect 1322 158 1374 170
rect 1322 100 1374 106
rect 1408 1088 1460 1094
rect 1408 1024 1460 1036
rect 1408 960 1460 972
rect 1408 904 1417 908
rect 1451 904 1460 908
rect 1408 896 1460 904
rect 1408 832 1417 844
rect 1451 832 1460 844
rect 1408 768 1417 780
rect 1451 768 1460 780
rect 1408 704 1417 716
rect 1451 704 1460 716
rect 1408 650 1460 652
rect 1408 616 1417 650
rect 1451 616 1460 650
rect 1408 578 1460 616
rect 1408 544 1417 578
rect 1451 544 1460 578
rect 1408 506 1460 544
rect 1408 472 1417 506
rect 1451 472 1460 506
rect 1408 434 1460 472
rect 1408 400 1417 434
rect 1451 400 1460 434
rect 1408 362 1460 400
rect 1408 328 1417 362
rect 1451 328 1460 362
rect 1408 290 1460 328
rect 1408 256 1417 290
rect 1451 256 1460 290
rect 1408 218 1460 256
rect 1408 184 1417 218
rect 1451 184 1460 218
rect 1408 146 1460 184
rect 1408 112 1417 146
rect 1451 112 1460 146
rect 1408 100 1460 112
rect 1494 1082 1546 1094
rect 1494 1048 1503 1082
rect 1537 1048 1546 1082
rect 1494 1010 1546 1048
rect 1494 976 1503 1010
rect 1537 976 1546 1010
rect 1494 938 1546 976
rect 1494 904 1503 938
rect 1537 904 1546 938
rect 1494 866 1546 904
rect 1494 832 1503 866
rect 1537 832 1546 866
rect 1494 794 1546 832
rect 1494 760 1503 794
rect 1537 760 1546 794
rect 1494 722 1546 760
rect 1494 688 1503 722
rect 1537 688 1546 722
rect 1494 650 1546 688
rect 1494 616 1503 650
rect 1537 616 1546 650
rect 1494 578 1546 616
rect 1494 544 1503 578
rect 1537 544 1546 578
rect 1494 542 1546 544
rect 1494 478 1503 490
rect 1537 478 1546 490
rect 1494 414 1503 426
rect 1537 414 1546 426
rect 1494 350 1503 362
rect 1537 350 1546 362
rect 1494 290 1546 298
rect 1494 286 1503 290
rect 1537 286 1546 290
rect 1494 222 1546 234
rect 1494 158 1546 170
rect 1494 100 1546 106
rect 1600 1082 1660 1280
rect 1600 1048 1614 1082
rect 1648 1048 1660 1082
rect 1600 1010 1660 1048
rect 1600 976 1614 1010
rect 1648 976 1660 1010
rect 1600 938 1660 976
rect 1600 904 1614 938
rect 1648 904 1660 938
rect 1600 866 1660 904
rect 1600 832 1614 866
rect 1648 832 1660 866
rect 1600 794 1660 832
rect 1600 760 1614 794
rect 1648 760 1660 794
rect 1600 722 1660 760
rect 1600 688 1614 722
rect 1648 688 1660 722
rect 1600 650 1660 688
rect 1600 616 1614 650
rect 1648 616 1660 650
rect 1600 578 1660 616
rect 1600 544 1614 578
rect 1648 544 1660 578
rect 1600 506 1660 544
rect 1600 472 1614 506
rect 1648 472 1660 506
rect 1600 434 1660 472
rect 1600 400 1614 434
rect 1648 400 1660 434
rect 1600 362 1660 400
rect 1600 328 1614 362
rect 1648 328 1660 362
rect 1600 290 1660 328
rect 1600 256 1614 290
rect 1648 256 1660 290
rect 1600 218 1660 256
rect 1600 184 1614 218
rect 1648 184 1660 218
rect 1600 146 1660 184
rect 1600 112 1614 146
rect 1648 112 1660 146
rect 545 54 747 66
rect 545 20 557 54
rect 591 20 629 54
rect 663 20 701 54
rect 735 20 747 54
rect 545 0 747 20
rect 820 -80 880 100
rect 939 54 1141 66
rect 939 20 951 54
rect 985 20 1023 54
rect 1057 20 1095 54
rect 1129 20 1141 54
rect 939 0 1141 20
rect 1200 -80 1260 100
rect 1333 54 1535 66
rect 1333 20 1345 54
rect 1379 20 1417 54
rect 1451 20 1489 54
rect 1523 20 1535 54
rect 1333 0 1535 20
rect 1600 -80 1660 112
rect 20 -100 1660 -80
rect 20 -180 120 -100
rect 400 -180 860 -100
rect 1580 -180 1660 -100
rect 20 -200 1660 -180
<< via1 >>
rect 160 1174 340 1240
rect 160 1160 163 1174
rect 163 1160 197 1174
rect 197 1160 235 1174
rect 235 1160 269 1174
rect 269 1160 307 1174
rect 307 1160 340 1174
rect 140 506 192 542
rect 140 490 149 506
rect 149 490 183 506
rect 183 490 192 506
rect 140 472 149 478
rect 149 472 183 478
rect 183 472 192 478
rect 140 434 192 472
rect 140 426 149 434
rect 149 426 183 434
rect 183 426 192 434
rect 140 400 149 414
rect 149 400 183 414
rect 183 400 192 414
rect 140 362 192 400
rect 140 328 149 350
rect 149 328 183 350
rect 183 328 192 350
rect 140 298 192 328
rect 140 256 149 286
rect 149 256 183 286
rect 183 256 192 286
rect 140 234 192 256
rect 140 218 192 222
rect 140 184 149 218
rect 149 184 183 218
rect 183 184 192 218
rect 140 170 192 184
rect 140 146 192 158
rect 140 112 149 146
rect 149 112 183 146
rect 183 112 192 146
rect 140 106 192 112
rect 226 1082 278 1088
rect 226 1048 235 1082
rect 235 1048 269 1082
rect 269 1048 278 1082
rect 226 1036 278 1048
rect 226 1010 278 1024
rect 226 976 235 1010
rect 235 976 269 1010
rect 269 976 278 1010
rect 226 972 278 976
rect 226 938 278 960
rect 226 908 235 938
rect 235 908 269 938
rect 269 908 278 938
rect 226 866 278 896
rect 226 844 235 866
rect 235 844 269 866
rect 269 844 278 866
rect 226 794 278 832
rect 226 780 235 794
rect 235 780 269 794
rect 269 780 278 794
rect 226 760 235 768
rect 235 760 269 768
rect 269 760 278 768
rect 226 722 278 760
rect 226 716 235 722
rect 235 716 269 722
rect 269 716 278 722
rect 226 688 235 704
rect 235 688 269 704
rect 269 688 278 704
rect 226 652 278 688
rect 312 506 364 542
rect 312 490 321 506
rect 321 490 355 506
rect 355 490 364 506
rect 312 472 321 478
rect 321 472 355 478
rect 355 472 364 478
rect 312 434 364 472
rect 312 426 321 434
rect 321 426 355 434
rect 355 426 364 434
rect 312 400 321 414
rect 321 400 355 414
rect 355 400 364 414
rect 312 362 364 400
rect 312 328 321 350
rect 321 328 355 350
rect 355 328 364 350
rect 312 298 364 328
rect 312 256 321 286
rect 321 256 355 286
rect 355 256 364 286
rect 312 234 364 256
rect 312 218 364 222
rect 312 184 321 218
rect 321 184 355 218
rect 355 184 364 218
rect 312 170 364 184
rect 312 146 364 158
rect 312 112 321 146
rect 321 112 355 146
rect 355 112 364 146
rect 312 106 364 112
rect 560 1174 740 1240
rect 560 1160 591 1174
rect 591 1160 629 1174
rect 629 1160 663 1174
rect 663 1160 701 1174
rect 701 1160 735 1174
rect 735 1160 740 1174
rect 960 1174 1140 1240
rect 960 1160 985 1174
rect 985 1160 1023 1174
rect 1023 1160 1057 1174
rect 1057 1160 1095 1174
rect 1095 1160 1129 1174
rect 1129 1160 1140 1174
rect 1340 1174 1520 1240
rect 1340 1160 1345 1174
rect 1345 1160 1379 1174
rect 1379 1160 1417 1174
rect 1417 1160 1451 1174
rect 1451 1160 1489 1174
rect 1489 1160 1520 1174
rect 534 506 586 542
rect 534 490 543 506
rect 543 490 577 506
rect 577 490 586 506
rect 534 472 543 478
rect 543 472 577 478
rect 577 472 586 478
rect 534 434 586 472
rect 534 426 543 434
rect 543 426 577 434
rect 577 426 586 434
rect 534 400 543 414
rect 543 400 577 414
rect 577 400 586 414
rect 534 362 586 400
rect 534 328 543 350
rect 543 328 577 350
rect 577 328 586 350
rect 534 298 586 328
rect 534 256 543 286
rect 543 256 577 286
rect 577 256 586 286
rect 534 234 586 256
rect 534 218 586 222
rect 534 184 543 218
rect 543 184 577 218
rect 577 184 586 218
rect 534 170 586 184
rect 534 146 586 158
rect 534 112 543 146
rect 543 112 577 146
rect 577 112 586 146
rect 534 106 586 112
rect 620 1082 672 1088
rect 620 1048 629 1082
rect 629 1048 663 1082
rect 663 1048 672 1082
rect 620 1036 672 1048
rect 620 1010 672 1024
rect 620 976 629 1010
rect 629 976 663 1010
rect 663 976 672 1010
rect 620 972 672 976
rect 620 938 672 960
rect 620 908 629 938
rect 629 908 663 938
rect 663 908 672 938
rect 620 866 672 896
rect 620 844 629 866
rect 629 844 663 866
rect 663 844 672 866
rect 620 794 672 832
rect 620 780 629 794
rect 629 780 663 794
rect 663 780 672 794
rect 620 760 629 768
rect 629 760 663 768
rect 663 760 672 768
rect 620 722 672 760
rect 620 716 629 722
rect 629 716 663 722
rect 663 716 672 722
rect 620 688 629 704
rect 629 688 663 704
rect 663 688 672 704
rect 620 652 672 688
rect 706 506 758 542
rect 706 490 715 506
rect 715 490 749 506
rect 749 490 758 506
rect 706 472 715 478
rect 715 472 749 478
rect 749 472 758 478
rect 706 434 758 472
rect 706 426 715 434
rect 715 426 749 434
rect 749 426 758 434
rect 706 400 715 414
rect 715 400 749 414
rect 749 400 758 414
rect 706 362 758 400
rect 706 328 715 350
rect 715 328 749 350
rect 749 328 758 350
rect 706 298 758 328
rect 706 256 715 286
rect 715 256 749 286
rect 749 256 758 286
rect 706 234 758 256
rect 706 218 758 222
rect 706 184 715 218
rect 715 184 749 218
rect 749 184 758 218
rect 706 170 758 184
rect 706 146 758 158
rect 706 112 715 146
rect 715 112 749 146
rect 749 112 758 146
rect 706 106 758 112
rect 928 506 980 542
rect 928 490 937 506
rect 937 490 971 506
rect 971 490 980 506
rect 928 472 937 478
rect 937 472 971 478
rect 971 472 980 478
rect 928 434 980 472
rect 928 426 937 434
rect 937 426 971 434
rect 971 426 980 434
rect 928 400 937 414
rect 937 400 971 414
rect 971 400 980 414
rect 928 362 980 400
rect 928 328 937 350
rect 937 328 971 350
rect 971 328 980 350
rect 928 298 980 328
rect 928 256 937 286
rect 937 256 971 286
rect 971 256 980 286
rect 928 234 980 256
rect 928 218 980 222
rect 928 184 937 218
rect 937 184 971 218
rect 971 184 980 218
rect 928 170 980 184
rect 928 146 980 158
rect 928 112 937 146
rect 937 112 971 146
rect 971 112 980 146
rect 928 106 980 112
rect 1014 1082 1066 1088
rect 1014 1048 1023 1082
rect 1023 1048 1057 1082
rect 1057 1048 1066 1082
rect 1014 1036 1066 1048
rect 1014 1010 1066 1024
rect 1014 976 1023 1010
rect 1023 976 1057 1010
rect 1057 976 1066 1010
rect 1014 972 1066 976
rect 1014 938 1066 960
rect 1014 908 1023 938
rect 1023 908 1057 938
rect 1057 908 1066 938
rect 1014 866 1066 896
rect 1014 844 1023 866
rect 1023 844 1057 866
rect 1057 844 1066 866
rect 1014 794 1066 832
rect 1014 780 1023 794
rect 1023 780 1057 794
rect 1057 780 1066 794
rect 1014 760 1023 768
rect 1023 760 1057 768
rect 1057 760 1066 768
rect 1014 722 1066 760
rect 1014 716 1023 722
rect 1023 716 1057 722
rect 1057 716 1066 722
rect 1014 688 1023 704
rect 1023 688 1057 704
rect 1057 688 1066 704
rect 1014 652 1066 688
rect 1100 506 1152 542
rect 1100 490 1109 506
rect 1109 490 1143 506
rect 1143 490 1152 506
rect 1100 472 1109 478
rect 1109 472 1143 478
rect 1143 472 1152 478
rect 1100 434 1152 472
rect 1100 426 1109 434
rect 1109 426 1143 434
rect 1143 426 1152 434
rect 1100 400 1109 414
rect 1109 400 1143 414
rect 1143 400 1152 414
rect 1100 362 1152 400
rect 1100 328 1109 350
rect 1109 328 1143 350
rect 1143 328 1152 350
rect 1100 298 1152 328
rect 1100 256 1109 286
rect 1109 256 1143 286
rect 1143 256 1152 286
rect 1100 234 1152 256
rect 1100 218 1152 222
rect 1100 184 1109 218
rect 1109 184 1143 218
rect 1143 184 1152 218
rect 1100 170 1152 184
rect 1100 146 1152 158
rect 1100 112 1109 146
rect 1109 112 1143 146
rect 1143 112 1152 146
rect 1100 106 1152 112
rect 1322 506 1374 542
rect 1322 490 1331 506
rect 1331 490 1365 506
rect 1365 490 1374 506
rect 1322 472 1331 478
rect 1331 472 1365 478
rect 1365 472 1374 478
rect 1322 434 1374 472
rect 1322 426 1331 434
rect 1331 426 1365 434
rect 1365 426 1374 434
rect 1322 400 1331 414
rect 1331 400 1365 414
rect 1365 400 1374 414
rect 1322 362 1374 400
rect 1322 328 1331 350
rect 1331 328 1365 350
rect 1365 328 1374 350
rect 1322 298 1374 328
rect 1322 256 1331 286
rect 1331 256 1365 286
rect 1365 256 1374 286
rect 1322 234 1374 256
rect 1322 218 1374 222
rect 1322 184 1331 218
rect 1331 184 1365 218
rect 1365 184 1374 218
rect 1322 170 1374 184
rect 1322 146 1374 158
rect 1322 112 1331 146
rect 1331 112 1365 146
rect 1365 112 1374 146
rect 1322 106 1374 112
rect 1408 1082 1460 1088
rect 1408 1048 1417 1082
rect 1417 1048 1451 1082
rect 1451 1048 1460 1082
rect 1408 1036 1460 1048
rect 1408 1010 1460 1024
rect 1408 976 1417 1010
rect 1417 976 1451 1010
rect 1451 976 1460 1010
rect 1408 972 1460 976
rect 1408 938 1460 960
rect 1408 908 1417 938
rect 1417 908 1451 938
rect 1451 908 1460 938
rect 1408 866 1460 896
rect 1408 844 1417 866
rect 1417 844 1451 866
rect 1451 844 1460 866
rect 1408 794 1460 832
rect 1408 780 1417 794
rect 1417 780 1451 794
rect 1451 780 1460 794
rect 1408 760 1417 768
rect 1417 760 1451 768
rect 1451 760 1460 768
rect 1408 722 1460 760
rect 1408 716 1417 722
rect 1417 716 1451 722
rect 1451 716 1460 722
rect 1408 688 1417 704
rect 1417 688 1451 704
rect 1451 688 1460 704
rect 1408 652 1460 688
rect 1494 506 1546 542
rect 1494 490 1503 506
rect 1503 490 1537 506
rect 1537 490 1546 506
rect 1494 472 1503 478
rect 1503 472 1537 478
rect 1537 472 1546 478
rect 1494 434 1546 472
rect 1494 426 1503 434
rect 1503 426 1537 434
rect 1537 426 1546 434
rect 1494 400 1503 414
rect 1503 400 1537 414
rect 1537 400 1546 414
rect 1494 362 1546 400
rect 1494 328 1503 350
rect 1503 328 1537 350
rect 1537 328 1546 350
rect 1494 298 1546 328
rect 1494 256 1503 286
rect 1503 256 1537 286
rect 1537 256 1546 286
rect 1494 234 1546 256
rect 1494 218 1546 222
rect 1494 184 1503 218
rect 1503 184 1537 218
rect 1537 184 1546 218
rect 1494 170 1546 184
rect 1494 146 1546 158
rect 1494 112 1503 146
rect 1503 112 1537 146
rect 1537 112 1546 146
rect 1494 106 1546 112
rect 120 -180 400 -100
rect 860 -180 1580 -100
<< metal2 >>
rect 140 1240 360 1260
rect 140 1160 160 1240
rect 340 1160 360 1240
rect 140 1140 360 1160
rect 540 1240 760 1260
rect 540 1160 560 1240
rect 740 1160 760 1240
rect 540 1140 760 1160
rect 940 1240 1160 1260
rect 940 1160 960 1240
rect 1140 1160 1160 1240
rect 940 1140 1160 1160
rect 1320 1240 1540 1260
rect 1320 1160 1340 1240
rect 1520 1160 1540 1240
rect 1320 1140 1540 1160
rect 0 1088 2000 1100
rect 0 1036 226 1088
rect 278 1036 620 1088
rect 672 1036 1014 1088
rect 1066 1036 1408 1088
rect 1460 1036 2000 1088
rect 0 1024 2000 1036
rect 0 972 226 1024
rect 278 972 620 1024
rect 672 972 1014 1024
rect 1066 972 1408 1024
rect 1460 972 2000 1024
rect 0 960 2000 972
rect 0 908 226 960
rect 278 908 620 960
rect 672 908 1014 960
rect 1066 908 1408 960
rect 1460 908 2000 960
rect 0 896 2000 908
rect 0 844 226 896
rect 278 844 620 896
rect 672 844 1014 896
rect 1066 844 1408 896
rect 1460 844 2000 896
rect 0 832 2000 844
rect 0 780 226 832
rect 278 780 620 832
rect 672 780 1014 832
rect 1066 780 1408 832
rect 1460 780 2000 832
rect 0 768 2000 780
rect 0 716 226 768
rect 278 716 620 768
rect 672 716 1014 768
rect 1066 716 1408 768
rect 1460 716 2000 768
rect 0 704 2000 716
rect 0 652 226 704
rect 278 652 620 704
rect 672 652 1014 704
rect 1066 652 1408 704
rect 1460 652 2000 704
rect 0 620 2000 652
rect 120 542 380 560
rect 120 490 140 542
rect 192 490 312 542
rect 364 490 380 542
rect 120 478 380 490
rect 120 426 140 478
rect 192 426 312 478
rect 364 426 380 478
rect 120 414 380 426
rect 120 362 140 414
rect 192 362 312 414
rect 364 362 380 414
rect 120 360 380 362
rect -60 350 380 360
rect -60 320 140 350
rect -60 20 -40 320
rect 80 298 140 320
rect 192 298 312 350
rect 364 298 380 350
rect 80 286 380 298
rect 80 234 140 286
rect 192 234 312 286
rect 364 234 380 286
rect 80 222 380 234
rect 80 170 140 222
rect 192 170 312 222
rect 364 170 380 222
rect 80 158 380 170
rect 80 106 140 158
rect 192 106 312 158
rect 364 106 380 158
rect 80 20 380 106
rect -60 0 380 20
rect 520 542 780 560
rect 520 490 534 542
rect 586 490 706 542
rect 758 490 780 542
rect 520 478 780 490
rect 520 426 534 478
rect 586 426 706 478
rect 758 426 780 478
rect 520 414 780 426
rect 520 362 534 414
rect 586 362 706 414
rect 758 362 780 414
rect 520 350 780 362
rect 520 298 534 350
rect 586 298 706 350
rect 758 298 780 350
rect 520 286 780 298
rect 520 234 534 286
rect 586 234 706 286
rect 758 234 780 286
rect 520 222 780 234
rect 520 170 534 222
rect 586 170 706 222
rect 758 170 780 222
rect 520 158 780 170
rect 520 106 534 158
rect 586 106 706 158
rect 758 106 780 158
rect 100 -100 420 -80
rect 100 -180 120 -100
rect 400 -180 420 -100
rect 100 -200 420 -180
rect 240 -920 400 -200
rect 520 -220 780 106
rect 920 542 1180 560
rect 920 490 928 542
rect 980 540 1100 542
rect 1152 540 1180 542
rect 920 478 940 490
rect 920 426 928 478
rect 920 414 940 426
rect 920 362 928 414
rect 920 350 940 362
rect 920 298 928 350
rect 920 286 940 298
rect 920 234 928 286
rect 920 222 940 234
rect 920 170 928 222
rect 920 158 940 170
rect 920 106 928 158
rect 1160 120 1180 540
rect 980 106 1100 120
rect 1152 106 1180 120
rect 920 80 1180 106
rect 1300 542 1560 560
rect 1300 490 1322 542
rect 1374 490 1494 542
rect 1546 490 1560 542
rect 1300 478 1560 490
rect 1300 426 1322 478
rect 1374 426 1494 478
rect 1546 426 1560 478
rect 1300 414 1560 426
rect 1300 362 1322 414
rect 1374 362 1494 414
rect 1546 362 1560 414
rect 1300 360 1560 362
rect 1300 350 1760 360
rect 1300 298 1322 350
rect 1374 298 1494 350
rect 1546 340 1760 350
rect 1546 298 1600 340
rect 1300 286 1600 298
rect 1300 234 1322 286
rect 1374 234 1494 286
rect 1546 234 1600 286
rect 1300 222 1600 234
rect 1300 170 1322 222
rect 1374 170 1494 222
rect 1546 170 1600 222
rect 1300 158 1600 170
rect 1300 106 1322 158
rect 1374 106 1494 158
rect 1546 106 1600 158
rect 1300 20 1600 106
rect 1740 20 1760 340
rect 1300 0 1760 20
rect 840 -100 1600 -80
rect 840 -180 860 -100
rect 1580 -180 1600 -100
rect 840 -200 1600 -180
rect 520 -380 540 -220
rect 760 -380 780 -220
rect 520 -400 780 -380
rect 1160 -920 1440 -200
rect 240 -1200 1440 -920
<< via2 >>
rect -40 20 80 320
rect 940 490 980 540
rect 980 490 1100 540
rect 1100 490 1152 540
rect 1152 490 1160 540
rect 940 478 1160 490
rect 940 426 980 478
rect 980 426 1100 478
rect 1100 426 1152 478
rect 1152 426 1160 478
rect 940 414 1160 426
rect 940 362 980 414
rect 980 362 1100 414
rect 1100 362 1152 414
rect 1152 362 1160 414
rect 940 350 1160 362
rect 940 298 980 350
rect 980 298 1100 350
rect 1100 298 1152 350
rect 1152 298 1160 350
rect 940 286 1160 298
rect 940 234 980 286
rect 980 234 1100 286
rect 1100 234 1152 286
rect 1152 234 1160 286
rect 940 222 1160 234
rect 940 170 980 222
rect 980 170 1100 222
rect 1100 170 1152 222
rect 1152 170 1160 222
rect 940 158 1160 170
rect 940 120 980 158
rect 980 120 1100 158
rect 1100 120 1152 158
rect 1152 120 1160 158
rect 1600 20 1740 340
rect 540 -380 760 -220
<< metal3 >>
rect 0 1320 1680 2400
rect 900 540 1180 1320
rect -60 320 100 400
rect -60 20 -40 320
rect 80 20 100 320
rect 900 120 940 540
rect 1160 120 1180 540
rect 900 100 1180 120
rect 1580 340 1760 360
rect -60 0 100 20
rect 1580 20 1600 340
rect 1740 20 1760 340
rect 1580 0 1760 20
rect -480 -880 100 0
rect 480 -220 780 -200
rect 480 -380 540 -220
rect 760 -360 780 -220
rect 760 -380 1060 -360
rect 480 -840 1060 -380
rect 1600 -1080 2480 0
<< mimcap >>
rect 40 2340 1640 2360
rect 40 1380 60 2340
rect 1620 1380 1640 2340
rect 40 1360 1640 1380
rect -440 -60 60 -40
rect -440 -820 -420 -60
rect 40 -820 60 -60
rect 1640 -60 2440 -40
rect 520 -420 1020 -400
rect 520 -780 540 -420
rect 1000 -780 1020 -420
rect 520 -800 1020 -780
rect -440 -840 60 -820
rect 1640 -1020 1660 -60
rect 2420 -1020 2440 -60
rect 1640 -1040 2440 -1020
<< mimcapcontact >>
rect 60 1380 1620 2340
rect -420 -820 40 -60
rect 540 -780 1000 -420
rect 1660 -1020 2420 -60
<< metal4 >>
rect 0 2340 1680 2400
rect 0 1660 60 2340
rect -640 1380 60 1660
rect 1620 1380 1680 2340
rect -640 1320 1680 1380
rect -640 400 -160 1320
rect -480 180 2220 400
rect -480 0 -160 180
rect -480 -60 100 0
rect -480 -820 -420 -60
rect 40 -820 100 -60
rect 840 -360 1100 180
rect -480 -880 100 -820
rect 480 -420 1100 -360
rect 480 -780 540 -420
rect 1000 -780 1100 -420
rect 480 -840 1100 -780
rect 1600 0 2220 180
rect 1600 -60 2480 0
rect 1600 -1020 1660 -60
rect 2420 -1020 2480 -60
rect 1600 -1080 2480 -1020
<< labels >>
rlabel metal2 1880 620 2000 1100 1 BOT
rlabel metal4 -640 400 -200 1660 1 TOP
rlabel metal2 240 -1200 1440 -920 1 SUB
rlabel metal2 140 1140 360 1260 1 G2
rlabel metal2 540 1140 760 1260 1 G1
rlabel metal2 940 1140 1160 1260 1 G8
rlabel metal2 1320 1140 1540 1260 1 G4
rlabel metal3 -60 -20 100 340 1 BOT_C2
rlabel metal3 1600 0 1760 360 1 BOT_C4
rlabel metal3 900 1260 1180 1320 1 BOT_C8
rlabel metal3 520 -400 780 -220 1 BOT_C1
<< end >>
