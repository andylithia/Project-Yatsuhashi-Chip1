magic
tech sky130B
magscale 1 2
timestamp 1660185098
<< nwell >>
rect 2700 3170 4010 3300
rect 2920 3160 4010 3170
rect 2660 1550 4010 3160
rect 2660 1430 2710 1550
rect 2660 1400 3130 1430
rect 3290 1400 4010 1550
rect 2660 1340 4010 1400
rect 2660 730 4270 1340
rect 2700 0 4270 730
<< locali >>
rect 2660 3200 2750 3240
rect 2660 3120 2750 3160
rect 2650 3040 2750 3080
rect 2650 2960 2750 3000
rect 2650 2880 2750 2920
rect 2650 2800 2750 2840
rect 2650 2720 2750 2760
rect 2650 2640 2750 2680
rect 2650 2560 2750 2600
rect 2650 2480 2750 2520
rect 2650 2400 2750 2440
rect 2650 2320 2750 2360
rect 2650 2240 2750 2280
rect 2650 2160 2750 2200
rect 2650 2080 2750 2120
rect 2650 2000 2750 2040
rect 2650 1920 2750 1960
rect 2650 1840 2750 1880
rect 2650 1760 2750 1800
rect 2650 1680 2750 1720
rect 2650 1600 2750 1640
rect 2650 1550 2750 1560
rect 2650 1520 2740 1550
rect 2720 1490 2800 1510
rect 2720 1480 2740 1490
rect 2650 1450 2740 1480
rect 2780 1450 2800 1490
rect 2650 1440 2800 1450
rect 2720 1430 2800 1440
rect 2650 1360 2750 1400
rect 2650 1330 2720 1360
rect 2650 1320 3960 1330
rect 3940 1280 3960 1320
rect 2650 1260 3960 1280
rect 2660 320 4240 360
rect 2650 310 4240 320
rect 4220 260 4240 310
rect 2580 150 2590 160
rect 2650 150 2660 160
rect 2580 140 2660 150
rect 2560 60 2660 140
<< viali >>
rect 50 160 110 3220
rect 2590 1320 2650 3220
rect 2740 1450 2780 1490
rect 2590 1280 3940 1320
rect 2590 310 2650 1280
rect 2590 260 4220 310
rect 2590 150 2650 260
<< metal1 >>
rect 40 3220 120 3240
rect 2580 3220 2660 3240
rect 2580 150 2590 3220
rect 2650 1330 2660 3220
rect 3170 3120 3280 3130
rect 3170 3040 3180 3120
rect 3270 3040 3280 3120
rect 3170 3030 3280 3040
rect 3400 3110 3820 3130
rect 3400 3050 3420 3110
rect 3800 3050 3820 3110
rect 3400 3030 3820 3050
rect 3170 2800 3280 2810
rect 3170 2720 3180 2800
rect 3270 2720 3280 2800
rect 3170 2710 3280 2720
rect 3400 2790 3820 2810
rect 3400 2730 3420 2790
rect 3800 2730 3820 2790
rect 3400 2710 3820 2730
rect 3170 2480 3280 2490
rect 3170 2400 3180 2480
rect 3270 2400 3280 2480
rect 3170 2390 3280 2400
rect 3400 2470 3820 2490
rect 3400 2410 3420 2470
rect 3800 2410 3820 2470
rect 3400 2390 3820 2410
rect 3170 2170 3280 2180
rect 3170 2090 3180 2170
rect 3270 2090 3280 2170
rect 3170 2080 3280 2090
rect 3400 2150 3820 2170
rect 3400 2090 3420 2150
rect 3800 2090 3820 2150
rect 3400 2070 3820 2090
rect 3170 1850 3280 1860
rect 3170 1770 3180 1850
rect 3270 1770 3280 1850
rect 3170 1760 3280 1770
rect 3400 1830 3820 1850
rect 3400 1770 3420 1830
rect 3800 1770 3820 1830
rect 3400 1750 3820 1770
rect 3400 1520 3820 1530
rect 3280 1510 3820 1520
rect 2720 1500 2800 1510
rect 2720 1440 2730 1500
rect 2790 1440 2800 1500
rect 3280 1460 3420 1510
rect 2720 1430 2800 1440
rect 3400 1450 3420 1460
rect 3800 1450 3820 1510
rect 3400 1430 3820 1450
rect 3930 1320 3960 1330
rect 3940 1280 3960 1320
rect 3930 1260 3960 1280
rect 2650 320 2660 1260
rect 2760 1150 2840 1210
rect 3080 1150 3160 1210
rect 3390 1150 3470 1210
rect 3710 1150 3790 1210
rect 4020 1150 4100 1210
rect 2700 1100 2780 1120
rect 2700 530 2710 1100
rect 2770 530 2780 1100
rect 2700 510 2780 530
rect 2820 1100 2900 1120
rect 2820 530 2830 1100
rect 2890 530 2900 1100
rect 2820 510 2900 530
rect 3010 1100 3090 1120
rect 3010 530 3020 1100
rect 3080 530 3090 1100
rect 3010 510 3090 530
rect 3140 1100 3220 1120
rect 3140 530 3150 1100
rect 3210 530 3220 1100
rect 3140 510 3220 530
rect 3340 1100 3420 1120
rect 3340 530 3350 1100
rect 3410 530 3420 1100
rect 3340 510 3420 530
rect 3450 1100 3530 1120
rect 3450 530 3460 1100
rect 3520 530 3530 1100
rect 3450 510 3530 530
rect 3650 1100 3730 1120
rect 3650 530 3660 1100
rect 3720 530 3730 1100
rect 3650 510 3730 530
rect 3770 1100 3850 1120
rect 3770 530 3780 1100
rect 3840 530 3850 1100
rect 3770 510 3850 530
rect 3970 1100 4040 1120
rect 3970 530 3980 1100
rect 3970 510 4040 530
rect 4080 1100 4160 1120
rect 4080 530 4090 1100
rect 4150 530 4160 1100
rect 4080 510 4160 530
rect 2760 470 2840 480
rect 2760 400 2770 470
rect 2830 400 2840 470
rect 2760 390 2840 400
rect 3080 470 3160 480
rect 3080 400 3090 470
rect 3150 400 3160 470
rect 3080 390 3160 400
rect 3390 470 3470 480
rect 3390 400 3400 470
rect 3460 400 3470 470
rect 3390 390 3470 400
rect 3710 470 3790 480
rect 3710 400 3720 470
rect 3780 400 3790 470
rect 3710 390 3790 400
rect 4020 470 4100 480
rect 4020 400 4030 470
rect 4090 400 4100 470
rect 4020 390 4100 400
rect 4220 260 4250 320
rect 2650 220 4250 260
rect 2650 150 2660 220
rect 2580 140 2660 150
rect 40 40 120 120
rect 2500 60 2660 140
rect 2580 40 2660 60
<< via1 >>
rect 40 160 50 3220
rect 50 160 110 3220
rect 110 160 120 3220
rect 40 120 120 160
rect 2590 1320 2650 3220
rect 3180 3040 3270 3120
rect 3420 3050 3800 3110
rect 3180 2720 3270 2800
rect 3420 2730 3800 2790
rect 3180 2400 3270 2480
rect 3420 2410 3800 2470
rect 3180 2090 3270 2170
rect 3420 2090 3800 2150
rect 3180 1770 3270 1850
rect 3420 1770 3800 1830
rect 2730 1490 2790 1500
rect 2730 1450 2740 1490
rect 2740 1450 2780 1490
rect 2780 1450 2790 1490
rect 2730 1440 2790 1450
rect 3420 1450 3800 1510
rect 2650 1320 3930 1330
rect 2590 1280 3930 1320
rect 2590 310 2650 1280
rect 2650 1260 3930 1280
rect 2710 530 2770 1100
rect 2830 530 2890 1100
rect 3020 530 3080 1100
rect 3150 530 3210 1100
rect 3350 530 3410 1100
rect 3460 530 3520 1100
rect 3660 530 3720 1100
rect 3780 530 3840 1100
rect 3980 530 4040 1100
rect 4090 530 4150 1100
rect 2770 400 2830 470
rect 3090 400 3150 470
rect 3400 400 3460 470
rect 3720 400 3780 470
rect 4030 400 4090 470
rect 2650 310 4220 320
rect 2590 260 4220 310
rect 2590 150 2650 260
<< metal2 >>
rect 40 3220 120 3240
rect 590 3190 2100 3340
rect 2580 3220 2660 3240
rect 2580 150 2590 3220
rect 2650 1510 2660 3220
rect 3170 3120 3280 3130
rect 3170 3040 3180 3120
rect 3270 3040 3280 3120
rect 3170 3030 3280 3040
rect 3400 3110 3820 3130
rect 3400 3050 3420 3110
rect 3800 3050 3820 3110
rect 3400 3030 3820 3050
rect 3400 2810 3500 3030
rect 3170 2800 3280 2810
rect 3170 2720 3180 2800
rect 3270 2720 3280 2800
rect 3170 2710 3280 2720
rect 3400 2790 3820 2810
rect 3400 2730 3420 2790
rect 3800 2730 3820 2790
rect 3400 2710 3820 2730
rect 3400 2490 3500 2710
rect 3170 2480 3280 2490
rect 3170 2400 3180 2480
rect 3270 2400 3280 2480
rect 3170 2390 3280 2400
rect 3400 2470 3820 2490
rect 3400 2410 3420 2470
rect 3800 2410 3820 2470
rect 3400 2390 3820 2410
rect 3170 2170 3280 2180
rect 3170 2090 3180 2170
rect 3270 2090 3280 2170
rect 3170 2080 3280 2090
rect 3400 2170 3500 2390
rect 3400 2150 3820 2170
rect 3400 2090 3420 2150
rect 3800 2090 3820 2150
rect 3400 2070 3820 2090
rect 3170 1850 3280 1860
rect 3170 1770 3180 1850
rect 3270 1770 3280 1850
rect 3170 1760 3280 1770
rect 3400 1850 3500 2070
rect 3400 1830 3820 1850
rect 3400 1770 3420 1830
rect 3800 1770 3820 1830
rect 3400 1750 3820 1770
rect 3400 1670 3500 1750
rect 2920 1630 3500 1670
rect 2920 1550 2930 1630
rect 3020 1550 3500 1630
rect 2920 1540 3500 1550
rect 3400 1530 3500 1540
rect 3400 1510 3820 1530
rect 2650 1500 2800 1510
rect 2650 1440 2730 1500
rect 2790 1440 2800 1500
rect 2650 1430 2800 1440
rect 3400 1450 3420 1510
rect 3800 1450 3820 1510
rect 3400 1430 3820 1450
rect 2650 1330 2660 1430
rect 3400 1420 3500 1430
rect 3930 1260 3960 1330
rect 2650 320 2660 1260
rect 2700 1100 2780 1120
rect 2700 530 2710 1100
rect 2770 530 2780 1100
rect 2700 510 2780 530
rect 2820 1100 2900 1120
rect 2820 530 2830 1100
rect 2890 580 2900 1100
rect 3010 1100 3090 1120
rect 2890 530 2980 580
rect 2820 510 2980 530
rect 3010 530 3020 1100
rect 3080 530 3090 1100
rect 3010 510 3090 530
rect 3140 1100 3220 1120
rect 3140 530 3150 1100
rect 3210 580 3220 1100
rect 3340 1100 3420 1120
rect 3210 530 3300 580
rect 3140 510 3300 530
rect 3340 530 3350 1100
rect 3410 530 3420 1100
rect 3340 510 3420 530
rect 3450 1100 3530 1120
rect 3450 530 3460 1100
rect 3520 580 3530 1100
rect 3650 1100 3730 1120
rect 3520 530 3610 580
rect 3450 510 3610 530
rect 3650 530 3660 1100
rect 3720 530 3730 1100
rect 3650 510 3730 530
rect 3770 1100 3850 1120
rect 3770 530 3780 1100
rect 3840 580 3850 1100
rect 3970 1100 4050 1120
rect 3840 530 3930 580
rect 3770 510 3930 530
rect 3970 530 3980 1100
rect 4040 530 4050 1100
rect 3970 510 4050 530
rect 4080 1100 4160 1120
rect 4080 530 4090 1100
rect 4150 580 4160 1100
rect 4150 530 4240 580
rect 4080 510 4240 530
rect 2760 470 2840 480
rect 2760 450 2770 470
rect 2740 440 2770 450
rect 2830 450 2840 470
rect 2900 450 2980 510
rect 3080 470 3160 480
rect 3080 450 3090 470
rect 2830 440 2860 450
rect 2740 360 2750 440
rect 2850 360 2860 440
rect 2740 350 2860 360
rect 2900 320 3020 450
rect 3060 440 3090 450
rect 3150 450 3160 470
rect 3220 450 3300 510
rect 3390 470 3470 480
rect 3390 450 3400 470
rect 3150 440 3180 450
rect 3060 360 3070 440
rect 3170 360 3180 440
rect 3060 350 3180 360
rect 3220 320 3340 450
rect 3370 440 3400 450
rect 3460 450 3470 470
rect 3530 450 3610 510
rect 3710 470 3790 480
rect 3710 450 3720 470
rect 3460 440 3490 450
rect 3370 360 3380 440
rect 3480 360 3490 440
rect 3370 350 3490 360
rect 3530 320 3650 450
rect 3690 440 3720 450
rect 3780 450 3790 470
rect 3850 450 3930 510
rect 4020 470 4100 480
rect 4020 450 4030 470
rect 3780 440 3810 450
rect 3690 360 3700 440
rect 3800 360 3810 440
rect 3690 350 3810 360
rect 3850 320 3970 450
rect 4000 440 4030 450
rect 4090 450 4100 470
rect 4160 450 4240 510
rect 4090 440 4120 450
rect 4000 360 4010 440
rect 4110 360 4120 440
rect 4000 350 4120 360
rect 4160 320 4280 450
rect 4220 260 4280 320
rect 2650 220 4280 260
rect 2650 150 2660 220
rect 2580 140 2660 150
rect 40 110 120 120
rect 2500 110 2660 140
rect 2900 110 3020 220
rect 3220 110 3340 220
rect 3530 110 3650 220
rect 3850 110 3970 220
rect 4160 110 4280 220
rect 40 40 4280 110
<< via2 >>
rect 3180 3040 3270 3120
rect 3180 2720 3270 2800
rect 3180 2400 3270 2480
rect 3180 2090 3270 2170
rect 3180 1770 3270 1850
rect 2930 1550 3020 1630
rect 2730 1440 2790 1500
rect 2710 530 2770 1100
rect 3020 530 3080 1100
rect 3350 530 3410 1100
rect 3660 530 3720 1100
rect 3980 530 4040 1100
rect 2750 400 2770 440
rect 2770 400 2830 440
rect 2830 400 2850 440
rect 2750 360 2850 400
rect 3070 400 3090 440
rect 3090 400 3150 440
rect 3150 400 3170 440
rect 3070 360 3170 400
rect 3380 400 3400 440
rect 3400 400 3460 440
rect 3460 400 3480 440
rect 3380 360 3480 400
rect 3700 400 3720 440
rect 3720 400 3780 440
rect 3780 400 3800 440
rect 3700 360 3800 400
rect 4010 400 4030 440
rect 4030 400 4090 440
rect 4090 400 4110 440
rect 4010 360 4110 400
<< metal3 >>
rect 3170 3120 3280 3130
rect 3170 3040 3180 3120
rect 3270 3040 3280 3120
rect 3170 3020 3280 3040
rect 2860 2950 3280 3020
rect 2860 2780 2940 2950
rect 2710 2710 2940 2780
rect 2700 2700 2940 2710
rect 3170 2800 3280 2810
rect 3170 2720 3180 2800
rect 3270 2720 3280 2800
rect 3170 2660 3280 2720
rect 3020 2590 3280 2660
rect 3020 2560 3100 2590
rect 2760 2490 3100 2560
rect 2760 2410 2840 2490
rect 2710 2330 2840 2410
rect 3170 2480 3280 2490
rect 3170 2400 3180 2480
rect 3270 2400 3280 2480
rect 3170 2350 3280 2400
rect 3170 2340 3680 2350
rect 2900 2270 3680 2340
rect 2900 2040 2980 2270
rect 3170 2240 3680 2270
rect 3170 2170 3280 2180
rect 3170 2090 3180 2170
rect 3270 2090 3280 2170
rect 3170 2070 3280 2090
rect 2710 1960 2980 2040
rect 3040 2000 3490 2070
rect 3040 1900 3110 2000
rect 3170 1960 3490 2000
rect 2710 1830 3110 1900
rect 3170 1850 3280 1870
rect 3170 1770 3180 1850
rect 3270 1770 3280 1850
rect 2710 1700 3280 1770
rect 2710 1630 3030 1640
rect 2710 1570 2930 1630
rect 2920 1550 2930 1570
rect 3020 1550 3030 1630
rect 2920 1540 3030 1550
rect 2720 1500 2800 1510
rect 2720 1440 2730 1500
rect 2790 1440 2800 1500
rect 2720 1430 2800 1440
rect 2340 1200 3090 1350
rect 3170 1320 3280 1700
rect 3380 1530 3490 1960
rect 3570 1770 3680 2240
rect 3570 1630 3840 1770
rect 3380 1410 3630 1530
rect 3170 1200 3420 1320
rect 2340 880 2490 1200
rect 2700 1100 2780 1120
rect 2700 650 2710 1100
rect 2550 530 2710 650
rect 2770 530 2780 1100
rect 2550 510 2780 530
rect 3010 1100 3090 1200
rect 3010 530 3020 1100
rect 3080 530 3090 1100
rect 3010 510 3090 530
rect 3340 1100 3420 1200
rect 3520 1220 3630 1410
rect 3730 1410 3840 1630
rect 3730 1310 4050 1410
rect 3520 1120 3730 1220
rect 3340 530 3350 1100
rect 3410 530 3420 1100
rect 3340 510 3420 530
rect 3650 1100 3730 1120
rect 3650 530 3660 1100
rect 3720 530 3730 1100
rect 3650 510 3730 530
rect 3970 1100 4050 1310
rect 3970 530 3980 1100
rect 4040 530 4050 1100
rect 3970 510 4050 530
rect 2740 440 2860 450
rect 2740 360 2750 440
rect 2850 360 2860 440
rect 2740 350 2860 360
rect 3060 440 3180 450
rect 3060 360 3070 440
rect 3170 360 3180 440
rect 3060 350 3180 360
rect 3370 440 3490 450
rect 3370 360 3380 440
rect 3480 360 3490 440
rect 3370 350 3490 360
rect 3690 440 3810 450
rect 3690 360 3700 440
rect 3800 360 3810 440
rect 3690 350 3810 360
rect 4000 440 4120 450
rect 4000 360 4010 440
rect 4110 360 4120 440
rect 4000 350 4120 360
use pmirror_pfet_64x_flat  pmirror_pfet_64x_flat_0
timestamp 1659903400
transform 1 0 140 0 1 920
box -140 -920 2590 2420
use sky130_fd_pr__pfet_01v8_Y3CBJH  sky130_fd_pr__pfet_01v8_Y3CBJH_0
timestamp 1659909041
transform 1 0 2800 0 1 817
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_Y3CBJH  sky130_fd_pr__pfet_01v8_Y3CBJH_1
timestamp 1659909041
transform 1 0 3115 0 1 818
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_Y3CBJH  sky130_fd_pr__pfet_01v8_Y3CBJH_2
timestamp 1659909041
transform 1 0 3430 0 1 819
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_Y3CBJH  sky130_fd_pr__pfet_01v8_Y3CBJH_3
timestamp 1659909041
transform 1 0 3745 0 1 819
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_Y3CBJH  sky130_fd_pr__pfet_01v8_Y3CBJH_4
timestamp 1659909041
transform 1 0 4060 0 1 819
box -211 -519 211 519
use sky130_fd_pr__res_xhigh_po_0p35_M33Z8U  sky130_fd_pr__res_xhigh_po_0p35_M33Z8U_0
timestamp 1659907243
transform 0 1 3337 -1 0 2287
box -1057 -657 1057 657
<< labels >>
rlabel metal3 2740 350 2860 450 1 G32
rlabel metal3 3060 350 3180 450 1 G16
rlabel metal3 3370 350 3490 450 1 G2
rlabel metal3 3690 350 3810 450 1 G4
rlabel metal3 4000 350 4120 450 1 G8
rlabel metal2 40 40 4280 110 1 VHI
rlabel metal2 590 3190 2100 3340 1 IOUT
rlabel metal3 2920 1540 3030 1640 1 IREF
<< end >>
