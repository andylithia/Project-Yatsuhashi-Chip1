magic
tech sky130B
magscale 1 2
timestamp 1659907584
<< error_p >>
rect -29 2471 29 2477
rect -29 2437 -17 2471
rect -29 2431 29 2437
rect -29 1743 29 1749
rect -29 1709 -17 1743
rect -29 1703 29 1709
rect -29 1635 29 1641
rect -29 1601 -17 1635
rect -29 1595 29 1601
rect -29 907 29 913
rect -29 873 -17 907
rect -29 867 29 873
rect -29 799 29 805
rect -29 765 -17 799
rect -29 759 29 765
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect -29 -805 29 -799
rect -29 -873 29 -867
rect -29 -907 -17 -873
rect -29 -913 29 -907
rect -29 -1601 29 -1595
rect -29 -1635 -17 -1601
rect -29 -1641 29 -1635
rect -29 -1709 29 -1703
rect -29 -1743 -17 -1709
rect -29 -1749 29 -1743
rect -29 -2437 29 -2431
rect -29 -2471 -17 -2437
rect -29 -2477 29 -2471
<< nwell >>
rect -211 -2609 211 2609
<< pmos >>
rect -15 1790 15 2390
rect -15 954 15 1554
rect -15 118 15 718
rect -15 -718 15 -118
rect -15 -1554 15 -954
rect -15 -2390 15 -1790
<< pdiff >>
rect -73 2378 -15 2390
rect -73 1802 -61 2378
rect -27 1802 -15 2378
rect -73 1790 -15 1802
rect 15 2378 73 2390
rect 15 1802 27 2378
rect 61 1802 73 2378
rect 15 1790 73 1802
rect -73 1542 -15 1554
rect -73 966 -61 1542
rect -27 966 -15 1542
rect -73 954 -15 966
rect 15 1542 73 1554
rect 15 966 27 1542
rect 61 966 73 1542
rect 15 954 73 966
rect -73 706 -15 718
rect -73 130 -61 706
rect -27 130 -15 706
rect -73 118 -15 130
rect 15 706 73 718
rect 15 130 27 706
rect 61 130 73 706
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -706 -61 -130
rect -27 -706 -15 -130
rect -73 -718 -15 -706
rect 15 -130 73 -118
rect 15 -706 27 -130
rect 61 -706 73 -130
rect 15 -718 73 -706
rect -73 -966 -15 -954
rect -73 -1542 -61 -966
rect -27 -1542 -15 -966
rect -73 -1554 -15 -1542
rect 15 -966 73 -954
rect 15 -1542 27 -966
rect 61 -1542 73 -966
rect 15 -1554 73 -1542
rect -73 -1802 -15 -1790
rect -73 -2378 -61 -1802
rect -27 -2378 -15 -1802
rect -73 -2390 -15 -2378
rect 15 -1802 73 -1790
rect 15 -2378 27 -1802
rect 61 -2378 73 -1802
rect 15 -2390 73 -2378
<< pdiffc >>
rect -61 1802 -27 2378
rect 27 1802 61 2378
rect -61 966 -27 1542
rect 27 966 61 1542
rect -61 130 -27 706
rect 27 130 61 706
rect -61 -706 -27 -130
rect 27 -706 61 -130
rect -61 -1542 -27 -966
rect 27 -1542 61 -966
rect -61 -2378 -27 -1802
rect 27 -2378 61 -1802
<< nsubdiff >>
rect -175 2539 -79 2573
rect 79 2539 175 2573
rect -175 2477 -141 2539
rect 141 2477 175 2539
rect -175 -2539 -141 -2477
rect 141 -2539 175 -2477
rect -175 -2573 -79 -2539
rect 79 -2573 175 -2539
<< nsubdiffcont >>
rect -79 2539 79 2573
rect -175 -2477 -141 2477
rect 141 -2477 175 2477
rect -79 -2573 79 -2539
<< poly >>
rect -33 2471 33 2487
rect -33 2437 -17 2471
rect 17 2437 33 2471
rect -33 2421 33 2437
rect -15 2390 15 2421
rect -15 1759 15 1790
rect -33 1743 33 1759
rect -33 1709 -17 1743
rect 17 1709 33 1743
rect -33 1693 33 1709
rect -33 1635 33 1651
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -33 1585 33 1601
rect -15 1554 15 1585
rect -15 923 15 954
rect -33 907 33 923
rect -33 873 -17 907
rect 17 873 33 907
rect -33 857 33 873
rect -33 799 33 815
rect -33 765 -17 799
rect 17 765 33 799
rect -33 749 33 765
rect -15 718 15 749
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -749 15 -718
rect -33 -765 33 -749
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -815 33 -799
rect -33 -873 33 -857
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -33 -923 33 -907
rect -15 -954 15 -923
rect -15 -1585 15 -1554
rect -33 -1601 33 -1585
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -33 -1651 33 -1635
rect -33 -1709 33 -1693
rect -33 -1743 -17 -1709
rect 17 -1743 33 -1709
rect -33 -1759 33 -1743
rect -15 -1790 15 -1759
rect -15 -2421 15 -2390
rect -33 -2437 33 -2421
rect -33 -2471 -17 -2437
rect 17 -2471 33 -2437
rect -33 -2487 33 -2471
<< polycont >>
rect -17 2437 17 2471
rect -17 1709 17 1743
rect -17 1601 17 1635
rect -17 873 17 907
rect -17 765 17 799
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -799 17 -765
rect -17 -907 17 -873
rect -17 -1635 17 -1601
rect -17 -1743 17 -1709
rect -17 -2471 17 -2437
<< locali >>
rect -175 2539 -79 2573
rect 79 2539 175 2573
rect -175 2477 -141 2539
rect 141 2477 175 2539
rect -33 2437 -17 2471
rect 17 2437 33 2471
rect -61 2378 -27 2394
rect -61 1786 -27 1802
rect 27 2378 61 2394
rect 27 1786 61 1802
rect -33 1709 -17 1743
rect 17 1709 33 1743
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -61 1542 -27 1558
rect -61 950 -27 966
rect 27 1542 61 1558
rect 27 950 61 966
rect -33 873 -17 907
rect 17 873 33 907
rect -33 765 -17 799
rect 17 765 33 799
rect -61 706 -27 722
rect -61 114 -27 130
rect 27 706 61 722
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -722 -27 -706
rect 27 -130 61 -114
rect 27 -722 61 -706
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -61 -966 -27 -950
rect -61 -1558 -27 -1542
rect 27 -966 61 -950
rect 27 -1558 61 -1542
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -33 -1743 -17 -1709
rect 17 -1743 33 -1709
rect -61 -1802 -27 -1786
rect -61 -2394 -27 -2378
rect 27 -1802 61 -1786
rect 27 -2394 61 -2378
rect -33 -2471 -17 -2437
rect 17 -2471 33 -2437
rect -175 -2539 -141 -2477
rect 141 -2539 175 -2477
rect -175 -2573 -79 -2539
rect 79 -2573 175 -2539
<< viali >>
rect -17 2437 17 2471
rect -61 1802 -27 2378
rect 27 1802 61 2378
rect -17 1709 17 1743
rect -17 1601 17 1635
rect -61 966 -27 1542
rect 27 966 61 1542
rect -17 873 17 907
rect -17 765 17 799
rect -61 130 -27 706
rect 27 130 61 706
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -706 -27 -130
rect 27 -706 61 -130
rect -17 -799 17 -765
rect -17 -907 17 -873
rect -61 -1542 -27 -966
rect 27 -1542 61 -966
rect -17 -1635 17 -1601
rect -17 -1743 17 -1709
rect -61 -2378 -27 -1802
rect 27 -2378 61 -1802
rect -17 -2471 17 -2437
<< metal1 >>
rect -29 2471 29 2477
rect -29 2437 -17 2471
rect 17 2437 29 2471
rect -29 2431 29 2437
rect -67 2378 -21 2390
rect -67 1802 -61 2378
rect -27 1802 -21 2378
rect -67 1790 -21 1802
rect 21 2378 67 2390
rect 21 1802 27 2378
rect 61 1802 67 2378
rect 21 1790 67 1802
rect -29 1743 29 1749
rect -29 1709 -17 1743
rect 17 1709 29 1743
rect -29 1703 29 1709
rect -29 1635 29 1641
rect -29 1601 -17 1635
rect 17 1601 29 1635
rect -29 1595 29 1601
rect -67 1542 -21 1554
rect -67 966 -61 1542
rect -27 966 -21 1542
rect -67 954 -21 966
rect 21 1542 67 1554
rect 21 966 27 1542
rect 61 966 67 1542
rect 21 954 67 966
rect -29 907 29 913
rect -29 873 -17 907
rect 17 873 29 907
rect -29 867 29 873
rect -29 799 29 805
rect -29 765 -17 799
rect 17 765 29 799
rect -29 759 29 765
rect -67 706 -21 718
rect -67 130 -61 706
rect -27 130 -21 706
rect -67 118 -21 130
rect 21 706 67 718
rect 21 130 27 706
rect 61 130 67 706
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -706 -61 -130
rect -27 -706 -21 -130
rect -67 -718 -21 -706
rect 21 -130 67 -118
rect 21 -706 27 -130
rect 61 -706 67 -130
rect 21 -718 67 -706
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -805 29 -799
rect -29 -873 29 -867
rect -29 -907 -17 -873
rect 17 -907 29 -873
rect -29 -913 29 -907
rect -67 -966 -21 -954
rect -67 -1542 -61 -966
rect -27 -1542 -21 -966
rect -67 -1554 -21 -1542
rect 21 -966 67 -954
rect 21 -1542 27 -966
rect 61 -1542 67 -966
rect 21 -1554 67 -1542
rect -29 -1601 29 -1595
rect -29 -1635 -17 -1601
rect 17 -1635 29 -1601
rect -29 -1641 29 -1635
rect -29 -1709 29 -1703
rect -29 -1743 -17 -1709
rect 17 -1743 29 -1709
rect -29 -1749 29 -1743
rect -67 -1802 -21 -1790
rect -67 -2378 -61 -1802
rect -27 -2378 -21 -1802
rect -67 -2390 -21 -2378
rect 21 -1802 67 -1790
rect 21 -2378 27 -1802
rect 61 -2378 67 -1802
rect 21 -2390 67 -2378
rect -29 -2437 29 -2431
rect -29 -2471 -17 -2437
rect 17 -2471 29 -2437
rect -29 -2477 29 -2471
<< properties >>
string FIXED_BBOX -158 -2556 158 2556
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.15 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
