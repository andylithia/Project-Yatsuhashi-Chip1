magic
tech sky130B
magscale 1 2
timestamp 1662654558
<< pwell >>
rect 2474 100 3088 1146
<< locali >>
rect 2880 980 2960 990
rect 2880 920 2890 980
rect 2950 920 2960 980
rect 2880 910 2960 920
rect 2660 330 2740 340
rect 2660 270 2670 330
rect 2730 270 2740 330
rect 2660 260 2740 270
<< viali >>
rect 2540 1080 3080 1120
rect 2890 920 2950 980
rect 2670 270 2730 330
<< metal1 >>
rect -600 1980 2900 2000
rect -600 1910 -450 1980
rect -250 1910 50 1980
rect 250 1910 550 1980
rect 750 1910 1050 1980
rect 1250 1910 1550 1980
rect 1750 1910 2050 1980
rect 2250 1910 2550 1980
rect 2750 1910 2900 1980
rect -600 1900 2900 1910
rect -600 1880 -480 1900
rect -220 1880 20 1900
rect 280 1880 520 1900
rect 780 1880 1020 1900
rect 1280 1880 1520 1900
rect 1780 1880 2020 1900
rect 2280 1880 2520 1900
rect 2780 1880 2900 1900
rect -600 1850 -500 1880
rect -600 1650 -580 1850
rect -510 1650 -500 1850
rect -600 1620 -500 1650
rect -200 1850 0 1880
rect -200 1650 -190 1850
rect -120 1650 -80 1850
rect -10 1650 0 1850
rect -200 1620 0 1650
rect 300 1850 500 1880
rect 300 1650 310 1850
rect 380 1650 420 1850
rect 490 1650 500 1850
rect 300 1620 500 1650
rect 800 1850 1000 1880
rect 800 1650 810 1850
rect 880 1650 920 1850
rect 990 1650 1000 1850
rect 800 1620 1000 1650
rect 1300 1850 1500 1880
rect 1300 1650 1310 1850
rect 1380 1650 1420 1850
rect 1490 1650 1500 1850
rect 1300 1620 1500 1650
rect 1800 1850 2000 1880
rect 1800 1650 1810 1850
rect 1880 1650 1920 1850
rect 1990 1650 2000 1850
rect 1800 1620 2000 1650
rect 2300 1850 2500 1880
rect 2300 1650 2310 1850
rect 2380 1650 2420 1850
rect 2490 1650 2500 1850
rect 2300 1620 2500 1650
rect 2800 1850 2900 1880
rect 2800 1650 2810 1850
rect 2880 1650 2900 1850
rect 2800 1620 2900 1650
rect -600 1600 -480 1620
rect -220 1600 20 1620
rect 280 1600 520 1620
rect 780 1600 1020 1620
rect 1280 1600 1520 1620
rect 1780 1600 2020 1620
rect 2280 1600 2520 1620
rect 2780 1600 2900 1620
rect -600 1590 2900 1600
rect -600 1520 -450 1590
rect -250 1520 50 1590
rect 250 1520 550 1590
rect 750 1520 1050 1590
rect 1250 1520 1550 1590
rect 1750 1520 2050 1590
rect 2250 1520 2550 1590
rect 2750 1520 2900 1590
rect -600 1500 2900 1520
rect -100 1400 3100 1500
rect 2500 1120 3100 1400
rect 2500 1080 2540 1120
rect 3080 1080 3100 1120
rect 2500 1060 3100 1080
rect 2870 990 3000 1000
rect 2870 910 2880 990
rect 2960 910 3000 990
rect 2870 900 3000 910
rect 2650 340 2750 350
rect 2650 260 2660 340
rect 2740 260 2750 340
rect 2650 250 2750 260
<< via1 >>
rect -450 1910 -250 1980
rect 50 1910 250 1980
rect 550 1910 750 1980
rect 1050 1910 1250 1980
rect 1550 1910 1750 1980
rect 2050 1910 2250 1980
rect 2550 1910 2750 1980
rect -580 1650 -510 1850
rect -190 1650 -120 1850
rect -80 1650 -10 1850
rect 310 1650 380 1850
rect 420 1650 490 1850
rect 810 1650 880 1850
rect 920 1650 990 1850
rect 1310 1650 1380 1850
rect 1420 1650 1490 1850
rect 1810 1650 1880 1850
rect 1920 1650 1990 1850
rect 2310 1650 2380 1850
rect 2420 1650 2490 1850
rect 2810 1650 2880 1850
rect -450 1520 -250 1590
rect 50 1520 250 1590
rect 550 1520 750 1590
rect 1050 1520 1250 1590
rect 1550 1520 1750 1590
rect 2050 1520 2250 1590
rect 2550 1520 2750 1590
rect 2880 980 2960 990
rect 2880 920 2890 980
rect 2890 920 2950 980
rect 2950 920 2960 980
rect 2880 910 2960 920
rect 2660 330 2740 340
rect 2660 270 2670 330
rect 2670 270 2730 330
rect 2730 270 2740 330
rect 2660 260 2740 270
<< metal2 >>
rect -460 1980 -240 2000
rect -460 1910 -450 1980
rect -250 1910 -240 1980
rect -460 1860 -240 1910
rect 40 1980 260 2000
rect 40 1910 50 1980
rect 250 1910 260 1980
rect 40 1860 260 1910
rect 540 1980 760 2000
rect 540 1910 550 1980
rect 750 1910 760 1980
rect 540 1860 760 1910
rect 1040 1980 1260 2000
rect 1040 1910 1050 1980
rect 1250 1910 1260 1980
rect 1040 1860 1260 1910
rect 1540 1980 1760 2000
rect 1540 1910 1550 1980
rect 1750 1910 1760 1980
rect 1540 1860 1760 1910
rect 2040 1980 2260 2000
rect 2040 1910 2050 1980
rect 2250 1910 2260 1980
rect 2040 1860 2260 1910
rect 2540 1980 2760 2000
rect 2540 1910 2550 1980
rect 2750 1910 2760 1980
rect 2540 1860 2760 1910
rect -600 1850 2900 1860
rect -600 1650 -580 1850
rect -510 1650 -190 1850
rect -120 1650 -80 1850
rect -10 1650 310 1850
rect 380 1650 420 1850
rect 490 1650 810 1850
rect 880 1650 920 1850
rect 990 1650 1310 1850
rect 1380 1650 1420 1850
rect 1490 1650 1810 1850
rect 1880 1650 1920 1850
rect 1990 1650 2310 1850
rect 2380 1650 2420 1850
rect 2490 1650 2810 1850
rect 2880 1650 2900 1850
rect -600 1640 2900 1650
rect -460 1590 -240 1640
rect -460 1520 -450 1590
rect -250 1520 -240 1590
rect -460 1500 -240 1520
rect 40 1590 260 1640
rect 40 1520 50 1590
rect 250 1520 260 1590
rect 40 1500 260 1520
rect 540 1590 760 1640
rect 540 1520 550 1590
rect 750 1520 760 1590
rect 540 1500 760 1520
rect 1040 1590 1260 1640
rect 1040 1520 1050 1590
rect 1250 1520 1260 1590
rect 1040 1500 1260 1520
rect 1540 1590 1760 1640
rect 1540 1520 1550 1590
rect 1750 1520 1760 1590
rect 1540 1500 1760 1520
rect 2040 1590 2260 1640
rect 2040 1520 2050 1590
rect 2250 1520 2260 1590
rect 2040 1500 2260 1520
rect 2540 1590 2760 1640
rect 2540 1520 2550 1590
rect 2750 1520 2760 1590
rect 2540 1500 2760 1520
rect -100 1400 2600 1500
rect -100 700 100 1400
rect 2400 700 2600 1400
rect 2770 990 2970 1000
rect 2770 910 2780 990
rect 2960 910 2970 990
rect 2770 900 2970 910
rect 2650 340 2850 350
rect 2650 260 2660 340
rect 2840 260 2850 340
rect 2650 250 2850 260
<< via2 >>
rect 2780 910 2880 990
rect 2880 910 2960 990
rect 980 220 1460 500
rect 2660 260 2740 340
rect 2740 260 2840 340
<< metal3 >>
rect 2420 990 2970 1100
rect 2420 910 2780 990
rect 2960 910 2970 990
rect 2420 900 2970 910
rect -650 530 500 790
rect 2420 760 2570 900
rect 2050 540 2570 760
rect 960 500 1520 540
rect 960 220 980 500
rect 1460 220 1520 500
rect 960 180 1520 220
rect 2650 340 2850 350
rect 2650 160 2660 340
rect 2840 160 2850 340
rect 2650 150 2850 160
<< via3 >>
rect 980 220 1460 500
rect 2660 260 2840 340
rect 2660 160 2840 260
<< metal4 >>
rect 960 500 2000 551
rect 960 220 980 500
rect 1460 220 2000 500
rect 960 30 2000 220
rect 600 -80 2000 30
rect 2650 340 2850 350
rect 2650 160 2660 340
rect 2840 160 2850 340
rect 2650 -80 2850 160
rect 600 -610 3840 -80
rect 600 -800 2000 -610
use RF_nfet_6xaM02W5p0L0p15  RF_nfet_6xaM02W5p0L0p15_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1662654558
transform 1 0 0 0 1 0
box 0 0 2474 1440
use sky130_fd_pr__res_generic_po_JFYRVD  sky130_fd_pr__res_generic_po_JFYRVD_0
timestamp 1659754026
transform 1 0 2857 0 1 623
box -307 -523 307 523
<< labels >>
rlabel metal4 600 -800 2000 -10 1 NDRAIN
rlabel metal3 -650 530 -300 790 1 NGATE
rlabel space -100 1390 2610 1500 1 NSOURCE
<< end >>
