** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/OSC_HF1.sch
**.subckt OSC_HF1
XM5 nop net7 GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=3
XM1 net1 net8 GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=3
Ltfm1 vsp net3 0.1n m=1
Ltfm2 net4 vsp 0.1n m=1
V1 net2 GND 1.8
I_starter net2 net1 PULSE(0 10n 1n 10p 10p 1n 2)
R2 nop net8 1 m=1
R3 net7 net1 1 m=1
Rs1 net1 net3 0.6 m=1
K1 Ltfm1 Ltfm2 0.5
Rload nop net1 120 m=1
Rs2 nop net4 0.6 m=1
C1 nop net1 20f m=1
C2 GND net1 30f m=1
C3 GND nop 30f m=1
XM1 net5 net6 net2 net2 sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20
XM2 vbgate vbgate net2 net2 sky130_fd_pr__pfet_01v8 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
I2 vbgate GND 1m
Lbias net5 vsp 0.5n m=1
R4 net6 vbgate 1k m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice ss
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice



.subckt sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=2.828e+12p pd=2.132e+07u as=4.242e+12p
+ ps=3.198e+07u w=5.05e+06u l=150000u
X1 SOURCE SUBSTRATE SUBSTRATE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.03e+12p
+ ps=2.14e+07u w=5.05e+06u l=150000u
X2 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X5 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends
.options savecurrents
.tran 1ps 20ns
.control
run
display
plot v(nop)
plot v(nmid)
* plot @I1[i]
fft v(nop)
plot db(nop)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
