magic
tech sky130B
magscale 1 2
timestamp 1659665733
<< locali >>
rect 33 -538 3371 -528
rect 33 -572 46 -538
rect 3351 -572 3371 -538
rect 33 -597 3371 -572
<< viali >>
rect 46 -572 3351 -538
<< metal1 >>
rect 321 517 395 526
rect 321 502 330 517
rect 273 461 330 502
rect 386 502 395 517
rect 516 517 584 523
rect 516 502 522 517
rect 386 461 522 502
rect 578 502 584 517
rect 708 517 776 523
rect 708 502 714 517
rect 578 461 714 502
rect 770 502 776 517
rect 900 517 968 523
rect 900 502 906 517
rect 770 461 906 502
rect 962 502 968 517
rect 1092 517 1160 523
rect 1092 502 1098 517
rect 962 461 1098 502
rect 1154 502 1160 517
rect 1284 517 1352 523
rect 1284 502 1290 517
rect 1154 461 1290 502
rect 1346 502 1352 517
rect 1476 517 1544 523
rect 1476 502 1482 517
rect 1346 461 1482 502
rect 1538 502 1544 517
rect 1668 517 1736 523
rect 1668 502 1674 517
rect 1538 461 1674 502
rect 1730 502 1736 517
rect 1857 517 1931 526
rect 1857 502 1866 517
rect 1730 461 1866 502
rect 1922 502 1931 517
rect 2052 517 2120 523
rect 2052 502 2058 517
rect 1922 461 2058 502
rect 2114 502 2120 517
rect 2244 517 2312 523
rect 2244 502 2250 517
rect 2114 461 2250 502
rect 2306 502 2312 517
rect 2436 517 2504 523
rect 2436 502 2442 517
rect 2306 461 2442 502
rect 2498 502 2504 517
rect 2628 517 2696 523
rect 2628 502 2634 517
rect 2498 461 2634 502
rect 2690 502 2696 517
rect 2820 517 2888 523
rect 2820 502 2826 517
rect 2690 461 2826 502
rect 2882 502 2888 517
rect 3012 517 3080 523
rect 3012 502 3018 517
rect 2882 461 3018 502
rect 3074 502 3080 517
rect 3204 517 3272 523
rect 3204 502 3210 517
rect 3074 461 3210 502
rect 3266 461 3272 517
rect 273 452 3229 461
rect 282 451 340 452
rect 474 451 532 452
rect 666 451 724 452
rect 858 451 916 452
rect 1050 451 1108 452
rect 1242 451 1300 452
rect 1434 451 1492 452
rect 1626 451 1684 452
rect 1818 451 1876 452
rect 2010 451 2068 452
rect 2202 451 2260 452
rect 2394 451 2452 452
rect 2586 451 2644 452
rect 2778 451 2836 452
rect 2970 451 3028 452
rect 3162 451 3220 452
rect 135 413 199 419
rect 135 -375 141 413
rect 193 -375 199 413
rect 135 -381 199 -375
rect 231 413 295 419
rect 231 -375 237 413
rect 289 -375 295 413
rect 231 -381 295 -375
rect 327 413 391 419
rect 327 -375 333 413
rect 385 -375 391 413
rect 327 -381 391 -375
rect 423 413 487 419
rect 423 -375 429 413
rect 481 -375 487 413
rect 423 -381 487 -375
rect 519 413 583 419
rect 519 -375 525 413
rect 577 -375 583 413
rect 519 -381 583 -375
rect 615 413 679 419
rect 615 -375 621 413
rect 673 -375 679 413
rect 615 -381 679 -375
rect 711 413 775 419
rect 711 -375 717 413
rect 769 -375 775 413
rect 711 -381 775 -375
rect 807 413 871 419
rect 807 -375 813 413
rect 865 -375 871 413
rect 807 -381 871 -375
rect 903 413 967 419
rect 903 -375 909 413
rect 961 -375 967 413
rect 903 -381 967 -375
rect 999 413 1063 419
rect 999 -375 1005 413
rect 1057 -375 1063 413
rect 999 -381 1063 -375
rect 1095 413 1159 419
rect 1095 -375 1101 413
rect 1153 -375 1159 413
rect 1095 -381 1159 -375
rect 1191 413 1255 419
rect 1191 -375 1197 413
rect 1249 -375 1255 413
rect 1191 -381 1255 -375
rect 1287 413 1351 419
rect 1287 -375 1293 413
rect 1345 -375 1351 413
rect 1287 -381 1351 -375
rect 1383 413 1447 419
rect 1383 -375 1389 413
rect 1441 -375 1447 413
rect 1383 -381 1447 -375
rect 1479 413 1543 419
rect 1479 -375 1485 413
rect 1537 -375 1543 413
rect 1479 -381 1543 -375
rect 1575 413 1639 419
rect 1575 -375 1581 413
rect 1633 -375 1639 413
rect 1575 -381 1639 -375
rect 1671 413 1735 419
rect 1671 -375 1677 413
rect 1729 -375 1735 413
rect 1671 -381 1735 -375
rect 1767 413 1831 419
rect 1767 -375 1773 413
rect 1825 -375 1831 413
rect 1767 -381 1831 -375
rect 1863 413 1927 419
rect 1863 -375 1869 413
rect 1921 -375 1927 413
rect 1863 -381 1927 -375
rect 1959 412 2023 419
rect 1959 -376 1965 412
rect 2017 -376 2023 412
rect 1959 -382 2023 -376
rect 2055 413 2119 419
rect 2055 -375 2061 413
rect 2113 -375 2119 413
rect 2055 -381 2119 -375
rect 2151 413 2215 419
rect 2151 -375 2157 413
rect 2209 -375 2215 413
rect 2151 -381 2215 -375
rect 2247 413 2311 419
rect 2247 -375 2253 413
rect 2305 -375 2311 413
rect 2247 -381 2311 -375
rect 2343 413 2407 419
rect 2343 -375 2349 413
rect 2401 -375 2407 413
rect 2343 -381 2407 -375
rect 2439 413 2503 419
rect 2439 -375 2445 413
rect 2497 -375 2503 413
rect 2439 -381 2503 -375
rect 2534 413 2598 419
rect 2534 -375 2540 413
rect 2592 -375 2598 413
rect 2534 -381 2598 -375
rect 2631 412 2695 419
rect 2631 -376 2637 412
rect 2689 -376 2695 412
rect 2631 -381 2695 -376
rect 2727 413 2791 419
rect 2727 -375 2733 413
rect 2785 -375 2791 413
rect 2727 -381 2791 -375
rect 2823 413 2887 419
rect 2823 -375 2829 413
rect 2881 -375 2887 413
rect 2823 -381 2887 -375
rect 2919 413 2983 419
rect 2919 -375 2925 413
rect 2977 -375 2983 413
rect 2919 -381 2983 -375
rect 3015 413 3079 419
rect 3015 -375 3021 413
rect 3073 -375 3079 413
rect 3015 -381 3079 -375
rect 3111 413 3175 419
rect 3111 -375 3117 413
rect 3169 -375 3175 413
rect 3111 -381 3175 -375
rect 3207 413 3271 419
rect 3207 -375 3213 413
rect 3265 -375 3271 413
rect 3207 -381 3271 -375
rect 186 -418 244 -413
rect 378 -418 436 -413
rect 570 -418 628 -413
rect 762 -418 820 -413
rect 954 -418 1012 -413
rect 1146 -418 1204 -413
rect 1338 -418 1396 -413
rect 1530 -418 1588 -413
rect 2121 -418 3271 -417
rect 182 -432 3271 -418
rect 182 -478 233 -432
rect 223 -488 233 -478
rect 289 -478 433 -432
rect 289 -488 298 -478
rect 423 -488 433 -478
rect 489 -478 623 -432
rect 489 -488 498 -478
rect 613 -488 623 -478
rect 679 -478 813 -432
rect 679 -488 688 -478
rect 803 -488 813 -478
rect 869 -478 1003 -432
rect 869 -488 878 -478
rect 993 -488 1003 -478
rect 1059 -478 1193 -432
rect 1059 -488 1068 -478
rect 1183 -488 1193 -478
rect 1249 -478 1383 -432
rect 1249 -488 1258 -478
rect 1373 -488 1383 -478
rect 1439 -478 1583 -432
rect 1439 -488 1448 -478
rect 1573 -488 1583 -478
rect 1639 -433 2156 -432
rect 1639 -478 1964 -433
rect 1639 -488 1648 -478
rect 224 -497 298 -488
rect 424 -497 498 -488
rect 614 -497 688 -488
rect 804 -497 878 -488
rect 994 -497 1068 -488
rect 1184 -497 1258 -488
rect 1374 -497 1448 -488
rect 1574 -497 1648 -488
rect 1955 -489 1964 -478
rect 2020 -478 2156 -433
rect 2020 -489 2029 -478
rect 1955 -498 2029 -489
rect 2147 -488 2156 -478
rect 2212 -478 2348 -432
rect 2212 -488 2221 -478
rect 2147 -497 2221 -488
rect 2339 -488 2348 -478
rect 2404 -478 2539 -432
rect 2404 -488 2413 -478
rect 2339 -497 2413 -488
rect 2459 -488 2539 -478
rect 2595 -478 2732 -432
rect 2595 -488 2604 -478
rect 2459 -497 2604 -488
rect 2678 -488 2732 -478
rect 2788 -478 2924 -432
rect 2788 -488 2797 -478
rect 2678 -497 2797 -488
rect 2825 -488 2924 -478
rect 2980 -478 3116 -432
rect 2980 -488 2989 -478
rect 2825 -497 2989 -488
rect 3107 -488 3116 -478
rect 3172 -477 3271 -432
rect 3172 -478 3266 -477
rect 3172 -488 3181 -478
rect 3107 -497 3181 -488
rect 33 -538 3411 -528
rect 33 -540 46 -538
rect 3351 -540 3411 -538
rect 33 -592 45 -540
rect 1821 -592 1869 -572
rect 33 -598 3411 -592
<< via1 >>
rect 330 461 386 517
rect 522 461 578 517
rect 714 461 770 517
rect 906 461 962 517
rect 1098 461 1154 517
rect 1290 461 1346 517
rect 1482 461 1538 517
rect 1674 461 1730 517
rect 1866 461 1922 517
rect 2058 461 2114 517
rect 2250 461 2306 517
rect 2442 461 2498 517
rect 2634 461 2690 517
rect 2826 461 2882 517
rect 3018 461 3074 517
rect 3210 461 3266 517
rect 141 -375 193 413
rect 237 -375 289 413
rect 333 -375 385 413
rect 429 -375 481 413
rect 525 -375 577 413
rect 621 -375 673 413
rect 717 -375 769 413
rect 813 -375 865 413
rect 909 -375 961 413
rect 1005 -375 1057 413
rect 1101 -375 1153 413
rect 1197 -375 1249 413
rect 1293 -375 1345 413
rect 1389 -375 1441 413
rect 1485 -375 1537 413
rect 1581 -375 1633 413
rect 1677 -375 1729 413
rect 1773 -375 1825 413
rect 1869 -375 1921 413
rect 1965 -376 2017 412
rect 2061 -375 2113 413
rect 2157 -375 2209 413
rect 2253 -375 2305 413
rect 2349 -375 2401 413
rect 2445 -375 2497 413
rect 2540 -375 2592 413
rect 2637 -376 2689 412
rect 2733 -375 2785 413
rect 2829 -375 2881 413
rect 2925 -375 2977 413
rect 3021 -375 3073 413
rect 3117 -375 3169 413
rect 3213 -375 3265 413
rect 233 -488 289 -432
rect 433 -488 489 -432
rect 623 -488 679 -432
rect 813 -488 869 -432
rect 1003 -488 1059 -432
rect 1193 -488 1249 -432
rect 1383 -488 1439 -432
rect 1583 -488 1639 -432
rect 1964 -489 2020 -433
rect 2156 -488 2212 -432
rect 2348 -488 2404 -432
rect 2539 -488 2595 -432
rect 2732 -488 2788 -432
rect 2924 -488 2980 -432
rect 3116 -488 3172 -432
rect 45 -572 46 -540
rect 46 -572 1821 -540
rect 1869 -572 3351 -540
rect 3351 -572 3411 -540
rect 45 -592 1821 -572
rect 1869 -592 3411 -572
<< metal2 >>
rect 231 648 3173 662
rect 231 592 243 648
rect 1623 592 1779 648
rect 3159 592 3173 648
rect 231 554 3173 592
rect 231 424 293 554
rect 321 517 395 526
rect 321 461 330 517
rect 386 461 395 517
rect 321 452 395 461
rect 423 424 485 554
rect 513 517 587 526
rect 513 461 522 517
rect 578 461 587 517
rect 513 452 587 461
rect 615 424 677 554
rect 705 517 779 526
rect 705 461 714 517
rect 770 461 779 517
rect 705 452 779 461
rect 807 424 869 554
rect 897 517 971 526
rect 897 461 906 517
rect 962 461 971 517
rect 897 452 971 461
rect 999 424 1061 554
rect 1089 517 1163 526
rect 1089 461 1098 517
rect 1154 461 1163 517
rect 1089 452 1163 461
rect 1191 424 1253 554
rect 1281 517 1355 526
rect 1281 461 1290 517
rect 1346 461 1355 517
rect 1281 452 1355 461
rect 1383 424 1445 554
rect 1473 517 1547 526
rect 1473 461 1482 517
rect 1538 461 1547 517
rect 1473 452 1547 461
rect 135 413 199 419
rect 135 -375 141 413
rect 193 -375 199 413
rect 135 -381 199 -375
rect 231 413 295 424
rect 231 -375 237 413
rect 289 -375 295 413
rect 231 -381 295 -375
rect 327 413 391 419
rect 327 -375 333 413
rect 385 -375 391 413
rect 135 -528 193 -381
rect 224 -432 298 -423
rect 224 -488 233 -432
rect 289 -488 298 -432
rect 224 -497 298 -488
rect 327 -528 391 -375
rect 423 413 487 424
rect 423 -375 429 413
rect 481 -375 487 413
rect 423 -381 487 -375
rect 519 413 583 419
rect 519 -375 525 413
rect 577 -375 583 413
rect 519 -388 583 -375
rect 615 413 679 424
rect 615 -375 621 413
rect 673 -375 679 413
rect 615 -381 679 -375
rect 711 413 775 419
rect 711 -375 717 413
rect 769 -375 775 413
rect 711 -388 775 -375
rect 807 413 871 424
rect 807 -375 813 413
rect 865 -375 871 413
rect 807 -381 871 -375
rect 903 413 967 419
rect 903 -375 909 413
rect 961 -375 967 413
rect 903 -388 967 -375
rect 999 413 1063 424
rect 999 -375 1005 413
rect 1057 -375 1063 413
rect 999 -381 1063 -375
rect 1095 413 1159 419
rect 1095 -375 1101 413
rect 1153 -375 1159 413
rect 1095 -388 1159 -375
rect 1191 413 1255 424
rect 1191 -375 1197 413
rect 1249 -375 1255 413
rect 1191 -381 1255 -375
rect 1287 413 1351 419
rect 1287 -375 1293 413
rect 1345 -375 1351 413
rect 1287 -388 1351 -375
rect 1383 413 1447 424
rect 1575 419 1637 554
rect 1665 517 1739 526
rect 1665 461 1674 517
rect 1730 461 1739 517
rect 1665 452 1739 461
rect 1767 424 1829 554
rect 1857 517 1931 526
rect 1857 461 1866 517
rect 1922 461 1931 517
rect 1857 452 1931 461
rect 1959 424 2021 554
rect 2049 517 2123 526
rect 2049 461 2058 517
rect 2114 461 2123 517
rect 2049 452 2123 461
rect 2151 424 2213 554
rect 2241 517 2315 526
rect 2241 461 2250 517
rect 2306 461 2315 517
rect 2241 452 2315 461
rect 2343 424 2405 554
rect 2433 517 2507 526
rect 2433 461 2442 517
rect 2498 461 2507 517
rect 2433 452 2507 461
rect 2535 424 2597 554
rect 2625 517 2699 526
rect 2625 461 2634 517
rect 2690 461 2699 517
rect 2625 452 2699 461
rect 2727 424 2789 554
rect 2817 517 2891 526
rect 2817 461 2826 517
rect 2882 461 2891 517
rect 2817 452 2891 461
rect 2919 424 2981 554
rect 3009 517 3083 526
rect 3009 461 3018 517
rect 3074 461 3083 517
rect 3009 452 3083 461
rect 1383 -375 1389 413
rect 1441 -375 1447 413
rect 1383 -381 1447 -375
rect 1479 413 1543 419
rect 1479 -375 1485 413
rect 1537 -375 1543 413
rect 424 -432 498 -423
rect 424 -488 433 -432
rect 489 -488 498 -432
rect 424 -497 498 -488
rect 526 -528 583 -388
rect 614 -432 688 -423
rect 614 -488 623 -432
rect 679 -488 688 -432
rect 614 -497 688 -488
rect 723 -528 775 -388
rect 804 -432 878 -423
rect 804 -488 813 -432
rect 869 -488 878 -432
rect 804 -497 878 -488
rect 913 -528 963 -388
rect 994 -432 1068 -423
rect 994 -488 1003 -432
rect 1059 -488 1068 -432
rect 994 -497 1068 -488
rect 1103 -528 1153 -388
rect 1184 -432 1258 -423
rect 1184 -488 1193 -432
rect 1249 -488 1258 -432
rect 1184 -497 1258 -488
rect 1287 -528 1343 -388
rect 1374 -432 1448 -423
rect 1374 -488 1383 -432
rect 1439 -488 1448 -432
rect 1374 -497 1448 -488
rect 1479 -528 1543 -375
rect 1575 413 1639 419
rect 1575 -375 1581 413
rect 1633 -375 1639 413
rect 1575 -381 1639 -375
rect 1671 413 1735 419
rect 1671 -375 1677 413
rect 1729 -375 1735 413
rect 1671 -388 1735 -375
rect 1767 413 1831 424
rect 1767 -375 1773 413
rect 1825 -375 1831 413
rect 1767 -381 1831 -375
rect 1863 413 1927 419
rect 1863 -375 1869 413
rect 1921 -375 1927 413
rect 1574 -432 1648 -423
rect 1574 -488 1583 -432
rect 1639 -488 1648 -432
rect 1574 -497 1648 -488
rect 1683 -528 1735 -388
rect 1863 -528 1927 -375
rect 1959 412 2023 424
rect 1959 -376 1965 412
rect 2017 -376 2023 412
rect 1959 -382 2023 -376
rect 2055 413 2119 419
rect 2055 -375 2061 413
rect 2113 -375 2119 413
rect 2055 -395 2119 -375
rect 2151 413 2215 424
rect 2151 -375 2157 413
rect 2209 -375 2215 413
rect 2151 -381 2215 -375
rect 2247 413 2311 419
rect 2247 -375 2253 413
rect 2305 -375 2311 413
rect 2247 -394 2311 -375
rect 2343 413 2407 424
rect 2535 419 2598 424
rect 2343 -375 2349 413
rect 2401 -375 2407 413
rect 2343 -381 2407 -375
rect 2439 413 2503 419
rect 2439 -375 2445 413
rect 2497 -375 2503 413
rect 2439 -394 2503 -375
rect 2534 413 2598 419
rect 2534 -375 2540 413
rect 2592 -375 2598 413
rect 2534 -381 2598 -375
rect 2631 412 2695 419
rect 2631 -376 2637 412
rect 2689 -376 2695 412
rect 2631 -381 2695 -376
rect 2727 413 2791 424
rect 2727 -375 2733 413
rect 2785 -375 2791 413
rect 2727 -381 2791 -375
rect 2823 413 2887 419
rect 2823 -375 2829 413
rect 2881 -375 2887 413
rect 2631 -394 2694 -381
rect 2823 -394 2887 -375
rect 2919 413 2983 424
rect 3111 419 3173 554
rect 3201 517 3275 526
rect 3201 461 3210 517
rect 3266 461 3275 517
rect 3201 452 3275 461
rect 2919 -375 2925 413
rect 2977 -375 2983 413
rect 2919 -381 2983 -375
rect 3015 413 3079 419
rect 3015 -375 3021 413
rect 3073 -375 3079 413
rect 3015 -394 3079 -375
rect 3111 413 3175 419
rect 3111 -375 3117 413
rect 3169 -375 3175 413
rect 3111 -381 3175 -375
rect 3207 413 3271 419
rect 3207 -375 3213 413
rect 3265 -375 3271 413
rect 3207 -394 3271 -375
rect 1955 -433 2029 -423
rect 1955 -489 1964 -433
rect 2020 -489 2029 -433
rect 1955 -498 2029 -489
rect 2057 -526 2119 -395
rect 2147 -432 2221 -422
rect 2147 -488 2156 -432
rect 2212 -488 2221 -432
rect 2147 -497 2221 -488
rect 2249 -525 2311 -394
rect 2339 -432 2413 -422
rect 2339 -488 2348 -432
rect 2404 -488 2413 -432
rect 2339 -497 2413 -488
rect 2055 -528 2119 -526
rect 2247 -528 2311 -525
rect 2441 -528 2502 -394
rect 2530 -432 2604 -422
rect 2530 -488 2539 -432
rect 2595 -488 2604 -432
rect 2530 -497 2604 -488
rect 2632 -525 2694 -394
rect 2723 -432 2797 -422
rect 2723 -488 2732 -432
rect 2788 -488 2797 -432
rect 2723 -497 2797 -488
rect 2825 -525 2887 -394
rect 2915 -432 2989 -422
rect 2915 -488 2924 -432
rect 2980 -488 2989 -432
rect 2915 -497 2989 -488
rect 3017 -525 3079 -394
rect 3107 -432 3181 -422
rect 3107 -488 3116 -432
rect 3172 -488 3181 -432
rect 3107 -497 3181 -488
rect 3209 -525 3271 -394
rect 2630 -528 2694 -525
rect 2823 -528 2887 -525
rect 3015 -528 3079 -525
rect 3207 -528 3271 -525
rect 33 -540 3429 -528
rect 33 -592 45 -540
rect 1821 -592 1869 -540
rect 3411 -592 3429 -540
rect 33 -598 3429 -592
<< via2 >>
rect 243 592 1623 648
rect 1779 592 3159 648
rect 330 461 386 517
rect 522 461 578 517
rect 714 461 770 517
rect 906 461 962 517
rect 1098 461 1154 517
rect 1290 461 1346 517
rect 1482 461 1538 517
rect 233 -488 289 -432
rect 1674 461 1730 517
rect 1866 461 1922 517
rect 2058 461 2114 517
rect 2250 461 2306 517
rect 2442 461 2498 517
rect 2634 461 2690 517
rect 2826 461 2882 517
rect 3018 461 3074 517
rect 433 -488 489 -432
rect 623 -488 679 -432
rect 813 -488 869 -432
rect 1003 -488 1059 -432
rect 1193 -488 1249 -432
rect 1383 -488 1439 -432
rect 1583 -488 1639 -432
rect 3210 461 3266 517
rect 1964 -489 2020 -433
rect 2156 -488 2212 -432
rect 2348 -488 2404 -432
rect 2539 -488 2595 -432
rect 2732 -488 2788 -432
rect 2924 -488 2980 -432
rect 3116 -488 3172 -432
<< metal3 >>
rect 231 648 3173 662
rect 231 592 243 648
rect 1623 592 1779 648
rect 3159 592 3173 648
rect 231 587 3173 592
rect 321 517 3350 526
rect 321 461 330 517
rect 386 461 522 517
rect 578 461 714 517
rect 770 461 906 517
rect 962 461 1098 517
rect 1154 461 1290 517
rect 1346 461 1482 517
rect 1538 461 1674 517
rect 1730 461 1866 517
rect 1922 461 2058 517
rect 2114 461 2250 517
rect 2306 461 2442 517
rect 2498 461 2634 517
rect 2690 461 2826 517
rect 2882 461 3018 517
rect 3074 461 3210 517
rect 3266 461 3350 517
rect 321 452 3350 461
rect 1573 446 1952 452
rect 3109 446 3350 452
rect 3289 -417 3350 446
rect 2121 -418 3350 -417
rect 223 -432 3350 -418
rect 223 -488 233 -432
rect 289 -488 433 -432
rect 489 -488 623 -432
rect 679 -488 813 -432
rect 869 -488 1003 -432
rect 1059 -488 1193 -432
rect 1249 -488 1383 -432
rect 1439 -488 1583 -432
rect 1639 -433 2156 -432
rect 1639 -488 1964 -433
rect 223 -489 1964 -488
rect 2020 -488 2156 -433
rect 2212 -488 2348 -432
rect 2404 -488 2539 -432
rect 2595 -488 2732 -432
rect 2788 -488 2924 -432
rect 2980 -488 3116 -432
rect 3172 -488 3350 -432
rect 2020 -489 3350 -488
rect 223 -497 3350 -489
rect 223 -498 2151 -497
use sky130_fd_pr__pfet_01v8_8D9A6L  sky130_fd_pr__pfet_01v8_8D9A6L_0
timestamp 1659664599
transform 1 0 1703 0 1 19
box -1703 -619 1703 619
<< labels >>
rlabel metal3 231 587 3173 662 1 D
rlabel metal3 3289 -497 3350 526 1 G
rlabel metal2 33 -598 3429 -528 1 SS
<< end >>
