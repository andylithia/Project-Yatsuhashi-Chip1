magic
tech sky130B
magscale 1 2
timestamp 1660519797
<< error_p >>
rect -33246 3206 -33226 3226
rect -33266 3186 -33246 3206
rect -33286 3166 -33266 3186
rect -33306 3146 -33286 3166
rect -33326 3126 -33306 3146
rect -33346 3106 -33326 3126
rect -33366 3086 -33346 3106
rect -33386 3066 -33366 3086
rect -33406 3046 -33386 3066
rect -33426 3026 -33406 3046
rect -33446 3006 -33426 3026
rect -33466 3000 -33446 3006
rect -33446 2986 -33426 3000
rect -33466 2966 -33446 2986
rect -33486 2946 -33466 2966
rect -33506 2926 -33486 2946
rect -33526 2906 -33506 2926
rect -33546 2886 -33526 2906
rect -33566 2866 -33546 2886
rect -33586 2846 -33566 2866
rect -33606 2826 -33586 2846
rect -33626 2806 -33606 2826
rect -33646 2786 -33626 2806
rect -33666 2766 -33646 2786
rect -33686 2746 -33666 2766
rect -32794 2754 -32774 2774
rect -33706 2726 -33686 2746
rect -32814 2734 -32794 2754
rect -33726 2706 -33706 2726
rect -32834 2714 -32814 2734
rect -33746 2686 -33726 2706
rect -32854 2694 -32834 2714
rect -33766 2666 -33746 2686
rect -32874 2674 -32854 2694
rect -33786 2646 -33766 2666
rect -32894 2654 -32874 2674
rect -33806 2626 -33786 2646
rect -32914 2634 -32894 2654
rect -33826 2606 -33806 2626
rect -32934 2614 -32914 2634
rect -33846 2586 -33826 2606
rect -32954 2594 -32934 2614
rect -33866 2566 -33846 2586
rect -32974 2574 -32954 2594
rect -33886 2546 -33866 2566
rect -32994 2554 -32974 2574
rect -33906 2526 -33886 2546
rect -33014 2534 -32994 2554
rect -33926 2506 -33906 2526
rect -33034 2514 -33014 2534
rect -33946 2486 -33926 2506
rect -33054 2494 -33034 2514
rect -33966 2466 -33946 2486
rect -33074 2474 -33054 2494
rect -33986 2446 -33966 2466
rect -33094 2454 -33074 2474
rect -34006 2426 -33986 2446
rect -33114 2434 -33094 2454
rect -34026 2406 -34006 2426
rect -33134 2414 -33114 2434
rect -34046 2386 -34026 2406
rect -33154 2394 -33134 2414
rect -34066 2366 -34046 2386
rect -33174 2374 -33154 2394
rect -34086 2346 -34066 2366
rect -33194 2354 -33174 2374
rect -34106 2326 -34086 2346
rect -33214 2334 -33194 2354
rect -34126 2306 -34106 2326
rect -33234 2314 -33214 2334
rect -34146 2286 -34126 2306
rect -33254 2294 -33234 2314
rect -34166 2266 -34146 2286
rect -33274 2274 -33254 2294
rect -34186 2246 -34166 2266
rect -33294 2254 -33274 2274
rect -34206 2226 -34186 2246
rect -33314 2234 -33294 2254
rect -34226 2206 -34206 2226
rect -33334 2214 -33314 2234
rect -34246 2186 -34226 2206
rect -33354 2194 -33334 2214
rect -34266 2166 -34246 2186
rect -33374 2174 -33354 2194
rect -34286 2146 -34266 2166
rect -33394 2154 -33374 2174
rect -34306 2126 -34286 2146
rect -33414 2134 -33394 2154
rect -34326 2106 -34306 2126
rect -33434 2114 -33414 2134
rect -34346 2086 -34326 2106
rect -33454 2094 -33434 2114
rect -34365 2067 -34346 2086
rect -33474 2074 -33454 2094
rect -34384 2048 -34365 2067
rect -33494 2054 -33474 2074
rect -34403 2029 -34384 2048
rect -33514 2034 -33494 2054
rect -34421 2011 -34403 2029
rect -33534 2014 -33514 2034
rect -34439 1993 -34421 2011
rect -33554 1994 -33534 2014
rect -34457 1975 -34439 1993
rect -34475 1957 -34457 1975
rect -33574 1974 -33554 1994
rect -34492 1940 -34475 1957
rect -33594 1954 -33574 1974
rect -34509 1923 -34492 1940
rect -33614 1934 -33594 1954
rect -34526 1906 -34509 1923
rect -33634 1914 -33614 1934
rect -34543 1889 -34526 1906
rect -33654 1894 -33634 1914
rect -34559 1873 -34543 1889
rect -34575 1857 -34559 1873
rect -34139 1860 -34120 1880
rect -33674 1874 -33654 1894
rect -34591 1841 -34575 1857
rect -33694 1854 -33674 1874
rect -34607 1825 -34591 1841
rect -33714 1834 -33694 1854
rect -34622 1810 -34607 1825
rect -34637 1795 -34622 1810
rect -34195 1803 -34177 1822
rect -33734 1814 -33714 1834
rect -34652 1780 -34637 1795
rect -33754 1794 -33734 1814
rect -34667 1765 -34652 1780
rect -33774 1774 -33754 1794
rect -34681 1751 -34667 1765
rect -33794 1754 -33774 1774
rect -34695 1737 -34681 1751
rect -34709 1723 -34695 1737
rect -34266 1731 -34249 1749
rect -33814 1734 -33794 1754
rect -34722 1710 -34709 1723
rect -33834 1714 -33814 1734
rect -34735 1697 -34722 1710
rect -34748 1684 -34735 1697
rect -33854 1694 -33834 1714
rect -34761 1671 -34748 1684
rect -34773 1659 -34761 1671
rect -34333 1663 -34317 1680
rect -33874 1674 -33854 1694
rect -33894 1661 -33874 1674
rect -34785 1647 -34773 1659
rect -33908 1654 -33874 1661
rect -34797 1635 -34785 1647
rect -33908 1641 -33889 1654
rect -34809 1623 -34797 1635
rect -34820 1612 -34809 1623
rect -33932 1615 -33913 1634
rect -34831 1601 -34820 1612
rect -34842 1590 -34831 1601
rect -34396 1599 -34381 1615
rect -33951 1603 -33932 1615
rect -33963 1596 -33932 1603
rect -34853 1579 -34842 1590
rect -33963 1584 -33945 1596
rect -34863 1569 -34853 1579
rect -34873 1559 -34863 1569
rect -33987 1559 -33969 1577
rect -34883 1549 -34873 1559
rect -34892 1540 -34883 1549
rect -34901 1531 -34892 1540
rect -34455 1539 -34441 1554
rect -34005 1541 -33987 1559
rect -34910 1522 -34901 1531
rect -34023 1530 -34005 1541
rect -34034 1523 -34005 1530
rect -34919 1513 -34910 1522
rect -34927 1505 -34919 1513
rect -34034 1512 -34017 1523
rect -34935 1497 -34927 1505
rect -34496 1497 -34483 1511
rect -34943 1489 -34935 1497
rect -34951 1481 -34943 1489
rect -34057 1488 -34040 1505
rect -34958 1474 -34951 1481
rect -34965 1467 -34958 1474
rect -34074 1471 -34057 1488
rect -34972 1460 -34965 1467
rect -34091 1461 -34074 1471
rect -34978 1454 -34972 1460
rect -34984 1448 -34978 1454
rect -34990 1442 -34984 1448
rect -34547 1445 -34535 1458
rect -34100 1454 -34074 1461
rect -34100 1444 -34084 1454
rect -34996 1436 -34990 1442
rect -35001 1431 -34996 1436
rect -35006 1426 -35001 1431
rect -35011 1421 -35006 1426
rect -34123 1421 -34107 1437
rect -35015 1417 -35011 1421
rect -35019 1413 -35015 1417
rect -35023 1409 -35019 1413
rect -35027 1405 -35023 1409
rect -35030 1402 -35027 1405
rect -35033 1399 -35030 1402
rect -35036 1396 -35033 1399
rect -34594 1397 -34583 1409
rect -34139 1405 -34123 1421
rect -34155 1397 -34139 1405
rect -35038 1394 -35036 1396
rect -35040 1392 -35038 1394
rect -35042 1390 -35040 1392
rect -35043 1389 -35042 1390
rect -34163 1389 -34139 1397
rect -35044 1388 -35043 1389
rect -35045 1387 -35044 1388
rect -35046 1386 -35045 1387
rect -35047 1385 -35046 1386
rect -34163 1381 -34148 1389
rect -34637 1353 -34627 1364
rect -34185 1358 -34170 1373
rect -34200 1343 -34185 1358
rect -34215 1337 -34200 1343
rect -34666 1323 -34657 1333
rect -34222 1328 -34200 1337
rect -34222 1322 -34208 1328
rect -34243 1299 -34229 1313
rect -34701 1287 -34693 1296
rect -34257 1294 -34243 1299
rect -34262 1285 -34243 1294
rect -34262 1280 -34249 1285
rect -34732 1255 -34725 1263
rect -34283 1258 -34270 1271
rect -34296 1245 -34283 1258
rect -34309 1242 -34296 1245
rect -34752 1234 -34746 1241
rect -34312 1232 -34296 1242
rect -34312 1229 -34300 1232
rect -34775 1210 -34770 1216
rect -34333 1207 -34321 1219
rect -34789 1195 -34785 1200
rect -34345 1195 -34333 1207
rect -34357 1194 -34345 1195
rect -34359 1183 -34345 1194
rect -34804 1179 -34801 1183
rect -34359 1182 -34348 1183
rect -34812 1170 -34810 1173
rect -34817 1164 -34816 1166
rect -34379 1160 -34368 1171
rect -34821 1159 -34501 1160
rect -34401 1149 -34391 1150
rect -34390 1149 -34379 1160
rect -34401 1138 -34390 1149
rect -34421 1120 -34411 1127
rect -34429 1117 -34411 1120
rect -34431 1110 -34420 1117
rect -34431 1107 -34421 1110
rect -34449 1088 -34440 1097
rect -34458 1084 -34449 1088
rect -34462 1079 -34449 1084
rect -34467 1075 -34454 1079
rect -34467 1070 -34458 1075
rect -34483 1053 -34475 1061
rect -34492 1045 -34483 1053
rect -34499 1037 -34491 1045
rect -34510 1029 -34504 1034
rect -34513 1027 -34504 1029
rect -34531 1021 -34530 1023
rect -34513 1022 -34506 1027
rect -34520 1015 -34513 1022
rect -34530 1008 -34525 1012
rect -34532 1006 -34525 1008
rect -34532 1002 -34526 1006
rect -34538 1001 -34532 1002
rect -34540 996 -34532 1001
rect -34546 993 -34538 996
rect -34548 987 -34545 991
rect -34544 990 -34538 993
rect -34554 979 -34549 984
rect -34559 974 -34554 979
rect -34567 965 -34563 969
rect -34571 961 -34567 965
rect -34575 957 -34571 961
rect -34581 950 -34578 953
rect -34584 947 -34581 950
rect -34588 942 -34586 944
rect -34590 940 -34588 942
rect -34592 937 -34591 938
rect -34593 936 -34592 937
rect -34594 935 -34593 936
rect -34595 934 -34594 935
rect -47842 -11958 -47800 -11680
rect -48120 -12000 -47800 -11958
rect -47616 -12226 -47574 -12184
<< metal4 >>
rect -48400 -24112 -34600 -24000
rect -48400 -27888 -48288 -24112
rect -44512 -27888 -38488 -24112
rect -34712 -27888 -34600 -24112
rect -48400 -28000 -34600 -27888
<< via4 >>
rect -48288 -27888 -44512 -24112
rect -38488 -27888 -34712 -24112
<< metal5 >>
rect -57600 2980 -33020 3000
tri -33020 2980 -33000 3000 nw
tri -33000 2980 -32980 3000 se
rect -32980 2980 -11620 3000
rect -57600 2960 -33040 2980
tri -33040 2960 -33020 2980 nw
tri -33020 2960 -33000 2980 se
rect -33000 2960 -11620 2980
rect -57600 2940 -33060 2960
tri -33060 2940 -33040 2960 nw
tri -33040 2940 -33020 2960 se
rect -33020 2940 -11620 2960
rect -57600 2920 -33080 2940
tri -33080 2920 -33060 2940 nw
tri -33060 2920 -33040 2940 se
rect -33040 2920 -11620 2940
rect -57600 2900 -33100 2920
tri -33100 2900 -33080 2920 nw
tri -33080 2900 -33060 2920 se
rect -33060 2900 -11620 2920
rect -57600 2880 -33120 2900
tri -33120 2880 -33100 2900 nw
tri -33100 2880 -33080 2900 se
rect -33080 2880 -11620 2900
rect -57600 2860 -33140 2880
tri -33140 2860 -33120 2880 nw
tri -33120 2860 -33100 2880 se
rect -33100 2860 -11620 2880
rect -57600 2840 -33160 2860
tri -33160 2840 -33140 2860 nw
tri -33140 2840 -33120 2860 se
rect -33120 2840 -11620 2860
rect -57600 2820 -33180 2840
tri -33180 2820 -33160 2840 nw
tri -33160 2820 -33140 2840 se
rect -33140 2820 -11620 2840
rect -57600 2800 -33200 2820
tri -33200 2800 -33180 2820 nw
tri -33180 2800 -33160 2820 se
rect -33160 2800 -11620 2820
rect -57600 2780 -33220 2800
tri -33220 2780 -33200 2800 nw
tri -33200 2780 -33180 2800 se
rect -33180 2780 -11620 2800
rect -57600 2760 -33240 2780
tri -33240 2760 -33220 2780 nw
tri -33220 2760 -33200 2780 se
rect -33200 2760 -11620 2780
rect -57600 2740 -33260 2760
tri -33260 2740 -33240 2760 nw
tri -33240 2740 -33220 2760 se
rect -33220 2740 -11620 2760
rect -57600 2720 -33280 2740
tri -33280 2720 -33260 2740 nw
tri -33260 2720 -33240 2740 se
rect -33240 2720 -11620 2740
rect -57600 2700 -33300 2720
tri -33300 2700 -33280 2720 nw
tri -33280 2700 -33260 2720 se
rect -33260 2700 -11620 2720
rect -57600 2680 -33320 2700
tri -33320 2680 -33300 2700 nw
tri -33300 2680 -33280 2700 se
rect -33280 2680 -11620 2700
rect -57600 2660 -33340 2680
tri -33340 2660 -33320 2680 nw
tri -33320 2660 -33300 2680 se
rect -33300 2660 -11620 2680
rect -57600 2640 -33360 2660
tri -33360 2640 -33340 2660 nw
tri -33340 2640 -33320 2660 se
rect -33320 2640 -11620 2660
rect -57600 2620 -33380 2640
tri -33380 2620 -33360 2640 nw
tri -33360 2620 -33340 2640 se
rect -33340 2620 -11620 2640
rect -57600 2600 -33400 2620
tri -33400 2600 -33380 2620 nw
tri -33380 2600 -33360 2620 se
rect -33360 2600 -11620 2620
rect -57600 2580 -33420 2600
tri -33420 2580 -33400 2600 nw
tri -33400 2580 -33380 2600 se
rect -33380 2580 -11620 2600
rect -57600 2560 -33440 2580
tri -33440 2560 -33420 2580 nw
tri -33420 2560 -33400 2580 se
rect -33400 2560 -11620 2580
rect -57600 2540 -33460 2560
tri -33460 2540 -33440 2560 nw
tri -33440 2540 -33420 2560 se
rect -33420 2540 -11620 2560
rect -57600 2520 -33480 2540
tri -33480 2520 -33460 2540 nw
tri -33460 2520 -33440 2540 se
rect -33440 2520 -11620 2540
rect -57600 2500 -33500 2520
tri -33500 2500 -33480 2520 nw
tri -33480 2500 -33460 2520 se
rect -33460 2500 -11620 2520
rect -57600 2480 -33520 2500
tri -33520 2480 -33500 2500 nw
tri -33500 2480 -33480 2500 se
rect -33480 2480 -11620 2500
rect -57600 2460 -33540 2480
tri -33540 2460 -33520 2480 nw
tri -33520 2460 -33500 2480 se
rect -33500 2460 -11620 2480
rect -57600 2440 -33560 2460
tri -33560 2440 -33540 2460 nw
tri -33540 2440 -33520 2460 se
rect -33520 2440 -11620 2460
rect -57600 2420 -33580 2440
tri -33580 2420 -33560 2440 nw
tri -33560 2420 -33540 2440 se
rect -33540 2420 -11620 2440
rect -57600 2400 -33600 2420
tri -33600 2400 -33580 2420 nw
tri -33580 2400 -33560 2420 se
rect -33560 2400 -11620 2420
rect -57600 2380 -33620 2400
tri -33620 2380 -33600 2400 nw
tri -33600 2380 -33580 2400 se
rect -33580 2380 -11620 2400
rect -57600 2360 -33640 2380
tri -33640 2360 -33620 2380 nw
tri -33620 2360 -33600 2380 se
rect -33600 2360 -11620 2380
rect -57600 2340 -33660 2360
tri -33660 2340 -33640 2360 nw
tri -33640 2340 -33620 2360 se
rect -33620 2340 -11620 2360
rect -57600 2320 -33680 2340
tri -33680 2320 -33660 2340 nw
tri -33660 2320 -33640 2340 se
rect -33640 2320 -11620 2340
rect -57600 2300 -33700 2320
tri -33700 2300 -33680 2320 nw
tri -33680 2300 -33660 2320 se
rect -33660 2300 -11620 2320
rect -57600 2280 -33720 2300
tri -33720 2280 -33700 2300 nw
tri -33700 2280 -33680 2300 se
rect -33680 2280 -11620 2300
rect -57600 2260 -33740 2280
tri -33740 2260 -33720 2280 nw
tri -33720 2260 -33700 2280 se
rect -33700 2260 -11620 2280
rect -57600 2240 -33760 2260
tri -33760 2240 -33740 2260 nw
tri -33740 2240 -33720 2260 se
rect -33720 2240 -11620 2260
rect -57600 2220 -33780 2240
tri -33780 2220 -33760 2240 nw
tri -33760 2220 -33740 2240 se
rect -33740 2220 -11620 2240
rect -57600 2200 -33800 2220
tri -33800 2200 -33780 2220 nw
tri -33780 2200 -33760 2220 se
rect -33760 2200 -11620 2220
rect -57600 2180 -33820 2200
tri -33820 2180 -33800 2200 nw
tri -33800 2180 -33780 2200 se
rect -33780 2180 -11620 2200
rect -57600 2160 -33840 2180
tri -33840 2160 -33820 2180 nw
tri -33820 2160 -33800 2180 se
rect -33800 2160 -11620 2180
rect -57600 2140 -33860 2160
tri -33860 2140 -33840 2160 nw
tri -33840 2140 -33820 2160 se
rect -33820 2140 -11620 2160
rect -57600 2120 -33880 2140
tri -33880 2120 -33860 2140 nw
tri -33860 2120 -33840 2140 se
rect -33840 2120 -11620 2140
rect -57600 2100 -33900 2120
tri -33900 2100 -33880 2120 nw
tri -33880 2100 -33860 2120 se
rect -33860 2100 -11620 2120
rect -57600 2080 -33920 2100
tri -33920 2080 -33900 2100 nw
tri -33900 2080 -33880 2100 se
rect -33880 2080 -11620 2100
rect -57600 2060 -33940 2080
tri -33940 2060 -33920 2080 nw
tri -33920 2060 -33900 2080 se
rect -33900 2060 -11620 2080
rect -57600 2040 -33960 2060
tri -33960 2040 -33940 2060 nw
tri -33940 2040 -33920 2060 se
rect -33920 2040 -11620 2060
rect -57600 2020 -33980 2040
tri -33980 2020 -33960 2040 nw
tri -33960 2020 -33940 2040 se
rect -33940 2020 -11620 2040
rect -57600 2000 -34000 2020
tri -34000 2000 -33980 2020 nw
tri -33980 2000 -33960 2020 se
rect -33960 2000 -11620 2020
rect -57600 1980 -34020 2000
tri -34020 1980 -34000 2000 nw
tri -34000 1980 -33980 2000 se
rect -33980 1980 -11620 2000
rect -57600 1960 -34040 1980
tri -34040 1960 -34020 1980 nw
tri -34020 1960 -34000 1980 se
rect -34000 1960 -11620 1980
rect -57600 1940 -34060 1960
tri -34060 1940 -34040 1960 nw
tri -34040 1940 -34020 1960 se
rect -34020 1940 -11620 1960
rect -57600 1920 -34080 1940
tri -34080 1920 -34060 1940 nw
tri -34060 1920 -34040 1940 se
rect -34040 1920 -11620 1940
rect -57600 1900 -34100 1920
tri -34100 1900 -34080 1920 nw
tri -34080 1900 -34060 1920 se
rect -34060 1900 -11620 1920
rect -57600 1880 -34120 1900
tri -34120 1880 -34100 1900 nw
tri -34100 1880 -34080 1900 se
rect -34080 1880 -11620 1900
rect -57600 1860 -34139 1880
tri -34139 1860 -34120 1880 nw
tri -34120 1860 -34100 1880 se
rect -34100 1860 -11620 1880
rect -57600 1841 -34158 1860
tri -34158 1841 -34139 1860 nw
tri -34139 1841 -34120 1860 se
rect -34120 1841 -11620 1860
rect -57600 1822 -34177 1841
tri -34177 1822 -34158 1841 nw
tri -34158 1822 -34139 1841 se
rect -34139 1822 -11620 1841
rect -57600 1803 -34195 1822
tri -34195 1803 -34177 1822 nw
tri -34177 1803 -34158 1822 se
rect -34158 1803 -11620 1822
rect -57600 1785 -34213 1803
tri -34213 1785 -34195 1803 nw
tri -34195 1785 -34177 1803 se
rect -34177 1785 -11620 1803
rect -57600 1767 -34231 1785
tri -34231 1767 -34213 1785 nw
tri -34213 1767 -34195 1785 se
rect -34195 1767 -11620 1785
rect -57600 1749 -34249 1767
tri -34249 1749 -34231 1767 nw
tri -34231 1749 -34213 1767 se
rect -34213 1749 -11620 1767
rect -57600 1731 -34266 1749
tri -34266 1731 -34249 1749 nw
tri -34249 1731 -34231 1749 se
rect -34231 1731 -11620 1749
rect -57600 1714 -34283 1731
tri -34283 1714 -34266 1731 nw
tri -34266 1714 -34249 1731 se
rect -34249 1714 -11620 1731
rect -57600 1697 -34300 1714
tri -34300 1697 -34283 1714 nw
tri -34283 1697 -34266 1714 se
rect -34266 1697 -11620 1714
rect -57600 1680 -34317 1697
tri -34317 1680 -34300 1697 nw
tri -34300 1680 -34283 1697 se
rect -34283 1680 -11620 1697
rect -57600 1663 -34333 1680
tri -34333 1663 -34317 1680 nw
tri -34317 1663 -34300 1680 se
rect -34300 1663 -11620 1680
rect -57600 1647 -34349 1663
tri -34349 1647 -34333 1663 nw
tri -34333 1647 -34317 1663 se
rect -34317 1647 -11620 1663
rect -57600 1631 -34365 1647
tri -34365 1631 -34349 1647 nw
tri -34349 1631 -34333 1647 se
rect -34333 1631 -11620 1647
rect -57600 1615 -34381 1631
tri -34381 1615 -34365 1631 nw
tri -34365 1615 -34349 1631 se
rect -34349 1615 -11620 1631
rect -57600 1599 -34396 1615
tri -34396 1599 -34381 1615 nw
tri -34381 1599 -34365 1615 se
rect -34365 1599 -11620 1615
rect -57600 1584 -34411 1599
tri -34411 1584 -34396 1599 nw
tri -34396 1584 -34381 1599 se
rect -34381 1584 -11620 1599
rect -57600 1569 -34426 1584
tri -34426 1569 -34411 1584 nw
tri -34411 1569 -34396 1584 se
rect -34396 1569 -11620 1584
rect -57600 1554 -34441 1569
tri -34441 1554 -34426 1569 nw
tri -34426 1554 -34411 1569 se
rect -34411 1554 -11620 1569
rect -57600 1539 -34455 1554
tri -34455 1539 -34441 1554 nw
tri -34441 1539 -34426 1554 se
rect -34426 1539 -11620 1554
rect -57600 1525 -34469 1539
tri -34469 1525 -34455 1539 nw
tri -34455 1525 -34441 1539 se
rect -34441 1525 -11620 1539
rect -57600 1511 -34483 1525
tri -34483 1511 -34469 1525 nw
tri -34469 1511 -34455 1525 se
rect -34455 1511 -11620 1525
rect -57600 1497 -34496 1511
tri -34496 1497 -34483 1511 nw
tri -34483 1497 -34469 1511 se
rect -34469 1497 -11620 1511
rect -57600 1484 -34509 1497
tri -34509 1484 -34496 1497 nw
tri -34496 1484 -34483 1497 se
rect -34483 1484 -11620 1497
rect -57600 1471 -34522 1484
tri -34522 1471 -34509 1484 nw
tri -34509 1471 -34496 1484 se
rect -34496 1471 -11620 1484
rect -57600 1458 -34535 1471
tri -34535 1458 -34522 1471 nw
tri -34522 1458 -34509 1471 se
rect -34509 1458 -11620 1471
rect -57600 1445 -34547 1458
tri -34547 1445 -34535 1458 nw
tri -34535 1445 -34522 1458 se
rect -34522 1445 -11620 1458
rect -57600 1433 -34559 1445
tri -34559 1433 -34547 1445 nw
tri -34547 1433 -34535 1445 se
rect -34535 1433 -11620 1445
rect -57600 1421 -34571 1433
tri -34571 1421 -34559 1433 nw
tri -34559 1421 -34547 1433 se
rect -34547 1421 -11620 1433
rect -57600 1409 -34583 1421
tri -34583 1409 -34571 1421 nw
tri -34571 1409 -34559 1421 se
rect -34559 1409 -11620 1421
rect -57600 1397 -34594 1409
tri -34594 1397 -34583 1409 nw
tri -34583 1397 -34571 1409 se
rect -34571 1397 -11620 1409
rect -57600 1386 -34605 1397
tri -34605 1386 -34594 1397 nw
tri -34594 1386 -34583 1397 se
rect -34583 1386 -11620 1397
rect -57600 1375 -34616 1386
tri -34616 1375 -34605 1386 nw
tri -34605 1375 -34594 1386 se
rect -34594 1375 -11620 1386
rect -57600 1364 -34627 1375
tri -34627 1364 -34616 1375 nw
tri -34616 1364 -34605 1375 se
rect -34605 1364 -11620 1375
rect -57600 1353 -34637 1364
tri -34637 1353 -34627 1364 nw
tri -34627 1353 -34616 1364 se
rect -34616 1353 -11620 1364
rect -57600 1343 -34647 1353
tri -34647 1343 -34637 1353 nw
tri -34637 1343 -34627 1353 se
rect -34627 1343 -11620 1353
rect -57600 1333 -34657 1343
tri -34657 1333 -34647 1343 nw
tri -34647 1333 -34637 1343 se
rect -34637 1333 -11620 1343
rect -57600 1323 -34666 1333
tri -34666 1323 -34657 1333 nw
tri -34657 1323 -34647 1333 se
rect -34647 1323 -11620 1333
rect -57600 1314 -34675 1323
tri -34675 1314 -34666 1323 nw
tri -34666 1314 -34657 1323 se
rect -34657 1314 -11620 1323
rect -57600 1305 -34684 1314
tri -34684 1305 -34675 1314 nw
tri -34675 1305 -34666 1314 se
rect -34666 1305 -11620 1314
rect -57600 1296 -34693 1305
tri -34693 1296 -34684 1305 nw
tri -34684 1296 -34675 1305 se
rect -34675 1296 -11620 1305
rect -57600 1287 -34701 1296
tri -34701 1287 -34693 1296 nw
tri -34693 1287 -34684 1296 se
rect -34684 1287 -11620 1296
rect -57600 1279 -34709 1287
tri -34709 1279 -34701 1287 nw
tri -34701 1279 -34693 1287 se
rect -34693 1279 -11620 1287
rect -57600 1271 -34717 1279
tri -34717 1271 -34709 1279 nw
tri -34709 1271 -34701 1279 se
rect -34701 1271 -11620 1279
rect -57600 1263 -34725 1271
tri -34725 1263 -34717 1271 nw
tri -34717 1263 -34709 1271 se
rect -34709 1263 -11620 1271
rect -57600 1255 -34732 1263
tri -34732 1255 -34725 1263 nw
tri -34725 1255 -34717 1263 se
rect -34717 1255 -11620 1263
rect -57600 1248 -34739 1255
tri -34739 1248 -34732 1255 nw
tri -34732 1248 -34725 1255 se
rect -34725 1248 -11620 1255
rect -57600 1241 -34746 1248
tri -34746 1241 -34739 1248 nw
tri -34739 1241 -34732 1248 se
rect -34732 1241 -11620 1248
rect -57600 1234 -34752 1241
tri -34752 1234 -34746 1241 nw
tri -34746 1234 -34739 1241 se
rect -34739 1234 -11620 1241
rect -57600 1228 -34758 1234
tri -34758 1228 -34752 1234 nw
tri -34752 1228 -34746 1234 se
rect -34746 1228 -11620 1234
rect -57600 1222 -34764 1228
tri -34764 1222 -34758 1228 nw
tri -34758 1222 -34752 1228 se
rect -34752 1222 -11620 1228
rect -57600 1216 -34770 1222
tri -34770 1216 -34764 1222 nw
tri -34764 1216 -34758 1222 se
rect -34758 1216 -11620 1222
rect -57600 1210 -34775 1216
tri -34775 1210 -34770 1216 nw
tri -34770 1210 -34764 1216 se
rect -34764 1210 -11620 1216
rect -57600 1205 -34780 1210
tri -34780 1205 -34775 1210 nw
tri -34775 1205 -34770 1210 se
rect -34770 1205 -11620 1210
rect -57600 1200 -34785 1205
tri -34785 1200 -34780 1205 nw
tri -34780 1200 -34775 1205 se
rect -34775 1200 -11620 1205
rect -57600 1195 -34789 1200
tri -34789 1195 -34785 1200 nw
tri -34785 1195 -34780 1200 se
rect -34780 1195 -11620 1200
rect -57600 1191 -34793 1195
tri -34793 1191 -34789 1195 nw
tri -34789 1191 -34785 1195 se
rect -34785 1191 -11620 1195
rect -57600 1187 -34797 1191
tri -34797 1187 -34793 1191 nw
tri -34793 1187 -34789 1191 se
rect -34789 1187 -11620 1191
rect -57600 1183 -34801 1187
tri -34801 1183 -34797 1187 nw
tri -34797 1183 -34793 1187 se
rect -34793 1183 -11620 1187
rect -57600 1179 -34804 1183
tri -34804 1179 -34801 1183 nw
tri -34801 1179 -34797 1183 se
rect -34797 1179 -11620 1183
rect -57600 1176 -34807 1179
tri -34807 1176 -34804 1179 nw
tri -34804 1176 -34801 1179 se
rect -34801 1176 -11620 1179
rect -57600 1173 -34810 1176
tri -34810 1173 -34807 1176 nw
tri -34807 1173 -34804 1176 se
rect -34804 1173 -11620 1176
rect -57600 1170 -34812 1173
tri -34812 1170 -34810 1173 nw
tri -34810 1170 -34807 1173 se
rect -34807 1170 -11620 1173
rect -57600 1168 -34814 1170
tri -34814 1168 -34812 1170 nw
tri -34812 1168 -34810 1170 se
rect -34810 1168 -11620 1170
rect -57600 1166 -34816 1168
tri -34816 1166 -34814 1168 nw
tri -34814 1166 -34812 1168 se
rect -34812 1166 -11620 1168
rect -57600 1164 -34817 1166
tri -34817 1164 -34816 1166 nw
tri -34816 1164 -34814 1166 se
rect -34814 1164 -11620 1166
rect -57600 1163 -34818 1164
tri -34818 1163 -34817 1164 nw
tri -34817 1163 -34816 1164 se
rect -34816 1163 -11620 1164
rect -57600 1162 -34819 1163
tri -34819 1162 -34818 1163 nw
tri -34818 1162 -34817 1163 se
rect -34817 1162 -11620 1163
rect -57600 1161 -34820 1162
tri -34820 1161 -34819 1162 nw
tri -34819 1161 -34818 1162 se
rect -34818 1161 -11620 1162
rect -57600 1159 -34821 1161
tri -34821 1160 -34820 1161 nw
tri -34820 1160 -34819 1161 se
rect -34819 1160 -11620 1161
tri -34821 1159 -34820 1160 se
rect -34820 1159 -11620 1160
rect -57600 906 -11620 1159
tri -11620 906 -9526 3000 sw
rect -57600 904 -9526 906
tri -9526 904 -9524 906 sw
rect -57600 -1000 -9524 904
tri -9524 -1000 -7620 904 sw
rect -57600 -1600 -31923 -1000
tri -31923 -1600 -31323 -1000 nw
tri -13277 -1600 -12677 -1000 ne
rect -12677 -1600 -7620 -1000
rect -57600 -2449 -32772 -1600
tri -32772 -2449 -31923 -1600 nw
tri -31923 -2449 -31074 -1600 se
rect -31074 -2449 -13526 -1600
tri -13526 -2449 -12677 -1600 sw
tri -12677 -2449 -11828 -1600 ne
rect -11828 -2449 -7620 -1600
rect -57600 -3298 -33621 -2449
tri -33621 -3298 -32772 -2449 nw
tri -32772 -3298 -31923 -2449 se
rect -31923 -3298 -12677 -2449
tri -12677 -3298 -11828 -2449 sw
tri -11828 -3298 -10979 -2449 ne
rect -10979 -3298 -7620 -2449
rect -57600 -3902 -34225 -3298
tri -34225 -3902 -33621 -3298 nw
tri -33376 -3902 -32772 -3298 se
rect -32772 -3902 -11828 -3298
tri -11828 -3902 -11224 -3298 sw
tri -10979 -3902 -10375 -3298 ne
rect -10375 -3902 -7620 -3298
rect -57600 -4751 -35074 -3902
tri -35074 -4751 -34225 -3902 nw
tri -34225 -4751 -33376 -3902 se
rect -33376 -4751 -11224 -3902
tri -11224 -4751 -10375 -3902 sw
tri -10375 -4751 -9526 -3902 ne
rect -9526 -4751 -7620 -3902
rect -57600 -5600 -35923 -4751
tri -35923 -5600 -35074 -4751 nw
tri -35074 -5600 -34225 -4751 se
rect -34225 -5600 -10375 -4751
tri -10375 -5600 -9526 -4751 sw
tri -9526 -5600 -8677 -4751 ne
rect -8677 -5600 -7620 -4751
tri -7620 -5600 -3020 -1000 sw
rect -57600 -6449 -36772 -5600
tri -36772 -6449 -35923 -5600 nw
tri -35923 -6449 -35074 -5600 se
rect -35074 -6449 -33543 -5600
rect -57600 -7298 -37621 -6449
tri -37621 -7298 -36772 -6449 nw
tri -36772 -7298 -35923 -6449 se
rect -35923 -7298 -33543 -6449
rect -57600 -8028 -38351 -7298
tri -38351 -8028 -37621 -7298 nw
tri -37502 -8028 -36772 -7298 se
rect -36772 -8028 -33543 -7298
rect -57600 -8877 -39200 -8028
tri -39200 -8877 -38351 -8028 nw
tri -38351 -8877 -37502 -8028 se
rect -37502 -8877 -33543 -8028
rect -57600 -9726 -40049 -8877
tri -40049 -9726 -39200 -8877 nw
tri -39200 -9726 -38351 -8877 se
rect -38351 -9726 -33543 -8877
tri -33543 -9726 -29417 -5600 nw
tri -15183 -9726 -11057 -5600 ne
rect -11057 -6449 -9526 -5600
tri -9526 -6449 -8677 -5600 sw
tri -8677 -6449 -7828 -5600 ne
rect -7828 -6449 -3020 -5600
rect -11057 -7298 -8677 -6449
tri -8677 -7298 -7828 -6449 sw
tri -7828 -7298 -6979 -6449 ne
rect -6979 -7298 -3020 -6449
rect -11057 -8028 -7828 -7298
tri -7828 -8028 -7098 -7298 sw
tri -6979 -8028 -6249 -7298 ne
rect -6249 -8028 -3020 -7298
rect -11057 -8877 -7098 -8028
tri -7098 -8877 -6249 -8028 sw
tri -6249 -8877 -5400 -8028 ne
rect -5400 -8877 -3020 -8028
rect -11057 -9726 -6249 -8877
tri -6249 -9726 -5400 -8877 sw
tri -5400 -9726 -4551 -8877 ne
rect -4551 -9726 -3020 -8877
tri -3020 -9726 1106 -5600 sw
rect -57600 -10575 -40898 -9726
tri -40898 -10575 -40049 -9726 nw
tri -40049 -10575 -39200 -9726 se
rect -39200 -10575 -35074 -9726
rect -57600 -11257 -41580 -10575
tri -41580 -11257 -40898 -10575 nw
tri -40731 -11257 -40049 -10575 se
rect -40049 -11257 -35074 -10575
tri -35074 -11257 -33543 -9726 nw
tri -11057 -11257 -9526 -9726 ne
rect -9526 -10575 -5400 -9726
tri -5400 -10575 -4551 -9726 sw
tri -4551 -10575 -3702 -9726 ne
rect -3702 -10575 1106 -9726
rect -9526 -11257 -4551 -10575
rect -57600 -11958 -42323 -11257
rect -57600 -12000 -47842 -11958
tri -47842 -12000 -47800 -11958 nw
rect -47800 -12000 -42323 -11958
tri -42323 -12000 -41580 -11257 nw
tri -41474 -12000 -40731 -11257 se
rect -40731 -12000 -35817 -11257
tri -35817 -12000 -35074 -11257 nw
tri -9526 -12000 -8783 -11257 ne
rect -8783 -11424 -4551 -11257
tri -4551 -11424 -3702 -10575 sw
tri -3702 -11424 -2853 -10575 ne
rect -2853 -11424 1106 -10575
rect -8783 -12000 -3702 -11424
rect -57600 -12849 -43172 -12000
tri -43172 -12849 -42323 -12000 nw
tri -42323 -12849 -41474 -12000 se
rect -41474 -12849 -39200 -12000
rect -57600 -12877 -43200 -12849
tri -43200 -12877 -43172 -12849 nw
tri -42351 -12877 -42323 -12849 se
rect -42323 -12877 -39200 -12849
rect -57600 -16000 -43800 -12877
tri -43800 -13477 -43200 -12877 nw
tri -42951 -13477 -42351 -12877 se
rect -42351 -13477 -39200 -12877
tri -43200 -13726 -42951 -13477 se
rect -42951 -13726 -39200 -13477
rect -57600 -24112 -44400 -24000
rect -57600 -27888 -48288 -24112
rect -44512 -27888 -44400 -24112
rect -57600 -28000 -44400 -27888
rect -43200 -28000 -39200 -13726
tri -39200 -15383 -35817 -12000 nw
tri -8783 -15383 -5400 -12000 ne
rect -5400 -12028 -3702 -12000
tri -3702 -12028 -3098 -11424 sw
tri -2853 -12028 -2249 -11424 ne
rect -2249 -11820 1106 -11424
tri 1106 -11820 3200 -9726 sw
rect -2249 -12028 3200 -11820
rect -5400 -12877 -3098 -12028
tri -3098 -12877 -2249 -12028 sw
tri -2249 -12877 -1400 -12028 ne
rect -1400 -12877 3200 -12028
rect -5400 -13477 -2249 -12877
tri -2249 -13477 -1649 -12877 sw
tri -1400 -13477 -800 -12877 ne
rect -5400 -13726 -1649 -13477
tri -1649 -13726 -1400 -13477 sw
rect -38600 -24112 -34600 -24000
tri -39200 -28000 -39070 -27870 sw
rect -38600 -27888 -38488 -24112
rect -34712 -27888 -34600 -24112
rect -38600 -28000 -34600 -27888
tri -34600 -28000 -32565 -25965 sw
tri -7435 -28000 -5400 -25965 se
rect -5400 -27622 -1400 -13726
rect -5400 -27870 -1648 -27622
tri -1648 -27870 -1400 -27622 nw
rect -5400 -28000 -2248 -27870
rect -43200 -28470 -39070 -28000
tri -39070 -28470 -38600 -28000 sw
tri -38222 -28470 -37752 -28000 ne
rect -37752 -28470 -32565 -28000
rect -43200 -29318 -38600 -28470
tri -38600 -29318 -37752 -28470 sw
tri -37752 -29318 -36904 -28470 ne
rect -36904 -29318 -32565 -28470
rect -43200 -29527 -37752 -29318
tri -43200 -31622 -41105 -29527 ne
rect -41105 -29926 -37752 -29527
tri -37752 -29926 -37144 -29318 sw
tri -36904 -29926 -36296 -29318 ne
rect -36296 -29926 -32565 -29318
rect -41105 -30774 -37144 -29926
tri -37144 -30774 -36296 -29926 sw
tri -36296 -30774 -35448 -29926 ne
rect -35448 -30774 -32565 -29926
rect -41105 -31622 -36296 -30774
tri -36296 -31622 -35448 -30774 sw
tri -35448 -31622 -34600 -30774 ne
rect -34600 -31622 -32565 -30774
tri -32565 -31622 -28943 -28000 sw
tri -8178 -28743 -7435 -28000 se
rect -7435 -28470 -2248 -28000
tri -2248 -28470 -1648 -27870 nw
tri -1400 -28470 -800 -27870 se
rect -800 -28470 3200 -12877
rect -7435 -28743 -2521 -28470
tri -2521 -28743 -2248 -28470 nw
tri -1673 -28743 -1400 -28470 se
rect -1400 -28743 3200 -28470
tri -11057 -31622 -8178 -28743 se
rect -8178 -29591 -3369 -28743
tri -3369 -29591 -2521 -28743 nw
tri -2521 -29591 -1673 -28743 se
rect -1673 -29527 3200 -28743
rect -1673 -29591 257 -29527
rect -8178 -29926 -3704 -29591
tri -3704 -29926 -3369 -29591 nw
tri -2856 -29926 -2521 -29591 se
rect -2521 -29926 257 -29591
rect -8178 -30774 -4552 -29926
tri -4552 -30774 -3704 -29926 nw
tri -3704 -30774 -2856 -29926 se
rect -2856 -30774 257 -29926
rect -8178 -31622 -5400 -30774
tri -5400 -31622 -4552 -30774 nw
tri -4552 -31622 -3704 -30774 se
rect -3704 -31622 257 -30774
tri -41105 -34400 -38327 -31622 ne
rect -38327 -32470 -35448 -31622
tri -35448 -32470 -34600 -31622 sw
tri -34600 -32470 -33752 -31622 ne
rect -33752 -32470 -28943 -31622
rect -38327 -33318 -34600 -32470
tri -34600 -33318 -33752 -32470 sw
tri -33752 -33318 -32904 -32470 ne
rect -32904 -33318 -28943 -32470
rect -38327 -33552 -33752 -33318
tri -33752 -33552 -33518 -33318 sw
tri -32904 -33552 -32670 -33318 ne
rect -32670 -33552 -28943 -33318
rect -38327 -34400 -33518 -33552
tri -33518 -34400 -32670 -33552 sw
tri -32670 -34400 -31822 -33552 ne
rect -31822 -34400 -28943 -33552
tri -28943 -34400 -26165 -31622 sw
tri -13835 -34400 -11057 -31622 se
rect -11057 -32470 -6248 -31622
tri -6248 -32470 -5400 -31622 nw
tri -5400 -32470 -4552 -31622 se
rect -4552 -32470 257 -31622
tri 257 -32470 3200 -29527 nw
rect -11057 -33318 -7096 -32470
tri -7096 -33318 -6248 -32470 nw
tri -6248 -33318 -5400 -32470 se
rect -5400 -33318 -800 -32470
rect -11057 -33552 -7330 -33318
tri -7330 -33552 -7096 -33318 nw
tri -6482 -33552 -6248 -33318 se
rect -6248 -33527 -800 -33318
tri -800 -33527 257 -32470 nw
rect -6248 -33552 -2521 -33527
rect -11057 -34400 -8178 -33552
tri -8178 -34400 -7330 -33552 nw
tri -7330 -34400 -6482 -33552 se
rect -6482 -34400 -2521 -33552
tri -38327 -39000 -33727 -34400 ne
rect -33727 -35248 -32670 -34400
tri -32670 -35248 -31822 -34400 sw
tri -31822 -35248 -30974 -34400 ne
rect -30974 -35248 -9026 -34400
tri -9026 -35248 -8178 -34400 nw
tri -8178 -35248 -7330 -34400 se
rect -7330 -35248 -2521 -34400
tri -2521 -35248 -800 -33527 nw
rect -33727 -36096 -31822 -35248
tri -31822 -36096 -30974 -35248 sw
tri -30974 -36096 -30126 -35248 ne
rect -30126 -36096 -9874 -35248
tri -9874 -36096 -9026 -35248 nw
tri -9026 -36096 -8178 -35248 se
rect -8178 -36096 -5400 -35248
rect -33727 -36704 -30974 -36096
tri -30974 -36704 -30366 -36096 sw
tri -30126 -36704 -29518 -36096 ne
rect -29518 -36704 -10482 -36096
tri -10482 -36704 -9874 -36096 nw
tri -9634 -36704 -9026 -36096 se
rect -9026 -36704 -5400 -36096
rect -33727 -37552 -30366 -36704
tri -30366 -37552 -29518 -36704 sw
tri -29518 -37552 -28670 -36704 ne
rect -28670 -37552 -11330 -36704
tri -11330 -37552 -10482 -36704 nw
tri -10482 -37552 -9634 -36704 se
rect -9634 -37552 -5400 -36704
rect -33727 -38400 -29518 -37552
tri -29518 -38400 -28670 -37552 sw
tri -28670 -38400 -27822 -37552 ne
rect -27822 -38400 -12178 -37552
tri -12178 -38400 -11330 -37552 nw
tri -11330 -38400 -10482 -37552 se
rect -10482 -38127 -5400 -37552
tri -5400 -38127 -2521 -35248 nw
rect -10482 -38400 -6273 -38127
rect -33727 -39000 -28670 -38400
tri -28670 -39000 -28070 -38400 sw
tri -11930 -39000 -11330 -38400 se
rect -11330 -39000 -6273 -38400
tri -6273 -39000 -5400 -38127 nw
tri -33727 -40905 -31822 -39000 ne
rect -31822 -40905 -8178 -39000
tri -8178 -40905 -6273 -39000 nw
tri -31822 -43000 -29727 -40905 ne
rect -29727 -43000 -10273 -40905
tri -10273 -43000 -8178 -40905 nw
<< end >>
