magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< nwell >>
rect -36 679 1484 1471
<< poly >>
rect 114 740 144 907
rect 81 674 144 740
rect 114 507 144 674
<< locali >>
rect 0 1397 1448 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1346 1297 1380 1397
rect 64 674 98 740
rect 704 724 738 1096
rect 704 690 755 724
rect 704 318 738 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1346 17 1380 104
rect 0 -17 1448 17
use sky130_sram_1r1w_24x128_8_contact_15  sky130_sram_1r1w_24x128_8_contact_15_0
timestamp 1661296025
transform 1 0 48 0 1 674
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_28  sky130_sram_1r1w_24x128_8_contact_28_0
timestamp 1661296025
transform 1 0 1338 0 1 1256
box -59 -43 109 125
use sky130_sram_1r1w_24x128_8_contact_29  sky130_sram_1r1w_24x128_8_contact_29_0
timestamp 1661296025
transform 1 0 1338 0 1 63
box -26 -26 76 108
use sky130_sram_1r1w_24x128_8_nmos_m11_w2_000_sli_dli_da_p  sky130_sram_1r1w_24x128_8_nmos_m11_w2_000_sli_dli_da_p_0
timestamp 1661296025
transform 1 0 54 0 1 51
box -26 -26 1256 456
use sky130_sram_1r1w_24x128_8_pmos_m11_w2_000_sli_dli_da_p  sky130_sram_1r1w_24x128_8_pmos_m11_w2_000_sli_dli_da_p_0
timestamp 1661296025
transform 1 0 54 0 1 963
box -59 -56 1289 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 738 707 738 707 4 Z
port 2 nsew
rlabel locali s 724 0 724 0 4 gnd
port 3 nsew
rlabel locali s 724 1414 724 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1448 1414
<< end >>
