** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/untitled-9.sch
**.subckt untitled-9
V1 net1 GND DC 0.9 AC 1
R1 n1 net1 1k m=1
XC1 n1 GND sky130_fd_pr__cap_mim_m3_1 W=1e7u L=1e6u MF=1 m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice ff
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice



.options savecurrents
.AC dec 1000 10M 10G
.control
run
display
plot v(n1)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
