* NGSPICE file created from flat3.ext - technology: sky130B

X0 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X1 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X2 captuner_complete_1_r_0/TOP RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__cap_mim_m3_2 l=4.4e+07u w=5e+07u
X3 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X5 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X6 captuner_complete_1_r_0/TOP captuner_complete_1_r_0/BOT_C1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2.5e+06u
X7 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X8 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X9 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X10 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X11 RF_nfet_12xW5p0L0p15_0/S captuner_complete_1_r_0/TOP sky130_fd_pr__cap_mim_m3_1 l=4.4e+07u w=5e+07u
X12 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__cap_mim_m3_2 l=7.5e+06u w=4.5e+06u
X13 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X14 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X15 BIAS_BOT RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__cap_mim_m3_2 l=1.15e+07u w=9.5e+06u
X16 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X17 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X18 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X19 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X20 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X21 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X22 RF_nfet_12xW5p0L0p15_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G sky130_fd_pr__cap_mim_m3_1 l=7.5e+06u w=4.5e+06u
X23 captuner_complete_1_r_0/BOT_C1 captuner_complete_1_r_0/G1 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X24 captuner_complete_1_r_0/BOT_C4 captuner_complete_1_r_0/G4 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X25 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
R0 RFB_MID RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S sky130_fd_pr__res_generic_po w=330000u l=1.28e+07u
X26 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X27 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S captuner_complete_1_r_0/G2 captuner_complete_1_r_0/BOT_C2 RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X28 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S captuner_complete_1_r_0/G8 captuner_complete_1_r_0/BOT_C8 RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X29 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X30 RF_nfet_12xW5p0L0p15_0/S BIAS_BOT sky130_fd_pr__cap_mim_m3_1 l=1.15e+07u w=9.5e+06u
X31 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X32 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X33 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X34 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X35 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X36 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X37 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X38 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X39 captuner_complete_1_r_0/TOP captuner_complete_1_r_0/BOT_C8 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=8e+06u
X40 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X41 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RFB_MID sky130_fd_pr__cap_mim_m3_2 l=2.05e+07u w=1.15e+07u
X42 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S captuner_complete_1_r_0/G1 captuner_complete_1_r_0/BOT_C1 RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X43 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S captuner_complete_1_r_0/G4 captuner_complete_1_r_0/BOT_C4 RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X44 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X45 captuner_complete_1_r_0/BOT_C8 captuner_complete_1_r_0/G8 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
R1 captuner_complete_1_r_0/TOP RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G sky130_fd_pr__res_generic_po w=330000u l=1.28e+07u
X46 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
R2 BIAS_BOT RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G sky130_fd_pr__res_generic_po w=330000u l=2.068e+07u
X47 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X48 RFB_MID RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G sky130_fd_pr__cap_mim_m3_1 l=2.05e+07u w=1.15e+07u
X49 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X50 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X51 captuner_complete_1_r_0/TOP captuner_complete_1_r_0/BOT_C4 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=4e+06u
X52 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X53 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X54 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X55 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X56 captuner_complete_1_r_0/TOP captuner_complete_1_r_0/BOT_C2 sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=2.5e+06u
X57 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X58 captuner_complete_1_r_0/BOT_C2 captuner_complete_1_r_0/G2 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X59 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
C0 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G 3.39fF
C1 captuner_complete_1_r_0/BOT_C1 captuner_complete_1_r_0/TOP 1.16fF
C2 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RFB_MID 40.06fF
C3 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G m5_n800_n3000# 1.17fF
C4 captuner_complete_1_r_0/BOT_C4 captuner_complete_1_r_0/TOP 2.60fF
C5 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S captuner_complete_1_r_0/BOT_C1 3.57fF
C6 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S 26.96fF
C7 captuner_complete_1_r_0/BOT_C4 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S 3.94fF
C8 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S captuner_complete_1_r_0/TOP 2.58fF
C9 captuner_complete_1_r_0/BOT_C8 captuner_complete_1_r_0/TOP 4.77fF
C10 captuner_complete_1_r_0/BOT_C2 captuner_complete_1_r_0/TOP 1.89fF
C11 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S m5_n800_n3000# 3.92fF
C12 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S 41.75fF
C13 captuner_complete_1_r_0/BOT_C8 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S 4.73fF
C14 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G 6.12fF
C15 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S captuner_complete_1_r_0/BOT_C2 3.54fF
C16 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G BIAS_BOT 2.13fF
C17 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S 14.77fF
C18 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G 3.11fF
C19 BIAS_BOT RF_nfet_12xW5p0L0p15_0/S 28.25fF $ **FLOATING
C20 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S 11.11fF $ **FLOATING
C21 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S 16.95fF $ **FLOATING
C22 RF_nfet_8xW5p0L0p15_1_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/S 23.70fF $ **FLOATING
C23 RFB_MID RF_nfet_12xW5p0L0p15_0/S 5.66fF $ **FLOATING
C24 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/D RF_nfet_12xW5p0L0p15_0/S 17.90fF $ **FLOATING
C25 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/G RF_nfet_12xW5p0L0p15_0/S 20.65fF $ **FLOATING
C26 captuner_complete_1_r_0/TOP RF_nfet_12xW5p0L0p15_0/S 432.32fF $ **FLOATING
C27 captuner_complete_1_r_0/BOT_C4 RF_nfet_12xW5p0L0p15_0/S 3.60fF $ **FLOATING
C28 captuner_complete_1_r_0/BOT_C8 RF_nfet_12xW5p0L0p15_0/S 3.33fF $ **FLOATING
C29 captuner_complete_1_r_0/BOT_C1 RF_nfet_12xW5p0L0p15_0/S 3.02fF $ **FLOATING
C30 RF_nfet_12xW5p0L0p15_0/sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0/S RF_nfet_12xW5p0L0p15_0/S 54.66fF $ **FLOATING
C31 captuner_complete_1_r_0/BOT_C2 RF_nfet_12xW5p0L0p15_0/S 3.12fF $ **FLOATING
C32 captuner_complete_1_r_0/G4 RF_nfet_12xW5p0L0p15_0/S 1.28fF $ **FLOATING
C33 captuner_complete_1_r_0/G8 RF_nfet_12xW5p0L0p15_0/S 1.10fF $ **FLOATING
C34 captuner_complete_1_r_0/G1 RF_nfet_12xW5p0L0p15_0/S 1.06fF $ **FLOATING
C35 captuner_complete_1_r_0/G2 RF_nfet_12xW5p0L0p15_0/S 1.29fF $ **FLOATING
