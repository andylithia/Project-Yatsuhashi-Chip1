magic
tech sky130B
magscale 1 2
timestamp 1661375332
<< metal1 >>
rect -2513 -1061 -2269 -1011
rect -2513 -1283 -2475 -1061
rect -2315 -1283 -2269 -1061
rect -2513 -1357 -2269 -1283
rect 162602 -1522 162846 -1472
rect -2485 -1854 -1961 -1677
rect 162602 -1744 162640 -1522
rect 162800 -1744 162846 -1522
rect 162602 -1818 162846 -1744
rect -2558 -2248 -1824 -1854
rect 162630 -2688 163154 -2138
<< via1 >>
rect -2475 -1283 -2315 -1061
rect 162640 -1744 162800 -1522
<< metal2 >>
rect -2505 -1061 -2281 -1027
rect -2505 -1283 -2475 -1061
rect -2315 -1283 -2281 -1061
rect -2505 -1307 -2281 -1283
rect 162610 -1522 162834 -1488
rect 162610 -1744 162640 -1522
rect 162800 -1744 162834 -1522
rect 162610 -1768 162834 -1744
<< via2 >>
rect -2475 -1279 -2321 -1061
rect 162640 -1740 162794 -1522
<< metal3 >>
rect -3600 -214 163800 -200
rect -3600 -1061 329732 -214
rect -3600 -1200 -2475 -1061
rect -2697 -1279 -2475 -1200
rect -2321 -1200 329732 -1061
rect -2321 -1279 -1857 -1200
rect 162332 -1214 329732 -1200
rect -2697 -1375 -1857 -1279
rect 162418 -1522 163258 -1214
rect 162418 -1740 162640 -1522
rect 162794 -1740 163258 -1522
rect 162418 -1836 163258 -1740
use sky130_fd_pr__res_generic_po_V3RDUA  sky130_fd_pr__res_generic_po_V3RDUA_0
timestamp 0
transform 1 0 162698 0 1 -1983
box -199 -404 199 404
use sky130_fd_pr__res_generic_po_V3RDUA  sky130_fd_pr__res_generic_po_V3RDUA_1
timestamp 0
transform 1 0 -2417 0 1 -1522
box -199 -404 199 404
<< labels >>
rlabel metal3 -3600 -1200 -2200 -200 1 A
rlabel metal3 162400 -1200 163800 -200 1 B
rlabel metal1 162636 -2688 163128 -2472 1 B1
rlabel metal1 -2464 -2180 -1924 -1978 1 A1
<< end >>
