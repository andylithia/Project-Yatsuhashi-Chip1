magic
tech sky130B
magscale 1 2
timestamp 1661315583
<< metal4 >>
rect -44100 -23712 -30900 -23600
rect -44100 -27088 -34388 -23712
rect -31012 -27088 -30900 -23712
rect -44100 -27200 -30900 -27088
<< via4 >>
rect -34388 -27088 -31012 -23712
<< metal5 >>
tri -36055 1400 -32455 5000 se
rect -32455 1400 -11745 5000
tri -11745 1400 -8145 5000 sw
tri -37667 -212 -36055 1400 se
rect -36055 800 -31564 1400
tri -31564 800 -30964 1400 nw
tri -13236 800 -12636 1400 ne
rect -12636 800 -8145 1400
rect -36055 -48 -32412 800
tri -32412 -48 -31564 800 nw
tri -31564 -48 -30716 800 se
rect -30716 -48 -13484 800
tri -13484 -48 -12636 800 sw
tri -12636 -48 -11788 800 ne
rect -11788 -48 -8145 800
rect -36055 -212 -32576 -48
tri -32576 -212 -32412 -48 nw
tri -31728 -212 -31564 -48 se
rect -31564 -212 -12636 -48
tri -39300 -1845 -37667 -212 se
rect -37667 -1060 -33424 -212
tri -33424 -1060 -32576 -212 nw
tri -32576 -1060 -31728 -212 se
rect -31728 -896 -12636 -212
tri -12636 -896 -11788 -48 sw
tri -11788 -896 -10940 -48 ne
rect -10940 -896 -8145 -48
rect -31728 -1060 -11788 -896
rect -37667 -1845 -34272 -1060
tri -40191 -2736 -39300 -1845 se
rect -39300 -1908 -34272 -1845
tri -34272 -1908 -33424 -1060 nw
tri -33424 -1908 -32576 -1060 se
rect -32576 -1104 -11788 -1060
tri -11788 -1104 -11580 -896 sw
tri -10940 -1104 -10732 -896 ne
rect -10732 -1104 -8145 -896
rect -32576 -1908 -11580 -1104
rect -39300 -2736 -35100 -1908
tri -35100 -2736 -34272 -1908 nw
tri -34252 -2736 -33424 -1908 se
rect -33424 -1952 -11580 -1908
tri -11580 -1952 -10732 -1104 sw
tri -10732 -1952 -9884 -1104 ne
rect -9884 -1952 -8145 -1104
rect -33424 -2736 -10732 -1952
tri -43500 -6045 -40191 -2736 se
rect -40191 -3584 -35948 -2736
tri -35948 -3584 -35100 -2736 nw
tri -34316 -2800 -34252 -2736 se
rect -34252 -2800 -10732 -2736
tri -10732 -2800 -9884 -1952 sw
tri -9884 -2800 -9036 -1952 ne
rect -9036 -2800 -8145 -1952
tri -8145 -2800 -3945 1400 sw
tri -35100 -3584 -34316 -2800 se
rect -34316 -3400 -29824 -2800
tri -29824 -3400 -29224 -2800 nw
tri -14976 -3400 -14376 -2800 ne
rect -14376 -3400 -9884 -2800
rect -34316 -3584 -30672 -3400
rect -40191 -4432 -36796 -3584
tri -36796 -4432 -35948 -3584 nw
tri -35948 -4432 -35100 -3584 se
rect -35100 -4248 -30672 -3584
tri -30672 -4248 -29824 -3400 nw
tri -29824 -4248 -28976 -3400 se
rect -28976 -4248 -15224 -3400
tri -15224 -4248 -14376 -3400 sw
tri -14376 -4248 -13528 -3400 ne
rect -13528 -3648 -9884 -3400
tri -9884 -3648 -9036 -2800 sw
tri -9036 -3648 -8188 -2800 ne
rect -8188 -3648 -3945 -2800
rect -13528 -4248 -9036 -3648
rect -35100 -4432 -31520 -4248
rect -40191 -5280 -37644 -4432
tri -37644 -5280 -36796 -4432 nw
tri -36796 -5280 -35948 -4432 se
rect -35948 -5096 -31520 -4432
tri -31520 -5096 -30672 -4248 nw
tri -30672 -5096 -29824 -4248 se
rect -29824 -5096 -14376 -4248
tri -14376 -5096 -13528 -4248 sw
tri -13528 -5096 -12680 -4248 ne
rect -12680 -4496 -9036 -4248
tri -9036 -4496 -8188 -3648 sw
tri -8188 -4496 -7340 -3648 ne
rect -7340 -4496 -3945 -3648
rect -12680 -5096 -8188 -4496
rect -35948 -5280 -31728 -5096
rect -40191 -5304 -37668 -5280
tri -37668 -5304 -37644 -5280 nw
tri -36820 -5304 -36796 -5280 se
rect -36796 -5304 -31728 -5280
tri -31728 -5304 -31520 -5096 nw
tri -30880 -5304 -30672 -5096 se
rect -30672 -5304 -13528 -5096
tri -13528 -5304 -13320 -5096 sw
tri -12680 -5304 -12472 -5096 ne
rect -12472 -5304 -8188 -5096
tri -8188 -5304 -7380 -4496 sw
tri -7340 -5304 -6532 -4496 ne
rect -6532 -5304 -3945 -4496
rect -40191 -6045 -38516 -5304
tri -44391 -6936 -43500 -6045 se
rect -43500 -6152 -38516 -6045
tri -38516 -6152 -37668 -5304 nw
tri -37668 -6152 -36820 -5304 se
rect -36820 -6152 -32576 -5304
tri -32576 -6152 -31728 -5304 nw
tri -31728 -6152 -30880 -5304 se
rect -30880 -6152 -13320 -5304
tri -13320 -6152 -12472 -5304 sw
tri -12472 -6152 -11624 -5304 ne
rect -11624 -6152 -7380 -5304
tri -7380 -6152 -6532 -5304 sw
tri -6532 -6152 -5684 -5304 ne
rect -5684 -6152 -3945 -5304
rect -43500 -6936 -39300 -6152
tri -39300 -6936 -38516 -6152 nw
tri -38452 -6936 -37668 -6152 se
rect -37668 -6936 -33424 -6152
tri -47100 -9645 -44391 -6936 se
rect -44391 -7784 -40148 -6936
tri -40148 -7784 -39300 -6936 nw
tri -39300 -7784 -38452 -6936 se
rect -38452 -7000 -33424 -6936
tri -33424 -7000 -32576 -6152 nw
tri -32576 -7000 -31728 -6152 se
rect -31728 -7000 -12472 -6152
tri -12472 -7000 -11624 -6152 sw
tri -11624 -7000 -10776 -6152 ne
rect -10776 -7000 -6532 -6152
tri -6532 -7000 -5684 -6152 sw
tri -5684 -7000 -4836 -6152 ne
rect -4836 -7000 -3945 -6152
tri -3945 -7000 255 -2800 sw
rect -38452 -7784 -34272 -7000
rect -44391 -8632 -40996 -7784
tri -40996 -8632 -40148 -7784 nw
tri -40148 -8632 -39300 -7784 se
rect -39300 -7848 -34272 -7784
tri -34272 -7848 -33424 -7000 nw
tri -33424 -7848 -32576 -7000 se
rect -39300 -8632 -35100 -7848
rect -44391 -8676 -41040 -8632
tri -41040 -8676 -40996 -8632 nw
tri -40192 -8676 -40148 -8632 se
rect -40148 -8676 -35100 -8632
tri -35100 -8676 -34272 -7848 nw
tri -34252 -8676 -33424 -7848 se
rect -33424 -8676 -32576 -7848
rect -44391 -9524 -41888 -8676
tri -41888 -9524 -41040 -8676 nw
tri -41040 -9524 -40192 -8676 se
rect -40192 -9524 -35948 -8676
tri -35948 -9524 -35100 -8676 nw
tri -35100 -9524 -34252 -8676 se
rect -34252 -9524 -32576 -8676
rect -44391 -9645 -42052 -9524
rect -47100 -9688 -42052 -9645
tri -42052 -9688 -41888 -9524 nw
tri -41204 -9688 -41040 -9524 se
rect -41040 -9688 -36796 -9524
rect -47100 -10536 -42900 -9688
tri -42900 -10536 -42052 -9688 nw
tri -42052 -10536 -41204 -9688 se
rect -41204 -10372 -36796 -9688
tri -36796 -10372 -35948 -9524 nw
tri -35948 -10372 -35100 -9524 se
rect -35100 -10372 -32576 -9524
rect -41204 -10536 -37644 -10372
rect -47100 -16400 -43500 -10536
tri -43500 -11136 -42900 -10536 nw
tri -42652 -11136 -42052 -10536 se
rect -42052 -11136 -37644 -10536
tri -42900 -11384 -42652 -11136 se
rect -42652 -11220 -37644 -11136
tri -37644 -11220 -36796 -10372 nw
tri -36796 -11220 -35948 -10372 se
rect -35948 -11220 -32576 -10372
rect -42652 -11243 -37667 -11220
tri -37667 -11243 -37644 -11220 nw
tri -36819 -11243 -36796 -11220 se
rect -36796 -11243 -32576 -11220
rect -42652 -11384 -38515 -11243
rect -42900 -12091 -38515 -11384
tri -38515 -12091 -37667 -11243 nw
tri -37667 -12091 -36819 -11243 se
rect -36819 -12091 -32576 -11243
tri -32576 -12091 -27485 -7000 nw
tri -16715 -12091 -11624 -7000 ne
tri -11624 -7848 -10776 -7000 sw
tri -10776 -7848 -9928 -7000 ne
rect -9928 -7848 -5684 -7000
tri -5684 -7848 -4836 -7000 sw
tri -4836 -7848 -3988 -7000 ne
rect -3988 -7848 255 -7000
rect -11624 -8676 -10776 -7848
tri -10776 -8676 -9948 -7848 sw
tri -9928 -8676 -9100 -7848 ne
rect -9100 -8676 -4836 -7848
tri -4836 -8676 -4008 -7848 sw
tri -3988 -8676 -3160 -7848 ne
rect -3160 -8676 255 -7848
rect -11624 -9524 -9948 -8676
tri -9948 -9524 -9100 -8676 sw
tri -9100 -9524 -8252 -8676 ne
rect -8252 -9524 -4008 -8676
tri -4008 -9524 -3160 -8676 sw
tri -3160 -9524 -2312 -8676 ne
rect -2312 -9524 255 -8676
rect -11624 -10372 -9100 -9524
tri -9100 -10372 -8252 -9524 sw
tri -8252 -10372 -7404 -9524 ne
rect -7404 -10372 -3160 -9524
tri -3160 -10372 -2312 -9524 sw
tri -2312 -10372 -1464 -9524 ne
rect -1464 -9645 255 -9524
tri 255 -9645 2900 -7000 sw
rect -1464 -10372 2900 -9645
rect -11624 -11220 -8252 -10372
tri -8252 -11220 -7404 -10372 sw
tri -7404 -11220 -6556 -10372 ne
rect -6556 -11136 -2312 -10372
tri -2312 -11136 -1548 -10372 sw
tri -1464 -11136 -700 -10372 ne
rect -6556 -11220 -1548 -11136
rect -11624 -11428 -7404 -11220
tri -7404 -11428 -7196 -11220 sw
tri -6556 -11428 -6348 -11220 ne
rect -6348 -11384 -1548 -11220
tri -1548 -11384 -1300 -11136 sw
rect -6348 -11428 -1300 -11384
rect -11624 -12091 -7196 -11428
rect -42900 -30694 -39300 -12091
tri -39300 -12876 -38515 -12091 nw
tri -38452 -12876 -37667 -12091 se
rect -37667 -12876 -35100 -12091
tri -38700 -13124 -38452 -12876 se
rect -38452 -13124 -35100 -12876
rect -38700 -28955 -35100 -13124
tri -35100 -14615 -32576 -12091 nw
tri -11624 -14615 -9100 -12091 ne
rect -9100 -12276 -7196 -12091
tri -7196 -12276 -6348 -11428 sw
tri -6348 -12276 -5500 -11428 ne
rect -5500 -12276 -1300 -11428
rect -9100 -13124 -6348 -12276
tri -6348 -13124 -5500 -12276 sw
tri -5500 -12876 -4900 -12276 ne
rect -34500 -23712 -30900 -23600
rect -34500 -27088 -34388 -23712
rect -31012 -27088 -30900 -23712
rect -34500 -28106 -30900 -27088
tri -35100 -28955 -34500 -28355 sw
tri -34500 -28955 -33651 -28106 ne
rect -33651 -28955 -30900 -28106
rect -38700 -29804 -34500 -28955
tri -34500 -29804 -33651 -28955 sw
tri -33651 -29804 -32802 -28955 ne
rect -32802 -29804 -30900 -28955
rect -38700 -29846 -33651 -29804
tri -39300 -30694 -38700 -30094 sw
tri -38700 -30694 -37852 -29846 ne
rect -37852 -30008 -33651 -29846
tri -33651 -30008 -33447 -29804 sw
tri -32802 -30008 -32598 -29804 ne
rect -32598 -30008 -30900 -29804
rect -37852 -30694 -33447 -30008
rect -42900 -30858 -38700 -30694
tri -38700 -30858 -38536 -30694 sw
tri -37852 -30858 -37688 -30694 ne
rect -37688 -30857 -33447 -30694
tri -33447 -30857 -32598 -30008 sw
tri -32598 -30857 -31749 -30008 ne
rect -31749 -30857 -30900 -30008
rect -37688 -30858 -32598 -30857
rect -42900 -31585 -38536 -30858
tri -42900 -31706 -42779 -31585 ne
rect -42779 -31706 -38536 -31585
tri -38536 -31706 -37688 -30858 sw
tri -37688 -31706 -36840 -30858 ne
rect -36840 -31706 -32598 -30858
tri -32598 -31706 -31749 -30857 sw
tri -31749 -31706 -30900 -30857 ne
tri -30900 -31706 -25809 -26615 sw
tri -10394 -27909 -9100 -26615 se
rect -9100 -27909 -5500 -13124
tri -14191 -31706 -10394 -27909 se
rect -10394 -28106 -5500 -27909
rect -10394 -28955 -6349 -28106
tri -6349 -28955 -5500 -28106 nw
tri -5500 -28955 -4900 -28355 se
rect -4900 -28955 -1300 -12276
rect -10394 -29804 -7198 -28955
tri -7198 -29804 -6349 -28955 nw
tri -6349 -29804 -5500 -28955 se
rect -5500 -29804 -1300 -28955
rect -10394 -30653 -8047 -29804
tri -8047 -30653 -7198 -29804 nw
tri -7198 -30653 -6349 -29804 se
rect -6349 -29846 -1300 -29804
rect -6349 -30653 -2148 -29846
rect -10394 -31302 -8696 -30653
tri -8696 -31302 -8047 -30653 nw
tri -7847 -31302 -7198 -30653 se
rect -7198 -30694 -2148 -30653
tri -2148 -30694 -1300 -29846 nw
tri -1300 -30694 -700 -30094 se
rect -700 -30694 2900 -10372
rect -7198 -31302 -2996 -30694
rect -10394 -31706 -9545 -31302
tri -42779 -36797 -37688 -31706 ne
tri -37688 -32554 -36840 -31706 sw
tri -36840 -32554 -35992 -31706 ne
rect -35992 -32554 -31749 -31706
rect -37688 -33402 -36840 -32554
tri -36840 -33402 -35992 -32554 sw
tri -35992 -33402 -35144 -32554 ne
rect -35144 -32555 -31749 -32554
tri -31749 -32555 -30900 -31706 sw
tri -30900 -32555 -30051 -31706 ne
rect -30051 -32555 -25809 -31706
rect -35144 -33000 -30900 -32555
tri -30900 -33000 -30455 -32555 sw
tri -30051 -33000 -29606 -32555 ne
rect -29606 -33000 -25809 -32555
tri -25809 -33000 -24515 -31706 sw
tri -15485 -33000 -14191 -31706 se
rect -14191 -32151 -9545 -31706
tri -9545 -32151 -8696 -31302 nw
tri -8696 -32151 -7847 -31302 se
rect -7847 -31542 -2996 -31302
tri -2996 -31542 -2148 -30694 nw
tri -2148 -31542 -1300 -30694 se
rect -1300 -31542 2900 -30694
rect -7847 -32151 -3607 -31542
rect -14191 -33000 -10394 -32151
tri -10394 -33000 -9545 -32151 nw
tri -9545 -33000 -8696 -32151 se
rect -8696 -32153 -3607 -32151
tri -3607 -32153 -2996 -31542 nw
tri -2759 -32153 -2148 -31542 se
rect -2148 -31585 2900 -31542
rect -2148 -32153 -700 -31585
rect -8696 -33000 -4455 -32153
rect -35144 -33402 -30455 -33000
rect -37688 -34250 -35992 -33402
tri -35992 -34250 -35144 -33402 sw
tri -35144 -34250 -34296 -33402 ne
rect -34296 -33849 -30455 -33402
tri -30455 -33849 -29606 -33000 sw
tri -29606 -33849 -28757 -33000 ne
rect -28757 -33849 -11243 -33000
tri -11243 -33849 -10394 -33000 nw
tri -10394 -33849 -9545 -33000 se
rect -9545 -33001 -4455 -33000
tri -4455 -33001 -3607 -32153 nw
tri -3607 -33001 -2759 -32153 se
rect -2759 -33001 -700 -32153
rect -9545 -33849 -5303 -33001
tri -5303 -33849 -4455 -33001 nw
tri -4455 -33849 -3607 -33001 se
rect -3607 -33849 -700 -33001
rect -34296 -34250 -29606 -33849
rect -37688 -34253 -35144 -34250
tri -35144 -34253 -35141 -34250 sw
tri -34296 -34253 -34293 -34250 ne
rect -34293 -34253 -29606 -34250
rect -37688 -35101 -35141 -34253
tri -35141 -35101 -34293 -34253 sw
tri -34293 -35101 -33445 -34253 ne
rect -33445 -34698 -29606 -34253
tri -29606 -34698 -28757 -33849 sw
tri -28757 -34698 -27908 -33849 ne
rect -27908 -34698 -12092 -33849
tri -12092 -34698 -11243 -33849 nw
tri -11243 -34698 -10394 -33849 se
rect -10394 -34697 -6151 -33849
tri -6151 -34697 -5303 -33849 nw
tri -5303 -34697 -4455 -33849 se
rect -4455 -34697 -700 -33849
rect -10394 -34698 -6999 -34697
rect -33445 -34902 -28757 -34698
tri -28757 -34902 -28553 -34698 sw
tri -27908 -34902 -27704 -34698 ne
rect -27704 -34902 -12296 -34698
tri -12296 -34902 -12092 -34698 nw
tri -11447 -34902 -11243 -34698 se
rect -11243 -34902 -6999 -34698
rect -33445 -35101 -28553 -34902
rect -37688 -35949 -34293 -35101
tri -34293 -35949 -33445 -35101 sw
tri -33445 -35949 -32597 -35101 ne
rect -32597 -35751 -28553 -35101
tri -28553 -35751 -27704 -34902 sw
tri -27704 -35751 -26855 -34902 ne
rect -26855 -35751 -13145 -34902
tri -13145 -35751 -12296 -34902 nw
tri -12296 -35751 -11447 -34902 se
rect -11447 -35545 -6999 -34902
tri -6999 -35545 -6151 -34697 nw
tri -6151 -35545 -5303 -34697 se
rect -5303 -35185 -700 -34697
tri -700 -35185 2900 -31585 nw
rect -11447 -35751 -7806 -35545
rect -32597 -35949 -27704 -35751
rect -37688 -36797 -33445 -35949
tri -33445 -36797 -32597 -35949 sw
tri -32597 -36797 -31749 -35949 ne
rect -31749 -36600 -27704 -35949
tri -27704 -36600 -26855 -35751 sw
tri -26855 -36600 -26006 -35751 ne
rect -26006 -36600 -13994 -35751
tri -13994 -36600 -13145 -35751 nw
tri -13145 -36600 -12296 -35751 se
rect -12296 -36352 -7806 -35751
tri -7806 -36352 -6999 -35545 nw
tri -6958 -36352 -6151 -35545 se
rect -6151 -36352 -5303 -35545
rect -12296 -36600 -8654 -36352
rect -31749 -36797 -26855 -36600
tri -37688 -41400 -33085 -36797 ne
rect -33085 -37645 -32597 -36797
tri -32597 -37645 -31749 -36797 sw
tri -31749 -37645 -30901 -36797 ne
rect -30901 -37200 -26855 -36797
tri -26855 -37200 -26255 -36600 sw
tri -13745 -37200 -13145 -36600 se
rect -13145 -37200 -8654 -36600
tri -8654 -37200 -7806 -36352 nw
tri -7806 -37200 -6958 -36352 se
rect -6958 -37200 -5303 -36352
rect -30901 -37645 -9502 -37200
rect -33085 -38493 -31749 -37645
tri -31749 -38493 -30901 -37645 sw
tri -30901 -38493 -30053 -37645 ne
rect -30053 -38048 -9502 -37645
tri -9502 -38048 -8654 -37200 nw
tri -8654 -38048 -7806 -37200 se
rect -7806 -38048 -5303 -37200
rect -30053 -38092 -9546 -38048
tri -9546 -38092 -9502 -38048 nw
tri -8698 -38092 -8654 -38048 se
rect -8654 -38092 -5303 -38048
rect -30053 -38493 -10394 -38092
rect -33085 -39104 -30901 -38493
tri -30901 -39104 -30290 -38493 sw
tri -30053 -39104 -29442 -38493 ne
rect -29442 -38940 -10394 -38493
tri -10394 -38940 -9546 -38092 nw
tri -9546 -38940 -8698 -38092 se
rect -8698 -38940 -5303 -38092
rect -29442 -39104 -11242 -38940
rect -33085 -39952 -30290 -39104
tri -30290 -39952 -29442 -39104 sw
tri -29442 -39952 -28594 -39104 ne
rect -28594 -39788 -11242 -39104
tri -11242 -39788 -10394 -38940 nw
tri -10394 -39788 -9546 -38940 se
rect -9546 -39788 -5303 -38940
tri -5303 -39788 -700 -35185 nw
rect -28594 -39952 -11406 -39788
tri -11406 -39952 -11242 -39788 nw
tri -10558 -39952 -10394 -39788 se
rect -33085 -40800 -29442 -39952
tri -29442 -40800 -28594 -39952 sw
tri -28594 -40800 -27746 -39952 ne
rect -27746 -40800 -12254 -39952
tri -12254 -40800 -11406 -39952 nw
tri -11406 -40800 -10558 -39952 se
rect -10558 -40800 -10394 -39952
rect -33085 -41400 -28594 -40800
tri -28594 -41400 -27994 -40800 sw
tri -12006 -41400 -11406 -40800 se
rect -11406 -41400 -10394 -40800
tri -33085 -45000 -29485 -41400 ne
rect -29485 -44879 -10394 -41400
tri -10394 -44879 -5303 -39788 nw
rect -29485 -45000 -10515 -44879
tri -10515 -45000 -10394 -44879 nw
<< end >>
