magic
tech sky130A
timestamp 0
<< end >>
