** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/untitled-7.sch
**.subckt untitled-7
V1 net2 GND 1
V2 net1 GND 1.8
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice ff
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice



.options savecurrents
* .tran 1ps 20ns
let vlim=1.8
.dc V1 0.1 1.8 0.1
.control
run
display
* print @m.xm1.msky130_fd_pr__nfet_05v0_nvt[id]
plot @v1[dc]/@r1[i]
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
