magic
tech sky130A
timestamp 1658635593
<< error_p >>
rect 345 311 352 547
rect 690 311 697 547
rect 1040 311 1042 547
rect 345 50 352 286
rect 690 50 697 286
rect 1040 50 1042 286
<< metal1 >>
rect 13 647 1015 705
rect 13 50 42 647
rect 80 615 260 620
rect 80 585 85 615
rect 115 585 125 615
rect 155 585 165 615
rect 195 585 205 615
rect 235 585 260 615
rect 80 564 260 585
rect 296 50 387 647
rect 427 615 607 620
rect 427 585 432 615
rect 462 585 472 615
rect 502 585 512 615
rect 542 585 552 615
rect 582 585 607 615
rect 427 564 607 585
rect 641 50 732 647
rect 770 615 950 620
rect 770 585 775 615
rect 805 585 815 615
rect 845 585 855 615
rect 885 585 895 615
rect 925 585 950 615
rect 770 564 950 585
rect 986 50 1015 647
rect 80 30 260 35
rect 80 0 85 30
rect 115 0 125 30
rect 155 0 165 30
rect 195 0 205 30
rect 235 0 260 30
rect 80 -21 260 0
rect 425 30 605 35
rect 425 0 430 30
rect 460 0 470 30
rect 500 0 510 30
rect 540 0 550 30
rect 580 0 605 30
rect 425 -21 605 0
rect 771 30 951 35
rect 771 0 776 30
rect 806 0 816 30
rect 846 0 856 30
rect 886 0 896 30
rect 926 0 951 30
rect 771 -21 951 0
<< via1 >>
rect 85 585 115 615
rect 125 585 155 615
rect 165 585 195 615
rect 205 585 235 615
rect 432 585 462 615
rect 472 585 502 615
rect 512 585 542 615
rect 552 585 582 615
rect 775 585 805 615
rect 815 585 845 615
rect 855 585 885 615
rect 895 585 925 615
rect 85 0 115 30
rect 125 0 155 30
rect 165 0 195 30
rect 205 0 235 30
rect 430 0 460 30
rect 470 0 500 30
rect 510 0 540 30
rect 550 0 580 30
rect 776 0 806 30
rect 816 0 846 30
rect 856 0 886 30
rect 896 0 926 30
<< metal2 >>
rect 80 575 85 615
rect 115 585 125 615
rect 155 605 165 615
rect 195 605 205 615
rect 235 605 260 615
rect 160 585 165 605
rect 115 575 130 585
rect 160 575 175 585
rect 205 575 220 585
rect 250 575 260 605
rect 80 570 260 575
rect 427 575 432 615
rect 462 585 472 615
rect 502 605 512 615
rect 542 605 552 615
rect 582 605 607 615
rect 507 585 512 605
rect 462 575 477 585
rect 507 575 522 585
rect 552 575 567 585
rect 597 575 607 605
rect 427 570 607 575
rect 770 575 775 615
rect 805 585 815 615
rect 845 605 855 615
rect 885 605 895 615
rect 925 605 950 615
rect 850 585 855 605
rect 805 575 820 585
rect 850 575 865 585
rect 895 575 910 585
rect 940 575 950 605
rect 770 570 950 575
rect 338 311 345 547
rect 683 311 690 547
rect 1028 311 1040 547
rect 338 50 345 286
rect 683 50 690 286
rect 1028 50 1040 286
rect 80 -10 85 30
rect 115 0 125 30
rect 155 20 165 30
rect 195 20 205 30
rect 235 20 260 30
rect 160 0 165 20
rect 115 -10 130 0
rect 160 -10 175 0
rect 205 -10 220 0
rect 250 -10 260 20
rect 80 -15 260 -10
rect 425 -10 430 30
rect 460 0 470 30
rect 500 20 510 30
rect 540 20 550 30
rect 580 20 605 30
rect 505 0 510 20
rect 460 -10 475 0
rect 505 -10 520 0
rect 550 -10 565 0
rect 595 -10 605 20
rect 425 -15 605 -10
rect 771 -10 776 30
rect 806 0 816 30
rect 846 20 856 30
rect 886 20 896 30
rect 926 20 951 30
rect 851 0 856 20
rect 806 -10 821 0
rect 851 -10 866 0
rect 896 -10 911 0
rect 941 -10 951 20
rect 771 -15 951 -10
<< via2 >>
rect 85 585 115 605
rect 130 585 155 605
rect 155 585 160 605
rect 175 585 195 605
rect 195 585 205 605
rect 220 585 235 605
rect 235 585 250 605
rect 85 575 115 585
rect 130 575 160 585
rect 175 575 205 585
rect 220 575 250 585
rect 432 585 462 605
rect 477 585 502 605
rect 502 585 507 605
rect 522 585 542 605
rect 542 585 552 605
rect 567 585 582 605
rect 582 585 597 605
rect 432 575 462 585
rect 477 575 507 585
rect 522 575 552 585
rect 567 575 597 585
rect 775 585 805 605
rect 820 585 845 605
rect 845 585 850 605
rect 865 585 885 605
rect 885 585 895 605
rect 910 585 925 605
rect 925 585 940 605
rect 775 575 805 585
rect 820 575 850 585
rect 865 575 895 585
rect 910 575 940 585
rect 85 0 115 20
rect 130 0 155 20
rect 155 0 160 20
rect 175 0 195 20
rect 195 0 205 20
rect 220 0 235 20
rect 235 0 250 20
rect 85 -10 115 0
rect 130 -10 160 0
rect 175 -10 205 0
rect 220 -10 250 0
rect 430 0 460 20
rect 475 0 500 20
rect 500 0 505 20
rect 520 0 540 20
rect 540 0 550 20
rect 565 0 580 20
rect 580 0 595 20
rect 430 -10 460 0
rect 475 -10 505 0
rect 520 -10 550 0
rect 565 -10 595 0
rect 776 0 806 20
rect 821 0 846 20
rect 846 0 851 20
rect 866 0 886 20
rect 886 0 896 20
rect 911 0 926 20
rect 926 0 941 20
rect 776 -10 806 0
rect 821 -10 851 0
rect 866 -10 896 0
rect 911 -10 941 0
<< metal3 >>
rect 80 605 90 610
rect 130 605 150 610
rect 190 605 210 610
rect 80 575 85 605
rect 205 575 210 605
rect 250 575 260 610
rect 80 570 260 575
rect 427 605 437 610
rect 477 605 497 610
rect 537 605 557 610
rect 427 575 432 605
rect 552 575 557 605
rect 597 575 607 610
rect 427 570 607 575
rect 770 605 780 610
rect 820 605 840 610
rect 880 605 900 610
rect 770 575 775 605
rect 895 575 900 605
rect 940 575 950 610
rect 770 570 950 575
rect 80 20 90 25
rect 130 20 150 25
rect 190 20 210 25
rect 80 -10 85 20
rect 205 -10 210 20
rect 250 -10 260 25
rect 80 -15 260 -10
rect 425 20 435 25
rect 475 20 495 25
rect 535 20 555 25
rect 425 -10 430 20
rect 550 -10 555 20
rect 595 -10 605 25
rect 425 -15 605 -10
rect 771 20 781 25
rect 821 20 841 25
rect 881 20 901 25
rect 771 -10 776 20
rect 896 -10 901 20
rect 941 -10 951 25
rect 771 -15 951 -10
<< via3 >>
rect 90 605 130 610
rect 150 605 190 610
rect 210 605 250 610
rect 90 575 115 605
rect 115 575 130 605
rect 150 575 160 605
rect 160 575 175 605
rect 175 575 190 605
rect 210 575 220 605
rect 220 575 250 605
rect 437 605 477 610
rect 497 605 537 610
rect 557 605 597 610
rect 437 575 462 605
rect 462 575 477 605
rect 497 575 507 605
rect 507 575 522 605
rect 522 575 537 605
rect 557 575 567 605
rect 567 575 597 605
rect 780 605 820 610
rect 840 605 880 610
rect 900 605 940 610
rect 780 575 805 605
rect 805 575 820 605
rect 840 575 850 605
rect 850 575 865 605
rect 865 575 880 605
rect 900 575 910 605
rect 910 575 940 605
rect 90 20 130 25
rect 150 20 190 25
rect 210 20 250 25
rect 90 -10 115 20
rect 115 -10 130 20
rect 150 -10 160 20
rect 160 -10 175 20
rect 175 -10 190 20
rect 210 -10 220 20
rect 220 -10 250 20
rect 435 20 475 25
rect 495 20 535 25
rect 555 20 595 25
rect 435 -10 460 20
rect 460 -10 475 20
rect 495 -10 505 20
rect 505 -10 520 20
rect 520 -10 535 20
rect 555 -10 565 20
rect 565 -10 595 20
rect 781 20 821 25
rect 841 20 881 25
rect 901 20 941 25
rect 781 -10 806 20
rect 806 -10 821 20
rect 841 -10 851 20
rect 851 -10 866 20
rect 866 -10 881 20
rect 901 -10 911 20
rect 911 -10 941 20
<< metal4 >>
rect 80 610 950 620
rect 80 575 90 610
rect 130 575 150 610
rect 190 575 210 610
rect 250 575 437 610
rect 477 575 497 610
rect 537 575 557 610
rect 597 575 780 610
rect 820 575 840 610
rect 880 575 900 610
rect 940 575 950 610
rect 80 555 950 575
rect 80 25 951 35
rect 80 -10 90 25
rect 130 -10 150 25
rect 190 -10 210 25
rect 250 -10 435 25
rect 475 -10 495 25
rect 535 -10 555 25
rect 595 -10 781 25
rect 821 -10 841 25
rect 881 -10 901 25
rect 941 -10 951 25
rect 80 -21 951 -10
rect 80 -30 950 -21
<< labels >>
rlabel metal2 1028 311 1040 547 0 D
port 1 n
rlabel metal2 1028 50 1040 286 0 S
port 2 n
<< end >>
