magic
tech sky130B
timestamp 1662171302
<< metal3 >>
rect 8097 61150 10597 62000
rect 34097 61150 36597 62000
rect 60097 61150 62597 62000
rect 82797 61150 85297 62000
rect 85447 61150 86547 62000
rect 86697 61150 87797 62000
rect 87947 61150 90447 62000
rect 108647 61150 111147 62000
rect 111297 61150 112397 62000
rect 112547 61150 113647 62000
rect 113797 61150 116297 62000
rect 159497 61150 161997 62000
rect 162147 61150 163247 62000
rect 163397 61150 164497 62000
rect 164647 61150 167147 62000
rect 206697 61150 209197 62000
rect 232697 61150 235197 62000
rect 255297 61170 257697 62000
rect 260297 61170 262697 62000
rect 283297 61150 285797 62000
rect 0 50121 850 52621
rect 291150 48992 292000 51492
rect 0 31921 830 34321
rect 291170 29892 292000 32292
rect 0 26921 830 29321
rect 291170 24892 292000 27292
rect 291760 4736 292400 4792
rect 291760 4145 292400 4201
rect 291760 3554 292400 3610
rect 291760 2963 292400 3019
rect 291760 2372 292400 2428
rect 291760 1781 292400 1837
rect 10000 0 10056 200
rect 12700 0 12756 200
rect 15400 0 15456 200
rect 18100 0 18156 200
rect 20800 0 20856 200
rect 23500 0 23556 200
rect 26200 0 26256 200
rect 28900 0 28956 200
rect 31600 0 31656 200
rect 34300 0 34356 200
rect 37000 0 37056 200
rect 39700 0 39756 200
rect 42400 0 42456 200
rect 45100 0 45156 200
rect 47800 0 47856 200
rect 50500 0 50556 200
rect 53200 0 53256 200
rect 55900 0 55956 200
rect 58600 0 58656 200
rect 61300 0 61356 200
rect 64000 0 64056 200
rect 66700 0 66756 200
rect 69400 0 69456 200
rect 72100 0 72156 200
rect 74800 0 74856 200
rect 77500 0 77556 200
rect 80200 0 80256 200
rect 82900 0 82956 200
rect 85600 0 85656 200
rect 88300 0 88356 200
rect 91000 0 91056 200
rect 93700 0 93756 200
rect 96400 0 96456 200
rect 99100 0 99156 200
rect 101800 0 101856 200
rect 104500 0 104556 200
rect 107200 0 107256 200
rect 109900 0 109956 200
rect 112600 0 112656 200
rect 115300 0 115356 200
rect 118000 0 118056 200
rect 120700 0 120756 200
rect 123400 0 123456 200
rect 126100 0 126156 200
rect 128800 0 128856 200
rect 131500 0 131556 200
rect 134200 0 134256 200
rect 136900 0 136956 200
rect 139600 0 139656 200
rect 142300 0 142356 200
rect 145000 0 145056 200
rect 147700 0 147756 200
rect 150400 0 150456 200
rect 153100 0 153156 200
rect 155800 0 155856 200
rect 158500 0 158556 200
rect 161200 0 161256 200
rect 163900 0 163956 200
rect 166600 0 166656 200
rect 169300 0 169356 200
rect 172000 0 172056 200
rect 174700 0 174756 200
rect 177400 0 177456 200
rect 180100 0 180156 200
rect 182800 0 182856 200
rect 185500 0 185556 200
rect 188200 0 188256 200
rect 190900 0 190956 200
rect 193600 0 193656 200
rect 196300 0 196356 200
rect 199000 0 199056 200
rect 201700 0 201756 200
rect 204400 0 204456 200
rect 207100 0 207156 200
rect 209800 0 209856 200
rect 212500 0 212556 200
rect 215200 0 215256 200
rect 217900 0 217956 200
rect 220600 0 220656 200
rect 223300 0 223356 200
rect 226000 0 226056 200
rect 228700 0 228756 200
rect 231400 0 231456 200
rect 234100 0 234156 200
rect 236800 0 236856 200
rect 239500 0 239556 200
rect 242200 0 242256 200
rect 244900 0 244956 200
rect 247600 0 247656 200
rect 250300 0 250356 200
rect 253000 0 253056 200
rect 255700 0 255756 200
<< metal4 >>
rect 3049 0 6899 400
rect 7229 0 11079 400
rect 12049 0 15899 400
rect 282049 0 285899 400
rect 286229 0 290079 400
<< labels >>
rlabel metal3 s 291760 1781 292400 1837 4 gpio_analog[6]
port 1 nsew
rlabel metal3 s 291760 2372 292400 2428 4 gpio_noesd[6]
port 2 nsew
rlabel metal3 s 291150 48992 292000 51492 4 io_analog[0]
port 3 nsew
rlabel metal3 s 283297 61150 285797 62000 4 io_analog[1]
port 4 nsew
rlabel metal3 s 232697 61150 235197 62000 4 io_analog[2]
port 5 nsew
rlabel metal3 s 206697 61150 209197 62000 4 io_analog[3]
port 6 nsew
rlabel metal3 s 159497 61150 161997 62000 4 io_analog[4]
port 7 nsew
rlabel metal3 s 163397 61150 164497 62000 4 io_clamp_high[0]
port 8 nsew
rlabel metal3 s 162147 61150 163247 62000 4 io_clamp_low[0]
port 9 nsew
rlabel metal3 s 291760 3554 292400 3610 4 io_in[13]
port 10 nsew
rlabel metal3 s 291760 2963 292400 3019 4 io_in_3v3[13]
port 11 nsew
rlabel metal3 s 291760 4736 292400 4792 4 io_oeb[13]
port 12 nsew
rlabel metal3 s 291760 4145 292400 4201 4 io_out[13]
port 13 nsew
rlabel metal3 s 291170 24892 292000 27292 4 vccd1
port 14 nsew
rlabel metal3 s 255297 61170 257697 62000 4 vssa1
port 15 nsew
rlabel metal3 s 86697 61150 87797 62000 4 io_clamp_high[2]
port 16 nsew
rlabel metal3 s 108647 61150 111147 62000 4 io_analog[5]
port 17 nsew
rlabel metal3 s 111297 61150 112397 62000 4 io_clamp_low[1]
port 18 nsew
rlabel metal3 s 85447 61150 86547 62000 4 io_clamp_low[2]
port 19 nsew
rlabel metal3 s 82797 61150 85297 62000 4 io_analog[6]
port 20 nsew
rlabel metal3 s 60097 61150 62597 62000 4 io_analog[7]
port 21 nsew
rlabel metal3 s 34097 61150 36597 62000 4 io_analog[8]
port 22 nsew
rlabel metal3 s 8097 61150 10597 62000 4 io_analog[9]
port 23 nsew
rlabel metal3 s 0 50121 850 52621 4 io_analog[10]
port 24 nsew
rlabel metal3 s 0 26921 830 29321 4 vccd2
port 25 nsew
rlabel metal3 s 112547 61150 113647 62000 4 io_clamp_high[1]
port 26 nsew
rlabel metal3 s 80200 0 80256 200 4 analog_la_out[26]
port 27 nsew
rlabel metal3 s 82900 0 82956 200 4 analog_la_out[27]
port 28 nsew
rlabel metal3 s 85600 0 85656 200 4 analog_la_out[28]
port 29 nsew
rlabel metal3 s 88300 0 88356 200 4 analog_la_out[29]
port 30 nsew
rlabel metal3 s 91000 0 91056 200 4 analog_la_in[0]
port 31 nsew
rlabel metal3 s 93700 0 93756 200 4 analog_la_in[1]
port 32 nsew
rlabel metal3 s 96400 0 96456 200 4 analog_la_in[2]
port 33 nsew
rlabel metal3 s 99100 0 99156 200 4 analog_la_in[3]
port 34 nsew
rlabel metal3 s 101800 0 101856 200 4 analog_la_in[4]
port 35 nsew
rlabel metal3 s 104500 0 104556 200 4 analog_la_in[5]
port 36 nsew
rlabel metal3 s 107200 0 107256 200 4 analog_la_in[6]
port 37 nsew
rlabel metal3 s 109900 0 109956 200 4 analog_la_in[7]
port 38 nsew
rlabel metal3 s 112600 0 112656 200 4 analog_la_in[8]
port 39 nsew
rlabel metal3 s 115300 0 115356 200 4 analog_la_in[9]
port 40 nsew
rlabel metal3 s 118000 0 118056 200 4 analog_la_in[10]
port 41 nsew
rlabel metal3 s 120700 0 120756 200 4 analog_la_in[11]
port 42 nsew
rlabel metal3 s 123400 0 123456 200 4 analog_la_in[12]
port 43 nsew
rlabel metal3 s 126100 0 126156 200 4 analog_la_in[13]
port 44 nsew
rlabel metal3 s 128800 0 128856 200 4 analog_la_in[14]
port 45 nsew
rlabel metal3 s 131500 0 131556 200 4 analog_la_in[15]
port 46 nsew
rlabel metal3 s 134200 0 134256 200 4 analog_la_in[16]
port 47 nsew
rlabel metal3 s 136900 0 136956 200 4 analog_la_in[17]
port 48 nsew
rlabel metal3 s 139600 0 139656 200 4 analog_la_in[18]
port 49 nsew
rlabel metal3 s 142300 0 142356 200 4 analog_la_in[19]
port 50 nsew
rlabel metal3 s 145000 0 145056 200 4 analog_la_in[20]
port 51 nsew
rlabel metal3 s 10000 0 10056 200 4 analog_la_out[0]
port 52 nsew
rlabel metal3 s 12700 0 12756 200 4 analog_la_out[1]
port 53 nsew
rlabel metal3 s 15400 0 15456 200 4 analog_la_out[2]
port 54 nsew
rlabel metal3 s 18100 0 18156 200 4 analog_la_out[3]
port 55 nsew
rlabel metal3 s 20800 0 20856 200 4 analog_la_out[4]
port 56 nsew
rlabel metal3 s 23500 0 23556 200 4 analog_la_out[5]
port 57 nsew
rlabel metal3 s 26200 0 26256 200 4 analog_la_out[6]
port 58 nsew
rlabel metal3 s 28900 0 28956 200 4 analog_la_out[7]
port 59 nsew
rlabel metal3 s 31600 0 31656 200 4 analog_la_out[8]
port 60 nsew
rlabel metal3 s 34300 0 34356 200 4 analog_la_out[9]
port 61 nsew
rlabel metal3 s 37000 0 37056 200 4 analog_la_out[10]
port 62 nsew
rlabel metal3 s 39700 0 39756 200 4 analog_la_out[11]
port 63 nsew
rlabel metal3 s 42400 0 42456 200 4 analog_la_out[12]
port 64 nsew
rlabel metal3 s 45100 0 45156 200 4 analog_la_out[13]
port 65 nsew
rlabel metal3 s 47800 0 47856 200 4 analog_la_out[14]
port 66 nsew
rlabel metal3 s 50500 0 50556 200 4 analog_la_out[15]
port 67 nsew
rlabel metal3 s 53200 0 53256 200 4 analog_la_out[16]
port 68 nsew
rlabel metal3 s 55900 0 55956 200 4 analog_la_out[17]
port 69 nsew
rlabel metal3 s 58600 0 58656 200 4 analog_la_out[18]
port 70 nsew
rlabel metal3 s 61300 0 61356 200 4 analog_la_out[19]
port 71 nsew
rlabel metal3 s 64000 0 64056 200 4 analog_la_out[20]
port 72 nsew
rlabel metal3 s 66700 0 66756 200 4 analog_la_out[21]
port 73 nsew
rlabel metal3 s 69400 0 69456 200 4 analog_la_out[22]
port 74 nsew
rlabel metal3 s 72100 0 72156 200 4 analog_la_out[23]
port 75 nsew
rlabel metal3 s 74800 0 74856 200 4 analog_la_out[24]
port 76 nsew
rlabel metal3 s 77500 0 77556 200 4 analog_la_out[25]
port 77 nsew
rlabel metal3 s 223300 0 223356 200 4 ctln[7]
port 78 nsew
rlabel metal3 s 226000 0 226056 200 4 ctln[8]
port 79 nsew
rlabel metal3 s 228700 0 228756 200 4 ctln[9]
port 80 nsew
rlabel metal3 s 231400 0 231456 200 4 trim[0]
port 81 nsew
rlabel metal3 s 234100 0 234156 200 4 trim[1]
port 82 nsew
rlabel metal3 s 236800 0 236856 200 4 trim[2]
port 83 nsew
rlabel metal3 s 239500 0 239556 200 4 trim[3]
port 84 nsew
rlabel metal3 s 242200 0 242256 200 4 trim[4]
port 85 nsew
rlabel metal3 s 244900 0 244956 200 4 trimb[0]
port 86 nsew
rlabel metal3 s 247600 0 247656 200 4 trimb[1]
port 87 nsew
rlabel metal3 s 250300 0 250356 200 4 trimb[2]
port 88 nsew
rlabel metal3 s 253000 0 253056 200 4 trimb[3]
port 89 nsew
rlabel metal3 s 255700 0 255756 200 4 trimb[4]
port 90 nsew
rlabel metal3 s 147700 0 147756 200 4 analog_la_in[21]
port 91 nsew
rlabel metal3 s 150400 0 150456 200 4 analog_la_in[22]
port 92 nsew
rlabel metal3 s 153100 0 153156 200 4 analog_la_in[23]
port 93 nsew
rlabel metal3 s 155800 0 155856 200 4 analog_la_in[24]
port 94 nsew
rlabel metal3 s 158500 0 158556 200 4 analog_la_in[25]
port 95 nsew
rlabel metal3 s 161200 0 161256 200 4 analog_la_in[26]
port 96 nsew
rlabel metal3 s 163900 0 163956 200 4 analog_la_in[27]
port 97 nsew
rlabel metal3 s 166600 0 166656 200 4 analog_la_in[28]
port 98 nsew
rlabel metal3 s 174700 0 174756 200 4 analog_la_in[29]
port 99 nsew
rlabel metal3 s 177400 0 177456 200 4 ctlp[0]
port 100 nsew
rlabel metal3 s 180100 0 180156 200 4 ctlp[1]
port 101 nsew
rlabel metal3 s 182800 0 182856 200 4 ctlp[2]
port 102 nsew
rlabel metal3 s 185500 0 185556 200 4 ctlp[3]
port 103 nsew
rlabel metal3 s 188200 0 188256 200 4 ctlp[4]
port 104 nsew
rlabel metal3 s 190900 0 190956 200 4 ctlp[5]
port 105 nsew
rlabel metal3 s 193600 0 193656 200 4 ctlp[6]
port 106 nsew
rlabel metal3 s 196300 0 196356 200 4 ctlp[7]
port 107 nsew
rlabel metal3 s 199000 0 199056 200 4 ctlp[8]
port 108 nsew
rlabel metal3 s 201700 0 201756 200 4 ctlp[9]
port 109 nsew
rlabel metal3 s 204400 0 204456 200 4 ctln[0]
port 110 nsew
rlabel metal3 s 207100 0 207156 200 4 ctln[1]
port 111 nsew
rlabel metal3 s 209800 0 209856 200 4 ctln[2]
port 112 nsew
rlabel metal3 s 212500 0 212556 200 4 ctln[3]
port 113 nsew
rlabel metal3 s 215200 0 215256 200 4 ctln[4]
port 114 nsew
rlabel metal3 s 217900 0 217956 200 4 ctln[5]
port 115 nsew
rlabel metal3 s 220600 0 220656 200 4 ctln[6]
port 116 nsew
rlabel metal4 s 286229 0 290079 400 4 vssa1
port 15 nsew
rlabel metal4 s 3049 0 6899 400 4 vdda2
port 117 nsew
rlabel metal4 s 7229 0 11079 400 4 vssd2
port 118 nsew
rlabel metal4 s 12049 0 15899 400 4 vssa2
port 119 nsew
rlabel metal4 s 282049 0 285899 400 4 vdda1
port 120 nsew
<< properties >>
string FIXED_BBOX 0 0 292000 62000
string path 2557.280 0.000 2557.280 2.000 
<< end >>
