magic
tech sky130B
timestamp 1659316836
<< metal1 >>
rect -1200 7650 8500 7700
rect -1200 -1950 -1150 7650
rect -650 7100 7950 7150
rect -650 6700 -100 7100
rect -650 6600 0 6700
rect 100 6600 400 7100
rect -650 6400 -600 6600
rect -200 6500 400 6600
rect -100 6400 400 6500
rect -650 6200 400 6400
rect -650 6100 500 6200
rect 600 6100 900 7100
rect -650 5900 -600 6100
rect 300 6000 900 6100
rect 400 5900 900 6000
rect -650 5700 900 5900
rect -650 5600 1000 5700
rect 1100 5600 1400 7100
rect -650 5400 -600 5600
rect 800 5500 1400 5600
rect 900 5400 1400 5500
rect -650 5200 1400 5400
rect -650 5100 1500 5200
rect 1600 5100 1900 7100
rect -650 4900 -600 5100
rect 1300 5000 1900 5100
rect 1400 4900 1900 5000
rect -650 4700 1900 4900
rect -650 4600 2000 4700
rect 2100 4600 2400 7100
rect -650 4400 -600 4600
rect 1800 4500 2400 4600
rect 1900 4400 2400 4500
rect -650 4200 2400 4400
rect -650 4100 2500 4200
rect 2600 4100 2900 7100
rect -650 3900 -600 4100
rect 2300 4000 2900 4100
rect 2400 3900 2900 4000
rect -650 3700 2900 3900
rect 3100 3700 3400 7100
rect 3600 4100 3900 7100
rect 4100 4600 4400 7100
rect 4600 5100 4900 7100
rect 5100 5600 5400 7100
rect 5600 6100 5900 7100
rect 6100 6600 6400 7100
rect 6600 7000 7200 7100
rect 6600 6900 7100 7000
rect 7900 6900 7950 7100
rect 6600 6700 7950 6900
rect 6500 6600 7950 6700
rect 6100 6500 6700 6600
rect 6100 6400 6600 6500
rect 7900 6400 7950 6600
rect 6100 6200 7950 6400
rect 6000 6100 7950 6200
rect 5600 6000 6200 6100
rect 5600 5900 6100 6000
rect 7900 5900 7950 6100
rect 5600 5700 7950 5900
rect 5500 5600 7950 5700
rect 5100 5500 5700 5600
rect 5100 5400 5600 5500
rect 7900 5400 7950 5600
rect 5100 5200 7950 5400
rect 5000 5100 7950 5200
rect 4600 5000 5200 5100
rect 4600 4900 5100 5000
rect 7900 4900 7950 5100
rect 4600 4700 7950 4900
rect 4500 4600 7950 4700
rect 4100 4500 4700 4600
rect 4100 4400 4600 4500
rect 7900 4400 7950 4600
rect 4100 4200 7950 4400
rect 4000 4100 7950 4200
rect 3600 4000 4200 4100
rect 3600 3900 4100 4000
rect 7900 3900 7950 4100
rect 3600 3700 7950 3900
rect -650 3650 7950 3700
rect 8450 3650 8500 7650
rect -650 3600 8500 3650
rect -650 3400 -600 3600
rect 2800 3400 3700 3600
rect -650 3100 3000 3400
rect -650 2900 -600 3100
rect 2800 2900 3000 3100
rect 3600 3100 7500 3400
rect 3600 2900 3700 3100
rect -650 2850 8500 2900
rect -650 2800 7950 2850
rect -650 2600 2900 2800
rect -650 2400 -600 2600
rect 2400 2500 2900 2600
rect 2300 2400 2900 2500
rect -650 2300 2500 2400
rect -650 2100 2400 2300
rect -650 1900 -600 2100
rect 1900 2000 2400 2100
rect 1800 1900 2400 2000
rect -650 1800 2000 1900
rect -650 1600 1900 1800
rect -650 1400 -600 1600
rect 1400 1500 1900 1600
rect 1300 1400 1900 1500
rect -650 1300 1500 1400
rect -650 1100 1400 1300
rect -650 900 -600 1100
rect 900 1000 1400 1100
rect 800 900 1400 1000
rect -650 800 1000 900
rect -650 600 900 800
rect -650 400 -600 600
rect 400 500 900 600
rect 300 400 900 500
rect -650 300 500 400
rect -650 100 400 300
rect -650 -100 -600 100
rect -100 0 400 100
rect -200 -100 400 0
rect -650 -200 0 -100
rect -650 -600 -100 -200
rect -650 -700 -500 -600
rect -650 -1400 -600 -700
rect -400 -1400 -100 -600
rect 100 -1400 400 -100
rect 600 -1400 900 400
rect 1100 -1400 1400 900
rect 1600 -1400 1900 1400
rect 2100 -1400 2400 1900
rect 2600 -1400 2900 2400
rect 3100 -1400 3400 2800
rect 3600 2600 7950 2800
rect 3600 2500 4100 2600
rect 3600 2400 4200 2500
rect 7900 2400 7950 2600
rect 3600 -1400 3900 2400
rect 4000 2300 7950 2400
rect 4100 2100 7950 2300
rect 4100 2000 4600 2100
rect 4100 1900 4700 2000
rect 7900 1900 7950 2100
rect 4100 -1400 4400 1900
rect 4500 1800 7950 1900
rect 4600 1600 7950 1800
rect 4600 1500 5100 1600
rect 4600 1400 5200 1500
rect 7900 1400 7950 1600
rect 4600 -1400 4900 1400
rect 5000 1300 7950 1400
rect 5100 1100 7950 1300
rect 5100 1000 5600 1100
rect 5100 900 5700 1000
rect 7900 900 7950 1100
rect 5100 -1400 5400 900
rect 5500 800 7950 900
rect 5600 600 7950 800
rect 5600 500 6100 600
rect 5600 400 6200 500
rect 7900 400 7950 600
rect 5600 -1400 5900 400
rect 6000 300 7950 400
rect 6100 100 7950 300
rect 6100 0 6600 100
rect 6100 -100 6700 0
rect 7900 -100 7950 100
rect 6100 -1400 6400 -100
rect 6500 -200 7950 -100
rect 6600 -400 7950 -200
rect 6600 -500 7100 -400
rect 6600 -600 7200 -500
rect 7900 -600 7950 -400
rect 6600 -1400 6900 -600
rect 7000 -700 7950 -600
rect 7100 -900 7950 -700
rect 7100 -1000 7600 -900
rect 7100 -1100 7700 -1000
rect 7100 -1400 7400 -1100
rect 7500 -1200 7800 -1100
rect 7900 -1200 7950 -900
rect 7600 -1300 7950 -1200
rect 7700 -1400 7950 -1300
rect -650 -1450 7950 -1400
rect 8450 -1950 8500 2850
rect -1200 -2000 8500 -1950
<< via1 >>
rect -1150 7150 8450 7650
rect -1150 -1450 -650 7150
rect 7950 3650 8450 7150
rect 3000 2900 3600 3400
rect 7950 -1450 8450 2850
rect -1150 -1950 8450 -1450
<< metal2 >>
rect -1200 7650 8500 7700
rect -1200 -1950 -1150 7650
rect -650 7100 7950 7150
rect -650 6700 -100 7100
rect -650 6600 0 6700
rect 100 6600 400 7100
rect -650 6400 -600 6600
rect -200 6500 400 6600
rect -100 6400 400 6500
rect -650 6200 400 6400
rect -650 6100 500 6200
rect 600 6100 900 7100
rect -650 5900 -600 6100
rect 300 6000 900 6100
rect 400 5900 900 6000
rect -650 5700 900 5900
rect -650 5600 1000 5700
rect 1100 5600 1400 7100
rect -650 5400 -600 5600
rect 800 5500 1400 5600
rect 900 5400 1400 5500
rect -650 5200 1400 5400
rect -650 5100 1500 5200
rect 1600 5100 1900 7100
rect -650 4900 -600 5100
rect 1300 5000 1900 5100
rect 1400 4900 1900 5000
rect -650 4700 1900 4900
rect -650 4600 2000 4700
rect 2100 4600 2400 7100
rect -650 4400 -600 4600
rect 1800 4500 2400 4600
rect 1900 4400 2400 4500
rect -650 4200 2400 4400
rect -650 4100 2500 4200
rect 2600 4100 2900 7100
rect -650 3900 -600 4100
rect 2300 4000 2900 4100
rect 2400 3900 2900 4000
rect -650 3700 2900 3900
rect 3100 3700 3400 7100
rect 3600 4100 3900 7100
rect 4100 4600 4400 7100
rect 4600 5100 4900 7100
rect 5100 5600 5400 7100
rect 5600 6100 5900 7100
rect 6100 6600 6400 7100
rect 6600 7000 7200 7100
rect 6600 6900 7100 7000
rect 7900 6900 7950 7100
rect 6600 6700 7950 6900
rect 6500 6600 7950 6700
rect 6100 6500 6700 6600
rect 6100 6400 6600 6500
rect 7900 6400 7950 6600
rect 6100 6200 7950 6400
rect 6000 6100 7950 6200
rect 5600 6000 6200 6100
rect 5600 5900 6100 6000
rect 7900 5900 7950 6100
rect 5600 5700 7950 5900
rect 5500 5600 7950 5700
rect 5100 5500 5700 5600
rect 5100 5400 5600 5500
rect 7900 5400 7950 5600
rect 5100 5200 7950 5400
rect 5000 5100 7950 5200
rect 4600 5000 5200 5100
rect 4600 4900 5100 5000
rect 7900 4900 7950 5100
rect 4600 4700 7950 4900
rect 4500 4600 7950 4700
rect 4100 4500 4700 4600
rect 4100 4400 4600 4500
rect 7900 4400 7950 4600
rect 4100 4200 7950 4400
rect 4000 4100 7950 4200
rect 3600 4000 4200 4100
rect 3600 3900 4100 4000
rect 7900 3900 7950 4100
rect 3600 3700 7950 3900
rect -650 3650 7950 3700
rect 8450 3650 8500 7650
rect -650 3600 8500 3650
rect -650 3400 -600 3600
rect 2800 3400 3700 3600
rect -650 3100 3000 3400
rect -650 2900 -600 3100
rect 2800 2900 3000 3100
rect 3600 3100 7500 3400
rect 3600 2900 3700 3100
rect -650 2850 8500 2900
rect -650 2800 7950 2850
rect -650 2600 2900 2800
rect -650 2400 -600 2600
rect 2400 2500 2900 2600
rect 2300 2400 2900 2500
rect -650 2300 2500 2400
rect -650 2100 2400 2300
rect -650 1900 -600 2100
rect 1900 2000 2400 2100
rect 1800 1900 2400 2000
rect -650 1800 2000 1900
rect -650 1600 1900 1800
rect -650 1400 -600 1600
rect 1400 1500 1900 1600
rect 1300 1400 1900 1500
rect -650 1300 1500 1400
rect -650 1100 1400 1300
rect -650 900 -600 1100
rect 900 1000 1400 1100
rect 800 900 1400 1000
rect -650 800 1000 900
rect -650 600 900 800
rect -650 400 -600 600
rect 400 500 900 600
rect 300 400 900 500
rect -650 300 500 400
rect -650 100 400 300
rect -650 -100 -600 100
rect -100 0 400 100
rect -200 -100 400 0
rect -650 -200 0 -100
rect -650 -600 -100 -200
rect -650 -700 -500 -600
rect -650 -1400 -600 -700
rect -400 -1400 -100 -600
rect 100 -1400 400 -100
rect 600 -1400 900 400
rect 1100 -1400 1400 900
rect 1600 -1400 1900 1400
rect 2100 -1400 2400 1900
rect 2600 -1400 2900 2400
rect 3100 -1400 3400 2800
rect 3600 2600 7950 2800
rect 3600 2500 4100 2600
rect 3600 2400 4200 2500
rect 7900 2400 7950 2600
rect 3600 -1400 3900 2400
rect 4000 2300 7950 2400
rect 4100 2100 7950 2300
rect 4100 2000 4600 2100
rect 4100 1900 4700 2000
rect 7900 1900 7950 2100
rect 4100 -1400 4400 1900
rect 4500 1800 7950 1900
rect 4600 1600 7950 1800
rect 4600 1500 5100 1600
rect 4600 1400 5200 1500
rect 7900 1400 7950 1600
rect 4600 -1400 4900 1400
rect 5000 1300 7950 1400
rect 5100 1100 7950 1300
rect 5100 1000 5600 1100
rect 5100 900 5700 1000
rect 7900 900 7950 1100
rect 5100 -1400 5400 900
rect 5500 800 7950 900
rect 5600 600 7950 800
rect 5600 500 6100 600
rect 5600 400 6200 500
rect 7900 400 7950 600
rect 5600 -1400 5900 400
rect 6000 300 7950 400
rect 6100 100 7950 300
rect 6100 0 6600 100
rect 6100 -100 6700 0
rect 7900 -100 7950 100
rect 6100 -1400 6400 -100
rect 6500 -200 7950 -100
rect 6600 -400 7950 -200
rect 6600 -500 7100 -400
rect 6600 -600 7200 -500
rect 7900 -600 7950 -400
rect 6600 -1400 6900 -600
rect 7000 -700 7950 -600
rect 7100 -900 7950 -700
rect 7100 -1000 7600 -900
rect 7100 -1100 7700 -1000
rect 7100 -1400 7400 -1100
rect 7500 -1200 7800 -1100
rect 7900 -1200 7950 -900
rect 7600 -1300 7950 -1200
rect 7700 -1400 7950 -1300
rect -650 -1450 7950 -1400
rect 8450 -1950 8500 2850
rect -1200 -2000 8500 -1950
<< via2 >>
rect -1150 7150 8450 7650
rect -1150 -1450 -650 7150
rect 7950 3650 8450 7150
rect 3000 2900 3600 3400
rect 7950 -1450 8450 2850
rect -1150 -1950 8450 -1450
<< metal3 >>
rect -1200 7650 8500 7700
rect -1200 -1950 -1150 7650
rect -650 7100 7950 7150
rect -650 6700 -100 7100
rect -650 6600 0 6700
rect 100 6600 400 7100
rect -650 6400 -600 6600
rect -200 6500 400 6600
rect -100 6400 400 6500
rect -650 6200 400 6400
rect -650 6100 500 6200
rect 600 6100 900 7100
rect -650 5900 -600 6100
rect 300 6000 900 6100
rect 400 5900 900 6000
rect -650 5700 900 5900
rect -650 5600 1000 5700
rect 1100 5600 1400 7100
rect -650 5400 -600 5600
rect 800 5500 1400 5600
rect 900 5400 1400 5500
rect -650 5200 1400 5400
rect -650 5100 1500 5200
rect 1600 5100 1900 7100
rect -650 4900 -600 5100
rect 1300 5000 1900 5100
rect 1400 4900 1900 5000
rect -650 4700 1900 4900
rect -650 4600 2000 4700
rect 2100 4600 2400 7100
rect -650 4400 -600 4600
rect 1800 4500 2400 4600
rect 1900 4400 2400 4500
rect -650 4200 2400 4400
rect -650 4100 2500 4200
rect 2600 4100 2900 7100
rect -650 3900 -600 4100
rect 2300 4000 2900 4100
rect 2400 3900 2900 4000
rect -650 3700 2900 3900
rect 3100 3700 3400 7100
rect 3600 4100 3900 7100
rect 4100 4600 4400 7100
rect 4600 5100 4900 7100
rect 5100 5600 5400 7100
rect 5600 6100 5900 7100
rect 6100 6600 6400 7100
rect 6600 7000 7200 7100
rect 6600 6900 7100 7000
rect 7900 6900 7950 7100
rect 6600 6700 7950 6900
rect 6500 6600 7950 6700
rect 6100 6500 6700 6600
rect 6100 6400 6600 6500
rect 7900 6400 7950 6600
rect 6100 6200 7950 6400
rect 6000 6100 7950 6200
rect 5600 6000 6200 6100
rect 5600 5900 6100 6000
rect 7900 5900 7950 6100
rect 5600 5700 7950 5900
rect 5500 5600 7950 5700
rect 5100 5500 5700 5600
rect 5100 5400 5600 5500
rect 7900 5400 7950 5600
rect 5100 5200 7950 5400
rect 5000 5100 7950 5200
rect 4600 5000 5200 5100
rect 4600 4900 5100 5000
rect 7900 4900 7950 5100
rect 4600 4700 7950 4900
rect 4500 4600 7950 4700
rect 4100 4500 4700 4600
rect 4100 4400 4600 4500
rect 7900 4400 7950 4600
rect 4100 4200 7950 4400
rect 4000 4100 7950 4200
rect 3600 4000 4200 4100
rect 3600 3900 4100 4000
rect 7900 3900 7950 4100
rect 3600 3700 7950 3900
rect -650 3650 7950 3700
rect 8450 3650 8500 7650
rect -650 3600 8500 3650
rect -650 3400 -600 3600
rect 2800 3400 3700 3600
rect -650 3100 3000 3400
rect -650 2900 -600 3100
rect 2800 2900 3000 3100
rect 3600 3100 7500 3400
rect 3600 2900 3700 3100
rect -650 2850 8500 2900
rect -650 2800 7950 2850
rect -650 2600 2900 2800
rect -650 2400 -600 2600
rect 2400 2500 2900 2600
rect 2300 2400 2900 2500
rect -650 2300 2500 2400
rect -650 2100 2400 2300
rect -650 1900 -600 2100
rect 1900 2000 2400 2100
rect 1800 1900 2400 2000
rect -650 1800 2000 1900
rect -650 1600 1900 1800
rect -650 1400 -600 1600
rect 1400 1500 1900 1600
rect 1300 1400 1900 1500
rect -650 1300 1500 1400
rect -650 1100 1400 1300
rect -650 900 -600 1100
rect 900 1000 1400 1100
rect 800 900 1400 1000
rect -650 800 1000 900
rect -650 600 900 800
rect -650 400 -600 600
rect 400 500 900 600
rect 300 400 900 500
rect -650 300 500 400
rect -650 100 400 300
rect -650 -100 -600 100
rect -100 0 400 100
rect -200 -100 400 0
rect -650 -200 0 -100
rect -650 -600 -100 -200
rect -650 -700 -500 -600
rect -650 -1400 -600 -700
rect -400 -1400 -100 -600
rect 100 -1400 400 -100
rect 600 -1400 900 400
rect 1100 -1400 1400 900
rect 1600 -1400 1900 1400
rect 2100 -1400 2400 1900
rect 2600 -1400 2900 2400
rect 3100 -1400 3400 2800
rect 3600 2600 7950 2800
rect 3600 2500 4100 2600
rect 3600 2400 4200 2500
rect 7900 2400 7950 2600
rect 3600 -1400 3900 2400
rect 4000 2300 7950 2400
rect 4100 2100 7950 2300
rect 4100 2000 4600 2100
rect 4100 1900 4700 2000
rect 7900 1900 7950 2100
rect 4100 -1400 4400 1900
rect 4500 1800 7950 1900
rect 4600 1600 7950 1800
rect 4600 1500 5100 1600
rect 4600 1400 5200 1500
rect 7900 1400 7950 1600
rect 4600 -1400 4900 1400
rect 5000 1300 7950 1400
rect 5100 1100 7950 1300
rect 5100 1000 5600 1100
rect 5100 900 5700 1000
rect 7900 900 7950 1100
rect 5100 -1400 5400 900
rect 5500 800 7950 900
rect 5600 600 7950 800
rect 5600 500 6100 600
rect 5600 400 6200 500
rect 7900 400 7950 600
rect 5600 -1400 5900 400
rect 6000 300 7950 400
rect 6100 100 7950 300
rect 6100 0 6600 100
rect 6100 -100 6700 0
rect 7900 -100 7950 100
rect 6100 -1400 6400 -100
rect 6500 -200 7950 -100
rect 6600 -400 7950 -200
rect 6600 -500 7100 -400
rect 6600 -600 7200 -500
rect 7900 -600 7950 -400
rect 6600 -1400 6900 -600
rect 7000 -700 7950 -600
rect 7100 -900 7950 -700
rect 7100 -1000 7600 -900
rect 7100 -1100 7700 -1000
rect 7100 -1400 7400 -1100
rect 7500 -1200 7800 -1100
rect 7900 -1200 7950 -900
rect 7600 -1300 7950 -1200
rect 7700 -1400 7950 -1300
rect -650 -1450 7950 -1400
rect 8450 -1950 8500 2850
rect -1200 -2000 8500 -1950
<< via3 >>
rect -1150 7150 8450 7650
rect -1150 -1450 -650 7150
rect 7950 3650 8450 7150
rect 3000 2900 3600 3400
rect 7950 -1450 8450 2850
rect -1150 -1950 8450 -1450
<< metal4 >>
rect -1200 7650 8500 7700
rect -1200 -1950 -1150 7650
rect -650 7100 7950 7150
rect -650 -1400 -600 7100
rect 7900 3650 7950 7100
rect 8450 3650 8500 7650
rect 7900 3600 8500 3650
rect 6800 3550 7650 3600
rect 2900 3400 3700 3500
rect 2900 2900 3000 3400
rect 3600 2900 3700 3400
rect 6800 2950 6850 3550
rect 7450 3500 7650 3550
rect 7450 3000 8700 3500
rect 7450 2950 7650 3000
rect 6800 2900 7650 2950
rect 2900 2800 3700 2900
rect 7900 2850 8500 2900
rect 7900 -1400 7950 2850
rect -650 -1450 7950 -1400
rect 8450 -1950 8500 2850
rect -1200 -2000 8500 -1950
<< via4 >>
rect 3000 2900 3600 3400
rect 6850 2950 7450 3550
<< metal5 >>
rect 0 6000 6500 6500
rect 0 -300 500 6000
rect 800 5200 5700 5700
rect 800 500 1300 5200
rect 1600 4400 4900 4900
rect 1600 1300 2100 4400
rect 2400 3400 3700 3500
rect 2400 2900 3000 3400
rect 3600 2900 3700 3400
rect 2400 2800 3700 2900
rect 2400 2100 2900 2800
rect 4400 2100 4900 4400
rect 2400 1600 4900 2100
rect 5200 1300 5700 5200
rect 1600 800 5700 1300
rect 6000 500 6500 6000
rect 800 0 6500 500
rect 6800 3550 7500 3600
rect 6800 2950 6850 3550
rect 7450 2950 7500 3550
rect 6800 2900 7500 2950
rect 6800 2850 7450 2900
rect 6800 2800 7400 2850
rect 6800 2750 7350 2800
rect 6800 -300 7300 2750
rect 0 -800 7300 -300
<< end >>
