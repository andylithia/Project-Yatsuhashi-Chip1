magic
tech sky130A
magscale 1 2
timestamp 1664325575
<< viali >>
rect 236 6432 4959 6470
rect 46 236 84 6280
rect 5054 236 5092 6280
rect 236 46 4902 84
<< metal1 >>
rect 30 6470 5110 6480
rect 30 6432 236 6470
rect 4959 6432 5110 6470
rect 30 6422 5110 6432
rect 30 6420 100 6422
rect 5040 6420 5110 6422
rect 232 6290 252 6390
rect 4886 6290 4906 6390
rect 165 6238 235 6258
rect 165 258 235 278
rect 323 6238 393 6258
rect 323 258 393 278
rect 481 6238 551 6258
rect 481 258 551 278
rect 639 6238 709 6258
rect 639 258 709 278
rect 797 6238 867 6258
rect 797 258 867 278
rect 955 6238 1025 6258
rect 955 258 1025 278
rect 1113 6238 1183 6258
rect 1113 258 1183 278
rect 1271 6238 1341 6258
rect 1271 258 1341 278
rect 1429 6238 1499 6258
rect 1429 258 1499 278
rect 1587 6238 1657 6258
rect 1587 258 1657 278
rect 1745 6238 1815 6258
rect 1745 258 1815 278
rect 1903 6238 1973 6258
rect 1903 258 1973 278
rect 2061 6238 2131 6258
rect 2061 258 2131 278
rect 2219 6238 2289 6258
rect 2219 258 2289 278
rect 2377 6238 2447 6258
rect 2377 258 2447 278
rect 2535 6238 2605 6258
rect 2535 258 2605 278
rect 2693 6238 2763 6258
rect 2693 258 2763 278
rect 2851 6238 2921 6258
rect 2851 258 2921 278
rect 3009 6238 3079 6258
rect 3009 258 3079 278
rect 3167 6238 3237 6258
rect 3167 258 3237 278
rect 3325 6238 3395 6258
rect 3325 258 3395 278
rect 3483 6238 3553 6258
rect 3483 258 3553 278
rect 3641 6238 3711 6258
rect 3641 258 3711 278
rect 3799 6238 3869 6258
rect 3799 258 3869 278
rect 3957 6238 4027 6258
rect 3957 258 4027 278
rect 4115 6238 4185 6258
rect 4115 258 4185 278
rect 4273 6238 4343 6258
rect 4273 258 4343 278
rect 4431 6238 4501 6258
rect 4431 258 4501 278
rect 4589 6238 4659 6258
rect 4589 258 4659 278
rect 4747 6238 4817 6258
rect 4747 258 4817 278
rect 4905 6238 4975 6258
rect 4905 258 4975 278
rect 232 126 252 226
rect 4886 126 4906 226
rect 30 94 100 100
rect 5040 94 5110 100
rect 30 84 5110 94
rect 30 46 236 84
rect 4902 46 5110 84
rect 30 30 5110 46
<< via1 >>
rect 30 6280 100 6420
rect 252 6290 4886 6390
rect 30 236 46 6280
rect 46 236 84 6280
rect 84 236 100 6280
rect 5040 6280 5110 6420
rect 165 278 235 6238
rect 323 278 393 6238
rect 481 278 551 6238
rect 639 278 709 6238
rect 797 278 867 6238
rect 955 278 1025 6238
rect 1113 278 1183 6238
rect 1271 278 1341 6238
rect 1429 278 1499 6238
rect 1587 278 1657 6238
rect 1745 278 1815 6238
rect 1903 278 1973 6238
rect 2061 278 2131 6238
rect 2219 278 2289 6238
rect 2377 278 2447 6238
rect 2535 278 2605 6238
rect 2693 278 2763 6238
rect 2851 278 2921 6238
rect 3009 278 3079 6238
rect 3167 278 3237 6238
rect 3325 278 3395 6238
rect 3483 278 3553 6238
rect 3641 278 3711 6238
rect 3799 278 3869 6238
rect 3957 278 4027 6238
rect 4115 278 4185 6238
rect 4273 278 4343 6238
rect 4431 278 4501 6238
rect 4589 278 4659 6238
rect 4747 278 4817 6238
rect 4905 278 4975 6238
rect 30 100 100 236
rect 5040 236 5054 6280
rect 5054 236 5092 6280
rect 5092 236 5110 6280
rect 252 126 4886 226
rect 5040 100 5110 236
<< metal2 >>
rect 30 6420 100 6480
rect 5040 6420 5110 6480
rect 232 6380 252 6390
rect 4886 6380 4906 6390
rect 232 6310 240 6380
rect 4900 6310 4906 6380
rect 232 6290 252 6310
rect 4886 6290 4906 6310
rect 165 6238 235 6258
rect 165 258 235 278
rect 323 6238 393 6258
rect 323 258 393 278
rect 481 6238 551 6258
rect 481 258 551 278
rect 639 6238 709 6258
rect 639 258 709 278
rect 797 6238 867 6258
rect 797 258 867 278
rect 955 6238 1025 6258
rect 955 258 1025 278
rect 1113 6238 1183 6258
rect 1113 258 1183 278
rect 1271 6238 1341 6258
rect 1271 258 1341 278
rect 1429 6238 1499 6258
rect 1429 258 1499 278
rect 1587 6238 1657 6258
rect 1587 258 1657 278
rect 1745 6238 1815 6258
rect 1745 258 1815 278
rect 1903 6238 1973 6258
rect 1903 258 1973 278
rect 2061 6238 2131 6258
rect 2061 258 2131 278
rect 2219 6238 2289 6258
rect 2219 258 2289 278
rect 2377 6238 2447 6258
rect 2377 258 2447 278
rect 2535 6238 2605 6258
rect 2535 258 2605 278
rect 2693 6238 2763 6258
rect 2693 258 2763 278
rect 2851 6238 2921 6258
rect 2851 258 2921 278
rect 3009 6238 3079 6258
rect 3009 258 3079 278
rect 3167 6238 3237 6258
rect 3167 258 3237 278
rect 3325 6238 3395 6258
rect 3325 258 3395 278
rect 3483 6238 3553 6258
rect 3483 258 3553 278
rect 3641 6238 3711 6258
rect 3641 258 3711 278
rect 3799 6238 3869 6258
rect 3799 258 3869 278
rect 3957 6238 4027 6258
rect 3957 258 4027 278
rect 4115 6238 4185 6258
rect 4115 258 4185 278
rect 4273 6238 4343 6258
rect 4273 258 4343 278
rect 4431 6238 4501 6258
rect 4431 258 4501 278
rect 4589 6238 4659 6258
rect 4589 258 4659 278
rect 4747 6238 4817 6258
rect 4747 258 4817 278
rect 4905 6238 4975 6258
rect 4905 258 4975 278
rect 232 210 252 226
rect 4886 210 4906 226
rect 232 140 240 210
rect 4890 140 4906 210
rect 232 126 252 140
rect 4886 126 4906 140
rect 30 30 100 100
rect 5040 30 5110 100
<< via2 >>
rect 240 6310 252 6380
rect 252 6310 4886 6380
rect 4886 6310 4900 6380
rect 170 810 230 5710
rect 328 810 388 5710
rect 486 810 546 5710
rect 644 810 704 5710
rect 802 810 862 5710
rect 960 810 1020 5710
rect 1118 810 1178 5710
rect 1276 810 1336 5710
rect 1434 810 1494 5710
rect 1592 810 1652 5710
rect 1750 810 1810 5710
rect 1908 810 1968 5710
rect 2066 810 2126 5710
rect 2224 810 2284 5710
rect 2382 810 2442 5710
rect 2540 810 2600 5710
rect 2698 810 2758 5710
rect 2856 810 2916 5710
rect 3014 810 3074 5710
rect 3172 810 3232 5710
rect 3330 810 3390 5710
rect 3488 810 3548 5710
rect 3646 810 3706 5710
rect 3804 810 3864 5710
rect 3962 810 4022 5710
rect 4120 810 4180 5710
rect 4278 810 4338 5710
rect 4436 810 4496 5710
rect 4594 810 4654 5710
rect 4752 810 4812 5710
rect 4910 810 4970 5710
rect 240 140 252 210
rect 252 140 4886 210
rect 4886 140 4890 210
<< metal3 >>
rect 100 6380 5100 6500
rect 100 6310 240 6380
rect 4900 6310 5100 6380
rect 100 6300 5100 6310
rect 323 6189 393 6190
rect 639 6189 709 6190
rect 955 6189 1025 6190
rect 1271 6189 1341 6190
rect 1587 6189 1657 6190
rect 1903 6189 1973 6190
rect 2219 6189 2289 6190
rect 2535 6189 2605 6190
rect 2851 6189 2921 6190
rect 3167 6189 3237 6190
rect 3483 6189 3553 6190
rect 3799 6189 3869 6190
rect 4115 6189 4185 6190
rect 4431 6189 4501 6190
rect 4747 6189 4817 6190
rect 160 5789 4980 6189
rect 165 5710 235 5720
rect 165 810 170 5710
rect 230 810 235 5710
rect 165 740 235 810
rect 323 5710 393 5789
rect 323 810 328 5710
rect 388 810 393 5710
rect 323 800 393 810
rect 481 5710 551 5720
rect 481 810 486 5710
rect 546 810 551 5710
rect 481 740 551 810
rect 639 5710 709 5789
rect 639 810 644 5710
rect 704 810 709 5710
rect 639 800 709 810
rect 797 5710 867 5720
rect 797 810 802 5710
rect 862 810 867 5710
rect 797 740 867 810
rect 955 5710 1025 5789
rect 955 810 960 5710
rect 1020 810 1025 5710
rect 955 800 1025 810
rect 1113 5710 1183 5720
rect 1113 810 1118 5710
rect 1178 810 1183 5710
rect 1113 740 1183 810
rect 1271 5710 1341 5789
rect 1271 810 1276 5710
rect 1336 810 1341 5710
rect 1271 800 1341 810
rect 1429 5710 1499 5720
rect 1429 810 1434 5710
rect 1494 810 1499 5710
rect 1429 740 1499 810
rect 1587 5710 1657 5789
rect 1587 810 1592 5710
rect 1652 810 1657 5710
rect 1587 800 1657 810
rect 1745 5710 1815 5720
rect 1745 810 1750 5710
rect 1810 810 1815 5710
rect 1745 740 1815 810
rect 1903 5710 1973 5789
rect 1903 810 1908 5710
rect 1968 810 1973 5710
rect 1903 800 1973 810
rect 2061 5710 2131 5720
rect 2061 810 2066 5710
rect 2126 810 2131 5710
rect 2061 740 2131 810
rect 2219 5710 2289 5789
rect 2535 5720 2605 5789
rect 2219 810 2224 5710
rect 2284 810 2289 5710
rect 2219 800 2289 810
rect 2377 5710 2447 5720
rect 2377 810 2382 5710
rect 2442 810 2447 5710
rect 2377 740 2447 810
rect 2535 5710 2606 5720
rect 2535 810 2540 5710
rect 2600 810 2606 5710
rect 2535 800 2606 810
rect 2693 5710 2763 5720
rect 2693 810 2698 5710
rect 2758 810 2763 5710
rect 2693 740 2763 810
rect 2851 5710 2921 5789
rect 2851 810 2856 5710
rect 2916 810 2921 5710
rect 2851 800 2921 810
rect 3009 5710 3079 5720
rect 3009 810 3014 5710
rect 3074 810 3079 5710
rect 3009 740 3079 810
rect 3167 5710 3237 5789
rect 3167 810 3172 5710
rect 3232 810 3237 5710
rect 3167 800 3237 810
rect 3325 5710 3395 5720
rect 3325 810 3330 5710
rect 3390 810 3395 5710
rect 3325 740 3395 810
rect 3483 5710 3553 5789
rect 3483 810 3488 5710
rect 3548 810 3553 5710
rect 3483 800 3553 810
rect 3641 5710 3711 5720
rect 3641 810 3646 5710
rect 3706 810 3711 5710
rect 3641 740 3711 810
rect 3799 5710 3869 5789
rect 3799 810 3804 5710
rect 3864 810 3869 5710
rect 3799 800 3869 810
rect 3957 5710 4027 5720
rect 3957 810 3962 5710
rect 4022 810 4027 5710
rect 3957 740 4027 810
rect 4115 5710 4185 5789
rect 4115 810 4120 5710
rect 4180 810 4185 5710
rect 4115 800 4185 810
rect 4273 5710 4343 5720
rect 4273 810 4278 5710
rect 4338 810 4343 5710
rect 4273 740 4343 810
rect 4431 5710 4501 5789
rect 4431 810 4436 5710
rect 4496 810 4501 5710
rect 4431 800 4501 810
rect 4589 5710 4659 5720
rect 4589 810 4594 5710
rect 4654 810 4659 5710
rect 4589 740 4659 810
rect 4747 5710 4817 5789
rect 4747 810 4752 5710
rect 4812 810 4817 5710
rect 4747 800 4817 810
rect 4905 5710 4975 5720
rect 4905 810 4910 5710
rect 4970 810 4975 5710
rect 4905 740 4975 810
rect 160 340 4980 740
rect 100 210 5100 230
rect 100 140 240 210
rect 4890 140 5100 210
rect 100 30 5100 140
use sky130_fd_pr__nfet_g5v0d10v5_UDPNFN  sky130_fd_pr__nfet_g5v0d10v5_UDPNFN_0
timestamp 1663719933
transform 1 0 2569 0 1 3258
box -2569 -3258 2569 3258
<< labels >>
rlabel metal2 30 6420 100 6480 1 SUB
rlabel metal3 140 6300 200 6500 1 G
rlabel metal3 160 5789 4980 6189 1 SD1
rlabel metal3 160 340 4980 740 1 SD2
<< end >>
