magic
tech sky130B
magscale 1 2
timestamp 1659107503
<< pwell >>
rect -500 3412 714 3420
rect -500 2220 860 3412
<< psubdiff >>
rect -490 3354 -420 3390
rect -490 3320 -470 3354
rect -436 3320 -420 3354
rect -490 3284 -420 3320
rect -490 3250 -470 3284
rect -436 3250 -420 3284
rect -490 3214 -420 3250
rect -490 3180 -470 3214
rect -436 3180 -420 3214
rect -490 3144 -420 3180
rect -490 3110 -470 3144
rect -436 3110 -420 3144
rect -490 3074 -420 3110
rect -490 3040 -470 3074
rect -436 3040 -420 3074
rect -490 3004 -420 3040
rect -490 2970 -470 3004
rect -436 2970 -420 3004
rect -490 2934 -420 2970
rect -490 2900 -470 2934
rect -436 2900 -420 2934
rect -490 2864 -420 2900
rect -490 2830 -470 2864
rect -436 2830 -420 2864
rect -490 2794 -420 2830
rect -490 2760 -470 2794
rect -436 2760 -420 2794
rect -490 2724 -420 2760
rect -490 2690 -470 2724
rect -436 2690 -420 2724
rect -490 2654 -420 2690
rect -490 2620 -470 2654
rect -436 2620 -420 2654
rect -490 2584 -420 2620
rect -490 2550 -470 2584
rect -436 2550 -420 2584
rect -490 2514 -420 2550
rect -490 2480 -470 2514
rect -436 2480 -420 2514
rect -490 2444 -420 2480
rect -490 2410 -470 2444
rect -436 2410 -420 2444
rect -490 2374 -420 2410
rect -490 2340 -470 2374
rect -436 2340 -420 2374
rect -490 2310 -420 2340
rect 780 3354 860 3390
rect 780 3320 800 3354
rect 834 3320 860 3354
rect 780 3284 860 3320
rect 780 3250 800 3284
rect 834 3250 860 3284
rect 780 3214 860 3250
rect 780 3180 800 3214
rect 834 3180 860 3214
rect 780 3144 860 3180
rect 780 3110 800 3144
rect 834 3110 860 3144
rect 780 3074 860 3110
rect 780 3040 800 3074
rect 834 3040 860 3074
rect 780 3004 860 3040
rect 780 2970 800 3004
rect 834 2970 860 3004
rect 780 2934 860 2970
rect 780 2900 800 2934
rect 834 2900 860 2934
rect 780 2864 860 2900
rect 780 2830 800 2864
rect 834 2830 860 2864
rect 780 2794 860 2830
rect 780 2760 800 2794
rect 834 2760 860 2794
rect 780 2724 860 2760
rect 780 2690 800 2724
rect 834 2690 860 2724
rect 780 2654 860 2690
rect 780 2620 800 2654
rect 834 2620 860 2654
rect 780 2584 860 2620
rect 780 2550 800 2584
rect 834 2550 860 2584
rect 780 2514 860 2550
rect 780 2480 800 2514
rect 834 2480 860 2514
rect 780 2444 860 2480
rect 780 2410 800 2444
rect 834 2410 860 2444
rect 780 2374 860 2410
rect 780 2340 800 2374
rect 834 2340 860 2374
rect 780 2310 860 2340
rect -490 2304 860 2310
rect -490 2270 -470 2304
rect -436 2284 800 2304
rect -436 2270 -400 2284
rect -490 2250 -400 2270
rect -366 2250 -330 2284
rect -296 2250 -260 2284
rect -226 2250 -190 2284
rect -156 2250 -120 2284
rect -86 2250 -50 2284
rect -16 2250 20 2284
rect 54 2250 90 2284
rect 124 2250 160 2284
rect 194 2250 230 2284
rect 264 2250 300 2284
rect 334 2250 370 2284
rect 404 2250 440 2284
rect 474 2250 510 2284
rect 544 2250 580 2284
rect 614 2250 650 2284
rect 684 2250 720 2284
rect 754 2270 800 2284
rect 834 2270 860 2304
rect 754 2250 860 2270
rect -490 2230 860 2250
<< psubdiffcont >>
rect -470 3320 -436 3354
rect -470 3250 -436 3284
rect -470 3180 -436 3214
rect -470 3110 -436 3144
rect -470 3040 -436 3074
rect -470 2970 -436 3004
rect -470 2900 -436 2934
rect -470 2830 -436 2864
rect -470 2760 -436 2794
rect -470 2690 -436 2724
rect -470 2620 -436 2654
rect -470 2550 -436 2584
rect -470 2480 -436 2514
rect -470 2410 -436 2444
rect -470 2340 -436 2374
rect 800 3320 834 3354
rect 800 3250 834 3284
rect 800 3180 834 3214
rect 800 3110 834 3144
rect 800 3040 834 3074
rect 800 2970 834 3004
rect 800 2900 834 2934
rect 800 2830 834 2864
rect 800 2760 834 2794
rect 800 2690 834 2724
rect 800 2620 834 2654
rect 800 2550 834 2584
rect 800 2480 834 2514
rect 800 2410 834 2444
rect 800 2340 834 2374
rect -470 2270 -436 2304
rect -400 2250 -366 2284
rect -330 2250 -296 2284
rect -260 2250 -226 2284
rect -190 2250 -156 2284
rect -120 2250 -86 2284
rect -50 2250 -16 2284
rect 20 2250 54 2284
rect 90 2250 124 2284
rect 160 2250 194 2284
rect 230 2250 264 2284
rect 300 2250 334 2284
rect 370 2250 404 2284
rect 440 2250 474 2284
rect 510 2250 544 2284
rect 580 2250 614 2284
rect 650 2250 684 2284
rect 720 2250 754 2284
rect 800 2270 834 2304
<< poly >>
rect -5 3479 17 3483
rect -5 3417 24 3479
rect 2 3413 24 3417
<< polycont >>
rect -316 3429 -282 3463
rect -44 3429 -10 3463
rect 24 3429 58 3463
rect 300 3429 334 3463
rect 368 3429 402 3463
<< locali >>
rect -332 3429 -316 3463
rect -282 3429 -44 3463
rect -10 3429 24 3463
rect 58 3429 300 3463
rect 334 3429 368 3463
rect 402 3429 714 3463
rect -480 3354 -430 3370
rect -480 3320 -470 3354
rect -436 3320 -430 3354
rect -480 3284 -430 3320
rect -480 3240 -470 3284
rect -436 3240 -430 3284
rect -480 3214 -430 3240
rect -480 3160 -470 3214
rect -436 3160 -430 3214
rect -480 3144 -430 3160
rect -480 3080 -470 3144
rect -436 3080 -430 3144
rect -480 3074 -430 3080
rect -480 3040 -470 3074
rect -436 3040 -430 3074
rect -480 3034 -430 3040
rect -480 2970 -470 3034
rect -436 2970 -430 3034
rect -480 2954 -430 2970
rect -480 2900 -470 2954
rect -436 2900 -430 2954
rect -480 2874 -430 2900
rect -480 2830 -470 2874
rect -436 2830 -430 2874
rect -480 2794 -430 2830
rect -480 2760 -470 2794
rect -436 2760 -430 2794
rect -480 2724 -430 2760
rect -480 2680 -470 2724
rect -436 2680 -430 2724
rect -480 2654 -430 2680
rect -480 2600 -470 2654
rect -436 2600 -430 2654
rect -480 2584 -430 2600
rect -480 2520 -470 2584
rect -436 2520 -430 2584
rect -480 2514 -430 2520
rect -480 2480 -470 2514
rect -436 2480 -430 2514
rect -480 2474 -430 2480
rect -480 2410 -470 2474
rect -436 2410 -430 2474
rect -480 2394 -430 2410
rect -480 2340 -470 2394
rect -436 2340 -430 2394
rect -480 2314 -430 2340
rect -480 2270 -470 2314
rect -436 2300 -430 2314
rect 790 3354 850 3370
rect 790 3320 800 3354
rect 834 3320 850 3354
rect 790 3284 850 3320
rect 790 3240 800 3284
rect 834 3240 850 3284
rect 790 3214 850 3240
rect 790 3160 800 3214
rect 834 3160 850 3214
rect 790 3144 850 3160
rect 790 3080 800 3144
rect 834 3080 850 3144
rect 790 3074 850 3080
rect 790 3040 800 3074
rect 834 3040 850 3074
rect 790 3034 850 3040
rect 790 2970 800 3034
rect 834 2970 850 3034
rect 790 2954 850 2970
rect 790 2900 800 2954
rect 834 2900 850 2954
rect 790 2874 850 2900
rect 790 2830 800 2874
rect 834 2830 850 2874
rect 790 2794 850 2830
rect 790 2760 800 2794
rect 834 2760 850 2794
rect 790 2724 850 2760
rect 790 2680 800 2724
rect 834 2680 850 2724
rect 790 2654 850 2680
rect 790 2600 800 2654
rect 834 2600 850 2654
rect 790 2584 850 2600
rect 790 2520 800 2584
rect 834 2520 850 2584
rect 790 2514 850 2520
rect 790 2480 800 2514
rect 834 2480 850 2514
rect 790 2474 850 2480
rect 790 2410 800 2474
rect 834 2410 850 2474
rect 790 2394 850 2410
rect 790 2340 800 2394
rect 834 2340 850 2394
rect 790 2314 850 2340
rect 790 2300 800 2314
rect -436 2284 800 2300
rect -436 2270 -400 2284
rect -480 2250 -400 2270
rect -356 2250 -330 2284
rect -276 2250 -260 2284
rect -196 2250 -190 2284
rect -156 2250 -150 2284
rect -86 2250 -70 2284
rect -16 2250 10 2284
rect 54 2250 90 2284
rect 124 2250 160 2284
rect 204 2250 230 2284
rect 284 2250 300 2284
rect 364 2250 370 2284
rect 404 2250 410 2284
rect 474 2250 490 2284
rect 544 2250 570 2284
rect 614 2250 650 2284
rect 684 2250 720 2284
rect 754 2270 800 2284
rect 834 2270 850 2314
rect 754 2250 850 2270
rect -480 2240 850 2250
<< viali >>
rect -470 3320 -436 3354
rect -470 3250 -436 3274
rect -470 3240 -436 3250
rect -470 3180 -436 3194
rect -470 3160 -436 3180
rect -470 3110 -436 3114
rect -470 3080 -436 3110
rect -470 3004 -436 3034
rect -470 3000 -436 3004
rect -470 2934 -436 2954
rect -470 2920 -436 2934
rect -470 2864 -436 2874
rect -470 2840 -436 2864
rect -470 2760 -436 2794
rect -470 2690 -436 2714
rect -470 2680 -436 2690
rect -470 2620 -436 2634
rect -470 2600 -436 2620
rect -470 2550 -436 2554
rect -470 2520 -436 2550
rect -470 2444 -436 2474
rect -470 2440 -436 2444
rect -470 2374 -436 2394
rect -470 2360 -436 2374
rect -470 2304 -436 2314
rect -470 2280 -436 2304
rect 800 3320 834 3354
rect 800 3250 834 3274
rect 800 3240 834 3250
rect 800 3180 834 3194
rect 800 3160 834 3180
rect 800 3110 834 3114
rect 800 3080 834 3110
rect 800 3004 834 3034
rect 800 3000 834 3004
rect 800 2934 834 2954
rect 800 2920 834 2934
rect 800 2864 834 2874
rect 800 2840 834 2864
rect 800 2760 834 2794
rect 800 2690 834 2714
rect 800 2680 834 2690
rect 800 2620 834 2634
rect 800 2600 834 2620
rect 800 2550 834 2554
rect 800 2520 834 2550
rect 800 2444 834 2474
rect 800 2440 834 2444
rect 800 2374 834 2394
rect 800 2360 834 2374
rect 800 2304 834 2314
rect -390 2250 -366 2284
rect -366 2250 -356 2284
rect -310 2250 -296 2284
rect -296 2250 -276 2284
rect -230 2250 -226 2284
rect -226 2250 -196 2284
rect -150 2250 -120 2284
rect -120 2250 -116 2284
rect -70 2250 -50 2284
rect -50 2250 -36 2284
rect 10 2250 20 2284
rect 20 2250 44 2284
rect 90 2250 124 2284
rect 170 2250 194 2284
rect 194 2250 204 2284
rect 250 2250 264 2284
rect 264 2250 284 2284
rect 330 2250 334 2284
rect 334 2250 364 2284
rect 410 2250 440 2284
rect 440 2250 444 2284
rect 490 2250 510 2284
rect 510 2250 524 2284
rect 570 2250 580 2284
rect 580 2250 604 2284
rect 650 2250 684 2284
rect 800 2280 834 2304
<< metal1 >>
rect -340 3520 710 3580
rect -5 3417 17 3483
rect -490 3380 -420 3390
rect 780 3380 850 3390
rect -490 3354 -310 3380
rect -490 3320 -470 3354
rect -436 3320 -310 3354
rect -490 3274 -310 3320
rect -490 3240 -470 3274
rect -436 3240 -310 3274
rect -490 3194 -310 3240
rect -490 3160 -470 3194
rect -436 3160 -310 3194
rect -490 3114 -310 3160
rect -490 3080 -470 3114
rect -436 3080 -310 3114
rect -490 3034 -310 3080
rect -490 3000 -470 3034
rect -436 3000 -310 3034
rect -490 2954 -310 3000
rect -490 2920 -470 2954
rect -436 2920 -310 2954
rect -490 2874 -310 2920
rect -490 2840 -470 2874
rect -436 2840 -310 2874
rect -490 2794 -310 2840
rect -490 2760 -470 2794
rect -436 2760 -310 2794
rect -490 2714 -310 2760
rect -490 2680 -470 2714
rect -436 2680 -310 2714
rect -490 2634 -310 2680
rect -490 2600 -470 2634
rect -436 2600 -310 2634
rect -490 2554 -310 2600
rect -490 2520 -470 2554
rect -436 2520 -310 2554
rect -490 2474 -310 2520
rect -490 2440 -470 2474
rect -436 2440 -310 2474
rect -490 2394 -310 2440
rect -490 2360 -470 2394
rect -436 2360 -310 2394
rect -490 2314 -310 2360
rect -490 2280 -470 2314
rect -436 2284 -310 2314
rect 680 3354 850 3380
rect 680 3320 800 3354
rect 834 3320 850 3354
rect 680 3274 850 3320
rect 680 3240 800 3274
rect 834 3240 850 3274
rect 680 3194 850 3240
rect 680 3160 800 3194
rect 834 3160 850 3194
rect 680 3114 850 3160
rect 680 3080 800 3114
rect 834 3080 850 3114
rect 680 3034 850 3080
rect 680 3000 800 3034
rect 834 3000 850 3034
rect 680 2954 850 3000
rect 680 2920 800 2954
rect 834 2920 850 2954
rect 680 2874 850 2920
rect 680 2840 800 2874
rect 834 2840 850 2874
rect 680 2794 850 2840
rect 680 2760 800 2794
rect 834 2760 850 2794
rect 680 2714 850 2760
rect 680 2680 800 2714
rect 834 2680 850 2714
rect 680 2634 850 2680
rect 680 2600 800 2634
rect 834 2600 850 2634
rect 680 2554 850 2600
rect 680 2520 800 2554
rect 834 2520 850 2554
rect 680 2474 850 2520
rect 680 2440 800 2474
rect 834 2440 850 2474
rect 680 2394 850 2440
rect 680 2360 800 2394
rect 834 2360 850 2394
rect 680 2314 850 2360
rect 680 2284 800 2314
rect -436 2280 -390 2284
rect -490 2250 -390 2280
rect -356 2250 -310 2284
rect 684 2280 800 2284
rect 834 2280 850 2314
rect 684 2250 850 2280
rect -490 2230 850 2250
rect -490 2210 -370 2230
<< metal2 >>
rect -340 3420 730 3500
use sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap  sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0
timestamp 1659107442
transform 1 0 -501 0 1 2289
box 100 -41 576 1290
use sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap  sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_1
timestamp 1659107442
transform 1 0 -157 0 1 2289
box 100 -41 576 1290
use sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap  sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_2
timestamp 1659107442
transform 1 0 187 0 1 2289
box 100 -41 576 1290
<< labels >>
rlabel metal1 -490 2210 -370 2230 1 S
rlabel metal1 -340 3520 -310 3580 1 G
rlabel metal2 -340 3420 -300 3500 1 SD
<< end >>
