magic
tech sky130B
timestamp 1662741506
<< metal4 >>
rect 0 -48580 60 0
rect 100 -48580 160 0
rect 200 -48580 260 0
rect 300 -48580 360 0
rect 400 -48580 460 0
rect 500 -48580 560 0
rect 600 -48580 660 0
rect 700 -48580 760 0
rect 800 -48580 860 0
rect 900 -38840 960 0
rect 1000 -38740 1060 0
rect 1100 -38640 1160 0
rect 1200 -38580 1260 0
rect 1300 -38490 1360 0
rect 1400 -5580 1460 0
rect 1500 -5580 1560 0
rect 1600 -5580 1660 0
rect 1700 -5580 1760 0
rect 1800 -5580 1860 0
rect 1900 -5580 1960 0
rect 2000 -5580 2060 0
rect 2100 -5580 2160 0
rect 2200 -5580 2260 0
rect 2300 -5580 2360 0
rect 2400 -5580 2460 0
rect 2500 -5580 2560 0
rect 2600 -5580 2660 0
rect 2700 -5580 2760 0
rect 2800 -5580 2860 0
rect 2900 -5580 2960 0
rect 3000 -5580 3060 0
rect 3100 -5580 3160 0
rect 3200 -5580 3260 0
rect 3300 -5580 3360 0
rect 3400 -5580 3460 0
rect 3500 -5580 3560 0
rect 3600 -5580 3660 0
rect 3700 -5580 3760 0
rect 3800 -5580 3860 0
rect 3900 -5580 3960 0
rect 4000 -5580 4060 0
rect 4100 -5580 4160 0
rect 4200 -5580 4260 0
rect 4300 -5580 4360 0
rect 4400 -5580 4460 0
rect 4500 -5580 4560 0
rect 4600 -5580 4660 0
rect 4700 -5580 4760 0
rect 4800 -5580 4860 0
rect 4900 -5580 4960 0
rect 5000 -5580 5060 0
rect 5100 -5580 5160 0
rect 5200 -5580 5260 0
rect 5300 -5580 5360 0
rect 5400 -5580 5460 0
rect 5500 -5580 5560 0
rect 5600 -5580 5660 0
rect 5700 -5580 5760 0
rect 5800 -5580 5860 0
rect 5900 -5580 5960 0
rect 6000 -5580 6060 0
rect 6100 -5580 6160 0
rect 6200 -5990 6260 0
rect 1400 -8270 1460 -6290
rect 1500 -8210 1560 -6300
rect 1600 -8160 1660 -6300
rect 1700 -8110 1760 -6300
rect 1800 -8060 1860 -6300
rect 1900 -8020 1960 -6300
rect 2000 -7970 2060 -6300
rect 2100 -7920 2160 -6300
rect 2200 -7870 2260 -6300
rect 2300 -7830 2360 -6300
rect 2400 -7780 2460 -6300
rect 2500 -7730 2560 -6300
rect 2600 -7680 2660 -6300
rect 2700 -7630 2760 -6300
rect 2800 -7580 2860 -6300
rect 2900 -7530 2960 -6300
rect 3000 -7490 3060 -6300
rect 3100 -7440 3160 -6300
rect 3200 -7390 3260 -6300
rect 3300 -7340 3360 -6300
rect 3400 -7290 3460 -6300
rect 4100 -7700 4160 -6300
rect 4200 -7930 4260 -6290
rect 1400 -9760 1460 -9090
rect 1500 -9760 1560 -9040
rect 1600 -9760 1660 -8990
rect 1700 -9760 1760 -8940
rect 1800 -9760 1860 -8880
rect 1900 -9760 1960 -8830
rect 2000 -9760 2060 -8780
rect 2100 -9760 2160 -8730
rect 2200 -9760 2260 -8680
rect 2300 -9760 2360 -8620
rect 2400 -9760 2460 -8570
rect 2500 -9760 2560 -8520
rect 2600 -9760 2660 -8470
rect 2700 -9760 2760 -8420
rect 2800 -9760 2860 -8360
rect 2900 -9760 2960 -8310
rect 3000 -9760 3060 -8260
rect 3100 -9760 3160 -8210
rect 3200 -9760 3260 -8160
rect 3300 -9760 3360 -8100
rect 3400 -9760 3460 -8050
rect 3500 -9760 3560 -8010
rect 4300 -8050 4360 -6300
rect 3600 -9760 3660 -8120
rect 4400 -8130 4460 -6300
rect 4500 -8190 4560 -6300
rect 4600 -8230 4660 -6300
rect 4700 -8260 4760 -6300
rect 4800 -8280 4860 -6300
rect 4900 -8280 4960 -6300
rect 5000 -8270 5060 -6300
rect 5100 -8240 5160 -6300
rect 5200 -8220 5260 -6300
rect 5300 -8160 5360 -6300
rect 5400 -8080 5460 -6300
rect 5500 -7960 5560 -6290
rect 5600 -7660 5660 -6310
rect 3700 -9760 3760 -8310
rect 3800 -9760 3860 -8450
rect 3900 -9760 3960 -8560
rect 4000 -9760 4060 -8650
rect 4100 -9760 4160 -8730
rect 4200 -9760 4260 -8780
rect 4300 -9760 4360 -8830
rect 4400 -9760 4460 -8870
rect 4500 -9760 4560 -8890
rect 4600 -9760 4660 -8910
rect 4700 -9760 4760 -8920
rect 4800 -9760 4860 -8930
rect 4900 -9760 4960 -8930
rect 5000 -9760 5060 -8920
rect 5100 -9760 5160 -8910
rect 5200 -9760 5260 -8900
rect 5300 -9760 5360 -8870
rect 5400 -9760 5460 -8830
rect 5500 -9760 5560 -8780
rect 5600 -9760 5660 -8730
rect 5700 -9760 5760 -8660
rect 5800 -9760 5860 -8560
rect 5900 -9760 5960 -8450
rect 6000 -9760 6060 -8310
rect 6100 -9760 6160 -8100
rect 6200 -9770 6260 -7560
rect 1400 -12370 1460 -10470
rect 1500 -11990 1560 -10470
rect 1600 -11740 1660 -10470
rect 1700 -11550 1760 -10470
rect 1800 -11390 1860 -10470
rect 1900 -11250 1960 -10470
rect 2000 -11160 2060 -10470
rect 2100 -11240 2160 -10470
rect 2200 -11330 2260 -10470
rect 2300 -11410 2360 -10470
rect 2400 -11500 2460 -10470
rect 2100 -13520 2160 -12370
rect 1400 -16690 1460 -13520
rect 2200 -13710 2260 -12090
rect 2300 -13820 2360 -11870
rect 2400 -13880 2460 -11740
rect 1500 -16380 1560 -13880
rect 2500 -13930 2560 -10470
rect 2600 -13940 2660 -10470
rect 2700 -13960 2760 -10470
rect 2800 -13960 2860 -10470
rect 2900 -13940 2960 -10470
rect 3000 -13920 3060 -10470
rect 3100 -13870 3160 -10470
rect 3200 -13790 3260 -10470
rect 3300 -13660 3360 -10470
rect 3400 -13420 3460 -10470
rect 3500 -12770 3560 -10470
rect 3600 -12310 3660 -10470
rect 3700 -12080 3760 -10470
rect 3800 -11910 3860 -10470
rect 3900 -11790 3960 -10470
rect 4000 -11690 4060 -10470
rect 4100 -11610 4160 -10470
rect 4200 -11540 4260 -10470
rect 4300 -11500 4360 -10470
rect 4400 -11450 4460 -10470
rect 4500 -11420 4560 -10470
rect 4600 -11410 4660 -10470
rect 4700 -11390 4760 -10470
rect 4800 -11380 4860 -10470
rect 4900 -11380 4960 -10470
rect 5000 -11390 5060 -10470
rect 5100 -11410 5160 -10470
rect 5200 -11410 5260 -10470
rect 5300 -11450 5360 -10470
rect 5400 -11480 5460 -10470
rect 5500 -11530 5560 -10470
rect 5600 -11580 5660 -10470
rect 5700 -11660 5760 -10470
rect 5800 -11740 5860 -10470
rect 5900 -11850 5960 -10470
rect 6000 -11980 6060 -10470
rect 1600 -16190 1660 -14080
rect 1700 -16060 1760 -14220
rect 1800 -15930 1860 -14330
rect 1900 -15830 1960 -14420
rect 2000 -15750 2060 -14480
rect 2100 -15670 2160 -14530
rect 2200 -15620 2260 -14570
rect 2300 -15560 2360 -14610
rect 2400 -15520 2460 -14630
rect 2500 -15500 2560 -14650
rect 2600 -15460 2660 -14660
rect 2700 -15450 2760 -14660
rect 2800 -15440 2860 -14660
rect 2900 -15420 2960 -14660
rect 3000 -15420 3060 -14650
rect 3100 -15420 3160 -14620
rect 3200 -15420 3260 -14590
rect 3300 -15420 3360 -14550
rect 3400 -15420 3460 -14500
rect 3500 -15420 3560 -14440
rect 3600 -15420 3660 -14360
rect 3700 -15420 3760 -14270
rect 3800 -15420 3860 -14170
rect 3900 -15420 3960 -13990
rect 4000 -15420 4060 -13760
rect 4100 -15420 4160 -13350
rect 4200 -15420 4260 -12690
rect 4300 -15420 4360 -12430
rect 4400 -15420 4460 -12300
rect 4500 -15420 4560 -12200
rect 4600 -15420 4660 -12140
rect 4700 -15420 4760 -12100
rect 4800 -15420 4860 -12090
rect 4900 -15420 4960 -12090
rect 5000 -15420 5060 -12100
rect 5100 -15420 5160 -12140
rect 5200 -15420 5260 -12180
rect 6100 -12190 6160 -10470
rect 5300 -13960 5360 -12240
rect 5400 -13760 5460 -12340
rect 5500 -13470 5560 -12510
rect 6200 -12530 6260 -10460
rect 5300 -15420 5360 -14190
rect 5400 -15420 5460 -14260
rect 5500 -15420 5560 -14330
rect 5600 -15420 5660 -14400
rect 5700 -15420 5760 -14470
rect 5800 -15420 5860 -14450
rect 5900 -15420 5960 -14290
rect 6000 -15420 6060 -14080
rect 6100 -15420 6160 -13840
rect 6200 -15430 6260 -13430
rect 2100 -17580 2160 -16700
rect 1400 -23340 1460 -17590
rect 2200 -17750 2260 -16530
rect 2300 -17860 2360 -16410
rect 1500 -23070 1560 -17900
rect 2400 -17940 2460 -16330
rect 2500 -18010 2560 -16270
rect 2600 -18060 2660 -16220
rect 2700 -18090 2760 -16180
rect 1600 -22910 1660 -18100
rect 2800 -18120 2860 -16150
rect 2900 -18130 2960 -16140
rect 3000 -18140 3060 -16130
rect 1700 -22780 1760 -18220
rect 1800 -22680 1860 -18350
rect 1900 -19390 1960 -18440
rect 2000 -19200 2060 -18540
rect 2100 -19010 2160 -18610
rect 2200 -18870 2260 -18590
rect 2300 -18770 2360 -18490
rect 2400 -18640 2460 -18430
rect 2500 -18570 2560 -18360
rect 2600 -18500 2660 -18310
rect 2700 -18460 2760 -18270
rect 2800 -18420 2860 -18230
rect 2900 -18420 2960 -18230
rect 3000 -18420 3060 -18200
rect 3100 -18460 3160 -16130
rect 3200 -18450 3260 -16120
rect 3300 -17950 3360 -16120
rect 3400 -17850 3460 -16120
rect 3500 -17700 3560 -16120
rect 3600 -17600 3660 -16120
rect 3700 -17500 3760 -16120
rect 3800 -17420 3860 -16120
rect 3900 -17350 3960 -16120
rect 4000 -17300 4060 -16120
rect 4100 -17250 4160 -16120
rect 4200 -17200 4260 -16120
rect 4300 -17170 4360 -16120
rect 4400 -17160 4460 -16120
rect 4500 -17200 4560 -16120
rect 4600 -17200 4660 -16120
rect 4700 -17210 4760 -16120
rect 4800 -17260 4860 -16120
rect 4900 -17310 4960 -16120
rect 5000 -17330 5060 -16120
rect 5100 -17200 5160 -16120
rect 5200 -17100 5260 -16120
rect 5300 -17020 5360 -16120
rect 5400 -16980 5460 -16120
rect 5500 -16980 5560 -16120
rect 5600 -16980 5660 -16120
rect 5700 -16940 5760 -16120
rect 5800 -16940 5860 -16120
rect 5900 -16940 5960 -16120
rect 6000 -16940 6060 -16120
rect 6100 -16980 6160 -16130
rect 6200 -16980 6260 -16100
rect 6300 -17010 6360 0
rect 6400 -17030 6460 0
rect 6500 -17030 6560 0
rect 6600 -17070 6660 0
rect 6700 -17120 6760 0
rect 1900 -19510 1960 -19450
rect 1900 -20300 1960 -20210
rect 1900 -22590 1960 -20360
rect 2100 -20390 2160 -19340
rect 2100 -20530 2160 -20450
rect 2000 -22530 2060 -20710
rect 2200 -20800 2260 -19150
rect 2100 -22470 2160 -20930
rect 2300 -20980 2360 -19010
rect 2200 -22430 2260 -21120
rect 2400 -21170 2460 -18910
rect 2300 -22410 2360 -21350
rect 2500 -21400 2560 -18790
rect 2600 -21540 2660 -18710
rect 2400 -22380 2460 -21540
rect 2500 -22370 2560 -21680
rect 2700 -21690 2760 -18650
rect 2800 -21790 2860 -18620
rect 2600 -22360 2660 -21830
rect 2900 -21930 2960 -18620
rect 2700 -22470 2760 -21930
rect 3000 -22070 3060 -18630
rect 2800 -22620 2860 -22070
rect 3100 -22130 3160 -18660
rect 3200 -22170 3260 -18660
rect 2900 -22720 2960 -22220
rect 3300 -22240 3360 -18580
rect 3000 -22860 3060 -22280
rect 3400 -22300 3460 -18180
rect 3100 -22960 3160 -22330
rect 3500 -22380 3560 -17980
rect 3600 -22410 3660 -17840
rect 3700 -22120 3760 -17750
rect 3800 -21800 3860 -17650
rect 3900 -21620 3960 -17550
rect 4000 -20730 4060 -17500
rect 4100 -20780 4160 -17450
rect 4200 -20880 4260 -17400
rect 4300 -20950 4360 -17370
rect 4400 -21020 4460 -17360
rect 4500 -20930 4560 -17400
rect 4600 -20740 4660 -17400
rect 4700 -20420 4760 -17410
rect 4800 -20230 4860 -17460
rect 4900 -20160 4960 -17550
rect 5000 -20160 5060 -17700
rect 5100 -20210 5160 -17690
rect 5200 -20260 5260 -17340
rect 5300 -20320 5360 -17240
rect 5400 -20380 5460 -17180
rect 4800 -20620 4860 -20560
rect 3800 -22400 3860 -22340
rect 2000 -23930 2060 -23490
rect 1400 -26560 1460 -24110
rect 2100 -24150 2160 -23280
rect 2200 -24250 2260 -23170
rect 2300 -24320 2360 -23110
rect 2400 -24360 2460 -23060
rect 1500 -26330 1560 -24370
rect 2500 -24380 2560 -23050
rect 2600 -24410 2660 -23020
rect 2700 -24420 2760 -23010
rect 2800 -24420 2860 -23010
rect 2900 -24420 2960 -23010
rect 3000 -24420 3060 -23010
rect 3100 -24420 3160 -23020
rect 3200 -24420 3260 -22630
rect 3500 -22760 3560 -22620
rect 3300 -24420 3360 -22880
rect 3600 -22940 3660 -22620
rect 3400 -24420 3460 -23100
rect 3700 -23130 3760 -22660
rect 3800 -23260 3860 -22460
rect 3500 -24420 3560 -23290
rect 3900 -23450 3960 -21980
rect 3600 -24420 3660 -23520
rect 4000 -23590 4060 -21750
rect 3700 -24420 3760 -23670
rect 4100 -23740 4160 -21470
rect 3800 -24420 3860 -23810
rect 4200 -23840 4260 -21110
rect 3900 -24540 3960 -23900
rect 4300 -23940 4360 -21170
rect 4400 -23990 4460 -21230
rect 4500 -21760 4560 -21210
rect 4600 -21430 4660 -21070
rect 4700 -21340 4760 -20880
rect 4800 -21340 4860 -20680
rect 4600 -22590 4660 -21940
rect 1600 -26170 1660 -24540
rect 1700 -26050 1760 -24660
rect 1800 -25970 1860 -24760
rect 1900 -25890 1960 -24840
rect 2000 -25830 2060 -24900
rect 2100 -25780 2160 -24960
rect 2200 -25730 2260 -25000
rect 2300 -25700 2360 -25020
rect 4000 -25030 4060 -24050
rect 2400 -25680 2460 -25050
rect 2500 -25660 2560 -25060
rect 2600 -25650 2660 -25070
rect 2700 -25640 2760 -25080
rect 2800 -25650 2860 -25090
rect 2900 -25680 2960 -25090
rect 3000 -25690 3060 -25090
rect 3100 -25710 3160 -25080
rect 3200 -25730 3260 -25080
rect 3300 -25750 3360 -25090
rect 3400 -25780 3460 -25090
rect 3500 -25820 3560 -25090
rect 3600 -25850 3660 -25080
rect 3700 -25900 3760 -25090
rect 3800 -25930 3860 -25090
rect 3900 -25980 3960 -25090
rect 4000 -26030 4060 -25090
rect 4100 -26070 4160 -24200
rect 4200 -26120 4260 -24300
rect 4300 -26170 4360 -25090
rect 4500 -25270 4560 -22720
rect 4700 -22860 4760 -21620
rect 4600 -23110 4660 -23050
rect 4400 -26220 4460 -25450
rect 4600 -25540 4660 -23170
rect 4800 -23180 4860 -21560
rect 4900 -23360 4960 -20420
rect 2000 -27200 2060 -26960
rect 1400 -30820 1460 -27440
rect 2100 -27460 2160 -26630
rect 2200 -27580 2260 -26510
rect 2300 -27670 2360 -26440
rect 1500 -30820 1560 -27700
rect 2400 -27720 2460 -26400
rect 2500 -27770 2560 -26360
rect 2600 -27780 2660 -26340
rect 2700 -27800 2760 -26330
rect 2800 -27800 2860 -26320
rect 2900 -27790 2960 -26320
rect 3000 -27780 3060 -26320
rect 3100 -27780 3160 -26350
rect 4500 -26360 4560 -25720
rect 4700 -25780 4760 -23360
rect 5000 -23460 5060 -20400
rect 5100 -23480 5160 -20420
rect 5500 -20440 5560 -17180
rect 5200 -23490 5260 -20470
rect 5600 -20490 5660 -17160
rect 5700 -20540 5760 -17140
rect 5300 -23430 5360 -20540
rect 5800 -20560 5860 -17140
rect 5900 -20590 5960 -17140
rect 5400 -23340 5460 -20590
rect 6000 -20630 6060 -17140
rect 6100 -20640 6160 -17150
rect 6800 -17170 6860 0
rect 6200 -20640 6260 -17180
rect 6300 -20610 6360 -17180
rect 6900 -17220 6960 0
rect 6400 -20590 6460 -17220
rect 6500 -20500 6560 -17230
rect 6600 -20440 6660 -17270
rect 7000 -17290 7060 0
rect 5500 -23280 5560 -20640
rect 5600 -23180 5660 -20690
rect 5700 -23130 5760 -20740
rect 5800 -23070 5860 -20770
rect 5900 -23030 5960 -20790
rect 6000 -23030 6060 -20790
rect 6100 -23030 6160 -20790
rect 6200 -23030 6260 -20790
rect 6300 -23030 6360 -20790
rect 6400 -23030 6460 -20790
rect 6500 -23030 6560 -20750
rect 6600 -23030 6660 -20680
rect 6700 -23060 6760 -17320
rect 7100 -17360 7160 0
rect 6800 -20460 6860 -17370
rect 7200 -17430 7260 0
rect 6900 -20010 6960 -17440
rect 7000 -19610 7060 -17520
rect 7100 -19380 7160 -17570
rect 7300 -17580 7360 0
rect 7200 -19140 7260 -17670
rect 7400 -17680 7460 0
rect 7300 -18960 7360 -17810
rect 7500 -17870 7560 0
rect 7500 -17990 7560 -17930
rect 7400 -18680 7460 -18270
rect 7600 -18580 7660 0
rect 7700 -18570 7760 0
rect 7800 -18460 7860 0
rect 7900 -18370 7960 0
rect 8000 -18330 8060 0
rect 8100 -18320 8160 0
rect 8200 -18290 8260 0
rect 8300 -18330 8360 0
rect 8400 -18340 8460 0
rect 8500 -18370 8560 0
rect 8600 -18440 8660 0
rect 7400 -18860 7460 -18740
rect 7600 -18910 7660 -18850
rect 7000 -21010 7060 -20190
rect 7100 -20990 7160 -19880
rect 7200 -20940 7260 -19510
rect 7300 -20900 7360 -19280
rect 7400 -20860 7460 -19100
rect 7500 -20860 7560 -19010
rect 7600 -20900 7660 -18990
rect 7700 -20900 7760 -18800
rect 7800 -20940 7860 -18680
rect 7900 -20940 7960 -18600
rect 8000 -20940 8060 -18530
rect 8100 -20940 8160 -18500
rect 8200 -20940 8260 -18490
rect 8300 -20910 8360 -18520
rect 8400 -20900 8460 -18530
rect 8700 -18580 8760 0
rect 8500 -20900 8560 -18580
rect 8800 -18680 8860 0
rect 8600 -20900 8660 -18720
rect 8900 -18820 8960 0
rect 8700 -20860 8760 -18820
rect 8800 -20820 8860 -18960
rect 9000 -19020 9060 0
rect 8900 -20760 8960 -19190
rect 9100 -19250 9160 0
rect 9000 -19440 9060 -19380
rect 9200 -19470 9260 0
rect 9000 -20680 9060 -19500
rect 6800 -23090 6860 -21060
rect 6900 -23120 6960 -21250
rect 7000 -23130 7060 -21250
rect 7100 -23140 7160 -21190
rect 7200 -23100 7260 -21150
rect 7300 -23030 7360 -21100
rect 7400 -21430 7460 -21050
rect 7500 -21420 7560 -21050
rect 7600 -21540 7660 -21100
rect 7400 -22950 7460 -21570
rect 7500 -22890 7560 -21670
rect 7700 -21770 7760 -21100
rect 7600 -22790 7660 -21940
rect 7800 -22560 7860 -21100
rect 3200 -27750 3260 -26390
rect 3300 -27710 3360 -26440
rect 3400 -27650 3460 -26500
rect 4600 -26590 4660 -25960
rect 4800 -26000 4860 -23500
rect 3500 -27560 3560 -26590
rect 3600 -27400 3660 -26740
rect 4700 -26820 4760 -26230
rect 4900 -26290 4960 -23600
rect 4200 -27020 4260 -26860
rect 1600 -30820 1660 -27870
rect 1700 -30820 1760 -27990
rect 1800 -30820 1860 -28090
rect 1900 -30820 1960 -28170
rect 2000 -30820 2060 -28230
rect 2100 -30790 2160 -28290
rect 2200 -28780 2260 -28330
rect 2300 -28780 2360 -28370
rect 2400 -28780 2460 -28410
rect 2500 -28780 2560 -28430
rect 2600 -28780 2660 -28450
rect 2700 -28780 2760 -28450
rect 2800 -28820 2860 -28450
rect 2900 -28860 2960 -28450
rect 3000 -28910 3060 -28450
rect 3100 -28960 3160 -28450
rect 3200 -29000 3260 -28450
rect 3300 -29050 3360 -28420
rect 3400 -29090 3460 -28400
rect 3500 -29140 3560 -28360
rect 3600 -29190 3660 -28320
rect 3700 -29240 3760 -28270
rect 3800 -29280 3860 -28190
rect 3900 -29330 3960 -28110
rect 4000 -29380 4060 -27990
rect 4100 -29420 4160 -27840
rect 4200 -29470 4260 -27510
rect 4300 -29520 4360 -26890
rect 2700 -29640 2760 -29580
rect 2800 -30820 2860 -29540
rect 4400 -29560 4460 -26950
rect 2900 -30820 2960 -29580
rect 4500 -29610 4560 -27000
rect 4800 -27050 4860 -26420
rect 5000 -26470 5060 -23660
rect 3000 -30820 3060 -29630
rect 4600 -29650 4660 -27050
rect 3100 -30820 3160 -29670
rect 4700 -29700 4760 -27110
rect 3200 -30820 3260 -29720
rect 4800 -29750 4860 -27150
rect 3300 -30820 3360 -29770
rect 4900 -29790 4960 -26600
rect 5100 -26660 5160 -23660
rect 3400 -30820 3460 -29820
rect 5000 -29840 5060 -26840
rect 5200 -26890 5260 -23660
rect 5300 -27030 5360 -23640
rect 3500 -30820 3560 -29860
rect 5100 -29890 5160 -27030
rect 3600 -30820 3660 -29910
rect 5200 -29940 5260 -27160
rect 5400 -27210 5460 -23580
rect 3700 -30820 3760 -29960
rect 5300 -29980 5360 -27350
rect 5500 -27400 5560 -23470
rect 5600 -27500 5660 -23420
rect 5700 -27350 5760 -23330
rect 5800 -27120 5860 -23280
rect 5900 -26840 5960 -23230
rect 6000 -26440 6060 -23230
rect 6100 -26410 6160 -23230
rect 6200 -26320 6260 -23230
rect 6300 -26300 6360 -23230
rect 6400 -26340 6460 -23230
rect 6500 -26390 6560 -23230
rect 6600 -26430 6660 -23230
rect 6700 -26460 6760 -23240
rect 6800 -26470 6860 -23290
rect 6900 -26470 6960 -23320
rect 7000 -26470 7060 -23320
rect 7100 -26470 7160 -23320
rect 7200 -26470 7260 -23300
rect 7300 -26470 7360 -23250
rect 7400 -26480 7460 -23150
rect 6000 -27290 6060 -27020
rect 6100 -27430 6160 -26620
rect 3800 -30820 3860 -30010
rect 5400 -30030 5460 -27540
rect 3900 -30820 3960 -30060
rect 5500 -30080 5560 -27720
rect 5700 -27820 5760 -27760
rect 4000 -30820 4060 -30100
rect 5600 -30120 5660 -27890
rect 4100 -30830 4160 -30150
rect 5700 -30170 5760 -27880
rect 1400 -38430 1460 -31490
rect 1500 -38350 1560 -31500
rect 1600 -38270 1660 -31500
rect 1700 -38210 1760 -31500
rect 1800 -38110 1860 -31500
rect 1900 -38060 1960 -31500
rect 2000 -37990 2060 -31490
rect 2100 -37900 2160 -31520
rect 2700 -31820 2760 -31760
rect 2200 -37840 2260 -31880
rect 2300 -37750 2360 -31880
rect 2400 -37690 2460 -31880
rect 2500 -37630 2560 -31880
rect 2600 -37540 2660 -31880
rect 2700 -37480 2760 -31880
rect 2800 -37420 2860 -31500
rect 2900 -37320 2960 -31500
rect 3000 -37260 3060 -31500
rect 3100 -37180 3160 -31500
rect 3200 -37110 3260 -31500
rect 3300 -37050 3360 -31500
rect 3400 -36960 3460 -31500
rect 3500 -36900 3560 -31500
rect 3600 -36820 3660 -31500
rect 3700 -36750 3760 -31500
rect 3800 -36680 3860 -31500
rect 3900 -36610 3960 -31500
rect 4000 -36530 4060 -31500
rect 4100 -36470 4160 -31490
rect 4200 -36370 4260 -30190
rect 5800 -30210 5860 -27480
rect 4300 -36310 4360 -30240
rect 5900 -30260 5960 -27480
rect 6200 -27580 6260 -26500
rect 4400 -36250 4460 -30290
rect 6000 -30300 6060 -27580
rect 4500 -36160 4560 -30330
rect 6100 -30350 6160 -27720
rect 6300 -27770 6360 -26500
rect 7500 -26510 7560 -23080
rect 7600 -26520 7660 -23030
rect 7700 -26520 7760 -22930
rect 7800 -24120 7860 -22700
rect 7900 -24180 7960 -21100
rect 8000 -24250 8060 -21140
rect 8100 -24250 8160 -21140
rect 8200 -24230 8260 -21130
rect 8300 -24180 8360 -21100
rect 8400 -24080 8460 -21100
rect 8500 -23980 8560 -21100
rect 8600 -23900 8660 -21080
rect 8700 -23830 8760 -21050
rect 8800 -23770 8860 -21020
rect 8900 -23670 8960 -20950
rect 9000 -23520 9060 -20890
rect 9100 -23120 9160 -19700
rect 9300 -19750 9360 0
rect 9400 -19890 9460 0
rect 9200 -20850 9260 -19890
rect 9300 -20360 9360 -20070
rect 9300 -20830 9360 -20750
rect 9200 -22680 9260 -21070
rect 9400 -21400 9460 -20540
rect 9500 -21830 9560 0
rect 9600 -22060 9660 0
rect 7800 -26510 7860 -24330
rect 7900 -26550 7960 -24410
rect 8000 -26560 8060 -24450
rect 8100 -26560 8160 -24450
rect 8200 -26560 8260 -24440
rect 8300 -26560 8360 -24380
rect 8400 -26560 8460 -24320
rect 8500 -26570 8560 -24220
rect 4600 -36100 4660 -30380
rect 6200 -30410 6260 -27870
rect 6400 -27910 6460 -26580
rect 8600 -26600 8660 -24120
rect 8700 -26600 8760 -24060
rect 4700 -36040 4760 -30430
rect 4800 -35940 4860 -30480
rect 4900 -35890 4960 -30520
rect 5000 -35820 5060 -30570
rect 5100 -35740 5160 -30620
rect 5200 -35680 5260 -30670
rect 5300 -35600 5360 -30710
rect 5400 -35560 5460 -30760
rect 5500 -35480 5560 -30810
rect 5600 -35430 5660 -30850
rect 5700 -35360 5760 -30900
rect 5800 -35310 5860 -30950
rect 5900 -35240 5960 -30990
rect 6000 -35180 6060 -31040
rect 6100 -35130 6160 -31090
rect 6200 -35070 6260 -31120
rect 6300 -35010 6360 -28050
rect 6500 -28100 6560 -26600
rect 8800 -26610 8860 -23980
rect 6400 -34960 6460 -28320
rect 6600 -28370 6660 -26620
rect 6500 -34900 6560 -28510
rect 6700 -28560 6760 -26630
rect 8900 -26650 8960 -23910
rect 9000 -26650 9060 -23810
rect 9100 -26650 9160 -23670
rect 9200 -26650 9260 -23390
rect 9300 -26650 9360 -22900
rect 9400 -26040 9460 -22360
rect 9500 -23250 9560 -22200
rect 9700 -22240 9760 0
rect 9600 -23320 9660 -22380
rect 9800 -22420 9860 0
rect 9900 -5480 9960 0
rect 10000 -4860 10060 0
rect 10100 -4800 10160 0
rect 10200 -4880 10260 0
rect 10300 -4940 10360 0
rect 10400 -5000 10460 0
rect 10500 -5050 10560 0
rect 9500 -25600 9560 -23670
rect 9700 -23850 9760 -22610
rect 9900 -22620 9960 -7310
rect 10100 -7750 10160 -5050
rect 6600 -34840 6660 -28690
rect 6800 -28790 6860 -26670
rect 6700 -34790 6760 -29020
rect 6900 -29110 6960 -26670
rect 6800 -34740 6860 -29290
rect 7000 -29340 7060 -26670
rect 6900 -34690 6960 -29510
rect 7100 -29560 7160 -26670
rect 7000 -34650 7060 -29790
rect 7200 -29830 7260 -26670
rect 7100 -34600 7160 -29980
rect 7300 -30030 7360 -26670
rect 7200 -34550 7260 -30160
rect 7400 -30250 7460 -26670
rect 7300 -34520 7360 -30400
rect 7500 -30450 7560 -26700
rect 7400 -34470 7460 -30670
rect 7600 -30720 7660 -26710
rect 7500 -34420 7560 -30850
rect 7700 -30910 7760 -26710
rect 7600 -34390 7660 -31040
rect 7800 -31090 7860 -26710
rect 7700 -34340 7760 -31270
rect 7900 -31280 7960 -26710
rect 8000 -31420 8060 -26710
rect 7800 -34290 7860 -31420
rect 7900 -34260 7960 -31560
rect 8100 -31570 8160 -26750
rect 8000 -34210 8060 -31700
rect 8200 -31710 8260 -26760
rect 8300 -31850 8360 -26750
rect 8100 -34170 8160 -31850
rect 8400 -31950 8460 -26750
rect 8200 -34130 8260 -31990
rect 8500 -32030 8560 -26760
rect 8600 -31890 8660 -26800
rect 8700 -31350 8760 -26800
rect 8800 -31310 8860 -26800
rect 8900 -31410 8960 -26840
rect 8700 -31470 8760 -31410
rect 9000 -31550 9060 -26840
rect 9100 -31650 9160 -26840
rect 8300 -34090 8360 -32100
rect 8400 -34050 8460 -32190
rect 8500 -34030 8560 -32290
rect 8600 -33990 8660 -32390
rect 8700 -33960 8760 -32380
rect 8800 -33920 8860 -31710
rect 8900 -33890 8960 -31690
rect 9200 -31750 9260 -26840
rect 9000 -33860 9060 -31790
rect 9300 -31850 9360 -26840
rect 9100 -33830 9160 -31890
rect 9400 -31950 9460 -26840
rect 9200 -33810 9260 -31990
rect 9500 -32050 9560 -26840
rect 9300 -33780 9360 -32090
rect 9600 -32150 9660 -25820
rect 9400 -33740 9460 -32190
rect 9700 -32250 9760 -24460
rect 9800 -24780 9860 -22800
rect 10000 -22890 10060 -8100
rect 10200 -8370 10260 -5090
rect 10600 -5100 10660 0
rect 10700 -5140 10760 0
rect 10300 -5570 10360 -5150
rect 10800 -5180 10860 0
rect 10400 -5700 10460 -5200
rect 10900 -5230 10960 0
rect 11000 -5250 11060 0
rect 10500 -5800 10560 -5250
rect 11100 -5280 11160 0
rect 10200 -8540 10260 -8480
rect 9900 -24770 9960 -23020
rect 10100 -23070 10160 -8780
rect 10300 -8950 10360 -5840
rect 10600 -5900 10660 -5300
rect 11200 -5320 11260 0
rect 11300 -5330 11360 0
rect 10700 -6000 10760 -5330
rect 11400 -5370 11460 0
rect 11500 -5360 11560 0
rect 10800 -6100 10860 -5380
rect 11600 -5400 11660 0
rect 11700 -5410 11760 0
rect 10500 -6850 10560 -6100
rect 10400 -7690 10460 -7630
rect 10200 -19630 10260 -9140
rect 10400 -9320 10460 -7750
rect 10600 -7990 10660 -6140
rect 10900 -6200 10960 -5430
rect 11800 -5440 11860 0
rect 11900 -5450 11960 0
rect 10300 -19600 10360 -9540
rect 10500 -9670 10560 -8260
rect 10700 -8530 10760 -6240
rect 10400 -9940 10460 -9880
rect 10400 -13070 10460 -10000
rect 10600 -10080 10660 -8750
rect 10800 -8980 10860 -6340
rect 11000 -6350 11060 -5460
rect 11100 -6440 11160 -5480
rect 12000 -5490 12060 0
rect 12100 -5490 12160 0
rect 10500 -12410 10560 -10220
rect 10700 -10310 10760 -9200
rect 10900 -9330 10960 -6490
rect 11200 -6550 11260 -5520
rect 10900 -9460 10960 -9400
rect 10600 -11840 10660 -10450
rect 10800 -10540 10860 -9560
rect 11000 -9650 11060 -6580
rect 11300 -6690 11360 -5520
rect 12200 -5530 12260 0
rect 12300 -5540 12360 0
rect 10700 -10750 10760 -10690
rect 10900 -10780 10960 -9830
rect 11100 -9970 11160 -6690
rect 10700 -11480 10760 -10810
rect 10800 -11240 10860 -10950
rect 11000 -11050 11060 -10110
rect 11200 -10210 11260 -6780
rect 11400 -6790 11460 -5560
rect 11500 -6890 11560 -5560
rect 12400 -5580 12460 0
rect 11300 -10300 11360 -6930
rect 11600 -7030 11660 -5600
rect 11400 -8160 11460 -7030
rect 11500 -8100 11560 -7170
rect 11700 -7180 11760 -5600
rect 12500 -5610 12560 0
rect 12600 -5640 12660 0
rect 11600 -8100 11660 -7270
rect 11800 -7280 11860 -5640
rect 11700 -8150 11760 -7410
rect 11900 -7420 11960 -5650
rect 12700 -5670 12760 0
rect 12000 -7560 12060 -5670
rect 11800 -8200 11860 -7560
rect 12100 -7700 12160 -5690
rect 12800 -5700 12860 0
rect 11400 -8280 11460 -8220
rect 11900 -8250 11960 -7700
rect 12000 -8300 12060 -7840
rect 12200 -7890 12260 -5700
rect 12900 -5710 12960 0
rect 12300 -8030 12360 -5740
rect 13000 -5750 13060 0
rect 13100 -5760 13160 0
rect 11400 -9040 11460 -8940
rect 11400 -10100 11460 -9100
rect 11600 -9120 11660 -8310
rect 12100 -8350 12160 -8030
rect 11500 -10030 11560 -9310
rect 11700 -9350 11760 -8350
rect 11600 -9970 11660 -9530
rect 11800 -9540 11860 -8400
rect 12200 -8410 12260 -8180
rect 12400 -8230 12460 -5780
rect 13200 -5800 13260 0
rect 13300 -5810 13360 0
rect 12300 -8430 12360 -8350
rect 12500 -8370 12560 -5820
rect 11700 -9930 11760 -9670
rect 11900 -9680 11960 -8450
rect 11800 -9930 11860 -9860
rect 12000 -9870 12060 -8500
rect 12600 -8550 12660 -5820
rect 13400 -5840 13460 0
rect 13500 -5850 13560 0
rect 11500 -10330 11560 -10260
rect 11100 -11230 11160 -10420
rect 11300 -10530 11360 -10360
rect 11200 -11460 11260 -10660
rect 11400 -10750 11460 -10410
rect 11600 -10470 11660 -10180
rect 10700 -11600 10760 -11540
rect 10400 -15470 10460 -15410
rect 10600 -15640 10660 -13690
rect 10400 -19520 10460 -15770
rect 10600 -16170 10660 -15700
rect 10500 -19330 10560 -16700
rect 10700 -17150 10760 -12800
rect 10600 -18400 10660 -18070
rect 10600 -19570 10660 -19510
rect 10700 -19590 10760 -19020
rect 10800 -19550 10860 -12310
rect 10900 -19510 10960 -11980
rect 11000 -19490 11060 -11710
rect 11100 -19410 11160 -11610
rect 11200 -19360 11260 -11520
rect 11300 -19290 11360 -10930
rect 11500 -11020 11560 -10610
rect 11700 -10620 11760 -10130
rect 11800 -10710 11860 -10100
rect 11600 -11160 11660 -10710
rect 11900 -10810 11960 -10080
rect 12000 -10850 12060 -10090
rect 12100 -10770 12160 -8560
rect 12200 -10580 12260 -8620
rect 12600 -8670 12660 -8610
rect 12300 -10440 12360 -8710
rect 12400 -10240 12460 -8850
rect 12700 -8870 12760 -5870
rect 13600 -5880 13660 0
rect 12500 -10110 12560 -9000
rect 12600 -9960 12660 -9100
rect 12800 -9140 12860 -5900
rect 13700 -5910 13760 0
rect 12700 -9830 12760 -9370
rect 12900 -9490 12960 -5910
rect 13800 -5930 13860 0
rect 13000 -9440 13060 -5950
rect 13100 -9290 13160 -5950
rect 13900 -5970 13960 0
rect 14000 -5990 14060 0
rect 13200 -9200 13260 -5990
rect 13300 -9050 13360 -6000
rect 14100 -6020 14160 0
rect 13400 -8950 13460 -6040
rect 14200 -6050 14260 0
rect 13500 -8800 13560 -6050
rect 13600 -8710 13660 -6080
rect 14300 -6100 14360 0
rect 13700 -8560 13760 -6110
rect 14400 -6120 14460 0
rect 13800 -8460 13860 -6130
rect 14500 -6150 14560 0
rect 13900 -8360 13960 -6170
rect 14000 -8300 14060 -6170
rect 14600 -6190 14660 0
rect 14100 -8210 14160 -6210
rect 14700 -6230 14760 0
rect 14200 -8110 14260 -6250
rect 14300 -8010 14360 -6270
rect 14800 -6280 14860 0
rect 14400 -7910 14460 -6310
rect 14900 -6330 14960 0
rect 14500 -7800 14560 -6350
rect 15000 -6380 15060 0
rect 14600 -7710 14660 -6390
rect 14700 -7600 14760 -6430
rect 15100 -6440 15160 0
rect 15200 -6440 15260 0
rect 15300 -6390 15360 0
rect 15400 -6320 15460 0
rect 15500 -6270 15560 0
rect 15600 -6220 15660 0
rect 15700 -6170 15760 0
rect 15800 -6120 15860 0
rect 15900 -6070 15960 0
rect 16000 -6020 16060 0
rect 16100 -5970 16160 0
rect 16200 -5930 16260 0
rect 16300 -5890 16360 0
rect 16400 -5840 16460 0
rect 16500 -5800 16560 0
rect 16600 -5760 16660 0
rect 16700 -5710 16760 0
rect 16800 -5680 16860 0
rect 16900 -5660 16960 0
rect 17000 -5620 17060 0
rect 17100 -5580 17160 0
rect 17200 -5580 17260 0
rect 17300 -5540 17360 0
rect 17400 -5520 17460 0
rect 17500 -5490 17560 0
rect 17600 -5460 17660 0
rect 17700 -5450 17760 0
rect 17800 -5420 17860 0
rect 17900 -5410 17960 0
rect 18000 -5400 18060 0
rect 18100 -5360 18160 0
rect 18200 -5360 18260 0
rect 18300 -5360 18360 0
rect 18400 -5340 18460 0
rect 18500 -5320 18560 0
rect 18600 -5320 18660 0
rect 18700 -5320 18760 0
rect 18800 -5320 18860 0
rect 18900 -5320 18960 0
rect 19000 -5320 19060 0
rect 19100 -5320 19160 0
rect 19200 -5320 19260 0
rect 19300 -5320 19360 0
rect 19400 -5320 19460 0
rect 19500 -5320 19560 0
rect 19600 -5320 19660 0
rect 19700 -5330 19760 0
rect 19800 -5370 19860 0
rect 19900 -5330 19960 0
rect 20000 -5320 20060 0
rect 20100 -5320 20160 0
rect 20200 -5290 20260 0
rect 20300 -5280 20360 0
rect 20400 -5280 20460 0
rect 20500 -5280 20560 0
rect 20600 -5270 20660 0
rect 20700 -5230 20760 0
rect 20800 -5230 20860 0
rect 20900 -5230 20960 0
rect 21000 -5230 21060 0
rect 21100 -5230 21160 0
rect 21200 -5230 21260 0
rect 21300 -5230 21360 0
rect 21400 -5230 21460 0
rect 21500 -5230 21560 0
rect 21600 -5230 21660 0
rect 21700 -5230 21760 0
rect 21800 -5230 21860 0
rect 21900 -5260 21960 0
rect 22000 -5280 22060 0
rect 22100 -5320 22160 0
rect 22200 -5320 22260 0
rect 22300 -5240 22360 0
rect 22400 -5100 22460 0
rect 22500 -4990 22560 0
rect 22600 -4860 22660 0
rect 22700 -4750 22760 0
rect 22800 -4610 22860 0
rect 22900 -4510 22960 0
rect 23000 -4410 23060 0
rect 23100 -4270 23160 0
rect 23200 -4170 23260 0
rect 23300 -4070 23360 0
rect 23400 -3970 23460 0
rect 23500 -3870 23560 0
rect 23600 -3770 23660 0
rect 23700 -3670 23760 0
rect 23800 -3570 23860 0
rect 23900 -3470 23960 0
rect 24000 -3370 24060 0
rect 24100 -3270 24160 0
rect 24200 -3170 24260 0
rect 24300 -3090 24360 0
rect 24400 -3020 24460 0
rect 24500 -3000 24560 0
rect 24600 -2930 24660 0
rect 14800 -7550 14860 -6480
rect 14900 -7450 14960 -6530
rect 15000 -7390 15060 -6580
rect 15100 -7320 15160 -6670
rect 11400 -12470 11460 -11200
rect 11500 -12110 11560 -11390
rect 11700 -11430 11760 -10850
rect 11800 -11330 11860 -10950
rect 11900 -11150 11960 -11050
rect 11600 -11880 11660 -11580
rect 11600 -12450 11660 -12290
rect 11400 -12630 11460 -12530
rect 11400 -12750 11460 -12690
rect 11500 -14020 11560 -13090
rect 11400 -19240 11460 -14160
rect 11500 -19160 11560 -14230
rect 11600 -19070 11660 -12510
rect 11700 -19140 11760 -12010
rect 10000 -24840 10060 -23210
rect 10200 -23310 10260 -19760
rect 9500 -33700 9560 -32290
rect 9800 -32350 9860 -24870
rect 10100 -24900 10160 -23490
rect 10300 -23540 10360 -19820
rect 9600 -33670 9660 -32390
rect 9900 -32430 9960 -24990
rect 10200 -25000 10260 -23670
rect 10400 -23770 10460 -19790
rect 9700 -33650 9760 -32490
rect 10000 -32500 10060 -25050
rect 10300 -25100 10360 -23900
rect 10500 -23990 10560 -19790
rect 10400 -24210 10460 -24150
rect 10600 -24260 10660 -19790
rect 10100 -32570 10160 -25140
rect 10400 -25200 10460 -24270
rect 9800 -33600 9860 -32580
rect 10200 -32640 10260 -25240
rect 10500 -25300 10560 -24410
rect 10700 -24500 10760 -19770
rect 9900 -33560 9960 -32640
rect 10300 -32720 10360 -25340
rect 10600 -25400 10660 -24640
rect 10800 -24730 10860 -19750
rect 10700 -25430 10760 -24910
rect 10900 -24960 10960 -19710
rect 10900 -25080 10960 -25020
rect 10000 -33520 10060 -32720
rect 10400 -32770 10460 -25440
rect 10800 -25480 10860 -25190
rect 11000 -25280 11060 -19680
rect 10100 -33490 10160 -32800
rect 10500 -32830 10560 -25540
rect 10900 -25550 10960 -25410
rect 11100 -25460 11160 -19630
rect 10200 -33460 10260 -32860
rect 10600 -32890 10660 -25640
rect 11200 -25650 11260 -19570
rect 10700 -32910 10760 -25740
rect 10300 -33410 10360 -32920
rect 10800 -32950 10860 -25840
rect 10900 -32960 10960 -25940
rect 11000 -32950 11060 -26040
rect 11300 -26050 11360 -19510
rect 10400 -33380 10460 -32970
rect 11100 -33000 11160 -26110
rect 11400 -26150 11460 -19450
rect 10500 -33350 10560 -33040
rect 10600 -33310 10660 -33090
rect 10700 -33300 10760 -33110
rect 10800 -33260 10860 -33150
rect 10900 -33220 10960 -33150
rect 11000 -33190 11060 -33130
rect 11100 -33170 11160 -33070
rect 11200 -33130 11260 -26200
rect 11500 -26250 11560 -19410
rect 11700 -19490 11760 -19280
rect 11300 -33110 11360 -26300
rect 11600 -26350 11660 -19670
rect 11800 -19770 11860 -11780
rect 11400 -33080 11460 -26400
rect 11500 -33040 11560 -26490
rect 11700 -26500 11760 -19950
rect 11900 -20040 11960 -11560
rect 11800 -26640 11860 -20220
rect 12000 -20270 12060 -11290
rect 12100 -14000 12160 -11140
rect 12200 -13940 12260 -10950
rect 12100 -14130 12160 -14070
rect 11600 -33020 11660 -26640
rect 11900 -26740 11960 -20410
rect 12100 -20460 12160 -14250
rect 12300 -14440 12360 -10720
rect 12200 -20600 12260 -14620
rect 12400 -14670 12460 -10580
rect 11700 -32990 11760 -26770
rect 11800 -32960 11860 -26880
rect 12000 -26890 12060 -20600
rect 12300 -20790 12360 -14800
rect 12500 -14850 12560 -10390
rect 12100 -26980 12160 -20790
rect 12400 -20930 12460 -14990
rect 12600 -15010 12660 -10250
rect 12700 -14920 12760 -10110
rect 12800 -14590 12860 -9960
rect 12900 -14410 12960 -9820
rect 13000 -14220 13060 -9680
rect 13100 -14150 13160 -9530
rect 13200 -14380 13260 -9430
rect 13300 -14470 13360 -9330
rect 11900 -32940 11960 -27020
rect 12000 -32910 12060 -27120
rect 12200 -27130 12260 -20930
rect 12500 -21070 12560 -15220
rect 12300 -27270 12360 -21070
rect 12100 -32870 12160 -27270
rect 12400 -27410 12460 -21210
rect 12600 -21220 12660 -15360
rect 12700 -21360 12760 -15440
rect 12200 -32860 12260 -27410
rect 12300 -32820 12360 -27550
rect 12500 -27560 12560 -21360
rect 12600 -27700 12660 -21450
rect 12800 -21460 12860 -15100
rect 12900 -21600 12960 -14830
rect 12400 -32780 12460 -27700
rect 12500 -32740 12560 -27880
rect 12700 -27890 12760 -21600
rect 12800 -28030 12860 -21740
rect 13000 -21750 13060 -14540
rect 12600 -32720 12660 -28030
rect 12900 -28170 12960 -21840
rect 13100 -21850 13160 -14530
rect 13400 -14570 13460 -9190
rect 13200 -21950 13260 -14610
rect 13500 -14640 13560 -9090
rect 12700 -32690 12760 -28170
rect 12800 -32660 12860 -28360
rect 13000 -28410 13060 -21980
rect 13300 -22050 13360 -14710
rect 13600 -14720 13660 -8950
rect 13700 -14780 13760 -8850
rect 13400 -18090 13460 -14790
rect 13800 -14830 13860 -8700
rect 13500 -17900 13560 -14870
rect 13900 -14900 13960 -8600
rect 13600 -17630 13660 -14930
rect 14000 -14950 14060 -8500
rect 13700 -17500 13760 -14990
rect 14100 -15010 14160 -8430
rect 14200 -15030 14260 -8340
rect 13800 -17430 13860 -15040
rect 14300 -15080 14360 -8250
rect 13900 -17320 13960 -15100
rect 14400 -15130 14460 -8130
rect 14000 -17230 14060 -15160
rect 14500 -15190 14560 -8050
rect 14100 -17130 14160 -15210
rect 14600 -15230 14660 -7950
rect 14700 -15190 14760 -7850
rect 14800 -14860 14860 -7750
rect 14900 -14630 14960 -7680
rect 15000 -10360 15060 -7590
rect 15100 -10150 15160 -7540
rect 15100 -11960 15160 -10620
rect 15000 -14360 15060 -12360
rect 15200 -12670 15260 -6730
rect 15100 -13090 15160 -12940
rect 15300 -13030 15360 -6790
rect 15100 -13910 15160 -13150
rect 15400 -13740 15460 -6690
rect 14200 -17030 14260 -15230
rect 14300 -16970 14360 -15280
rect 14400 -16870 14460 -15330
rect 14500 -16820 14560 -15390
rect 14600 -16760 14660 -15410
rect 14700 -16700 14760 -15440
rect 14800 -16630 14860 -15360
rect 14900 -16580 14960 -15090
rect 15000 -16530 15060 -14770
rect 15100 -16500 15160 -14540
rect 15200 -16450 15260 -14180
rect 15300 -16420 15360 -13930
rect 15500 -14060 15560 -6650
rect 15400 -16400 15460 -14240
rect 15600 -14330 15660 -6570
rect 15500 -16320 15560 -14600
rect 15700 -14650 15760 -6520
rect 15600 -16290 15660 -14790
rect 15800 -14890 15860 -6480
rect 15700 -16300 15760 -15020
rect 15900 -15070 15960 -6430
rect 15800 -16360 15860 -15210
rect 16000 -15250 16060 -6380
rect 15900 -16450 15960 -15440
rect 16100 -15490 16160 -6300
rect 16000 -16460 16060 -15620
rect 16200 -15670 16260 -6260
rect 16300 -15810 16360 -6220
rect 16100 -16500 16160 -15810
rect 16200 -16580 16260 -15960
rect 16400 -15970 16460 -6170
rect 16500 -16020 16560 -6130
rect 16600 -15500 16660 -6080
rect 16700 -15430 16760 -6040
rect 16800 -15580 16860 -6000
rect 16900 -15720 16960 -5960
rect 17000 -15860 17060 -5920
rect 16300 -16670 16360 -16100
rect 16700 -16220 16760 -15930
rect 15200 -17120 15260 -17060
rect 13100 -28320 13160 -22090
rect 13400 -22150 13460 -18340
rect 13200 -28200 13260 -22190
rect 13500 -22290 13560 -18330
rect 13300 -28170 13360 -22290
rect 13600 -22350 13660 -18280
rect 12900 -32650 12960 -28590
rect 13100 -28690 13160 -28380
rect 13400 -28390 13460 -22430
rect 13700 -22450 13760 -18200
rect 13000 -32610 13060 -28860
rect 13200 -29000 13260 -28460
rect 13500 -28470 13560 -22480
rect 13800 -22510 13860 -18180
rect 13600 -28550 13660 -22590
rect 13900 -22600 13960 -18400
rect 13300 -29150 13360 -28590
rect 13100 -32600 13160 -29250
rect 13200 -32560 13260 -29720
rect 13300 -32550 13360 -30020
rect 13400 -32520 13460 -30000
rect 13500 -32490 13560 -28810
rect 13600 -32460 13660 -28840
rect 13700 -29370 13760 -22670
rect 14000 -22700 14060 -18580
rect 13800 -28660 13860 -22740
rect 14100 -22760 14160 -18540
rect 14200 -18680 14260 -18180
rect 14300 -18630 14360 -17950
rect 14400 -18650 14460 -17760
rect 14500 -18720 14560 -17620
rect 13900 -28390 13960 -22840
rect 14200 -22850 14260 -18750
rect 14600 -18810 14660 -17520
rect 14300 -22900 14360 -18830
rect 14000 -28110 14060 -22900
rect 14400 -22940 14460 -18860
rect 14100 -27840 14160 -22970
rect 14500 -22990 14560 -18960
rect 14600 -23010 14660 -18970
rect 14700 -22930 14760 -17420
rect 14800 -19000 14860 -17350
rect 14900 -18380 14960 -17260
rect 15000 -18190 15060 -17230
rect 15100 -18040 15160 -17330
rect 15300 -17390 15360 -17010
rect 15200 -17900 15260 -17570
rect 15300 -17800 15360 -17610
rect 15400 -17700 15460 -16970
rect 15500 -17640 15560 -16920
rect 15600 -17580 15660 -16880
rect 15700 -17540 15760 -16840
rect 15800 -17500 15860 -16830
rect 15900 -17470 15960 -16830
rect 16000 -17460 16060 -16830
rect 16100 -17430 16160 -16830
rect 16400 -16910 16460 -16240
rect 16200 -17420 16260 -16910
rect 16500 -17060 16560 -16380
rect 16300 -17420 16360 -17060
rect 16400 -17460 16460 -17200
rect 16600 -17210 16660 -16530
rect 16500 -17460 16560 -17320
rect 16600 -17470 16660 -17270
rect 16700 -17510 16760 -16570
rect 16800 -17550 16860 -15880
rect 17100 -15960 17160 -5890
rect 16900 -17600 16960 -16000
rect 17200 -16060 17260 -5860
rect 15000 -18710 15060 -18550
rect 14800 -22830 14860 -19080
rect 15000 -19170 15060 -18770
rect 15000 -19350 15060 -19230
rect 14900 -22730 14960 -19530
rect 15100 -19620 15160 -18330
rect 15000 -22630 15060 -19760
rect 15200 -19770 15260 -18140
rect 15100 -22490 15160 -19910
rect 15300 -19950 15360 -18040
rect 15400 -20050 15460 -17940
rect 15500 -18040 15560 -17850
rect 15600 -17990 15660 -17780
rect 15200 -22340 15260 -20090
rect 15500 -20150 15560 -18130
rect 15700 -18180 15760 -17730
rect 15600 -20250 15660 -18310
rect 15800 -18370 15860 -17700
rect 15900 -18500 15960 -17660
rect 15300 -22250 15360 -20320
rect 15700 -20330 15760 -18500
rect 16000 -18650 16060 -17660
rect 15800 -20380 15860 -18650
rect 16100 -18830 16160 -17620
rect 15900 -20420 15960 -18830
rect 16000 -20470 16060 -18970
rect 16200 -18980 16260 -17620
rect 16300 -19120 16360 -17610
rect 15400 -22100 15460 -20470
rect 16100 -20510 16160 -19120
rect 16400 -19270 16460 -17640
rect 17000 -17650 17060 -16100
rect 17300 -16160 17360 -5820
rect 16200 -19860 16260 -19270
rect 16500 -19370 16560 -17660
rect 16300 -19810 16360 -19400
rect 16600 -19450 16660 -17670
rect 17100 -17700 17160 -16200
rect 17400 -16260 17460 -5780
rect 16700 -19500 16760 -17710
rect 16800 -17910 16860 -17750
rect 17200 -17770 17260 -16300
rect 17500 -16330 17560 -5750
rect 16900 -17900 16960 -17800
rect 16800 -19510 16860 -18030
rect 17000 -18130 17060 -17850
rect 17300 -17860 17360 -16400
rect 17600 -16420 17660 -5730
rect 16900 -19510 16960 -18350
rect 17100 -18450 17160 -17920
rect 17400 -17960 17460 -16490
rect 17700 -16500 17760 -5720
rect 17000 -19510 17060 -18630
rect 17200 -18720 17260 -18000
rect 17500 -18060 17560 -16560
rect 17800 -16570 17860 -5690
rect 17900 -16640 17960 -5680
rect 17100 -19490 17160 -18900
rect 17300 -19160 17360 -18100
rect 17600 -18200 17660 -16650
rect 16400 -19790 16460 -19510
rect 16500 -19770 16560 -19580
rect 16600 -19730 16660 -19650
rect 16200 -20550 16260 -19960
rect 16300 -20550 16360 -20010
rect 16400 -20590 16460 -19990
rect 16500 -20600 16560 -19960
rect 16600 -20600 16660 -19920
rect 16700 -20570 16760 -19880
rect 16800 -20550 16860 -19850
rect 16900 -20510 16960 -19840
rect 17000 -20490 17060 -19800
rect 17100 -20440 17160 -19730
rect 17200 -20390 17260 -19630
rect 17300 -20330 17360 -19350
rect 17400 -20230 17460 -18200
rect 17700 -18340 17760 -16710
rect 18000 -16720 18060 -5650
rect 18100 -16760 18160 -5650
rect 17500 -20130 17560 -18350
rect 17600 -19990 17660 -18530
rect 17800 -18580 17860 -16770
rect 18200 -16810 18260 -5600
rect 18300 -16810 18360 -5600
rect 18400 -16810 18460 -5590
rect 18500 -16700 18560 -5580
rect 18600 -16550 18660 -5690
rect 18700 -16460 18760 -5700
rect 18800 -11170 18860 -5740
rect 18900 -11140 18960 -5730
rect 19000 -11380 19060 -5740
rect 19100 -6130 19160 -5780
rect 19200 -6060 19260 -5780
rect 19300 -6020 19360 -5790
rect 19400 -5980 19460 -5820
rect 19500 -5940 19560 -5820
rect 19600 -5930 19660 -5870
rect 18800 -16320 18860 -11410
rect 18900 -16070 18960 -11690
rect 19100 -11740 19160 -6300
rect 19200 -11880 19260 -6270
rect 19000 -15850 19060 -12000
rect 19300 -12070 19360 -6230
rect 19400 -12250 19460 -6180
rect 19100 -15580 19160 -12410
rect 19500 -12440 19560 -6150
rect 19300 -12760 19360 -12490
rect 19200 -15000 19260 -13130
rect 19400 -13520 19460 -12570
rect 19600 -12630 19660 -6120
rect 19400 -13670 19460 -13590
rect 19400 -13940 19460 -13880
rect 19400 -14480 19460 -14420
rect 19400 -14750 19460 -14590
rect 19400 -14920 19460 -14840
rect 19200 -15210 19260 -15060
rect 17700 -19760 17760 -18710
rect 17900 -18850 17960 -16870
rect 18000 -18920 18060 -16920
rect 18100 -18620 18160 -16970
rect 18200 -18430 18260 -17010
rect 18300 -18340 18360 -17050
rect 18400 -18290 18460 -17020
rect 18500 -18250 18560 -17050
rect 18600 -18290 18660 -16830
rect 18700 -18340 18760 -16700
rect 18800 -18490 18860 -16590
rect 18900 -18630 18960 -16450
rect 19000 -18640 19060 -16260
rect 19100 -18550 19160 -16030
rect 19200 -18580 19260 -15710
rect 19300 -17290 19360 -15440
rect 19400 -17060 19460 -14980
rect 19500 -16880 19560 -12760
rect 19700 -12770 19760 -6080
rect 19800 -12960 19860 -6070
rect 19600 -16730 19660 -12960
rect 19900 -13100 19960 -6020
rect 19700 -15330 19760 -13100
rect 20000 -13240 20060 -5990
rect 19800 -15280 19860 -13240
rect 20100 -13390 20160 -5950
rect 19900 -15240 19960 -13430
rect 20000 -15190 20060 -13570
rect 20200 -13580 20260 -5910
rect 20100 -15110 20160 -13670
rect 20300 -13680 20360 -5880
rect 20400 -13750 20460 -5850
rect 20500 -13340 20560 -5820
rect 20600 -13310 20660 -5790
rect 20700 -13410 20760 -5770
rect 20500 -13520 20560 -13460
rect 20800 -13470 20860 -5730
rect 20900 -13520 20960 -5710
rect 21000 -13550 21060 -5690
rect 21100 -7700 21160 -5650
rect 21200 -7480 21260 -5650
rect 21300 -7240 21360 -5620
rect 21400 -7060 21460 -5600
rect 21500 -6870 21560 -5600
rect 21600 -6550 21660 -5600
rect 21700 -6320 21760 -5570
rect 21800 -6130 21860 -5560
rect 21900 -5900 21960 -5560
rect 22000 -5670 22060 -5570
rect 21300 -7840 21360 -7650
rect 21100 -13600 21160 -8010
rect 20200 -15040 20260 -13810
rect 20300 -15050 20360 -13960
rect 20700 -14030 20760 -13630
rect 21200 -13650 21260 -8020
rect 21300 -8770 21360 -7910
rect 21400 -8760 21460 -7420
rect 21500 -8820 21560 -7190
rect 21600 -7950 21660 -7000
rect 21700 -7670 21760 -6770
rect 21800 -7400 21860 -6450
rect 21900 -7170 21960 -6270
rect 22000 -6890 22060 -6040
rect 22100 -6660 22160 -5850
rect 22200 -6470 22260 -5660
rect 22300 -6290 22360 -5530
rect 22400 -6140 22460 -5380
rect 22500 -6000 22560 -5230
rect 22600 -5900 22660 -5140
rect 22700 -5760 22760 -4990
rect 22800 -5610 22860 -4890
rect 22900 -5510 22960 -4760
rect 23000 -5330 23060 -4650
rect 23100 -5140 23160 -4550
rect 23200 -5040 23260 -4410
rect 23300 -4860 23360 -4310
rect 23400 -4750 23460 -4210
rect 23500 -4610 23560 -4110
rect 23600 -4510 23660 -4010
rect 23700 -4360 23760 -3910
rect 23800 -4260 23860 -3810
rect 23900 -4170 23960 -3710
rect 24000 -4070 24060 -3610
rect 24100 -4000 24160 -3510
rect 24200 -3950 24260 -3410
rect 24300 -3680 24360 -3310
rect 24400 -3640 24460 -3250
rect 24300 -3900 24360 -3740
rect 21800 -7930 21860 -7850
rect 21600 -8070 21660 -8010
rect 21700 -8540 21760 -8260
rect 21300 -13680 21360 -8910
rect 21600 -8920 21660 -8690
rect 20400 -15020 20460 -14060
rect 20500 -14980 20560 -14140
rect 20600 -14900 20660 -14180
rect 20700 -14850 20760 -14130
rect 20800 -14830 20860 -13680
rect 21400 -13730 21460 -8970
rect 21700 -9020 21760 -8650
rect 20900 -14780 20960 -13730
rect 21000 -14750 21060 -13750
rect 21500 -13760 21560 -9060
rect 21800 -9120 21860 -7990
rect 21600 -13810 21660 -9170
rect 21900 -9220 21960 -7570
rect 21100 -14720 21160 -13810
rect 21700 -13850 21760 -9260
rect 22000 -9320 22060 -7300
rect 21200 -14680 21260 -13860
rect 21300 -14640 21360 -13880
rect 21800 -13890 21860 -9360
rect 22100 -9420 22160 -7070
rect 21900 -13920 21960 -9460
rect 21400 -14590 21460 -13930
rect 22000 -13970 22060 -9560
rect 22200 -9570 22260 -6800
rect 22300 -8500 22360 -6610
rect 22400 -8140 22460 -6470
rect 22500 -7820 22560 -6270
rect 22600 -7550 22660 -6140
rect 22700 -7410 22760 -6040
rect 22800 -7270 22860 -5900
rect 22900 -7160 22960 -5750
rect 23000 -7150 23060 -5600
rect 23100 -7200 23160 -5470
rect 22600 -7670 22660 -7610
rect 22300 -8690 22360 -8630
rect 22500 -9300 22560 -8320
rect 22300 -9700 22360 -9300
rect 22400 -9680 22460 -9440
rect 21500 -14590 21560 -13970
rect 22100 -13990 22160 -9700
rect 22500 -9710 22560 -9480
rect 22600 -9790 22660 -8010
rect 21600 -14550 21660 -14000
rect 22200 -14020 22260 -9800
rect 22700 -9850 22760 -7780
rect 22800 -9310 22860 -7550
rect 22900 -9280 22960 -7400
rect 23000 -9400 23060 -7390
rect 23200 -7520 23260 -5280
rect 22800 -9900 22860 -9440
rect 23100 -9510 23160 -7740
rect 23300 -8050 23360 -5130
rect 23400 -8060 23460 -5030
rect 23500 -7970 23560 -4890
rect 23600 -7900 23660 -4750
rect 23700 -7850 23760 -4650
rect 23800 -7800 23860 -4500
rect 23900 -7730 23960 -4400
rect 24000 -7630 24060 -4300
rect 24100 -7720 24160 -4200
rect 22900 -9980 22960 -9590
rect 23200 -9610 23260 -8410
rect 23300 -9710 23360 -8430
rect 23400 -9760 23460 -8260
rect 21700 -14550 21760 -14040
rect 22300 -14070 22360 -9990
rect 22600 -10140 22660 -9990
rect 21800 -14530 21860 -14090
rect 22400 -14110 22460 -10140
rect 21900 -14500 21960 -14120
rect 22500 -14150 22560 -10280
rect 22700 -10290 22760 -10050
rect 23000 -10060 23060 -9820
rect 23500 -9860 23560 -8200
rect 23100 -10060 23160 -10000
rect 23300 -10060 23360 -9920
rect 23600 -9960 23660 -8130
rect 22800 -10430 22860 -10130
rect 22000 -14470 22060 -14150
rect 22600 -14180 22660 -10440
rect 22100 -14460 22160 -14190
rect 22700 -14200 22760 -10610
rect 22900 -10620 22960 -10200
rect 22200 -14460 22260 -14230
rect 22800 -14240 22860 -10750
rect 23000 -10760 23060 -10260
rect 23400 -10290 23460 -10000
rect 23700 -10020 23760 -8050
rect 22900 -14240 22960 -10890
rect 23100 -10900 23160 -10360
rect 22300 -14460 22360 -14260
rect 23000 -14280 23060 -11040
rect 23200 -11050 23260 -10420
rect 23100 -14290 23160 -11180
rect 23300 -11190 23360 -10510
rect 23200 -14300 23260 -11320
rect 23400 -11330 23460 -10480
rect 22400 -14450 22460 -14310
rect 23300 -14330 23360 -11470
rect 23500 -11520 23560 -10090
rect 23800 -10120 23860 -8000
rect 23900 -10150 23960 -7970
rect 24000 -9590 24060 -8380
rect 24200 -8650 24260 -4150
rect 24300 -4210 24360 -4150
rect 24000 -10150 24060 -9840
rect 24100 -10010 24160 -9770
rect 24200 -9880 24260 -9490
rect 24300 -9650 24360 -4270
rect 24500 -5490 24560 -3230
rect 24700 -3360 24760 0
rect 24400 -9200 24460 -6000
rect 24600 -6740 24660 -3540
rect 24800 -3720 24860 0
rect 24500 -9520 24560 -9420
rect 23400 -14330 23460 -11610
rect 23600 -11660 23660 -10160
rect 23700 -11800 23760 -10260
rect 23500 -14330 23560 -11800
rect 23800 -11940 23860 -10320
rect 22500 -14420 22560 -14350
rect 22600 -14420 22660 -14360
rect 23600 -14370 23660 -11940
rect 23700 -14370 23760 -12090
rect 23900 -12130 23960 -10410
rect 24100 -10420 24160 -10300
rect 24200 -10520 24260 -10150
rect 23800 -14370 23860 -12270
rect 24000 -12280 24060 -10560
rect 24300 -10660 24360 -10010
rect 24100 -12420 24160 -10660
rect 24400 -10800 24460 -9780
rect 23900 -14370 23960 -12420
rect 24000 -14370 24060 -12600
rect 24200 -12610 24260 -10800
rect 24300 -12750 24360 -10940
rect 24500 -10950 24560 -9580
rect 24100 -14370 24160 -12750
rect 24400 -12890 24460 -11090
rect 24600 -11140 24660 -8360
rect 24200 -14370 24260 -12890
rect 24500 -13040 24560 -11230
rect 24700 -11280 24760 -4040
rect 24900 -4170 24960 0
rect 24800 -11420 24860 -4390
rect 25000 -4530 25060 0
rect 24300 -14370 24360 -13040
rect 24600 -13180 24660 -11420
rect 24400 -14370 24460 -13180
rect 24700 -13280 24760 -11560
rect 24900 -11610 24960 -4710
rect 25100 -4810 25160 0
rect 25000 -5040 25060 -4980
rect 25000 -11750 25060 -5100
rect 25200 -5210 25260 0
rect 24500 -14370 24560 -13280
rect 24800 -13420 24860 -11750
rect 25100 -11890 25160 -5350
rect 25300 -5440 25360 0
rect 24600 -14370 24660 -13420
rect 24900 -13610 24960 -11890
rect 24700 -14370 24760 -13610
rect 25000 -13750 25060 -12080
rect 25200 -12130 25260 -5620
rect 25400 -5670 25460 0
rect 25300 -5910 25360 -5850
rect 25500 -5940 25560 0
rect 24800 -14370 24860 -13750
rect 24900 -14330 24960 -13890
rect 25100 -13900 25160 -12260
rect 25300 -12270 25360 -5970
rect 25200 -14000 25260 -12410
rect 25000 -14320 25060 -14020
rect 25300 -14100 25360 -12480
rect 25100 -14200 25160 -14140
rect 25400 -14160 25460 -6210
rect 25600 -6310 25660 0
rect 22700 -14460 22760 -14400
rect 22800 -14460 22860 -14400
rect 23800 -14630 23860 -14570
rect 23900 -14640 23960 -14570
rect 24000 -14680 24060 -14570
rect 24100 -14710 24160 -14570
rect 24200 -15050 24260 -14570
rect 24300 -15180 24360 -14570
rect 19700 -15850 19760 -15530
rect 19700 -16630 19760 -16010
rect 19800 -16530 19860 -16080
rect 19900 -16430 19960 -15980
rect 20000 -16330 20060 -15930
rect 20100 -16280 20160 -15860
rect 20200 -16220 20260 -15810
rect 20300 -16170 20360 -15760
rect 20400 -16140 20460 -15710
rect 20500 -16110 20560 -15660
rect 20600 -16070 20660 -15610
rect 20700 -16060 20760 -15560
rect 20800 -16030 20860 -15530
rect 20900 -16030 20960 -15480
rect 21000 -16030 21060 -15440
rect 21100 -16030 21160 -15400
rect 21200 -16030 21260 -15390
rect 21300 -16030 21360 -15350
rect 21400 -16030 21460 -15350
rect 21500 -16070 21560 -15680
rect 21600 -16070 21660 -15740
rect 21700 -16110 21760 -15280
rect 21800 -16150 21860 -15270
rect 21900 -16180 21960 -15220
rect 19400 -17590 19460 -17520
rect 19400 -17710 19460 -17650
rect 19400 -18100 19460 -17840
rect 19300 -18550 19360 -18310
rect 19500 -18410 19560 -17190
rect 19600 -18590 19660 -17010
rect 17800 -19360 17860 -19160
rect 15500 -21950 15560 -20610
rect 15600 -21810 15660 -20760
rect 16000 -20770 16060 -20680
rect 15700 -21710 15760 -20810
rect 16100 -20830 16160 -20710
rect 16200 -20890 16260 -20750
rect 15800 -21570 15860 -20910
rect 16300 -20950 16360 -20750
rect 16400 -20990 16460 -20770
rect 16500 -21010 16560 -20790
rect 15900 -21380 15960 -21010
rect 16600 -21040 16660 -20780
rect 16000 -21240 16060 -21060
rect 16700 -21080 16760 -20750
rect 16800 -21080 16860 -20750
rect 16900 -21120 16960 -20720
rect 14200 -27560 14260 -23050
rect 14300 -27420 14360 -23100
rect 14400 -27280 14460 -23170
rect 14500 -27180 14560 -23220
rect 14600 -27070 14660 -23270
rect 14700 -26980 14760 -23210
rect 14800 -26900 14860 -23070
rect 14900 -26730 14960 -22970
rect 15000 -26580 15060 -22870
rect 15100 -26490 15160 -22770
rect 15200 -26340 15260 -22630
rect 15300 -26160 15360 -22480
rect 15400 -26020 15460 -22380
rect 15500 -25830 15560 -22240
rect 15600 -25640 15660 -22100
rect 15700 -25500 15760 -21950
rect 15800 -25350 15860 -21850
rect 15900 -24990 15960 -21700
rect 16000 -24810 16060 -21560
rect 16100 -24590 16160 -21370
rect 16200 -24590 16260 -21180
rect 16300 -24590 16360 -21140
rect 17000 -21150 17060 -20700
rect 17100 -21160 17160 -20640
rect 16400 -23930 16460 -21180
rect 17200 -21200 17260 -20590
rect 16500 -23440 16560 -21220
rect 16600 -23160 16660 -21230
rect 17300 -21240 17360 -20530
rect 17400 -21260 17460 -20470
rect 16700 -22940 16760 -21270
rect 16800 -22700 16860 -21280
rect 17500 -21290 17560 -20370
rect 17600 -21300 17660 -20270
rect 16900 -22560 16960 -21310
rect 17000 -22460 17060 -21330
rect 17700 -21340 17760 -20130
rect 17800 -21340 17860 -19930
rect 17100 -22400 17160 -21360
rect 17900 -21380 17960 -19660
rect 18000 -21380 18060 -19190
rect 17200 -22340 17260 -21400
rect 18100 -21420 18160 -19170
rect 18200 -21430 18260 -18970
rect 17300 -22300 17360 -21440
rect 17400 -22250 17460 -21450
rect 18300 -21470 18360 -18750
rect 18400 -21470 18460 -18660
rect 18500 -21470 18560 -18660
rect 17500 -22220 17560 -21490
rect 17600 -22190 17660 -21490
rect 18600 -21510 18660 -18720
rect 18700 -21510 18760 -18830
rect 18800 -21510 18860 -18900
rect 18900 -21510 18960 -18920
rect 19000 -21510 19060 -18920
rect 19100 -20450 19160 -18920
rect 19200 -20420 19260 -18880
rect 19300 -20470 19360 -18830
rect 19400 -20510 19460 -18680
rect 19500 -20480 19560 -18720
rect 19700 -18780 19760 -16870
rect 19800 -18880 19860 -16770
rect 19600 -20380 19660 -18920
rect 19700 -20290 19760 -19010
rect 19900 -19020 19960 -16670
rect 20000 -19080 20060 -16570
rect 19100 -21510 19160 -20580
rect 19200 -21510 19260 -20650
rect 19300 -21510 19360 -20660
rect 19400 -21510 19460 -20700
rect 19500 -21510 19560 -20660
rect 19600 -21510 19660 -20630
rect 19700 -21510 19760 -20520
rect 19800 -21510 19860 -19160
rect 20100 -19180 20160 -16490
rect 20200 -19220 20260 -16440
rect 19900 -21480 19960 -19220
rect 20300 -19300 20360 -16370
rect 20000 -21470 20060 -19320
rect 20400 -19340 20460 -16340
rect 20100 -21470 20160 -19380
rect 20500 -19400 20560 -16290
rect 20600 -19420 20660 -16270
rect 20200 -21470 20260 -19450
rect 20700 -19460 20760 -16230
rect 20800 -19480 20860 -16220
rect 20300 -21460 20360 -19500
rect 20900 -19510 20960 -16220
rect 21000 -19510 21060 -16220
rect 21100 -19510 21160 -16220
rect 21200 -19510 21260 -16220
rect 21300 -19510 21360 -16220
rect 21400 -19510 21460 -16220
rect 22000 -16230 22060 -15220
rect 21500 -19510 21560 -16250
rect 21600 -19460 21660 -16270
rect 22100 -16290 22160 -15220
rect 21700 -16460 21760 -16310
rect 22200 -16350 22260 -15220
rect 21800 -16650 21860 -16350
rect 21700 -19450 21760 -16880
rect 21900 -17150 21960 -16380
rect 22300 -16420 22360 -15220
rect 21800 -19420 21860 -17320
rect 22000 -17460 22060 -16440
rect 21900 -19370 21960 -17690
rect 22100 -17740 22160 -16500
rect 22400 -16510 22460 -15220
rect 22000 -19320 22060 -17910
rect 22200 -17920 22260 -16580
rect 22500 -16610 22560 -15220
rect 22300 -18060 22360 -16650
rect 22600 -16710 22660 -15220
rect 22100 -19270 22160 -18060
rect 22400 -18110 22460 -16750
rect 22700 -16850 22760 -15200
rect 22200 -19220 22260 -18200
rect 22300 -19130 22360 -18280
rect 22400 -19070 22460 -18310
rect 22500 -18970 22560 -16860
rect 22600 -18820 22660 -16990
rect 22800 -17000 22860 -15220
rect 22700 -18640 22760 -17180
rect 22900 -17230 22960 -15220
rect 22800 -18450 22860 -17360
rect 23000 -17500 23060 -15220
rect 22900 -18050 22960 -17770
rect 23100 -17880 23160 -15230
rect 24400 -15240 24460 -14570
rect 23200 -17840 23260 -15290
rect 23300 -17690 23360 -15510
rect 23500 -15610 23560 -15330
rect 24500 -15340 24560 -14570
rect 23400 -17500 23460 -15790
rect 23600 -15970 23660 -15350
rect 23500 -17190 23560 -16280
rect 20400 -21420 20460 -19550
rect 20500 -21400 20560 -19580
rect 20600 -21340 20660 -19620
rect 20700 -21290 20760 -19660
rect 20800 -21230 20860 -19670
rect 20900 -21180 20960 -19700
rect 21000 -21110 21060 -19700
rect 21100 -21030 21160 -19700
rect 21200 -20960 21260 -19700
rect 21300 -20900 21360 -19700
rect 21400 -20810 21460 -19700
rect 21500 -20750 21560 -19700
rect 21600 -20700 21660 -19660
rect 21700 -20600 21760 -19660
rect 21800 -20540 21860 -19620
rect 21900 -20480 21960 -19580
rect 22000 -20380 22060 -19530
rect 22100 -20330 22160 -19480
rect 22200 -20240 22260 -19420
rect 22300 -20170 22360 -19370
rect 22400 -20100 22460 -19280
rect 22500 -20010 22560 -19210
rect 22600 -19950 22660 -19060
rect 22700 -19860 22760 -18960
rect 22800 -19800 22860 -18780
rect 22900 -19700 22960 -18590
rect 23000 -19630 23060 -18320
rect 23100 -19540 23160 -18110
rect 23200 -19440 23260 -18070
rect 23300 -19390 23360 -17970
rect 23400 -19290 23460 -17880
rect 23500 -19190 23560 -17650
rect 23600 -19040 23660 -17340
rect 23700 -18940 23760 -15390
rect 24600 -15400 24660 -14570
rect 23800 -18800 23860 -15410
rect 23900 -18680 23960 -15460
rect 24700 -15500 24760 -14570
rect 24500 -15740 24560 -15650
rect 24000 -18600 24060 -17200
rect 24100 -17420 24160 -17050
rect 24200 -17400 24260 -16770
rect 24200 -18180 24260 -17600
rect 24300 -19320 24360 -16540
rect 23300 -19650 23360 -19590
rect 21100 -21460 21160 -21300
rect 21200 -21450 21260 -21230
rect 17700 -22160 17760 -21530
rect 17800 -22120 17860 -21530
rect 21400 -21550 21460 -21390
rect 21500 -21550 21560 -21070
rect 21600 -21300 21660 -20970
rect 21700 -21110 21760 -20830
rect 21800 -20890 21860 -20800
rect 21800 -21550 21860 -21250
rect 21900 -21550 21960 -21020
rect 22000 -21500 22060 -20790
rect 22100 -21240 22160 -20610
rect 22200 -20970 22260 -20460
rect 22300 -20690 22360 -20370
rect 22400 -20500 22460 -20330
rect 22200 -21450 22260 -21380
rect 22300 -21470 22360 -21100
rect 22400 -21430 22460 -20870
rect 22500 -21400 22560 -20640
rect 22600 -21100 22660 -20410
rect 22700 -20810 22760 -20180
rect 22800 -20590 22860 -20010
rect 22900 -20360 22960 -19940
rect 23000 -20070 23060 -19840
rect 23100 -19870 23160 -19810
rect 23300 -19950 23360 -19890
rect 22800 -21060 22860 -21000
rect 22600 -21220 22660 -21160
rect 22800 -21330 22860 -21120
rect 22900 -21290 22960 -20720
rect 23000 -21040 23060 -20530
rect 23100 -20810 23160 -20310
rect 23200 -20490 23260 -19990
rect 23300 -20200 23360 -20010
rect 24400 -20360 24460 -16310
rect 24500 -20440 24560 -15940
rect 24600 -20260 24660 -15610
rect 24700 -20150 24760 -15610
rect 24800 -20020 24860 -14560
rect 24900 -19920 24960 -14530
rect 25000 -19820 25060 -14500
rect 25100 -19720 25160 -14480
rect 25200 -19580 25260 -14350
rect 25300 -19390 25360 -14350
rect 25400 -19290 25460 -14350
rect 25500 -19340 25560 -6440
rect 25700 -6530 25760 0
rect 25800 -6680 25860 0
rect 25600 -19500 25660 -6710
rect 25900 -6770 25960 0
rect 26000 -6870 26060 0
rect 26100 -6930 26160 0
rect 26200 -7030 26260 0
rect 24500 -20700 24560 -20510
rect 23200 -21160 23260 -20940
rect 23300 -21140 23360 -20790
rect 24600 -20800 24660 -20430
rect 23400 -21030 23460 -20880
rect 24700 -20900 24760 -20440
rect 24800 -20980 24860 -20280
rect 24900 -21030 24960 -20160
rect 25000 -21110 25060 -20060
rect 17900 -22110 17960 -21570
rect 18000 -22070 18060 -21570
rect 18100 -22040 18160 -21600
rect 18200 -22030 18260 -21620
rect 18300 -21990 18360 -21660
rect 18400 -21990 18460 -21660
rect 18500 -21950 18560 -21660
rect 18600 -21950 18660 -21700
rect 18700 -21900 18760 -21710
rect 18800 -21900 18860 -21710
rect 18900 -21860 18960 -21710
rect 19000 -21850 19060 -21700
rect 19100 -21810 19160 -21710
rect 19200 -21810 19260 -21710
rect 19300 -21770 19360 -21710
rect 19400 -21780 19460 -21710
rect 19500 -21820 19560 -21710
rect 19600 -21970 19660 -21710
rect 19700 -21950 19760 -21710
rect 19800 -21920 19860 -21700
rect 19900 -21890 19960 -21660
rect 20000 -21850 20060 -21660
rect 20100 -21810 20160 -21710
rect 20200 -21770 20260 -21710
rect 20300 -21770 20360 -21710
rect 16500 -24590 16560 -24200
rect 16600 -24590 16660 -23700
rect 16700 -24570 16760 -23350
rect 16800 -23490 16860 -23110
rect 16900 -23420 16960 -22880
rect 17000 -23200 17060 -22700
rect 17100 -23140 17160 -22600
rect 17200 -23070 17260 -22550
rect 17300 -23020 17360 -22500
rect 17400 -22970 17460 -22450
rect 17500 -22910 17560 -22420
rect 17600 -22860 17660 -22370
rect 17700 -22810 17760 -22350
rect 17800 -22770 17860 -22320
rect 17900 -22730 17960 -22280
rect 18000 -22690 18060 -22270
rect 18100 -22660 18160 -22230
rect 18200 -22610 18260 -22230
rect 18300 -22590 18360 -22190
rect 18400 -22530 18460 -22170
rect 18500 -22480 18560 -22140
rect 18600 -22430 18660 -22140
rect 18700 -22410 18760 -22100
rect 18800 -22360 18860 -22080
rect 18900 -22330 18960 -22060
rect 19000 -22280 19060 -22020
rect 19100 -22220 19160 -22010
rect 19200 -22170 19260 -21980
rect 19300 -22120 19360 -21970
rect 19400 -22080 19460 -21980
rect 17200 -23340 17260 -23280
rect 17300 -23330 17360 -23220
rect 17400 -23290 17460 -23170
rect 17500 -23260 17560 -23120
rect 17600 -23240 17660 -23070
rect 17700 -23200 17760 -23020
rect 17800 -23160 17860 -22970
rect 17900 -23130 17960 -22930
rect 18000 -23120 18060 -22890
rect 18100 -23080 18160 -22870
rect 18200 -23080 18260 -22810
rect 18300 -23080 18360 -22760
rect 18400 -23060 18460 -22730
rect 18500 -23030 18560 -22690
rect 18600 -23040 18660 -22630
rect 18700 -23030 18760 -22610
rect 18800 -22990 18860 -22560
rect 18900 -22980 18960 -22530
rect 19000 -22950 19060 -22480
rect 19100 -22950 19160 -22430
rect 19200 -22910 19260 -22380
rect 19300 -22900 19360 -22330
rect 19400 -22900 19460 -22280
rect 19500 -22900 19560 -22230
rect 19600 -22860 19660 -22200
rect 19700 -22860 19760 -22150
rect 19800 -22820 19860 -22120
rect 19900 -22820 19960 -22070
rect 20000 -22820 20060 -22050
rect 20100 -22810 20160 -22010
rect 20200 -22750 20260 -21970
rect 20300 -22560 20360 -21940
rect 20400 -22380 20460 -21910
rect 20500 -22130 20560 -21880
rect 20600 -21990 20660 -21840
rect 20700 -21910 20760 -21830
rect 20800 -21880 20860 -21810
rect 21100 -22020 21160 -21710
rect 20500 -22560 20560 -22500
rect 20600 -22550 20660 -22320
rect 20700 -22500 20760 -22180
rect 20800 -22280 20860 -22100
rect 21100 -22290 21160 -22080
rect 21200 -22250 21260 -21700
rect 21300 -22200 21360 -21710
rect 21400 -22160 21460 -21750
rect 21500 -22120 21560 -21750
rect 21600 -22040 21660 -21750
rect 21700 -21990 21760 -21750
rect 21800 -21940 21860 -21750
rect 21900 -21900 21960 -21730
rect 22000 -21850 22060 -21710
rect 22100 -21800 22160 -21700
rect 22200 -21750 22260 -21660
rect 22300 -21730 22360 -21670
rect 20400 -22940 20460 -22880
rect 20400 -23060 20460 -23000
rect 16800 -24590 16860 -23710
rect 16900 -24560 16960 -23620
rect 17000 -24550 17060 -23580
rect 17100 -24490 17160 -23560
rect 17200 -24390 17260 -23530
rect 17300 -24290 17360 -23520
rect 17400 -24190 17460 -23490
rect 17500 -23610 17560 -23450
rect 17600 -23510 17660 -23410
rect 17700 -23510 17760 -23390
rect 17800 -23470 17860 -23360
rect 17900 -23550 17960 -23320
rect 15600 -26280 15660 -26180
rect 15700 -26240 15760 -26040
rect 15800 -26160 15860 -25950
rect 15900 -26110 15960 -25840
rect 16000 -26040 16060 -25750
rect 16100 -25990 16160 -25600
rect 16200 -25940 16260 -25500
rect 16300 -25860 16360 -25440
rect 16400 -25810 16460 -25340
rect 16500 -25770 16560 -25240
rect 16600 -25720 16660 -25150
rect 16700 -25640 16760 -25080
rect 16800 -25600 16860 -24990
rect 16900 -25520 16960 -24890
rect 17000 -25460 17060 -24830
rect 17100 -25400 17160 -24730
rect 17200 -25330 17260 -24630
rect 17300 -25260 17360 -24570
rect 17400 -25190 17460 -24470
rect 17500 -25130 17560 -24370
rect 17600 -25040 17660 -24230
rect 17700 -24980 17760 -24000
rect 17800 -24920 17860 -23810
rect 17900 -24850 17960 -23610
rect 18000 -24780 18060 -23310
rect 18100 -24710 18160 -23270
rect 18200 -24650 18260 -23270
rect 18300 -23940 18360 -23270
rect 18400 -23800 18460 -23230
rect 18500 -23700 18560 -23230
rect 18600 -23600 18660 -23230
rect 18700 -23540 18760 -23230
rect 18800 -23440 18860 -23190
rect 18900 -23390 18960 -23150
rect 19000 -23300 19060 -23140
rect 19100 -23230 19160 -23140
rect 19200 -23170 19260 -23110
rect 20400 -23230 20460 -23150
rect 18400 -24400 18460 -24120
rect 18500 -24630 18560 -23940
rect 13800 -30950 13860 -30630
rect 13900 -31170 13960 -29010
rect 14000 -31120 14060 -28550
rect 14100 -31010 14160 -28250
rect 14200 -30950 14260 -27970
rect 14300 -30860 14360 -27710
rect 14400 -30800 14460 -27560
rect 14500 -30730 14560 -27410
rect 14600 -30650 14660 -27310
rect 14700 -30580 14760 -27260
rect 14800 -30530 14860 -27160
rect 14900 -30470 14960 -27100
rect 15000 -30350 15060 -26960
rect 15100 -30300 15160 -26860
rect 15200 -30260 15260 -26790
rect 15300 -30170 15360 -26700
rect 15400 -30100 15460 -26630
rect 15500 -30050 15560 -26550
rect 15600 -29980 15660 -26490
rect 15700 -29910 15760 -26440
rect 15800 -29860 15860 -26380
rect 15900 -29810 15960 -26310
rect 16000 -29760 16060 -26270
rect 16100 -29730 16160 -26190
rect 16200 -29690 16260 -26140
rect 16300 -29650 16360 -26090
rect 16400 -29620 16460 -26020
rect 16500 -29570 16560 -25970
rect 16600 -29550 16660 -25920
rect 16700 -29500 16760 -25870
rect 16800 -29440 16860 -25800
rect 16900 -29380 16960 -25750
rect 17000 -29330 17060 -25670
rect 17100 -29270 17160 -25600
rect 17200 -29220 17260 -25550
rect 17300 -29160 17360 -25490
rect 17400 -29070 17460 -25410
rect 17500 -26610 17560 -25340
rect 17600 -26470 17660 -25280
rect 17700 -26370 17760 -25190
rect 17800 -26270 17860 -25130
rect 17900 -26170 17960 -25070
rect 18000 -26130 18060 -25010
rect 18100 -26190 18160 -24930
rect 18200 -25960 18260 -24860
rect 18300 -25730 18360 -24790
rect 18400 -25460 18460 -24770
rect 18600 -24820 18660 -23840
rect 18700 -24960 18760 -23760
rect 18500 -25100 18560 -24960
rect 18800 -25100 18860 -23680
rect 17700 -26840 17760 -26610
rect 17800 -26750 17860 -26500
rect 17900 -26570 17960 -26410
rect 18000 -26430 18060 -26370
rect 17500 -28960 17560 -26950
rect 17600 -28860 17660 -27060
rect 17700 -28770 17760 -27050
rect 17800 -28660 17860 -26990
rect 17900 -28520 17960 -26890
rect 18000 -28380 18060 -26750
rect 18100 -28200 18160 -26560
rect 18200 -28000 18260 -26370
rect 18300 -27820 18360 -26140
rect 18400 -27590 18460 -25870
rect 18500 -27390 18560 -25640
rect 18600 -27080 18660 -25370
rect 18700 -26680 18760 -25250
rect 18900 -25290 18960 -23590
rect 19000 -25320 19060 -23530
rect 19100 -25290 19160 -23450
rect 19200 -25260 19260 -23380
rect 19300 -25210 19360 -23320
rect 19400 -25160 19460 -23260
rect 19500 -25120 19560 -23230
rect 19600 -25090 19660 -23260
rect 19700 -25040 19760 -23270
rect 19800 -25010 19860 -23280
rect 19900 -24960 19960 -23320
rect 20000 -24900 20060 -23330
rect 20100 -24760 20160 -23460
rect 20200 -24490 20260 -23560
rect 18800 -26410 18860 -25430
rect 18900 -25780 18960 -25540
rect 19400 -25560 19460 -25500
rect 17100 -29630 17160 -29480
rect 13700 -32430 13760 -31530
rect 13800 -32390 13860 -31510
rect 13900 -32350 13960 -31410
rect 14000 -32330 14060 -31330
rect 14100 -32270 14160 -31250
rect 14200 -32220 14260 -31150
rect 14300 -32200 14360 -31100
rect 14400 -32140 14460 -31000
rect 14500 -32120 14560 -30940
rect 14600 -32080 14660 -30880
rect 14700 -32040 14760 -30810
rect 14800 -32010 14860 -30730
rect 14900 -31990 14960 -30690
rect 15000 -31940 15060 -30770
rect 15200 -30990 15260 -30460
rect 15100 -31860 15160 -31220
rect 15300 -31400 15360 -30400
rect 15200 -31860 15260 -31710
rect 15400 -31940 15460 -30330
rect 15200 -32010 15260 -31950
rect 1400 -38700 1460 -38620
rect 1500 -38670 1560 -38570
rect 1600 -38620 1660 -38470
rect 1700 -38600 1760 -38410
rect 1800 -38550 1860 -38340
rect 1900 -38490 1960 -38260
rect 2000 -38450 2060 -38200
rect 2100 -38420 2160 -38120
rect 2200 -38390 2260 -38050
rect 2300 -38350 2360 -37990
rect 2400 -38350 2460 -37900
rect 2500 -38310 2560 -37830
rect 2600 -38310 2660 -37770
rect 2700 -38310 2760 -37690
rect 2800 -38310 2860 -37620
rect 2900 -38260 2960 -37560
rect 3000 -38270 3060 -37470
rect 3100 -38270 3160 -37410
rect 3200 -38270 3260 -37330
rect 3300 -38270 3360 -37260
rect 3400 -38270 3460 -37190
rect 3500 -38270 3560 -37120
rect 3600 -38260 3660 -37040
rect 3700 -38230 3760 -36980
rect 3800 -38220 3860 -36900
rect 3900 -38220 3960 -36830
rect 4000 -38220 4060 -36760
rect 4100 -38220 4160 -36670
rect 4200 -38220 4260 -36620
rect 4300 -38220 4360 -36520
rect 4400 -38180 4460 -36460
rect 4500 -38180 4560 -36380
rect 4600 -38180 4660 -36300
rect 4700 -38170 4760 -36240
rect 4800 -38130 4860 -36160
rect 4900 -38140 4960 -36090
rect 5000 -38130 5060 -36030
rect 5100 -38090 5160 -35970
rect 5200 -38090 5260 -35870
rect 5300 -38060 5360 -35820
rect 5400 -38050 5460 -35760
rect 5500 -38050 5560 -35710
rect 5600 -38030 5660 -35630
rect 5700 -38000 5760 -35580
rect 5800 -38000 5860 -35510
rect 5900 -38010 5960 -35460
rect 6000 -38000 6060 -35390
rect 6100 -37960 6160 -35340
rect 6200 -37960 6260 -35290
rect 6300 -37960 6360 -35220
rect 6400 -37920 6460 -35160
rect 6500 -37910 6560 -35120
rect 6600 -37870 6660 -35050
rect 6700 -37870 6760 -34990
rect 6800 -37830 6860 -34950
rect 6900 -37800 6960 -34900
rect 7000 -37790 7060 -34850
rect 7100 -37750 7160 -34800
rect 7200 -37720 7260 -34750
rect 7300 -37700 7360 -34720
rect 7400 -37660 7460 -34670
rect 7500 -37640 7560 -34620
rect 7600 -37610 7660 -34560
rect 7700 -37580 7760 -34540
rect 7800 -37570 7860 -34490
rect 7900 -37530 7960 -34460
rect 8000 -37490 8060 -34410
rect 8100 -37470 8160 -34370
rect 8200 -37420 8260 -34330
rect 8300 -37390 8360 -34290
rect 8400 -37350 8460 -34260
rect 8500 -37310 8560 -34200
rect 8600 -37270 8660 -34180
rect 8700 -37230 8760 -34150
rect 8800 -37180 8860 -34120
rect 8900 -37150 8960 -34100
rect 9000 -37130 9060 -34060
rect 9100 -37080 9160 -34030
rect 9200 -37040 9260 -33980
rect 9300 -37000 9360 -33960
rect 9400 -36960 9460 -33940
rect 9500 -36920 9560 -33900
rect 9600 -36870 9660 -33880
rect 9700 -36820 9760 -33820
rect 9800 -36770 9860 -33800
rect 9900 -36740 9960 -33760
rect 10000 -36690 10060 -33720
rect 10100 -36650 10160 -33690
rect 10200 -36600 10260 -33640
rect 10300 -36540 10360 -33610
rect 10400 -36490 10460 -33580
rect 10500 -36420 10560 -33550
rect 10600 -36370 10660 -33510
rect 10700 -36300 10760 -33480
rect 10800 -36250 10860 -33450
rect 10900 -36180 10960 -33410
rect 11000 -36110 11060 -33400
rect 11100 -36050 11160 -33370
rect 11200 -35990 11260 -33330
rect 11300 -35910 11360 -33290
rect 11400 -35840 11460 -33280
rect 11500 -35770 11560 -33240
rect 11600 -35700 11660 -33200
rect 11700 -35630 11760 -33190
rect 11800 -35570 11860 -33160
rect 11900 -35390 11960 -33120
rect 12000 -35250 12060 -33110
rect 12100 -35050 12160 -33070
rect 12200 -34910 12260 -33030
rect 12300 -34770 12360 -33020
rect 12400 -34630 12460 -32980
rect 12500 -34530 12560 -32950
rect 12600 -34430 12660 -32930
rect 12700 -34280 12760 -32890
rect 12800 -34180 12860 -32850
rect 12900 -34080 12960 -32840
rect 13000 -33980 13060 -32800
rect 13100 -33880 13160 -32780
rect 13200 -33780 13260 -32760
rect 13300 -33680 13360 -32720
rect 13400 -33580 13460 -32720
rect 13500 -33480 13560 -32680
rect 13600 -33380 13660 -32660
rect 13700 -33240 13760 -32630
rect 13800 -33140 13860 -32590
rect 13900 -33040 13960 -32550
rect 14000 -32940 14060 -32530
rect 14100 -32840 14160 -32470
rect 14200 -32740 14260 -32430
rect 14300 -32640 14360 -32380
rect 14400 -32540 14460 -32350
rect 14500 -32440 14560 -32320
rect 14600 -32350 14660 -32290
rect 11500 -36050 11560 -35990
rect 10900 -37990 10960 -37930
rect 900 -48580 960 -39020
rect 1000 -48580 1060 -39020
rect 1100 -48580 1160 -38980
rect 1200 -48580 1260 -38980
rect 1300 -48580 1360 -38980
rect 1400 -48580 1460 -39030
rect 1500 -48580 1560 -39060
rect 1600 -48580 1660 -39080
rect 1700 -48580 1760 -39120
rect 1800 -48580 1860 -39160
rect 1900 -48580 1960 -39160
rect 2000 -48580 2060 -39200
rect 2100 -48580 2160 -39200
rect 2200 -48580 2260 -39230
rect 2300 -48580 2360 -39250
rect 2400 -48580 2460 -39280
rect 2500 -48580 2560 -39310
rect 2600 -48580 2660 -39330
rect 2700 -48580 2760 -39340
rect 2800 -48580 2860 -39380
rect 2900 -48580 2960 -39380
rect 3000 -48580 3060 -39420
rect 3100 -48580 3160 -39460
rect 3200 -48580 3260 -39490
rect 3300 -48580 3360 -39510
rect 3400 -48580 3460 -39520
rect 3500 -48580 3560 -39550
rect 3600 -48580 3660 -39550
rect 3700 -48580 3760 -39550
rect 3800 -48580 3860 -39570
rect 3900 -48580 3960 -39590
rect 4000 -44410 4060 -39590
rect 4100 -43700 4160 -39590
rect 4200 -43120 4260 -39590
rect 4300 -42540 4360 -39590
rect 4400 -42270 4460 -39590
rect 4500 -42000 4560 -39550
rect 4600 -41710 4660 -39550
rect 4700 -41400 4760 -39550
rect 4800 -41170 4860 -39550
rect 4900 -40900 4960 -39510
rect 5000 -40580 5060 -39510
rect 5100 -40350 5160 -39500
rect 5200 -40080 5260 -39460
rect 5300 -39810 5360 -39420
rect 5400 -39610 5460 -39380
rect 5500 -39450 5560 -39390
rect 7100 -44090 7160 -44030
rect 7200 -44060 7260 -43950
rect 7300 -44050 7360 -43870
rect 7400 -44010 7460 -43810
rect 7500 -43990 7560 -43710
rect 7600 -43970 7660 -43620
rect 7700 -43960 7760 -43520
rect 7800 -43920 7860 -43420
rect 7900 -43900 7960 -43320
rect 8000 -43870 8060 -43220
rect 8100 -43840 8160 -43120
rect 8200 -43820 8260 -42980
rect 8300 -43790 8360 -42830
rect 8400 -43760 8460 -42690
rect 8500 -43750 8560 -42500
rect 8600 -43710 8660 -42270
rect 8700 -43670 8760 -42080
rect 8800 -43620 8860 -41900
rect 8900 -43530 8960 -41670
rect 9000 -43530 9060 -41480
rect 7700 -44190 7760 -44130
rect 4000 -48580 4060 -45380
rect 4100 -48580 4160 -45360
rect 4200 -48580 4260 -45350
rect 4300 -48580 4360 -45300
rect 4400 -48580 4460 -45330
rect 4500 -48580 4560 -45340
rect 4600 -48580 4660 -45340
rect 4700 -48580 4760 -45340
rect 4800 -48580 4860 -45300
rect 4900 -48580 4960 -45290
rect 5000 -48580 5060 -45290
rect 5100 -48580 5160 -45300
rect 5200 -48580 5260 -45250
rect 5300 -48580 5360 -45250
rect 5400 -48580 5460 -45220
rect 5500 -48580 5560 -45210
rect 5600 -48580 5660 -45210
rect 5700 -48580 5760 -45160
rect 5800 -48580 5860 -45160
rect 5900 -48580 5960 -45160
rect 6000 -48580 6060 -45160
rect 6100 -48580 6160 -45160
rect 6200 -48580 6260 -45120
rect 6300 -48580 6360 -45080
rect 6400 -48580 6460 -45070
rect 6500 -48580 6560 -45040
rect 6600 -48580 6660 -44990
rect 6700 -48580 6760 -44950
rect 6800 -48580 6860 -44910
rect 6900 -48580 6960 -44860
rect 7000 -48580 7060 -44830
rect 7100 -48580 7160 -44780
rect 7200 -48580 7260 -44730
rect 7300 -48580 7360 -44660
rect 7400 -48580 7460 -44600
rect 7500 -48580 7560 -44540
rect 7600 -48580 7660 -44470
rect 7700 -48580 7760 -44400
rect 7800 -48580 7860 -44350
rect 7900 -48580 7960 -44300
rect 8000 -45550 8060 -44090
rect 8100 -45190 8160 -44040
rect 8200 -44910 8260 -44000
rect 8300 -44680 8360 -43990
rect 8400 -44360 8460 -43950
rect 8500 -44180 8560 -43940
rect 8600 -43990 8660 -43910
rect 8200 -45470 8260 -45370
rect 8000 -45760 8060 -45610
rect 8000 -48580 8060 -45890
rect 8100 -48580 8160 -45900
rect 8200 -48580 8260 -45530
rect 8300 -48580 8360 -45090
rect 8400 -48580 8460 -44820
rect 8500 -48580 8560 -44590
rect 8600 -48580 8660 -44320
rect 8700 -48580 8760 -44130
rect 8800 -48580 8860 -43990
rect 8900 -48580 8960 -43840
rect 9000 -48580 9060 -43700
rect 9100 -48580 9160 -41290
rect 9200 -48580 9260 -41100
rect 9300 -48580 9360 -40910
rect 9400 -48580 9460 -40730
rect 9500 -48580 9560 -40550
rect 9600 -48580 9660 -40360
rect 9700 -48580 9760 -40170
rect 9800 -48580 9860 -40030
rect 9900 -48580 9960 -39840
rect 10000 -48580 10060 -39690
rect 10100 -48580 10160 -39510
rect 10200 -48580 10260 -39360
rect 10300 -39860 10360 -39230
rect 10400 -39290 10460 -39230
rect 10400 -42310 10460 -40380
rect 10300 -48580 10360 -42700
rect 10500 -43060 10560 -39550
rect 10400 -43390 10460 -43330
rect 10400 -48580 10460 -43580
rect 10600 -43900 10660 -38920
rect 10500 -48580 10560 -44170
rect 10700 -44390 10760 -38560
rect 10600 -48580 10660 -44610
rect 10800 -44840 10860 -38290
rect 10700 -48580 10760 -45060
rect 10900 -45330 10960 -38050
rect 10900 -45530 10960 -45390
rect 10800 -48580 10860 -45820
rect 10900 -48580 10960 -45900
rect 11000 -48580 11060 -37650
rect 11100 -48580 11160 -37420
rect 11200 -48580 11260 -37190
rect 11300 -48580 11360 -36920
rect 11400 -48580 11460 -36710
rect 11500 -48580 11560 -36510
rect 11600 -48580 11660 -36270
rect 11700 -48580 11760 -36080
rect 11800 -48580 11860 -35940
rect 11900 -48580 11960 -35750
rect 12000 -48580 12060 -35520
rect 12100 -48580 12160 -35380
rect 12200 -48580 12260 -35190
rect 12300 -48580 12360 -35050
rect 12400 -48580 12460 -34910
rect 12500 -48580 12560 -34810
rect 12600 -48580 12660 -34660
rect 12700 -48580 12760 -34570
rect 12800 -48580 12860 -34420
rect 12900 -48580 12960 -34320
rect 13000 -48580 13060 -34220
rect 13100 -48580 13160 -34120
rect 13200 -48580 13260 -34020
rect 13300 -48580 13360 -33920
rect 13400 -48580 13460 -33820
rect 13500 -48580 13560 -33720
rect 13600 -48580 13660 -33630
rect 13700 -48580 13760 -33470
rect 13800 -48580 13860 -33380
rect 13900 -48580 13960 -33280
rect 14000 -48580 14060 -33180
rect 14100 -48580 14160 -33080
rect 14200 -48580 14260 -32980
rect 14300 -48580 14360 -32880
rect 14400 -48580 14460 -32780
rect 14500 -48580 14560 -32680
rect 14600 -48580 14660 -32580
rect 14700 -48580 14760 -32480
rect 14800 -48580 14860 -32380
rect 14900 -48580 14960 -32280
rect 15000 -48580 15060 -32200
rect 15100 -48580 15160 -32200
rect 15200 -48580 15260 -32160
rect 15300 -48580 15360 -32160
rect 15500 -32300 15560 -30250
rect 15400 -48580 15460 -32430
rect 15600 -32570 15660 -30190
rect 15500 -48580 15560 -32750
rect 15700 -32900 15760 -30130
rect 15800 -31850 15860 -30060
rect 15900 -32000 15960 -30010
rect 15800 -32210 15860 -32140
rect 15600 -48580 15660 -33020
rect 15800 -33030 15860 -32270
rect 16000 -32360 16060 -29960
rect 16000 -32480 16060 -32420
rect 16000 -32650 16060 -32540
rect 16000 -32830 16060 -32770
rect 16000 -32950 16060 -32890
rect 16000 -33110 16060 -33050
rect 16000 -33230 16060 -33170
rect 15700 -48580 15760 -33260
rect 15800 -48580 15860 -33400
rect 15900 -48580 15960 -33450
rect 16000 -48580 16060 -33290
rect 16100 -48580 16160 -29930
rect 16200 -48580 16260 -29890
rect 16300 -48580 16360 -29850
rect 16400 -48580 16460 -29810
rect 16500 -48580 16560 -29770
rect 16600 -48580 16660 -29750
rect 16700 -48580 16760 -29700
rect 16800 -48580 16860 -29650
rect 16900 -48580 16960 -29630
rect 17000 -48580 17060 -29810
rect 17200 -29950 17260 -29420
rect 17100 -48580 17160 -30130
rect 17300 -30260 17360 -29360
rect 17200 -30530 17260 -30470
rect 17200 -48580 17260 -30590
rect 17400 -30660 17460 -29280
rect 17300 -48580 17360 -30850
rect 17500 -30990 17560 -29210
rect 17400 -48580 17460 -31160
rect 17600 -31260 17660 -29110
rect 17500 -31510 17560 -31450
rect 17500 -48580 17560 -31570
rect 17700 -31580 17760 -29010
rect 17700 -31700 17760 -31640
rect 17600 -48580 17660 -31840
rect 17800 -31940 17860 -28910
rect 17700 -48580 17760 -32120
rect 17900 -32210 17960 -28800
rect 17800 -48580 17860 -32350
rect 18000 -32440 18060 -28660
rect 17900 -48580 17960 -32670
rect 18100 -32760 18160 -28520
rect 18000 -48580 18060 -32900
rect 18200 -32990 18260 -28330
rect 18100 -48580 18160 -33120
rect 18300 -33180 18360 -28190
rect 18200 -48580 18260 -33360
rect 18400 -33450 18460 -27950
rect 18300 -48580 18360 -33590
rect 18500 -33680 18560 -27770
rect 18400 -48580 18460 -33820
rect 18600 -33870 18660 -27540
rect 18500 -48580 18560 -34000
rect 18700 -34060 18760 -27300
rect 18800 -34240 18860 -26900
rect 18600 -45320 18660 -34240
rect 18700 -45220 18760 -34380
rect 18900 -34430 18960 -26750
rect 19000 -34520 19060 -26620
rect 18800 -45120 18860 -34520
rect 19100 -34670 19160 -26260
rect 18900 -45050 18960 -34710
rect 19200 -34770 19260 -26020
rect 19000 -44960 19060 -34810
rect 19300 -34820 19360 -25750
rect 19400 -34860 19460 -25620
rect 19100 -44910 19160 -34890
rect 19200 -44810 19260 -34970
rect 19300 -44750 19360 -35020
rect 19400 -44650 19460 -35020
rect 19500 -44550 19560 -25340
rect 19600 -44450 19660 -25290
rect 19700 -44350 19760 -25240
rect 19800 -44210 19860 -25220
rect 19900 -44070 19960 -25160
rect 20000 -37520 20060 -25110
rect 20100 -37380 20160 -25040
rect 20200 -33100 20260 -24900
rect 20300 -29390 20360 -26010
rect 20500 -26450 20560 -22800
rect 20600 -26440 20660 -22750
rect 20700 -26370 20760 -22700
rect 20800 -26300 20860 -22660
rect 20900 -26220 20960 -22620
rect 21000 -26160 21060 -22570
rect 21100 -26070 21160 -22520
rect 21200 -25970 21260 -22450
rect 21300 -25470 21360 -22410
rect 21400 -25160 21460 -22370
rect 21500 -24930 21560 -22320
rect 21600 -24740 21660 -22270
rect 21700 -23380 21760 -22220
rect 21800 -22890 21860 -22170
rect 21900 -22520 21960 -22100
rect 22000 -22250 22060 -22050
rect 22100 -22110 22160 -22000
rect 22200 -22050 22260 -21990
rect 21800 -24470 21860 -24040
rect 21300 -25870 21360 -25790
rect 21500 -26000 21560 -25300
rect 20400 -28900 20460 -26730
rect 20500 -28540 20560 -26690
rect 20600 -28180 20660 -26640
rect 20700 -27950 20760 -26580
rect 20800 -27720 20860 -26520
rect 20900 -27530 20960 -26450
rect 21000 -27340 21060 -26360
rect 21100 -27200 21160 -26310
rect 21200 -27010 21260 -26190
rect 21300 -26660 21360 -26120
rect 20500 -29460 20560 -29130
rect 20600 -29400 20660 -28720
rect 20700 -29300 20760 -28400
rect 20800 -29200 20860 -28080
rect 20900 -29100 20960 -27850
rect 21000 -29040 21060 -27670
rect 21100 -28940 21160 -27480
rect 21200 -28880 21260 -27340
rect 21300 -28790 21360 -27150
rect 21400 -28720 21460 -26970
rect 21500 -28630 21560 -26600
rect 21600 -28560 21660 -25060
rect 21700 -28570 21760 -24880
rect 20300 -32610 20360 -29930
rect 20400 -32380 20460 -29870
rect 20500 -32060 20560 -29730
rect 20600 -31750 20660 -29630
rect 20700 -31520 20760 -29530
rect 20800 -31240 20860 -29430
rect 20900 -30920 20960 -29340
rect 21000 -30600 21060 -29240
rect 21100 -30290 21160 -29240
rect 21300 -29380 21360 -29060
rect 21100 -30850 21160 -30790
rect 20900 -31040 20960 -30980
rect 20400 -32860 20460 -32800
rect 20300 -34610 20360 -33460
rect 20200 -37190 20260 -34830
rect 20400 -35060 20460 -32920
rect 20400 -35210 20460 -35120
rect 20300 -36700 20360 -35460
rect 20500 -35590 20560 -32520
rect 20400 -36250 20460 -35770
rect 20400 -36980 20460 -36920
rect 20300 -37510 20360 -37330
rect 20400 -37430 20460 -37060
rect 20500 -37370 20560 -36520
rect 20600 -37270 20660 -32240
rect 20700 -37180 20760 -31980
rect 20800 -37110 20860 -31660
rect 20900 -37040 20960 -31420
rect 21000 -36960 21060 -31150
rect 21100 -36900 21160 -30910
rect 21200 -36850 21260 -30470
rect 20000 -43970 20060 -37850
rect 20100 -43820 20160 -37840
rect 20200 -43730 20260 -37790
rect 20300 -43570 20360 -37720
rect 20400 -43440 20460 -37670
rect 20500 -43290 20560 -37570
rect 20600 -43100 20660 -37510
rect 20700 -42960 20760 -37410
rect 20800 -42780 20860 -37310
rect 20900 -42590 20960 -37250
rect 21000 -42400 21060 -37200
rect 21100 -42220 21160 -37300
rect 21300 -37430 21360 -30110
rect 21400 -37580 21460 -28920
rect 21200 -42030 21260 -37580
rect 21500 -37720 21560 -28910
rect 21700 -28960 21760 -28760
rect 21600 -29200 21660 -29140
rect 21300 -41790 21360 -37720
rect 21600 -37860 21660 -29260
rect 21800 -29320 21860 -24690
rect 21400 -41610 21460 -37860
rect 21700 -37960 21760 -29500
rect 21900 -29550 21960 -23110
rect 21500 -41430 21560 -38000
rect 21600 -41190 21660 -38100
rect 21800 -38110 21860 -29730
rect 22000 -29820 22060 -22710
rect 21900 -38200 21960 -29960
rect 22100 -30060 22160 -22430
rect 21700 -41000 21760 -38250
rect 22000 -38310 22060 -30280
rect 22200 -30370 22260 -22250
rect 21800 -40820 21860 -38350
rect 22100 -38410 22160 -30550
rect 22300 -30650 22360 -22150
rect 21900 -40590 21960 -38440
rect 22200 -38510 22260 -30780
rect 22400 -30870 22460 -22050
rect 22000 -40310 22060 -38550
rect 22300 -38610 22360 -31040
rect 22500 -31100 22560 -22000
rect 22100 -40010 22160 -38650
rect 22400 -38710 22460 -31240
rect 22600 -31300 22660 -21940
rect 22700 -31370 22760 -21890
rect 22800 -31250 22860 -21850
rect 22900 -31110 22960 -21900
rect 23000 -30920 23060 -22450
rect 23100 -30770 23160 -22440
rect 23200 -30670 23260 -22120
rect 23300 -30600 23360 -21980
rect 23400 -30520 23460 -21830
rect 23500 -30470 23560 -21690
rect 23600 -30430 23660 -21590
rect 23700 -30350 23760 -21490
rect 23800 -30290 23860 -21410
rect 23900 -30210 23960 -21340
rect 24000 -30130 24060 -21290
rect 24100 -30040 24160 -21240
rect 24200 -29930 24260 -21190
rect 24300 -29830 24360 -21180
rect 24400 -29730 24460 -21140
rect 24500 -29640 24560 -21140
rect 24600 -29530 24660 -21140
rect 24700 -29480 24760 -21140
rect 25100 -21190 25160 -19960
rect 24800 -29380 24860 -21190
rect 25200 -21220 25260 -19820
rect 24900 -29300 24960 -21250
rect 25300 -21280 25360 -19720
rect 25000 -29220 25060 -21350
rect 25100 -29120 25160 -21450
rect 25200 -29020 25260 -21550
rect 25400 -21590 25460 -19590
rect 25500 -21680 25560 -19620
rect 25700 -19760 25760 -7040
rect 26300 -7100 26360 0
rect 26000 -7280 26060 -7220
rect 26400 -7230 26460 0
rect 25600 -21640 25660 -19940
rect 25800 -20040 25860 -7310
rect 26000 -7410 26060 -7340
rect 25700 -21640 25760 -20270
rect 25900 -20390 25960 -7540
rect 26100 -7670 26160 -7340
rect 26500 -7380 26560 0
rect 26000 -7880 26060 -7820
rect 26200 -7940 26260 -7400
rect 25800 -21680 25860 -20580
rect 26000 -20760 26060 -7940
rect 26200 -8060 26260 -8000
rect 26100 -21160 26160 -8170
rect 26300 -8320 26360 -7500
rect 26600 -7520 26660 0
rect 26200 -21110 26260 -8530
rect 26400 -8750 26460 -7600
rect 26700 -7620 26760 0
rect 26300 -21000 26360 -8980
rect 26500 -9200 26560 -7700
rect 26800 -7720 26860 0
rect 26500 -9380 26560 -9320
rect 26500 -9500 26560 -9440
rect 26400 -11670 26460 -9950
rect 26400 -20950 26460 -11920
rect 26500 -20850 26560 -11910
rect 26600 -12120 26660 -7800
rect 26900 -7820 26960 0
rect 26700 -12140 26760 -7900
rect 27000 -7920 27060 0
rect 26600 -20750 26660 -12290
rect 26800 -12330 26860 -8000
rect 27100 -8020 27160 0
rect 26900 -12600 26960 -8100
rect 27200 -8120 27260 0
rect 26700 -20650 26760 -12610
rect 26900 -12720 26960 -12660
rect 26800 -20550 26860 -12870
rect 27000 -12970 27060 -8200
rect 27300 -8220 27360 0
rect 26900 -20450 26960 -13130
rect 27100 -13190 27160 -8350
rect 27400 -8360 27460 0
rect 27000 -20310 27060 -13330
rect 27200 -13430 27260 -8440
rect 27500 -8460 27560 0
rect 27100 -20080 27160 -13650
rect 27200 -19840 27260 -13710
rect 27300 -19640 27360 -8540
rect 27600 -8640 27660 0
rect 27400 -13980 27460 -8690
rect 27700 -8790 27760 0
rect 27500 -13990 27560 -8830
rect 27800 -8940 27860 0
rect 27300 -20230 27360 -19980
rect 25900 -21700 25960 -21240
rect 26000 -21730 26060 -21360
rect 26100 -21730 26160 -21320
rect 26200 -21770 26260 -21310
rect 26300 -21810 26360 -21240
rect 25300 -28920 25360 -22130
rect 25400 -28780 25460 -22100
rect 25500 -28590 25560 -21920
rect 25600 -28450 25660 -21840
rect 25700 -28170 25760 -21840
rect 26400 -21860 26460 -21150
rect 25800 -27990 25860 -21880
rect 25900 -27960 25960 -21880
rect 26000 -23530 26060 -21920
rect 26100 -23460 26160 -21930
rect 26500 -21950 26560 -21090
rect 26200 -23410 26260 -21970
rect 26300 -23380 26360 -22010
rect 26400 -23370 26460 -22090
rect 26600 -22140 26660 -20990
rect 26700 -22210 26760 -20890
rect 26800 -22210 26860 -20790
rect 26900 -22220 26960 -20690
rect 26500 -23340 26560 -22240
rect 27000 -22280 27060 -20590
rect 27100 -22290 27160 -20660
rect 27400 -20770 27460 -14170
rect 27600 -14310 27660 -8970
rect 27900 -9000 27960 0
rect 28000 -8120 28060 0
rect 28100 -7720 28160 0
rect 28200 -7620 28260 0
rect 28300 -7560 28360 0
rect 28400 -7510 28460 0
rect 28500 -7480 28560 0
rect 28600 -7430 28660 0
rect 28700 -7400 28760 0
rect 28800 -7350 28860 0
rect 28900 -7310 28960 0
rect 29000 -7250 29060 0
rect 29100 -7230 29160 0
rect 29200 -7180 29260 0
rect 29300 -7120 29360 0
rect 29400 -7070 29460 0
rect 29500 -6800 29560 0
rect 29600 -6490 29660 0
rect 29700 -6260 29760 0
rect 29800 -5890 29860 0
rect 29900 -5590 29960 0
rect 30000 -5380 30060 0
rect 30100 -5160 30160 0
rect 30200 -4930 30260 0
rect 30300 -4650 30360 0
rect 30400 -4420 30460 0
rect 30500 -4190 30560 0
rect 30600 -4050 30660 0
rect 30700 -3860 30760 0
rect 30800 -3630 30860 0
rect 30900 -3490 30960 0
rect 31000 -3340 31060 0
rect 31100 -3160 31160 0
rect 31200 -3020 31260 0
rect 31300 -2870 31360 0
rect 31400 -2720 31460 0
rect 31500 -2580 31560 0
rect 31600 -2490 31660 0
rect 31700 -2340 31760 0
rect 31800 -2240 31860 0
rect 31900 -2140 31960 0
rect 32000 -2030 32060 0
rect 32100 -1940 32160 0
rect 32200 -1840 32260 0
rect 32300 -1740 32360 0
rect 32400 -1640 32460 0
rect 32500 -1580 32560 0
rect 32600 -1480 32660 0
rect 32700 -1390 32760 0
rect 32800 -1280 32860 0
rect 32900 -1270 32960 0
rect 33000 -1350 33060 0
rect 33100 -1400 33160 0
rect 33200 -1480 33260 0
rect 33300 -1540 33360 0
rect 33400 -1620 33460 0
rect 29900 -7390 29960 -7290
rect 28500 -8570 28560 -8510
rect 28600 -8530 28660 -8280
rect 28700 -8380 28760 -8140
rect 28800 -8240 28860 -7990
rect 28900 -8100 28960 -7850
rect 29000 -7960 29060 -7750
rect 29100 -7810 29160 -7650
rect 29200 -7720 29260 -7570
rect 28400 -8720 28460 -8660
rect 28500 -8690 28560 -8630
rect 29800 -8750 29860 -8390
rect 29900 -8710 29960 -7500
rect 30000 -8620 30060 -6880
rect 30100 -8160 30160 -6520
rect 30200 -7490 30260 -6210
rect 30300 -6960 30360 -5840
rect 30400 -6470 30460 -5570
rect 30500 -6060 30560 -5340
rect 30600 -5700 30660 -5080
rect 30700 -5470 30760 -4830
rect 30800 -5070 30860 -4650
rect 30900 -4840 30960 -4470
rect 31000 -4650 31060 -4230
rect 31100 -4460 31160 -4090
rect 31200 -4230 31260 -3900
rect 31300 -4040 31360 -3720
rect 31400 -3900 31460 -3570
rect 31500 -3710 31560 -3430
rect 31600 -3620 31660 -3290
rect 31700 -3470 31760 -3100
rect 31800 -3290 31860 -3000
rect 31900 -3140 31960 -2860
rect 32000 -3000 32060 -2710
rect 32100 -2850 32160 -2610
rect 32200 -2710 32260 -2470
rect 32300 -2610 32360 -2370
rect 32400 -2510 32460 -2270
rect 32500 -2370 32560 -2170
rect 32600 -2270 32660 -2070
rect 32700 -2210 32760 -1970
rect 32800 -2100 32860 -1870
rect 32900 -2020 32960 -1770
rect 33000 -2030 33060 -1720
rect 33100 -2170 33160 -1650
rect 33200 -2230 33260 -1680
rect 33500 -1700 33560 0
rect 30700 -6100 30760 -5830
rect 30800 -6070 30860 -5610
rect 30900 -6020 30960 -5340
rect 31000 -5970 31060 -4980
rect 31100 -5940 31160 -4780
rect 31200 -5890 31260 -4600
rect 31300 -5860 31360 -4360
rect 31400 -5810 31460 -4180
rect 31500 -5790 31560 -4040
rect 31600 -5750 31660 -3850
rect 31700 -5710 31760 -3750
rect 31800 -5670 31860 -3560
rect 31900 -5650 31960 -3430
rect 32000 -5620 32060 -3280
rect 32100 -5580 32160 -3130
rect 32200 -5570 32260 -2990
rect 32300 -5540 32360 -2850
rect 32400 -5530 32460 -2750
rect 32500 -5500 32560 -2650
rect 32600 -5500 32660 -2510
rect 32700 -5490 32760 -2400
rect 32800 -5450 32860 -2340
rect 32900 -5450 32960 -2270
rect 33000 -5450 33060 -2310
rect 33300 -2330 33360 -1750
rect 33600 -1800 33660 0
rect 33100 -5410 33160 -2370
rect 33400 -2430 33460 -1840
rect 33700 -1900 33760 0
rect 33200 -5410 33260 -2470
rect 33500 -2530 33560 -1940
rect 33800 -2040 33860 0
rect 33300 -5370 33360 -2570
rect 33600 -2630 33660 -2040
rect 33900 -2140 33960 0
rect 33400 -5360 33460 -2670
rect 33700 -2720 33760 -2180
rect 34000 -2280 34060 0
rect 33500 -5360 33560 -2770
rect 33800 -2820 33860 -2280
rect 34100 -2390 34160 0
rect 33600 -5320 33660 -2870
rect 33900 -2920 33960 -2420
rect 34200 -2530 34260 0
rect 33700 -5320 33760 -2970
rect 34000 -3020 34060 -2530
rect 33800 -5320 33860 -3070
rect 34100 -3140 34160 -2620
rect 34300 -2630 34360 0
rect 34400 -2730 34460 0
rect 33900 -5320 33960 -3170
rect 34000 -5320 34060 -3260
rect 34200 -3270 34260 -2770
rect 34500 -2830 34560 0
rect 34300 -3370 34360 -2870
rect 34600 -2970 34660 0
rect 34100 -5320 34160 -3410
rect 34400 -3470 34460 -2970
rect 34700 -3070 34760 0
rect 34200 -5310 34260 -3510
rect 34500 -3570 34560 -3110
rect 34800 -3180 34860 0
rect 34300 -5280 34360 -3610
rect 34600 -3670 34660 -3210
rect 34400 -5280 34460 -3710
rect 34700 -3770 34760 -3310
rect 34900 -3320 34960 0
rect 35000 -3410 35060 0
rect 34500 -5280 34560 -3810
rect 34800 -3870 34860 -3460
rect 35100 -3510 35160 0
rect 34600 -5270 34660 -3910
rect 34900 -3970 34960 -3560
rect 35200 -3660 35260 0
rect 34700 -5230 34760 -4010
rect 35000 -4070 35060 -3660
rect 35300 -3760 35360 0
rect 34800 -5230 34860 -4110
rect 35100 -4210 35160 -3800
rect 35400 -3860 35460 0
rect 34900 -5230 34960 -4250
rect 35200 -4310 35260 -3900
rect 35500 -3960 35560 0
rect 35000 -5230 35060 -4350
rect 35300 -4450 35360 -4000
rect 35600 -4060 35660 0
rect 35100 -5210 35160 -4450
rect 35400 -4550 35460 -4100
rect 35700 -4160 35760 0
rect 35200 -5190 35260 -4600
rect 35500 -4700 35560 -4200
rect 35800 -4300 35860 0
rect 35300 -5190 35360 -4700
rect 35600 -4800 35660 -4340
rect 35900 -4400 35960 0
rect 35400 -5230 35460 -4840
rect 35700 -4940 35760 -4440
rect 36000 -4500 36060 0
rect 35500 -5230 35560 -4940
rect 35600 -5240 35660 -5080
rect 35800 -5090 35860 -4540
rect 36100 -4600 36160 0
rect 35900 -5180 35960 -4640
rect 36200 -4700 36260 0
rect 35700 -5260 35760 -5180
rect 36000 -5290 36060 -4740
rect 36300 -4840 36360 0
rect 36100 -5430 36160 -4840
rect 36400 -4940 36460 0
rect 36200 -5440 36260 -4980
rect 36300 -5400 36360 -5080
rect 36500 -5090 36560 0
rect 36600 -5230 36660 0
rect 36400 -5360 36460 -5230
rect 36700 -5300 36760 0
rect 36800 -5280 36860 0
rect 36900 -5280 36960 0
rect 37000 -5280 37060 0
rect 37100 -5250 37160 0
rect 37200 -5230 37260 0
rect 37300 -5230 37360 0
rect 37400 -5230 37460 0
rect 37500 -5200 37560 0
rect 37600 -5190 37660 0
rect 37700 -5190 37760 0
rect 37800 -5190 37860 0
rect 37900 -5190 37960 0
rect 38000 -5190 38060 0
rect 38100 -5170 38160 0
rect 38200 -5120 38260 0
rect 38300 -5060 38360 0
rect 38400 -5020 38460 0
rect 38500 -4970 38560 0
rect 38600 -4940 38660 0
rect 38700 -4910 38760 0
rect 38800 -4880 38860 0
rect 38900 -4840 38960 0
rect 39000 -4800 39060 0
rect 39100 -4780 39160 0
rect 39200 -4750 39260 0
rect 39300 -4720 39360 0
rect 39400 -4710 39460 0
rect 39500 -4670 39560 0
rect 39600 -4670 39660 0
rect 39700 -4630 39760 0
rect 39800 -4620 39860 0
rect 39900 -4590 39960 0
rect 40000 -4580 40060 0
rect 40100 -4560 40160 0
rect 40200 -4540 40260 0
rect 40300 -4540 40360 0
rect 40400 -4520 40460 0
rect 40500 -4490 40560 0
rect 40600 -4490 40660 0
rect 40700 -4480 40760 0
rect 40800 -4450 40860 0
rect 40900 -4450 40960 0
rect 41000 -4450 41060 0
rect 41100 -4450 41160 0
rect 41200 -4410 41260 0
rect 41300 -4410 41360 0
rect 41400 -4410 41460 0
rect 41500 -4410 41560 0
rect 41600 -4410 41660 0
rect 41700 -4410 41760 0
rect 41800 -4370 41860 0
rect 41900 -4360 41960 0
rect 42000 -4360 42060 0
rect 42100 -4360 42160 0
rect 42200 -4360 42260 0
rect 42300 -4360 42360 0
rect 42400 -4360 42460 0
rect 42500 -4360 42560 0
rect 42600 -4360 42660 0
rect 42700 -4360 42760 0
rect 42800 -4360 42860 0
rect 42900 -4360 42960 0
rect 43000 -4360 43060 0
rect 43100 -4360 43160 0
rect 43200 -4360 43260 0
rect 43300 -4360 43360 0
rect 43400 -4400 43460 0
rect 43500 -4410 43560 0
rect 43600 -4410 43660 0
rect 43700 -4410 43760 0
rect 43800 -4410 43860 0
rect 43900 -4410 43960 0
rect 44000 -4430 44060 0
rect 44100 -4450 44160 0
rect 44200 -4450 44260 0
rect 44300 -4450 44360 0
rect 44400 -4480 44460 0
rect 44500 -4490 44560 0
rect 44600 -4490 44660 0
rect 44700 -4520 44760 0
rect 44800 -4540 44860 0
rect 44900 -4540 44960 0
rect 45000 -4580 45060 0
rect 45100 -4580 45160 0
rect 45200 -4620 45260 0
rect 45300 -4620 45360 0
rect 45400 -4650 45460 0
rect 45500 -4670 45560 0
rect 45600 -4710 45660 0
rect 45700 -4710 45760 0
rect 45800 -4750 45860 0
rect 45900 -4820 45960 0
rect 38800 -5630 38860 -5540
rect 38900 -5620 38960 -5490
rect 39000 -5660 39060 -5440
rect 39100 -5650 39160 -5390
rect 39200 -5620 39260 -5350
rect 39300 -5590 39360 -5310
rect 39400 -5570 39460 -5290
rect 39500 -5540 39560 -5260
rect 39600 -5510 39660 -5220
rect 39700 -5490 39760 -5180
rect 39800 -5450 39860 -5170
rect 39900 -5420 39960 -5130
rect 40000 -5410 40060 -5120
rect 40100 -5410 40160 -5090
rect 40200 -5360 40260 -5080
rect 40300 -5360 40360 -5040
rect 40400 -5320 40460 -5040
rect 40500 -5320 40560 -5020
rect 40600 -5320 40660 -4990
rect 40700 -5280 40760 -4990
rect 40800 -5280 40860 -4980
rect 40900 -5270 40960 -4950
rect 41000 -5230 41060 -4950
rect 41100 -5230 41160 -4950
rect 41200 -5240 41260 -4910
rect 41300 -5230 41360 -4910
rect 41400 -5190 41460 -4910
rect 41500 -5190 41560 -4910
rect 41600 -5190 41660 -4910
rect 41700 -5150 41760 -4870
rect 41800 -5150 41860 -4860
rect 41900 -5150 41960 -4860
rect 42000 -5150 42060 -4860
rect 42100 -5130 42160 -4860
rect 42200 -5100 42260 -4860
rect 42300 -5100 42360 -4860
rect 42400 -5100 42460 -4860
rect 42500 -5100 42560 -4860
rect 42600 -5100 42660 -4860
rect 42700 -5060 42760 -4860
rect 42800 -5060 42860 -4860
rect 42900 -5060 42960 -4860
rect 43000 -5060 43060 -4860
rect 43100 -5060 43160 -4860
rect 43200 -5060 43260 -4860
rect 43300 -5060 43360 -4860
rect 43400 -5060 43460 -4860
rect 43500 -5060 43560 -4900
rect 43600 -5060 43660 -4910
rect 43700 -5060 43760 -4910
rect 43800 -5060 43860 -4910
rect 43900 -5060 43960 -4910
rect 44000 -5060 44060 -4910
rect 44100 -5060 44160 -4950
rect 44200 -5060 44260 -4950
rect 44300 -5060 44360 -4950
rect 44400 -5060 44460 -4960
rect 44500 -5070 44560 -5000
rect 44600 -5100 44660 -4990
rect 44700 -5100 44760 -5000
rect 44800 -5100 44860 -5040
rect 44900 -5140 44960 -5040
rect 45000 -5170 45060 -5040
rect 39600 -5800 39660 -5690
rect 39700 -5850 39760 -5680
rect 39800 -5900 39860 -5650
rect 30400 -6590 30460 -6530
rect 30300 -8400 30360 -8260
rect 30400 -8340 30460 -8050
rect 30500 -8270 30560 -7990
rect 30600 -8180 30660 -7890
rect 30700 -8080 30760 -7800
rect 30800 -8030 30860 -7700
rect 30900 -7930 30960 -7640
rect 31000 -7840 31060 -7550
rect 31100 -7770 31160 -7450
rect 31200 -7670 31260 -7390
rect 31300 -7610 31360 -7330
rect 31400 -7530 31460 -7230
rect 31500 -7460 31560 -7170
rect 31600 -7400 31660 -7120
rect 31700 -7340 31760 -7070
rect 31800 -7290 31860 -7020
rect 31900 -7230 31960 -6990
rect 32000 -7170 32060 -6940
rect 32100 -7100 32160 -6880
rect 32200 -7050 32260 -6830
rect 32300 -7000 32360 -6790
rect 32400 -6950 32460 -6740
rect 32500 -6890 32560 -6690
rect 32600 -6850 32660 -6650
rect 32700 -6800 32760 -6610
rect 32800 -6750 32860 -6570
rect 32900 -6700 32960 -6530
rect 33000 -6650 33060 -6480
rect 33100 -6620 33160 -6450
rect 33200 -6570 33260 -6430
rect 33300 -6520 33360 -6390
rect 33400 -6490 33460 -6350
rect 33500 -6440 33560 -6300
rect 33600 -6410 33660 -6260
rect 33700 -6360 33760 -6240
rect 33800 -6320 33860 -6210
rect 33900 -6270 33960 -6170
rect 34000 -6230 34060 -6130
rect 34100 -6190 34160 -6100
rect 34200 -6160 34260 -6050
rect 34300 -6130 34360 -6030
rect 34400 -6080 34460 -5990
rect 34500 -6050 34560 -5960
rect 34600 -6010 34660 -5950
rect 34700 -5970 34760 -5910
rect 39900 -5950 39960 -5620
rect 40000 -6020 40060 -5600
rect 40100 -6070 40160 -5600
rect 40200 -6120 40260 -5560
rect 40300 -6190 40360 -5560
rect 40400 -6270 40460 -5520
rect 40500 -6340 40560 -5520
rect 40600 -6410 40660 -5510
rect 40700 -6500 40760 -5470
rect 40800 -6550 40860 -5470
rect 40900 -6650 40960 -5450
rect 41000 -6710 41060 -5430
rect 30100 -8600 30160 -8540
rect 27200 -22330 27260 -21110
rect 27400 -21240 27460 -20930
rect 27300 -22340 27360 -21600
rect 27500 -21830 27560 -14490
rect 27700 -14620 27760 -9190
rect 27600 -21880 27660 -14800
rect 27800 -14940 27860 -9390
rect 27700 -15310 27760 -15150
rect 27700 -18910 27760 -15370
rect 27900 -15700 27960 -9580
rect 27800 -18510 27860 -16050
rect 28000 -16540 28060 -9810
rect 27900 -17970 27960 -16980
rect 27900 -18830 27960 -18740
rect 27700 -19040 27760 -18970
rect 27700 -21480 27760 -19420
rect 27800 -21120 27860 -19230
rect 27900 -20670 27960 -18890
rect 28000 -20040 28060 -18280
rect 28100 -19420 28160 -10080
rect 28200 -18890 28260 -10350
rect 28300 -18270 28360 -10580
rect 28400 -16770 28460 -10940
rect 28500 -15630 28560 -11310
rect 28600 -15070 28660 -11670
rect 28700 -12230 28760 -12130
rect 28700 -15090 28760 -12290
rect 28900 -12530 28960 -12470
rect 29000 -12520 29060 -12460
rect 28800 -15620 28860 -12740
rect 28500 -17480 28560 -17420
rect 28500 -17670 28560 -17540
rect 28600 -17590 28660 -15810
rect 28700 -17130 28760 -15810
rect 28900 -16410 28960 -13100
rect 29100 -13220 29160 -12700
rect 29200 -13110 29260 -12430
rect 29300 -12870 29360 -12110
rect 29400 -12600 29460 -11880
rect 29500 -12410 29560 -11690
rect 29600 -12190 29660 -11460
rect 29700 -12000 29760 -11270
rect 29800 -11810 29860 -11130
rect 29900 -11620 29960 -10980
rect 30000 -11480 30060 -10800
rect 30100 -11290 30160 -10660
rect 30200 -11150 30260 -10520
rect 30300 -11010 30360 -10370
rect 30400 -10860 30460 -10230
rect 30500 -10720 30560 -10130
rect 30600 -10570 30660 -9980
rect 30700 -10430 30760 -9890
rect 30800 -10330 30860 -9790
rect 30900 -10190 30960 -9650
rect 31000 -10090 31060 -9550
rect 31100 -9940 31160 -9440
rect 31200 -9850 31260 -9350
rect 31300 -9750 31360 -9240
rect 31400 -9650 31460 -9150
rect 31500 -9550 31560 -9090
rect 31600 -9450 31660 -8990
rect 31700 -9340 31760 -8890
rect 31800 -9240 31860 -8820
rect 31900 -9150 31960 -8730
rect 32000 -9060 32060 -8650
rect 32100 -8990 32160 -8570
rect 32200 -8890 32260 -8510
rect 32300 -8830 32360 -8440
rect 32400 -8740 32460 -8360
rect 32500 -8660 32560 -8300
rect 32600 -8580 32660 -8220
rect 32700 -8520 32760 -8170
rect 32800 -8450 32860 -8100
rect 32900 -8370 32960 -8040
rect 33000 -8310 33060 -7990
rect 33100 -8250 33160 -7930
rect 33200 -8180 33260 -7870
rect 33300 -8110 33360 -7810
rect 33400 -8060 33460 -7760
rect 33500 -7990 33560 -7710
rect 33600 -7930 33660 -7660
rect 33700 -7890 33760 -7610
rect 33800 -7840 33860 -7560
rect 33900 -7790 33960 -7520
rect 34000 -7740 34060 -7480
rect 34100 -7680 34160 -7430
rect 34200 -7640 34260 -7390
rect 34300 -7580 34360 -7350
rect 34400 -7540 34460 -7300
rect 34500 -7510 34560 -7280
rect 34600 -7460 34660 -7250
rect 34700 -7430 34760 -7220
rect 34800 -7380 34860 -7180
rect 34900 -7360 34960 -7140
rect 35000 -7320 35060 -7120
rect 35100 -7280 35160 -7080
rect 35200 -7240 35260 -7040
rect 35300 -7220 35360 -7030
rect 35400 -7190 35460 -7000
rect 35500 -7160 35560 -6970
rect 35600 -7140 35660 -6950
rect 35700 -7100 35760 -6920
rect 35800 -7070 35860 -6910
rect 35900 -7060 35960 -6870
rect 36000 -7050 36060 -6870
rect 36100 -7020 36160 -6850
rect 36200 -7010 36260 -6820
rect 36300 -6970 36360 -6820
rect 36400 -6980 36460 -6780
rect 36500 -6950 36560 -6780
rect 36600 -6930 36660 -6780
rect 36700 -6930 36760 -6770
rect 36800 -6900 36860 -6730
rect 36900 -6890 36960 -6740
rect 37000 -6890 37060 -6730
rect 37100 -6890 37160 -6730
rect 37200 -6890 37260 -6730
rect 37300 -6890 37360 -6730
rect 37400 -6870 37460 -6730
rect 37500 -6840 37560 -6730
rect 37600 -6840 37660 -6730
rect 37700 -6840 37760 -6730
rect 37800 -6840 37860 -6730
rect 37900 -6850 37960 -6730
rect 38000 -6890 38060 -6730
rect 38100 -6890 38160 -6730
rect 38200 -6890 38260 -6730
rect 38300 -6890 38360 -6730
rect 38400 -6890 38460 -6740
rect 38500 -6910 38560 -6780
rect 38600 -6930 38660 -6780
rect 38700 -6930 38760 -6780
rect 41100 -6790 41160 -5430
rect 38800 -6930 38860 -6800
rect 38900 -6970 38960 -6820
rect 39000 -6970 39060 -6820
rect 41200 -6860 41260 -5430
rect 39100 -7010 39160 -6870
rect 39200 -7020 39260 -6870
rect 39300 -7050 39360 -6900
rect 39400 -7060 39460 -6910
rect 41300 -6930 41360 -5400
rect 39500 -7080 39560 -6950
rect 39600 -7110 39660 -6960
rect 39700 -7150 39760 -7000
rect 41400 -7020 41460 -5380
rect 39800 -7160 39860 -7020
rect 39900 -7190 39960 -7050
rect 40000 -7230 40060 -7080
rect 41500 -7120 41560 -5390
rect 40100 -7270 40160 -7120
rect 40200 -7300 40260 -7150
rect 40300 -7330 40360 -7180
rect 41600 -7190 41660 -5380
rect 40400 -7380 40460 -7230
rect 40500 -7410 40560 -7260
rect 41700 -7280 41760 -5340
rect 40600 -7460 40660 -7310
rect 40700 -7500 40760 -7360
rect 41800 -7370 41860 -5340
rect 40800 -7530 40860 -7400
rect 40900 -7580 40960 -7460
rect 41900 -7480 41960 -5340
rect 41000 -7630 41060 -7510
rect 42000 -7540 42060 -5340
rect 41100 -7680 41160 -7560
rect 41200 -7730 41260 -7610
rect 42100 -7630 42160 -5300
rect 41300 -7790 41360 -7650
rect 42200 -7730 42260 -5300
rect 41400 -7850 41460 -7730
rect 41500 -7900 41560 -7780
rect 42300 -7830 42360 -5300
rect 41600 -7960 41660 -7850
rect 41700 -8020 41760 -7910
rect 42000 -7940 42060 -7880
rect 41800 -8100 41860 -7970
rect 42100 -7980 42160 -7880
rect 42400 -7930 42460 -5300
rect 41900 -8180 41960 -8060
rect 42200 -8080 42260 -7970
rect 42500 -8030 42560 -5300
rect 42600 -8100 42660 -5300
rect 42000 -8230 42060 -8120
rect 42100 -8280 42160 -8220
rect 42700 -8230 42760 -5260
rect 42200 -8380 42260 -8280
rect 42500 -8310 42560 -8230
rect 42800 -8330 42860 -5250
rect 42300 -8440 42360 -8370
rect 42900 -8430 42960 -5250
rect 43000 -8530 43060 -5260
rect 43100 -8630 43160 -5260
rect 43200 -8710 43260 -5250
rect 43300 -8690 43360 -5250
rect 43400 -8540 43460 -5260
rect 43500 -8440 43560 -5250
rect 43600 -8340 43660 -5250
rect 43700 -8150 43760 -5250
rect 43800 -8010 43860 -5250
rect 43900 -7830 43960 -5260
rect 44000 -7590 44060 -5260
rect 44100 -7410 44160 -5260
rect 44200 -7180 44260 -5260
rect 44300 -6950 44360 -5260
rect 44400 -6540 44460 -5250
rect 44500 -6270 44560 -5260
rect 44600 -6040 44660 -5300
rect 44700 -5680 44760 -5300
rect 44800 -5400 44860 -5310
rect 43400 -9060 43460 -8820
rect 43500 -9210 43560 -8680
rect 43600 -9270 43660 -8580
rect 43700 -9150 43760 -8440
rect 43800 -9060 43860 -8290
rect 43900 -8910 43960 -8150
rect 44000 -8770 44060 -7960
rect 44100 -8580 44160 -7770
rect 44200 -8440 44260 -7540
rect 44300 -8250 44360 -7310
rect 44400 -8020 44460 -7090
rect 44500 -7840 44560 -6810
rect 44600 -7660 44660 -6450
rect 44700 -7420 44760 -6180
rect 44800 -7190 44860 -5950
rect 44900 -6910 44960 -5580
rect 45000 -6690 45060 -5400
rect 45100 -6320 45160 -5080
rect 45200 -6050 45260 -5080
rect 45300 -5780 45360 -5120
rect 45400 -5410 45460 -5130
rect 45200 -6530 45260 -6470
rect 43700 -9540 43760 -9440
rect 43800 -9720 43860 -9340
rect 43900 -9890 43960 -9200
rect 44000 -10050 44060 -9050
rect 44100 -10240 44160 -8910
rect 44200 -10430 44260 -8720
rect 44300 -10620 44360 -8580
rect 44100 -10760 44160 -10660
rect 44200 -10970 44260 -10750
rect 44400 -10800 44460 -8390
rect 44300 -10990 44360 -10930
rect 44500 -10990 44560 -8210
rect 44600 -11310 44660 -7970
rect 44700 -11620 44760 -7790
rect 44800 -12030 44860 -7550
rect 44900 -12610 44960 -7320
rect 45000 -13010 45060 -7100
rect 28900 -16730 28960 -16470
rect 28700 -17310 28760 -17190
rect 28900 -17280 28960 -16790
rect 29000 -17190 29060 -13500
rect 45100 -13640 45160 -6820
rect 29100 -16860 29160 -14220
rect 29200 -16190 29260 -14700
rect 32800 -16510 32860 -15320
rect 32900 -16580 32960 -14440
rect 33000 -16630 33060 -13930
rect 36200 -14340 36260 -14280
rect 33100 -16680 33160 -15300
rect 33200 -16730 33260 -15350
rect 33300 -16760 33360 -15310
rect 33400 -16800 33460 -15310
rect 33500 -16840 33560 -15310
rect 33600 -16860 33660 -15310
rect 33700 -16900 33760 -15310
rect 33800 -16940 33860 -15340
rect 33900 -16970 33960 -15350
rect 34000 -16980 34060 -15390
rect 34100 -17020 34160 -15400
rect 34200 -17030 34260 -15440
rect 34300 -17040 34360 -15480
rect 34400 -17070 34460 -15550
rect 35600 -15590 35660 -15480
rect 34500 -17100 34560 -15600
rect 34600 -17110 34660 -15660
rect 34700 -17150 34760 -15700
rect 34800 -17160 34860 -15700
rect 34900 -17190 34960 -15690
rect 35000 -17200 35060 -15660
rect 35100 -17240 35160 -15660
rect 35200 -17240 35260 -15660
rect 32800 -17420 32860 -17240
rect 35300 -17280 35360 -15660
rect 32900 -17410 32960 -17280
rect 35400 -17290 35460 -15680
rect 35500 -17320 35560 -15780
rect 35600 -17330 35660 -15800
rect 35700 -17330 35760 -15260
rect 35800 -15700 35860 -15070
rect 35900 -15520 35960 -14880
rect 36000 -15190 36060 -14700
rect 36100 -14920 36160 -14510
rect 36200 -14520 36260 -14410
rect 36200 -14640 36260 -14580
rect 33000 -17390 33060 -17330
rect 35800 -17350 35860 -15860
rect 35900 -17380 35960 -15870
rect 36000 -17370 36060 -15820
rect 36100 -17400 36160 -15750
rect 32800 -18720 32860 -17750
rect 32900 -20000 32960 -17750
rect 28000 -20220 28060 -20100
rect 28900 -20380 28960 -20320
rect 27900 -21420 27960 -21340
rect 27700 -21600 27760 -21540
rect 27400 -22370 27460 -22180
rect 27600 -22440 27660 -22380
rect 26600 -23230 26660 -22460
rect 26800 -23290 26860 -22460
rect 26900 -23300 26960 -22490
rect 27000 -23370 27060 -22490
rect 26000 -26870 26060 -23700
rect 26100 -26820 26160 -23750
rect 26200 -26730 26260 -23610
rect 26300 -26660 26360 -23580
rect 26400 -26560 26460 -23550
rect 26500 -26470 26560 -23530
rect 26600 -26400 26660 -23540
rect 26700 -26310 26760 -23500
rect 26800 -26240 26860 -23490
rect 26900 -26150 26960 -23500
rect 27100 -23560 27160 -22490
rect 27700 -22500 27760 -22060
rect 27000 -25920 27060 -23690
rect 27200 -23870 27260 -22510
rect 27200 -23990 27260 -23930
rect 27200 -24120 27260 -24050
rect 27200 -24240 27260 -24180
rect 27200 -25850 27260 -25610
rect 27000 -26040 27060 -25980
rect 26700 -26680 26760 -26550
rect 22200 -39760 22260 -38750
rect 22500 -38810 22560 -31430
rect 22300 -39400 22360 -38840
rect 22600 -38860 22660 -31700
rect 22400 -39180 22460 -38950
rect 22700 -38960 22760 -31720
rect 22500 -39060 22560 -39000
rect 22800 -39040 22860 -31570
rect 22900 -39110 22960 -31390
rect 23000 -39170 23060 -31240
rect 22300 -39520 22360 -39460
rect 20700 -43360 20760 -43290
rect 18600 -48580 18660 -45470
rect 18700 -48580 18760 -45460
rect 18800 -48580 18860 -45360
rect 18900 -48580 18960 -45260
rect 19000 -48580 19060 -45200
rect 19100 -48580 19160 -45100
rect 19200 -48580 19260 -45030
rect 19300 -48580 19360 -44960
rect 19400 -48580 19460 -44900
rect 19500 -48580 19560 -44790
rect 19600 -48580 19660 -44690
rect 19700 -48580 19760 -44590
rect 19800 -48580 19860 -44490
rect 19900 -48580 19960 -44340
rect 20000 -48580 20060 -44210
rect 20100 -48580 20160 -44110
rect 20200 -48580 20260 -43960
rect 20300 -48580 20360 -43860
rect 20400 -48580 20460 -43720
rect 20500 -48580 20560 -43570
rect 20600 -48580 20660 -43560
rect 20800 -43590 20860 -43100
rect 20700 -48580 20760 -43730
rect 20900 -43780 20960 -42910
rect 20800 -48580 20860 -43910
rect 21000 -43920 21060 -42770
rect 20900 -48580 20960 -44060
rect 21100 -44120 21160 -42560
rect 21000 -48580 21060 -44250
rect 21200 -44260 21260 -42350
rect 21300 -44350 21360 -42160
rect 21100 -48580 21160 -44390
rect 21400 -44490 21460 -41980
rect 21200 -48580 21260 -44500
rect 21500 -44640 21560 -41750
rect 21300 -48580 21360 -44640
rect 21600 -44740 21660 -41560
rect 21400 -48580 21460 -44780
rect 21700 -44880 21760 -41370
rect 21500 -48580 21560 -44880
rect 21600 -48580 21660 -45020
rect 21800 -45030 21860 -41160
rect 21900 -45130 21960 -40950
rect 21700 -48580 21760 -45170
rect 22000 -45220 22060 -40770
rect 22100 -45230 22160 -40540
rect 22200 -45230 22260 -40180
rect 22300 -45230 22360 -39900
rect 21800 -48580 21860 -45270
rect 21900 -48580 21960 -45370
rect 22000 -48580 22060 -45420
rect 22100 -48580 22160 -45430
rect 22200 -48580 22260 -45430
rect 22300 -48580 22360 -45380
rect 22400 -48580 22460 -39620
rect 22500 -48580 22560 -39310
rect 22600 -48580 22660 -39180
rect 22700 -48580 22760 -39190
rect 23100 -39230 23160 -31060
rect 22800 -48580 22860 -39260
rect 23200 -39310 23260 -30910
rect 22900 -48580 22960 -39320
rect 23000 -48580 23060 -39370
rect 23300 -39390 23360 -30810
rect 23100 -48580 23160 -39460
rect 23400 -39480 23460 -30750
rect 23200 -48580 23260 -39520
rect 23500 -39560 23560 -30680
rect 23600 -39500 23660 -30630
rect 23700 -39400 23760 -30580
rect 23800 -39300 23860 -30500
rect 23900 -39200 23960 -30430
rect 24000 -39060 24060 -30360
rect 24100 -38870 24160 -30270
rect 24200 -38680 24260 -30180
rect 24300 -38540 24360 -30070
rect 24400 -38350 24460 -29980
rect 24500 -38160 24560 -29870
rect 24600 -38130 24660 -29770
rect 24700 -38050 24760 -29680
rect 24800 -38100 24860 -29620
rect 24900 -38150 24960 -29520
rect 25000 -38250 25060 -29450
rect 23300 -48580 23360 -39630
rect 23400 -48580 23460 -39730
rect 23500 -48580 23560 -39770
rect 23600 -48580 23660 -39740
rect 23700 -48580 23760 -39640
rect 23800 -48580 23860 -39540
rect 23900 -48580 23960 -39440
rect 24000 -48580 24060 -39340
rect 24100 -48580 24160 -39200
rect 24200 -48580 24260 -39010
rect 24300 -48580 24360 -38820
rect 24400 -48580 24460 -38680
rect 24500 -48580 24560 -38490
rect 24600 -48580 24660 -38300
rect 24700 -48580 24760 -38250
rect 24800 -48580 24860 -38290
rect 25100 -38400 25160 -29360
rect 24900 -48580 24960 -38400
rect 25200 -38420 25260 -29260
rect 25300 -38160 25360 -29160
rect 25400 -37880 25460 -29060
rect 25500 -37610 25560 -28920
rect 25600 -30490 25660 -28730
rect 25700 -30500 25760 -28590
rect 25800 -30520 25860 -28400
rect 25600 -37110 25660 -30740
rect 25900 -30970 25960 -28120
rect 25700 -36880 25760 -30970
rect 26000 -31120 26060 -27060
rect 26100 -29350 26160 -27030
rect 26200 -28900 26260 -26960
rect 26300 -28450 26360 -26890
rect 26400 -27730 26460 -26800
rect 26500 -27030 26560 -26770
rect 26700 -27120 26760 -26800
rect 26800 -27130 26860 -26450
rect 26900 -27180 26960 -26390
rect 27000 -27240 27060 -26290
rect 27100 -27280 27160 -26150
rect 27200 -27330 27260 -25910
rect 27300 -27360 27360 -22530
rect 27400 -27420 27460 -22570
rect 27800 -22590 27860 -21790
rect 27500 -27440 27560 -22590
rect 27600 -27490 27660 -22640
rect 27900 -22650 27960 -21480
rect 28000 -22710 28060 -21110
rect 27700 -27540 27760 -22720
rect 27800 -27590 27860 -22800
rect 28100 -22850 28160 -21180
rect 28400 -21300 28460 -21240
rect 27900 -27660 27960 -22860
rect 28000 -27720 28060 -22950
rect 28200 -22960 28260 -21320
rect 28300 -23050 28360 -21460
rect 28100 -27780 28160 -23090
rect 28400 -23150 28460 -21620
rect 28200 -27870 28260 -23190
rect 28500 -23240 28560 -21620
rect 28300 -27890 28360 -23290
rect 28600 -23310 28660 -21210
rect 28400 -27610 28460 -23390
rect 28700 -23410 28760 -21020
rect 28500 -27290 28560 -23450
rect 28800 -23520 28860 -20750
rect 28900 -23540 28960 -20440
rect 29000 -23440 29060 -20110
rect 29100 -23350 29160 -20210
rect 29200 -23240 29260 -20450
rect 29300 -23150 29360 -20640
rect 29400 -23050 29460 -20830
rect 29500 -22990 29560 -20930
rect 29600 -22890 29660 -21030
rect 29700 -22790 29760 -21050
rect 29800 -22600 29860 -21010
rect 29900 -22500 29960 -20960
rect 30000 -22470 30060 -20810
rect 30100 -22470 30160 -20620
rect 30200 -22470 30260 -20340
rect 30300 -22470 30360 -20250
rect 33000 -20260 33060 -17790
rect 33100 -20320 33160 -17790
rect 33200 -20380 33260 -17830
rect 35800 -17840 35860 -17750
rect 33300 -20460 33360 -17850
rect 30400 -20540 30460 -20480
rect 30400 -22470 30460 -20600
rect 33000 -20670 33060 -20500
rect 30500 -22470 30560 -20790
rect 30600 -22470 30660 -20930
rect 33000 -20970 33060 -20730
rect 30700 -22470 30760 -21120
rect 30800 -22470 30860 -21310
rect 30900 -22470 30960 -21500
rect 33100 -21530 33160 -20530
rect 33400 -20540 33460 -17880
rect 33500 -20600 33560 -17880
rect 33600 -20650 33660 -17920
rect 33200 -21430 33260 -20660
rect 33700 -20720 33760 -17920
rect 33800 -20800 33860 -17950
rect 33500 -21070 33560 -20840
rect 33900 -20850 33960 -17960
rect 31000 -22470 31060 -21680
rect 31100 -22470 31160 -21870
rect 31200 -22470 31260 -22010
rect 31300 -22470 31360 -22110
rect 31400 -22470 31460 -22290
rect 31500 -22510 31560 -22450
rect 32000 -22570 32060 -22370
rect 32100 -22630 32160 -22360
rect 28600 -27020 28660 -23550
rect 28700 -26680 28760 -23660
rect 29100 -23730 29160 -23580
rect 28900 -23970 28960 -23910
rect 28800 -26300 28860 -24180
rect 29000 -24390 29060 -23890
rect 28900 -25770 28960 -24720
rect 28900 -26550 28960 -26490
rect 26200 -30650 26260 -29920
rect 26100 -31200 26160 -30880
rect 26300 -31150 26360 -29080
rect 25800 -36650 25860 -31370
rect 26000 -31640 26060 -31470
rect 25900 -36290 25960 -31910
rect 26100 -32210 26160 -31500
rect 26000 -32620 26060 -32560
rect 26000 -32750 26060 -32680
rect 26000 -35530 26060 -32810
rect 26200 -32840 26260 -31600
rect 26200 -33000 26260 -32900
rect 26200 -33170 26260 -33060
rect 26200 -33290 26260 -33230
rect 26200 -35300 26260 -35130
rect 26200 -35470 26260 -35410
rect 26000 -35650 26060 -35590
rect 26000 -35770 26060 -35710
rect 26200 -36050 26260 -35530
rect 26300 -36030 26360 -31670
rect 26400 -35570 26460 -28680
rect 26500 -35300 26560 -28220
rect 26600 -34990 26660 -28190
rect 26700 -34580 26760 -28240
rect 28400 -28250 28460 -28020
rect 26800 -34250 26860 -28280
rect 26900 -33900 26960 -28300
rect 27000 -33670 27060 -28330
rect 27100 -33440 27160 -28370
rect 27200 -33210 27260 -28410
rect 27300 -32980 27360 -28460
rect 27400 -32530 27460 -28510
rect 27500 -31780 27560 -28550
rect 27600 -30980 27660 -28610
rect 27700 -29840 27760 -28680
rect 27800 -29080 27860 -28760
rect 27700 -30070 27760 -29930
rect 27700 -30190 27760 -30130
rect 26100 -36140 26160 -36080
rect 25600 -37320 25660 -37260
rect 25300 -38280 25360 -38220
rect 25000 -48580 25060 -38540
rect 25100 -48580 25160 -38730
rect 25200 -48580 25260 -38850
rect 25300 -48580 25360 -38780
rect 25400 -48580 25460 -38380
rect 25500 -48580 25560 -38090
rect 25600 -48580 25660 -37780
rect 25700 -48580 25760 -37640
rect 25800 -48580 25860 -37450
rect 25900 -48580 25960 -37220
rect 26000 -48580 26060 -37080
rect 26100 -48580 26160 -36850
rect 26200 -48580 26260 -36580
rect 26300 -45720 26360 -36580
rect 26400 -45670 26460 -36680
rect 26500 -45610 26560 -36820
rect 26600 -45530 26660 -36910
rect 26700 -45480 26760 -37060
rect 26800 -45350 26860 -37200
rect 26900 -45270 26960 -37340
rect 27000 -45200 27060 -37500
rect 27100 -45150 27160 -37680
rect 27200 -45080 27260 -37860
rect 27500 -38060 27560 -35280
rect 27300 -45030 27360 -38060
rect 27600 -38290 27660 -33960
rect 27400 -44980 27460 -38370
rect 27500 -44920 27560 -38430
rect 27700 -38470 27760 -33380
rect 27800 -38610 27860 -32840
rect 27600 -44860 27660 -38610
rect 27700 -44800 27760 -38750
rect 27900 -38800 27960 -32130
rect 27800 -44740 27860 -38940
rect 28000 -38990 28060 -30680
rect 27900 -44680 27960 -39130
rect 28100 -39180 28160 -29890
rect 28000 -44640 28060 -39310
rect 28200 -39360 28260 -29180
rect 28100 -44570 28160 -39550
rect 28300 -39590 28360 -28560
rect 28200 -41750 28260 -39730
rect 28400 -39780 28460 -28540
rect 28300 -41770 28360 -39910
rect 28500 -39970 28560 -27840
rect 28200 -44480 28260 -41950
rect 28400 -42040 28460 -40150
rect 28600 -40200 28660 -27480
rect 28300 -44400 28360 -42180
rect 28500 -42270 28560 -40380
rect 28700 -40430 28760 -27160
rect 28600 -42310 28660 -40610
rect 28800 -40700 28860 -26880
rect 28700 -42360 28760 -40860
rect 28900 -40940 28960 -26610
rect 28800 -42430 28860 -41160
rect 29000 -41250 29060 -26070
rect 28400 -44280 28460 -42460
rect 28900 -42490 28960 -41430
rect 29100 -41530 29160 -23920
rect 29000 -42570 29060 -41700
rect 29200 -41890 29260 -23480
rect 29200 -42050 29260 -41990
rect 28500 -44210 28560 -42640
rect 28700 -42740 28760 -42620
rect 28600 -44130 28660 -42870
rect 28800 -42960 28860 -42640
rect 29100 -42650 29160 -42200
rect 29300 -42420 29360 -23380
rect 28700 -43200 28760 -43140
rect 28700 -44050 28760 -43260
rect 28900 -43280 28960 -42700
rect 28800 -43970 28860 -43550
rect 29000 -43690 29060 -42800
rect 29100 -43790 29160 -42850
rect 29200 -43740 29260 -42900
rect 29300 -43670 29360 -42900
rect 29400 -43600 29460 -23280
rect 29500 -43530 29560 -23200
rect 29600 -43460 29660 -23130
rect 29700 -43390 29760 -23030
rect 29800 -43320 29860 -22930
rect 29900 -43240 29960 -22830
rect 30000 -43170 30060 -22750
rect 30100 -43100 30160 -22680
rect 30200 -43030 30260 -22660
rect 30300 -42950 30360 -22660
rect 30400 -28130 30460 -22660
rect 30500 -28200 30560 -22660
rect 30600 -28250 30660 -22670
rect 30700 -28290 30760 -22710
rect 30800 -28340 30860 -22710
rect 30400 -42880 30460 -28350
rect 30900 -28400 30960 -22710
rect 30500 -42800 30560 -28400
rect 31000 -28450 31060 -22710
rect 30600 -42730 30660 -28450
rect 31100 -28500 31160 -22710
rect 30700 -42660 30760 -28500
rect 31200 -28520 31260 -22710
rect 30800 -42580 30860 -28550
rect 31300 -28570 31360 -22750
rect 30900 -42500 30960 -28600
rect 31400 -28630 31460 -22750
rect 31000 -42430 31060 -28650
rect 31500 -28680 31560 -22750
rect 31100 -42350 31160 -28710
rect 31200 -42280 31260 -28720
rect 31600 -28730 31660 -22750
rect 31700 -28770 31760 -22770
rect 31800 -25520 31860 -22850
rect 31900 -25560 31960 -22870
rect 31300 -34600 31360 -28780
rect 31800 -28820 31860 -25790
rect 32000 -25800 32060 -22800
rect 32100 -25890 32160 -22790
rect 31400 -34450 31460 -28830
rect 31900 -28870 31960 -25930
rect 32200 -25990 32260 -22440
rect 31500 -34300 31560 -28880
rect 32000 -28920 32060 -26030
rect 32300 -26100 32360 -22590
rect 31600 -34210 31660 -28930
rect 32100 -28980 32160 -26130
rect 32400 -26190 32460 -22690
rect 33300 -22700 33360 -22220
rect 31700 -34110 31760 -28980
rect 31800 -33960 31860 -29030
rect 32200 -29040 32260 -26230
rect 32500 -26290 32560 -22740
rect 31900 -33870 31960 -29080
rect 32300 -29090 32360 -26330
rect 32600 -26390 32660 -22810
rect 33300 -22830 33360 -22770
rect 32000 -33770 32060 -29130
rect 32400 -29150 32460 -26430
rect 32700 -26490 32760 -22880
rect 33300 -22960 33360 -22900
rect 32100 -33670 32160 -29180
rect 32500 -29200 32560 -26530
rect 32800 -26590 32860 -22960
rect 33400 -22990 33460 -21850
rect 32200 -33570 32260 -29240
rect 32600 -29260 32660 -26630
rect 32300 -33460 32360 -29300
rect 32700 -29320 32760 -26730
rect 32900 -26740 32960 -23010
rect 33500 -23030 33560 -21370
rect 33600 -23070 33660 -20880
rect 34000 -20900 34060 -17960
rect 33000 -26830 33060 -23070
rect 33700 -23120 33760 -20930
rect 34100 -20940 34160 -17970
rect 32400 -33360 32460 -29350
rect 32800 -29380 32860 -26880
rect 33100 -26930 33160 -23150
rect 33800 -23160 33860 -21000
rect 34200 -21020 34260 -18010
rect 33900 -23210 33960 -21050
rect 34300 -21070 34360 -18010
rect 32500 -33310 32560 -29410
rect 32900 -29440 32960 -26980
rect 32600 -33210 32660 -29470
rect 33000 -29490 33060 -27070
rect 33200 -27080 33260 -23230
rect 34000 -23260 34060 -21100
rect 34400 -21110 34460 -18010
rect 34500 -21160 34560 -18010
rect 33300 -27180 33360 -23290
rect 34100 -23340 34160 -21170
rect 32700 -33130 32760 -29520
rect 33100 -29560 33160 -27220
rect 33400 -27320 33460 -23360
rect 34200 -23380 34260 -21220
rect 34600 -21240 34660 -18010
rect 34700 -21260 34760 -18010
rect 34300 -23430 34360 -21270
rect 34800 -21320 34860 -18050
rect 32800 -33050 32860 -29590
rect 33200 -29640 33260 -27360
rect 32900 -32960 32960 -29640
rect 33300 -29700 33360 -27460
rect 33500 -27470 33560 -23440
rect 34400 -23490 34460 -21320
rect 34900 -21380 34960 -18050
rect 33600 -27610 33660 -23500
rect 33000 -32900 33060 -29710
rect 33400 -29760 33460 -27610
rect 33700 -27750 33760 -23560
rect 34000 -23580 34060 -23500
rect 33100 -32820 33160 -29790
rect 33200 -32750 33260 -29840
rect 33500 -29860 33560 -27750
rect 33300 -32680 33360 -29910
rect 33600 -29920 33660 -27890
rect 33800 -27900 33860 -23650
rect 34100 -23670 34160 -23540
rect 34500 -23560 34560 -21390
rect 35000 -21420 35060 -18050
rect 33900 -27990 33960 -23710
rect 34200 -23730 34260 -23590
rect 34600 -23610 34660 -21440
rect 35100 -21460 35160 -18050
rect 33400 -32630 33460 -30000
rect 33700 -30010 33760 -27990
rect 34000 -28130 34060 -23810
rect 34300 -23820 34360 -23640
rect 34700 -23680 34760 -21470
rect 35200 -21510 35260 -18050
rect 34400 -23880 34460 -23710
rect 34800 -23760 34860 -21520
rect 35300 -21560 35360 -18050
rect 33500 -32560 33560 -30070
rect 33800 -30110 33860 -28130
rect 34100 -28280 34160 -23890
rect 33600 -32480 33660 -30150
rect 33700 -32410 33760 -30250
rect 33800 -32360 33860 -30350
rect 33900 -32300 33960 -28280
rect 34000 -32240 34060 -28420
rect 34200 -28430 34260 -23960
rect 34500 -23980 34560 -23760
rect 34900 -23800 34960 -21580
rect 35400 -21600 35460 -18050
rect 34100 -32190 34160 -28560
rect 34300 -28570 34360 -24060
rect 34600 -24080 34660 -23830
rect 35000 -23870 35060 -21620
rect 35500 -21640 35560 -18050
rect 35600 -21670 35660 -18050
rect 34400 -28710 34460 -24150
rect 34700 -24160 34760 -23900
rect 35100 -23920 35160 -21670
rect 35700 -21720 35760 -18010
rect 34200 -32130 34260 -28710
rect 34300 -32070 34360 -28850
rect 34500 -28860 34560 -24220
rect 34800 -24240 34860 -23960
rect 35200 -23990 35260 -21720
rect 34600 -28950 34660 -24320
rect 34900 -24340 34960 -24010
rect 35300 -24040 35360 -21750
rect 35800 -21770 35860 -18010
rect 34400 -32020 34460 -28990
rect 34500 -31960 34560 -29090
rect 34700 -29100 34760 -24410
rect 35000 -24430 35060 -24070
rect 35400 -24140 35460 -21790
rect 35900 -21800 35960 -17700
rect 36000 -21770 36060 -17650
rect 36100 -21770 36160 -17570
rect 36200 -21770 36260 -15670
rect 36300 -21770 36360 -15620
rect 36400 -21770 36460 -15550
rect 36500 -21770 36560 -15450
rect 36600 -20340 36660 -15390
rect 36700 -20330 36760 -15300
rect 36800 -20360 36860 -15200
rect 36900 -20380 36960 -15100
rect 37000 -15930 37060 -15060
rect 37000 -20380 37060 -16140
rect 37100 -20420 37160 -16180
rect 37200 -20420 37260 -16180
rect 37300 -20420 37360 -16180
rect 37400 -20430 37460 -16200
rect 37500 -20490 37560 -16220
rect 36700 -20690 36760 -20560
rect 36800 -20800 36860 -20560
rect 36900 -20810 36960 -20580
rect 37000 -20750 37060 -20570
rect 37100 -20710 37160 -20600
rect 36600 -21730 36660 -20840
rect 36700 -21730 36760 -20920
rect 36800 -21720 36860 -20980
rect 36900 -21680 36960 -21000
rect 37000 -21680 37060 -20960
rect 37100 -21660 37160 -20910
rect 37200 -21640 37260 -20850
rect 37300 -21640 37360 -20780
rect 37400 -21600 37460 -20710
rect 37500 -21590 37560 -20630
rect 37600 -21550 37660 -16220
rect 37700 -21550 37760 -16220
rect 37800 -21510 37860 -16250
rect 39800 -16290 39860 -16230
rect 37900 -21510 37960 -16300
rect 38000 -21470 38060 -16350
rect 38100 -21440 38160 -16360
rect 38200 -21420 38260 -16400
rect 38300 -21420 38360 -16400
rect 38400 -21380 38460 -16440
rect 38500 -21350 38560 -16490
rect 38600 -21330 38660 -16540
rect 38700 -21300 38760 -16590
rect 38800 -21290 38860 -16620
rect 38900 -18040 38960 -16610
rect 39000 -18030 39060 -16650
rect 39100 -18040 39160 -16660
rect 39200 -18070 39260 -16660
rect 39300 -18110 39360 -16650
rect 39400 -18120 39460 -16620
rect 39500 -18150 39560 -16600
rect 39600 -18160 39660 -16540
rect 38900 -21250 38960 -18170
rect 39700 -18200 39760 -16390
rect 39800 -18200 39860 -16350
rect 39900 -18200 39960 -16750
rect 40000 -18210 40060 -16700
rect 40100 -18250 40160 -16620
rect 40200 -18250 40260 -16550
rect 40300 -18250 40360 -16480
rect 40400 -18250 40460 -16430
rect 40500 -18250 40560 -16380
rect 40600 -18250 40660 -16310
rect 40700 -18250 40760 -16260
rect 40800 -18250 40860 -16180
rect 40900 -18250 40960 -16110
rect 41000 -18250 41060 -16010
rect 41100 -18250 41160 -15910
rect 41200 -16920 41260 -15850
rect 44400 -16300 44460 -16240
rect 41200 -18220 41260 -17310
rect 41300 -18200 41360 -17310
rect 41400 -18160 41460 -17270
rect 41500 -18010 41560 -17250
rect 41600 -17860 41660 -17220
rect 41700 -17640 41760 -17170
rect 41800 -17410 41860 -17130
rect 41900 -17170 41960 -17110
rect 43600 -18320 43660 -18070
rect 43700 -18250 43760 -17580
rect 43800 -18160 43860 -17390
rect 43900 -18010 43960 -17200
rect 44000 -17860 44060 -17060
rect 44100 -17590 44160 -16920
rect 44200 -17360 44260 -16670
rect 44300 -17040 44360 -16500
rect 44400 -16530 44460 -16370
rect 39000 -21240 39060 -18450
rect 39100 -21200 39160 -18510
rect 39200 -21180 39260 -18560
rect 39300 -21160 39360 -18630
rect 39400 -21120 39460 -18680
rect 41100 -18690 41160 -18620
rect 41200 -18700 41260 -18630
rect 39500 -21070 39560 -18710
rect 39600 -21020 39660 -18760
rect 39700 -20980 39760 -18800
rect 39800 -20900 39860 -18860
rect 39900 -20830 39960 -18880
rect 40000 -20780 40060 -18920
rect 40100 -20670 40160 -18920
rect 40200 -20580 40260 -18960
rect 40300 -20380 40360 -18960
rect 40400 -20290 40460 -18960
rect 40500 -20140 40560 -18990
rect 40600 -20000 40660 -19010
rect 40700 -19900 40760 -19010
rect 40800 -19720 40860 -19010
rect 40900 -19530 40960 -19050
rect 41000 -19250 41060 -19050
rect 43400 -19620 43460 -19140
rect 43500 -19580 43560 -18710
rect 43600 -19510 43660 -18660
rect 43700 -19460 43760 -18610
rect 43800 -19400 43860 -18520
rect 43900 -19340 43960 -18510
rect 44000 -19290 44060 -18460
rect 44100 -19240 44160 -18350
rect 44200 -19180 44260 -18220
rect 44300 -19130 44360 -18060
rect 44400 -19080 44460 -17970
rect 44500 -19030 44560 -17820
rect 44600 -18980 44660 -17670
rect 44700 -18930 44760 -17490
rect 44800 -18880 44860 -17310
rect 44900 -18840 44960 -16820
rect 45000 -18780 45060 -16360
rect 45100 -18730 45160 -15750
rect 45200 -18690 45260 -6590
rect 45300 -18650 45360 -6230
rect 45400 -18600 45460 -5960
rect 45500 -18570 45560 -5680
rect 45600 -18520 45660 -5280
rect 45700 -18480 45760 -5010
rect 45800 -18440 45860 -4950
rect 45900 -18410 45960 -4880
rect 46000 -18370 46060 0
rect 46100 -18330 46160 0
rect 46200 -18300 46260 0
rect 46300 -18400 46360 0
rect 46400 -18500 46460 0
rect 46500 -18630 46560 0
rect 46600 -18770 46660 0
rect 46700 -18900 46760 0
rect 46800 -19000 46860 0
rect 46900 -19170 46960 0
rect 47000 -19300 47060 0
rect 47100 -19430 47160 0
rect 47200 -19520 47260 0
rect 47300 -19690 47360 0
rect 47400 -19850 47460 0
rect 47500 -17980 47560 0
rect 47600 -17980 47660 0
rect 47700 -17970 47760 0
rect 47800 -17960 47860 0
rect 47900 -17960 47960 0
rect 48000 -17960 48060 0
rect 48100 -17980 48160 0
rect 48200 -17980 48260 0
rect 48300 -17980 48360 0
rect 48400 -11890 48460 0
rect 48500 -11890 48560 0
rect 48600 -11890 48660 0
rect 48700 -11890 48760 0
rect 48800 -11890 48860 0
rect 48900 -11890 48960 0
rect 49000 -11890 49060 0
rect 49100 -11890 49160 0
rect 49200 -11890 49260 0
rect 49300 -11890 49360 0
rect 49400 -11890 49460 0
rect 49500 -11890 49560 0
rect 49600 -11890 49660 0
rect 49700 -11890 49760 0
rect 49800 -11890 49860 0
rect 49900 -11890 49960 0
rect 50000 -11890 50060 0
rect 50100 -11890 50160 0
rect 50200 -11890 50260 0
rect 50300 -11890 50360 0
rect 50400 -11890 50460 0
rect 50500 -11890 50560 0
rect 50600 -11890 50660 0
rect 50700 -11890 50760 0
rect 50800 -11890 50860 0
rect 50900 -11890 50960 0
rect 51000 -11890 51060 0
rect 51100 -11890 51160 0
rect 51200 -11890 51260 0
rect 51300 -11890 51360 0
rect 51400 -11890 51460 0
rect 51500 -11890 51560 0
rect 51600 -11890 51660 0
rect 51700 -11890 51760 0
rect 51800 -11890 51860 0
rect 51900 -11890 51960 0
rect 52000 -11890 52060 0
rect 52100 -11890 52160 0
rect 52200 -11890 52260 0
rect 52300 -11890 52360 0
rect 52400 -11890 52460 0
rect 52500 -11890 52560 0
rect 52600 -11890 52660 0
rect 52700 -11890 52760 0
rect 52800 -11890 52860 0
rect 52900 -11890 52960 0
rect 53000 -11890 53060 0
rect 48400 -17030 48460 -12610
rect 49100 -12670 49160 -12530
rect 48500 -17030 48560 -12740
rect 49200 -12810 49260 -12520
rect 48600 -17030 48660 -12880
rect 49300 -12950 49360 -12520
rect 48700 -17030 48760 -13010
rect 49400 -13080 49460 -12530
rect 48800 -17030 48860 -13150
rect 48900 -17020 48960 -13210
rect 48400 -18020 48460 -17670
rect 48500 -18040 48560 -17660
rect 48600 -18080 48660 -17660
rect 48700 -18120 48760 -17660
rect 34800 -29200 34860 -24480
rect 35100 -24510 35160 -24150
rect 35500 -24200 35560 -22300
rect 34600 -31910 34660 -29240
rect 34900 -29340 34960 -24580
rect 35200 -24590 35260 -24200
rect 35600 -24260 35660 -22450
rect 36700 -22460 36760 -22400
rect 36800 -22490 36860 -22200
rect 34700 -31870 34760 -29340
rect 35000 -29450 35060 -24680
rect 35300 -24690 35360 -24270
rect 34800 -31820 34860 -29480
rect 34900 -31770 34960 -29620
rect 35100 -29630 35160 -24780
rect 35400 -24790 35460 -24340
rect 35700 -24350 35760 -22510
rect 35800 -24400 35860 -22560
rect 35200 -29730 35260 -24880
rect 35500 -24890 35560 -24410
rect 35000 -31720 35060 -29750
rect 35100 -31670 35160 -29860
rect 35300 -29910 35360 -24970
rect 35600 -24990 35660 -24490
rect 35900 -24500 35960 -22590
rect 35700 -25050 35760 -24550
rect 36000 -24560 36060 -22620
rect 36100 -24620 36160 -22620
rect 36200 -24480 36260 -22670
rect 36300 -24160 36360 -22720
rect 36400 -23590 36460 -22750
rect 36500 -23010 36560 -22780
rect 36900 -23030 36960 -22060
rect 35400 -30100 35460 -25120
rect 35800 -25200 35860 -24630
rect 36200 -24640 36260 -24580
rect 35200 -31620 35260 -30100
rect 35300 -31570 35360 -30240
rect 35500 -30300 35560 -25220
rect 35900 -25290 35960 -24710
rect 35600 -30430 35660 -25320
rect 36000 -25390 36060 -24770
rect 36400 -24860 36460 -24300
rect 35400 -31530 35460 -30430
rect 35500 -31490 35560 -30580
rect 35700 -30620 35760 -25420
rect 36100 -25540 36160 -24860
rect 35600 -31480 35660 -30760
rect 35800 -30810 35860 -25560
rect 35700 -31480 35760 -30940
rect 35900 -30950 35960 -25660
rect 36200 -25680 36260 -24920
rect 36500 -24930 36560 -23890
rect 36300 -25780 36360 -25010
rect 36600 -25020 36660 -23290
rect 37000 -23340 37060 -21960
rect 35800 -31480 35860 -31090
rect 36000 -31140 36060 -25810
rect 36100 -31250 36160 -25910
rect 36400 -25970 36460 -25070
rect 36700 -25090 36760 -23360
rect 37100 -24100 37160 -21840
rect 37200 -22640 37260 -21840
rect 37300 -22650 37360 -21830
rect 37400 -22690 37460 -21790
rect 37500 -22730 37560 -21790
rect 37600 -22730 37660 -21750
rect 37700 -22770 37760 -21750
rect 37800 -22790 37860 -21710
rect 37900 -22810 37960 -21700
rect 38000 -22850 38060 -21660
rect 36800 -25090 36860 -24290
rect 37200 -24500 37260 -22850
rect 38100 -22860 38160 -21650
rect 36200 -31100 36260 -26050
rect 36500 -26110 36560 -25170
rect 36300 -30910 36360 -26150
rect 36600 -26250 36660 -25230
rect 36400 -30720 36460 -26290
rect 36700 -26440 36760 -25330
rect 36500 -30540 36560 -26440
rect 36800 -26550 36860 -25410
rect 36600 -29870 36660 -26620
rect 36700 -29250 36760 -26810
rect 36800 -28540 36860 -26990
rect 37100 -27010 37160 -26690
rect 37100 -27360 37160 -27300
rect 36600 -30940 36660 -30790
rect 36700 -30870 36760 -30530
rect 36800 -30800 36860 -30170
rect 36900 -30750 36960 -29500
rect 37000 -30700 37060 -28270
rect 37100 -30650 37160 -27710
rect 37200 -30600 37260 -25940
rect 37300 -30550 37360 -22880
rect 37400 -30500 37460 -22880
rect 38200 -22890 38260 -21620
rect 38300 -22900 38360 -21580
rect 38400 -22900 38460 -21580
rect 38500 -22920 38560 -21540
rect 37500 -30450 37560 -22930
rect 37600 -30380 37660 -22930
rect 38600 -22950 38660 -21530
rect 38700 -22950 38760 -21490
rect 38800 -22960 38860 -21480
rect 37700 -30330 37760 -22960
rect 38900 -22990 38960 -21450
rect 37800 -30260 37860 -22990
rect 37900 -30180 37960 -23010
rect 39000 -23020 39060 -21410
rect 38000 -30120 38060 -23020
rect 38100 -30040 38160 -23050
rect 38200 -29970 38260 -23060
rect 39100 -23080 39160 -21400
rect 38300 -29920 38360 -23100
rect 38400 -29870 38460 -23100
rect 38500 -29820 38560 -23100
rect 38600 -29780 38660 -23140
rect 38700 -29740 38760 -23140
rect 38800 -29690 38860 -23140
rect 38900 -29580 38960 -23190
rect 39200 -23270 39260 -21380
rect 39000 -29390 39060 -23320
rect 39300 -23420 39360 -21350
rect 39100 -29200 39160 -23420
rect 39400 -23560 39460 -21320
rect 39200 -28970 39260 -23560
rect 39500 -23600 39560 -21280
rect 39600 -23640 39660 -21240
rect 39700 -23690 39760 -21200
rect 39300 -23770 39360 -23700
rect 39800 -23730 39860 -21410
rect 39900 -23150 39960 -22100
rect 42500 -22670 42560 -22560
rect 39900 -23700 39960 -23210
rect 39300 -28610 39360 -24090
rect 39500 -24150 39560 -23880
rect 39400 -28250 39460 -24330
rect 39600 -24380 39660 -23850
rect 39500 -27800 39560 -24550
rect 39700 -24640 39760 -23900
rect 40100 -23940 40160 -23780
rect 39600 -27080 39660 -24870
rect 39800 -25050 39860 -23950
rect 39600 -27200 39660 -27140
rect 39200 -29460 39260 -29340
rect 39300 -29420 39360 -29150
rect 39400 -29370 39460 -28910
rect 39500 -29340 39560 -28430
rect 39600 -29300 39660 -28020
rect 39700 -29290 39760 -27530
rect 39800 -29260 39860 -26090
rect 39900 -29290 39960 -24000
rect 40200 -24020 40260 -23680
rect 40300 -24030 40360 -23630
rect 40400 -24040 40460 -23480
rect 40000 -29370 40060 -24090
rect 40100 -29260 40160 -24160
rect 40200 -29190 40260 -24250
rect 40500 -24310 40560 -23380
rect 40300 -28740 40360 -24330
rect 40600 -24410 40660 -23280
rect 40400 -28470 40460 -24450
rect 40700 -24510 40760 -23140
rect 40500 -28200 40560 -24560
rect 40600 -27750 40660 -24650
rect 40800 -24660 40860 -23050
rect 40900 -24800 40960 -22900
rect 40700 -27380 40760 -24800
rect 41000 -24900 41060 -22770
rect 40800 -26940 40860 -24900
rect 40900 -26540 40960 -25040
rect 41100 -25050 41160 -22800
rect 41000 -26080 41060 -25180
rect 41200 -25190 41260 -22990
rect 41300 -25330 41360 -23180
rect 41100 -25950 41160 -25330
rect 40800 -27730 40860 -27610
rect 40600 -27870 40660 -27810
rect 35900 -31470 35960 -31280
rect 31700 -34450 31760 -34340
rect 31800 -34390 31860 -34200
rect 31900 -34300 31960 -34110
rect 32000 -34240 32060 -34000
rect 32100 -34140 32160 -33910
rect 32200 -34090 32260 -33810
rect 32300 -34030 32360 -33710
rect 32400 -33930 32460 -33610
rect 32500 -33880 32560 -33510
rect 32600 -33780 32660 -33450
rect 32700 -33720 32760 -33350
rect 32800 -33660 32860 -33250
rect 32900 -33600 32960 -33190
rect 33000 -33520 33060 -33120
rect 33100 -33450 33160 -33040
rect 33200 -33400 33260 -32970
rect 33300 -33340 33360 -32900
rect 33400 -33280 33460 -32830
rect 33500 -33210 33560 -32770
rect 33600 -33160 33660 -32710
rect 33700 -33080 33760 -32640
rect 33800 -33040 33860 -32560
rect 33900 -32990 33960 -32510
rect 34000 -32940 34060 -32440
rect 34100 -32880 34160 -32390
rect 34200 -32830 34260 -32340
rect 34300 -32780 34360 -32280
rect 34400 -32740 34460 -32220
rect 34500 -32710 34560 -32170
rect 34600 -32650 34660 -32120
rect 34700 -32610 34760 -32070
rect 34800 -32560 34860 -32020
rect 34900 -32510 34960 -31980
rect 35000 -32460 35060 -31920
rect 35100 -32390 35160 -31870
rect 31300 -42200 31360 -34850
rect 31400 -38500 31460 -34850
rect 31500 -38310 31560 -34800
rect 31600 -38040 31660 -34730
rect 31700 -37770 31760 -34660
rect 31800 -37400 31860 -34600
rect 31900 -37170 31960 -34510
rect 32000 -36940 32060 -34440
rect 32100 -36630 32160 -34380
rect 32200 -36400 32260 -34290
rect 32300 -36160 32360 -34220
rect 32400 -35940 32460 -34160
rect 32500 -35710 32560 -34080
rect 32600 -35520 32660 -34020
rect 32700 -35330 32760 -33940
rect 32800 -35140 32860 -33860
rect 32900 -34960 32960 -33810
rect 33000 -34810 33060 -33750
rect 33100 -34660 33160 -33680
rect 33200 -34530 33260 -33600
rect 33300 -34380 33360 -33540
rect 33400 -34240 33460 -33480
rect 33500 -34100 33560 -33420
rect 33600 -34000 33660 -33360
rect 33700 -33850 33760 -33310
rect 33800 -33750 33860 -33240
rect 33900 -33650 33960 -33190
rect 34000 -33510 34060 -33140
rect 34100 -33410 34160 -33090
rect 34200 -33310 34260 -33040
rect 34300 -33160 34360 -32980
rect 34400 -33060 34460 -32940
rect 34500 -33020 34560 -32960
rect 31800 -37520 31860 -37460
rect 31400 -42120 31460 -38560
rect 31500 -42050 31560 -38630
rect 31600 -41960 31660 -38490
rect 31700 -41880 31760 -38220
rect 31800 -41810 31860 -37950
rect 31900 -41730 31960 -37630
rect 32000 -41650 32060 -37310
rect 32100 -41570 32160 -37080
rect 32200 -41490 32260 -36850
rect 32300 -41410 32360 -36580
rect 32400 -41320 32460 -36300
rect 32500 -41370 32560 -36120
rect 32600 -41520 32660 -35890
rect 32700 -41660 32760 -35660
rect 32800 -41830 32860 -35470
rect 32900 -41990 32960 -35280
rect 33000 -42140 33060 -35090
rect 33100 -42290 33160 -34950
rect 33200 -42420 33260 -34810
rect 29500 -45320 29560 -45250
rect 26300 -48580 26360 -45890
rect 26400 -48580 26460 -46030
rect 26500 -48580 26560 -46070
rect 26600 -48580 26660 -45990
rect 26700 -46020 26760 -45940
rect 26800 -45970 26860 -45900
rect 26700 -48580 26760 -46250
rect 26800 -48580 26860 -46220
rect 26900 -46280 26960 -46220
rect 26900 -48580 26960 -46400
rect 27000 -48580 27060 -46430
rect 27100 -48580 27160 -46390
rect 27200 -46520 27260 -46390
rect 27200 -48580 27260 -46710
rect 27300 -48580 27360 -46710
rect 27400 -48580 27460 -46660
rect 27500 -48580 27560 -46600
rect 27600 -48580 27660 -46540
rect 27700 -48580 27760 -46470
rect 27800 -48580 27860 -46390
rect 27900 -48580 27960 -46330
rect 28000 -48580 28060 -46270
rect 28100 -48580 28160 -46180
rect 28200 -48580 28260 -46110
rect 28300 -48580 28360 -46060
rect 28400 -48580 28460 -45960
rect 28500 -48580 28560 -45900
rect 28600 -48580 28660 -45820
rect 28700 -48580 28760 -45750
rect 28800 -48580 28860 -45690
rect 28900 -48580 28960 -45640
rect 29000 -48580 29060 -45630
rect 29100 -48580 29160 -45560
rect 29200 -48580 29260 -45490
rect 29300 -48580 29360 -45440
rect 29400 -48580 29460 -45530
rect 29500 -48580 29560 -45770
rect 29600 -48580 29660 -45190
rect 29700 -48580 29760 -45090
rect 29800 -48580 29860 -44980
rect 29900 -48580 29960 -44910
rect 30000 -48580 30060 -44860
rect 30100 -48580 30160 -44800
rect 30200 -48580 30260 -44730
rect 30300 -48580 30360 -44670
rect 30400 -48580 30460 -44600
rect 30500 -48580 30560 -44540
rect 30600 -48580 30660 -44470
rect 30700 -48580 30760 -44390
rect 30800 -48580 30860 -44320
rect 30900 -48580 30960 -44250
rect 31000 -48580 31060 -44170
rect 31100 -48580 31160 -44100
rect 31200 -48580 31260 -44030
rect 31300 -48580 31360 -43960
rect 31400 -48580 31460 -43900
rect 31500 -48580 31560 -43830
rect 31600 -48580 31660 -43770
rect 31700 -48580 31760 -43690
rect 31800 -48580 31860 -43620
rect 31900 -48580 31960 -43540
rect 32000 -48580 32060 -43460
rect 32100 -48580 32160 -43390
rect 32200 -48580 32260 -43310
rect 32300 -48580 32360 -43240
rect 32400 -48580 32460 -43150
rect 32500 -48580 32560 -43080
rect 32600 -48580 32660 -43000
rect 32700 -48580 32760 -42920
rect 32800 -48580 32860 -42850
rect 32900 -48580 32960 -42760
rect 33000 -48580 33060 -42680
rect 33100 -48580 33160 -42600
rect 33200 -48580 33260 -42520
rect 33300 -48580 33360 -34670
rect 33400 -48580 33460 -34520
rect 33500 -48580 33560 -34380
rect 33600 -48580 33660 -34280
rect 33700 -48580 33760 -34130
rect 33800 -48580 33860 -33990
rect 33900 -48580 33960 -33890
rect 34000 -48580 34060 -33750
rect 34100 -48580 34160 -33650
rect 34200 -39810 34260 -33550
rect 34300 -39730 34360 -33450
rect 34400 -39630 34460 -33310
rect 34500 -39540 34560 -33200
rect 34600 -39450 34660 -33110
rect 34700 -39380 34760 -33010
rect 34800 -39280 34860 -32860
rect 34900 -39200 34960 -32760
rect 35000 -39100 35060 -32680
rect 35100 -39020 35160 -32610
rect 35200 -38920 35260 -31820
rect 35300 -38840 35360 -31770
rect 35400 -38740 35460 -31750
rect 35500 -38660 35560 -31690
rect 35600 -38560 35660 -31670
rect 35700 -38400 35760 -31690
rect 35800 -38350 35860 -31790
rect 35900 -38280 35960 -31770
rect 36000 -38200 36060 -31630
rect 36100 -38100 36160 -31610
rect 36200 -38000 36260 -31460
rect 36300 -37880 36360 -31380
rect 36400 -37770 36460 -31310
rect 36500 -37670 36560 -31240
rect 36600 -37570 36660 -31150
rect 36700 -37530 36760 -31090
rect 36800 -37410 36860 -31020
rect 36900 -37230 36960 -30940
rect 37000 -37170 37060 -30900
rect 37100 -37100 37160 -30850
rect 37200 -37010 37260 -30800
rect 37300 -36880 37360 -30750
rect 37400 -36750 37460 -30700
rect 37500 -36670 37560 -30650
rect 37600 -36570 37660 -30590
rect 37700 -36520 37760 -30540
rect 37800 -36460 37860 -30480
rect 37900 -36360 37960 -30410
rect 38000 -36260 38060 -30320
rect 38100 -36170 38160 -30270
rect 38200 -36060 38260 -30190
rect 38300 -35970 38360 -30120
rect 38400 -35870 38460 -30070
rect 38500 -35760 38560 -30020
rect 38600 -35660 38660 -29980
rect 38700 -35560 38760 -29940
rect 38800 -35470 38860 -29890
rect 38900 -35350 38960 -29840
rect 39000 -35240 39060 -29800
rect 39100 -35140 39160 -29750
rect 39200 -31670 39260 -29690
rect 39300 -30220 39360 -29620
rect 39400 -30040 39460 -29580
rect 39400 -30550 39460 -30490
rect 39400 -30670 39460 -30610
rect 39200 -35020 39260 -33260
rect 39300 -34920 39360 -32630
rect 39400 -34830 39460 -30970
rect 39500 -34730 39560 -29540
rect 39600 -34630 39660 -29500
rect 39700 -34530 39760 -29460
rect 39800 -34420 39860 -29450
rect 39900 -34300 39960 -29430
rect 40000 -34210 40060 -29500
rect 40200 -29590 40260 -29390
rect 40100 -34090 40160 -29770
rect 40300 -29860 40360 -29330
rect 40200 -33980 40260 -30040
rect 40400 -30090 40460 -29010
rect 40500 -30150 40560 -28650
rect 40600 -30200 40660 -28380
rect 40700 -28950 40760 -28060
rect 40800 -28910 40860 -27790
rect 40900 -28840 40960 -27160
rect 41000 -28820 41060 -26760
rect 41100 -28780 41160 -26400
rect 41200 -28780 41260 -25470
rect 41400 -25480 41460 -23280
rect 41500 -25620 41560 -23420
rect 41300 -28740 41360 -25620
rect 41600 -25760 41660 -23520
rect 41400 -28730 41460 -25760
rect 41700 -25860 41760 -23660
rect 41500 -28730 41560 -25860
rect 41800 -26000 41860 -23760
rect 41600 -28690 41660 -26000
rect 41900 -26100 41960 -23880
rect 41700 -28690 41760 -26140
rect 42000 -26200 42060 -23760
rect 41800 -28690 41860 -26250
rect 42100 -26300 42160 -23610
rect 41900 -28670 41960 -26340
rect 42200 -26400 42260 -23420
rect 42000 -28690 42060 -26450
rect 42100 -28690 42160 -26540
rect 42300 -26550 42360 -23200
rect 42200 -28730 42260 -26680
rect 42400 -26690 42460 -22970
rect 42500 -26880 42560 -22730
rect 42300 -28740 42360 -26880
rect 42600 -27020 42660 -22340
rect 40800 -30220 40860 -29220
rect 40900 -30280 40960 -29170
rect 40300 -33880 40360 -30320
rect 40400 -33760 40460 -30590
rect 40900 -30810 40960 -30460
rect 40500 -33670 40560 -30910
rect 40600 -31040 40660 -30970
rect 40600 -33550 40660 -31100
rect 40700 -33450 40760 -31410
rect 40800 -33330 40860 -31730
rect 41000 -32000 41060 -29020
rect 40900 -32510 40960 -32310
rect 41100 -32570 41160 -28970
rect 40900 -33220 40960 -32570
rect 41100 -32800 41160 -32740
rect 41200 -32850 41260 -28970
rect 41300 -32780 41360 -28930
rect 41400 -32670 41460 -28930
rect 41500 -32740 41560 -28910
rect 41600 -32850 41660 -28890
rect 41700 -32970 41760 -28890
rect 41000 -33110 41060 -33020
rect 41800 -33100 41860 -28890
rect 41900 -33240 41960 -28850
rect 42000 -33380 42060 -28850
rect 42100 -33510 42160 -28890
rect 42400 -28910 42460 -27020
rect 42200 -33640 42260 -28910
rect 42200 -33960 42260 -33790
rect 42300 -33930 42360 -28930
rect 42400 -33840 42460 -28970
rect 34200 -48580 34260 -39900
rect 34300 -48580 34360 -40040
rect 34400 -48580 34460 -40180
rect 34500 -48580 34560 -40310
rect 34600 -48580 34660 -40460
rect 34700 -48580 34760 -40590
rect 34800 -48580 34860 -40730
rect 35400 -40740 35460 -40680
rect 34900 -48580 34960 -40860
rect 35000 -48580 35060 -40980
rect 35100 -48580 35160 -40920
rect 35200 -48580 35260 -40830
rect 35300 -48580 35360 -40740
rect 35400 -48580 35460 -40840
rect 35500 -48580 35560 -40740
rect 35600 -48580 35660 -40720
rect 35700 -48580 35760 -40670
rect 35800 -48580 35860 -40570
rect 35900 -48580 35960 -40470
rect 36000 -48580 36060 -40370
rect 36100 -48580 36160 -40270
rect 36200 -48580 36260 -40170
rect 36300 -48580 36360 -40070
rect 36400 -48580 36460 -39970
rect 36500 -48580 36560 -39900
rect 36600 -48580 36660 -39810
rect 36700 -48580 36760 -39710
rect 36800 -48580 36860 -39640
rect 36900 -48580 36960 -39560
rect 37000 -48580 37060 -39470
rect 37100 -48580 37160 -39400
rect 37200 -48580 37260 -39300
rect 37300 -48580 37360 -39200
rect 37400 -48580 37460 -39100
rect 37500 -48580 37560 -39000
rect 37600 -48580 37660 -38900
rect 37700 -48580 37760 -38800
rect 37800 -48580 37860 -38750
rect 37900 -48580 37960 -38640
rect 38000 -48580 38060 -38550
rect 38100 -48580 38160 -38470
rect 38200 -48580 38260 -38390
rect 38300 -48580 38360 -38290
rect 38400 -48580 38460 -38190
rect 38500 -48580 38560 -38090
rect 38600 -48580 38660 -37990
rect 38700 -48580 38760 -37890
rect 38800 -48580 38860 -37790
rect 38900 -48580 38960 -37650
rect 39000 -48580 39060 -37590
rect 39100 -48580 39160 -37470
rect 39200 -48580 39260 -37350
rect 39300 -48580 39360 -37250
rect 39400 -48580 39460 -37150
rect 39500 -48580 39560 -37050
rect 39600 -48580 39660 -36950
rect 39700 -48580 39760 -36850
rect 39800 -48580 39860 -36710
rect 39900 -48580 39960 -36610
rect 40000 -48580 40060 -36500
rect 40100 -48580 40160 -36400
rect 40200 -48580 40260 -36300
rect 40300 -48580 40360 -36210
rect 40400 -48580 40460 -36150
rect 40500 -48580 40560 -36050
rect 40600 -48580 40660 -35950
rect 40700 -48580 40760 -35850
rect 40800 -48580 40860 -35750
rect 40900 -48580 40960 -35610
rect 41000 -48580 41060 -35510
rect 41100 -48580 41160 -35410
rect 41200 -48580 41260 -35260
rect 41300 -48580 41360 -35170
rect 41400 -48580 41460 -35160
rect 41600 -35250 41660 -34860
rect 41500 -48580 41560 -35510
rect 41700 -35700 41760 -34770
rect 41600 -35980 41660 -35920
rect 41600 -48580 41660 -36040
rect 41800 -36100 41860 -34700
rect 41800 -36220 41860 -36160
rect 41800 -36370 41860 -36280
rect 41900 -36770 41960 -34610
rect 42000 -36710 42060 -34510
rect 41700 -48580 41760 -36810
rect 41800 -48580 41860 -36860
rect 41900 -48580 41960 -36910
rect 42100 -37100 42160 -34410
rect 42000 -48580 42060 -37460
rect 42200 -37680 42260 -34310
rect 42100 -48580 42160 -37950
rect 42300 -38210 42360 -34160
rect 42200 -48580 42260 -38520
rect 42400 -38880 42460 -34020
rect 42300 -39300 42360 -39240
rect 42300 -39460 42360 -39380
rect 42300 -48580 42360 -39520
rect 42500 -39620 42560 -27160
rect 42700 -27170 42760 -22160
rect 42500 -39740 42560 -39680
rect 42500 -39930 42560 -39800
rect 42400 -48580 42460 -40290
rect 42600 -40640 42660 -27300
rect 42800 -27350 42860 -22090
rect 42500 -48580 42560 -40960
rect 42700 -41220 42760 -27490
rect 42900 -27540 42960 -22020
rect 42800 -31030 42860 -27680
rect 43000 -27730 43060 -21970
rect 43100 -27860 43160 -21910
rect 42900 -30920 42960 -27860
rect 43200 -28050 43260 -21850
rect 43000 -30790 43060 -28050
rect 43100 -30660 43160 -28190
rect 43300 -28240 43360 -21790
rect 43200 -30550 43260 -28380
rect 43400 -28390 43460 -21730
rect 43300 -30430 43360 -28520
rect 43500 -28530 43560 -21670
rect 43500 -28650 43560 -28590
rect 43400 -30300 43460 -28760
rect 43600 -28810 43660 -21620
rect 43500 -30180 43560 -28930
rect 43600 -29230 43660 -28910
rect 43700 -29160 43760 -21560
rect 43600 -30070 43660 -29300
rect 43800 -29350 43860 -21500
rect 43700 -29950 43760 -29490
rect 43900 -29530 43960 -21450
rect 44000 -29530 44060 -21390
rect 44100 -29440 44160 -21340
rect 44200 -29310 44260 -21280
rect 44300 -29180 44360 -21230
rect 44400 -29040 44460 -21180
rect 44500 -28910 44560 -21120
rect 44600 -28790 44660 -21080
rect 44700 -28660 44760 -21020
rect 44800 -28520 44860 -20970
rect 44900 -28380 44960 -20920
rect 45000 -28260 45060 -20870
rect 45100 -28120 45160 -20830
rect 45200 -27980 45260 -20790
rect 45300 -27840 45360 -20740
rect 45400 -27710 45460 -20690
rect 45500 -27580 45560 -20640
rect 45600 -27440 45660 -20600
rect 45700 -27290 45760 -20570
rect 45800 -27150 45860 -20520
rect 45900 -27000 45960 -20480
rect 46000 -26860 46060 -20440
rect 46100 -26720 46160 -20400
rect 46200 -26580 46260 -20360
rect 46300 -26410 46360 -20320
rect 46400 -26270 46460 -20280
rect 46500 -26120 46560 -20250
rect 46600 -25970 46660 -20220
rect 46700 -25810 46760 -20190
rect 46800 -25660 46860 -20160
rect 46900 -25510 46960 -20130
rect 47000 -25350 47060 -20090
rect 47100 -25170 47160 -20070
rect 47200 -25010 47260 -20050
rect 47300 -24860 47360 -20030
rect 47400 -24720 47460 -20010
rect 47500 -24840 47560 -18160
rect 48800 -18170 48860 -17660
rect 48900 -18230 48960 -17660
rect 47600 -25000 47660 -18300
rect 49000 -18310 49060 -13210
rect 49100 -18410 49160 -13200
rect 47700 -25120 47760 -18430
rect 49200 -18530 49260 -13210
rect 47800 -25290 47860 -18590
rect 49300 -18620 49360 -13210
rect 47900 -25400 47960 -18720
rect 49400 -18870 49460 -13210
rect 48000 -25530 48060 -18890
rect 49500 -19030 49560 -12530
rect 48100 -25770 48160 -19040
rect 48200 -23250 48260 -19190
rect 49600 -19210 49660 -12530
rect 48300 -23060 48360 -19320
rect 49600 -19330 49660 -19270
rect 48400 -20660 48460 -19450
rect 49700 -19530 49760 -12530
rect 49800 -17020 49860 -12530
rect 49900 -17030 49960 -12530
rect 50000 -17030 50060 -12530
rect 50100 -17030 50160 -12530
rect 50200 -17030 50260 -12520
rect 50300 -17030 50360 -12520
rect 50400 -17030 50460 -12520
rect 50500 -17030 50560 -12520
rect 50600 -17030 50660 -12520
rect 50700 -17030 50760 -12520
rect 50800 -17030 50860 -12520
rect 50900 -17030 50960 -12520
rect 51000 -14240 51060 -12520
rect 51100 -14240 51160 -12520
rect 51200 -14240 51260 -12520
rect 51300 -14240 51360 -12520
rect 51400 -14240 51460 -12520
rect 51500 -14240 51560 -12520
rect 51000 -17030 51060 -16210
rect 51100 -17030 51160 -16210
rect 51200 -17030 51260 -16210
rect 51300 -17030 51360 -16210
rect 51400 -17030 51460 -16210
rect 51500 -17030 51560 -16210
rect 51600 -17030 51660 -12520
rect 51700 -17030 51760 -12520
rect 51800 -17030 51860 -12520
rect 51900 -17030 51960 -12520
rect 52000 -17030 52060 -12520
rect 52100 -17030 52160 -12520
rect 52200 -17030 52260 -12520
rect 52300 -17030 52360 -12520
rect 52400 -17030 52460 -12520
rect 52500 -17030 52560 -12520
rect 52600 -17030 52660 -12520
rect 52700 -17030 52760 -12520
rect 52800 -17030 52860 -12520
rect 52900 -17030 52960 -12530
rect 53000 -17030 53060 -12530
rect 48500 -20660 48560 -19580
rect 48600 -20660 48660 -19710
rect 48700 -20660 48760 -19850
rect 49800 -19890 49860 -17670
rect 49900 -19100 49960 -17660
rect 50000 -18960 50060 -17660
rect 50100 -18880 50160 -17660
rect 50200 -18810 50260 -17660
rect 50300 -18750 50360 -17660
rect 50400 -18710 50460 -17660
rect 50500 -18680 50560 -17660
rect 50600 -18660 50660 -17660
rect 50700 -18640 50760 -17660
rect 50800 -18640 50860 -17660
rect 50900 -18640 50960 -17660
rect 51000 -18640 51060 -17660
rect 51100 -18640 51160 -17660
rect 51200 -18640 51260 -17660
rect 51300 -18640 51360 -17660
rect 51400 -18640 51460 -17660
rect 51500 -18640 51560 -17660
rect 51600 -18640 51660 -17660
rect 51700 -18640 51760 -17660
rect 51800 -18640 51860 -17660
rect 51900 -18640 51960 -17660
rect 52000 -18640 52060 -17660
rect 52100 -18640 52160 -17660
rect 52200 -18640 52260 -17660
rect 52300 -18640 52360 -17660
rect 52400 -18640 52460 -17660
rect 52500 -18640 52560 -17660
rect 52600 -18640 52660 -17660
rect 52700 -18640 52760 -17660
rect 52800 -18640 52860 -17660
rect 52900 -18640 52960 -17660
rect 53000 -18640 53060 -17670
rect 48800 -20650 48860 -19990
rect 48900 -20680 48960 -20030
rect 48900 -20800 48960 -20740
rect 48400 -22850 48460 -21310
rect 48500 -22630 48560 -21310
rect 48600 -22410 48660 -21310
rect 48700 -22190 48760 -21310
rect 48800 -21950 48860 -21230
rect 48900 -21680 48960 -20860
rect 49000 -21400 49060 -20070
rect 49100 -21090 49160 -20120
rect 49200 -20760 49260 -20190
rect 49300 -20330 49360 -20270
rect 49900 -20380 49960 -19280
rect 43800 -29820 43860 -29680
rect 44800 -31130 44860 -30840
rect 42600 -48580 42660 -41490
rect 42800 -41850 42860 -31300
rect 42800 -41980 42860 -41920
rect 42700 -48580 42760 -42550
rect 42900 -43040 42960 -31430
rect 42800 -48580 42860 -43560
rect 43000 -44100 43060 -31580
rect 42900 -48580 42960 -44490
rect 43100 -44970 43160 -31700
rect 43000 -48580 43060 -46210
rect 43200 -47480 43260 -31840
rect 43100 -48580 43160 -47550
rect 43200 -48580 43260 -47540
rect 43300 -48580 43360 -31960
rect 43400 -48580 43460 -32110
rect 43500 -48580 43560 -32230
rect 43600 -48580 43660 -32340
rect 43700 -48580 43760 -32330
rect 43800 -48580 43860 -32160
rect 43900 -48580 43960 -32030
rect 44000 -48580 44060 -31900
rect 44100 -48580 44160 -31770
rect 44200 -48580 44260 -31630
rect 44300 -48580 44360 -31500
rect 44400 -48580 44460 -31370
rect 44500 -48580 44560 -31240
rect 44600 -48580 44660 -31160
rect 44700 -48580 44760 -31270
rect 44900 -31320 44960 -30710
rect 44800 -48580 44860 -31460
rect 45000 -31510 45060 -30580
rect 44900 -48580 44960 -31640
rect 45100 -31740 45160 -30440
rect 45000 -48580 45060 -31880
rect 45200 -31890 45260 -30280
rect 45100 -48580 45160 -32060
rect 45300 -32110 45360 -30140
rect 45200 -48580 45260 -32250
rect 45400 -32330 45460 -30020
rect 45500 -32360 45560 -29880
rect 45300 -48580 45360 -32530
rect 45400 -48580 45460 -32670
rect 45600 -32720 45660 -29740
rect 45500 -48580 45560 -32850
rect 45700 -32860 45760 -29600
rect 45800 -33000 45860 -29480
rect 45600 -48580 45660 -33000
rect 45700 -48580 45760 -33140
rect 45900 -33190 45960 -29350
rect 45800 -48580 45860 -33370
rect 46000 -33380 46060 -29200
rect 45900 -48580 45960 -33510
rect 46100 -33560 46160 -29060
rect 46000 -48580 46060 -33700
rect 46200 -33750 46260 -28920
rect 46100 -48580 46160 -33930
rect 46300 -33990 46360 -28800
rect 46200 -48580 46260 -34120
rect 46400 -34170 46460 -28640
rect 46300 -48580 46360 -34310
rect 46500 -34350 46560 -28510
rect 46400 -48580 46460 -34540
rect 46600 -34630 46660 -28360
rect 46500 -48580 46560 -34760
rect 46700 -34820 46760 -28210
rect 46600 -48580 46660 -34990
rect 46800 -35040 46860 -28070
rect 46700 -48580 46760 -35180
rect 46900 -35320 46960 -27920
rect 46800 -48580 46860 -35460
rect 47000 -35510 47060 -27780
rect 46900 -48580 46960 -35690
rect 47100 -35740 47160 -27620
rect 47000 -48580 47060 -35880
rect 47200 -35960 47260 -27480
rect 47100 -48580 47160 -36190
rect 47300 -36290 47360 -27320
rect 47200 -48580 47260 -36420
rect 47400 -36520 47460 -27160
rect 47300 -48580 47360 -36650
rect 47500 -36700 47560 -27000
rect 47400 -48580 47460 -36890
rect 47600 -36940 47660 -26850
rect 47600 -37060 47660 -37000
rect 47500 -48580 47560 -37160
rect 47700 -37250 47760 -26700
rect 47600 -48580 47660 -37390
rect 47800 -37480 47860 -26530
rect 47700 -48580 47760 -37660
rect 47900 -37750 47960 -26360
rect 47800 -48580 47860 -38020
rect 48000 -38210 48060 -26190
rect 47900 -48580 47960 -38430
rect 48100 -38610 48160 -26030
rect 48000 -48580 48060 -38780
rect 48200 -38970 48260 -23340
rect 48100 -39220 48160 -39160
rect 48100 -48580 48160 -39280
rect 48300 -39420 48360 -23510
rect 48400 -30760 48460 -23670
rect 48500 -30760 48560 -23830
rect 48600 -30750 48660 -24010
rect 48700 -30760 48760 -24150
rect 48800 -30760 48860 -24310
rect 48900 -30760 48960 -24460
rect 49000 -30760 49060 -24310
rect 49100 -30760 49160 -24100
rect 49200 -30760 49260 -23850
rect 49300 -30760 49360 -23600
rect 49400 -30760 49460 -23330
rect 49500 -30760 49560 -23140
rect 49600 -30760 49660 -22910
rect 49700 -23370 49760 -22680
rect 49800 -23080 49860 -22410
rect 49900 -22860 49960 -22140
rect 50000 -22670 50060 -19630
rect 50100 -19970 50160 -19910
rect 50100 -22490 50160 -20030
rect 50300 -20070 50360 -19860
rect 50400 -20350 50460 -19590
rect 50200 -22190 50260 -20440
rect 50500 -20460 50560 -19470
rect 50600 -20540 50660 -19400
rect 50700 -20590 50760 -19350
rect 50800 -20630 50860 -19310
rect 50900 -20640 50960 -19290
rect 51000 -20650 51060 -19280
rect 51100 -20660 51160 -19270
rect 51200 -20660 51260 -19270
rect 51300 -20660 51360 -19270
rect 51400 -20660 51460 -19270
rect 51500 -20660 51560 -19270
rect 51600 -20660 51660 -19270
rect 51700 -20660 51760 -19270
rect 51800 -20660 51860 -19270
rect 51900 -20660 51960 -19270
rect 52000 -20660 52060 -19270
rect 52100 -20660 52160 -19270
rect 52200 -20660 52260 -19270
rect 52300 -20660 52360 -19270
rect 52400 -20660 52460 -19270
rect 52500 -20660 52560 -19270
rect 52600 -20660 52660 -19270
rect 52700 -20660 52760 -19270
rect 52800 -20660 52860 -19270
rect 52900 -20660 52960 -19270
rect 53000 -20660 53060 -19270
rect 50300 -22250 50360 -21310
rect 50400 -22340 50460 -21310
rect 50500 -22430 50560 -21310
rect 49700 -26480 49760 -23600
rect 50300 -23700 50360 -23030
rect 50400 -23860 50460 -22750
rect 50500 -23940 50560 -22590
rect 50600 -23970 50660 -21310
rect 50700 -23990 50760 -21310
rect 50800 -23970 50860 -21310
rect 50900 -23900 50960 -21310
rect 51000 -23760 51060 -21310
rect 51100 -22900 51160 -21310
rect 51200 -22510 51260 -21310
rect 51300 -22330 51360 -21310
rect 51400 -22220 51460 -21310
rect 51500 -22150 51560 -21310
rect 51600 -22100 51660 -21310
rect 51700 -22060 51760 -21310
rect 51800 -22030 51860 -21310
rect 51900 -22020 51960 -21310
rect 52000 -22000 52060 -21310
rect 52100 -22000 52160 -21310
rect 52200 -22020 52260 -21310
rect 52300 -22030 52360 -21310
rect 52400 -22070 52460 -21310
rect 52500 -22110 52560 -21310
rect 52600 -22180 52660 -21310
rect 52700 -22270 52760 -21310
rect 52800 -22390 52860 -21310
rect 52900 -22550 52960 -21310
rect 49800 -26030 49860 -24020
rect 49900 -25830 49960 -24210
rect 50000 -25700 50060 -24340
rect 50100 -25600 50160 -24440
rect 50200 -25540 50260 -24510
rect 50300 -25500 50360 -24550
rect 50400 -25470 50460 -24590
rect 50500 -25430 50560 -24620
rect 50600 -25430 50660 -24620
rect 50700 -25420 50760 -24630
rect 50800 -25420 50860 -24620
rect 50900 -25420 50960 -24610
rect 51000 -25420 51060 -24580
rect 51100 -25420 51160 -24540
rect 51200 -25420 51260 -24480
rect 51300 -25420 51360 -24400
rect 51400 -25420 51460 -24280
rect 51500 -25420 51560 -24120
rect 51600 -25420 51660 -23800
rect 51700 -25420 51760 -22890
rect 51800 -25420 51860 -22730
rect 51900 -25420 51960 -22670
rect 52000 -25420 52060 -22660
rect 52100 -24380 52160 -22660
rect 52200 -24250 52260 -22680
rect 52300 -24120 52360 -22730
rect 53000 -22810 53060 -21310
rect 52400 -23920 52460 -22870
rect 52500 -23420 52560 -23250
rect 52100 -25420 52160 -24440
rect 52200 -25420 52260 -24520
rect 52300 -25420 52360 -24620
rect 52400 -25420 52460 -24720
rect 52500 -25420 52560 -24810
rect 52600 -25420 52660 -24720
rect 52700 -25420 52760 -24580
rect 52800 -25420 52860 -24430
rect 52900 -25420 52960 -24230
rect 53000 -25420 53060 -23950
rect 49700 -29690 49760 -27000
rect 50300 -27140 50360 -26390
rect 50400 -27320 50460 -26190
rect 49800 -29360 49860 -27450
rect 49900 -29190 49960 -27630
rect 50000 -29060 50060 -27770
rect 50100 -28970 50160 -27870
rect 50200 -28900 50260 -27820
rect 50300 -28850 50360 -27690
rect 50400 -28810 50460 -27560
rect 50500 -28780 50560 -26110
rect 50600 -28760 50660 -26070
rect 50700 -28740 50760 -26060
rect 50800 -28730 50860 -26060
rect 50900 -28730 50960 -26060
rect 51000 -28730 51060 -26060
rect 51100 -28730 51160 -26080
rect 51700 -27300 51760 -26060
rect 51800 -27420 51860 -26060
rect 51900 -27470 51960 -26060
rect 52000 -27480 52060 -26060
rect 52100 -27480 52160 -26070
rect 52200 -27460 52260 -26100
rect 52800 -26140 52860 -26060
rect 52300 -27400 52360 -26140
rect 52400 -27290 52460 -26220
rect 52900 -26230 52960 -26060
rect 53000 -26390 53060 -26060
rect 52500 -26980 52560 -26590
rect 51200 -28730 51260 -27500
rect 51300 -28730 51360 -27700
rect 51400 -28730 51460 -27820
rect 51500 -28730 51560 -27910
rect 51600 -28730 51660 -27980
rect 51700 -28730 51760 -28020
rect 51800 -28730 51860 -28060
rect 51900 -28730 51960 -28080
rect 52000 -28730 52060 -28100
rect 52100 -28730 52160 -28100
rect 52200 -28730 52260 -28090
rect 52300 -28730 52360 -28070
rect 52400 -28730 52460 -28050
rect 52500 -28730 52560 -28000
rect 52600 -28730 52660 -27940
rect 52700 -28730 52760 -27860
rect 52800 -28730 52860 -27770
rect 52900 -28730 52960 -27630
rect 53000 -28730 53060 -27420
rect 49700 -30760 49760 -29970
rect 50300 -30180 50360 -29970
rect 49800 -30760 49860 -30360
rect 50400 -30450 50460 -29690
rect 49900 -30760 49960 -30530
rect 50500 -30560 50560 -29570
rect 50000 -30750 50060 -30630
rect 50600 -30640 50660 -29490
rect 50700 -30690 50760 -29440
rect 50800 -30730 50860 -29410
rect 50900 -30740 50960 -29390
rect 51000 -30750 51060 -29370
rect 51100 -30760 51160 -29370
rect 51200 -30760 51260 -29370
rect 51300 -30760 51360 -29370
rect 51400 -30760 51460 -29370
rect 51500 -30760 51560 -29370
rect 51600 -30760 51660 -29370
rect 51700 -30760 51760 -29370
rect 51800 -30760 51860 -29370
rect 51900 -30760 51960 -29370
rect 52000 -30760 52060 -29370
rect 52100 -30760 52160 -29370
rect 52200 -30760 52260 -29370
rect 52300 -30760 52360 -29370
rect 52400 -30760 52460 -29370
rect 52500 -30760 52560 -29370
rect 52600 -30760 52660 -29370
rect 52700 -30760 52760 -29370
rect 52800 -30760 52860 -29370
rect 52900 -30750 52960 -29370
rect 53000 -30750 53060 -29370
rect 48200 -48580 48260 -39600
rect 48400 -39780 48460 -31410
rect 48300 -48580 48360 -39960
rect 48500 -40140 48560 -31410
rect 48400 -40440 48460 -40380
rect 48400 -48580 48460 -40500
rect 48600 -40580 48660 -31410
rect 48600 -40790 48660 -40640
rect 48500 -48580 48560 -41030
rect 48700 -41340 48760 -31410
rect 48800 -39380 48860 -31410
rect 48900 -39380 48960 -31410
rect 49000 -39380 49060 -31410
rect 49100 -39380 49160 -31410
rect 49200 -39380 49260 -31410
rect 49300 -39380 49360 -31410
rect 49400 -39380 49460 -31410
rect 49500 -39380 49560 -31410
rect 49600 -39380 49660 -31410
rect 49700 -36820 49760 -31410
rect 49800 -32340 49860 -31410
rect 49900 -32350 49960 -31410
rect 50000 -32350 50060 -31410
rect 50100 -32350 50160 -31410
rect 50200 -32350 50260 -31410
rect 50300 -32350 50360 -31410
rect 50400 -32350 50460 -31410
rect 50500 -32350 50560 -31410
rect 50600 -32350 50660 -31410
rect 50700 -32350 50760 -31410
rect 50800 -32350 50860 -31410
rect 50900 -32350 50960 -31410
rect 51000 -32350 51060 -31410
rect 51100 -32350 51160 -31410
rect 51200 -32350 51260 -31410
rect 51300 -32350 51360 -31410
rect 51400 -32350 51460 -31410
rect 51500 -32350 51560 -31410
rect 51600 -32350 51660 -31410
rect 51700 -32350 51760 -31410
rect 51800 -32350 51860 -31410
rect 51900 -32350 51960 -31410
rect 52000 -32350 52060 -31410
rect 52100 -32350 52160 -31410
rect 52200 -32350 52260 -31410
rect 52300 -32350 52360 -31410
rect 52400 -32350 52460 -31410
rect 52500 -32350 52560 -31410
rect 52600 -32350 52660 -31410
rect 52700 -32350 52760 -31410
rect 52800 -32350 52860 -31410
rect 52900 -32350 52960 -31410
rect 53000 -32340 53060 -31410
rect 49800 -34360 49860 -32980
rect 49900 -34370 49960 -32980
rect 50000 -34370 50060 -32980
rect 50100 -34370 50160 -32980
rect 50200 -34370 50260 -32980
rect 50300 -34370 50360 -32980
rect 50400 -34370 50460 -32980
rect 50500 -34370 50560 -32980
rect 50600 -34370 50660 -32980
rect 50700 -34370 50760 -32980
rect 50800 -34370 50860 -32980
rect 50900 -34370 50960 -32980
rect 51000 -34370 51060 -32980
rect 51100 -34370 51160 -32980
rect 51200 -34370 51260 -32980
rect 51300 -34370 51360 -32980
rect 51400 -34370 51460 -32980
rect 51500 -34370 51560 -32980
rect 51600 -34370 51660 -32980
rect 51700 -34370 51760 -32980
rect 51800 -34350 51860 -32990
rect 51900 -34350 51960 -33010
rect 52000 -34320 52060 -33030
rect 52700 -33070 52760 -33010
rect 52100 -34280 52160 -33070
rect 52200 -34220 52260 -33130
rect 52800 -33150 52860 -32980
rect 52300 -34130 52360 -33220
rect 52900 -33280 52960 -32980
rect 52400 -33990 52460 -33360
rect 53000 -33480 53060 -32980
rect 49800 -36340 49860 -35020
rect 49900 -36150 49960 -35020
rect 50000 -35970 50060 -35020
rect 50100 -35830 50160 -35020
rect 50200 -35880 50260 -35020
rect 50300 -35960 50360 -35020
rect 50400 -36050 50460 -35020
rect 50500 -36130 50560 -35020
rect 49700 -39360 49760 -37340
rect 50300 -37420 50360 -36750
rect 50400 -37570 50460 -36470
rect 50500 -37650 50560 -36300
rect 50600 -37680 50660 -35020
rect 50700 -37700 50760 -35020
rect 50800 -37680 50860 -35020
rect 50900 -37610 50960 -35020
rect 51000 -37470 51060 -35020
rect 51100 -36640 51160 -35020
rect 51200 -36210 51260 -35020
rect 51300 -36040 51360 -35020
rect 51400 -35930 51460 -35020
rect 51500 -35860 51560 -35020
rect 51600 -35810 51660 -35020
rect 51700 -35770 51760 -35020
rect 51800 -35740 51860 -35020
rect 51900 -35730 51960 -35020
rect 52000 -35710 52060 -35010
rect 52100 -35710 52160 -34990
rect 52200 -35730 52260 -34980
rect 52300 -35740 52360 -34950
rect 52400 -35780 52460 -34930
rect 52500 -35820 52560 -34880
rect 52600 -35890 52660 -34810
rect 52700 -35980 52760 -34720
rect 52800 -36100 52860 -34610
rect 52900 -36270 52960 -34490
rect 49800 -38870 49860 -37730
rect 49900 -38880 49960 -37920
rect 50000 -38880 50060 -38050
rect 50100 -38870 50160 -38150
rect 50200 -39360 50260 -38210
rect 50300 -39380 50360 -38260
rect 50400 -39380 50460 -38290
rect 50500 -39380 50560 -38330
rect 50600 -39380 50660 -38330
rect 50700 -39380 50760 -38330
rect 50800 -39380 50860 -38330
rect 50900 -39380 50960 -38320
rect 51000 -39380 51060 -38290
rect 51100 -39380 51160 -38250
rect 51200 -39380 51260 -38190
rect 51300 -39380 51360 -38110
rect 51400 -39380 51460 -37990
rect 51500 -39380 51560 -37830
rect 51600 -39380 51660 -37500
rect 51700 -39380 51760 -36600
rect 51800 -39380 51860 -36440
rect 51900 -39380 51960 -36380
rect 52000 -39380 52060 -36370
rect 52100 -38080 52160 -36370
rect 52200 -37960 52260 -36390
rect 52300 -37830 52360 -36450
rect 53000 -36530 53060 -34290
rect 52400 -37630 52460 -36560
rect 52500 -37130 52560 -36960
rect 52100 -39380 52160 -38140
rect 52200 -39380 52260 -38230
rect 52300 -39360 52360 -38330
rect 52400 -39300 52460 -38440
rect 52500 -38880 52560 -38520
rect 52600 -38880 52660 -38430
rect 52700 -38880 52760 -38300
rect 52800 -38880 52860 -38130
rect 52900 -38880 52960 -37940
rect 53000 -38870 53060 -37670
rect 48600 -41840 48660 -41640
rect 48700 -42250 48760 -41620
rect 48600 -48580 48660 -42520
rect 48800 -42770 48860 -39810
rect 48700 -48580 48760 -43090
rect 48900 -43540 48960 -40030
rect 48800 -48580 48860 -44510
rect 49000 -44820 49060 -40030
rect 48900 -48580 48960 -45100
rect 49100 -45350 49160 -40030
rect 49200 -43610 49260 -40030
rect 49300 -43660 49360 -40030
rect 49400 -43710 49460 -40030
rect 49500 -43760 49560 -40030
rect 49600 -43810 49660 -40030
rect 49700 -42050 49760 -40040
rect 49800 -41570 49860 -40360
rect 49900 -41370 49960 -40360
rect 50000 -41230 50060 -40360
rect 50100 -41140 50160 -40370
rect 50200 -41080 50260 -40040
rect 50300 -41030 50360 -40030
rect 50400 -41000 50460 -40030
rect 50500 -40970 50560 -40030
rect 50600 -40960 50660 -40030
rect 50700 -40960 50760 -40030
rect 50800 -40960 50860 -40030
rect 50900 -40960 50960 -40030
rect 51000 -40960 51060 -40030
rect 51100 -40960 51160 -40030
rect 51200 -40960 51260 -40030
rect 51300 -40960 51360 -40030
rect 51400 -40960 51460 -40030
rect 51500 -40960 51560 -40030
rect 51600 -40960 51660 -40030
rect 51700 -40960 51760 -40030
rect 51800 -40960 51860 -40030
rect 51900 -40960 51960 -40030
rect 52000 -40960 52060 -40030
rect 52100 -40960 52160 -40030
rect 52200 -40960 52260 -40030
rect 52300 -40960 52360 -40020
rect 52400 -40960 52460 -40000
rect 52500 -40960 52560 -39990
rect 52600 -40960 52660 -39950
rect 52700 -40960 52760 -39900
rect 52800 -40960 52860 -39820
rect 52900 -40960 52960 -39700
rect 53000 -40950 53060 -39500
rect 49700 -43860 49760 -42540
rect 50300 -42690 50360 -41920
rect 50400 -42850 50460 -41720
rect 49000 -48580 49060 -45660
rect 49100 -48580 49160 -46690
rect 49200 -48580 49260 -43860
rect 49800 -43910 49860 -42990
rect 49900 -43960 49960 -43160
rect 50000 -44010 50060 -43300
rect 50100 -44060 50160 -43400
rect 50200 -44110 50260 -43360
rect 50300 -44170 50360 -43230
rect 50400 -44220 50460 -43100
rect 50500 -44270 50560 -41650
rect 50600 -44320 50660 -41600
rect 49300 -48580 49360 -44340
rect 50700 -44370 50760 -41590
rect 49400 -46040 49460 -44380
rect 50800 -44420 50860 -41590
rect 49500 -45370 49560 -44430
rect 50900 -44470 50960 -41600
rect 49600 -45320 49660 -44480
rect 51000 -44520 51060 -41590
rect 49700 -45270 49760 -44530
rect 51100 -44570 51160 -41610
rect 51700 -42850 51760 -41600
rect 51800 -42950 51860 -41600
rect 51900 -43010 51960 -41600
rect 52000 -43020 52060 -41600
rect 52100 -43020 52160 -41600
rect 52200 -43000 52260 -41640
rect 52800 -41680 52860 -41600
rect 52300 -42940 52360 -41680
rect 52900 -41760 52960 -41590
rect 52400 -42830 52460 -41760
rect 53000 -41930 53060 -41600
rect 52500 -42510 52560 -42120
rect 49800 -45220 49860 -44570
rect 51200 -44580 51260 -43050
rect 51300 -44580 51360 -43240
rect 51400 -44580 51460 -43360
rect 51500 -44580 51560 -43440
rect 51600 -44580 51660 -43510
rect 51700 -44580 51760 -43560
rect 51800 -44580 51860 -43600
rect 51900 -44580 51960 -43610
rect 52000 -44580 52060 -43640
rect 52100 -44580 52160 -43640
rect 52200 -44580 52260 -43630
rect 52300 -44580 52360 -43600
rect 52400 -44580 52460 -43580
rect 52500 -44580 52560 -43540
rect 52600 -44580 52660 -43480
rect 52700 -44580 52760 -43400
rect 52800 -44580 52860 -43300
rect 52900 -44580 52960 -43170
rect 53000 -44580 53060 -42960
rect 49900 -45180 49960 -44630
rect 50000 -45130 50060 -44670
rect 50100 -45080 50160 -44720
rect 50200 -45030 50260 -44770
rect 50300 -44980 50360 -44820
rect 50400 -44930 50460 -44860
rect 49400 -48580 49460 -46100
rect 49500 -48580 49560 -46040
rect 49600 -48580 49660 -45990
rect 49700 -48580 49760 -45940
rect 49800 -48580 49860 -45890
rect 49900 -48580 49960 -45840
rect 50000 -48580 50060 -45780
rect 50100 -48580 50160 -45740
rect 50200 -48580 50260 -45690
rect 50300 -48580 50360 -45640
rect 50400 -48580 50460 -45580
rect 50500 -48580 50560 -45530
rect 50600 -48580 50660 -45480
rect 50700 -48580 50760 -45430
rect 50800 -48580 50860 -45380
rect 50900 -48580 50960 -45330
rect 51000 -48580 51060 -45270
rect 51100 -48580 51160 -45230
rect 51200 -48580 51260 -45210
rect 51300 -48580 51360 -45210
rect 51400 -48580 51460 -45210
rect 51500 -48580 51560 -45210
rect 51600 -48580 51660 -45210
rect 51700 -48580 51760 -45210
rect 51800 -48580 51860 -45210
rect 51900 -48580 51960 -45210
rect 52000 -48580 52060 -45210
rect 52100 -48580 52160 -45210
rect 52200 -48580 52260 -45210
rect 52300 -48580 52360 -45210
rect 52400 -48580 52460 -45210
rect 52500 -48580 52560 -45210
rect 52600 -48580 52660 -45210
rect 52700 -48580 52760 -45210
rect 52800 -48580 52860 -45210
rect 52900 -48580 52960 -45210
rect 53000 -48580 53060 -45220
rect 53100 -48580 53160 0
rect 53200 -48580 53260 0
rect 53300 -48580 53360 0
rect 53400 -48580 53460 0
rect 53500 -48580 53560 0
rect 53600 -48580 53660 0
rect 53700 -48580 53760 0
rect 53800 -48580 53860 0
rect 53900 -48580 53960 0
rect 54000 -48580 54060 0
rect 54100 -48580 54160 0
rect 54200 -48580 54260 0
rect 54300 -48580 54360 0
rect 54400 -48580 54460 0
rect 54500 -48580 54560 0
rect 54600 -48580 54660 0
rect 54700 -48580 54760 0
rect 54800 -48580 54860 0
rect 54900 -48580 54960 0
<< end >>
