magic
tech sky130B
magscale 1 2
timestamp 1659841776
<< error_p >>
rect 2138 3513 2196 3519
rect 2256 3513 2314 3519
rect 2374 3513 2432 3519
rect 2492 3513 2550 3519
rect 2610 3513 2668 3519
rect 2728 3513 2786 3519
rect 2846 3513 2904 3519
rect 2964 3513 3022 3519
rect 3082 3513 3140 3519
rect 3200 3513 3258 3519
rect 3318 3513 3376 3519
rect 3436 3513 3494 3519
rect 3554 3513 3612 3519
rect 3672 3513 3730 3519
rect 3790 3513 3848 3519
rect 3908 3513 3966 3519
rect 4026 3513 4084 3519
rect 4144 3513 4202 3519
rect 4262 3513 4320 3519
rect 4380 3513 4438 3519
rect 4498 3513 4556 3519
rect 4616 3513 4674 3519
rect 4734 3513 4792 3519
rect 4852 3513 4910 3519
rect 4970 3513 5028 3519
rect 5088 3513 5146 3519
rect 2138 3479 2150 3513
rect 2256 3479 2268 3513
rect 2374 3479 2386 3513
rect 2492 3479 2504 3513
rect 2610 3479 2622 3513
rect 2728 3479 2740 3513
rect 2846 3479 2858 3513
rect 2964 3479 2976 3513
rect 3082 3479 3094 3513
rect 3200 3479 3212 3513
rect 3318 3479 3330 3513
rect 3436 3479 3448 3513
rect 3554 3479 3566 3513
rect 3672 3479 3684 3513
rect 3790 3479 3802 3513
rect 3908 3479 3920 3513
rect 4026 3479 4038 3513
rect 4144 3479 4156 3513
rect 4262 3479 4274 3513
rect 4380 3479 4392 3513
rect 4498 3479 4510 3513
rect 4616 3479 4628 3513
rect 4734 3479 4746 3513
rect 4852 3479 4864 3513
rect 4970 3479 4982 3513
rect 5088 3479 5100 3513
rect 2138 3473 2196 3479
rect 2256 3473 2314 3479
rect 2374 3473 2432 3479
rect 2492 3473 2550 3479
rect 2610 3473 2668 3479
rect 2728 3473 2786 3479
rect 2846 3473 2904 3479
rect 2964 3473 3022 3479
rect 3082 3473 3140 3479
rect 3200 3473 3258 3479
rect 3318 3473 3376 3479
rect 3436 3473 3494 3479
rect 3554 3473 3612 3479
rect 3672 3473 3730 3479
rect 3790 3473 3848 3479
rect 3908 3473 3966 3479
rect 4026 3473 4084 3479
rect 4144 3473 4202 3479
rect 4262 3473 4320 3479
rect 4380 3473 4438 3479
rect 4498 3473 4556 3479
rect 4616 3473 4674 3479
rect 4734 3473 4792 3479
rect 4852 3473 4910 3479
rect 4970 3473 5028 3479
rect 5088 3473 5146 3479
rect 2138 3185 2196 3191
rect 2256 3185 2314 3191
rect 2374 3185 2432 3191
rect 2492 3185 2550 3191
rect 2610 3185 2668 3191
rect 2728 3185 2786 3191
rect 2846 3185 2904 3191
rect 2964 3185 3022 3191
rect 3082 3185 3140 3191
rect 3200 3185 3258 3191
rect 3318 3185 3376 3191
rect 3436 3185 3494 3191
rect 3554 3185 3612 3191
rect 3672 3185 3730 3191
rect 3790 3185 3848 3191
rect 3908 3185 3966 3191
rect 4026 3185 4084 3191
rect 4144 3185 4202 3191
rect 4262 3185 4320 3191
rect 4380 3185 4438 3191
rect 4498 3185 4556 3191
rect 4616 3185 4674 3191
rect 4734 3185 4792 3191
rect 4852 3185 4910 3191
rect 4970 3185 5028 3191
rect 5088 3185 5146 3191
rect 2138 3151 2150 3185
rect 2256 3151 2268 3185
rect 2374 3151 2386 3185
rect 2492 3151 2504 3185
rect 2610 3151 2622 3185
rect 2728 3151 2740 3185
rect 2846 3151 2858 3185
rect 2964 3151 2976 3185
rect 3082 3151 3094 3185
rect 3200 3151 3212 3185
rect 3318 3151 3330 3185
rect 3436 3151 3448 3185
rect 3554 3151 3566 3185
rect 3672 3151 3684 3185
rect 3790 3151 3802 3185
rect 3908 3151 3920 3185
rect 4026 3151 4038 3185
rect 4144 3151 4156 3185
rect 4262 3151 4274 3185
rect 4380 3151 4392 3185
rect 4498 3151 4510 3185
rect 4616 3151 4628 3185
rect 4734 3151 4746 3185
rect 4852 3151 4864 3185
rect 4970 3151 4982 3185
rect 5088 3151 5100 3185
rect 2138 3145 2196 3151
rect 2256 3145 2314 3151
rect 2374 3145 2432 3151
rect 2492 3145 2550 3151
rect 2610 3145 2668 3151
rect 2728 3145 2786 3151
rect 2846 3145 2904 3151
rect 2964 3145 3022 3151
rect 3082 3145 3140 3151
rect 3200 3145 3258 3151
rect 3318 3145 3376 3151
rect 3436 3145 3494 3151
rect 3554 3145 3612 3151
rect 3672 3145 3730 3151
rect 3790 3145 3848 3151
rect 3908 3145 3966 3151
rect 4026 3145 4084 3151
rect 4144 3145 4202 3151
rect 4262 3145 4320 3151
rect 4380 3145 4438 3151
rect 4498 3145 4556 3151
rect 4616 3145 4674 3151
rect 4734 3145 4792 3151
rect 4852 3145 4910 3151
rect 4970 3145 5028 3151
rect 5088 3145 5146 3151
rect 2138 3077 2196 3083
rect 2256 3077 2314 3083
rect 2374 3077 2432 3083
rect 2492 3077 2550 3083
rect 2610 3077 2668 3083
rect 2728 3077 2786 3083
rect 2846 3077 2904 3083
rect 2964 3077 3022 3083
rect 3082 3077 3140 3083
rect 3200 3077 3258 3083
rect 3318 3077 3376 3083
rect 3436 3077 3494 3083
rect 3554 3077 3612 3083
rect 3672 3077 3730 3083
rect 3790 3077 3848 3083
rect 3908 3077 3966 3083
rect 4026 3077 4084 3083
rect 4144 3077 4202 3083
rect 4262 3077 4320 3083
rect 4380 3077 4438 3083
rect 4498 3077 4556 3083
rect 4616 3077 4674 3083
rect 4734 3077 4792 3083
rect 4852 3077 4910 3083
rect 4970 3077 5028 3083
rect 5088 3077 5146 3083
rect 2138 3043 2150 3077
rect 2256 3043 2268 3077
rect 2374 3043 2386 3077
rect 2492 3043 2504 3077
rect 2610 3043 2622 3077
rect 2728 3043 2740 3077
rect 2846 3043 2858 3077
rect 2964 3043 2976 3077
rect 3082 3043 3094 3077
rect 3200 3043 3212 3077
rect 3318 3043 3330 3077
rect 3436 3043 3448 3077
rect 3554 3043 3566 3077
rect 3672 3043 3684 3077
rect 3790 3043 3802 3077
rect 3908 3043 3920 3077
rect 4026 3043 4038 3077
rect 4144 3043 4156 3077
rect 4262 3043 4274 3077
rect 4380 3043 4392 3077
rect 4498 3043 4510 3077
rect 4616 3043 4628 3077
rect 4734 3043 4746 3077
rect 4852 3043 4864 3077
rect 4970 3043 4982 3077
rect 5088 3043 5100 3077
rect 2138 3037 2196 3043
rect 2256 3037 2314 3043
rect 2374 3037 2432 3043
rect 2492 3037 2550 3043
rect 2610 3037 2668 3043
rect 2728 3037 2786 3043
rect 2846 3037 2904 3043
rect 2964 3037 3022 3043
rect 3082 3037 3140 3043
rect 3200 3037 3258 3043
rect 3318 3037 3376 3043
rect 3436 3037 3494 3043
rect 3554 3037 3612 3043
rect 3672 3037 3730 3043
rect 3790 3037 3848 3043
rect 3908 3037 3966 3043
rect 4026 3037 4084 3043
rect 4144 3037 4202 3043
rect 4262 3037 4320 3043
rect 4380 3037 4438 3043
rect 4498 3037 4556 3043
rect 4616 3037 4674 3043
rect 4734 3037 4792 3043
rect 4852 3037 4910 3043
rect 4970 3037 5028 3043
rect 5088 3037 5146 3043
rect 2138 2749 2196 2755
rect 2256 2749 2314 2755
rect 2374 2749 2432 2755
rect 2492 2749 2550 2755
rect 2610 2749 2668 2755
rect 2728 2749 2786 2755
rect 2846 2749 2904 2755
rect 2964 2749 3022 2755
rect 3082 2749 3140 2755
rect 3200 2749 3258 2755
rect 3318 2749 3376 2755
rect 3436 2749 3494 2755
rect 3554 2749 3612 2755
rect 3672 2749 3730 2755
rect 3790 2749 3848 2755
rect 3908 2749 3966 2755
rect 4026 2749 4084 2755
rect 4144 2749 4202 2755
rect 4262 2749 4320 2755
rect 4380 2749 4438 2755
rect 4498 2749 4556 2755
rect 4616 2749 4674 2755
rect 4734 2749 4792 2755
rect 4852 2749 4910 2755
rect 4970 2749 5028 2755
rect 5088 2749 5146 2755
rect 2138 2715 2150 2749
rect 2256 2715 2268 2749
rect 2374 2715 2386 2749
rect 2492 2715 2504 2749
rect 2610 2715 2622 2749
rect 2728 2715 2740 2749
rect 2846 2715 2858 2749
rect 2964 2715 2976 2749
rect 3082 2715 3094 2749
rect 3200 2715 3212 2749
rect 3318 2715 3330 2749
rect 3436 2715 3448 2749
rect 3554 2715 3566 2749
rect 3672 2715 3684 2749
rect 3790 2715 3802 2749
rect 3908 2715 3920 2749
rect 4026 2715 4038 2749
rect 4144 2715 4156 2749
rect 4262 2715 4274 2749
rect 4380 2715 4392 2749
rect 4498 2715 4510 2749
rect 4616 2715 4628 2749
rect 4734 2715 4746 2749
rect 4852 2715 4864 2749
rect 4970 2715 4982 2749
rect 5088 2715 5100 2749
rect 2138 2709 2196 2715
rect 2256 2709 2314 2715
rect 2374 2709 2432 2715
rect 2492 2709 2550 2715
rect 2610 2709 2668 2715
rect 2728 2709 2786 2715
rect 2846 2709 2904 2715
rect 2964 2709 3022 2715
rect 3082 2709 3140 2715
rect 3200 2709 3258 2715
rect 3318 2709 3376 2715
rect 3436 2709 3494 2715
rect 3554 2709 3612 2715
rect 3672 2709 3730 2715
rect 3790 2709 3848 2715
rect 3908 2709 3966 2715
rect 4026 2709 4084 2715
rect 4144 2709 4202 2715
rect 4262 2709 4320 2715
rect 4380 2709 4438 2715
rect 4498 2709 4556 2715
rect 4616 2709 4674 2715
rect 4734 2709 4792 2715
rect 4852 2709 4910 2715
rect 4970 2709 5028 2715
rect 5088 2709 5146 2715
rect 2138 2641 2196 2647
rect 2256 2641 2314 2647
rect 2374 2641 2432 2647
rect 2492 2641 2550 2647
rect 2610 2641 2668 2647
rect 2728 2641 2786 2647
rect 2846 2641 2904 2647
rect 2964 2641 3022 2647
rect 3082 2641 3140 2647
rect 3200 2641 3258 2647
rect 3318 2641 3376 2647
rect 3436 2641 3494 2647
rect 3554 2641 3612 2647
rect 3672 2641 3730 2647
rect 3790 2641 3848 2647
rect 3908 2641 3966 2647
rect 4026 2641 4084 2647
rect 4144 2641 4202 2647
rect 4262 2641 4320 2647
rect 4380 2641 4438 2647
rect 4498 2641 4556 2647
rect 4616 2641 4674 2647
rect 4734 2641 4792 2647
rect 4852 2641 4910 2647
rect 4970 2641 5028 2647
rect 5088 2641 5146 2647
rect 2138 2607 2150 2641
rect 2256 2607 2268 2641
rect 2374 2607 2386 2641
rect 2492 2607 2504 2641
rect 2610 2607 2622 2641
rect 2728 2607 2740 2641
rect 2846 2607 2858 2641
rect 2964 2607 2976 2641
rect 3082 2607 3094 2641
rect 3200 2607 3212 2641
rect 3318 2607 3330 2641
rect 3436 2607 3448 2641
rect 3554 2607 3566 2641
rect 3672 2607 3684 2641
rect 3790 2607 3802 2641
rect 3908 2607 3920 2641
rect 4026 2607 4038 2641
rect 4144 2607 4156 2641
rect 4262 2607 4274 2641
rect 4380 2607 4392 2641
rect 4498 2607 4510 2641
rect 4616 2607 4628 2641
rect 4734 2607 4746 2641
rect 4852 2607 4864 2641
rect 4970 2607 4982 2641
rect 5088 2607 5100 2641
rect 2138 2601 2196 2607
rect 2256 2601 2314 2607
rect 2374 2601 2432 2607
rect 2492 2601 2550 2607
rect 2610 2601 2668 2607
rect 2728 2601 2786 2607
rect 2846 2601 2904 2607
rect 2964 2601 3022 2607
rect 3082 2601 3140 2607
rect 3200 2601 3258 2607
rect 3318 2601 3376 2607
rect 3436 2601 3494 2607
rect 3554 2601 3612 2607
rect 3672 2601 3730 2607
rect 3790 2601 3848 2607
rect 3908 2601 3966 2607
rect 4026 2601 4084 2607
rect 4144 2601 4202 2607
rect 4262 2601 4320 2607
rect 4380 2601 4438 2607
rect 4498 2601 4556 2607
rect 4616 2601 4674 2607
rect 4734 2601 4792 2607
rect 4852 2601 4910 2607
rect 4970 2601 5028 2607
rect 5088 2601 5146 2607
rect 2138 2313 2196 2319
rect 2256 2313 2314 2319
rect 2374 2313 2432 2319
rect 2492 2313 2550 2319
rect 2610 2313 2668 2319
rect 2728 2313 2786 2319
rect 2846 2313 2904 2319
rect 2964 2313 3022 2319
rect 3082 2313 3140 2319
rect 3200 2313 3258 2319
rect 3318 2313 3376 2319
rect 3436 2313 3494 2319
rect 3554 2313 3612 2319
rect 3672 2313 3730 2319
rect 3790 2313 3848 2319
rect 3908 2313 3966 2319
rect 4026 2313 4084 2319
rect 4144 2313 4202 2319
rect 4262 2313 4320 2319
rect 4380 2313 4438 2319
rect 4498 2313 4556 2319
rect 4616 2313 4674 2319
rect 4734 2313 4792 2319
rect 4852 2313 4910 2319
rect 4970 2313 5028 2319
rect 5088 2313 5146 2319
rect 2138 2279 2150 2313
rect 2256 2279 2268 2313
rect 2374 2279 2386 2313
rect 2492 2279 2504 2313
rect 2610 2279 2622 2313
rect 2728 2279 2740 2313
rect 2846 2279 2858 2313
rect 2964 2279 2976 2313
rect 3082 2279 3094 2313
rect 3200 2279 3212 2313
rect 3318 2279 3330 2313
rect 3436 2279 3448 2313
rect 3554 2279 3566 2313
rect 3672 2279 3684 2313
rect 3790 2279 3802 2313
rect 3908 2279 3920 2313
rect 4026 2279 4038 2313
rect 4144 2279 4156 2313
rect 4262 2279 4274 2313
rect 4380 2279 4392 2313
rect 4498 2279 4510 2313
rect 4616 2279 4628 2313
rect 4734 2279 4746 2313
rect 4852 2279 4864 2313
rect 4970 2279 4982 2313
rect 5088 2279 5100 2313
rect 2138 2273 2196 2279
rect 2256 2273 2314 2279
rect 2374 2273 2432 2279
rect 2492 2273 2550 2279
rect 2610 2273 2668 2279
rect 2728 2273 2786 2279
rect 2846 2273 2904 2279
rect 2964 2273 3022 2279
rect 3082 2273 3140 2279
rect 3200 2273 3258 2279
rect 3318 2273 3376 2279
rect 3436 2273 3494 2279
rect 3554 2273 3612 2279
rect 3672 2273 3730 2279
rect 3790 2273 3848 2279
rect 3908 2273 3966 2279
rect 4026 2273 4084 2279
rect 4144 2273 4202 2279
rect 4262 2273 4320 2279
rect 4380 2273 4438 2279
rect 4498 2273 4556 2279
rect 4616 2273 4674 2279
rect 4734 2273 4792 2279
rect 4852 2273 4910 2279
rect 4970 2273 5028 2279
rect 5088 2273 5146 2279
use sky130_fd_pr__pfet_01v8_4XGD6H  sky130_fd_pr__pfet_01v8_4XGD6H_0
timestamp 1659841776
transform 1 0 3642 0 1 2896
box -1701 -755 1701 755
<< end >>
