magic
tech sky130B
magscale 1 2
timestamp 1659840519
<< error_p >>
rect -2743 617 -2685 623
rect -2625 617 -2567 623
rect -2507 617 -2449 623
rect -2389 617 -2331 623
rect -2271 617 -2213 623
rect -2153 617 -2095 623
rect -2035 617 -1977 623
rect -1917 617 -1859 623
rect -1799 617 -1741 623
rect -1681 617 -1623 623
rect -1563 617 -1505 623
rect -1445 617 -1387 623
rect -1327 617 -1269 623
rect -1209 617 -1151 623
rect -1091 617 -1033 623
rect -973 617 -915 623
rect -855 617 -797 623
rect -737 617 -679 623
rect -619 617 -561 623
rect -501 617 -443 623
rect -383 617 -325 623
rect -265 617 -207 623
rect -147 617 -89 623
rect -29 617 29 623
rect 89 617 147 623
rect 207 617 265 623
rect 325 617 383 623
rect 443 617 501 623
rect 561 617 619 623
rect 679 617 737 623
rect 797 617 855 623
rect 915 617 973 623
rect 1033 617 1091 623
rect 1151 617 1209 623
rect 1269 617 1327 623
rect 1387 617 1445 623
rect 1505 617 1563 623
rect 1623 617 1681 623
rect 1741 617 1799 623
rect 1859 617 1917 623
rect 1977 617 2035 623
rect 2095 617 2153 623
rect 2213 617 2271 623
rect 2331 617 2389 623
rect 2449 617 2507 623
rect 2567 617 2625 623
rect 2685 617 2743 623
rect -2743 583 -2731 617
rect -2625 583 -2613 617
rect -2507 583 -2495 617
rect -2389 583 -2377 617
rect -2271 583 -2259 617
rect -2153 583 -2141 617
rect -2035 583 -2023 617
rect -1917 583 -1905 617
rect -1799 583 -1787 617
rect -1681 583 -1669 617
rect -1563 583 -1551 617
rect -1445 583 -1433 617
rect -1327 583 -1315 617
rect -1209 583 -1197 617
rect -1091 583 -1079 617
rect -973 583 -961 617
rect -855 583 -843 617
rect -737 583 -725 617
rect -619 583 -607 617
rect -501 583 -489 617
rect -383 583 -371 617
rect -265 583 -253 617
rect -147 583 -135 617
rect -29 583 -17 617
rect 89 583 101 617
rect 207 583 219 617
rect 325 583 337 617
rect 443 583 455 617
rect 561 583 573 617
rect 679 583 691 617
rect 797 583 809 617
rect 915 583 927 617
rect 1033 583 1045 617
rect 1151 583 1163 617
rect 1269 583 1281 617
rect 1387 583 1399 617
rect 1505 583 1517 617
rect 1623 583 1635 617
rect 1741 583 1753 617
rect 1859 583 1871 617
rect 1977 583 1989 617
rect 2095 583 2107 617
rect 2213 583 2225 617
rect 2331 583 2343 617
rect 2449 583 2461 617
rect 2567 583 2579 617
rect 2685 583 2697 617
rect -2743 577 -2685 583
rect -2625 577 -2567 583
rect -2507 577 -2449 583
rect -2389 577 -2331 583
rect -2271 577 -2213 583
rect -2153 577 -2095 583
rect -2035 577 -1977 583
rect -1917 577 -1859 583
rect -1799 577 -1741 583
rect -1681 577 -1623 583
rect -1563 577 -1505 583
rect -1445 577 -1387 583
rect -1327 577 -1269 583
rect -1209 577 -1151 583
rect -1091 577 -1033 583
rect -973 577 -915 583
rect -855 577 -797 583
rect -737 577 -679 583
rect -619 577 -561 583
rect -501 577 -443 583
rect -383 577 -325 583
rect -265 577 -207 583
rect -147 577 -89 583
rect -29 577 29 583
rect 89 577 147 583
rect 207 577 265 583
rect 325 577 383 583
rect 443 577 501 583
rect 561 577 619 583
rect 679 577 737 583
rect 797 577 855 583
rect 915 577 973 583
rect 1033 577 1091 583
rect 1151 577 1209 583
rect 1269 577 1327 583
rect 1387 577 1445 583
rect 1505 577 1563 583
rect 1623 577 1681 583
rect 1741 577 1799 583
rect 1859 577 1917 583
rect 1977 577 2035 583
rect 2095 577 2153 583
rect 2213 577 2271 583
rect 2331 577 2389 583
rect 2449 577 2507 583
rect 2567 577 2625 583
rect 2685 577 2743 583
rect -2743 289 -2685 295
rect -2625 289 -2567 295
rect -2507 289 -2449 295
rect -2389 289 -2331 295
rect -2271 289 -2213 295
rect -2153 289 -2095 295
rect -2035 289 -1977 295
rect -1917 289 -1859 295
rect -1799 289 -1741 295
rect -1681 289 -1623 295
rect -1563 289 -1505 295
rect -1445 289 -1387 295
rect -1327 289 -1269 295
rect -1209 289 -1151 295
rect -1091 289 -1033 295
rect -973 289 -915 295
rect -855 289 -797 295
rect -737 289 -679 295
rect -619 289 -561 295
rect -501 289 -443 295
rect -383 289 -325 295
rect -265 289 -207 295
rect -147 289 -89 295
rect -29 289 29 295
rect 89 289 147 295
rect 207 289 265 295
rect 325 289 383 295
rect 443 289 501 295
rect 561 289 619 295
rect 679 289 737 295
rect 797 289 855 295
rect 915 289 973 295
rect 1033 289 1091 295
rect 1151 289 1209 295
rect 1269 289 1327 295
rect 1387 289 1445 295
rect 1505 289 1563 295
rect 1623 289 1681 295
rect 1741 289 1799 295
rect 1859 289 1917 295
rect 1977 289 2035 295
rect 2095 289 2153 295
rect 2213 289 2271 295
rect 2331 289 2389 295
rect 2449 289 2507 295
rect 2567 289 2625 295
rect 2685 289 2743 295
rect -2743 255 -2731 289
rect -2625 255 -2613 289
rect -2507 255 -2495 289
rect -2389 255 -2377 289
rect -2271 255 -2259 289
rect -2153 255 -2141 289
rect -2035 255 -2023 289
rect -1917 255 -1905 289
rect -1799 255 -1787 289
rect -1681 255 -1669 289
rect -1563 255 -1551 289
rect -1445 255 -1433 289
rect -1327 255 -1315 289
rect -1209 255 -1197 289
rect -1091 255 -1079 289
rect -973 255 -961 289
rect -855 255 -843 289
rect -737 255 -725 289
rect -619 255 -607 289
rect -501 255 -489 289
rect -383 255 -371 289
rect -265 255 -253 289
rect -147 255 -135 289
rect -29 255 -17 289
rect 89 255 101 289
rect 207 255 219 289
rect 325 255 337 289
rect 443 255 455 289
rect 561 255 573 289
rect 679 255 691 289
rect 797 255 809 289
rect 915 255 927 289
rect 1033 255 1045 289
rect 1151 255 1163 289
rect 1269 255 1281 289
rect 1387 255 1399 289
rect 1505 255 1517 289
rect 1623 255 1635 289
rect 1741 255 1753 289
rect 1859 255 1871 289
rect 1977 255 1989 289
rect 2095 255 2107 289
rect 2213 255 2225 289
rect 2331 255 2343 289
rect 2449 255 2461 289
rect 2567 255 2579 289
rect 2685 255 2697 289
rect -2743 249 -2685 255
rect -2625 249 -2567 255
rect -2507 249 -2449 255
rect -2389 249 -2331 255
rect -2271 249 -2213 255
rect -2153 249 -2095 255
rect -2035 249 -1977 255
rect -1917 249 -1859 255
rect -1799 249 -1741 255
rect -1681 249 -1623 255
rect -1563 249 -1505 255
rect -1445 249 -1387 255
rect -1327 249 -1269 255
rect -1209 249 -1151 255
rect -1091 249 -1033 255
rect -973 249 -915 255
rect -855 249 -797 255
rect -737 249 -679 255
rect -619 249 -561 255
rect -501 249 -443 255
rect -383 249 -325 255
rect -265 249 -207 255
rect -147 249 -89 255
rect -29 249 29 255
rect 89 249 147 255
rect 207 249 265 255
rect 325 249 383 255
rect 443 249 501 255
rect 561 249 619 255
rect 679 249 737 255
rect 797 249 855 255
rect 915 249 973 255
rect 1033 249 1091 255
rect 1151 249 1209 255
rect 1269 249 1327 255
rect 1387 249 1445 255
rect 1505 249 1563 255
rect 1623 249 1681 255
rect 1741 249 1799 255
rect 1859 249 1917 255
rect 1977 249 2035 255
rect 2095 249 2153 255
rect 2213 249 2271 255
rect 2331 249 2389 255
rect 2449 249 2507 255
rect 2567 249 2625 255
rect 2685 249 2743 255
rect -2743 181 -2685 187
rect -2625 181 -2567 187
rect -2507 181 -2449 187
rect -2389 181 -2331 187
rect -2271 181 -2213 187
rect -2153 181 -2095 187
rect -2035 181 -1977 187
rect -1917 181 -1859 187
rect -1799 181 -1741 187
rect -1681 181 -1623 187
rect -1563 181 -1505 187
rect -1445 181 -1387 187
rect -1327 181 -1269 187
rect -1209 181 -1151 187
rect -1091 181 -1033 187
rect -973 181 -915 187
rect -855 181 -797 187
rect -737 181 -679 187
rect -619 181 -561 187
rect -501 181 -443 187
rect -383 181 -325 187
rect -265 181 -207 187
rect -147 181 -89 187
rect -29 181 29 187
rect 89 181 147 187
rect 207 181 265 187
rect 325 181 383 187
rect 443 181 501 187
rect 561 181 619 187
rect 679 181 737 187
rect 797 181 855 187
rect 915 181 973 187
rect 1033 181 1091 187
rect 1151 181 1209 187
rect 1269 181 1327 187
rect 1387 181 1445 187
rect 1505 181 1563 187
rect 1623 181 1681 187
rect 1741 181 1799 187
rect 1859 181 1917 187
rect 1977 181 2035 187
rect 2095 181 2153 187
rect 2213 181 2271 187
rect 2331 181 2389 187
rect 2449 181 2507 187
rect 2567 181 2625 187
rect 2685 181 2743 187
rect -2743 147 -2731 181
rect -2625 147 -2613 181
rect -2507 147 -2495 181
rect -2389 147 -2377 181
rect -2271 147 -2259 181
rect -2153 147 -2141 181
rect -2035 147 -2023 181
rect -1917 147 -1905 181
rect -1799 147 -1787 181
rect -1681 147 -1669 181
rect -1563 147 -1551 181
rect -1445 147 -1433 181
rect -1327 147 -1315 181
rect -1209 147 -1197 181
rect -1091 147 -1079 181
rect -973 147 -961 181
rect -855 147 -843 181
rect -737 147 -725 181
rect -619 147 -607 181
rect -501 147 -489 181
rect -383 147 -371 181
rect -265 147 -253 181
rect -147 147 -135 181
rect -29 147 -17 181
rect 89 147 101 181
rect 207 147 219 181
rect 325 147 337 181
rect 443 147 455 181
rect 561 147 573 181
rect 679 147 691 181
rect 797 147 809 181
rect 915 147 927 181
rect 1033 147 1045 181
rect 1151 147 1163 181
rect 1269 147 1281 181
rect 1387 147 1399 181
rect 1505 147 1517 181
rect 1623 147 1635 181
rect 1741 147 1753 181
rect 1859 147 1871 181
rect 1977 147 1989 181
rect 2095 147 2107 181
rect 2213 147 2225 181
rect 2331 147 2343 181
rect 2449 147 2461 181
rect 2567 147 2579 181
rect 2685 147 2697 181
rect -2743 141 -2685 147
rect -2625 141 -2567 147
rect -2507 141 -2449 147
rect -2389 141 -2331 147
rect -2271 141 -2213 147
rect -2153 141 -2095 147
rect -2035 141 -1977 147
rect -1917 141 -1859 147
rect -1799 141 -1741 147
rect -1681 141 -1623 147
rect -1563 141 -1505 147
rect -1445 141 -1387 147
rect -1327 141 -1269 147
rect -1209 141 -1151 147
rect -1091 141 -1033 147
rect -973 141 -915 147
rect -855 141 -797 147
rect -737 141 -679 147
rect -619 141 -561 147
rect -501 141 -443 147
rect -383 141 -325 147
rect -265 141 -207 147
rect -147 141 -89 147
rect -29 141 29 147
rect 89 141 147 147
rect 207 141 265 147
rect 325 141 383 147
rect 443 141 501 147
rect 561 141 619 147
rect 679 141 737 147
rect 797 141 855 147
rect 915 141 973 147
rect 1033 141 1091 147
rect 1151 141 1209 147
rect 1269 141 1327 147
rect 1387 141 1445 147
rect 1505 141 1563 147
rect 1623 141 1681 147
rect 1741 141 1799 147
rect 1859 141 1917 147
rect 1977 141 2035 147
rect 2095 141 2153 147
rect 2213 141 2271 147
rect 2331 141 2389 147
rect 2449 141 2507 147
rect 2567 141 2625 147
rect 2685 141 2743 147
rect -2743 -147 -2685 -141
rect -2625 -147 -2567 -141
rect -2507 -147 -2449 -141
rect -2389 -147 -2331 -141
rect -2271 -147 -2213 -141
rect -2153 -147 -2095 -141
rect -2035 -147 -1977 -141
rect -1917 -147 -1859 -141
rect -1799 -147 -1741 -141
rect -1681 -147 -1623 -141
rect -1563 -147 -1505 -141
rect -1445 -147 -1387 -141
rect -1327 -147 -1269 -141
rect -1209 -147 -1151 -141
rect -1091 -147 -1033 -141
rect -973 -147 -915 -141
rect -855 -147 -797 -141
rect -737 -147 -679 -141
rect -619 -147 -561 -141
rect -501 -147 -443 -141
rect -383 -147 -325 -141
rect -265 -147 -207 -141
rect -147 -147 -89 -141
rect -29 -147 29 -141
rect 89 -147 147 -141
rect 207 -147 265 -141
rect 325 -147 383 -141
rect 443 -147 501 -141
rect 561 -147 619 -141
rect 679 -147 737 -141
rect 797 -147 855 -141
rect 915 -147 973 -141
rect 1033 -147 1091 -141
rect 1151 -147 1209 -141
rect 1269 -147 1327 -141
rect 1387 -147 1445 -141
rect 1505 -147 1563 -141
rect 1623 -147 1681 -141
rect 1741 -147 1799 -141
rect 1859 -147 1917 -141
rect 1977 -147 2035 -141
rect 2095 -147 2153 -141
rect 2213 -147 2271 -141
rect 2331 -147 2389 -141
rect 2449 -147 2507 -141
rect 2567 -147 2625 -141
rect 2685 -147 2743 -141
rect -2743 -181 -2731 -147
rect -2625 -181 -2613 -147
rect -2507 -181 -2495 -147
rect -2389 -181 -2377 -147
rect -2271 -181 -2259 -147
rect -2153 -181 -2141 -147
rect -2035 -181 -2023 -147
rect -1917 -181 -1905 -147
rect -1799 -181 -1787 -147
rect -1681 -181 -1669 -147
rect -1563 -181 -1551 -147
rect -1445 -181 -1433 -147
rect -1327 -181 -1315 -147
rect -1209 -181 -1197 -147
rect -1091 -181 -1079 -147
rect -973 -181 -961 -147
rect -855 -181 -843 -147
rect -737 -181 -725 -147
rect -619 -181 -607 -147
rect -501 -181 -489 -147
rect -383 -181 -371 -147
rect -265 -181 -253 -147
rect -147 -181 -135 -147
rect -29 -181 -17 -147
rect 89 -181 101 -147
rect 207 -181 219 -147
rect 325 -181 337 -147
rect 443 -181 455 -147
rect 561 -181 573 -147
rect 679 -181 691 -147
rect 797 -181 809 -147
rect 915 -181 927 -147
rect 1033 -181 1045 -147
rect 1151 -181 1163 -147
rect 1269 -181 1281 -147
rect 1387 -181 1399 -147
rect 1505 -181 1517 -147
rect 1623 -181 1635 -147
rect 1741 -181 1753 -147
rect 1859 -181 1871 -147
rect 1977 -181 1989 -147
rect 2095 -181 2107 -147
rect 2213 -181 2225 -147
rect 2331 -181 2343 -147
rect 2449 -181 2461 -147
rect 2567 -181 2579 -147
rect 2685 -181 2697 -147
rect -2743 -187 -2685 -181
rect -2625 -187 -2567 -181
rect -2507 -187 -2449 -181
rect -2389 -187 -2331 -181
rect -2271 -187 -2213 -181
rect -2153 -187 -2095 -181
rect -2035 -187 -1977 -181
rect -1917 -187 -1859 -181
rect -1799 -187 -1741 -181
rect -1681 -187 -1623 -181
rect -1563 -187 -1505 -181
rect -1445 -187 -1387 -181
rect -1327 -187 -1269 -181
rect -1209 -187 -1151 -181
rect -1091 -187 -1033 -181
rect -973 -187 -915 -181
rect -855 -187 -797 -181
rect -737 -187 -679 -181
rect -619 -187 -561 -181
rect -501 -187 -443 -181
rect -383 -187 -325 -181
rect -265 -187 -207 -181
rect -147 -187 -89 -181
rect -29 -187 29 -181
rect 89 -187 147 -181
rect 207 -187 265 -181
rect 325 -187 383 -181
rect 443 -187 501 -181
rect 561 -187 619 -181
rect 679 -187 737 -181
rect 797 -187 855 -181
rect 915 -187 973 -181
rect 1033 -187 1091 -181
rect 1151 -187 1209 -181
rect 1269 -187 1327 -181
rect 1387 -187 1445 -181
rect 1505 -187 1563 -181
rect 1623 -187 1681 -181
rect 1741 -187 1799 -181
rect 1859 -187 1917 -181
rect 1977 -187 2035 -181
rect 2095 -187 2153 -181
rect 2213 -187 2271 -181
rect 2331 -187 2389 -181
rect 2449 -187 2507 -181
rect 2567 -187 2625 -181
rect 2685 -187 2743 -181
rect -2743 -255 -2685 -249
rect -2625 -255 -2567 -249
rect -2507 -255 -2449 -249
rect -2389 -255 -2331 -249
rect -2271 -255 -2213 -249
rect -2153 -255 -2095 -249
rect -2035 -255 -1977 -249
rect -1917 -255 -1859 -249
rect -1799 -255 -1741 -249
rect -1681 -255 -1623 -249
rect -1563 -255 -1505 -249
rect -1445 -255 -1387 -249
rect -1327 -255 -1269 -249
rect -1209 -255 -1151 -249
rect -1091 -255 -1033 -249
rect -973 -255 -915 -249
rect -855 -255 -797 -249
rect -737 -255 -679 -249
rect -619 -255 -561 -249
rect -501 -255 -443 -249
rect -383 -255 -325 -249
rect -265 -255 -207 -249
rect -147 -255 -89 -249
rect -29 -255 29 -249
rect 89 -255 147 -249
rect 207 -255 265 -249
rect 325 -255 383 -249
rect 443 -255 501 -249
rect 561 -255 619 -249
rect 679 -255 737 -249
rect 797 -255 855 -249
rect 915 -255 973 -249
rect 1033 -255 1091 -249
rect 1151 -255 1209 -249
rect 1269 -255 1327 -249
rect 1387 -255 1445 -249
rect 1505 -255 1563 -249
rect 1623 -255 1681 -249
rect 1741 -255 1799 -249
rect 1859 -255 1917 -249
rect 1977 -255 2035 -249
rect 2095 -255 2153 -249
rect 2213 -255 2271 -249
rect 2331 -255 2389 -249
rect 2449 -255 2507 -249
rect 2567 -255 2625 -249
rect 2685 -255 2743 -249
rect -2743 -289 -2731 -255
rect -2625 -289 -2613 -255
rect -2507 -289 -2495 -255
rect -2389 -289 -2377 -255
rect -2271 -289 -2259 -255
rect -2153 -289 -2141 -255
rect -2035 -289 -2023 -255
rect -1917 -289 -1905 -255
rect -1799 -289 -1787 -255
rect -1681 -289 -1669 -255
rect -1563 -289 -1551 -255
rect -1445 -289 -1433 -255
rect -1327 -289 -1315 -255
rect -1209 -289 -1197 -255
rect -1091 -289 -1079 -255
rect -973 -289 -961 -255
rect -855 -289 -843 -255
rect -737 -289 -725 -255
rect -619 -289 -607 -255
rect -501 -289 -489 -255
rect -383 -289 -371 -255
rect -265 -289 -253 -255
rect -147 -289 -135 -255
rect -29 -289 -17 -255
rect 89 -289 101 -255
rect 207 -289 219 -255
rect 325 -289 337 -255
rect 443 -289 455 -255
rect 561 -289 573 -255
rect 679 -289 691 -255
rect 797 -289 809 -255
rect 915 -289 927 -255
rect 1033 -289 1045 -255
rect 1151 -289 1163 -255
rect 1269 -289 1281 -255
rect 1387 -289 1399 -255
rect 1505 -289 1517 -255
rect 1623 -289 1635 -255
rect 1741 -289 1753 -255
rect 1859 -289 1871 -255
rect 1977 -289 1989 -255
rect 2095 -289 2107 -255
rect 2213 -289 2225 -255
rect 2331 -289 2343 -255
rect 2449 -289 2461 -255
rect 2567 -289 2579 -255
rect 2685 -289 2697 -255
rect -2743 -295 -2685 -289
rect -2625 -295 -2567 -289
rect -2507 -295 -2449 -289
rect -2389 -295 -2331 -289
rect -2271 -295 -2213 -289
rect -2153 -295 -2095 -289
rect -2035 -295 -1977 -289
rect -1917 -295 -1859 -289
rect -1799 -295 -1741 -289
rect -1681 -295 -1623 -289
rect -1563 -295 -1505 -289
rect -1445 -295 -1387 -289
rect -1327 -295 -1269 -289
rect -1209 -295 -1151 -289
rect -1091 -295 -1033 -289
rect -973 -295 -915 -289
rect -855 -295 -797 -289
rect -737 -295 -679 -289
rect -619 -295 -561 -289
rect -501 -295 -443 -289
rect -383 -295 -325 -289
rect -265 -295 -207 -289
rect -147 -295 -89 -289
rect -29 -295 29 -289
rect 89 -295 147 -289
rect 207 -295 265 -289
rect 325 -295 383 -289
rect 443 -295 501 -289
rect 561 -295 619 -289
rect 679 -295 737 -289
rect 797 -295 855 -289
rect 915 -295 973 -289
rect 1033 -295 1091 -289
rect 1151 -295 1209 -289
rect 1269 -295 1327 -289
rect 1387 -295 1445 -289
rect 1505 -295 1563 -289
rect 1623 -295 1681 -289
rect 1741 -295 1799 -289
rect 1859 -295 1917 -289
rect 1977 -295 2035 -289
rect 2095 -295 2153 -289
rect 2213 -295 2271 -289
rect 2331 -295 2389 -289
rect 2449 -295 2507 -289
rect 2567 -295 2625 -289
rect 2685 -295 2743 -289
rect -2743 -583 -2685 -577
rect -2625 -583 -2567 -577
rect -2507 -583 -2449 -577
rect -2389 -583 -2331 -577
rect -2271 -583 -2213 -577
rect -2153 -583 -2095 -577
rect -2035 -583 -1977 -577
rect -1917 -583 -1859 -577
rect -1799 -583 -1741 -577
rect -1681 -583 -1623 -577
rect -1563 -583 -1505 -577
rect -1445 -583 -1387 -577
rect -1327 -583 -1269 -577
rect -1209 -583 -1151 -577
rect -1091 -583 -1033 -577
rect -973 -583 -915 -577
rect -855 -583 -797 -577
rect -737 -583 -679 -577
rect -619 -583 -561 -577
rect -501 -583 -443 -577
rect -383 -583 -325 -577
rect -265 -583 -207 -577
rect -147 -583 -89 -577
rect -29 -583 29 -577
rect 89 -583 147 -577
rect 207 -583 265 -577
rect 325 -583 383 -577
rect 443 -583 501 -577
rect 561 -583 619 -577
rect 679 -583 737 -577
rect 797 -583 855 -577
rect 915 -583 973 -577
rect 1033 -583 1091 -577
rect 1151 -583 1209 -577
rect 1269 -583 1327 -577
rect 1387 -583 1445 -577
rect 1505 -583 1563 -577
rect 1623 -583 1681 -577
rect 1741 -583 1799 -577
rect 1859 -583 1917 -577
rect 1977 -583 2035 -577
rect 2095 -583 2153 -577
rect 2213 -583 2271 -577
rect 2331 -583 2389 -577
rect 2449 -583 2507 -577
rect 2567 -583 2625 -577
rect 2685 -583 2743 -577
rect -2743 -617 -2731 -583
rect -2625 -617 -2613 -583
rect -2507 -617 -2495 -583
rect -2389 -617 -2377 -583
rect -2271 -617 -2259 -583
rect -2153 -617 -2141 -583
rect -2035 -617 -2023 -583
rect -1917 -617 -1905 -583
rect -1799 -617 -1787 -583
rect -1681 -617 -1669 -583
rect -1563 -617 -1551 -583
rect -1445 -617 -1433 -583
rect -1327 -617 -1315 -583
rect -1209 -617 -1197 -583
rect -1091 -617 -1079 -583
rect -973 -617 -961 -583
rect -855 -617 -843 -583
rect -737 -617 -725 -583
rect -619 -617 -607 -583
rect -501 -617 -489 -583
rect -383 -617 -371 -583
rect -265 -617 -253 -583
rect -147 -617 -135 -583
rect -29 -617 -17 -583
rect 89 -617 101 -583
rect 207 -617 219 -583
rect 325 -617 337 -583
rect 443 -617 455 -583
rect 561 -617 573 -583
rect 679 -617 691 -583
rect 797 -617 809 -583
rect 915 -617 927 -583
rect 1033 -617 1045 -583
rect 1151 -617 1163 -583
rect 1269 -617 1281 -583
rect 1387 -617 1399 -583
rect 1505 -617 1517 -583
rect 1623 -617 1635 -583
rect 1741 -617 1753 -583
rect 1859 -617 1871 -583
rect 1977 -617 1989 -583
rect 2095 -617 2107 -583
rect 2213 -617 2225 -583
rect 2331 -617 2343 -583
rect 2449 -617 2461 -583
rect 2567 -617 2579 -583
rect 2685 -617 2697 -583
rect -2743 -623 -2685 -617
rect -2625 -623 -2567 -617
rect -2507 -623 -2449 -617
rect -2389 -623 -2331 -617
rect -2271 -623 -2213 -617
rect -2153 -623 -2095 -617
rect -2035 -623 -1977 -617
rect -1917 -623 -1859 -617
rect -1799 -623 -1741 -617
rect -1681 -623 -1623 -617
rect -1563 -623 -1505 -617
rect -1445 -623 -1387 -617
rect -1327 -623 -1269 -617
rect -1209 -623 -1151 -617
rect -1091 -623 -1033 -617
rect -973 -623 -915 -617
rect -855 -623 -797 -617
rect -737 -623 -679 -617
rect -619 -623 -561 -617
rect -501 -623 -443 -617
rect -383 -623 -325 -617
rect -265 -623 -207 -617
rect -147 -623 -89 -617
rect -29 -623 29 -617
rect 89 -623 147 -617
rect 207 -623 265 -617
rect 325 -623 383 -617
rect 443 -623 501 -617
rect 561 -623 619 -617
rect 679 -623 737 -617
rect 797 -623 855 -617
rect 915 -623 973 -617
rect 1033 -623 1091 -617
rect 1151 -623 1209 -617
rect 1269 -623 1327 -617
rect 1387 -623 1445 -617
rect 1505 -623 1563 -617
rect 1623 -623 1681 -617
rect 1741 -623 1799 -617
rect 1859 -623 1917 -617
rect 1977 -623 2035 -617
rect 2095 -623 2153 -617
rect 2213 -623 2271 -617
rect 2331 -623 2389 -617
rect 2449 -623 2507 -617
rect 2567 -623 2625 -617
rect 2685 -623 2743 -617
<< nwell >>
rect -2940 -755 2940 755
<< pmos >>
rect -2744 336 -2684 536
rect -2626 336 -2566 536
rect -2508 336 -2448 536
rect -2390 336 -2330 536
rect -2272 336 -2212 536
rect -2154 336 -2094 536
rect -2036 336 -1976 536
rect -1918 336 -1858 536
rect -1800 336 -1740 536
rect -1682 336 -1622 536
rect -1564 336 -1504 536
rect -1446 336 -1386 536
rect -1328 336 -1268 536
rect -1210 336 -1150 536
rect -1092 336 -1032 536
rect -974 336 -914 536
rect -856 336 -796 536
rect -738 336 -678 536
rect -620 336 -560 536
rect -502 336 -442 536
rect -384 336 -324 536
rect -266 336 -206 536
rect -148 336 -88 536
rect -30 336 30 536
rect 88 336 148 536
rect 206 336 266 536
rect 324 336 384 536
rect 442 336 502 536
rect 560 336 620 536
rect 678 336 738 536
rect 796 336 856 536
rect 914 336 974 536
rect 1032 336 1092 536
rect 1150 336 1210 536
rect 1268 336 1328 536
rect 1386 336 1446 536
rect 1504 336 1564 536
rect 1622 336 1682 536
rect 1740 336 1800 536
rect 1858 336 1918 536
rect 1976 336 2036 536
rect 2094 336 2154 536
rect 2212 336 2272 536
rect 2330 336 2390 536
rect 2448 336 2508 536
rect 2566 336 2626 536
rect 2684 336 2744 536
rect -2744 -100 -2684 100
rect -2626 -100 -2566 100
rect -2508 -100 -2448 100
rect -2390 -100 -2330 100
rect -2272 -100 -2212 100
rect -2154 -100 -2094 100
rect -2036 -100 -1976 100
rect -1918 -100 -1858 100
rect -1800 -100 -1740 100
rect -1682 -100 -1622 100
rect -1564 -100 -1504 100
rect -1446 -100 -1386 100
rect -1328 -100 -1268 100
rect -1210 -100 -1150 100
rect -1092 -100 -1032 100
rect -974 -100 -914 100
rect -856 -100 -796 100
rect -738 -100 -678 100
rect -620 -100 -560 100
rect -502 -100 -442 100
rect -384 -100 -324 100
rect -266 -100 -206 100
rect -148 -100 -88 100
rect -30 -100 30 100
rect 88 -100 148 100
rect 206 -100 266 100
rect 324 -100 384 100
rect 442 -100 502 100
rect 560 -100 620 100
rect 678 -100 738 100
rect 796 -100 856 100
rect 914 -100 974 100
rect 1032 -100 1092 100
rect 1150 -100 1210 100
rect 1268 -100 1328 100
rect 1386 -100 1446 100
rect 1504 -100 1564 100
rect 1622 -100 1682 100
rect 1740 -100 1800 100
rect 1858 -100 1918 100
rect 1976 -100 2036 100
rect 2094 -100 2154 100
rect 2212 -100 2272 100
rect 2330 -100 2390 100
rect 2448 -100 2508 100
rect 2566 -100 2626 100
rect 2684 -100 2744 100
rect -2744 -536 -2684 -336
rect -2626 -536 -2566 -336
rect -2508 -536 -2448 -336
rect -2390 -536 -2330 -336
rect -2272 -536 -2212 -336
rect -2154 -536 -2094 -336
rect -2036 -536 -1976 -336
rect -1918 -536 -1858 -336
rect -1800 -536 -1740 -336
rect -1682 -536 -1622 -336
rect -1564 -536 -1504 -336
rect -1446 -536 -1386 -336
rect -1328 -536 -1268 -336
rect -1210 -536 -1150 -336
rect -1092 -536 -1032 -336
rect -974 -536 -914 -336
rect -856 -536 -796 -336
rect -738 -536 -678 -336
rect -620 -536 -560 -336
rect -502 -536 -442 -336
rect -384 -536 -324 -336
rect -266 -536 -206 -336
rect -148 -536 -88 -336
rect -30 -536 30 -336
rect 88 -536 148 -336
rect 206 -536 266 -336
rect 324 -536 384 -336
rect 442 -536 502 -336
rect 560 -536 620 -336
rect 678 -536 738 -336
rect 796 -536 856 -336
rect 914 -536 974 -336
rect 1032 -536 1092 -336
rect 1150 -536 1210 -336
rect 1268 -536 1328 -336
rect 1386 -536 1446 -336
rect 1504 -536 1564 -336
rect 1622 -536 1682 -336
rect 1740 -536 1800 -336
rect 1858 -536 1918 -336
rect 1976 -536 2036 -336
rect 2094 -536 2154 -336
rect 2212 -536 2272 -336
rect 2330 -536 2390 -336
rect 2448 -536 2508 -336
rect 2566 -536 2626 -336
rect 2684 -536 2744 -336
<< pdiff >>
rect -2802 524 -2744 536
rect -2802 348 -2790 524
rect -2756 348 -2744 524
rect -2802 336 -2744 348
rect -2684 524 -2626 536
rect -2684 348 -2672 524
rect -2638 348 -2626 524
rect -2684 336 -2626 348
rect -2566 524 -2508 536
rect -2566 348 -2554 524
rect -2520 348 -2508 524
rect -2566 336 -2508 348
rect -2448 524 -2390 536
rect -2448 348 -2436 524
rect -2402 348 -2390 524
rect -2448 336 -2390 348
rect -2330 524 -2272 536
rect -2330 348 -2318 524
rect -2284 348 -2272 524
rect -2330 336 -2272 348
rect -2212 524 -2154 536
rect -2212 348 -2200 524
rect -2166 348 -2154 524
rect -2212 336 -2154 348
rect -2094 524 -2036 536
rect -2094 348 -2082 524
rect -2048 348 -2036 524
rect -2094 336 -2036 348
rect -1976 524 -1918 536
rect -1976 348 -1964 524
rect -1930 348 -1918 524
rect -1976 336 -1918 348
rect -1858 524 -1800 536
rect -1858 348 -1846 524
rect -1812 348 -1800 524
rect -1858 336 -1800 348
rect -1740 524 -1682 536
rect -1740 348 -1728 524
rect -1694 348 -1682 524
rect -1740 336 -1682 348
rect -1622 524 -1564 536
rect -1622 348 -1610 524
rect -1576 348 -1564 524
rect -1622 336 -1564 348
rect -1504 524 -1446 536
rect -1504 348 -1492 524
rect -1458 348 -1446 524
rect -1504 336 -1446 348
rect -1386 524 -1328 536
rect -1386 348 -1374 524
rect -1340 348 -1328 524
rect -1386 336 -1328 348
rect -1268 524 -1210 536
rect -1268 348 -1256 524
rect -1222 348 -1210 524
rect -1268 336 -1210 348
rect -1150 524 -1092 536
rect -1150 348 -1138 524
rect -1104 348 -1092 524
rect -1150 336 -1092 348
rect -1032 524 -974 536
rect -1032 348 -1020 524
rect -986 348 -974 524
rect -1032 336 -974 348
rect -914 524 -856 536
rect -914 348 -902 524
rect -868 348 -856 524
rect -914 336 -856 348
rect -796 524 -738 536
rect -796 348 -784 524
rect -750 348 -738 524
rect -796 336 -738 348
rect -678 524 -620 536
rect -678 348 -666 524
rect -632 348 -620 524
rect -678 336 -620 348
rect -560 524 -502 536
rect -560 348 -548 524
rect -514 348 -502 524
rect -560 336 -502 348
rect -442 524 -384 536
rect -442 348 -430 524
rect -396 348 -384 524
rect -442 336 -384 348
rect -324 524 -266 536
rect -324 348 -312 524
rect -278 348 -266 524
rect -324 336 -266 348
rect -206 524 -148 536
rect -206 348 -194 524
rect -160 348 -148 524
rect -206 336 -148 348
rect -88 524 -30 536
rect -88 348 -76 524
rect -42 348 -30 524
rect -88 336 -30 348
rect 30 524 88 536
rect 30 348 42 524
rect 76 348 88 524
rect 30 336 88 348
rect 148 524 206 536
rect 148 348 160 524
rect 194 348 206 524
rect 148 336 206 348
rect 266 524 324 536
rect 266 348 278 524
rect 312 348 324 524
rect 266 336 324 348
rect 384 524 442 536
rect 384 348 396 524
rect 430 348 442 524
rect 384 336 442 348
rect 502 524 560 536
rect 502 348 514 524
rect 548 348 560 524
rect 502 336 560 348
rect 620 524 678 536
rect 620 348 632 524
rect 666 348 678 524
rect 620 336 678 348
rect 738 524 796 536
rect 738 348 750 524
rect 784 348 796 524
rect 738 336 796 348
rect 856 524 914 536
rect 856 348 868 524
rect 902 348 914 524
rect 856 336 914 348
rect 974 524 1032 536
rect 974 348 986 524
rect 1020 348 1032 524
rect 974 336 1032 348
rect 1092 524 1150 536
rect 1092 348 1104 524
rect 1138 348 1150 524
rect 1092 336 1150 348
rect 1210 524 1268 536
rect 1210 348 1222 524
rect 1256 348 1268 524
rect 1210 336 1268 348
rect 1328 524 1386 536
rect 1328 348 1340 524
rect 1374 348 1386 524
rect 1328 336 1386 348
rect 1446 524 1504 536
rect 1446 348 1458 524
rect 1492 348 1504 524
rect 1446 336 1504 348
rect 1564 524 1622 536
rect 1564 348 1576 524
rect 1610 348 1622 524
rect 1564 336 1622 348
rect 1682 524 1740 536
rect 1682 348 1694 524
rect 1728 348 1740 524
rect 1682 336 1740 348
rect 1800 524 1858 536
rect 1800 348 1812 524
rect 1846 348 1858 524
rect 1800 336 1858 348
rect 1918 524 1976 536
rect 1918 348 1930 524
rect 1964 348 1976 524
rect 1918 336 1976 348
rect 2036 524 2094 536
rect 2036 348 2048 524
rect 2082 348 2094 524
rect 2036 336 2094 348
rect 2154 524 2212 536
rect 2154 348 2166 524
rect 2200 348 2212 524
rect 2154 336 2212 348
rect 2272 524 2330 536
rect 2272 348 2284 524
rect 2318 348 2330 524
rect 2272 336 2330 348
rect 2390 524 2448 536
rect 2390 348 2402 524
rect 2436 348 2448 524
rect 2390 336 2448 348
rect 2508 524 2566 536
rect 2508 348 2520 524
rect 2554 348 2566 524
rect 2508 336 2566 348
rect 2626 524 2684 536
rect 2626 348 2638 524
rect 2672 348 2684 524
rect 2626 336 2684 348
rect 2744 524 2802 536
rect 2744 348 2756 524
rect 2790 348 2802 524
rect 2744 336 2802 348
rect -2802 88 -2744 100
rect -2802 -88 -2790 88
rect -2756 -88 -2744 88
rect -2802 -100 -2744 -88
rect -2684 88 -2626 100
rect -2684 -88 -2672 88
rect -2638 -88 -2626 88
rect -2684 -100 -2626 -88
rect -2566 88 -2508 100
rect -2566 -88 -2554 88
rect -2520 -88 -2508 88
rect -2566 -100 -2508 -88
rect -2448 88 -2390 100
rect -2448 -88 -2436 88
rect -2402 -88 -2390 88
rect -2448 -100 -2390 -88
rect -2330 88 -2272 100
rect -2330 -88 -2318 88
rect -2284 -88 -2272 88
rect -2330 -100 -2272 -88
rect -2212 88 -2154 100
rect -2212 -88 -2200 88
rect -2166 -88 -2154 88
rect -2212 -100 -2154 -88
rect -2094 88 -2036 100
rect -2094 -88 -2082 88
rect -2048 -88 -2036 88
rect -2094 -100 -2036 -88
rect -1976 88 -1918 100
rect -1976 -88 -1964 88
rect -1930 -88 -1918 88
rect -1976 -100 -1918 -88
rect -1858 88 -1800 100
rect -1858 -88 -1846 88
rect -1812 -88 -1800 88
rect -1858 -100 -1800 -88
rect -1740 88 -1682 100
rect -1740 -88 -1728 88
rect -1694 -88 -1682 88
rect -1740 -100 -1682 -88
rect -1622 88 -1564 100
rect -1622 -88 -1610 88
rect -1576 -88 -1564 88
rect -1622 -100 -1564 -88
rect -1504 88 -1446 100
rect -1504 -88 -1492 88
rect -1458 -88 -1446 88
rect -1504 -100 -1446 -88
rect -1386 88 -1328 100
rect -1386 -88 -1374 88
rect -1340 -88 -1328 88
rect -1386 -100 -1328 -88
rect -1268 88 -1210 100
rect -1268 -88 -1256 88
rect -1222 -88 -1210 88
rect -1268 -100 -1210 -88
rect -1150 88 -1092 100
rect -1150 -88 -1138 88
rect -1104 -88 -1092 88
rect -1150 -100 -1092 -88
rect -1032 88 -974 100
rect -1032 -88 -1020 88
rect -986 -88 -974 88
rect -1032 -100 -974 -88
rect -914 88 -856 100
rect -914 -88 -902 88
rect -868 -88 -856 88
rect -914 -100 -856 -88
rect -796 88 -738 100
rect -796 -88 -784 88
rect -750 -88 -738 88
rect -796 -100 -738 -88
rect -678 88 -620 100
rect -678 -88 -666 88
rect -632 -88 -620 88
rect -678 -100 -620 -88
rect -560 88 -502 100
rect -560 -88 -548 88
rect -514 -88 -502 88
rect -560 -100 -502 -88
rect -442 88 -384 100
rect -442 -88 -430 88
rect -396 -88 -384 88
rect -442 -100 -384 -88
rect -324 88 -266 100
rect -324 -88 -312 88
rect -278 -88 -266 88
rect -324 -100 -266 -88
rect -206 88 -148 100
rect -206 -88 -194 88
rect -160 -88 -148 88
rect -206 -100 -148 -88
rect -88 88 -30 100
rect -88 -88 -76 88
rect -42 -88 -30 88
rect -88 -100 -30 -88
rect 30 88 88 100
rect 30 -88 42 88
rect 76 -88 88 88
rect 30 -100 88 -88
rect 148 88 206 100
rect 148 -88 160 88
rect 194 -88 206 88
rect 148 -100 206 -88
rect 266 88 324 100
rect 266 -88 278 88
rect 312 -88 324 88
rect 266 -100 324 -88
rect 384 88 442 100
rect 384 -88 396 88
rect 430 -88 442 88
rect 384 -100 442 -88
rect 502 88 560 100
rect 502 -88 514 88
rect 548 -88 560 88
rect 502 -100 560 -88
rect 620 88 678 100
rect 620 -88 632 88
rect 666 -88 678 88
rect 620 -100 678 -88
rect 738 88 796 100
rect 738 -88 750 88
rect 784 -88 796 88
rect 738 -100 796 -88
rect 856 88 914 100
rect 856 -88 868 88
rect 902 -88 914 88
rect 856 -100 914 -88
rect 974 88 1032 100
rect 974 -88 986 88
rect 1020 -88 1032 88
rect 974 -100 1032 -88
rect 1092 88 1150 100
rect 1092 -88 1104 88
rect 1138 -88 1150 88
rect 1092 -100 1150 -88
rect 1210 88 1268 100
rect 1210 -88 1222 88
rect 1256 -88 1268 88
rect 1210 -100 1268 -88
rect 1328 88 1386 100
rect 1328 -88 1340 88
rect 1374 -88 1386 88
rect 1328 -100 1386 -88
rect 1446 88 1504 100
rect 1446 -88 1458 88
rect 1492 -88 1504 88
rect 1446 -100 1504 -88
rect 1564 88 1622 100
rect 1564 -88 1576 88
rect 1610 -88 1622 88
rect 1564 -100 1622 -88
rect 1682 88 1740 100
rect 1682 -88 1694 88
rect 1728 -88 1740 88
rect 1682 -100 1740 -88
rect 1800 88 1858 100
rect 1800 -88 1812 88
rect 1846 -88 1858 88
rect 1800 -100 1858 -88
rect 1918 88 1976 100
rect 1918 -88 1930 88
rect 1964 -88 1976 88
rect 1918 -100 1976 -88
rect 2036 88 2094 100
rect 2036 -88 2048 88
rect 2082 -88 2094 88
rect 2036 -100 2094 -88
rect 2154 88 2212 100
rect 2154 -88 2166 88
rect 2200 -88 2212 88
rect 2154 -100 2212 -88
rect 2272 88 2330 100
rect 2272 -88 2284 88
rect 2318 -88 2330 88
rect 2272 -100 2330 -88
rect 2390 88 2448 100
rect 2390 -88 2402 88
rect 2436 -88 2448 88
rect 2390 -100 2448 -88
rect 2508 88 2566 100
rect 2508 -88 2520 88
rect 2554 -88 2566 88
rect 2508 -100 2566 -88
rect 2626 88 2684 100
rect 2626 -88 2638 88
rect 2672 -88 2684 88
rect 2626 -100 2684 -88
rect 2744 88 2802 100
rect 2744 -88 2756 88
rect 2790 -88 2802 88
rect 2744 -100 2802 -88
rect -2802 -348 -2744 -336
rect -2802 -524 -2790 -348
rect -2756 -524 -2744 -348
rect -2802 -536 -2744 -524
rect -2684 -348 -2626 -336
rect -2684 -524 -2672 -348
rect -2638 -524 -2626 -348
rect -2684 -536 -2626 -524
rect -2566 -348 -2508 -336
rect -2566 -524 -2554 -348
rect -2520 -524 -2508 -348
rect -2566 -536 -2508 -524
rect -2448 -348 -2390 -336
rect -2448 -524 -2436 -348
rect -2402 -524 -2390 -348
rect -2448 -536 -2390 -524
rect -2330 -348 -2272 -336
rect -2330 -524 -2318 -348
rect -2284 -524 -2272 -348
rect -2330 -536 -2272 -524
rect -2212 -348 -2154 -336
rect -2212 -524 -2200 -348
rect -2166 -524 -2154 -348
rect -2212 -536 -2154 -524
rect -2094 -348 -2036 -336
rect -2094 -524 -2082 -348
rect -2048 -524 -2036 -348
rect -2094 -536 -2036 -524
rect -1976 -348 -1918 -336
rect -1976 -524 -1964 -348
rect -1930 -524 -1918 -348
rect -1976 -536 -1918 -524
rect -1858 -348 -1800 -336
rect -1858 -524 -1846 -348
rect -1812 -524 -1800 -348
rect -1858 -536 -1800 -524
rect -1740 -348 -1682 -336
rect -1740 -524 -1728 -348
rect -1694 -524 -1682 -348
rect -1740 -536 -1682 -524
rect -1622 -348 -1564 -336
rect -1622 -524 -1610 -348
rect -1576 -524 -1564 -348
rect -1622 -536 -1564 -524
rect -1504 -348 -1446 -336
rect -1504 -524 -1492 -348
rect -1458 -524 -1446 -348
rect -1504 -536 -1446 -524
rect -1386 -348 -1328 -336
rect -1386 -524 -1374 -348
rect -1340 -524 -1328 -348
rect -1386 -536 -1328 -524
rect -1268 -348 -1210 -336
rect -1268 -524 -1256 -348
rect -1222 -524 -1210 -348
rect -1268 -536 -1210 -524
rect -1150 -348 -1092 -336
rect -1150 -524 -1138 -348
rect -1104 -524 -1092 -348
rect -1150 -536 -1092 -524
rect -1032 -348 -974 -336
rect -1032 -524 -1020 -348
rect -986 -524 -974 -348
rect -1032 -536 -974 -524
rect -914 -348 -856 -336
rect -914 -524 -902 -348
rect -868 -524 -856 -348
rect -914 -536 -856 -524
rect -796 -348 -738 -336
rect -796 -524 -784 -348
rect -750 -524 -738 -348
rect -796 -536 -738 -524
rect -678 -348 -620 -336
rect -678 -524 -666 -348
rect -632 -524 -620 -348
rect -678 -536 -620 -524
rect -560 -348 -502 -336
rect -560 -524 -548 -348
rect -514 -524 -502 -348
rect -560 -536 -502 -524
rect -442 -348 -384 -336
rect -442 -524 -430 -348
rect -396 -524 -384 -348
rect -442 -536 -384 -524
rect -324 -348 -266 -336
rect -324 -524 -312 -348
rect -278 -524 -266 -348
rect -324 -536 -266 -524
rect -206 -348 -148 -336
rect -206 -524 -194 -348
rect -160 -524 -148 -348
rect -206 -536 -148 -524
rect -88 -348 -30 -336
rect -88 -524 -76 -348
rect -42 -524 -30 -348
rect -88 -536 -30 -524
rect 30 -348 88 -336
rect 30 -524 42 -348
rect 76 -524 88 -348
rect 30 -536 88 -524
rect 148 -348 206 -336
rect 148 -524 160 -348
rect 194 -524 206 -348
rect 148 -536 206 -524
rect 266 -348 324 -336
rect 266 -524 278 -348
rect 312 -524 324 -348
rect 266 -536 324 -524
rect 384 -348 442 -336
rect 384 -524 396 -348
rect 430 -524 442 -348
rect 384 -536 442 -524
rect 502 -348 560 -336
rect 502 -524 514 -348
rect 548 -524 560 -348
rect 502 -536 560 -524
rect 620 -348 678 -336
rect 620 -524 632 -348
rect 666 -524 678 -348
rect 620 -536 678 -524
rect 738 -348 796 -336
rect 738 -524 750 -348
rect 784 -524 796 -348
rect 738 -536 796 -524
rect 856 -348 914 -336
rect 856 -524 868 -348
rect 902 -524 914 -348
rect 856 -536 914 -524
rect 974 -348 1032 -336
rect 974 -524 986 -348
rect 1020 -524 1032 -348
rect 974 -536 1032 -524
rect 1092 -348 1150 -336
rect 1092 -524 1104 -348
rect 1138 -524 1150 -348
rect 1092 -536 1150 -524
rect 1210 -348 1268 -336
rect 1210 -524 1222 -348
rect 1256 -524 1268 -348
rect 1210 -536 1268 -524
rect 1328 -348 1386 -336
rect 1328 -524 1340 -348
rect 1374 -524 1386 -348
rect 1328 -536 1386 -524
rect 1446 -348 1504 -336
rect 1446 -524 1458 -348
rect 1492 -524 1504 -348
rect 1446 -536 1504 -524
rect 1564 -348 1622 -336
rect 1564 -524 1576 -348
rect 1610 -524 1622 -348
rect 1564 -536 1622 -524
rect 1682 -348 1740 -336
rect 1682 -524 1694 -348
rect 1728 -524 1740 -348
rect 1682 -536 1740 -524
rect 1800 -348 1858 -336
rect 1800 -524 1812 -348
rect 1846 -524 1858 -348
rect 1800 -536 1858 -524
rect 1918 -348 1976 -336
rect 1918 -524 1930 -348
rect 1964 -524 1976 -348
rect 1918 -536 1976 -524
rect 2036 -348 2094 -336
rect 2036 -524 2048 -348
rect 2082 -524 2094 -348
rect 2036 -536 2094 -524
rect 2154 -348 2212 -336
rect 2154 -524 2166 -348
rect 2200 -524 2212 -348
rect 2154 -536 2212 -524
rect 2272 -348 2330 -336
rect 2272 -524 2284 -348
rect 2318 -524 2330 -348
rect 2272 -536 2330 -524
rect 2390 -348 2448 -336
rect 2390 -524 2402 -348
rect 2436 -524 2448 -348
rect 2390 -536 2448 -524
rect 2508 -348 2566 -336
rect 2508 -524 2520 -348
rect 2554 -524 2566 -348
rect 2508 -536 2566 -524
rect 2626 -348 2684 -336
rect 2626 -524 2638 -348
rect 2672 -524 2684 -348
rect 2626 -536 2684 -524
rect 2744 -348 2802 -336
rect 2744 -524 2756 -348
rect 2790 -524 2802 -348
rect 2744 -536 2802 -524
<< pdiffc >>
rect -2790 348 -2756 524
rect -2672 348 -2638 524
rect -2554 348 -2520 524
rect -2436 348 -2402 524
rect -2318 348 -2284 524
rect -2200 348 -2166 524
rect -2082 348 -2048 524
rect -1964 348 -1930 524
rect -1846 348 -1812 524
rect -1728 348 -1694 524
rect -1610 348 -1576 524
rect -1492 348 -1458 524
rect -1374 348 -1340 524
rect -1256 348 -1222 524
rect -1138 348 -1104 524
rect -1020 348 -986 524
rect -902 348 -868 524
rect -784 348 -750 524
rect -666 348 -632 524
rect -548 348 -514 524
rect -430 348 -396 524
rect -312 348 -278 524
rect -194 348 -160 524
rect -76 348 -42 524
rect 42 348 76 524
rect 160 348 194 524
rect 278 348 312 524
rect 396 348 430 524
rect 514 348 548 524
rect 632 348 666 524
rect 750 348 784 524
rect 868 348 902 524
rect 986 348 1020 524
rect 1104 348 1138 524
rect 1222 348 1256 524
rect 1340 348 1374 524
rect 1458 348 1492 524
rect 1576 348 1610 524
rect 1694 348 1728 524
rect 1812 348 1846 524
rect 1930 348 1964 524
rect 2048 348 2082 524
rect 2166 348 2200 524
rect 2284 348 2318 524
rect 2402 348 2436 524
rect 2520 348 2554 524
rect 2638 348 2672 524
rect 2756 348 2790 524
rect -2790 -88 -2756 88
rect -2672 -88 -2638 88
rect -2554 -88 -2520 88
rect -2436 -88 -2402 88
rect -2318 -88 -2284 88
rect -2200 -88 -2166 88
rect -2082 -88 -2048 88
rect -1964 -88 -1930 88
rect -1846 -88 -1812 88
rect -1728 -88 -1694 88
rect -1610 -88 -1576 88
rect -1492 -88 -1458 88
rect -1374 -88 -1340 88
rect -1256 -88 -1222 88
rect -1138 -88 -1104 88
rect -1020 -88 -986 88
rect -902 -88 -868 88
rect -784 -88 -750 88
rect -666 -88 -632 88
rect -548 -88 -514 88
rect -430 -88 -396 88
rect -312 -88 -278 88
rect -194 -88 -160 88
rect -76 -88 -42 88
rect 42 -88 76 88
rect 160 -88 194 88
rect 278 -88 312 88
rect 396 -88 430 88
rect 514 -88 548 88
rect 632 -88 666 88
rect 750 -88 784 88
rect 868 -88 902 88
rect 986 -88 1020 88
rect 1104 -88 1138 88
rect 1222 -88 1256 88
rect 1340 -88 1374 88
rect 1458 -88 1492 88
rect 1576 -88 1610 88
rect 1694 -88 1728 88
rect 1812 -88 1846 88
rect 1930 -88 1964 88
rect 2048 -88 2082 88
rect 2166 -88 2200 88
rect 2284 -88 2318 88
rect 2402 -88 2436 88
rect 2520 -88 2554 88
rect 2638 -88 2672 88
rect 2756 -88 2790 88
rect -2790 -524 -2756 -348
rect -2672 -524 -2638 -348
rect -2554 -524 -2520 -348
rect -2436 -524 -2402 -348
rect -2318 -524 -2284 -348
rect -2200 -524 -2166 -348
rect -2082 -524 -2048 -348
rect -1964 -524 -1930 -348
rect -1846 -524 -1812 -348
rect -1728 -524 -1694 -348
rect -1610 -524 -1576 -348
rect -1492 -524 -1458 -348
rect -1374 -524 -1340 -348
rect -1256 -524 -1222 -348
rect -1138 -524 -1104 -348
rect -1020 -524 -986 -348
rect -902 -524 -868 -348
rect -784 -524 -750 -348
rect -666 -524 -632 -348
rect -548 -524 -514 -348
rect -430 -524 -396 -348
rect -312 -524 -278 -348
rect -194 -524 -160 -348
rect -76 -524 -42 -348
rect 42 -524 76 -348
rect 160 -524 194 -348
rect 278 -524 312 -348
rect 396 -524 430 -348
rect 514 -524 548 -348
rect 632 -524 666 -348
rect 750 -524 784 -348
rect 868 -524 902 -348
rect 986 -524 1020 -348
rect 1104 -524 1138 -348
rect 1222 -524 1256 -348
rect 1340 -524 1374 -348
rect 1458 -524 1492 -348
rect 1576 -524 1610 -348
rect 1694 -524 1728 -348
rect 1812 -524 1846 -348
rect 1930 -524 1964 -348
rect 2048 -524 2082 -348
rect 2166 -524 2200 -348
rect 2284 -524 2318 -348
rect 2402 -524 2436 -348
rect 2520 -524 2554 -348
rect 2638 -524 2672 -348
rect 2756 -524 2790 -348
<< nsubdiff >>
rect -2904 685 -2808 719
rect 2808 685 2904 719
rect -2904 623 -2870 685
rect 2870 623 2904 685
rect -2904 -685 -2870 -623
rect 2870 -685 2904 -623
rect -2904 -719 -2808 -685
rect 2808 -719 2904 -685
<< nsubdiffcont >>
rect -2808 685 2808 719
rect -2904 -623 -2870 623
rect 2870 -623 2904 623
rect -2808 -719 2808 -685
<< poly >>
rect -2747 617 -2681 633
rect -2747 583 -2731 617
rect -2697 583 -2681 617
rect -2747 567 -2681 583
rect -2629 617 -2563 633
rect -2629 583 -2613 617
rect -2579 583 -2563 617
rect -2629 567 -2563 583
rect -2511 617 -2445 633
rect -2511 583 -2495 617
rect -2461 583 -2445 617
rect -2511 567 -2445 583
rect -2393 617 -2327 633
rect -2393 583 -2377 617
rect -2343 583 -2327 617
rect -2393 567 -2327 583
rect -2275 617 -2209 633
rect -2275 583 -2259 617
rect -2225 583 -2209 617
rect -2275 567 -2209 583
rect -2157 617 -2091 633
rect -2157 583 -2141 617
rect -2107 583 -2091 617
rect -2157 567 -2091 583
rect -2039 617 -1973 633
rect -2039 583 -2023 617
rect -1989 583 -1973 617
rect -2039 567 -1973 583
rect -1921 617 -1855 633
rect -1921 583 -1905 617
rect -1871 583 -1855 617
rect -1921 567 -1855 583
rect -1803 617 -1737 633
rect -1803 583 -1787 617
rect -1753 583 -1737 617
rect -1803 567 -1737 583
rect -1685 617 -1619 633
rect -1685 583 -1669 617
rect -1635 583 -1619 617
rect -1685 567 -1619 583
rect -1567 617 -1501 633
rect -1567 583 -1551 617
rect -1517 583 -1501 617
rect -1567 567 -1501 583
rect -1449 617 -1383 633
rect -1449 583 -1433 617
rect -1399 583 -1383 617
rect -1449 567 -1383 583
rect -1331 617 -1265 633
rect -1331 583 -1315 617
rect -1281 583 -1265 617
rect -1331 567 -1265 583
rect -1213 617 -1147 633
rect -1213 583 -1197 617
rect -1163 583 -1147 617
rect -1213 567 -1147 583
rect -1095 617 -1029 633
rect -1095 583 -1079 617
rect -1045 583 -1029 617
rect -1095 567 -1029 583
rect -977 617 -911 633
rect -977 583 -961 617
rect -927 583 -911 617
rect -977 567 -911 583
rect -859 617 -793 633
rect -859 583 -843 617
rect -809 583 -793 617
rect -859 567 -793 583
rect -741 617 -675 633
rect -741 583 -725 617
rect -691 583 -675 617
rect -741 567 -675 583
rect -623 617 -557 633
rect -623 583 -607 617
rect -573 583 -557 617
rect -623 567 -557 583
rect -505 617 -439 633
rect -505 583 -489 617
rect -455 583 -439 617
rect -505 567 -439 583
rect -387 617 -321 633
rect -387 583 -371 617
rect -337 583 -321 617
rect -387 567 -321 583
rect -269 617 -203 633
rect -269 583 -253 617
rect -219 583 -203 617
rect -269 567 -203 583
rect -151 617 -85 633
rect -151 583 -135 617
rect -101 583 -85 617
rect -151 567 -85 583
rect -33 617 33 633
rect -33 583 -17 617
rect 17 583 33 617
rect -33 567 33 583
rect 85 617 151 633
rect 85 583 101 617
rect 135 583 151 617
rect 85 567 151 583
rect 203 617 269 633
rect 203 583 219 617
rect 253 583 269 617
rect 203 567 269 583
rect 321 617 387 633
rect 321 583 337 617
rect 371 583 387 617
rect 321 567 387 583
rect 439 617 505 633
rect 439 583 455 617
rect 489 583 505 617
rect 439 567 505 583
rect 557 617 623 633
rect 557 583 573 617
rect 607 583 623 617
rect 557 567 623 583
rect 675 617 741 633
rect 675 583 691 617
rect 725 583 741 617
rect 675 567 741 583
rect 793 617 859 633
rect 793 583 809 617
rect 843 583 859 617
rect 793 567 859 583
rect 911 617 977 633
rect 911 583 927 617
rect 961 583 977 617
rect 911 567 977 583
rect 1029 617 1095 633
rect 1029 583 1045 617
rect 1079 583 1095 617
rect 1029 567 1095 583
rect 1147 617 1213 633
rect 1147 583 1163 617
rect 1197 583 1213 617
rect 1147 567 1213 583
rect 1265 617 1331 633
rect 1265 583 1281 617
rect 1315 583 1331 617
rect 1265 567 1331 583
rect 1383 617 1449 633
rect 1383 583 1399 617
rect 1433 583 1449 617
rect 1383 567 1449 583
rect 1501 617 1567 633
rect 1501 583 1517 617
rect 1551 583 1567 617
rect 1501 567 1567 583
rect 1619 617 1685 633
rect 1619 583 1635 617
rect 1669 583 1685 617
rect 1619 567 1685 583
rect 1737 617 1803 633
rect 1737 583 1753 617
rect 1787 583 1803 617
rect 1737 567 1803 583
rect 1855 617 1921 633
rect 1855 583 1871 617
rect 1905 583 1921 617
rect 1855 567 1921 583
rect 1973 617 2039 633
rect 1973 583 1989 617
rect 2023 583 2039 617
rect 1973 567 2039 583
rect 2091 617 2157 633
rect 2091 583 2107 617
rect 2141 583 2157 617
rect 2091 567 2157 583
rect 2209 617 2275 633
rect 2209 583 2225 617
rect 2259 583 2275 617
rect 2209 567 2275 583
rect 2327 617 2393 633
rect 2327 583 2343 617
rect 2377 583 2393 617
rect 2327 567 2393 583
rect 2445 617 2511 633
rect 2445 583 2461 617
rect 2495 583 2511 617
rect 2445 567 2511 583
rect 2563 617 2629 633
rect 2563 583 2579 617
rect 2613 583 2629 617
rect 2563 567 2629 583
rect 2681 617 2747 633
rect 2681 583 2697 617
rect 2731 583 2747 617
rect 2681 567 2747 583
rect -2744 536 -2684 567
rect -2626 536 -2566 567
rect -2508 536 -2448 567
rect -2390 536 -2330 567
rect -2272 536 -2212 567
rect -2154 536 -2094 567
rect -2036 536 -1976 567
rect -1918 536 -1858 567
rect -1800 536 -1740 567
rect -1682 536 -1622 567
rect -1564 536 -1504 567
rect -1446 536 -1386 567
rect -1328 536 -1268 567
rect -1210 536 -1150 567
rect -1092 536 -1032 567
rect -974 536 -914 567
rect -856 536 -796 567
rect -738 536 -678 567
rect -620 536 -560 567
rect -502 536 -442 567
rect -384 536 -324 567
rect -266 536 -206 567
rect -148 536 -88 567
rect -30 536 30 567
rect 88 536 148 567
rect 206 536 266 567
rect 324 536 384 567
rect 442 536 502 567
rect 560 536 620 567
rect 678 536 738 567
rect 796 536 856 567
rect 914 536 974 567
rect 1032 536 1092 567
rect 1150 536 1210 567
rect 1268 536 1328 567
rect 1386 536 1446 567
rect 1504 536 1564 567
rect 1622 536 1682 567
rect 1740 536 1800 567
rect 1858 536 1918 567
rect 1976 536 2036 567
rect 2094 536 2154 567
rect 2212 536 2272 567
rect 2330 536 2390 567
rect 2448 536 2508 567
rect 2566 536 2626 567
rect 2684 536 2744 567
rect -2744 305 -2684 336
rect -2626 305 -2566 336
rect -2508 305 -2448 336
rect -2390 305 -2330 336
rect -2272 305 -2212 336
rect -2154 305 -2094 336
rect -2036 305 -1976 336
rect -1918 305 -1858 336
rect -1800 305 -1740 336
rect -1682 305 -1622 336
rect -1564 305 -1504 336
rect -1446 305 -1386 336
rect -1328 305 -1268 336
rect -1210 305 -1150 336
rect -1092 305 -1032 336
rect -974 305 -914 336
rect -856 305 -796 336
rect -738 305 -678 336
rect -620 305 -560 336
rect -502 305 -442 336
rect -384 305 -324 336
rect -266 305 -206 336
rect -148 305 -88 336
rect -30 305 30 336
rect 88 305 148 336
rect 206 305 266 336
rect 324 305 384 336
rect 442 305 502 336
rect 560 305 620 336
rect 678 305 738 336
rect 796 305 856 336
rect 914 305 974 336
rect 1032 305 1092 336
rect 1150 305 1210 336
rect 1268 305 1328 336
rect 1386 305 1446 336
rect 1504 305 1564 336
rect 1622 305 1682 336
rect 1740 305 1800 336
rect 1858 305 1918 336
rect 1976 305 2036 336
rect 2094 305 2154 336
rect 2212 305 2272 336
rect 2330 305 2390 336
rect 2448 305 2508 336
rect 2566 305 2626 336
rect 2684 305 2744 336
rect -2747 289 -2681 305
rect -2747 255 -2731 289
rect -2697 255 -2681 289
rect -2747 239 -2681 255
rect -2629 289 -2563 305
rect -2629 255 -2613 289
rect -2579 255 -2563 289
rect -2629 239 -2563 255
rect -2511 289 -2445 305
rect -2511 255 -2495 289
rect -2461 255 -2445 289
rect -2511 239 -2445 255
rect -2393 289 -2327 305
rect -2393 255 -2377 289
rect -2343 255 -2327 289
rect -2393 239 -2327 255
rect -2275 289 -2209 305
rect -2275 255 -2259 289
rect -2225 255 -2209 289
rect -2275 239 -2209 255
rect -2157 289 -2091 305
rect -2157 255 -2141 289
rect -2107 255 -2091 289
rect -2157 239 -2091 255
rect -2039 289 -1973 305
rect -2039 255 -2023 289
rect -1989 255 -1973 289
rect -2039 239 -1973 255
rect -1921 289 -1855 305
rect -1921 255 -1905 289
rect -1871 255 -1855 289
rect -1921 239 -1855 255
rect -1803 289 -1737 305
rect -1803 255 -1787 289
rect -1753 255 -1737 289
rect -1803 239 -1737 255
rect -1685 289 -1619 305
rect -1685 255 -1669 289
rect -1635 255 -1619 289
rect -1685 239 -1619 255
rect -1567 289 -1501 305
rect -1567 255 -1551 289
rect -1517 255 -1501 289
rect -1567 239 -1501 255
rect -1449 289 -1383 305
rect -1449 255 -1433 289
rect -1399 255 -1383 289
rect -1449 239 -1383 255
rect -1331 289 -1265 305
rect -1331 255 -1315 289
rect -1281 255 -1265 289
rect -1331 239 -1265 255
rect -1213 289 -1147 305
rect -1213 255 -1197 289
rect -1163 255 -1147 289
rect -1213 239 -1147 255
rect -1095 289 -1029 305
rect -1095 255 -1079 289
rect -1045 255 -1029 289
rect -1095 239 -1029 255
rect -977 289 -911 305
rect -977 255 -961 289
rect -927 255 -911 289
rect -977 239 -911 255
rect -859 289 -793 305
rect -859 255 -843 289
rect -809 255 -793 289
rect -859 239 -793 255
rect -741 289 -675 305
rect -741 255 -725 289
rect -691 255 -675 289
rect -741 239 -675 255
rect -623 289 -557 305
rect -623 255 -607 289
rect -573 255 -557 289
rect -623 239 -557 255
rect -505 289 -439 305
rect -505 255 -489 289
rect -455 255 -439 289
rect -505 239 -439 255
rect -387 289 -321 305
rect -387 255 -371 289
rect -337 255 -321 289
rect -387 239 -321 255
rect -269 289 -203 305
rect -269 255 -253 289
rect -219 255 -203 289
rect -269 239 -203 255
rect -151 289 -85 305
rect -151 255 -135 289
rect -101 255 -85 289
rect -151 239 -85 255
rect -33 289 33 305
rect -33 255 -17 289
rect 17 255 33 289
rect -33 239 33 255
rect 85 289 151 305
rect 85 255 101 289
rect 135 255 151 289
rect 85 239 151 255
rect 203 289 269 305
rect 203 255 219 289
rect 253 255 269 289
rect 203 239 269 255
rect 321 289 387 305
rect 321 255 337 289
rect 371 255 387 289
rect 321 239 387 255
rect 439 289 505 305
rect 439 255 455 289
rect 489 255 505 289
rect 439 239 505 255
rect 557 289 623 305
rect 557 255 573 289
rect 607 255 623 289
rect 557 239 623 255
rect 675 289 741 305
rect 675 255 691 289
rect 725 255 741 289
rect 675 239 741 255
rect 793 289 859 305
rect 793 255 809 289
rect 843 255 859 289
rect 793 239 859 255
rect 911 289 977 305
rect 911 255 927 289
rect 961 255 977 289
rect 911 239 977 255
rect 1029 289 1095 305
rect 1029 255 1045 289
rect 1079 255 1095 289
rect 1029 239 1095 255
rect 1147 289 1213 305
rect 1147 255 1163 289
rect 1197 255 1213 289
rect 1147 239 1213 255
rect 1265 289 1331 305
rect 1265 255 1281 289
rect 1315 255 1331 289
rect 1265 239 1331 255
rect 1383 289 1449 305
rect 1383 255 1399 289
rect 1433 255 1449 289
rect 1383 239 1449 255
rect 1501 289 1567 305
rect 1501 255 1517 289
rect 1551 255 1567 289
rect 1501 239 1567 255
rect 1619 289 1685 305
rect 1619 255 1635 289
rect 1669 255 1685 289
rect 1619 239 1685 255
rect 1737 289 1803 305
rect 1737 255 1753 289
rect 1787 255 1803 289
rect 1737 239 1803 255
rect 1855 289 1921 305
rect 1855 255 1871 289
rect 1905 255 1921 289
rect 1855 239 1921 255
rect 1973 289 2039 305
rect 1973 255 1989 289
rect 2023 255 2039 289
rect 1973 239 2039 255
rect 2091 289 2157 305
rect 2091 255 2107 289
rect 2141 255 2157 289
rect 2091 239 2157 255
rect 2209 289 2275 305
rect 2209 255 2225 289
rect 2259 255 2275 289
rect 2209 239 2275 255
rect 2327 289 2393 305
rect 2327 255 2343 289
rect 2377 255 2393 289
rect 2327 239 2393 255
rect 2445 289 2511 305
rect 2445 255 2461 289
rect 2495 255 2511 289
rect 2445 239 2511 255
rect 2563 289 2629 305
rect 2563 255 2579 289
rect 2613 255 2629 289
rect 2563 239 2629 255
rect 2681 289 2747 305
rect 2681 255 2697 289
rect 2731 255 2747 289
rect 2681 239 2747 255
rect -2747 181 -2681 197
rect -2747 147 -2731 181
rect -2697 147 -2681 181
rect -2747 131 -2681 147
rect -2629 181 -2563 197
rect -2629 147 -2613 181
rect -2579 147 -2563 181
rect -2629 131 -2563 147
rect -2511 181 -2445 197
rect -2511 147 -2495 181
rect -2461 147 -2445 181
rect -2511 131 -2445 147
rect -2393 181 -2327 197
rect -2393 147 -2377 181
rect -2343 147 -2327 181
rect -2393 131 -2327 147
rect -2275 181 -2209 197
rect -2275 147 -2259 181
rect -2225 147 -2209 181
rect -2275 131 -2209 147
rect -2157 181 -2091 197
rect -2157 147 -2141 181
rect -2107 147 -2091 181
rect -2157 131 -2091 147
rect -2039 181 -1973 197
rect -2039 147 -2023 181
rect -1989 147 -1973 181
rect -2039 131 -1973 147
rect -1921 181 -1855 197
rect -1921 147 -1905 181
rect -1871 147 -1855 181
rect -1921 131 -1855 147
rect -1803 181 -1737 197
rect -1803 147 -1787 181
rect -1753 147 -1737 181
rect -1803 131 -1737 147
rect -1685 181 -1619 197
rect -1685 147 -1669 181
rect -1635 147 -1619 181
rect -1685 131 -1619 147
rect -1567 181 -1501 197
rect -1567 147 -1551 181
rect -1517 147 -1501 181
rect -1567 131 -1501 147
rect -1449 181 -1383 197
rect -1449 147 -1433 181
rect -1399 147 -1383 181
rect -1449 131 -1383 147
rect -1331 181 -1265 197
rect -1331 147 -1315 181
rect -1281 147 -1265 181
rect -1331 131 -1265 147
rect -1213 181 -1147 197
rect -1213 147 -1197 181
rect -1163 147 -1147 181
rect -1213 131 -1147 147
rect -1095 181 -1029 197
rect -1095 147 -1079 181
rect -1045 147 -1029 181
rect -1095 131 -1029 147
rect -977 181 -911 197
rect -977 147 -961 181
rect -927 147 -911 181
rect -977 131 -911 147
rect -859 181 -793 197
rect -859 147 -843 181
rect -809 147 -793 181
rect -859 131 -793 147
rect -741 181 -675 197
rect -741 147 -725 181
rect -691 147 -675 181
rect -741 131 -675 147
rect -623 181 -557 197
rect -623 147 -607 181
rect -573 147 -557 181
rect -623 131 -557 147
rect -505 181 -439 197
rect -505 147 -489 181
rect -455 147 -439 181
rect -505 131 -439 147
rect -387 181 -321 197
rect -387 147 -371 181
rect -337 147 -321 181
rect -387 131 -321 147
rect -269 181 -203 197
rect -269 147 -253 181
rect -219 147 -203 181
rect -269 131 -203 147
rect -151 181 -85 197
rect -151 147 -135 181
rect -101 147 -85 181
rect -151 131 -85 147
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect 85 181 151 197
rect 85 147 101 181
rect 135 147 151 181
rect 85 131 151 147
rect 203 181 269 197
rect 203 147 219 181
rect 253 147 269 181
rect 203 131 269 147
rect 321 181 387 197
rect 321 147 337 181
rect 371 147 387 181
rect 321 131 387 147
rect 439 181 505 197
rect 439 147 455 181
rect 489 147 505 181
rect 439 131 505 147
rect 557 181 623 197
rect 557 147 573 181
rect 607 147 623 181
rect 557 131 623 147
rect 675 181 741 197
rect 675 147 691 181
rect 725 147 741 181
rect 675 131 741 147
rect 793 181 859 197
rect 793 147 809 181
rect 843 147 859 181
rect 793 131 859 147
rect 911 181 977 197
rect 911 147 927 181
rect 961 147 977 181
rect 911 131 977 147
rect 1029 181 1095 197
rect 1029 147 1045 181
rect 1079 147 1095 181
rect 1029 131 1095 147
rect 1147 181 1213 197
rect 1147 147 1163 181
rect 1197 147 1213 181
rect 1147 131 1213 147
rect 1265 181 1331 197
rect 1265 147 1281 181
rect 1315 147 1331 181
rect 1265 131 1331 147
rect 1383 181 1449 197
rect 1383 147 1399 181
rect 1433 147 1449 181
rect 1383 131 1449 147
rect 1501 181 1567 197
rect 1501 147 1517 181
rect 1551 147 1567 181
rect 1501 131 1567 147
rect 1619 181 1685 197
rect 1619 147 1635 181
rect 1669 147 1685 181
rect 1619 131 1685 147
rect 1737 181 1803 197
rect 1737 147 1753 181
rect 1787 147 1803 181
rect 1737 131 1803 147
rect 1855 181 1921 197
rect 1855 147 1871 181
rect 1905 147 1921 181
rect 1855 131 1921 147
rect 1973 181 2039 197
rect 1973 147 1989 181
rect 2023 147 2039 181
rect 1973 131 2039 147
rect 2091 181 2157 197
rect 2091 147 2107 181
rect 2141 147 2157 181
rect 2091 131 2157 147
rect 2209 181 2275 197
rect 2209 147 2225 181
rect 2259 147 2275 181
rect 2209 131 2275 147
rect 2327 181 2393 197
rect 2327 147 2343 181
rect 2377 147 2393 181
rect 2327 131 2393 147
rect 2445 181 2511 197
rect 2445 147 2461 181
rect 2495 147 2511 181
rect 2445 131 2511 147
rect 2563 181 2629 197
rect 2563 147 2579 181
rect 2613 147 2629 181
rect 2563 131 2629 147
rect 2681 181 2747 197
rect 2681 147 2697 181
rect 2731 147 2747 181
rect 2681 131 2747 147
rect -2744 100 -2684 131
rect -2626 100 -2566 131
rect -2508 100 -2448 131
rect -2390 100 -2330 131
rect -2272 100 -2212 131
rect -2154 100 -2094 131
rect -2036 100 -1976 131
rect -1918 100 -1858 131
rect -1800 100 -1740 131
rect -1682 100 -1622 131
rect -1564 100 -1504 131
rect -1446 100 -1386 131
rect -1328 100 -1268 131
rect -1210 100 -1150 131
rect -1092 100 -1032 131
rect -974 100 -914 131
rect -856 100 -796 131
rect -738 100 -678 131
rect -620 100 -560 131
rect -502 100 -442 131
rect -384 100 -324 131
rect -266 100 -206 131
rect -148 100 -88 131
rect -30 100 30 131
rect 88 100 148 131
rect 206 100 266 131
rect 324 100 384 131
rect 442 100 502 131
rect 560 100 620 131
rect 678 100 738 131
rect 796 100 856 131
rect 914 100 974 131
rect 1032 100 1092 131
rect 1150 100 1210 131
rect 1268 100 1328 131
rect 1386 100 1446 131
rect 1504 100 1564 131
rect 1622 100 1682 131
rect 1740 100 1800 131
rect 1858 100 1918 131
rect 1976 100 2036 131
rect 2094 100 2154 131
rect 2212 100 2272 131
rect 2330 100 2390 131
rect 2448 100 2508 131
rect 2566 100 2626 131
rect 2684 100 2744 131
rect -2744 -131 -2684 -100
rect -2626 -131 -2566 -100
rect -2508 -131 -2448 -100
rect -2390 -131 -2330 -100
rect -2272 -131 -2212 -100
rect -2154 -131 -2094 -100
rect -2036 -131 -1976 -100
rect -1918 -131 -1858 -100
rect -1800 -131 -1740 -100
rect -1682 -131 -1622 -100
rect -1564 -131 -1504 -100
rect -1446 -131 -1386 -100
rect -1328 -131 -1268 -100
rect -1210 -131 -1150 -100
rect -1092 -131 -1032 -100
rect -974 -131 -914 -100
rect -856 -131 -796 -100
rect -738 -131 -678 -100
rect -620 -131 -560 -100
rect -502 -131 -442 -100
rect -384 -131 -324 -100
rect -266 -131 -206 -100
rect -148 -131 -88 -100
rect -30 -131 30 -100
rect 88 -131 148 -100
rect 206 -131 266 -100
rect 324 -131 384 -100
rect 442 -131 502 -100
rect 560 -131 620 -100
rect 678 -131 738 -100
rect 796 -131 856 -100
rect 914 -131 974 -100
rect 1032 -131 1092 -100
rect 1150 -131 1210 -100
rect 1268 -131 1328 -100
rect 1386 -131 1446 -100
rect 1504 -131 1564 -100
rect 1622 -131 1682 -100
rect 1740 -131 1800 -100
rect 1858 -131 1918 -100
rect 1976 -131 2036 -100
rect 2094 -131 2154 -100
rect 2212 -131 2272 -100
rect 2330 -131 2390 -100
rect 2448 -131 2508 -100
rect 2566 -131 2626 -100
rect 2684 -131 2744 -100
rect -2747 -147 -2681 -131
rect -2747 -181 -2731 -147
rect -2697 -181 -2681 -147
rect -2747 -197 -2681 -181
rect -2629 -147 -2563 -131
rect -2629 -181 -2613 -147
rect -2579 -181 -2563 -147
rect -2629 -197 -2563 -181
rect -2511 -147 -2445 -131
rect -2511 -181 -2495 -147
rect -2461 -181 -2445 -147
rect -2511 -197 -2445 -181
rect -2393 -147 -2327 -131
rect -2393 -181 -2377 -147
rect -2343 -181 -2327 -147
rect -2393 -197 -2327 -181
rect -2275 -147 -2209 -131
rect -2275 -181 -2259 -147
rect -2225 -181 -2209 -147
rect -2275 -197 -2209 -181
rect -2157 -147 -2091 -131
rect -2157 -181 -2141 -147
rect -2107 -181 -2091 -147
rect -2157 -197 -2091 -181
rect -2039 -147 -1973 -131
rect -2039 -181 -2023 -147
rect -1989 -181 -1973 -147
rect -2039 -197 -1973 -181
rect -1921 -147 -1855 -131
rect -1921 -181 -1905 -147
rect -1871 -181 -1855 -147
rect -1921 -197 -1855 -181
rect -1803 -147 -1737 -131
rect -1803 -181 -1787 -147
rect -1753 -181 -1737 -147
rect -1803 -197 -1737 -181
rect -1685 -147 -1619 -131
rect -1685 -181 -1669 -147
rect -1635 -181 -1619 -147
rect -1685 -197 -1619 -181
rect -1567 -147 -1501 -131
rect -1567 -181 -1551 -147
rect -1517 -181 -1501 -147
rect -1567 -197 -1501 -181
rect -1449 -147 -1383 -131
rect -1449 -181 -1433 -147
rect -1399 -181 -1383 -147
rect -1449 -197 -1383 -181
rect -1331 -147 -1265 -131
rect -1331 -181 -1315 -147
rect -1281 -181 -1265 -147
rect -1331 -197 -1265 -181
rect -1213 -147 -1147 -131
rect -1213 -181 -1197 -147
rect -1163 -181 -1147 -147
rect -1213 -197 -1147 -181
rect -1095 -147 -1029 -131
rect -1095 -181 -1079 -147
rect -1045 -181 -1029 -147
rect -1095 -197 -1029 -181
rect -977 -147 -911 -131
rect -977 -181 -961 -147
rect -927 -181 -911 -147
rect -977 -197 -911 -181
rect -859 -147 -793 -131
rect -859 -181 -843 -147
rect -809 -181 -793 -147
rect -859 -197 -793 -181
rect -741 -147 -675 -131
rect -741 -181 -725 -147
rect -691 -181 -675 -147
rect -741 -197 -675 -181
rect -623 -147 -557 -131
rect -623 -181 -607 -147
rect -573 -181 -557 -147
rect -623 -197 -557 -181
rect -505 -147 -439 -131
rect -505 -181 -489 -147
rect -455 -181 -439 -147
rect -505 -197 -439 -181
rect -387 -147 -321 -131
rect -387 -181 -371 -147
rect -337 -181 -321 -147
rect -387 -197 -321 -181
rect -269 -147 -203 -131
rect -269 -181 -253 -147
rect -219 -181 -203 -147
rect -269 -197 -203 -181
rect -151 -147 -85 -131
rect -151 -181 -135 -147
rect -101 -181 -85 -147
rect -151 -197 -85 -181
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
rect 85 -147 151 -131
rect 85 -181 101 -147
rect 135 -181 151 -147
rect 85 -197 151 -181
rect 203 -147 269 -131
rect 203 -181 219 -147
rect 253 -181 269 -147
rect 203 -197 269 -181
rect 321 -147 387 -131
rect 321 -181 337 -147
rect 371 -181 387 -147
rect 321 -197 387 -181
rect 439 -147 505 -131
rect 439 -181 455 -147
rect 489 -181 505 -147
rect 439 -197 505 -181
rect 557 -147 623 -131
rect 557 -181 573 -147
rect 607 -181 623 -147
rect 557 -197 623 -181
rect 675 -147 741 -131
rect 675 -181 691 -147
rect 725 -181 741 -147
rect 675 -197 741 -181
rect 793 -147 859 -131
rect 793 -181 809 -147
rect 843 -181 859 -147
rect 793 -197 859 -181
rect 911 -147 977 -131
rect 911 -181 927 -147
rect 961 -181 977 -147
rect 911 -197 977 -181
rect 1029 -147 1095 -131
rect 1029 -181 1045 -147
rect 1079 -181 1095 -147
rect 1029 -197 1095 -181
rect 1147 -147 1213 -131
rect 1147 -181 1163 -147
rect 1197 -181 1213 -147
rect 1147 -197 1213 -181
rect 1265 -147 1331 -131
rect 1265 -181 1281 -147
rect 1315 -181 1331 -147
rect 1265 -197 1331 -181
rect 1383 -147 1449 -131
rect 1383 -181 1399 -147
rect 1433 -181 1449 -147
rect 1383 -197 1449 -181
rect 1501 -147 1567 -131
rect 1501 -181 1517 -147
rect 1551 -181 1567 -147
rect 1501 -197 1567 -181
rect 1619 -147 1685 -131
rect 1619 -181 1635 -147
rect 1669 -181 1685 -147
rect 1619 -197 1685 -181
rect 1737 -147 1803 -131
rect 1737 -181 1753 -147
rect 1787 -181 1803 -147
rect 1737 -197 1803 -181
rect 1855 -147 1921 -131
rect 1855 -181 1871 -147
rect 1905 -181 1921 -147
rect 1855 -197 1921 -181
rect 1973 -147 2039 -131
rect 1973 -181 1989 -147
rect 2023 -181 2039 -147
rect 1973 -197 2039 -181
rect 2091 -147 2157 -131
rect 2091 -181 2107 -147
rect 2141 -181 2157 -147
rect 2091 -197 2157 -181
rect 2209 -147 2275 -131
rect 2209 -181 2225 -147
rect 2259 -181 2275 -147
rect 2209 -197 2275 -181
rect 2327 -147 2393 -131
rect 2327 -181 2343 -147
rect 2377 -181 2393 -147
rect 2327 -197 2393 -181
rect 2445 -147 2511 -131
rect 2445 -181 2461 -147
rect 2495 -181 2511 -147
rect 2445 -197 2511 -181
rect 2563 -147 2629 -131
rect 2563 -181 2579 -147
rect 2613 -181 2629 -147
rect 2563 -197 2629 -181
rect 2681 -147 2747 -131
rect 2681 -181 2697 -147
rect 2731 -181 2747 -147
rect 2681 -197 2747 -181
rect -2747 -255 -2681 -239
rect -2747 -289 -2731 -255
rect -2697 -289 -2681 -255
rect -2747 -305 -2681 -289
rect -2629 -255 -2563 -239
rect -2629 -289 -2613 -255
rect -2579 -289 -2563 -255
rect -2629 -305 -2563 -289
rect -2511 -255 -2445 -239
rect -2511 -289 -2495 -255
rect -2461 -289 -2445 -255
rect -2511 -305 -2445 -289
rect -2393 -255 -2327 -239
rect -2393 -289 -2377 -255
rect -2343 -289 -2327 -255
rect -2393 -305 -2327 -289
rect -2275 -255 -2209 -239
rect -2275 -289 -2259 -255
rect -2225 -289 -2209 -255
rect -2275 -305 -2209 -289
rect -2157 -255 -2091 -239
rect -2157 -289 -2141 -255
rect -2107 -289 -2091 -255
rect -2157 -305 -2091 -289
rect -2039 -255 -1973 -239
rect -2039 -289 -2023 -255
rect -1989 -289 -1973 -255
rect -2039 -305 -1973 -289
rect -1921 -255 -1855 -239
rect -1921 -289 -1905 -255
rect -1871 -289 -1855 -255
rect -1921 -305 -1855 -289
rect -1803 -255 -1737 -239
rect -1803 -289 -1787 -255
rect -1753 -289 -1737 -255
rect -1803 -305 -1737 -289
rect -1685 -255 -1619 -239
rect -1685 -289 -1669 -255
rect -1635 -289 -1619 -255
rect -1685 -305 -1619 -289
rect -1567 -255 -1501 -239
rect -1567 -289 -1551 -255
rect -1517 -289 -1501 -255
rect -1567 -305 -1501 -289
rect -1449 -255 -1383 -239
rect -1449 -289 -1433 -255
rect -1399 -289 -1383 -255
rect -1449 -305 -1383 -289
rect -1331 -255 -1265 -239
rect -1331 -289 -1315 -255
rect -1281 -289 -1265 -255
rect -1331 -305 -1265 -289
rect -1213 -255 -1147 -239
rect -1213 -289 -1197 -255
rect -1163 -289 -1147 -255
rect -1213 -305 -1147 -289
rect -1095 -255 -1029 -239
rect -1095 -289 -1079 -255
rect -1045 -289 -1029 -255
rect -1095 -305 -1029 -289
rect -977 -255 -911 -239
rect -977 -289 -961 -255
rect -927 -289 -911 -255
rect -977 -305 -911 -289
rect -859 -255 -793 -239
rect -859 -289 -843 -255
rect -809 -289 -793 -255
rect -859 -305 -793 -289
rect -741 -255 -675 -239
rect -741 -289 -725 -255
rect -691 -289 -675 -255
rect -741 -305 -675 -289
rect -623 -255 -557 -239
rect -623 -289 -607 -255
rect -573 -289 -557 -255
rect -623 -305 -557 -289
rect -505 -255 -439 -239
rect -505 -289 -489 -255
rect -455 -289 -439 -255
rect -505 -305 -439 -289
rect -387 -255 -321 -239
rect -387 -289 -371 -255
rect -337 -289 -321 -255
rect -387 -305 -321 -289
rect -269 -255 -203 -239
rect -269 -289 -253 -255
rect -219 -289 -203 -255
rect -269 -305 -203 -289
rect -151 -255 -85 -239
rect -151 -289 -135 -255
rect -101 -289 -85 -255
rect -151 -305 -85 -289
rect -33 -255 33 -239
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect -33 -305 33 -289
rect 85 -255 151 -239
rect 85 -289 101 -255
rect 135 -289 151 -255
rect 85 -305 151 -289
rect 203 -255 269 -239
rect 203 -289 219 -255
rect 253 -289 269 -255
rect 203 -305 269 -289
rect 321 -255 387 -239
rect 321 -289 337 -255
rect 371 -289 387 -255
rect 321 -305 387 -289
rect 439 -255 505 -239
rect 439 -289 455 -255
rect 489 -289 505 -255
rect 439 -305 505 -289
rect 557 -255 623 -239
rect 557 -289 573 -255
rect 607 -289 623 -255
rect 557 -305 623 -289
rect 675 -255 741 -239
rect 675 -289 691 -255
rect 725 -289 741 -255
rect 675 -305 741 -289
rect 793 -255 859 -239
rect 793 -289 809 -255
rect 843 -289 859 -255
rect 793 -305 859 -289
rect 911 -255 977 -239
rect 911 -289 927 -255
rect 961 -289 977 -255
rect 911 -305 977 -289
rect 1029 -255 1095 -239
rect 1029 -289 1045 -255
rect 1079 -289 1095 -255
rect 1029 -305 1095 -289
rect 1147 -255 1213 -239
rect 1147 -289 1163 -255
rect 1197 -289 1213 -255
rect 1147 -305 1213 -289
rect 1265 -255 1331 -239
rect 1265 -289 1281 -255
rect 1315 -289 1331 -255
rect 1265 -305 1331 -289
rect 1383 -255 1449 -239
rect 1383 -289 1399 -255
rect 1433 -289 1449 -255
rect 1383 -305 1449 -289
rect 1501 -255 1567 -239
rect 1501 -289 1517 -255
rect 1551 -289 1567 -255
rect 1501 -305 1567 -289
rect 1619 -255 1685 -239
rect 1619 -289 1635 -255
rect 1669 -289 1685 -255
rect 1619 -305 1685 -289
rect 1737 -255 1803 -239
rect 1737 -289 1753 -255
rect 1787 -289 1803 -255
rect 1737 -305 1803 -289
rect 1855 -255 1921 -239
rect 1855 -289 1871 -255
rect 1905 -289 1921 -255
rect 1855 -305 1921 -289
rect 1973 -255 2039 -239
rect 1973 -289 1989 -255
rect 2023 -289 2039 -255
rect 1973 -305 2039 -289
rect 2091 -255 2157 -239
rect 2091 -289 2107 -255
rect 2141 -289 2157 -255
rect 2091 -305 2157 -289
rect 2209 -255 2275 -239
rect 2209 -289 2225 -255
rect 2259 -289 2275 -255
rect 2209 -305 2275 -289
rect 2327 -255 2393 -239
rect 2327 -289 2343 -255
rect 2377 -289 2393 -255
rect 2327 -305 2393 -289
rect 2445 -255 2511 -239
rect 2445 -289 2461 -255
rect 2495 -289 2511 -255
rect 2445 -305 2511 -289
rect 2563 -255 2629 -239
rect 2563 -289 2579 -255
rect 2613 -289 2629 -255
rect 2563 -305 2629 -289
rect 2681 -255 2747 -239
rect 2681 -289 2697 -255
rect 2731 -289 2747 -255
rect 2681 -305 2747 -289
rect -2744 -336 -2684 -305
rect -2626 -336 -2566 -305
rect -2508 -336 -2448 -305
rect -2390 -336 -2330 -305
rect -2272 -336 -2212 -305
rect -2154 -336 -2094 -305
rect -2036 -336 -1976 -305
rect -1918 -336 -1858 -305
rect -1800 -336 -1740 -305
rect -1682 -336 -1622 -305
rect -1564 -336 -1504 -305
rect -1446 -336 -1386 -305
rect -1328 -336 -1268 -305
rect -1210 -336 -1150 -305
rect -1092 -336 -1032 -305
rect -974 -336 -914 -305
rect -856 -336 -796 -305
rect -738 -336 -678 -305
rect -620 -336 -560 -305
rect -502 -336 -442 -305
rect -384 -336 -324 -305
rect -266 -336 -206 -305
rect -148 -336 -88 -305
rect -30 -336 30 -305
rect 88 -336 148 -305
rect 206 -336 266 -305
rect 324 -336 384 -305
rect 442 -336 502 -305
rect 560 -336 620 -305
rect 678 -336 738 -305
rect 796 -336 856 -305
rect 914 -336 974 -305
rect 1032 -336 1092 -305
rect 1150 -336 1210 -305
rect 1268 -336 1328 -305
rect 1386 -336 1446 -305
rect 1504 -336 1564 -305
rect 1622 -336 1682 -305
rect 1740 -336 1800 -305
rect 1858 -336 1918 -305
rect 1976 -336 2036 -305
rect 2094 -336 2154 -305
rect 2212 -336 2272 -305
rect 2330 -336 2390 -305
rect 2448 -336 2508 -305
rect 2566 -336 2626 -305
rect 2684 -336 2744 -305
rect -2744 -567 -2684 -536
rect -2626 -567 -2566 -536
rect -2508 -567 -2448 -536
rect -2390 -567 -2330 -536
rect -2272 -567 -2212 -536
rect -2154 -567 -2094 -536
rect -2036 -567 -1976 -536
rect -1918 -567 -1858 -536
rect -1800 -567 -1740 -536
rect -1682 -567 -1622 -536
rect -1564 -567 -1504 -536
rect -1446 -567 -1386 -536
rect -1328 -567 -1268 -536
rect -1210 -567 -1150 -536
rect -1092 -567 -1032 -536
rect -974 -567 -914 -536
rect -856 -567 -796 -536
rect -738 -567 -678 -536
rect -620 -567 -560 -536
rect -502 -567 -442 -536
rect -384 -567 -324 -536
rect -266 -567 -206 -536
rect -148 -567 -88 -536
rect -30 -567 30 -536
rect 88 -567 148 -536
rect 206 -567 266 -536
rect 324 -567 384 -536
rect 442 -567 502 -536
rect 560 -567 620 -536
rect 678 -567 738 -536
rect 796 -567 856 -536
rect 914 -567 974 -536
rect 1032 -567 1092 -536
rect 1150 -567 1210 -536
rect 1268 -567 1328 -536
rect 1386 -567 1446 -536
rect 1504 -567 1564 -536
rect 1622 -567 1682 -536
rect 1740 -567 1800 -536
rect 1858 -567 1918 -536
rect 1976 -567 2036 -536
rect 2094 -567 2154 -536
rect 2212 -567 2272 -536
rect 2330 -567 2390 -536
rect 2448 -567 2508 -536
rect 2566 -567 2626 -536
rect 2684 -567 2744 -536
rect -2747 -583 -2681 -567
rect -2747 -617 -2731 -583
rect -2697 -617 -2681 -583
rect -2747 -633 -2681 -617
rect -2629 -583 -2563 -567
rect -2629 -617 -2613 -583
rect -2579 -617 -2563 -583
rect -2629 -633 -2563 -617
rect -2511 -583 -2445 -567
rect -2511 -617 -2495 -583
rect -2461 -617 -2445 -583
rect -2511 -633 -2445 -617
rect -2393 -583 -2327 -567
rect -2393 -617 -2377 -583
rect -2343 -617 -2327 -583
rect -2393 -633 -2327 -617
rect -2275 -583 -2209 -567
rect -2275 -617 -2259 -583
rect -2225 -617 -2209 -583
rect -2275 -633 -2209 -617
rect -2157 -583 -2091 -567
rect -2157 -617 -2141 -583
rect -2107 -617 -2091 -583
rect -2157 -633 -2091 -617
rect -2039 -583 -1973 -567
rect -2039 -617 -2023 -583
rect -1989 -617 -1973 -583
rect -2039 -633 -1973 -617
rect -1921 -583 -1855 -567
rect -1921 -617 -1905 -583
rect -1871 -617 -1855 -583
rect -1921 -633 -1855 -617
rect -1803 -583 -1737 -567
rect -1803 -617 -1787 -583
rect -1753 -617 -1737 -583
rect -1803 -633 -1737 -617
rect -1685 -583 -1619 -567
rect -1685 -617 -1669 -583
rect -1635 -617 -1619 -583
rect -1685 -633 -1619 -617
rect -1567 -583 -1501 -567
rect -1567 -617 -1551 -583
rect -1517 -617 -1501 -583
rect -1567 -633 -1501 -617
rect -1449 -583 -1383 -567
rect -1449 -617 -1433 -583
rect -1399 -617 -1383 -583
rect -1449 -633 -1383 -617
rect -1331 -583 -1265 -567
rect -1331 -617 -1315 -583
rect -1281 -617 -1265 -583
rect -1331 -633 -1265 -617
rect -1213 -583 -1147 -567
rect -1213 -617 -1197 -583
rect -1163 -617 -1147 -583
rect -1213 -633 -1147 -617
rect -1095 -583 -1029 -567
rect -1095 -617 -1079 -583
rect -1045 -617 -1029 -583
rect -1095 -633 -1029 -617
rect -977 -583 -911 -567
rect -977 -617 -961 -583
rect -927 -617 -911 -583
rect -977 -633 -911 -617
rect -859 -583 -793 -567
rect -859 -617 -843 -583
rect -809 -617 -793 -583
rect -859 -633 -793 -617
rect -741 -583 -675 -567
rect -741 -617 -725 -583
rect -691 -617 -675 -583
rect -741 -633 -675 -617
rect -623 -583 -557 -567
rect -623 -617 -607 -583
rect -573 -617 -557 -583
rect -623 -633 -557 -617
rect -505 -583 -439 -567
rect -505 -617 -489 -583
rect -455 -617 -439 -583
rect -505 -633 -439 -617
rect -387 -583 -321 -567
rect -387 -617 -371 -583
rect -337 -617 -321 -583
rect -387 -633 -321 -617
rect -269 -583 -203 -567
rect -269 -617 -253 -583
rect -219 -617 -203 -583
rect -269 -633 -203 -617
rect -151 -583 -85 -567
rect -151 -617 -135 -583
rect -101 -617 -85 -583
rect -151 -633 -85 -617
rect -33 -583 33 -567
rect -33 -617 -17 -583
rect 17 -617 33 -583
rect -33 -633 33 -617
rect 85 -583 151 -567
rect 85 -617 101 -583
rect 135 -617 151 -583
rect 85 -633 151 -617
rect 203 -583 269 -567
rect 203 -617 219 -583
rect 253 -617 269 -583
rect 203 -633 269 -617
rect 321 -583 387 -567
rect 321 -617 337 -583
rect 371 -617 387 -583
rect 321 -633 387 -617
rect 439 -583 505 -567
rect 439 -617 455 -583
rect 489 -617 505 -583
rect 439 -633 505 -617
rect 557 -583 623 -567
rect 557 -617 573 -583
rect 607 -617 623 -583
rect 557 -633 623 -617
rect 675 -583 741 -567
rect 675 -617 691 -583
rect 725 -617 741 -583
rect 675 -633 741 -617
rect 793 -583 859 -567
rect 793 -617 809 -583
rect 843 -617 859 -583
rect 793 -633 859 -617
rect 911 -583 977 -567
rect 911 -617 927 -583
rect 961 -617 977 -583
rect 911 -633 977 -617
rect 1029 -583 1095 -567
rect 1029 -617 1045 -583
rect 1079 -617 1095 -583
rect 1029 -633 1095 -617
rect 1147 -583 1213 -567
rect 1147 -617 1163 -583
rect 1197 -617 1213 -583
rect 1147 -633 1213 -617
rect 1265 -583 1331 -567
rect 1265 -617 1281 -583
rect 1315 -617 1331 -583
rect 1265 -633 1331 -617
rect 1383 -583 1449 -567
rect 1383 -617 1399 -583
rect 1433 -617 1449 -583
rect 1383 -633 1449 -617
rect 1501 -583 1567 -567
rect 1501 -617 1517 -583
rect 1551 -617 1567 -583
rect 1501 -633 1567 -617
rect 1619 -583 1685 -567
rect 1619 -617 1635 -583
rect 1669 -617 1685 -583
rect 1619 -633 1685 -617
rect 1737 -583 1803 -567
rect 1737 -617 1753 -583
rect 1787 -617 1803 -583
rect 1737 -633 1803 -617
rect 1855 -583 1921 -567
rect 1855 -617 1871 -583
rect 1905 -617 1921 -583
rect 1855 -633 1921 -617
rect 1973 -583 2039 -567
rect 1973 -617 1989 -583
rect 2023 -617 2039 -583
rect 1973 -633 2039 -617
rect 2091 -583 2157 -567
rect 2091 -617 2107 -583
rect 2141 -617 2157 -583
rect 2091 -633 2157 -617
rect 2209 -583 2275 -567
rect 2209 -617 2225 -583
rect 2259 -617 2275 -583
rect 2209 -633 2275 -617
rect 2327 -583 2393 -567
rect 2327 -617 2343 -583
rect 2377 -617 2393 -583
rect 2327 -633 2393 -617
rect 2445 -583 2511 -567
rect 2445 -617 2461 -583
rect 2495 -617 2511 -583
rect 2445 -633 2511 -617
rect 2563 -583 2629 -567
rect 2563 -617 2579 -583
rect 2613 -617 2629 -583
rect 2563 -633 2629 -617
rect 2681 -583 2747 -567
rect 2681 -617 2697 -583
rect 2731 -617 2747 -583
rect 2681 -633 2747 -617
<< polycont >>
rect -2731 583 -2697 617
rect -2613 583 -2579 617
rect -2495 583 -2461 617
rect -2377 583 -2343 617
rect -2259 583 -2225 617
rect -2141 583 -2107 617
rect -2023 583 -1989 617
rect -1905 583 -1871 617
rect -1787 583 -1753 617
rect -1669 583 -1635 617
rect -1551 583 -1517 617
rect -1433 583 -1399 617
rect -1315 583 -1281 617
rect -1197 583 -1163 617
rect -1079 583 -1045 617
rect -961 583 -927 617
rect -843 583 -809 617
rect -725 583 -691 617
rect -607 583 -573 617
rect -489 583 -455 617
rect -371 583 -337 617
rect -253 583 -219 617
rect -135 583 -101 617
rect -17 583 17 617
rect 101 583 135 617
rect 219 583 253 617
rect 337 583 371 617
rect 455 583 489 617
rect 573 583 607 617
rect 691 583 725 617
rect 809 583 843 617
rect 927 583 961 617
rect 1045 583 1079 617
rect 1163 583 1197 617
rect 1281 583 1315 617
rect 1399 583 1433 617
rect 1517 583 1551 617
rect 1635 583 1669 617
rect 1753 583 1787 617
rect 1871 583 1905 617
rect 1989 583 2023 617
rect 2107 583 2141 617
rect 2225 583 2259 617
rect 2343 583 2377 617
rect 2461 583 2495 617
rect 2579 583 2613 617
rect 2697 583 2731 617
rect -2731 255 -2697 289
rect -2613 255 -2579 289
rect -2495 255 -2461 289
rect -2377 255 -2343 289
rect -2259 255 -2225 289
rect -2141 255 -2107 289
rect -2023 255 -1989 289
rect -1905 255 -1871 289
rect -1787 255 -1753 289
rect -1669 255 -1635 289
rect -1551 255 -1517 289
rect -1433 255 -1399 289
rect -1315 255 -1281 289
rect -1197 255 -1163 289
rect -1079 255 -1045 289
rect -961 255 -927 289
rect -843 255 -809 289
rect -725 255 -691 289
rect -607 255 -573 289
rect -489 255 -455 289
rect -371 255 -337 289
rect -253 255 -219 289
rect -135 255 -101 289
rect -17 255 17 289
rect 101 255 135 289
rect 219 255 253 289
rect 337 255 371 289
rect 455 255 489 289
rect 573 255 607 289
rect 691 255 725 289
rect 809 255 843 289
rect 927 255 961 289
rect 1045 255 1079 289
rect 1163 255 1197 289
rect 1281 255 1315 289
rect 1399 255 1433 289
rect 1517 255 1551 289
rect 1635 255 1669 289
rect 1753 255 1787 289
rect 1871 255 1905 289
rect 1989 255 2023 289
rect 2107 255 2141 289
rect 2225 255 2259 289
rect 2343 255 2377 289
rect 2461 255 2495 289
rect 2579 255 2613 289
rect 2697 255 2731 289
rect -2731 147 -2697 181
rect -2613 147 -2579 181
rect -2495 147 -2461 181
rect -2377 147 -2343 181
rect -2259 147 -2225 181
rect -2141 147 -2107 181
rect -2023 147 -1989 181
rect -1905 147 -1871 181
rect -1787 147 -1753 181
rect -1669 147 -1635 181
rect -1551 147 -1517 181
rect -1433 147 -1399 181
rect -1315 147 -1281 181
rect -1197 147 -1163 181
rect -1079 147 -1045 181
rect -961 147 -927 181
rect -843 147 -809 181
rect -725 147 -691 181
rect -607 147 -573 181
rect -489 147 -455 181
rect -371 147 -337 181
rect -253 147 -219 181
rect -135 147 -101 181
rect -17 147 17 181
rect 101 147 135 181
rect 219 147 253 181
rect 337 147 371 181
rect 455 147 489 181
rect 573 147 607 181
rect 691 147 725 181
rect 809 147 843 181
rect 927 147 961 181
rect 1045 147 1079 181
rect 1163 147 1197 181
rect 1281 147 1315 181
rect 1399 147 1433 181
rect 1517 147 1551 181
rect 1635 147 1669 181
rect 1753 147 1787 181
rect 1871 147 1905 181
rect 1989 147 2023 181
rect 2107 147 2141 181
rect 2225 147 2259 181
rect 2343 147 2377 181
rect 2461 147 2495 181
rect 2579 147 2613 181
rect 2697 147 2731 181
rect -2731 -181 -2697 -147
rect -2613 -181 -2579 -147
rect -2495 -181 -2461 -147
rect -2377 -181 -2343 -147
rect -2259 -181 -2225 -147
rect -2141 -181 -2107 -147
rect -2023 -181 -1989 -147
rect -1905 -181 -1871 -147
rect -1787 -181 -1753 -147
rect -1669 -181 -1635 -147
rect -1551 -181 -1517 -147
rect -1433 -181 -1399 -147
rect -1315 -181 -1281 -147
rect -1197 -181 -1163 -147
rect -1079 -181 -1045 -147
rect -961 -181 -927 -147
rect -843 -181 -809 -147
rect -725 -181 -691 -147
rect -607 -181 -573 -147
rect -489 -181 -455 -147
rect -371 -181 -337 -147
rect -253 -181 -219 -147
rect -135 -181 -101 -147
rect -17 -181 17 -147
rect 101 -181 135 -147
rect 219 -181 253 -147
rect 337 -181 371 -147
rect 455 -181 489 -147
rect 573 -181 607 -147
rect 691 -181 725 -147
rect 809 -181 843 -147
rect 927 -181 961 -147
rect 1045 -181 1079 -147
rect 1163 -181 1197 -147
rect 1281 -181 1315 -147
rect 1399 -181 1433 -147
rect 1517 -181 1551 -147
rect 1635 -181 1669 -147
rect 1753 -181 1787 -147
rect 1871 -181 1905 -147
rect 1989 -181 2023 -147
rect 2107 -181 2141 -147
rect 2225 -181 2259 -147
rect 2343 -181 2377 -147
rect 2461 -181 2495 -147
rect 2579 -181 2613 -147
rect 2697 -181 2731 -147
rect -2731 -289 -2697 -255
rect -2613 -289 -2579 -255
rect -2495 -289 -2461 -255
rect -2377 -289 -2343 -255
rect -2259 -289 -2225 -255
rect -2141 -289 -2107 -255
rect -2023 -289 -1989 -255
rect -1905 -289 -1871 -255
rect -1787 -289 -1753 -255
rect -1669 -289 -1635 -255
rect -1551 -289 -1517 -255
rect -1433 -289 -1399 -255
rect -1315 -289 -1281 -255
rect -1197 -289 -1163 -255
rect -1079 -289 -1045 -255
rect -961 -289 -927 -255
rect -843 -289 -809 -255
rect -725 -289 -691 -255
rect -607 -289 -573 -255
rect -489 -289 -455 -255
rect -371 -289 -337 -255
rect -253 -289 -219 -255
rect -135 -289 -101 -255
rect -17 -289 17 -255
rect 101 -289 135 -255
rect 219 -289 253 -255
rect 337 -289 371 -255
rect 455 -289 489 -255
rect 573 -289 607 -255
rect 691 -289 725 -255
rect 809 -289 843 -255
rect 927 -289 961 -255
rect 1045 -289 1079 -255
rect 1163 -289 1197 -255
rect 1281 -289 1315 -255
rect 1399 -289 1433 -255
rect 1517 -289 1551 -255
rect 1635 -289 1669 -255
rect 1753 -289 1787 -255
rect 1871 -289 1905 -255
rect 1989 -289 2023 -255
rect 2107 -289 2141 -255
rect 2225 -289 2259 -255
rect 2343 -289 2377 -255
rect 2461 -289 2495 -255
rect 2579 -289 2613 -255
rect 2697 -289 2731 -255
rect -2731 -617 -2697 -583
rect -2613 -617 -2579 -583
rect -2495 -617 -2461 -583
rect -2377 -617 -2343 -583
rect -2259 -617 -2225 -583
rect -2141 -617 -2107 -583
rect -2023 -617 -1989 -583
rect -1905 -617 -1871 -583
rect -1787 -617 -1753 -583
rect -1669 -617 -1635 -583
rect -1551 -617 -1517 -583
rect -1433 -617 -1399 -583
rect -1315 -617 -1281 -583
rect -1197 -617 -1163 -583
rect -1079 -617 -1045 -583
rect -961 -617 -927 -583
rect -843 -617 -809 -583
rect -725 -617 -691 -583
rect -607 -617 -573 -583
rect -489 -617 -455 -583
rect -371 -617 -337 -583
rect -253 -617 -219 -583
rect -135 -617 -101 -583
rect -17 -617 17 -583
rect 101 -617 135 -583
rect 219 -617 253 -583
rect 337 -617 371 -583
rect 455 -617 489 -583
rect 573 -617 607 -583
rect 691 -617 725 -583
rect 809 -617 843 -583
rect 927 -617 961 -583
rect 1045 -617 1079 -583
rect 1163 -617 1197 -583
rect 1281 -617 1315 -583
rect 1399 -617 1433 -583
rect 1517 -617 1551 -583
rect 1635 -617 1669 -583
rect 1753 -617 1787 -583
rect 1871 -617 1905 -583
rect 1989 -617 2023 -583
rect 2107 -617 2141 -583
rect 2225 -617 2259 -583
rect 2343 -617 2377 -583
rect 2461 -617 2495 -583
rect 2579 -617 2613 -583
rect 2697 -617 2731 -583
<< locali >>
rect -2904 685 -2808 719
rect 2808 685 2904 719
rect -2904 623 -2870 685
rect 2870 623 2904 685
rect -2747 583 -2731 617
rect -2697 583 -2681 617
rect -2629 583 -2613 617
rect -2579 583 -2563 617
rect -2511 583 -2495 617
rect -2461 583 -2445 617
rect -2393 583 -2377 617
rect -2343 583 -2327 617
rect -2275 583 -2259 617
rect -2225 583 -2209 617
rect -2157 583 -2141 617
rect -2107 583 -2091 617
rect -2039 583 -2023 617
rect -1989 583 -1973 617
rect -1921 583 -1905 617
rect -1871 583 -1855 617
rect -1803 583 -1787 617
rect -1753 583 -1737 617
rect -1685 583 -1669 617
rect -1635 583 -1619 617
rect -1567 583 -1551 617
rect -1517 583 -1501 617
rect -1449 583 -1433 617
rect -1399 583 -1383 617
rect -1331 583 -1315 617
rect -1281 583 -1265 617
rect -1213 583 -1197 617
rect -1163 583 -1147 617
rect -1095 583 -1079 617
rect -1045 583 -1029 617
rect -977 583 -961 617
rect -927 583 -911 617
rect -859 583 -843 617
rect -809 583 -793 617
rect -741 583 -725 617
rect -691 583 -675 617
rect -623 583 -607 617
rect -573 583 -557 617
rect -505 583 -489 617
rect -455 583 -439 617
rect -387 583 -371 617
rect -337 583 -321 617
rect -269 583 -253 617
rect -219 583 -203 617
rect -151 583 -135 617
rect -101 583 -85 617
rect -33 583 -17 617
rect 17 583 33 617
rect 85 583 101 617
rect 135 583 151 617
rect 203 583 219 617
rect 253 583 269 617
rect 321 583 337 617
rect 371 583 387 617
rect 439 583 455 617
rect 489 583 505 617
rect 557 583 573 617
rect 607 583 623 617
rect 675 583 691 617
rect 725 583 741 617
rect 793 583 809 617
rect 843 583 859 617
rect 911 583 927 617
rect 961 583 977 617
rect 1029 583 1045 617
rect 1079 583 1095 617
rect 1147 583 1163 617
rect 1197 583 1213 617
rect 1265 583 1281 617
rect 1315 583 1331 617
rect 1383 583 1399 617
rect 1433 583 1449 617
rect 1501 583 1517 617
rect 1551 583 1567 617
rect 1619 583 1635 617
rect 1669 583 1685 617
rect 1737 583 1753 617
rect 1787 583 1803 617
rect 1855 583 1871 617
rect 1905 583 1921 617
rect 1973 583 1989 617
rect 2023 583 2039 617
rect 2091 583 2107 617
rect 2141 583 2157 617
rect 2209 583 2225 617
rect 2259 583 2275 617
rect 2327 583 2343 617
rect 2377 583 2393 617
rect 2445 583 2461 617
rect 2495 583 2511 617
rect 2563 583 2579 617
rect 2613 583 2629 617
rect 2681 583 2697 617
rect 2731 583 2747 617
rect -2790 524 -2756 540
rect -2790 332 -2756 348
rect -2672 524 -2638 540
rect -2672 332 -2638 348
rect -2554 524 -2520 540
rect -2554 332 -2520 348
rect -2436 524 -2402 540
rect -2436 332 -2402 348
rect -2318 524 -2284 540
rect -2318 332 -2284 348
rect -2200 524 -2166 540
rect -2200 332 -2166 348
rect -2082 524 -2048 540
rect -2082 332 -2048 348
rect -1964 524 -1930 540
rect -1964 332 -1930 348
rect -1846 524 -1812 540
rect -1846 332 -1812 348
rect -1728 524 -1694 540
rect -1728 332 -1694 348
rect -1610 524 -1576 540
rect -1610 332 -1576 348
rect -1492 524 -1458 540
rect -1492 332 -1458 348
rect -1374 524 -1340 540
rect -1374 332 -1340 348
rect -1256 524 -1222 540
rect -1256 332 -1222 348
rect -1138 524 -1104 540
rect -1138 332 -1104 348
rect -1020 524 -986 540
rect -1020 332 -986 348
rect -902 524 -868 540
rect -902 332 -868 348
rect -784 524 -750 540
rect -784 332 -750 348
rect -666 524 -632 540
rect -666 332 -632 348
rect -548 524 -514 540
rect -548 332 -514 348
rect -430 524 -396 540
rect -430 332 -396 348
rect -312 524 -278 540
rect -312 332 -278 348
rect -194 524 -160 540
rect -194 332 -160 348
rect -76 524 -42 540
rect -76 332 -42 348
rect 42 524 76 540
rect 42 332 76 348
rect 160 524 194 540
rect 160 332 194 348
rect 278 524 312 540
rect 278 332 312 348
rect 396 524 430 540
rect 396 332 430 348
rect 514 524 548 540
rect 514 332 548 348
rect 632 524 666 540
rect 632 332 666 348
rect 750 524 784 540
rect 750 332 784 348
rect 868 524 902 540
rect 868 332 902 348
rect 986 524 1020 540
rect 986 332 1020 348
rect 1104 524 1138 540
rect 1104 332 1138 348
rect 1222 524 1256 540
rect 1222 332 1256 348
rect 1340 524 1374 540
rect 1340 332 1374 348
rect 1458 524 1492 540
rect 1458 332 1492 348
rect 1576 524 1610 540
rect 1576 332 1610 348
rect 1694 524 1728 540
rect 1694 332 1728 348
rect 1812 524 1846 540
rect 1812 332 1846 348
rect 1930 524 1964 540
rect 1930 332 1964 348
rect 2048 524 2082 540
rect 2048 332 2082 348
rect 2166 524 2200 540
rect 2166 332 2200 348
rect 2284 524 2318 540
rect 2284 332 2318 348
rect 2402 524 2436 540
rect 2402 332 2436 348
rect 2520 524 2554 540
rect 2520 332 2554 348
rect 2638 524 2672 540
rect 2638 332 2672 348
rect 2756 524 2790 540
rect 2756 332 2790 348
rect -2747 255 -2731 289
rect -2697 255 -2681 289
rect -2629 255 -2613 289
rect -2579 255 -2563 289
rect -2511 255 -2495 289
rect -2461 255 -2445 289
rect -2393 255 -2377 289
rect -2343 255 -2327 289
rect -2275 255 -2259 289
rect -2225 255 -2209 289
rect -2157 255 -2141 289
rect -2107 255 -2091 289
rect -2039 255 -2023 289
rect -1989 255 -1973 289
rect -1921 255 -1905 289
rect -1871 255 -1855 289
rect -1803 255 -1787 289
rect -1753 255 -1737 289
rect -1685 255 -1669 289
rect -1635 255 -1619 289
rect -1567 255 -1551 289
rect -1517 255 -1501 289
rect -1449 255 -1433 289
rect -1399 255 -1383 289
rect -1331 255 -1315 289
rect -1281 255 -1265 289
rect -1213 255 -1197 289
rect -1163 255 -1147 289
rect -1095 255 -1079 289
rect -1045 255 -1029 289
rect -977 255 -961 289
rect -927 255 -911 289
rect -859 255 -843 289
rect -809 255 -793 289
rect -741 255 -725 289
rect -691 255 -675 289
rect -623 255 -607 289
rect -573 255 -557 289
rect -505 255 -489 289
rect -455 255 -439 289
rect -387 255 -371 289
rect -337 255 -321 289
rect -269 255 -253 289
rect -219 255 -203 289
rect -151 255 -135 289
rect -101 255 -85 289
rect -33 255 -17 289
rect 17 255 33 289
rect 85 255 101 289
rect 135 255 151 289
rect 203 255 219 289
rect 253 255 269 289
rect 321 255 337 289
rect 371 255 387 289
rect 439 255 455 289
rect 489 255 505 289
rect 557 255 573 289
rect 607 255 623 289
rect 675 255 691 289
rect 725 255 741 289
rect 793 255 809 289
rect 843 255 859 289
rect 911 255 927 289
rect 961 255 977 289
rect 1029 255 1045 289
rect 1079 255 1095 289
rect 1147 255 1163 289
rect 1197 255 1213 289
rect 1265 255 1281 289
rect 1315 255 1331 289
rect 1383 255 1399 289
rect 1433 255 1449 289
rect 1501 255 1517 289
rect 1551 255 1567 289
rect 1619 255 1635 289
rect 1669 255 1685 289
rect 1737 255 1753 289
rect 1787 255 1803 289
rect 1855 255 1871 289
rect 1905 255 1921 289
rect 1973 255 1989 289
rect 2023 255 2039 289
rect 2091 255 2107 289
rect 2141 255 2157 289
rect 2209 255 2225 289
rect 2259 255 2275 289
rect 2327 255 2343 289
rect 2377 255 2393 289
rect 2445 255 2461 289
rect 2495 255 2511 289
rect 2563 255 2579 289
rect 2613 255 2629 289
rect 2681 255 2697 289
rect 2731 255 2747 289
rect -2747 147 -2731 181
rect -2697 147 -2681 181
rect -2629 147 -2613 181
rect -2579 147 -2563 181
rect -2511 147 -2495 181
rect -2461 147 -2445 181
rect -2393 147 -2377 181
rect -2343 147 -2327 181
rect -2275 147 -2259 181
rect -2225 147 -2209 181
rect -2157 147 -2141 181
rect -2107 147 -2091 181
rect -2039 147 -2023 181
rect -1989 147 -1973 181
rect -1921 147 -1905 181
rect -1871 147 -1855 181
rect -1803 147 -1787 181
rect -1753 147 -1737 181
rect -1685 147 -1669 181
rect -1635 147 -1619 181
rect -1567 147 -1551 181
rect -1517 147 -1501 181
rect -1449 147 -1433 181
rect -1399 147 -1383 181
rect -1331 147 -1315 181
rect -1281 147 -1265 181
rect -1213 147 -1197 181
rect -1163 147 -1147 181
rect -1095 147 -1079 181
rect -1045 147 -1029 181
rect -977 147 -961 181
rect -927 147 -911 181
rect -859 147 -843 181
rect -809 147 -793 181
rect -741 147 -725 181
rect -691 147 -675 181
rect -623 147 -607 181
rect -573 147 -557 181
rect -505 147 -489 181
rect -455 147 -439 181
rect -387 147 -371 181
rect -337 147 -321 181
rect -269 147 -253 181
rect -219 147 -203 181
rect -151 147 -135 181
rect -101 147 -85 181
rect -33 147 -17 181
rect 17 147 33 181
rect 85 147 101 181
rect 135 147 151 181
rect 203 147 219 181
rect 253 147 269 181
rect 321 147 337 181
rect 371 147 387 181
rect 439 147 455 181
rect 489 147 505 181
rect 557 147 573 181
rect 607 147 623 181
rect 675 147 691 181
rect 725 147 741 181
rect 793 147 809 181
rect 843 147 859 181
rect 911 147 927 181
rect 961 147 977 181
rect 1029 147 1045 181
rect 1079 147 1095 181
rect 1147 147 1163 181
rect 1197 147 1213 181
rect 1265 147 1281 181
rect 1315 147 1331 181
rect 1383 147 1399 181
rect 1433 147 1449 181
rect 1501 147 1517 181
rect 1551 147 1567 181
rect 1619 147 1635 181
rect 1669 147 1685 181
rect 1737 147 1753 181
rect 1787 147 1803 181
rect 1855 147 1871 181
rect 1905 147 1921 181
rect 1973 147 1989 181
rect 2023 147 2039 181
rect 2091 147 2107 181
rect 2141 147 2157 181
rect 2209 147 2225 181
rect 2259 147 2275 181
rect 2327 147 2343 181
rect 2377 147 2393 181
rect 2445 147 2461 181
rect 2495 147 2511 181
rect 2563 147 2579 181
rect 2613 147 2629 181
rect 2681 147 2697 181
rect 2731 147 2747 181
rect -2790 88 -2756 104
rect -2790 -104 -2756 -88
rect -2672 88 -2638 104
rect -2672 -104 -2638 -88
rect -2554 88 -2520 104
rect -2554 -104 -2520 -88
rect -2436 88 -2402 104
rect -2436 -104 -2402 -88
rect -2318 88 -2284 104
rect -2318 -104 -2284 -88
rect -2200 88 -2166 104
rect -2200 -104 -2166 -88
rect -2082 88 -2048 104
rect -2082 -104 -2048 -88
rect -1964 88 -1930 104
rect -1964 -104 -1930 -88
rect -1846 88 -1812 104
rect -1846 -104 -1812 -88
rect -1728 88 -1694 104
rect -1728 -104 -1694 -88
rect -1610 88 -1576 104
rect -1610 -104 -1576 -88
rect -1492 88 -1458 104
rect -1492 -104 -1458 -88
rect -1374 88 -1340 104
rect -1374 -104 -1340 -88
rect -1256 88 -1222 104
rect -1256 -104 -1222 -88
rect -1138 88 -1104 104
rect -1138 -104 -1104 -88
rect -1020 88 -986 104
rect -1020 -104 -986 -88
rect -902 88 -868 104
rect -902 -104 -868 -88
rect -784 88 -750 104
rect -784 -104 -750 -88
rect -666 88 -632 104
rect -666 -104 -632 -88
rect -548 88 -514 104
rect -548 -104 -514 -88
rect -430 88 -396 104
rect -430 -104 -396 -88
rect -312 88 -278 104
rect -312 -104 -278 -88
rect -194 88 -160 104
rect -194 -104 -160 -88
rect -76 88 -42 104
rect -76 -104 -42 -88
rect 42 88 76 104
rect 42 -104 76 -88
rect 160 88 194 104
rect 160 -104 194 -88
rect 278 88 312 104
rect 278 -104 312 -88
rect 396 88 430 104
rect 396 -104 430 -88
rect 514 88 548 104
rect 514 -104 548 -88
rect 632 88 666 104
rect 632 -104 666 -88
rect 750 88 784 104
rect 750 -104 784 -88
rect 868 88 902 104
rect 868 -104 902 -88
rect 986 88 1020 104
rect 986 -104 1020 -88
rect 1104 88 1138 104
rect 1104 -104 1138 -88
rect 1222 88 1256 104
rect 1222 -104 1256 -88
rect 1340 88 1374 104
rect 1340 -104 1374 -88
rect 1458 88 1492 104
rect 1458 -104 1492 -88
rect 1576 88 1610 104
rect 1576 -104 1610 -88
rect 1694 88 1728 104
rect 1694 -104 1728 -88
rect 1812 88 1846 104
rect 1812 -104 1846 -88
rect 1930 88 1964 104
rect 1930 -104 1964 -88
rect 2048 88 2082 104
rect 2048 -104 2082 -88
rect 2166 88 2200 104
rect 2166 -104 2200 -88
rect 2284 88 2318 104
rect 2284 -104 2318 -88
rect 2402 88 2436 104
rect 2402 -104 2436 -88
rect 2520 88 2554 104
rect 2520 -104 2554 -88
rect 2638 88 2672 104
rect 2638 -104 2672 -88
rect 2756 88 2790 104
rect 2756 -104 2790 -88
rect -2747 -181 -2731 -147
rect -2697 -181 -2681 -147
rect -2629 -181 -2613 -147
rect -2579 -181 -2563 -147
rect -2511 -181 -2495 -147
rect -2461 -181 -2445 -147
rect -2393 -181 -2377 -147
rect -2343 -181 -2327 -147
rect -2275 -181 -2259 -147
rect -2225 -181 -2209 -147
rect -2157 -181 -2141 -147
rect -2107 -181 -2091 -147
rect -2039 -181 -2023 -147
rect -1989 -181 -1973 -147
rect -1921 -181 -1905 -147
rect -1871 -181 -1855 -147
rect -1803 -181 -1787 -147
rect -1753 -181 -1737 -147
rect -1685 -181 -1669 -147
rect -1635 -181 -1619 -147
rect -1567 -181 -1551 -147
rect -1517 -181 -1501 -147
rect -1449 -181 -1433 -147
rect -1399 -181 -1383 -147
rect -1331 -181 -1315 -147
rect -1281 -181 -1265 -147
rect -1213 -181 -1197 -147
rect -1163 -181 -1147 -147
rect -1095 -181 -1079 -147
rect -1045 -181 -1029 -147
rect -977 -181 -961 -147
rect -927 -181 -911 -147
rect -859 -181 -843 -147
rect -809 -181 -793 -147
rect -741 -181 -725 -147
rect -691 -181 -675 -147
rect -623 -181 -607 -147
rect -573 -181 -557 -147
rect -505 -181 -489 -147
rect -455 -181 -439 -147
rect -387 -181 -371 -147
rect -337 -181 -321 -147
rect -269 -181 -253 -147
rect -219 -181 -203 -147
rect -151 -181 -135 -147
rect -101 -181 -85 -147
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect 85 -181 101 -147
rect 135 -181 151 -147
rect 203 -181 219 -147
rect 253 -181 269 -147
rect 321 -181 337 -147
rect 371 -181 387 -147
rect 439 -181 455 -147
rect 489 -181 505 -147
rect 557 -181 573 -147
rect 607 -181 623 -147
rect 675 -181 691 -147
rect 725 -181 741 -147
rect 793 -181 809 -147
rect 843 -181 859 -147
rect 911 -181 927 -147
rect 961 -181 977 -147
rect 1029 -181 1045 -147
rect 1079 -181 1095 -147
rect 1147 -181 1163 -147
rect 1197 -181 1213 -147
rect 1265 -181 1281 -147
rect 1315 -181 1331 -147
rect 1383 -181 1399 -147
rect 1433 -181 1449 -147
rect 1501 -181 1517 -147
rect 1551 -181 1567 -147
rect 1619 -181 1635 -147
rect 1669 -181 1685 -147
rect 1737 -181 1753 -147
rect 1787 -181 1803 -147
rect 1855 -181 1871 -147
rect 1905 -181 1921 -147
rect 1973 -181 1989 -147
rect 2023 -181 2039 -147
rect 2091 -181 2107 -147
rect 2141 -181 2157 -147
rect 2209 -181 2225 -147
rect 2259 -181 2275 -147
rect 2327 -181 2343 -147
rect 2377 -181 2393 -147
rect 2445 -181 2461 -147
rect 2495 -181 2511 -147
rect 2563 -181 2579 -147
rect 2613 -181 2629 -147
rect 2681 -181 2697 -147
rect 2731 -181 2747 -147
rect -2747 -289 -2731 -255
rect -2697 -289 -2681 -255
rect -2629 -289 -2613 -255
rect -2579 -289 -2563 -255
rect -2511 -289 -2495 -255
rect -2461 -289 -2445 -255
rect -2393 -289 -2377 -255
rect -2343 -289 -2327 -255
rect -2275 -289 -2259 -255
rect -2225 -289 -2209 -255
rect -2157 -289 -2141 -255
rect -2107 -289 -2091 -255
rect -2039 -289 -2023 -255
rect -1989 -289 -1973 -255
rect -1921 -289 -1905 -255
rect -1871 -289 -1855 -255
rect -1803 -289 -1787 -255
rect -1753 -289 -1737 -255
rect -1685 -289 -1669 -255
rect -1635 -289 -1619 -255
rect -1567 -289 -1551 -255
rect -1517 -289 -1501 -255
rect -1449 -289 -1433 -255
rect -1399 -289 -1383 -255
rect -1331 -289 -1315 -255
rect -1281 -289 -1265 -255
rect -1213 -289 -1197 -255
rect -1163 -289 -1147 -255
rect -1095 -289 -1079 -255
rect -1045 -289 -1029 -255
rect -977 -289 -961 -255
rect -927 -289 -911 -255
rect -859 -289 -843 -255
rect -809 -289 -793 -255
rect -741 -289 -725 -255
rect -691 -289 -675 -255
rect -623 -289 -607 -255
rect -573 -289 -557 -255
rect -505 -289 -489 -255
rect -455 -289 -439 -255
rect -387 -289 -371 -255
rect -337 -289 -321 -255
rect -269 -289 -253 -255
rect -219 -289 -203 -255
rect -151 -289 -135 -255
rect -101 -289 -85 -255
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect 85 -289 101 -255
rect 135 -289 151 -255
rect 203 -289 219 -255
rect 253 -289 269 -255
rect 321 -289 337 -255
rect 371 -289 387 -255
rect 439 -289 455 -255
rect 489 -289 505 -255
rect 557 -289 573 -255
rect 607 -289 623 -255
rect 675 -289 691 -255
rect 725 -289 741 -255
rect 793 -289 809 -255
rect 843 -289 859 -255
rect 911 -289 927 -255
rect 961 -289 977 -255
rect 1029 -289 1045 -255
rect 1079 -289 1095 -255
rect 1147 -289 1163 -255
rect 1197 -289 1213 -255
rect 1265 -289 1281 -255
rect 1315 -289 1331 -255
rect 1383 -289 1399 -255
rect 1433 -289 1449 -255
rect 1501 -289 1517 -255
rect 1551 -289 1567 -255
rect 1619 -289 1635 -255
rect 1669 -289 1685 -255
rect 1737 -289 1753 -255
rect 1787 -289 1803 -255
rect 1855 -289 1871 -255
rect 1905 -289 1921 -255
rect 1973 -289 1989 -255
rect 2023 -289 2039 -255
rect 2091 -289 2107 -255
rect 2141 -289 2157 -255
rect 2209 -289 2225 -255
rect 2259 -289 2275 -255
rect 2327 -289 2343 -255
rect 2377 -289 2393 -255
rect 2445 -289 2461 -255
rect 2495 -289 2511 -255
rect 2563 -289 2579 -255
rect 2613 -289 2629 -255
rect 2681 -289 2697 -255
rect 2731 -289 2747 -255
rect -2790 -348 -2756 -332
rect -2790 -540 -2756 -524
rect -2672 -348 -2638 -332
rect -2672 -540 -2638 -524
rect -2554 -348 -2520 -332
rect -2554 -540 -2520 -524
rect -2436 -348 -2402 -332
rect -2436 -540 -2402 -524
rect -2318 -348 -2284 -332
rect -2318 -540 -2284 -524
rect -2200 -348 -2166 -332
rect -2200 -540 -2166 -524
rect -2082 -348 -2048 -332
rect -2082 -540 -2048 -524
rect -1964 -348 -1930 -332
rect -1964 -540 -1930 -524
rect -1846 -348 -1812 -332
rect -1846 -540 -1812 -524
rect -1728 -348 -1694 -332
rect -1728 -540 -1694 -524
rect -1610 -348 -1576 -332
rect -1610 -540 -1576 -524
rect -1492 -348 -1458 -332
rect -1492 -540 -1458 -524
rect -1374 -348 -1340 -332
rect -1374 -540 -1340 -524
rect -1256 -348 -1222 -332
rect -1256 -540 -1222 -524
rect -1138 -348 -1104 -332
rect -1138 -540 -1104 -524
rect -1020 -348 -986 -332
rect -1020 -540 -986 -524
rect -902 -348 -868 -332
rect -902 -540 -868 -524
rect -784 -348 -750 -332
rect -784 -540 -750 -524
rect -666 -348 -632 -332
rect -666 -540 -632 -524
rect -548 -348 -514 -332
rect -548 -540 -514 -524
rect -430 -348 -396 -332
rect -430 -540 -396 -524
rect -312 -348 -278 -332
rect -312 -540 -278 -524
rect -194 -348 -160 -332
rect -194 -540 -160 -524
rect -76 -348 -42 -332
rect -76 -540 -42 -524
rect 42 -348 76 -332
rect 42 -540 76 -524
rect 160 -348 194 -332
rect 160 -540 194 -524
rect 278 -348 312 -332
rect 278 -540 312 -524
rect 396 -348 430 -332
rect 396 -540 430 -524
rect 514 -348 548 -332
rect 514 -540 548 -524
rect 632 -348 666 -332
rect 632 -540 666 -524
rect 750 -348 784 -332
rect 750 -540 784 -524
rect 868 -348 902 -332
rect 868 -540 902 -524
rect 986 -348 1020 -332
rect 986 -540 1020 -524
rect 1104 -348 1138 -332
rect 1104 -540 1138 -524
rect 1222 -348 1256 -332
rect 1222 -540 1256 -524
rect 1340 -348 1374 -332
rect 1340 -540 1374 -524
rect 1458 -348 1492 -332
rect 1458 -540 1492 -524
rect 1576 -348 1610 -332
rect 1576 -540 1610 -524
rect 1694 -348 1728 -332
rect 1694 -540 1728 -524
rect 1812 -348 1846 -332
rect 1812 -540 1846 -524
rect 1930 -348 1964 -332
rect 1930 -540 1964 -524
rect 2048 -348 2082 -332
rect 2048 -540 2082 -524
rect 2166 -348 2200 -332
rect 2166 -540 2200 -524
rect 2284 -348 2318 -332
rect 2284 -540 2318 -524
rect 2402 -348 2436 -332
rect 2402 -540 2436 -524
rect 2520 -348 2554 -332
rect 2520 -540 2554 -524
rect 2638 -348 2672 -332
rect 2638 -540 2672 -524
rect 2756 -348 2790 -332
rect 2756 -540 2790 -524
rect -2747 -617 -2731 -583
rect -2697 -617 -2681 -583
rect -2629 -617 -2613 -583
rect -2579 -617 -2563 -583
rect -2511 -617 -2495 -583
rect -2461 -617 -2445 -583
rect -2393 -617 -2377 -583
rect -2343 -617 -2327 -583
rect -2275 -617 -2259 -583
rect -2225 -617 -2209 -583
rect -2157 -617 -2141 -583
rect -2107 -617 -2091 -583
rect -2039 -617 -2023 -583
rect -1989 -617 -1973 -583
rect -1921 -617 -1905 -583
rect -1871 -617 -1855 -583
rect -1803 -617 -1787 -583
rect -1753 -617 -1737 -583
rect -1685 -617 -1669 -583
rect -1635 -617 -1619 -583
rect -1567 -617 -1551 -583
rect -1517 -617 -1501 -583
rect -1449 -617 -1433 -583
rect -1399 -617 -1383 -583
rect -1331 -617 -1315 -583
rect -1281 -617 -1265 -583
rect -1213 -617 -1197 -583
rect -1163 -617 -1147 -583
rect -1095 -617 -1079 -583
rect -1045 -617 -1029 -583
rect -977 -617 -961 -583
rect -927 -617 -911 -583
rect -859 -617 -843 -583
rect -809 -617 -793 -583
rect -741 -617 -725 -583
rect -691 -617 -675 -583
rect -623 -617 -607 -583
rect -573 -617 -557 -583
rect -505 -617 -489 -583
rect -455 -617 -439 -583
rect -387 -617 -371 -583
rect -337 -617 -321 -583
rect -269 -617 -253 -583
rect -219 -617 -203 -583
rect -151 -617 -135 -583
rect -101 -617 -85 -583
rect -33 -617 -17 -583
rect 17 -617 33 -583
rect 85 -617 101 -583
rect 135 -617 151 -583
rect 203 -617 219 -583
rect 253 -617 269 -583
rect 321 -617 337 -583
rect 371 -617 387 -583
rect 439 -617 455 -583
rect 489 -617 505 -583
rect 557 -617 573 -583
rect 607 -617 623 -583
rect 675 -617 691 -583
rect 725 -617 741 -583
rect 793 -617 809 -583
rect 843 -617 859 -583
rect 911 -617 927 -583
rect 961 -617 977 -583
rect 1029 -617 1045 -583
rect 1079 -617 1095 -583
rect 1147 -617 1163 -583
rect 1197 -617 1213 -583
rect 1265 -617 1281 -583
rect 1315 -617 1331 -583
rect 1383 -617 1399 -583
rect 1433 -617 1449 -583
rect 1501 -617 1517 -583
rect 1551 -617 1567 -583
rect 1619 -617 1635 -583
rect 1669 -617 1685 -583
rect 1737 -617 1753 -583
rect 1787 -617 1803 -583
rect 1855 -617 1871 -583
rect 1905 -617 1921 -583
rect 1973 -617 1989 -583
rect 2023 -617 2039 -583
rect 2091 -617 2107 -583
rect 2141 -617 2157 -583
rect 2209 -617 2225 -583
rect 2259 -617 2275 -583
rect 2327 -617 2343 -583
rect 2377 -617 2393 -583
rect 2445 -617 2461 -583
rect 2495 -617 2511 -583
rect 2563 -617 2579 -583
rect 2613 -617 2629 -583
rect 2681 -617 2697 -583
rect 2731 -617 2747 -583
rect -2904 -685 -2870 -623
rect 2870 -685 2904 -623
rect -2904 -719 -2808 -685
rect 2808 -719 2904 -685
<< viali >>
rect -2731 583 -2697 617
rect -2613 583 -2579 617
rect -2495 583 -2461 617
rect -2377 583 -2343 617
rect -2259 583 -2225 617
rect -2141 583 -2107 617
rect -2023 583 -1989 617
rect -1905 583 -1871 617
rect -1787 583 -1753 617
rect -1669 583 -1635 617
rect -1551 583 -1517 617
rect -1433 583 -1399 617
rect -1315 583 -1281 617
rect -1197 583 -1163 617
rect -1079 583 -1045 617
rect -961 583 -927 617
rect -843 583 -809 617
rect -725 583 -691 617
rect -607 583 -573 617
rect -489 583 -455 617
rect -371 583 -337 617
rect -253 583 -219 617
rect -135 583 -101 617
rect -17 583 17 617
rect 101 583 135 617
rect 219 583 253 617
rect 337 583 371 617
rect 455 583 489 617
rect 573 583 607 617
rect 691 583 725 617
rect 809 583 843 617
rect 927 583 961 617
rect 1045 583 1079 617
rect 1163 583 1197 617
rect 1281 583 1315 617
rect 1399 583 1433 617
rect 1517 583 1551 617
rect 1635 583 1669 617
rect 1753 583 1787 617
rect 1871 583 1905 617
rect 1989 583 2023 617
rect 2107 583 2141 617
rect 2225 583 2259 617
rect 2343 583 2377 617
rect 2461 583 2495 617
rect 2579 583 2613 617
rect 2697 583 2731 617
rect -2790 348 -2756 524
rect -2672 348 -2638 524
rect -2554 348 -2520 524
rect -2436 348 -2402 524
rect -2318 348 -2284 524
rect -2200 348 -2166 524
rect -2082 348 -2048 524
rect -1964 348 -1930 524
rect -1846 348 -1812 524
rect -1728 348 -1694 524
rect -1610 348 -1576 524
rect -1492 348 -1458 524
rect -1374 348 -1340 524
rect -1256 348 -1222 524
rect -1138 348 -1104 524
rect -1020 348 -986 524
rect -902 348 -868 524
rect -784 348 -750 524
rect -666 348 -632 524
rect -548 348 -514 524
rect -430 348 -396 524
rect -312 348 -278 524
rect -194 348 -160 524
rect -76 348 -42 524
rect 42 348 76 524
rect 160 348 194 524
rect 278 348 312 524
rect 396 348 430 524
rect 514 348 548 524
rect 632 348 666 524
rect 750 348 784 524
rect 868 348 902 524
rect 986 348 1020 524
rect 1104 348 1138 524
rect 1222 348 1256 524
rect 1340 348 1374 524
rect 1458 348 1492 524
rect 1576 348 1610 524
rect 1694 348 1728 524
rect 1812 348 1846 524
rect 1930 348 1964 524
rect 2048 348 2082 524
rect 2166 348 2200 524
rect 2284 348 2318 524
rect 2402 348 2436 524
rect 2520 348 2554 524
rect 2638 348 2672 524
rect 2756 348 2790 524
rect -2731 255 -2697 289
rect -2613 255 -2579 289
rect -2495 255 -2461 289
rect -2377 255 -2343 289
rect -2259 255 -2225 289
rect -2141 255 -2107 289
rect -2023 255 -1989 289
rect -1905 255 -1871 289
rect -1787 255 -1753 289
rect -1669 255 -1635 289
rect -1551 255 -1517 289
rect -1433 255 -1399 289
rect -1315 255 -1281 289
rect -1197 255 -1163 289
rect -1079 255 -1045 289
rect -961 255 -927 289
rect -843 255 -809 289
rect -725 255 -691 289
rect -607 255 -573 289
rect -489 255 -455 289
rect -371 255 -337 289
rect -253 255 -219 289
rect -135 255 -101 289
rect -17 255 17 289
rect 101 255 135 289
rect 219 255 253 289
rect 337 255 371 289
rect 455 255 489 289
rect 573 255 607 289
rect 691 255 725 289
rect 809 255 843 289
rect 927 255 961 289
rect 1045 255 1079 289
rect 1163 255 1197 289
rect 1281 255 1315 289
rect 1399 255 1433 289
rect 1517 255 1551 289
rect 1635 255 1669 289
rect 1753 255 1787 289
rect 1871 255 1905 289
rect 1989 255 2023 289
rect 2107 255 2141 289
rect 2225 255 2259 289
rect 2343 255 2377 289
rect 2461 255 2495 289
rect 2579 255 2613 289
rect 2697 255 2731 289
rect -2731 147 -2697 181
rect -2613 147 -2579 181
rect -2495 147 -2461 181
rect -2377 147 -2343 181
rect -2259 147 -2225 181
rect -2141 147 -2107 181
rect -2023 147 -1989 181
rect -1905 147 -1871 181
rect -1787 147 -1753 181
rect -1669 147 -1635 181
rect -1551 147 -1517 181
rect -1433 147 -1399 181
rect -1315 147 -1281 181
rect -1197 147 -1163 181
rect -1079 147 -1045 181
rect -961 147 -927 181
rect -843 147 -809 181
rect -725 147 -691 181
rect -607 147 -573 181
rect -489 147 -455 181
rect -371 147 -337 181
rect -253 147 -219 181
rect -135 147 -101 181
rect -17 147 17 181
rect 101 147 135 181
rect 219 147 253 181
rect 337 147 371 181
rect 455 147 489 181
rect 573 147 607 181
rect 691 147 725 181
rect 809 147 843 181
rect 927 147 961 181
rect 1045 147 1079 181
rect 1163 147 1197 181
rect 1281 147 1315 181
rect 1399 147 1433 181
rect 1517 147 1551 181
rect 1635 147 1669 181
rect 1753 147 1787 181
rect 1871 147 1905 181
rect 1989 147 2023 181
rect 2107 147 2141 181
rect 2225 147 2259 181
rect 2343 147 2377 181
rect 2461 147 2495 181
rect 2579 147 2613 181
rect 2697 147 2731 181
rect -2790 -88 -2756 88
rect -2672 -88 -2638 88
rect -2554 -88 -2520 88
rect -2436 -88 -2402 88
rect -2318 -88 -2284 88
rect -2200 -88 -2166 88
rect -2082 -88 -2048 88
rect -1964 -88 -1930 88
rect -1846 -88 -1812 88
rect -1728 -88 -1694 88
rect -1610 -88 -1576 88
rect -1492 -88 -1458 88
rect -1374 -88 -1340 88
rect -1256 -88 -1222 88
rect -1138 -88 -1104 88
rect -1020 -88 -986 88
rect -902 -88 -868 88
rect -784 -88 -750 88
rect -666 -88 -632 88
rect -548 -88 -514 88
rect -430 -88 -396 88
rect -312 -88 -278 88
rect -194 -88 -160 88
rect -76 -88 -42 88
rect 42 -88 76 88
rect 160 -88 194 88
rect 278 -88 312 88
rect 396 -88 430 88
rect 514 -88 548 88
rect 632 -88 666 88
rect 750 -88 784 88
rect 868 -88 902 88
rect 986 -88 1020 88
rect 1104 -88 1138 88
rect 1222 -88 1256 88
rect 1340 -88 1374 88
rect 1458 -88 1492 88
rect 1576 -88 1610 88
rect 1694 -88 1728 88
rect 1812 -88 1846 88
rect 1930 -88 1964 88
rect 2048 -88 2082 88
rect 2166 -88 2200 88
rect 2284 -88 2318 88
rect 2402 -88 2436 88
rect 2520 -88 2554 88
rect 2638 -88 2672 88
rect 2756 -88 2790 88
rect -2731 -181 -2697 -147
rect -2613 -181 -2579 -147
rect -2495 -181 -2461 -147
rect -2377 -181 -2343 -147
rect -2259 -181 -2225 -147
rect -2141 -181 -2107 -147
rect -2023 -181 -1989 -147
rect -1905 -181 -1871 -147
rect -1787 -181 -1753 -147
rect -1669 -181 -1635 -147
rect -1551 -181 -1517 -147
rect -1433 -181 -1399 -147
rect -1315 -181 -1281 -147
rect -1197 -181 -1163 -147
rect -1079 -181 -1045 -147
rect -961 -181 -927 -147
rect -843 -181 -809 -147
rect -725 -181 -691 -147
rect -607 -181 -573 -147
rect -489 -181 -455 -147
rect -371 -181 -337 -147
rect -253 -181 -219 -147
rect -135 -181 -101 -147
rect -17 -181 17 -147
rect 101 -181 135 -147
rect 219 -181 253 -147
rect 337 -181 371 -147
rect 455 -181 489 -147
rect 573 -181 607 -147
rect 691 -181 725 -147
rect 809 -181 843 -147
rect 927 -181 961 -147
rect 1045 -181 1079 -147
rect 1163 -181 1197 -147
rect 1281 -181 1315 -147
rect 1399 -181 1433 -147
rect 1517 -181 1551 -147
rect 1635 -181 1669 -147
rect 1753 -181 1787 -147
rect 1871 -181 1905 -147
rect 1989 -181 2023 -147
rect 2107 -181 2141 -147
rect 2225 -181 2259 -147
rect 2343 -181 2377 -147
rect 2461 -181 2495 -147
rect 2579 -181 2613 -147
rect 2697 -181 2731 -147
rect -2731 -289 -2697 -255
rect -2613 -289 -2579 -255
rect -2495 -289 -2461 -255
rect -2377 -289 -2343 -255
rect -2259 -289 -2225 -255
rect -2141 -289 -2107 -255
rect -2023 -289 -1989 -255
rect -1905 -289 -1871 -255
rect -1787 -289 -1753 -255
rect -1669 -289 -1635 -255
rect -1551 -289 -1517 -255
rect -1433 -289 -1399 -255
rect -1315 -289 -1281 -255
rect -1197 -289 -1163 -255
rect -1079 -289 -1045 -255
rect -961 -289 -927 -255
rect -843 -289 -809 -255
rect -725 -289 -691 -255
rect -607 -289 -573 -255
rect -489 -289 -455 -255
rect -371 -289 -337 -255
rect -253 -289 -219 -255
rect -135 -289 -101 -255
rect -17 -289 17 -255
rect 101 -289 135 -255
rect 219 -289 253 -255
rect 337 -289 371 -255
rect 455 -289 489 -255
rect 573 -289 607 -255
rect 691 -289 725 -255
rect 809 -289 843 -255
rect 927 -289 961 -255
rect 1045 -289 1079 -255
rect 1163 -289 1197 -255
rect 1281 -289 1315 -255
rect 1399 -289 1433 -255
rect 1517 -289 1551 -255
rect 1635 -289 1669 -255
rect 1753 -289 1787 -255
rect 1871 -289 1905 -255
rect 1989 -289 2023 -255
rect 2107 -289 2141 -255
rect 2225 -289 2259 -255
rect 2343 -289 2377 -255
rect 2461 -289 2495 -255
rect 2579 -289 2613 -255
rect 2697 -289 2731 -255
rect -2790 -524 -2756 -348
rect -2672 -524 -2638 -348
rect -2554 -524 -2520 -348
rect -2436 -524 -2402 -348
rect -2318 -524 -2284 -348
rect -2200 -524 -2166 -348
rect -2082 -524 -2048 -348
rect -1964 -524 -1930 -348
rect -1846 -524 -1812 -348
rect -1728 -524 -1694 -348
rect -1610 -524 -1576 -348
rect -1492 -524 -1458 -348
rect -1374 -524 -1340 -348
rect -1256 -524 -1222 -348
rect -1138 -524 -1104 -348
rect -1020 -524 -986 -348
rect -902 -524 -868 -348
rect -784 -524 -750 -348
rect -666 -524 -632 -348
rect -548 -524 -514 -348
rect -430 -524 -396 -348
rect -312 -524 -278 -348
rect -194 -524 -160 -348
rect -76 -524 -42 -348
rect 42 -524 76 -348
rect 160 -524 194 -348
rect 278 -524 312 -348
rect 396 -524 430 -348
rect 514 -524 548 -348
rect 632 -524 666 -348
rect 750 -524 784 -348
rect 868 -524 902 -348
rect 986 -524 1020 -348
rect 1104 -524 1138 -348
rect 1222 -524 1256 -348
rect 1340 -524 1374 -348
rect 1458 -524 1492 -348
rect 1576 -524 1610 -348
rect 1694 -524 1728 -348
rect 1812 -524 1846 -348
rect 1930 -524 1964 -348
rect 2048 -524 2082 -348
rect 2166 -524 2200 -348
rect 2284 -524 2318 -348
rect 2402 -524 2436 -348
rect 2520 -524 2554 -348
rect 2638 -524 2672 -348
rect 2756 -524 2790 -348
rect -2731 -617 -2697 -583
rect -2613 -617 -2579 -583
rect -2495 -617 -2461 -583
rect -2377 -617 -2343 -583
rect -2259 -617 -2225 -583
rect -2141 -617 -2107 -583
rect -2023 -617 -1989 -583
rect -1905 -617 -1871 -583
rect -1787 -617 -1753 -583
rect -1669 -617 -1635 -583
rect -1551 -617 -1517 -583
rect -1433 -617 -1399 -583
rect -1315 -617 -1281 -583
rect -1197 -617 -1163 -583
rect -1079 -617 -1045 -583
rect -961 -617 -927 -583
rect -843 -617 -809 -583
rect -725 -617 -691 -583
rect -607 -617 -573 -583
rect -489 -617 -455 -583
rect -371 -617 -337 -583
rect -253 -617 -219 -583
rect -135 -617 -101 -583
rect -17 -617 17 -583
rect 101 -617 135 -583
rect 219 -617 253 -583
rect 337 -617 371 -583
rect 455 -617 489 -583
rect 573 -617 607 -583
rect 691 -617 725 -583
rect 809 -617 843 -583
rect 927 -617 961 -583
rect 1045 -617 1079 -583
rect 1163 -617 1197 -583
rect 1281 -617 1315 -583
rect 1399 -617 1433 -583
rect 1517 -617 1551 -583
rect 1635 -617 1669 -583
rect 1753 -617 1787 -583
rect 1871 -617 1905 -583
rect 1989 -617 2023 -583
rect 2107 -617 2141 -583
rect 2225 -617 2259 -583
rect 2343 -617 2377 -583
rect 2461 -617 2495 -583
rect 2579 -617 2613 -583
rect 2697 -617 2731 -583
<< metal1 >>
rect -2743 617 -2685 623
rect -2743 583 -2731 617
rect -2697 583 -2685 617
rect -2743 577 -2685 583
rect -2625 617 -2567 623
rect -2625 583 -2613 617
rect -2579 583 -2567 617
rect -2625 577 -2567 583
rect -2507 617 -2449 623
rect -2507 583 -2495 617
rect -2461 583 -2449 617
rect -2507 577 -2449 583
rect -2389 617 -2331 623
rect -2389 583 -2377 617
rect -2343 583 -2331 617
rect -2389 577 -2331 583
rect -2271 617 -2213 623
rect -2271 583 -2259 617
rect -2225 583 -2213 617
rect -2271 577 -2213 583
rect -2153 617 -2095 623
rect -2153 583 -2141 617
rect -2107 583 -2095 617
rect -2153 577 -2095 583
rect -2035 617 -1977 623
rect -2035 583 -2023 617
rect -1989 583 -1977 617
rect -2035 577 -1977 583
rect -1917 617 -1859 623
rect -1917 583 -1905 617
rect -1871 583 -1859 617
rect -1917 577 -1859 583
rect -1799 617 -1741 623
rect -1799 583 -1787 617
rect -1753 583 -1741 617
rect -1799 577 -1741 583
rect -1681 617 -1623 623
rect -1681 583 -1669 617
rect -1635 583 -1623 617
rect -1681 577 -1623 583
rect -1563 617 -1505 623
rect -1563 583 -1551 617
rect -1517 583 -1505 617
rect -1563 577 -1505 583
rect -1445 617 -1387 623
rect -1445 583 -1433 617
rect -1399 583 -1387 617
rect -1445 577 -1387 583
rect -1327 617 -1269 623
rect -1327 583 -1315 617
rect -1281 583 -1269 617
rect -1327 577 -1269 583
rect -1209 617 -1151 623
rect -1209 583 -1197 617
rect -1163 583 -1151 617
rect -1209 577 -1151 583
rect -1091 617 -1033 623
rect -1091 583 -1079 617
rect -1045 583 -1033 617
rect -1091 577 -1033 583
rect -973 617 -915 623
rect -973 583 -961 617
rect -927 583 -915 617
rect -973 577 -915 583
rect -855 617 -797 623
rect -855 583 -843 617
rect -809 583 -797 617
rect -855 577 -797 583
rect -737 617 -679 623
rect -737 583 -725 617
rect -691 583 -679 617
rect -737 577 -679 583
rect -619 617 -561 623
rect -619 583 -607 617
rect -573 583 -561 617
rect -619 577 -561 583
rect -501 617 -443 623
rect -501 583 -489 617
rect -455 583 -443 617
rect -501 577 -443 583
rect -383 617 -325 623
rect -383 583 -371 617
rect -337 583 -325 617
rect -383 577 -325 583
rect -265 617 -207 623
rect -265 583 -253 617
rect -219 583 -207 617
rect -265 577 -207 583
rect -147 617 -89 623
rect -147 583 -135 617
rect -101 583 -89 617
rect -147 577 -89 583
rect -29 617 29 623
rect -29 583 -17 617
rect 17 583 29 617
rect -29 577 29 583
rect 89 617 147 623
rect 89 583 101 617
rect 135 583 147 617
rect 89 577 147 583
rect 207 617 265 623
rect 207 583 219 617
rect 253 583 265 617
rect 207 577 265 583
rect 325 617 383 623
rect 325 583 337 617
rect 371 583 383 617
rect 325 577 383 583
rect 443 617 501 623
rect 443 583 455 617
rect 489 583 501 617
rect 443 577 501 583
rect 561 617 619 623
rect 561 583 573 617
rect 607 583 619 617
rect 561 577 619 583
rect 679 617 737 623
rect 679 583 691 617
rect 725 583 737 617
rect 679 577 737 583
rect 797 617 855 623
rect 797 583 809 617
rect 843 583 855 617
rect 797 577 855 583
rect 915 617 973 623
rect 915 583 927 617
rect 961 583 973 617
rect 915 577 973 583
rect 1033 617 1091 623
rect 1033 583 1045 617
rect 1079 583 1091 617
rect 1033 577 1091 583
rect 1151 617 1209 623
rect 1151 583 1163 617
rect 1197 583 1209 617
rect 1151 577 1209 583
rect 1269 617 1327 623
rect 1269 583 1281 617
rect 1315 583 1327 617
rect 1269 577 1327 583
rect 1387 617 1445 623
rect 1387 583 1399 617
rect 1433 583 1445 617
rect 1387 577 1445 583
rect 1505 617 1563 623
rect 1505 583 1517 617
rect 1551 583 1563 617
rect 1505 577 1563 583
rect 1623 617 1681 623
rect 1623 583 1635 617
rect 1669 583 1681 617
rect 1623 577 1681 583
rect 1741 617 1799 623
rect 1741 583 1753 617
rect 1787 583 1799 617
rect 1741 577 1799 583
rect 1859 617 1917 623
rect 1859 583 1871 617
rect 1905 583 1917 617
rect 1859 577 1917 583
rect 1977 617 2035 623
rect 1977 583 1989 617
rect 2023 583 2035 617
rect 1977 577 2035 583
rect 2095 617 2153 623
rect 2095 583 2107 617
rect 2141 583 2153 617
rect 2095 577 2153 583
rect 2213 617 2271 623
rect 2213 583 2225 617
rect 2259 583 2271 617
rect 2213 577 2271 583
rect 2331 617 2389 623
rect 2331 583 2343 617
rect 2377 583 2389 617
rect 2331 577 2389 583
rect 2449 617 2507 623
rect 2449 583 2461 617
rect 2495 583 2507 617
rect 2449 577 2507 583
rect 2567 617 2625 623
rect 2567 583 2579 617
rect 2613 583 2625 617
rect 2567 577 2625 583
rect 2685 617 2743 623
rect 2685 583 2697 617
rect 2731 583 2743 617
rect 2685 577 2743 583
rect -2796 524 -2750 536
rect -2796 348 -2790 524
rect -2756 348 -2750 524
rect -2796 336 -2750 348
rect -2678 524 -2632 536
rect -2678 348 -2672 524
rect -2638 348 -2632 524
rect -2678 336 -2632 348
rect -2560 524 -2514 536
rect -2560 348 -2554 524
rect -2520 348 -2514 524
rect -2560 336 -2514 348
rect -2442 524 -2396 536
rect -2442 348 -2436 524
rect -2402 348 -2396 524
rect -2442 336 -2396 348
rect -2324 524 -2278 536
rect -2324 348 -2318 524
rect -2284 348 -2278 524
rect -2324 336 -2278 348
rect -2206 524 -2160 536
rect -2206 348 -2200 524
rect -2166 348 -2160 524
rect -2206 336 -2160 348
rect -2088 524 -2042 536
rect -2088 348 -2082 524
rect -2048 348 -2042 524
rect -2088 336 -2042 348
rect -1970 524 -1924 536
rect -1970 348 -1964 524
rect -1930 348 -1924 524
rect -1970 336 -1924 348
rect -1852 524 -1806 536
rect -1852 348 -1846 524
rect -1812 348 -1806 524
rect -1852 336 -1806 348
rect -1734 524 -1688 536
rect -1734 348 -1728 524
rect -1694 348 -1688 524
rect -1734 336 -1688 348
rect -1616 524 -1570 536
rect -1616 348 -1610 524
rect -1576 348 -1570 524
rect -1616 336 -1570 348
rect -1498 524 -1452 536
rect -1498 348 -1492 524
rect -1458 348 -1452 524
rect -1498 336 -1452 348
rect -1380 524 -1334 536
rect -1380 348 -1374 524
rect -1340 348 -1334 524
rect -1380 336 -1334 348
rect -1262 524 -1216 536
rect -1262 348 -1256 524
rect -1222 348 -1216 524
rect -1262 336 -1216 348
rect -1144 524 -1098 536
rect -1144 348 -1138 524
rect -1104 348 -1098 524
rect -1144 336 -1098 348
rect -1026 524 -980 536
rect -1026 348 -1020 524
rect -986 348 -980 524
rect -1026 336 -980 348
rect -908 524 -862 536
rect -908 348 -902 524
rect -868 348 -862 524
rect -908 336 -862 348
rect -790 524 -744 536
rect -790 348 -784 524
rect -750 348 -744 524
rect -790 336 -744 348
rect -672 524 -626 536
rect -672 348 -666 524
rect -632 348 -626 524
rect -672 336 -626 348
rect -554 524 -508 536
rect -554 348 -548 524
rect -514 348 -508 524
rect -554 336 -508 348
rect -436 524 -390 536
rect -436 348 -430 524
rect -396 348 -390 524
rect -436 336 -390 348
rect -318 524 -272 536
rect -318 348 -312 524
rect -278 348 -272 524
rect -318 336 -272 348
rect -200 524 -154 536
rect -200 348 -194 524
rect -160 348 -154 524
rect -200 336 -154 348
rect -82 524 -36 536
rect -82 348 -76 524
rect -42 348 -36 524
rect -82 336 -36 348
rect 36 524 82 536
rect 36 348 42 524
rect 76 348 82 524
rect 36 336 82 348
rect 154 524 200 536
rect 154 348 160 524
rect 194 348 200 524
rect 154 336 200 348
rect 272 524 318 536
rect 272 348 278 524
rect 312 348 318 524
rect 272 336 318 348
rect 390 524 436 536
rect 390 348 396 524
rect 430 348 436 524
rect 390 336 436 348
rect 508 524 554 536
rect 508 348 514 524
rect 548 348 554 524
rect 508 336 554 348
rect 626 524 672 536
rect 626 348 632 524
rect 666 348 672 524
rect 626 336 672 348
rect 744 524 790 536
rect 744 348 750 524
rect 784 348 790 524
rect 744 336 790 348
rect 862 524 908 536
rect 862 348 868 524
rect 902 348 908 524
rect 862 336 908 348
rect 980 524 1026 536
rect 980 348 986 524
rect 1020 348 1026 524
rect 980 336 1026 348
rect 1098 524 1144 536
rect 1098 348 1104 524
rect 1138 348 1144 524
rect 1098 336 1144 348
rect 1216 524 1262 536
rect 1216 348 1222 524
rect 1256 348 1262 524
rect 1216 336 1262 348
rect 1334 524 1380 536
rect 1334 348 1340 524
rect 1374 348 1380 524
rect 1334 336 1380 348
rect 1452 524 1498 536
rect 1452 348 1458 524
rect 1492 348 1498 524
rect 1452 336 1498 348
rect 1570 524 1616 536
rect 1570 348 1576 524
rect 1610 348 1616 524
rect 1570 336 1616 348
rect 1688 524 1734 536
rect 1688 348 1694 524
rect 1728 348 1734 524
rect 1688 336 1734 348
rect 1806 524 1852 536
rect 1806 348 1812 524
rect 1846 348 1852 524
rect 1806 336 1852 348
rect 1924 524 1970 536
rect 1924 348 1930 524
rect 1964 348 1970 524
rect 1924 336 1970 348
rect 2042 524 2088 536
rect 2042 348 2048 524
rect 2082 348 2088 524
rect 2042 336 2088 348
rect 2160 524 2206 536
rect 2160 348 2166 524
rect 2200 348 2206 524
rect 2160 336 2206 348
rect 2278 524 2324 536
rect 2278 348 2284 524
rect 2318 348 2324 524
rect 2278 336 2324 348
rect 2396 524 2442 536
rect 2396 348 2402 524
rect 2436 348 2442 524
rect 2396 336 2442 348
rect 2514 524 2560 536
rect 2514 348 2520 524
rect 2554 348 2560 524
rect 2514 336 2560 348
rect 2632 524 2678 536
rect 2632 348 2638 524
rect 2672 348 2678 524
rect 2632 336 2678 348
rect 2750 524 2796 536
rect 2750 348 2756 524
rect 2790 348 2796 524
rect 2750 336 2796 348
rect -2743 289 -2685 295
rect -2743 255 -2731 289
rect -2697 255 -2685 289
rect -2743 249 -2685 255
rect -2625 289 -2567 295
rect -2625 255 -2613 289
rect -2579 255 -2567 289
rect -2625 249 -2567 255
rect -2507 289 -2449 295
rect -2507 255 -2495 289
rect -2461 255 -2449 289
rect -2507 249 -2449 255
rect -2389 289 -2331 295
rect -2389 255 -2377 289
rect -2343 255 -2331 289
rect -2389 249 -2331 255
rect -2271 289 -2213 295
rect -2271 255 -2259 289
rect -2225 255 -2213 289
rect -2271 249 -2213 255
rect -2153 289 -2095 295
rect -2153 255 -2141 289
rect -2107 255 -2095 289
rect -2153 249 -2095 255
rect -2035 289 -1977 295
rect -2035 255 -2023 289
rect -1989 255 -1977 289
rect -2035 249 -1977 255
rect -1917 289 -1859 295
rect -1917 255 -1905 289
rect -1871 255 -1859 289
rect -1917 249 -1859 255
rect -1799 289 -1741 295
rect -1799 255 -1787 289
rect -1753 255 -1741 289
rect -1799 249 -1741 255
rect -1681 289 -1623 295
rect -1681 255 -1669 289
rect -1635 255 -1623 289
rect -1681 249 -1623 255
rect -1563 289 -1505 295
rect -1563 255 -1551 289
rect -1517 255 -1505 289
rect -1563 249 -1505 255
rect -1445 289 -1387 295
rect -1445 255 -1433 289
rect -1399 255 -1387 289
rect -1445 249 -1387 255
rect -1327 289 -1269 295
rect -1327 255 -1315 289
rect -1281 255 -1269 289
rect -1327 249 -1269 255
rect -1209 289 -1151 295
rect -1209 255 -1197 289
rect -1163 255 -1151 289
rect -1209 249 -1151 255
rect -1091 289 -1033 295
rect -1091 255 -1079 289
rect -1045 255 -1033 289
rect -1091 249 -1033 255
rect -973 289 -915 295
rect -973 255 -961 289
rect -927 255 -915 289
rect -973 249 -915 255
rect -855 289 -797 295
rect -855 255 -843 289
rect -809 255 -797 289
rect -855 249 -797 255
rect -737 289 -679 295
rect -737 255 -725 289
rect -691 255 -679 289
rect -737 249 -679 255
rect -619 289 -561 295
rect -619 255 -607 289
rect -573 255 -561 289
rect -619 249 -561 255
rect -501 289 -443 295
rect -501 255 -489 289
rect -455 255 -443 289
rect -501 249 -443 255
rect -383 289 -325 295
rect -383 255 -371 289
rect -337 255 -325 289
rect -383 249 -325 255
rect -265 289 -207 295
rect -265 255 -253 289
rect -219 255 -207 289
rect -265 249 -207 255
rect -147 289 -89 295
rect -147 255 -135 289
rect -101 255 -89 289
rect -147 249 -89 255
rect -29 289 29 295
rect -29 255 -17 289
rect 17 255 29 289
rect -29 249 29 255
rect 89 289 147 295
rect 89 255 101 289
rect 135 255 147 289
rect 89 249 147 255
rect 207 289 265 295
rect 207 255 219 289
rect 253 255 265 289
rect 207 249 265 255
rect 325 289 383 295
rect 325 255 337 289
rect 371 255 383 289
rect 325 249 383 255
rect 443 289 501 295
rect 443 255 455 289
rect 489 255 501 289
rect 443 249 501 255
rect 561 289 619 295
rect 561 255 573 289
rect 607 255 619 289
rect 561 249 619 255
rect 679 289 737 295
rect 679 255 691 289
rect 725 255 737 289
rect 679 249 737 255
rect 797 289 855 295
rect 797 255 809 289
rect 843 255 855 289
rect 797 249 855 255
rect 915 289 973 295
rect 915 255 927 289
rect 961 255 973 289
rect 915 249 973 255
rect 1033 289 1091 295
rect 1033 255 1045 289
rect 1079 255 1091 289
rect 1033 249 1091 255
rect 1151 289 1209 295
rect 1151 255 1163 289
rect 1197 255 1209 289
rect 1151 249 1209 255
rect 1269 289 1327 295
rect 1269 255 1281 289
rect 1315 255 1327 289
rect 1269 249 1327 255
rect 1387 289 1445 295
rect 1387 255 1399 289
rect 1433 255 1445 289
rect 1387 249 1445 255
rect 1505 289 1563 295
rect 1505 255 1517 289
rect 1551 255 1563 289
rect 1505 249 1563 255
rect 1623 289 1681 295
rect 1623 255 1635 289
rect 1669 255 1681 289
rect 1623 249 1681 255
rect 1741 289 1799 295
rect 1741 255 1753 289
rect 1787 255 1799 289
rect 1741 249 1799 255
rect 1859 289 1917 295
rect 1859 255 1871 289
rect 1905 255 1917 289
rect 1859 249 1917 255
rect 1977 289 2035 295
rect 1977 255 1989 289
rect 2023 255 2035 289
rect 1977 249 2035 255
rect 2095 289 2153 295
rect 2095 255 2107 289
rect 2141 255 2153 289
rect 2095 249 2153 255
rect 2213 289 2271 295
rect 2213 255 2225 289
rect 2259 255 2271 289
rect 2213 249 2271 255
rect 2331 289 2389 295
rect 2331 255 2343 289
rect 2377 255 2389 289
rect 2331 249 2389 255
rect 2449 289 2507 295
rect 2449 255 2461 289
rect 2495 255 2507 289
rect 2449 249 2507 255
rect 2567 289 2625 295
rect 2567 255 2579 289
rect 2613 255 2625 289
rect 2567 249 2625 255
rect 2685 289 2743 295
rect 2685 255 2697 289
rect 2731 255 2743 289
rect 2685 249 2743 255
rect -2743 181 -2685 187
rect -2743 147 -2731 181
rect -2697 147 -2685 181
rect -2743 141 -2685 147
rect -2625 181 -2567 187
rect -2625 147 -2613 181
rect -2579 147 -2567 181
rect -2625 141 -2567 147
rect -2507 181 -2449 187
rect -2507 147 -2495 181
rect -2461 147 -2449 181
rect -2507 141 -2449 147
rect -2389 181 -2331 187
rect -2389 147 -2377 181
rect -2343 147 -2331 181
rect -2389 141 -2331 147
rect -2271 181 -2213 187
rect -2271 147 -2259 181
rect -2225 147 -2213 181
rect -2271 141 -2213 147
rect -2153 181 -2095 187
rect -2153 147 -2141 181
rect -2107 147 -2095 181
rect -2153 141 -2095 147
rect -2035 181 -1977 187
rect -2035 147 -2023 181
rect -1989 147 -1977 181
rect -2035 141 -1977 147
rect -1917 181 -1859 187
rect -1917 147 -1905 181
rect -1871 147 -1859 181
rect -1917 141 -1859 147
rect -1799 181 -1741 187
rect -1799 147 -1787 181
rect -1753 147 -1741 181
rect -1799 141 -1741 147
rect -1681 181 -1623 187
rect -1681 147 -1669 181
rect -1635 147 -1623 181
rect -1681 141 -1623 147
rect -1563 181 -1505 187
rect -1563 147 -1551 181
rect -1517 147 -1505 181
rect -1563 141 -1505 147
rect -1445 181 -1387 187
rect -1445 147 -1433 181
rect -1399 147 -1387 181
rect -1445 141 -1387 147
rect -1327 181 -1269 187
rect -1327 147 -1315 181
rect -1281 147 -1269 181
rect -1327 141 -1269 147
rect -1209 181 -1151 187
rect -1209 147 -1197 181
rect -1163 147 -1151 181
rect -1209 141 -1151 147
rect -1091 181 -1033 187
rect -1091 147 -1079 181
rect -1045 147 -1033 181
rect -1091 141 -1033 147
rect -973 181 -915 187
rect -973 147 -961 181
rect -927 147 -915 181
rect -973 141 -915 147
rect -855 181 -797 187
rect -855 147 -843 181
rect -809 147 -797 181
rect -855 141 -797 147
rect -737 181 -679 187
rect -737 147 -725 181
rect -691 147 -679 181
rect -737 141 -679 147
rect -619 181 -561 187
rect -619 147 -607 181
rect -573 147 -561 181
rect -619 141 -561 147
rect -501 181 -443 187
rect -501 147 -489 181
rect -455 147 -443 181
rect -501 141 -443 147
rect -383 181 -325 187
rect -383 147 -371 181
rect -337 147 -325 181
rect -383 141 -325 147
rect -265 181 -207 187
rect -265 147 -253 181
rect -219 147 -207 181
rect -265 141 -207 147
rect -147 181 -89 187
rect -147 147 -135 181
rect -101 147 -89 181
rect -147 141 -89 147
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect 89 181 147 187
rect 89 147 101 181
rect 135 147 147 181
rect 89 141 147 147
rect 207 181 265 187
rect 207 147 219 181
rect 253 147 265 181
rect 207 141 265 147
rect 325 181 383 187
rect 325 147 337 181
rect 371 147 383 181
rect 325 141 383 147
rect 443 181 501 187
rect 443 147 455 181
rect 489 147 501 181
rect 443 141 501 147
rect 561 181 619 187
rect 561 147 573 181
rect 607 147 619 181
rect 561 141 619 147
rect 679 181 737 187
rect 679 147 691 181
rect 725 147 737 181
rect 679 141 737 147
rect 797 181 855 187
rect 797 147 809 181
rect 843 147 855 181
rect 797 141 855 147
rect 915 181 973 187
rect 915 147 927 181
rect 961 147 973 181
rect 915 141 973 147
rect 1033 181 1091 187
rect 1033 147 1045 181
rect 1079 147 1091 181
rect 1033 141 1091 147
rect 1151 181 1209 187
rect 1151 147 1163 181
rect 1197 147 1209 181
rect 1151 141 1209 147
rect 1269 181 1327 187
rect 1269 147 1281 181
rect 1315 147 1327 181
rect 1269 141 1327 147
rect 1387 181 1445 187
rect 1387 147 1399 181
rect 1433 147 1445 181
rect 1387 141 1445 147
rect 1505 181 1563 187
rect 1505 147 1517 181
rect 1551 147 1563 181
rect 1505 141 1563 147
rect 1623 181 1681 187
rect 1623 147 1635 181
rect 1669 147 1681 181
rect 1623 141 1681 147
rect 1741 181 1799 187
rect 1741 147 1753 181
rect 1787 147 1799 181
rect 1741 141 1799 147
rect 1859 181 1917 187
rect 1859 147 1871 181
rect 1905 147 1917 181
rect 1859 141 1917 147
rect 1977 181 2035 187
rect 1977 147 1989 181
rect 2023 147 2035 181
rect 1977 141 2035 147
rect 2095 181 2153 187
rect 2095 147 2107 181
rect 2141 147 2153 181
rect 2095 141 2153 147
rect 2213 181 2271 187
rect 2213 147 2225 181
rect 2259 147 2271 181
rect 2213 141 2271 147
rect 2331 181 2389 187
rect 2331 147 2343 181
rect 2377 147 2389 181
rect 2331 141 2389 147
rect 2449 181 2507 187
rect 2449 147 2461 181
rect 2495 147 2507 181
rect 2449 141 2507 147
rect 2567 181 2625 187
rect 2567 147 2579 181
rect 2613 147 2625 181
rect 2567 141 2625 147
rect 2685 181 2743 187
rect 2685 147 2697 181
rect 2731 147 2743 181
rect 2685 141 2743 147
rect -2796 88 -2750 100
rect -2796 -88 -2790 88
rect -2756 -88 -2750 88
rect -2796 -100 -2750 -88
rect -2678 88 -2632 100
rect -2678 -88 -2672 88
rect -2638 -88 -2632 88
rect -2678 -100 -2632 -88
rect -2560 88 -2514 100
rect -2560 -88 -2554 88
rect -2520 -88 -2514 88
rect -2560 -100 -2514 -88
rect -2442 88 -2396 100
rect -2442 -88 -2436 88
rect -2402 -88 -2396 88
rect -2442 -100 -2396 -88
rect -2324 88 -2278 100
rect -2324 -88 -2318 88
rect -2284 -88 -2278 88
rect -2324 -100 -2278 -88
rect -2206 88 -2160 100
rect -2206 -88 -2200 88
rect -2166 -88 -2160 88
rect -2206 -100 -2160 -88
rect -2088 88 -2042 100
rect -2088 -88 -2082 88
rect -2048 -88 -2042 88
rect -2088 -100 -2042 -88
rect -1970 88 -1924 100
rect -1970 -88 -1964 88
rect -1930 -88 -1924 88
rect -1970 -100 -1924 -88
rect -1852 88 -1806 100
rect -1852 -88 -1846 88
rect -1812 -88 -1806 88
rect -1852 -100 -1806 -88
rect -1734 88 -1688 100
rect -1734 -88 -1728 88
rect -1694 -88 -1688 88
rect -1734 -100 -1688 -88
rect -1616 88 -1570 100
rect -1616 -88 -1610 88
rect -1576 -88 -1570 88
rect -1616 -100 -1570 -88
rect -1498 88 -1452 100
rect -1498 -88 -1492 88
rect -1458 -88 -1452 88
rect -1498 -100 -1452 -88
rect -1380 88 -1334 100
rect -1380 -88 -1374 88
rect -1340 -88 -1334 88
rect -1380 -100 -1334 -88
rect -1262 88 -1216 100
rect -1262 -88 -1256 88
rect -1222 -88 -1216 88
rect -1262 -100 -1216 -88
rect -1144 88 -1098 100
rect -1144 -88 -1138 88
rect -1104 -88 -1098 88
rect -1144 -100 -1098 -88
rect -1026 88 -980 100
rect -1026 -88 -1020 88
rect -986 -88 -980 88
rect -1026 -100 -980 -88
rect -908 88 -862 100
rect -908 -88 -902 88
rect -868 -88 -862 88
rect -908 -100 -862 -88
rect -790 88 -744 100
rect -790 -88 -784 88
rect -750 -88 -744 88
rect -790 -100 -744 -88
rect -672 88 -626 100
rect -672 -88 -666 88
rect -632 -88 -626 88
rect -672 -100 -626 -88
rect -554 88 -508 100
rect -554 -88 -548 88
rect -514 -88 -508 88
rect -554 -100 -508 -88
rect -436 88 -390 100
rect -436 -88 -430 88
rect -396 -88 -390 88
rect -436 -100 -390 -88
rect -318 88 -272 100
rect -318 -88 -312 88
rect -278 -88 -272 88
rect -318 -100 -272 -88
rect -200 88 -154 100
rect -200 -88 -194 88
rect -160 -88 -154 88
rect -200 -100 -154 -88
rect -82 88 -36 100
rect -82 -88 -76 88
rect -42 -88 -36 88
rect -82 -100 -36 -88
rect 36 88 82 100
rect 36 -88 42 88
rect 76 -88 82 88
rect 36 -100 82 -88
rect 154 88 200 100
rect 154 -88 160 88
rect 194 -88 200 88
rect 154 -100 200 -88
rect 272 88 318 100
rect 272 -88 278 88
rect 312 -88 318 88
rect 272 -100 318 -88
rect 390 88 436 100
rect 390 -88 396 88
rect 430 -88 436 88
rect 390 -100 436 -88
rect 508 88 554 100
rect 508 -88 514 88
rect 548 -88 554 88
rect 508 -100 554 -88
rect 626 88 672 100
rect 626 -88 632 88
rect 666 -88 672 88
rect 626 -100 672 -88
rect 744 88 790 100
rect 744 -88 750 88
rect 784 -88 790 88
rect 744 -100 790 -88
rect 862 88 908 100
rect 862 -88 868 88
rect 902 -88 908 88
rect 862 -100 908 -88
rect 980 88 1026 100
rect 980 -88 986 88
rect 1020 -88 1026 88
rect 980 -100 1026 -88
rect 1098 88 1144 100
rect 1098 -88 1104 88
rect 1138 -88 1144 88
rect 1098 -100 1144 -88
rect 1216 88 1262 100
rect 1216 -88 1222 88
rect 1256 -88 1262 88
rect 1216 -100 1262 -88
rect 1334 88 1380 100
rect 1334 -88 1340 88
rect 1374 -88 1380 88
rect 1334 -100 1380 -88
rect 1452 88 1498 100
rect 1452 -88 1458 88
rect 1492 -88 1498 88
rect 1452 -100 1498 -88
rect 1570 88 1616 100
rect 1570 -88 1576 88
rect 1610 -88 1616 88
rect 1570 -100 1616 -88
rect 1688 88 1734 100
rect 1688 -88 1694 88
rect 1728 -88 1734 88
rect 1688 -100 1734 -88
rect 1806 88 1852 100
rect 1806 -88 1812 88
rect 1846 -88 1852 88
rect 1806 -100 1852 -88
rect 1924 88 1970 100
rect 1924 -88 1930 88
rect 1964 -88 1970 88
rect 1924 -100 1970 -88
rect 2042 88 2088 100
rect 2042 -88 2048 88
rect 2082 -88 2088 88
rect 2042 -100 2088 -88
rect 2160 88 2206 100
rect 2160 -88 2166 88
rect 2200 -88 2206 88
rect 2160 -100 2206 -88
rect 2278 88 2324 100
rect 2278 -88 2284 88
rect 2318 -88 2324 88
rect 2278 -100 2324 -88
rect 2396 88 2442 100
rect 2396 -88 2402 88
rect 2436 -88 2442 88
rect 2396 -100 2442 -88
rect 2514 88 2560 100
rect 2514 -88 2520 88
rect 2554 -88 2560 88
rect 2514 -100 2560 -88
rect 2632 88 2678 100
rect 2632 -88 2638 88
rect 2672 -88 2678 88
rect 2632 -100 2678 -88
rect 2750 88 2796 100
rect 2750 -88 2756 88
rect 2790 -88 2796 88
rect 2750 -100 2796 -88
rect -2743 -147 -2685 -141
rect -2743 -181 -2731 -147
rect -2697 -181 -2685 -147
rect -2743 -187 -2685 -181
rect -2625 -147 -2567 -141
rect -2625 -181 -2613 -147
rect -2579 -181 -2567 -147
rect -2625 -187 -2567 -181
rect -2507 -147 -2449 -141
rect -2507 -181 -2495 -147
rect -2461 -181 -2449 -147
rect -2507 -187 -2449 -181
rect -2389 -147 -2331 -141
rect -2389 -181 -2377 -147
rect -2343 -181 -2331 -147
rect -2389 -187 -2331 -181
rect -2271 -147 -2213 -141
rect -2271 -181 -2259 -147
rect -2225 -181 -2213 -147
rect -2271 -187 -2213 -181
rect -2153 -147 -2095 -141
rect -2153 -181 -2141 -147
rect -2107 -181 -2095 -147
rect -2153 -187 -2095 -181
rect -2035 -147 -1977 -141
rect -2035 -181 -2023 -147
rect -1989 -181 -1977 -147
rect -2035 -187 -1977 -181
rect -1917 -147 -1859 -141
rect -1917 -181 -1905 -147
rect -1871 -181 -1859 -147
rect -1917 -187 -1859 -181
rect -1799 -147 -1741 -141
rect -1799 -181 -1787 -147
rect -1753 -181 -1741 -147
rect -1799 -187 -1741 -181
rect -1681 -147 -1623 -141
rect -1681 -181 -1669 -147
rect -1635 -181 -1623 -147
rect -1681 -187 -1623 -181
rect -1563 -147 -1505 -141
rect -1563 -181 -1551 -147
rect -1517 -181 -1505 -147
rect -1563 -187 -1505 -181
rect -1445 -147 -1387 -141
rect -1445 -181 -1433 -147
rect -1399 -181 -1387 -147
rect -1445 -187 -1387 -181
rect -1327 -147 -1269 -141
rect -1327 -181 -1315 -147
rect -1281 -181 -1269 -147
rect -1327 -187 -1269 -181
rect -1209 -147 -1151 -141
rect -1209 -181 -1197 -147
rect -1163 -181 -1151 -147
rect -1209 -187 -1151 -181
rect -1091 -147 -1033 -141
rect -1091 -181 -1079 -147
rect -1045 -181 -1033 -147
rect -1091 -187 -1033 -181
rect -973 -147 -915 -141
rect -973 -181 -961 -147
rect -927 -181 -915 -147
rect -973 -187 -915 -181
rect -855 -147 -797 -141
rect -855 -181 -843 -147
rect -809 -181 -797 -147
rect -855 -187 -797 -181
rect -737 -147 -679 -141
rect -737 -181 -725 -147
rect -691 -181 -679 -147
rect -737 -187 -679 -181
rect -619 -147 -561 -141
rect -619 -181 -607 -147
rect -573 -181 -561 -147
rect -619 -187 -561 -181
rect -501 -147 -443 -141
rect -501 -181 -489 -147
rect -455 -181 -443 -147
rect -501 -187 -443 -181
rect -383 -147 -325 -141
rect -383 -181 -371 -147
rect -337 -181 -325 -147
rect -383 -187 -325 -181
rect -265 -147 -207 -141
rect -265 -181 -253 -147
rect -219 -181 -207 -147
rect -265 -187 -207 -181
rect -147 -147 -89 -141
rect -147 -181 -135 -147
rect -101 -181 -89 -147
rect -147 -187 -89 -181
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
rect 89 -147 147 -141
rect 89 -181 101 -147
rect 135 -181 147 -147
rect 89 -187 147 -181
rect 207 -147 265 -141
rect 207 -181 219 -147
rect 253 -181 265 -147
rect 207 -187 265 -181
rect 325 -147 383 -141
rect 325 -181 337 -147
rect 371 -181 383 -147
rect 325 -187 383 -181
rect 443 -147 501 -141
rect 443 -181 455 -147
rect 489 -181 501 -147
rect 443 -187 501 -181
rect 561 -147 619 -141
rect 561 -181 573 -147
rect 607 -181 619 -147
rect 561 -187 619 -181
rect 679 -147 737 -141
rect 679 -181 691 -147
rect 725 -181 737 -147
rect 679 -187 737 -181
rect 797 -147 855 -141
rect 797 -181 809 -147
rect 843 -181 855 -147
rect 797 -187 855 -181
rect 915 -147 973 -141
rect 915 -181 927 -147
rect 961 -181 973 -147
rect 915 -187 973 -181
rect 1033 -147 1091 -141
rect 1033 -181 1045 -147
rect 1079 -181 1091 -147
rect 1033 -187 1091 -181
rect 1151 -147 1209 -141
rect 1151 -181 1163 -147
rect 1197 -181 1209 -147
rect 1151 -187 1209 -181
rect 1269 -147 1327 -141
rect 1269 -181 1281 -147
rect 1315 -181 1327 -147
rect 1269 -187 1327 -181
rect 1387 -147 1445 -141
rect 1387 -181 1399 -147
rect 1433 -181 1445 -147
rect 1387 -187 1445 -181
rect 1505 -147 1563 -141
rect 1505 -181 1517 -147
rect 1551 -181 1563 -147
rect 1505 -187 1563 -181
rect 1623 -147 1681 -141
rect 1623 -181 1635 -147
rect 1669 -181 1681 -147
rect 1623 -187 1681 -181
rect 1741 -147 1799 -141
rect 1741 -181 1753 -147
rect 1787 -181 1799 -147
rect 1741 -187 1799 -181
rect 1859 -147 1917 -141
rect 1859 -181 1871 -147
rect 1905 -181 1917 -147
rect 1859 -187 1917 -181
rect 1977 -147 2035 -141
rect 1977 -181 1989 -147
rect 2023 -181 2035 -147
rect 1977 -187 2035 -181
rect 2095 -147 2153 -141
rect 2095 -181 2107 -147
rect 2141 -181 2153 -147
rect 2095 -187 2153 -181
rect 2213 -147 2271 -141
rect 2213 -181 2225 -147
rect 2259 -181 2271 -147
rect 2213 -187 2271 -181
rect 2331 -147 2389 -141
rect 2331 -181 2343 -147
rect 2377 -181 2389 -147
rect 2331 -187 2389 -181
rect 2449 -147 2507 -141
rect 2449 -181 2461 -147
rect 2495 -181 2507 -147
rect 2449 -187 2507 -181
rect 2567 -147 2625 -141
rect 2567 -181 2579 -147
rect 2613 -181 2625 -147
rect 2567 -187 2625 -181
rect 2685 -147 2743 -141
rect 2685 -181 2697 -147
rect 2731 -181 2743 -147
rect 2685 -187 2743 -181
rect -2743 -255 -2685 -249
rect -2743 -289 -2731 -255
rect -2697 -289 -2685 -255
rect -2743 -295 -2685 -289
rect -2625 -255 -2567 -249
rect -2625 -289 -2613 -255
rect -2579 -289 -2567 -255
rect -2625 -295 -2567 -289
rect -2507 -255 -2449 -249
rect -2507 -289 -2495 -255
rect -2461 -289 -2449 -255
rect -2507 -295 -2449 -289
rect -2389 -255 -2331 -249
rect -2389 -289 -2377 -255
rect -2343 -289 -2331 -255
rect -2389 -295 -2331 -289
rect -2271 -255 -2213 -249
rect -2271 -289 -2259 -255
rect -2225 -289 -2213 -255
rect -2271 -295 -2213 -289
rect -2153 -255 -2095 -249
rect -2153 -289 -2141 -255
rect -2107 -289 -2095 -255
rect -2153 -295 -2095 -289
rect -2035 -255 -1977 -249
rect -2035 -289 -2023 -255
rect -1989 -289 -1977 -255
rect -2035 -295 -1977 -289
rect -1917 -255 -1859 -249
rect -1917 -289 -1905 -255
rect -1871 -289 -1859 -255
rect -1917 -295 -1859 -289
rect -1799 -255 -1741 -249
rect -1799 -289 -1787 -255
rect -1753 -289 -1741 -255
rect -1799 -295 -1741 -289
rect -1681 -255 -1623 -249
rect -1681 -289 -1669 -255
rect -1635 -289 -1623 -255
rect -1681 -295 -1623 -289
rect -1563 -255 -1505 -249
rect -1563 -289 -1551 -255
rect -1517 -289 -1505 -255
rect -1563 -295 -1505 -289
rect -1445 -255 -1387 -249
rect -1445 -289 -1433 -255
rect -1399 -289 -1387 -255
rect -1445 -295 -1387 -289
rect -1327 -255 -1269 -249
rect -1327 -289 -1315 -255
rect -1281 -289 -1269 -255
rect -1327 -295 -1269 -289
rect -1209 -255 -1151 -249
rect -1209 -289 -1197 -255
rect -1163 -289 -1151 -255
rect -1209 -295 -1151 -289
rect -1091 -255 -1033 -249
rect -1091 -289 -1079 -255
rect -1045 -289 -1033 -255
rect -1091 -295 -1033 -289
rect -973 -255 -915 -249
rect -973 -289 -961 -255
rect -927 -289 -915 -255
rect -973 -295 -915 -289
rect -855 -255 -797 -249
rect -855 -289 -843 -255
rect -809 -289 -797 -255
rect -855 -295 -797 -289
rect -737 -255 -679 -249
rect -737 -289 -725 -255
rect -691 -289 -679 -255
rect -737 -295 -679 -289
rect -619 -255 -561 -249
rect -619 -289 -607 -255
rect -573 -289 -561 -255
rect -619 -295 -561 -289
rect -501 -255 -443 -249
rect -501 -289 -489 -255
rect -455 -289 -443 -255
rect -501 -295 -443 -289
rect -383 -255 -325 -249
rect -383 -289 -371 -255
rect -337 -289 -325 -255
rect -383 -295 -325 -289
rect -265 -255 -207 -249
rect -265 -289 -253 -255
rect -219 -289 -207 -255
rect -265 -295 -207 -289
rect -147 -255 -89 -249
rect -147 -289 -135 -255
rect -101 -289 -89 -255
rect -147 -295 -89 -289
rect -29 -255 29 -249
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -295 29 -289
rect 89 -255 147 -249
rect 89 -289 101 -255
rect 135 -289 147 -255
rect 89 -295 147 -289
rect 207 -255 265 -249
rect 207 -289 219 -255
rect 253 -289 265 -255
rect 207 -295 265 -289
rect 325 -255 383 -249
rect 325 -289 337 -255
rect 371 -289 383 -255
rect 325 -295 383 -289
rect 443 -255 501 -249
rect 443 -289 455 -255
rect 489 -289 501 -255
rect 443 -295 501 -289
rect 561 -255 619 -249
rect 561 -289 573 -255
rect 607 -289 619 -255
rect 561 -295 619 -289
rect 679 -255 737 -249
rect 679 -289 691 -255
rect 725 -289 737 -255
rect 679 -295 737 -289
rect 797 -255 855 -249
rect 797 -289 809 -255
rect 843 -289 855 -255
rect 797 -295 855 -289
rect 915 -255 973 -249
rect 915 -289 927 -255
rect 961 -289 973 -255
rect 915 -295 973 -289
rect 1033 -255 1091 -249
rect 1033 -289 1045 -255
rect 1079 -289 1091 -255
rect 1033 -295 1091 -289
rect 1151 -255 1209 -249
rect 1151 -289 1163 -255
rect 1197 -289 1209 -255
rect 1151 -295 1209 -289
rect 1269 -255 1327 -249
rect 1269 -289 1281 -255
rect 1315 -289 1327 -255
rect 1269 -295 1327 -289
rect 1387 -255 1445 -249
rect 1387 -289 1399 -255
rect 1433 -289 1445 -255
rect 1387 -295 1445 -289
rect 1505 -255 1563 -249
rect 1505 -289 1517 -255
rect 1551 -289 1563 -255
rect 1505 -295 1563 -289
rect 1623 -255 1681 -249
rect 1623 -289 1635 -255
rect 1669 -289 1681 -255
rect 1623 -295 1681 -289
rect 1741 -255 1799 -249
rect 1741 -289 1753 -255
rect 1787 -289 1799 -255
rect 1741 -295 1799 -289
rect 1859 -255 1917 -249
rect 1859 -289 1871 -255
rect 1905 -289 1917 -255
rect 1859 -295 1917 -289
rect 1977 -255 2035 -249
rect 1977 -289 1989 -255
rect 2023 -289 2035 -255
rect 1977 -295 2035 -289
rect 2095 -255 2153 -249
rect 2095 -289 2107 -255
rect 2141 -289 2153 -255
rect 2095 -295 2153 -289
rect 2213 -255 2271 -249
rect 2213 -289 2225 -255
rect 2259 -289 2271 -255
rect 2213 -295 2271 -289
rect 2331 -255 2389 -249
rect 2331 -289 2343 -255
rect 2377 -289 2389 -255
rect 2331 -295 2389 -289
rect 2449 -255 2507 -249
rect 2449 -289 2461 -255
rect 2495 -289 2507 -255
rect 2449 -295 2507 -289
rect 2567 -255 2625 -249
rect 2567 -289 2579 -255
rect 2613 -289 2625 -255
rect 2567 -295 2625 -289
rect 2685 -255 2743 -249
rect 2685 -289 2697 -255
rect 2731 -289 2743 -255
rect 2685 -295 2743 -289
rect -2796 -348 -2750 -336
rect -2796 -524 -2790 -348
rect -2756 -524 -2750 -348
rect -2796 -536 -2750 -524
rect -2678 -348 -2632 -336
rect -2678 -524 -2672 -348
rect -2638 -524 -2632 -348
rect -2678 -536 -2632 -524
rect -2560 -348 -2514 -336
rect -2560 -524 -2554 -348
rect -2520 -524 -2514 -348
rect -2560 -536 -2514 -524
rect -2442 -348 -2396 -336
rect -2442 -524 -2436 -348
rect -2402 -524 -2396 -348
rect -2442 -536 -2396 -524
rect -2324 -348 -2278 -336
rect -2324 -524 -2318 -348
rect -2284 -524 -2278 -348
rect -2324 -536 -2278 -524
rect -2206 -348 -2160 -336
rect -2206 -524 -2200 -348
rect -2166 -524 -2160 -348
rect -2206 -536 -2160 -524
rect -2088 -348 -2042 -336
rect -2088 -524 -2082 -348
rect -2048 -524 -2042 -348
rect -2088 -536 -2042 -524
rect -1970 -348 -1924 -336
rect -1970 -524 -1964 -348
rect -1930 -524 -1924 -348
rect -1970 -536 -1924 -524
rect -1852 -348 -1806 -336
rect -1852 -524 -1846 -348
rect -1812 -524 -1806 -348
rect -1852 -536 -1806 -524
rect -1734 -348 -1688 -336
rect -1734 -524 -1728 -348
rect -1694 -524 -1688 -348
rect -1734 -536 -1688 -524
rect -1616 -348 -1570 -336
rect -1616 -524 -1610 -348
rect -1576 -524 -1570 -348
rect -1616 -536 -1570 -524
rect -1498 -348 -1452 -336
rect -1498 -524 -1492 -348
rect -1458 -524 -1452 -348
rect -1498 -536 -1452 -524
rect -1380 -348 -1334 -336
rect -1380 -524 -1374 -348
rect -1340 -524 -1334 -348
rect -1380 -536 -1334 -524
rect -1262 -348 -1216 -336
rect -1262 -524 -1256 -348
rect -1222 -524 -1216 -348
rect -1262 -536 -1216 -524
rect -1144 -348 -1098 -336
rect -1144 -524 -1138 -348
rect -1104 -524 -1098 -348
rect -1144 -536 -1098 -524
rect -1026 -348 -980 -336
rect -1026 -524 -1020 -348
rect -986 -524 -980 -348
rect -1026 -536 -980 -524
rect -908 -348 -862 -336
rect -908 -524 -902 -348
rect -868 -524 -862 -348
rect -908 -536 -862 -524
rect -790 -348 -744 -336
rect -790 -524 -784 -348
rect -750 -524 -744 -348
rect -790 -536 -744 -524
rect -672 -348 -626 -336
rect -672 -524 -666 -348
rect -632 -524 -626 -348
rect -672 -536 -626 -524
rect -554 -348 -508 -336
rect -554 -524 -548 -348
rect -514 -524 -508 -348
rect -554 -536 -508 -524
rect -436 -348 -390 -336
rect -436 -524 -430 -348
rect -396 -524 -390 -348
rect -436 -536 -390 -524
rect -318 -348 -272 -336
rect -318 -524 -312 -348
rect -278 -524 -272 -348
rect -318 -536 -272 -524
rect -200 -348 -154 -336
rect -200 -524 -194 -348
rect -160 -524 -154 -348
rect -200 -536 -154 -524
rect -82 -348 -36 -336
rect -82 -524 -76 -348
rect -42 -524 -36 -348
rect -82 -536 -36 -524
rect 36 -348 82 -336
rect 36 -524 42 -348
rect 76 -524 82 -348
rect 36 -536 82 -524
rect 154 -348 200 -336
rect 154 -524 160 -348
rect 194 -524 200 -348
rect 154 -536 200 -524
rect 272 -348 318 -336
rect 272 -524 278 -348
rect 312 -524 318 -348
rect 272 -536 318 -524
rect 390 -348 436 -336
rect 390 -524 396 -348
rect 430 -524 436 -348
rect 390 -536 436 -524
rect 508 -348 554 -336
rect 508 -524 514 -348
rect 548 -524 554 -348
rect 508 -536 554 -524
rect 626 -348 672 -336
rect 626 -524 632 -348
rect 666 -524 672 -348
rect 626 -536 672 -524
rect 744 -348 790 -336
rect 744 -524 750 -348
rect 784 -524 790 -348
rect 744 -536 790 -524
rect 862 -348 908 -336
rect 862 -524 868 -348
rect 902 -524 908 -348
rect 862 -536 908 -524
rect 980 -348 1026 -336
rect 980 -524 986 -348
rect 1020 -524 1026 -348
rect 980 -536 1026 -524
rect 1098 -348 1144 -336
rect 1098 -524 1104 -348
rect 1138 -524 1144 -348
rect 1098 -536 1144 -524
rect 1216 -348 1262 -336
rect 1216 -524 1222 -348
rect 1256 -524 1262 -348
rect 1216 -536 1262 -524
rect 1334 -348 1380 -336
rect 1334 -524 1340 -348
rect 1374 -524 1380 -348
rect 1334 -536 1380 -524
rect 1452 -348 1498 -336
rect 1452 -524 1458 -348
rect 1492 -524 1498 -348
rect 1452 -536 1498 -524
rect 1570 -348 1616 -336
rect 1570 -524 1576 -348
rect 1610 -524 1616 -348
rect 1570 -536 1616 -524
rect 1688 -348 1734 -336
rect 1688 -524 1694 -348
rect 1728 -524 1734 -348
rect 1688 -536 1734 -524
rect 1806 -348 1852 -336
rect 1806 -524 1812 -348
rect 1846 -524 1852 -348
rect 1806 -536 1852 -524
rect 1924 -348 1970 -336
rect 1924 -524 1930 -348
rect 1964 -524 1970 -348
rect 1924 -536 1970 -524
rect 2042 -348 2088 -336
rect 2042 -524 2048 -348
rect 2082 -524 2088 -348
rect 2042 -536 2088 -524
rect 2160 -348 2206 -336
rect 2160 -524 2166 -348
rect 2200 -524 2206 -348
rect 2160 -536 2206 -524
rect 2278 -348 2324 -336
rect 2278 -524 2284 -348
rect 2318 -524 2324 -348
rect 2278 -536 2324 -524
rect 2396 -348 2442 -336
rect 2396 -524 2402 -348
rect 2436 -524 2442 -348
rect 2396 -536 2442 -524
rect 2514 -348 2560 -336
rect 2514 -524 2520 -348
rect 2554 -524 2560 -348
rect 2514 -536 2560 -524
rect 2632 -348 2678 -336
rect 2632 -524 2638 -348
rect 2672 -524 2678 -348
rect 2632 -536 2678 -524
rect 2750 -348 2796 -336
rect 2750 -524 2756 -348
rect 2790 -524 2796 -348
rect 2750 -536 2796 -524
rect -2743 -583 -2685 -577
rect -2743 -617 -2731 -583
rect -2697 -617 -2685 -583
rect -2743 -623 -2685 -617
rect -2625 -583 -2567 -577
rect -2625 -617 -2613 -583
rect -2579 -617 -2567 -583
rect -2625 -623 -2567 -617
rect -2507 -583 -2449 -577
rect -2507 -617 -2495 -583
rect -2461 -617 -2449 -583
rect -2507 -623 -2449 -617
rect -2389 -583 -2331 -577
rect -2389 -617 -2377 -583
rect -2343 -617 -2331 -583
rect -2389 -623 -2331 -617
rect -2271 -583 -2213 -577
rect -2271 -617 -2259 -583
rect -2225 -617 -2213 -583
rect -2271 -623 -2213 -617
rect -2153 -583 -2095 -577
rect -2153 -617 -2141 -583
rect -2107 -617 -2095 -583
rect -2153 -623 -2095 -617
rect -2035 -583 -1977 -577
rect -2035 -617 -2023 -583
rect -1989 -617 -1977 -583
rect -2035 -623 -1977 -617
rect -1917 -583 -1859 -577
rect -1917 -617 -1905 -583
rect -1871 -617 -1859 -583
rect -1917 -623 -1859 -617
rect -1799 -583 -1741 -577
rect -1799 -617 -1787 -583
rect -1753 -617 -1741 -583
rect -1799 -623 -1741 -617
rect -1681 -583 -1623 -577
rect -1681 -617 -1669 -583
rect -1635 -617 -1623 -583
rect -1681 -623 -1623 -617
rect -1563 -583 -1505 -577
rect -1563 -617 -1551 -583
rect -1517 -617 -1505 -583
rect -1563 -623 -1505 -617
rect -1445 -583 -1387 -577
rect -1445 -617 -1433 -583
rect -1399 -617 -1387 -583
rect -1445 -623 -1387 -617
rect -1327 -583 -1269 -577
rect -1327 -617 -1315 -583
rect -1281 -617 -1269 -583
rect -1327 -623 -1269 -617
rect -1209 -583 -1151 -577
rect -1209 -617 -1197 -583
rect -1163 -617 -1151 -583
rect -1209 -623 -1151 -617
rect -1091 -583 -1033 -577
rect -1091 -617 -1079 -583
rect -1045 -617 -1033 -583
rect -1091 -623 -1033 -617
rect -973 -583 -915 -577
rect -973 -617 -961 -583
rect -927 -617 -915 -583
rect -973 -623 -915 -617
rect -855 -583 -797 -577
rect -855 -617 -843 -583
rect -809 -617 -797 -583
rect -855 -623 -797 -617
rect -737 -583 -679 -577
rect -737 -617 -725 -583
rect -691 -617 -679 -583
rect -737 -623 -679 -617
rect -619 -583 -561 -577
rect -619 -617 -607 -583
rect -573 -617 -561 -583
rect -619 -623 -561 -617
rect -501 -583 -443 -577
rect -501 -617 -489 -583
rect -455 -617 -443 -583
rect -501 -623 -443 -617
rect -383 -583 -325 -577
rect -383 -617 -371 -583
rect -337 -617 -325 -583
rect -383 -623 -325 -617
rect -265 -583 -207 -577
rect -265 -617 -253 -583
rect -219 -617 -207 -583
rect -265 -623 -207 -617
rect -147 -583 -89 -577
rect -147 -617 -135 -583
rect -101 -617 -89 -583
rect -147 -623 -89 -617
rect -29 -583 29 -577
rect -29 -617 -17 -583
rect 17 -617 29 -583
rect -29 -623 29 -617
rect 89 -583 147 -577
rect 89 -617 101 -583
rect 135 -617 147 -583
rect 89 -623 147 -617
rect 207 -583 265 -577
rect 207 -617 219 -583
rect 253 -617 265 -583
rect 207 -623 265 -617
rect 325 -583 383 -577
rect 325 -617 337 -583
rect 371 -617 383 -583
rect 325 -623 383 -617
rect 443 -583 501 -577
rect 443 -617 455 -583
rect 489 -617 501 -583
rect 443 -623 501 -617
rect 561 -583 619 -577
rect 561 -617 573 -583
rect 607 -617 619 -583
rect 561 -623 619 -617
rect 679 -583 737 -577
rect 679 -617 691 -583
rect 725 -617 737 -583
rect 679 -623 737 -617
rect 797 -583 855 -577
rect 797 -617 809 -583
rect 843 -617 855 -583
rect 797 -623 855 -617
rect 915 -583 973 -577
rect 915 -617 927 -583
rect 961 -617 973 -583
rect 915 -623 973 -617
rect 1033 -583 1091 -577
rect 1033 -617 1045 -583
rect 1079 -617 1091 -583
rect 1033 -623 1091 -617
rect 1151 -583 1209 -577
rect 1151 -617 1163 -583
rect 1197 -617 1209 -583
rect 1151 -623 1209 -617
rect 1269 -583 1327 -577
rect 1269 -617 1281 -583
rect 1315 -617 1327 -583
rect 1269 -623 1327 -617
rect 1387 -583 1445 -577
rect 1387 -617 1399 -583
rect 1433 -617 1445 -583
rect 1387 -623 1445 -617
rect 1505 -583 1563 -577
rect 1505 -617 1517 -583
rect 1551 -617 1563 -583
rect 1505 -623 1563 -617
rect 1623 -583 1681 -577
rect 1623 -617 1635 -583
rect 1669 -617 1681 -583
rect 1623 -623 1681 -617
rect 1741 -583 1799 -577
rect 1741 -617 1753 -583
rect 1787 -617 1799 -583
rect 1741 -623 1799 -617
rect 1859 -583 1917 -577
rect 1859 -617 1871 -583
rect 1905 -617 1917 -583
rect 1859 -623 1917 -617
rect 1977 -583 2035 -577
rect 1977 -617 1989 -583
rect 2023 -617 2035 -583
rect 1977 -623 2035 -617
rect 2095 -583 2153 -577
rect 2095 -617 2107 -583
rect 2141 -617 2153 -583
rect 2095 -623 2153 -617
rect 2213 -583 2271 -577
rect 2213 -617 2225 -583
rect 2259 -617 2271 -583
rect 2213 -623 2271 -617
rect 2331 -583 2389 -577
rect 2331 -617 2343 -583
rect 2377 -617 2389 -583
rect 2331 -623 2389 -617
rect 2449 -583 2507 -577
rect 2449 -617 2461 -583
rect 2495 -617 2507 -583
rect 2449 -623 2507 -617
rect 2567 -583 2625 -577
rect 2567 -617 2579 -583
rect 2613 -617 2625 -583
rect 2567 -623 2625 -617
rect 2685 -583 2743 -577
rect 2685 -617 2697 -583
rect 2731 -617 2743 -583
rect 2685 -623 2743 -617
<< properties >>
string FIXED_BBOX -2887 -702 2887 702
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.3 m 3 nf 47 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
