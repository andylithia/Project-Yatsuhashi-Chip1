magic
tech sky130B
magscale 1 2
timestamp 1659144393
<< error_s >>
rect -170 1968 -155 1969
rect -198 1940 -183 1941
rect -198 1860 -180 1940
rect -170 1860 -152 1968
rect -4500 1750 -3930 1790
rect -4400 1670 -4250 1710
rect -4400 1590 -4250 1630
rect -4500 1510 -3930 1550
<< metal1 >>
rect -1250 1750 -1240 1810
rect -210 1750 -200 1810
rect -1250 1740 -200 1750
rect 310 1500 2660 1510
rect -1210 1410 -160 1420
rect -1210 1350 -1200 1410
rect -170 1350 -160 1410
rect 310 1390 320 1500
rect 2640 1390 2660 1500
rect 310 1380 2660 1390
rect -1210 1340 -160 1350
<< via1 >>
rect -1240 1750 -210 1810
rect 340 1710 2660 1820
rect -1200 1350 -170 1410
rect 320 1390 2640 1500
<< metal2 >>
rect -170 1990 0 2010
rect -170 1870 -160 1990
rect -10 1870 0 1990
rect -170 1860 0 1870
rect -1250 1820 2670 1830
rect -1250 1810 100 1820
rect -1250 1750 -1240 1810
rect -210 1750 100 1810
rect -1250 1720 100 1750
rect 250 1720 340 1820
rect -1250 1710 340 1720
rect 2660 1710 2670 1820
rect -1250 1690 2670 1710
rect 310 1500 2660 1510
rect 310 1490 320 1500
rect -10 1480 320 1490
rect -1210 1470 320 1480
rect -1210 1410 -160 1470
rect -1210 1350 -1200 1410
rect -170 1370 -160 1410
rect -10 1390 320 1470
rect 2640 1390 2660 1500
rect -10 1380 2660 1390
rect -10 1370 0 1380
rect -170 1360 0 1370
rect -170 1350 -130 1360
rect -1210 1340 -130 1350
rect 60 1330 260 1340
rect 60 1310 100 1330
rect -150 1230 100 1310
rect 250 1230 260 1330
rect -150 1220 260 1230
<< via2 >>
rect -160 1870 -10 1990
rect 100 1720 250 1820
rect -160 1370 -10 1470
rect 100 1230 250 1330
<< metal3 >>
rect -170 1990 110 2030
rect -170 1870 -160 1990
rect -10 1910 110 1990
rect -10 1870 0 1910
rect -170 1470 0 1870
rect -170 1370 -160 1470
rect -10 1370 0 1470
rect -170 1360 0 1370
rect 90 1820 260 1830
rect 90 1720 100 1820
rect 250 1720 260 1820
rect 90 1330 260 1720
rect 90 1250 100 1330
rect 70 1230 100 1250
rect 250 1230 260 1330
rect 70 1160 260 1230
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659107503
transform 1 0 -870 0 1 -2200
box -500 2210 860 3580
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_1
timestamp 1659107503
transform 1 0 -910 0 -1 5360
box -500 2210 860 3580
use RF_pfet_28xW5p0L0p15  RF_pfet_28xW5p0L0p15_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659106999
transform 1 0 -980 0 1 100
box 980 -100 3880 1386
use RF_pfet_28xW5p0L0p15  RF_pfet_28xW5p0L0p15_1
timestamp 1659106999
transform 1 0 -962 0 -1 3090
box 980 -100 3880 1386
use captuner_complete_1  captuner_complete_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659144393
transform -1 0 -4800 0 1 -550
box -3300 1000 -300 3400
use square_ind_1p12n_5GHz  square_ind_1p12n_5GHz_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1659057364
transform 0 1 3940 -1 0 4478
box 0 -800 20000 20000
<< end >>
