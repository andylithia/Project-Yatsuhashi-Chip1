magic
tech sky130B
timestamp 1659501465
<< metal1 >>
rect 0 140 1000 150
rect 0 105 75 140
rect 175 105 325 140
rect 425 105 575 140
rect 675 105 825 140
rect 925 105 1000 140
rect 0 100 1000 105
rect 0 90 60 100
rect 190 90 310 100
rect 440 90 560 100
rect 690 90 810 100
rect 940 90 1000 100
rect 0 75 50 90
rect 0 -25 10 75
rect 45 -25 50 75
rect 0 -40 50 -25
rect 200 75 300 90
rect 200 -25 205 75
rect 240 -25 260 75
rect 295 -25 300 75
rect 200 -40 300 -25
rect 450 75 550 90
rect 450 -25 455 75
rect 490 -25 510 75
rect 545 -25 550 75
rect 450 -40 550 -25
rect 700 75 800 90
rect 700 -25 705 75
rect 740 -25 760 75
rect 795 -25 800 75
rect 700 -40 800 -25
rect 950 75 1000 90
rect 950 -25 955 75
rect 990 -25 1000 75
rect 950 -40 1000 -25
rect 0 -50 60 -40
rect 190 -50 310 -40
rect 440 -50 560 -40
rect 690 -50 810 -40
rect 940 -50 1000 -40
rect 0 -55 1000 -50
rect 0 -90 75 -55
rect 175 -90 325 -55
rect 425 -90 575 -55
rect 675 -90 825 -55
rect 925 -90 1000 -55
rect 0 -110 1000 -90
rect 0 -145 75 -110
rect 175 -145 325 -110
rect 425 -145 575 -110
rect 675 -145 825 -110
rect 925 -145 1000 -110
rect 0 -150 1000 -145
rect 0 -160 60 -150
rect 190 -160 310 -150
rect 440 -160 560 -150
rect 690 -160 810 -150
rect 940 -160 1000 -150
rect 0 -175 50 -160
rect 0 -275 10 -175
rect 45 -275 50 -175
rect 0 -290 50 -275
rect 200 -175 300 -160
rect 200 -275 205 -175
rect 240 -275 260 -175
rect 295 -275 300 -175
rect 200 -290 300 -275
rect 450 -175 550 -160
rect 450 -275 455 -175
rect 490 -275 510 -175
rect 545 -275 550 -175
rect 450 -290 550 -275
rect 700 -175 800 -160
rect 700 -275 705 -175
rect 740 -275 760 -175
rect 795 -275 800 -175
rect 700 -290 800 -275
rect 950 -175 1000 -160
rect 950 -275 955 -175
rect 990 -275 1000 -175
rect 950 -290 1000 -275
rect 0 -300 60 -290
rect 190 -300 310 -290
rect 440 -300 560 -290
rect 690 -300 810 -290
rect 940 -300 1000 -290
rect 0 -305 1000 -300
rect 0 -340 75 -305
rect 175 -340 325 -305
rect 425 -340 575 -305
rect 675 -340 825 -305
rect 925 -340 1000 -305
rect 0 -360 1000 -340
rect 0 -395 75 -360
rect 175 -395 325 -360
rect 425 -395 575 -360
rect 675 -395 825 -360
rect 925 -395 1000 -360
rect 0 -400 1000 -395
rect 0 -410 60 -400
rect 190 -410 310 -400
rect 440 -410 560 -400
rect 690 -410 810 -400
rect 940 -410 1000 -400
rect 0 -425 50 -410
rect 0 -525 10 -425
rect 45 -525 50 -425
rect 0 -540 50 -525
rect 200 -425 300 -410
rect 200 -525 205 -425
rect 240 -525 260 -425
rect 295 -525 300 -425
rect 200 -540 300 -525
rect 450 -425 550 -410
rect 450 -525 455 -425
rect 490 -525 510 -425
rect 545 -525 550 -425
rect 450 -540 550 -525
rect 700 -425 800 -410
rect 700 -525 705 -425
rect 740 -525 760 -425
rect 795 -525 800 -425
rect 700 -540 800 -525
rect 950 -425 1000 -410
rect 950 -525 955 -425
rect 990 -525 1000 -425
rect 950 -540 1000 -525
rect 0 -550 60 -540
rect 190 -550 310 -540
rect 440 -550 560 -540
rect 690 -550 810 -540
rect 940 -550 1000 -540
rect 0 -555 1000 -550
rect 0 -590 75 -555
rect 175 -590 325 -555
rect 425 -590 575 -555
rect 675 -590 825 -555
rect 925 -590 1000 -555
rect 0 -610 1000 -590
rect 0 -645 75 -610
rect 175 -645 325 -610
rect 425 -645 575 -610
rect 675 -645 825 -610
rect 925 -645 1000 -610
rect 0 -650 1000 -645
rect 0 -660 60 -650
rect 190 -660 310 -650
rect 440 -660 560 -650
rect 690 -660 810 -650
rect 940 -660 1000 -650
rect 0 -675 50 -660
rect 0 -775 10 -675
rect 45 -775 50 -675
rect 0 -790 50 -775
rect 200 -675 300 -660
rect 200 -775 205 -675
rect 240 -775 260 -675
rect 295 -775 300 -675
rect 200 -790 300 -775
rect 450 -675 550 -660
rect 450 -775 455 -675
rect 490 -775 510 -675
rect 545 -775 550 -675
rect 450 -790 550 -775
rect 700 -675 800 -660
rect 700 -775 705 -675
rect 740 -775 760 -675
rect 795 -775 800 -675
rect 700 -790 800 -775
rect 950 -675 1000 -660
rect 950 -775 955 -675
rect 990 -775 1000 -675
rect 950 -790 1000 -775
rect 0 -800 60 -790
rect 190 -800 310 -790
rect 440 -800 560 -790
rect 690 -800 810 -790
rect 940 -800 1000 -790
rect 0 -805 1000 -800
rect 0 -840 75 -805
rect 175 -840 325 -805
rect 425 -840 575 -805
rect 675 -840 825 -805
rect 925 -840 1000 -805
rect 0 -850 1000 -840
<< via1 >>
rect 75 105 175 140
rect 325 105 425 140
rect 575 105 675 140
rect 825 105 925 140
rect 10 -25 45 75
rect 205 -25 240 75
rect 260 -25 295 75
rect 455 -25 490 75
rect 510 -25 545 75
rect 705 -25 740 75
rect 760 -25 795 75
rect 955 -25 990 75
rect 75 -90 175 -55
rect 325 -90 425 -55
rect 575 -90 675 -55
rect 825 -90 925 -55
rect 75 -145 175 -110
rect 325 -145 425 -110
rect 575 -145 675 -110
rect 825 -145 925 -110
rect 10 -275 45 -175
rect 205 -275 240 -175
rect 260 -275 295 -175
rect 455 -275 490 -175
rect 510 -275 545 -175
rect 705 -275 740 -175
rect 760 -275 795 -175
rect 955 -275 990 -175
rect 75 -340 175 -305
rect 325 -340 425 -305
rect 575 -340 675 -305
rect 825 -340 925 -305
rect 75 -395 175 -360
rect 325 -395 425 -360
rect 575 -395 675 -360
rect 825 -395 925 -360
rect 10 -525 45 -425
rect 205 -525 240 -425
rect 260 -525 295 -425
rect 455 -525 490 -425
rect 510 -525 545 -425
rect 705 -525 740 -425
rect 760 -525 795 -425
rect 955 -525 990 -425
rect 75 -590 175 -555
rect 325 -590 425 -555
rect 575 -590 675 -555
rect 825 -590 925 -555
rect 75 -645 175 -610
rect 325 -645 425 -610
rect 575 -645 675 -610
rect 825 -645 925 -610
rect 10 -775 45 -675
rect 205 -775 240 -675
rect 260 -775 295 -675
rect 455 -775 490 -675
rect 510 -775 545 -675
rect 705 -775 740 -675
rect 760 -775 795 -675
rect 955 -775 990 -675
rect 75 -840 175 -805
rect 325 -840 425 -805
rect 575 -840 675 -805
rect 825 -840 925 -805
<< metal2 >>
rect 70 140 180 150
rect 70 105 75 140
rect 175 105 180 140
rect 70 80 180 105
rect 320 140 430 150
rect 320 105 325 140
rect 425 105 430 140
rect 320 80 430 105
rect 570 140 680 150
rect 570 105 575 140
rect 675 105 680 140
rect 570 80 680 105
rect 820 140 930 150
rect 820 105 825 140
rect 925 105 930 140
rect 820 80 930 105
rect 0 75 1000 80
rect 0 -25 10 75
rect 45 -25 205 75
rect 240 -25 260 75
rect 295 -25 455 75
rect 490 -25 510 75
rect 545 -25 705 75
rect 740 -25 760 75
rect 795 -25 955 75
rect 990 -25 1000 75
rect 0 -30 1000 -25
rect 70 -55 180 -30
rect 70 -90 75 -55
rect 175 -90 180 -55
rect 70 -110 180 -90
rect 70 -145 75 -110
rect 175 -145 180 -110
rect 70 -170 180 -145
rect 320 -55 430 -30
rect 320 -90 325 -55
rect 425 -90 430 -55
rect 320 -110 430 -90
rect 320 -145 325 -110
rect 425 -145 430 -110
rect 320 -170 430 -145
rect 570 -55 680 -30
rect 570 -90 575 -55
rect 675 -90 680 -55
rect 570 -110 680 -90
rect 570 -145 575 -110
rect 675 -145 680 -110
rect 570 -170 680 -145
rect 820 -55 930 -30
rect 820 -90 825 -55
rect 925 -90 930 -55
rect 820 -110 930 -90
rect 820 -145 825 -110
rect 925 -145 930 -110
rect 820 -170 930 -145
rect 0 -175 1000 -170
rect 0 -275 10 -175
rect 45 -275 205 -175
rect 240 -275 260 -175
rect 295 -275 455 -175
rect 490 -275 510 -175
rect 545 -275 705 -175
rect 740 -275 760 -175
rect 795 -275 955 -175
rect 990 -275 1000 -175
rect 0 -280 1000 -275
rect 70 -305 180 -280
rect 70 -340 75 -305
rect 175 -340 180 -305
rect 70 -360 180 -340
rect 70 -395 75 -360
rect 175 -395 180 -360
rect 70 -420 180 -395
rect 320 -305 430 -280
rect 320 -340 325 -305
rect 425 -340 430 -305
rect 320 -360 430 -340
rect 320 -395 325 -360
rect 425 -395 430 -360
rect 320 -420 430 -395
rect 570 -305 680 -280
rect 570 -340 575 -305
rect 675 -340 680 -305
rect 570 -360 680 -340
rect 570 -395 575 -360
rect 675 -395 680 -360
rect 570 -420 680 -395
rect 820 -305 930 -280
rect 820 -340 825 -305
rect 925 -340 930 -305
rect 820 -360 930 -340
rect 820 -395 825 -360
rect 925 -395 930 -360
rect 820 -420 930 -395
rect 0 -425 1000 -420
rect 0 -525 10 -425
rect 45 -525 205 -425
rect 240 -525 260 -425
rect 295 -525 455 -425
rect 490 -525 510 -425
rect 545 -525 705 -425
rect 740 -525 760 -425
rect 795 -525 955 -425
rect 990 -525 1000 -425
rect 0 -530 1000 -525
rect 70 -555 180 -530
rect 70 -590 75 -555
rect 175 -590 180 -555
rect 70 -610 180 -590
rect 70 -645 75 -610
rect 175 -645 180 -610
rect 70 -670 180 -645
rect 320 -555 430 -530
rect 320 -590 325 -555
rect 425 -590 430 -555
rect 320 -610 430 -590
rect 320 -645 325 -610
rect 425 -645 430 -610
rect 320 -670 430 -645
rect 570 -555 680 -530
rect 570 -590 575 -555
rect 675 -590 680 -555
rect 570 -610 680 -590
rect 570 -645 575 -610
rect 675 -645 680 -610
rect 570 -670 680 -645
rect 820 -555 930 -530
rect 820 -590 825 -555
rect 925 -590 930 -555
rect 820 -610 930 -590
rect 820 -645 825 -610
rect 925 -645 930 -610
rect 820 -670 930 -645
rect 0 -675 1000 -670
rect 0 -775 10 -675
rect 45 -775 205 -675
rect 240 -775 260 -675
rect 295 -775 455 -675
rect 490 -775 510 -675
rect 545 -775 705 -675
rect 740 -775 760 -675
rect 795 -775 955 -675
rect 990 -775 1000 -675
rect 0 -780 1000 -775
rect 70 -805 180 -780
rect 70 -840 75 -805
rect 175 -840 180 -805
rect 70 -850 180 -840
rect 320 -805 430 -780
rect 320 -840 325 -805
rect 425 -840 430 -805
rect 320 -850 430 -840
rect 570 -805 680 -780
rect 570 -840 575 -805
rect 675 -840 680 -805
rect 570 -850 680 -840
rect 820 -805 930 -780
rect 820 -840 825 -805
rect 925 -840 930 -805
rect 820 -850 930 -840
<< via2 >>
rect 75 105 175 140
rect 325 105 425 140
rect 575 105 675 140
rect 825 105 925 140
rect 10 -25 45 75
rect 205 -25 240 75
rect 260 -25 295 75
rect 455 -25 490 75
rect 510 -25 545 75
rect 705 -25 740 75
rect 760 -25 795 75
rect 955 -25 990 75
rect 75 -90 175 -55
rect 75 -145 175 -110
rect 325 -90 425 -55
rect 325 -145 425 -110
rect 575 -90 675 -55
rect 575 -145 675 -110
rect 825 -90 925 -55
rect 825 -145 925 -110
rect 10 -275 45 -175
rect 205 -275 240 -175
rect 260 -275 295 -175
rect 455 -275 490 -175
rect 510 -275 545 -175
rect 705 -275 740 -175
rect 760 -275 795 -175
rect 955 -275 990 -175
rect 75 -340 175 -305
rect 75 -395 175 -360
rect 325 -340 425 -305
rect 325 -395 425 -360
rect 575 -340 675 -305
rect 575 -395 675 -360
rect 825 -340 925 -305
rect 825 -395 925 -360
rect 10 -525 45 -425
rect 205 -525 240 -425
rect 260 -525 295 -425
rect 455 -525 490 -425
rect 510 -525 545 -425
rect 705 -525 740 -425
rect 760 -525 795 -425
rect 955 -525 990 -425
rect 75 -590 175 -555
rect 75 -645 175 -610
rect 325 -590 425 -555
rect 325 -645 425 -610
rect 575 -590 675 -555
rect 575 -645 675 -610
rect 825 -590 925 -555
rect 825 -645 925 -610
rect 10 -775 45 -675
rect 205 -775 240 -675
rect 260 -775 295 -675
rect 455 -775 490 -675
rect 510 -775 545 -675
rect 705 -775 740 -675
rect 760 -775 795 -675
rect 955 -775 990 -675
rect 75 -840 175 -805
rect 325 -840 425 -805
rect 575 -840 675 -805
rect 825 -840 925 -805
<< metal3 >>
rect 0 140 1000 150
rect 0 105 75 140
rect 175 105 325 140
rect 425 105 575 140
rect 675 105 825 140
rect 925 105 1000 140
rect 0 100 1000 105
rect 0 90 60 100
rect 190 90 310 100
rect 440 90 560 100
rect 690 90 810 100
rect 940 90 1000 100
rect 0 75 50 90
rect 0 -25 10 75
rect 45 -25 50 75
rect 0 -40 50 -25
rect 200 75 300 90
rect 200 -25 205 75
rect 240 -25 260 75
rect 295 -25 300 75
rect 200 -40 300 -25
rect 450 75 550 90
rect 450 -25 455 75
rect 490 -25 510 75
rect 545 -25 550 75
rect 450 -40 550 -25
rect 700 75 800 90
rect 700 -25 705 75
rect 740 -25 760 75
rect 795 -25 800 75
rect 700 -40 800 -25
rect 950 75 1000 90
rect 950 -25 955 75
rect 990 -25 1000 75
rect 950 -40 1000 -25
rect 0 -50 60 -40
rect 190 -50 310 -40
rect 440 -50 560 -40
rect 690 -50 810 -40
rect 940 -50 1000 -40
rect 0 -55 200 -50
rect 0 -90 75 -55
rect 175 -90 200 -55
rect 0 -110 200 -90
rect 0 -145 75 -110
rect 175 -145 200 -110
rect 0 -150 200 -145
rect 300 -55 450 -50
rect 300 -90 325 -55
rect 425 -90 450 -55
rect 300 -110 450 -90
rect 300 -145 325 -110
rect 425 -145 450 -110
rect 300 -150 450 -145
rect 550 -55 700 -50
rect 550 -90 575 -55
rect 675 -90 700 -55
rect 550 -110 700 -90
rect 550 -145 575 -110
rect 675 -145 700 -110
rect 550 -150 700 -145
rect 800 -55 1000 -50
rect 800 -90 825 -55
rect 925 -90 1000 -55
rect 800 -110 1000 -90
rect 800 -145 825 -110
rect 925 -145 1000 -110
rect 800 -150 1000 -145
rect 0 -160 60 -150
rect 190 -160 310 -150
rect 440 -160 560 -150
rect 690 -160 810 -150
rect 940 -160 1000 -150
rect 0 -175 50 -160
rect 0 -275 10 -175
rect 45 -275 50 -175
rect 0 -290 50 -275
rect 200 -175 300 -160
rect 200 -275 205 -175
rect 240 -275 260 -175
rect 295 -275 300 -175
rect 200 -290 300 -275
rect 450 -175 550 -160
rect 450 -275 455 -175
rect 490 -275 510 -175
rect 545 -275 550 -175
rect 450 -290 550 -275
rect 700 -175 800 -160
rect 700 -275 705 -175
rect 740 -275 760 -175
rect 795 -275 800 -175
rect 700 -290 800 -275
rect 950 -175 1000 -160
rect 950 -275 955 -175
rect 990 -275 1000 -175
rect 950 -290 1000 -275
rect 0 -300 60 -290
rect 190 -300 310 -290
rect 440 -300 560 -290
rect 690 -300 810 -290
rect 940 -300 1000 -290
rect 0 -305 200 -300
rect 0 -340 75 -305
rect 175 -340 200 -305
rect 0 -360 200 -340
rect 0 -395 75 -360
rect 175 -395 200 -360
rect 0 -400 200 -395
rect 300 -305 450 -300
rect 300 -340 325 -305
rect 425 -340 450 -305
rect 300 -360 450 -340
rect 300 -395 325 -360
rect 425 -395 450 -360
rect 300 -400 450 -395
rect 550 -305 700 -300
rect 550 -340 575 -305
rect 675 -340 700 -305
rect 550 -360 700 -340
rect 550 -395 575 -360
rect 675 -395 700 -360
rect 550 -400 700 -395
rect 800 -305 1000 -300
rect 800 -340 825 -305
rect 925 -340 1000 -305
rect 800 -360 1000 -340
rect 800 -395 825 -360
rect 925 -395 1000 -360
rect 800 -400 1000 -395
rect 0 -410 60 -400
rect 190 -410 310 -400
rect 440 -410 560 -400
rect 690 -410 810 -400
rect 940 -410 1000 -400
rect 0 -425 50 -410
rect 0 -525 10 -425
rect 45 -525 50 -425
rect 0 -540 50 -525
rect 200 -425 300 -410
rect 200 -525 205 -425
rect 240 -525 260 -425
rect 295 -525 300 -425
rect 200 -540 300 -525
rect 450 -425 550 -410
rect 450 -525 455 -425
rect 490 -525 510 -425
rect 545 -525 550 -425
rect 450 -540 550 -525
rect 700 -425 800 -410
rect 700 -525 705 -425
rect 740 -525 760 -425
rect 795 -525 800 -425
rect 700 -540 800 -525
rect 950 -425 1000 -410
rect 950 -525 955 -425
rect 990 -525 1000 -425
rect 950 -540 1000 -525
rect 0 -550 60 -540
rect 190 -550 310 -540
rect 440 -550 560 -540
rect 690 -550 810 -540
rect 940 -550 1000 -540
rect 0 -555 200 -550
rect 0 -590 75 -555
rect 175 -590 200 -555
rect 0 -610 200 -590
rect 0 -645 75 -610
rect 175 -645 200 -610
rect 0 -650 200 -645
rect 300 -555 450 -550
rect 300 -590 325 -555
rect 425 -590 450 -555
rect 300 -610 450 -590
rect 300 -645 325 -610
rect 425 -645 450 -610
rect 300 -650 450 -645
rect 550 -555 700 -550
rect 550 -590 575 -555
rect 675 -590 700 -555
rect 550 -610 700 -590
rect 550 -645 575 -610
rect 675 -645 700 -610
rect 550 -650 700 -645
rect 800 -555 1000 -550
rect 800 -590 825 -555
rect 925 -590 1000 -555
rect 800 -610 1000 -590
rect 800 -645 825 -610
rect 925 -645 1000 -610
rect 800 -650 1000 -645
rect 0 -660 60 -650
rect 190 -660 310 -650
rect 440 -660 560 -650
rect 690 -660 810 -650
rect 940 -660 1000 -650
rect 0 -675 50 -660
rect 0 -775 10 -675
rect 45 -775 50 -675
rect 0 -790 50 -775
rect 200 -675 300 -660
rect 200 -775 205 -675
rect 240 -775 260 -675
rect 295 -775 300 -675
rect 200 -790 300 -775
rect 450 -675 550 -660
rect 450 -775 455 -675
rect 490 -775 510 -675
rect 545 -775 550 -675
rect 450 -790 550 -775
rect 700 -675 800 -660
rect 700 -775 705 -675
rect 740 -775 760 -675
rect 795 -775 800 -675
rect 700 -790 800 -775
rect 950 -675 1000 -660
rect 950 -775 955 -675
rect 990 -775 1000 -675
rect 950 -790 1000 -775
rect 0 -800 60 -790
rect 190 -800 310 -790
rect 440 -800 560 -790
rect 690 -800 810 -790
rect 940 -800 1000 -790
rect 0 -805 1000 -800
rect 0 -840 75 -805
rect 175 -840 325 -805
rect 425 -840 575 -805
rect 675 -840 825 -805
rect 925 -840 1000 -805
rect 0 -850 1000 -840
<< via3 >>
rect 200 -150 300 -50
rect 450 -150 550 -50
rect 700 -150 800 -50
rect 200 -400 300 -300
rect 450 -400 550 -300
rect 700 -400 800 -300
rect 200 -650 300 -550
rect 450 -650 550 -550
rect 700 -650 800 -550
<< metal4 >>
rect 260 -30 740 150
rect 180 -50 820 -30
rect 180 -110 200 -50
rect 0 -150 200 -110
rect 300 -150 450 -50
rect 550 -150 700 -50
rect 800 -110 820 -50
rect 800 -150 1000 -110
rect 0 -300 1000 -150
rect 0 -400 200 -300
rect 300 -400 450 -300
rect 550 -400 700 -300
rect 800 -400 1000 -300
rect 0 -550 1000 -400
rect 0 -590 200 -550
rect 180 -650 200 -590
rect 300 -650 450 -550
rect 550 -650 700 -550
rect 800 -590 1000 -550
rect 800 -650 820 -590
rect 180 -670 820 -650
rect 260 -850 740 -670
<< end >>
