** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/zptest.sch
**.subckt zptest
V1 net6 GND 1.8
V2 net9 GND dc 0 ac 1 portnum 1 z0 50
V3 net8 GND dc 0 ac 1 portnum 2 z0 50
Ldeg3 net2 net1 0.5n m=1
C2 net3 net9 1n m=1
R1 vgate1 vbias1 2k m=1
C4 net3 GND 50f m=1
Ldeg1 vgate1 net4 2n m=1
Ldeg4 net4 net3 1n m=1
C6 net4 GND 50f m=1
R2 net5 net6 2k m=1
I0 GND vbias1 1m
Ldeg2 net19 net7 3n m=1
XM5 n_ds1 vgate1 net2 net1 sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=6
XM1 vbias1 vbias1 GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
XM2 net7 net5 n_ds1 net1 sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=6
XC5 net7 net10 sky130_fd_pr__cap_mim_m3_1 W=5 L=1 MF=1 m=1
XC10 net7 net11 sky130_fd_pr__cap_mim_m3_1 W=5 L=2 MF=1 m=1
XC9 net7 net12 sky130_fd_pr__cap_mim_m3_1 W=5 L=4 MF=1 m=1
XC11 net7 net13 sky130_fd_pr__cap_mim_m3_1 W=5 L=8 MF=1 m=1
XM3 net10 net6 GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
XM4 net11 net6 GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
XM6 net12 net6 GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
XM7 net13 GND GND GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
XC12 net8 net7 sky130_fd_pr__cap_mim_m3_1 W=10 L=6 MF=1 m=1
XC1 net5 GND sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=1 m=1
XC7 vbias1 GND sky130_fd_pr__cap_mim_m3_1 W=20 L=10 MF=1 m=1
XC13 vgate1 net14 sky130_fd_pr__cap_mim_m3_1 W=7 L=1 MF=1 m=1
XC14 vgate1 net15 sky130_fd_pr__cap_mim_m3_1 W=7 L=2 MF=1 m=1
XC15 vgate1 net16 sky130_fd_pr__cap_mim_m3_1 W=7 L=4 MF=1 m=1
XC16 vgate1 net17 sky130_fd_pr__cap_mim_m3_1 W=7 L=8 MF=1 m=1
XM8 net14 net6 net2 GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
XM9 net15 net6 net2 GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
XM10 net16 net6 net2 GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
XM11 net17 GND net2 GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
Ldeg5 net18 net19 2n m=1
R3 net18 net6 5 m=1
C3 net19 GND 10p m=1
Ldeg6 net20 GND 2n m=1
R4 net20 net1 5 m=1
C8 net1 GND 10p m=1
R5 net21 net7 2k m=1
XC17 net21 vgate1 sky130_fd_pr__cap_mim_m3_1 W=10 L=100 MF=1 m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice



.subckt sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=2.828e+12p pd=2.132e+07u as=4.242e+12p
+ ps=3.198e+07u w=5.05e+06u l=150000u
X1 SOURCE SUBSTRATE SUBSTRATE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.03e+12p
+ ps=2.14e+07u w=5.05e+06u l=150000u
X2 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X5 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends
.sp dec 1000 1e9 10e9 1
* .ac dec 1000 0.01e9 100e9
.control
run
display

let S11 = S_1_1
let S21 = S_2_1
let S12 = S_1_2
let S22 = S_2_2

* Stability
let delta=S11*S22-S12*S21
let K    = (1-mag(S11)^2-mag(S22)^2+mag(delta)^2)/(2*mag(S12*S21))
let mu   = (1-mag(S11)^2)/(mag(S22-conj(S11)*delta)+mag(S21*S12))

let z11=50*(1+s_1_1)/(1-s_1_1)
let z22=50*(1+s_2_2)/(1-s_2_2)
plot real(z11) real(z22)
plot imag(z11) imag(z22)
plot db(S_1_1) db(S_2_2) db(S_2_1)

plot mag(delta)
plot (K)
plot (mu)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
