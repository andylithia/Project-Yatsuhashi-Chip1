* NGSPICE file created from ./CLASSE/cascode_2.ext - technology: sky130A

X0 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X1 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X2 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X3 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X4 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X5 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X6 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X7 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X8 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X9 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X10 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X11 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X12 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X13 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X14 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X15 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X16 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X17 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X18 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X19 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X20 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X21 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X22 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X23 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X24 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X25 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X26 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X27 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X28 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X29 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X30 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X31 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X32 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X33 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X34 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X35 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X36 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X37 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X38 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X39 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X40 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X41 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X42 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X43 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X44 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X45 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X46 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X47 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X48 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X49 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X50 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X51 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X52 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X53 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X54 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X55 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X56 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X57 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X58 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X59 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X60 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X61 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X62 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X63 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X64 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X65 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X66 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X67 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X68 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X69 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X70 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X71 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X72 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X73 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X74 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X75 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X76 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X77 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X78 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X79 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X80 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X81 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X82 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X83 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X84 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X85 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X86 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X87 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X88 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X89 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X90 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X91 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X92 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X93 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X94 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X95 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X96 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X97 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X98 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X99 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X100 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X101 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X102 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X103 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X104 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X105 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X106 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X107 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X108 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X109 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X110 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X111 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X112 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X113 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X114 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X115 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X116 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X117 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X118 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X119 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X120 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X121 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X122 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X123 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X124 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X125 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X126 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X127 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X128 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X129 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X130 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X131 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X132 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X133 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X134 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X135 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X136 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X137 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X138 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X139 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X140 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X141 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X142 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X143 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X144 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X145 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X146 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X147 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X148 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X149 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X150 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X151 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X152 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X153 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X154 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X155 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X156 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X157 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X158 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X159 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X160 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X161 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X162 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X163 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X164 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X165 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X166 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X167 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X168 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X169 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X170 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X171 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X172 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X173 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X174 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X175 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X176 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X177 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X178 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X179 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X180 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X181 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X182 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X183 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X184 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X185 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X186 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X187 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X188 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X189 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X190 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X191 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X192 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X193 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X194 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X195 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X196 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X197 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X198 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X199 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X200 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X201 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X202 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X203 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X204 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X205 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X206 SD1L G12L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X207 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X208 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X209 SD3L G12L SD1L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X210 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X211 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X212 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X213 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X214 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X215 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X216 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X217 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X218 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X219 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X220 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X221 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X222 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X223 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X224 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X225 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X226 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X227 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X228 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X229 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X230 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X231 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X232 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X233 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X234 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X235 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X236 SD1R G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X237 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X238 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X239 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G12R SD1R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X240 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X241 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X242 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X243 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X244 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X245 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X246 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X247 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X248 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X249 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X250 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X251 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X252 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X253 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X254 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X255 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X256 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X257 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X258 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X259 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X260 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X261 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X262 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X263 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X264 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X265 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X266 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X267 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X268 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X269 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X270 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X271 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X272 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X273 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X274 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X275 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X276 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X277 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X278 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X279 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X280 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X281 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X282 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X283 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X284 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X285 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X286 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X287 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X288 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X289 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X290 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X291 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X292 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X293 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X294 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X295 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X296 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X297 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X298 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X299 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X300 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X301 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X302 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X303 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X304 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X305 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X306 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X307 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X308 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X309 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X310 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X311 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X312 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X313 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X314 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X315 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X316 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X317 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X318 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X319 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X320 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X321 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X322 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X323 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X324 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X325 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X326 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X327 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X328 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X329 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X330 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X331 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X332 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X333 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X334 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X335 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X336 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X337 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X338 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X339 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X340 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X341 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X342 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X343 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X344 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X345 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X346 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X347 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X348 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X349 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X350 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X351 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X352 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X353 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X354 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X355 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X356 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X357 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X358 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X359 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X360 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X361 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X362 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X363 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X364 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X365 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X366 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X367 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X368 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X369 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X370 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X371 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X372 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X373 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X374 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X375 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X376 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X377 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X378 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X379 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X380 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X381 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X382 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X383 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X384 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X385 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X386 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X387 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X388 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X389 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X390 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X391 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X392 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X393 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X394 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X395 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X396 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X397 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X398 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X399 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X400 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X401 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X402 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X403 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X404 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X405 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X406 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X407 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X408 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X409 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X410 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X411 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X412 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X413 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X414 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X415 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X416 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X417 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X418 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X419 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X420 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X421 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X422 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X423 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X424 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X425 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X426 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X427 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X428 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X429 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X430 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X431 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X432 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X433 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X434 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X435 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X436 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X437 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X438 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X439 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X440 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X441 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X442 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X443 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X444 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X445 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X446 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X447 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X448 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X449 SD3L G23L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X450 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X451 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X452 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X453 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X454 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X455 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X456 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X457 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X458 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X459 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X460 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X461 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X462 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X463 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X464 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X465 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X466 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X467 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X468 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X469 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X470 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X471 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X472 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X473 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X474 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X475 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X476 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X477 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X478 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X479 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X480 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X481 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X482 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X483 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X484 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X485 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X486 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X487 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X488 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X489 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X490 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X491 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X492 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X493 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X494 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X495 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X496 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X497 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X498 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X499 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X500 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X501 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X502 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X503 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X504 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X505 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X506 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X507 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X508 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X509 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X510 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X511 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X512 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X513 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X514 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X515 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X516 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X517 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X518 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X519 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X520 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X521 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X522 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X523 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X524 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X525 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X526 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X527 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X528 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X529 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X530 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X531 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X532 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X533 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X534 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X535 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X536 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X537 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X538 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X539 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X540 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X541 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X542 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X543 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X544 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X545 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X546 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X547 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X548 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X549 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X550 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X551 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X552 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X553 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X554 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X555 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X556 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X557 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X558 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X559 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X560 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X561 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X562 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X563 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X564 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X565 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X566 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X567 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X568 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X569 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X570 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X571 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X572 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X573 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X574 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X575 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X576 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X577 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X578 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X579 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X580 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X581 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X582 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X583 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X584 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X585 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X586 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X587 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X588 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X589 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X590 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X591 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X592 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X593 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X594 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X595 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X596 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X597 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X598 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X599 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X600 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X601 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X602 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X603 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X604 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X605 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X606 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X607 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X608 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X609 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X610 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X611 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X612 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X613 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X614 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X615 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X616 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X617 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X618 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X619 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X620 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X621 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X622 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X623 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X624 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X625 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X626 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X627 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X628 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X629 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X630 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X631 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X632 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X633 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X634 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X635 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X636 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X637 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X638 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X639 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X640 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X641 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X642 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X643 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X644 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X645 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X646 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X647 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X648 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X649 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X650 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X651 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X652 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X653 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X654 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X655 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X656 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X657 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X658 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X659 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X660 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X661 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X662 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X663 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X664 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X665 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X666 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X667 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X668 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X669 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X670 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X671 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X672 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X673 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X674 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X675 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X676 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X677 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X678 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X679 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X680 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X681 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X682 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X683 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X684 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X685 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X686 SD3L G34L SD4L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X687 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X688 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X689 SD4L G34L SD3L VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X690 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X691 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X692 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X693 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X694 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X695 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X696 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X697 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X698 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X699 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X700 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X701 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X702 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X703 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X704 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X705 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X706 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X707 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X708 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X709 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X710 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X711 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X712 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X713 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X714 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X715 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X716 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R SD4R VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X717 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X718 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X719 SD4R G34R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
C0 G23L NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 14.42fF
C1 SD1L SD3L 675.49fF
C2 G12R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 80.61fF
C3 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 670.04fF
C4 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34L 14.42fF
C5 G12L NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 17.62fF
C6 G34R G34L 29.94fF
C7 SD3L NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 157.48fF
C8 SD3L G34L 86.11fF
C9 G23L G23R 29.94fF
C10 SD1L NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 43.91fF
C11 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 SD4L 36.59fF
C12 SD4L G34R 13.55fF
C13 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23R 80.93fF
C14 SD3L SD4L 675.30fF
C15 G23R SD3L 31.85fF
C16 SD1R G12R 83.48fF
C17 G12L SD1R 16.09fF
C18 SD4L G34L 77.89fF
C19 SD1R SD3L 37.13fF
C20 G23R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 82.64fF
C21 SD1R SD1L 57.82fF
C22 SD1R NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 670.56fF
C23 SD4R NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 670.23fF
C24 SD4R G34R 77.97fF
C25 SD4R SD3L 38.75fF
C26 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G23L 17.96fF
C27 G12L G12R 29.94fF
C28 G23L SD3L 164.25fF
C29 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 G34R 82.64fF
C30 SD4R G34L 14.16fF
C31 G12R SD3L 13.55fF
C32 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 SD3L 158.68fF
C33 G12L SD3L 78.01fF
C34 SD3L G34R 18.13fF
C35 SD1L G12R 16.11fF
C36 G12L SD1L 81.48fF
C37 SD4R SD4L 61.24fF
C38 SD4R VSUBS 45.52fF $ **FLOATING
C39 G34R VSUBS 75.89fF $ **FLOATING
C40 SD4L VSUBS 34.69fF $ **FLOATING
C41 G34L VSUBS 75.93fF $ **FLOATING
C42 G23R VSUBS 75.89fF $ **FLOATING
C43 G23L VSUBS 75.93fF $ **FLOATING
C44 NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 VSUBS 91.15fF $ **FLOATING
C45 NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 VSUBS 90.81fF $ **FLOATING
C46 G12R VSUBS 75.89fF $ **FLOATING
C47 SD3L VSUBS 149.14fF $ **FLOATING
C48 G12L VSUBS 75.93fF $ **FLOATING
C49 SD1R VSUBS 50.84fF $ **FLOATING
C50 SD1L VSUBS 45.19fF $ **FLOATING
