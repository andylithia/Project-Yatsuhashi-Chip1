magic
tech sky130B
magscale 1 2
timestamp 1660524432
<< locali >>
rect 678 9488 1320 9522
rect 582 7778 1224 7812
<< metal1 >>
rect 660 9550 1320 9560
rect 660 9490 670 9550
rect 1310 9490 1320 9550
rect 660 9480 1320 9490
rect 540 9410 600 9450
rect 540 7850 600 7890
rect 630 9410 690 9450
rect 630 7850 690 7890
rect 730 9410 790 9450
rect 730 7850 790 7890
rect 830 9410 890 9450
rect 830 7850 890 7890
rect 920 9410 980 9450
rect 920 7850 980 7890
rect 1020 9410 1080 9450
rect 1020 7850 1080 7890
rect 1110 9410 1170 9450
rect 1110 7850 1170 7890
rect 1210 9410 1270 9450
rect 1210 7850 1270 7890
rect 1310 9410 1370 9450
rect 1310 7850 1370 7890
rect 570 7810 1230 7820
rect 570 7750 580 7810
rect 1220 7750 1230 7810
rect 570 7740 1230 7750
rect 0 7580 200 7600
rect 0 7120 20 7580
rect 180 7120 200 7580
rect 10200 7580 10400 7600
rect 10200 7420 10220 7580
rect 10380 7420 10400 7580
rect 10200 7400 10400 7420
rect 0 7100 200 7120
rect 0 6480 200 6500
rect 0 6120 20 6480
rect 180 6120 200 6480
rect 0 6100 200 6120
rect 10200 380 10400 400
rect 10200 220 10220 380
rect 10380 220 10400 380
rect 10200 200 10400 220
<< via1 >>
rect 670 9490 1310 9550
rect 540 7890 600 9410
rect 630 7890 690 9410
rect 730 7890 790 9410
rect 830 7890 890 9410
rect 920 7890 980 9410
rect 1020 7890 1080 9410
rect 1110 7890 1170 9410
rect 1210 7890 1270 9410
rect 1310 7890 1370 9410
rect 580 7750 1220 7810
rect 20 7120 180 7580
rect 10220 7420 10380 7580
rect 20 6120 180 6480
rect 10220 220 10380 380
<< metal2 >>
rect 630 9550 1320 9560
rect 630 9490 670 9550
rect 1310 9490 1320 9550
rect 630 9480 1320 9490
rect 540 9410 600 9450
rect 540 7850 600 7890
rect 630 9410 690 9480
rect 630 7820 690 7890
rect 730 9410 790 9450
rect 730 7850 790 7890
rect 830 9410 890 9480
rect 830 7820 890 7890
rect 920 9410 980 9450
rect 920 7850 980 7890
rect 1020 9410 1080 9480
rect 1020 7820 1080 7890
rect 1110 9410 1170 9450
rect 1110 7850 1170 7890
rect 1210 9410 1270 9480
rect 1210 7820 1270 7890
rect 1310 9410 1370 9450
rect 1310 7850 1370 7890
rect 570 7810 1270 7820
rect 570 7750 580 7810
rect 1220 7750 1270 7810
rect 570 7740 1270 7750
rect 0 7580 200 7600
rect 0 7120 20 7580
rect 180 7120 200 7580
rect 10200 7580 10400 7600
rect 10200 7420 10220 7580
rect 10380 7420 10400 7580
rect 10200 7400 10400 7420
rect 0 7100 200 7120
rect 0 6480 200 6500
rect 0 6120 20 6480
rect 180 6120 200 6480
rect 0 6100 200 6120
rect 10200 380 10400 400
rect 10200 220 10220 380
rect 10380 220 10400 380
rect 10200 200 10400 220
<< via2 >>
rect 670 9490 1310 9550
rect 540 8270 600 9030
rect 730 8270 790 9030
rect 920 8270 980 9030
rect 1110 8270 1170 9030
rect 1310 8270 1370 9030
rect 580 7750 1220 7810
rect 20 7120 180 7580
rect 10220 7420 10380 7580
rect 20 6120 180 6480
rect 10220 220 10380 380
<< metal3 >>
rect -1600 12400 1000 12600
rect -1600 11800 -1400 12400
rect 800 11800 1000 12400
rect -1600 11400 1000 11800
rect -1600 9560 400 11400
rect -1600 9550 1320 9560
rect -1600 9490 670 9550
rect 1310 9490 1320 9550
rect -1600 9480 1320 9490
rect -8000 8400 -4000 8600
rect -8000 6000 -7800 8400
rect -4200 7200 -4000 8400
rect -1600 7920 420 9480
rect 1440 9050 1620 9060
rect 520 9030 1620 9050
rect 520 8270 540 9030
rect 600 8980 730 9030
rect 600 8700 620 8980
rect 710 8700 730 8980
rect 600 8620 730 8700
rect 600 8320 620 8620
rect 710 8320 730 8620
rect 600 8270 730 8320
rect 790 8980 920 9030
rect 790 8700 810 8980
rect 900 8700 920 8980
rect 790 8620 920 8700
rect 790 8320 810 8620
rect 900 8320 920 8620
rect 790 8270 920 8320
rect 980 8980 1110 9030
rect 980 8700 1000 8980
rect 1090 8700 1110 8980
rect 980 8620 1110 8700
rect 980 8320 1000 8620
rect 1090 8320 1110 8620
rect 980 8270 1110 8320
rect 1170 8980 1310 9030
rect 1170 8700 1190 8980
rect 1290 8700 1310 8980
rect 1170 8620 1310 8700
rect 1170 8320 1190 8620
rect 1290 8320 1310 8620
rect 1170 8270 1310 8320
rect 1370 8980 1620 9030
rect 1370 8700 1390 8980
rect 1460 8700 1620 8980
rect 1370 8620 1620 8700
rect 1370 8320 1390 8620
rect 1460 8320 1620 8620
rect 1370 8270 1620 8320
rect 520 8250 1620 8270
rect 1440 8240 1620 8250
rect -1600 7740 -1580 7920
rect -20 7820 420 7920
rect -20 7810 1230 7820
rect -20 7750 580 7810
rect 1220 7750 1230 7810
rect -20 7740 1230 7750
rect -1600 7720 200 7740
rect 0 7580 200 7720
rect 1460 7640 1620 8240
rect -4200 6400 -200 7200
rect 0 7120 20 7580
rect 180 7120 200 7580
rect 10200 7580 11200 7600
rect 10200 7420 10220 7580
rect 10380 7420 11200 7580
rect 10200 7400 11200 7420
rect 0 7100 200 7120
rect -100 6480 200 6500
rect -100 6400 20 6480
rect -4200 6120 20 6400
rect 180 6120 200 6480
rect -4200 6000 200 6120
rect -8000 5800 200 6000
rect -1600 2400 200 5800
rect 11000 400 11200 7400
rect 10200 380 11200 400
rect 10200 220 10220 380
rect 10380 220 11200 380
rect 10200 200 11200 220
rect 11000 -200 11200 200
rect 9800 -300 11200 -200
rect 4000 -500 9000 -400
rect 4000 -3700 8500 -500
rect 8900 -3700 9000 -500
rect 9800 -700 9900 -300
rect 11100 -700 11200 -300
rect 9800 -800 11200 -700
rect 4000 -3800 9000 -3700
<< via3 >>
rect -1400 11800 800 12400
rect -7800 6000 -4200 8400
rect -1580 7740 -20 7920
rect 8500 -3700 8900 -500
rect 9900 -700 11100 -300
<< mimcap >>
rect -1560 11340 360 11360
rect -1560 8100 -1540 11340
rect 340 8100 360 11340
rect -1560 8080 360 8100
rect 4100 -600 7900 -500
rect 4100 -3600 4200 -600
rect 7800 -3600 7900 -600
rect 4100 -3700 7900 -3600
<< mimcapcontact >>
rect -1540 8100 340 11340
rect 4200 -3600 7800 -600
<< metal4 >>
rect -1600 12400 1000 20400
rect -1600 11800 -1400 12400
rect 800 11800 1000 12400
rect -1600 11600 1000 11800
rect -1600 11340 400 11400
rect -8000 8400 -4000 8600
rect -8000 6000 -7800 8400
rect -4200 6000 -4000 8400
rect -1600 8100 -1540 11340
rect 340 8100 400 11340
rect -1600 8020 400 8100
rect -1600 7920 0 7940
rect -1600 7740 -1580 7920
rect -20 7740 0 7920
rect -1600 7580 -1560 7740
rect -40 7580 0 7740
rect -1600 7540 0 7580
rect -8000 5800 -4000 6000
rect 10200 1800 17800 6000
rect 3700 -400 4400 400
rect 9800 -300 11200 -200
rect 3700 -600 8000 -400
rect 3700 -3400 4200 -600
rect 4000 -3600 4200 -3400
rect 7800 -3600 8000 -600
rect 4000 -3800 8000 -3600
rect 8400 -500 9000 -400
rect 8400 -3700 8500 -500
rect 8900 -3700 9000 -500
rect 9800 -1100 9900 -300
rect 11100 -1100 11200 -300
rect 9800 -1200 11200 -1100
rect 8400 -3800 9000 -3700
rect 11800 -17800 16400 1800
rect 11800 -41000 12000 -17800
rect 16200 -41000 16400 -17800
rect 11800 -41200 16400 -41000
<< via4 >>
rect -1400 11800 800 12400
rect -7800 6000 -4200 8400
rect -1560 7740 -40 7920
rect -1560 7580 -40 7740
rect 8500 -3700 8900 -500
rect 9900 -700 11100 -300
rect 9900 -1100 11100 -700
rect 12000 -41000 16200 -17800
<< mimcap2 >>
rect -1560 11340 360 11360
rect -1560 8100 -1540 11340
rect 340 8100 360 11340
rect -1560 8080 360 8100
rect 4100 -600 7900 -500
rect 4100 -3600 4200 -600
rect 7800 -3600 7900 -600
rect 4100 -3700 7900 -3600
<< mimcap2contact >>
rect -1540 8100 340 11340
rect 4200 -3600 7800 -600
<< metal5 >>
rect -23000 47000 17000 48000
rect -23000 16000 -22000 47000
rect 16000 33000 17000 47000
rect 16000 32000 71000 33000
rect -1600 18400 1000 21000
rect -1600 12400 1000 12600
rect -1600 11800 -1400 12400
rect 800 11800 1000 12400
rect -1600 11400 1000 11800
rect -1600 11340 400 11400
rect -8000 8400 -4000 10600
rect -8000 6000 -7800 8400
rect -4200 6000 -4000 8400
rect -1600 8100 -1540 11340
rect 340 8100 400 11340
rect -1600 8020 400 8100
rect -1600 7920 0 8020
rect -1600 7580 -1560 7920
rect -40 7580 0 7920
rect 2400 7600 9800 9000
rect -1600 7540 0 7580
rect -8000 5800 -4000 6000
rect 70000 5000 71000 32000
rect 9000 -300 11200 -200
rect 9000 -400 9900 -300
rect 4000 -500 9900 -400
rect 4000 -600 8500 -500
rect 4000 -3600 4200 -600
rect 7800 -3600 8500 -600
rect 4000 -3700 8500 -3600
rect 8900 -1100 9900 -500
rect 11100 -1100 11200 -300
rect 8900 -1200 11200 -1100
rect 8900 -3700 9000 -1200
rect 4000 -3800 9000 -3700
rect 66000 -9000 71000 5000
rect 64000 -11000 71000 -9000
rect 11800 -17800 16400 -17600
rect 7000 -42000 8000 -26000
rect 11800 -41000 12000 -17800
rect 16200 -41000 16400 -17800
rect 70000 -26000 71000 -11000
rect 11800 -41200 16400 -41000
rect 20000 -27000 71000 -26000
rect 20000 -42000 21000 -27000
use PA_core_1  PA_core_1_0
timestamp 1660307541
transform 0 -1 10000 1 0 700
box -700 -500 7196 10000
use octa_ind_3t_140_160_flat  octa_ind_3t_140_160_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1660524083
transform 0 -1 -23000 1 0 47900
box -39300 -34000 -5300 -6000
use octa_ind_thick_1p8n_flat  octa_ind_thick_1p8n_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1659752630
transform -1 0 20600 0 -1 -16800
box -51300 -45000 3200 5000
use sky130_fd_pr__nfet_01v8_6H2JGK  sky130_fd_pr__nfet_01v8_6H2JGK_0
timestamp 1660448881
transform 1 0 951 0 1 8650
box -551 -1010 551 1010
use sky130_fd_pr__res_high_po_0p35_ZE2H5K  sky130_fd_pr__res_high_po_0p35_ZE2H5K_0
timestamp 1660277336
transform 1 0 101 0 1 6798
box -201 -898 201 898
<< labels >>
rlabel metal5 8000 -2400 9000 -400 1 VGATE_CAS
rlabel metal3 420 9480 1320 9560 1 IREF_L
<< end >>
