magic
tech sky130B
magscale 1 2
timestamp 1661738380
<< metal4 >>
rect -31600 -22112 -26600 -22000
rect -31600 -23888 -28488 -22112
rect -26712 -23888 -26600 -22112
rect -31600 -24000 -26600 -23888
<< via4 >>
rect -28488 -23888 -26712 -22112
<< metal5 >>
tri -27401 -12100 -25401 -10100 se
rect -25401 -12100 -17199 -10100
tri -17199 -12100 -15199 -10100 sw
tri -30048 -14747 -27401 -12100 se
tri -31200 -15899 -30048 -14747 se
rect -30048 -14929 -27401 -14747
tri -27401 -14929 -24572 -12100 nw
tri -18028 -14929 -15199 -12100 ne
tri -15199 -13899 -13400 -12100 sw
rect -15199 -14929 -13400 -13899
rect -30048 -15899 -29200 -14929
rect -31200 -25711 -29200 -15899
tri -29200 -16728 -27401 -14929 nw
tri -15199 -16728 -13400 -14929 ne
tri -13400 -15899 -11400 -13899 sw
rect -28600 -22112 -26600 -22000
rect -28600 -23888 -28488 -22112
rect -26712 -23888 -26600 -22112
rect -28600 -24862 -26600 -23888
tri -29200 -25711 -28600 -25111 sw
tri -28600 -25711 -27751 -24862 ne
rect -27751 -25711 -26600 -24862
rect -31200 -25939 -28600 -25711
tri -31200 -26862 -30277 -25939 ne
rect -30277 -26013 -28600 -25939
tri -28600 -26013 -28298 -25711 sw
tri -27751 -26013 -27449 -25711 ne
rect -27449 -26013 -26600 -25711
rect -30277 -26862 -28298 -26013
tri -28298 -26862 -27449 -26013 sw
tri -27449 -26862 -26600 -26013 ne
tri -26600 -26862 -23772 -24034 sw
tri -14438 -25072 -13400 -24034 se
rect -13400 -24862 -11400 -15899
rect -13400 -25072 -11649 -24862
tri -16228 -26862 -14438 -25072 se
rect -14438 -25111 -11649 -25072
tri -11649 -25111 -11400 -24862 nw
rect -14438 -25921 -12459 -25111
tri -12459 -25921 -11649 -25111 nw
tri -11610 -25921 -10800 -25111 se
rect -10800 -25921 -8800 -23800
rect -14438 -26770 -13308 -25921
tri -13308 -26770 -12459 -25921 nw
tri -12459 -26770 -11610 -25921 se
rect -11610 -25939 -8800 -25921
rect -14438 -26862 -13589 -26770
tri -30277 -29690 -27449 -26862 ne
tri -27449 -27711 -26600 -26862 sw
tri -26600 -27711 -25751 -26862 ne
rect -25751 -27711 -23772 -26862
rect -27449 -27900 -26600 -27711
tri -26600 -27900 -26411 -27711 sw
tri -25751 -27900 -25562 -27711 ne
rect -25562 -27900 -23772 -27711
tri -23772 -27900 -22734 -26862 sw
tri -17266 -27900 -16228 -26862 se
rect -16228 -27051 -13589 -26862
tri -13589 -27051 -13308 -26770 nw
tri -12740 -27051 -12459 -26770 se
rect -12459 -27051 -11610 -26770
rect -16228 -27900 -14438 -27051
tri -14438 -27900 -13589 -27051 nw
tri -13589 -27900 -12740 -27051 se
rect -12740 -27900 -11610 -27051
rect -27449 -28749 -26411 -27900
tri -26411 -28749 -25562 -27900 sw
tri -25562 -28749 -24713 -27900 ne
rect -24713 -28749 -15287 -27900
tri -15287 -28749 -14438 -27900 nw
tri -14438 -28749 -13589 -27900 se
rect -13589 -28749 -11610 -27900
tri -11610 -28749 -8800 -25939 nw
rect -27449 -28841 -25562 -28749
tri -25562 -28841 -25470 -28749 sw
tri -24713 -28841 -24621 -28749 ne
rect -24621 -28841 -15379 -28749
tri -15379 -28841 -15287 -28749 nw
tri -14530 -28841 -14438 -28749 se
rect -27449 -29690 -25470 -28841
tri -25470 -29690 -24621 -28841 sw
tri -24621 -29690 -23772 -28841 ne
rect -23772 -29690 -16228 -28841
tri -16228 -29690 -15379 -28841 nw
tri -15379 -29690 -14530 -28841 se
rect -14530 -29690 -14438 -28841
tri -27449 -32500 -24639 -29690 ne
rect -24639 -30500 -24621 -29690
tri -24621 -30500 -23811 -29690 sw
tri -23772 -29900 -23562 -29690 ne
rect -23562 -29900 -16438 -29690
tri -16438 -29900 -16228 -29690 nw
tri -16189 -30500 -15379 -29690 se
rect -15379 -30500 -14438 -29690
rect -24639 -31577 -14438 -30500
tri -14438 -31577 -11610 -28749 nw
rect -24639 -32500 -15361 -31577
tri -15361 -32500 -14438 -31577 nw
<< comment >>
rect -33800 -18000 -33700 -17900
rect -31900 -18000 -31800 -17900
<< end >>
