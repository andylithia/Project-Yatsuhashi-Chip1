magic
tech sky130A
magscale 1 2
timestamp 1658291242
<< pwell >>
rect -612 -719 612 719
<< nmos >>
rect -416 109 -296 509
rect -238 109 -118 509
rect -60 109 60 509
rect 118 109 238 509
rect 296 109 416 509
rect -416 -509 -296 -109
rect -238 -509 -118 -109
rect -60 -509 60 -109
rect 118 -509 238 -109
rect 296 -509 416 -109
<< ndiff >>
rect -474 497 -416 509
rect -474 121 -462 497
rect -428 121 -416 497
rect -474 109 -416 121
rect -296 497 -238 509
rect -296 121 -284 497
rect -250 121 -238 497
rect -296 109 -238 121
rect -118 497 -60 509
rect -118 121 -106 497
rect -72 121 -60 497
rect -118 109 -60 121
rect 60 497 118 509
rect 60 121 72 497
rect 106 121 118 497
rect 60 109 118 121
rect 238 497 296 509
rect 238 121 250 497
rect 284 121 296 497
rect 238 109 296 121
rect 416 497 474 509
rect 416 121 428 497
rect 462 121 474 497
rect 416 109 474 121
rect -474 -121 -416 -109
rect -474 -497 -462 -121
rect -428 -497 -416 -121
rect -474 -509 -416 -497
rect -296 -121 -238 -109
rect -296 -497 -284 -121
rect -250 -497 -238 -121
rect -296 -509 -238 -497
rect -118 -121 -60 -109
rect -118 -497 -106 -121
rect -72 -497 -60 -121
rect -118 -509 -60 -497
rect 60 -121 118 -109
rect 60 -497 72 -121
rect 106 -497 118 -121
rect 60 -509 118 -497
rect 238 -121 296 -109
rect 238 -497 250 -121
rect 284 -497 296 -121
rect 238 -509 296 -497
rect 416 -121 474 -109
rect 416 -497 428 -121
rect 462 -497 474 -121
rect 416 -509 474 -497
<< ndiffc >>
rect -462 121 -428 497
rect -284 121 -250 497
rect -106 121 -72 497
rect 72 121 106 497
rect 250 121 284 497
rect 428 121 462 497
rect -462 -497 -428 -121
rect -284 -497 -250 -121
rect -106 -497 -72 -121
rect 72 -497 106 -121
rect 250 -497 284 -121
rect 428 -497 462 -121
<< psubdiff >>
rect -576 649 -480 683
rect 480 649 576 683
rect -576 587 -542 649
rect 542 587 576 649
rect -576 -649 -542 -587
rect 542 -649 576 -587
rect -576 -683 -480 -649
rect 480 -683 576 -649
<< psubdiffcont >>
rect -480 649 480 683
rect -576 -587 -542 587
rect 542 -587 576 587
rect -480 -683 480 -649
<< poly >>
rect -416 581 -296 597
rect -416 547 -400 581
rect -312 547 -296 581
rect -416 509 -296 547
rect -238 581 -118 597
rect -238 547 -222 581
rect -134 547 -118 581
rect -238 509 -118 547
rect -60 581 60 597
rect -60 547 -44 581
rect 44 547 60 581
rect -60 509 60 547
rect 118 581 238 597
rect 118 547 134 581
rect 222 547 238 581
rect 118 509 238 547
rect 296 581 416 597
rect 296 547 312 581
rect 400 547 416 581
rect 296 509 416 547
rect -416 71 -296 109
rect -416 37 -400 71
rect -312 37 -296 71
rect -416 21 -296 37
rect -238 71 -118 109
rect -238 37 -222 71
rect -134 37 -118 71
rect -238 21 -118 37
rect -60 71 60 109
rect -60 37 -44 71
rect 44 37 60 71
rect -60 21 60 37
rect 118 71 238 109
rect 118 37 134 71
rect 222 37 238 71
rect 118 21 238 37
rect 296 71 416 109
rect 296 37 312 71
rect 400 37 416 71
rect 296 21 416 37
rect -416 -37 -296 -21
rect -416 -71 -400 -37
rect -312 -71 -296 -37
rect -416 -109 -296 -71
rect -238 -37 -118 -21
rect -238 -71 -222 -37
rect -134 -71 -118 -37
rect -238 -109 -118 -71
rect -60 -37 60 -21
rect -60 -71 -44 -37
rect 44 -71 60 -37
rect -60 -109 60 -71
rect 118 -37 238 -21
rect 118 -71 134 -37
rect 222 -71 238 -37
rect 118 -109 238 -71
rect 296 -37 416 -21
rect 296 -71 312 -37
rect 400 -71 416 -37
rect 296 -109 416 -71
rect -416 -547 -296 -509
rect -416 -581 -400 -547
rect -312 -581 -296 -547
rect -416 -597 -296 -581
rect -238 -547 -118 -509
rect -238 -581 -222 -547
rect -134 -581 -118 -547
rect -238 -597 -118 -581
rect -60 -547 60 -509
rect -60 -581 -44 -547
rect 44 -581 60 -547
rect -60 -597 60 -581
rect 118 -547 238 -509
rect 118 -581 134 -547
rect 222 -581 238 -547
rect 118 -597 238 -581
rect 296 -547 416 -509
rect 296 -581 312 -547
rect 400 -581 416 -547
rect 296 -597 416 -581
<< polycont >>
rect -400 547 -312 581
rect -222 547 -134 581
rect -44 547 44 581
rect 134 547 222 581
rect 312 547 400 581
rect -400 37 -312 71
rect -222 37 -134 71
rect -44 37 44 71
rect 134 37 222 71
rect 312 37 400 71
rect -400 -71 -312 -37
rect -222 -71 -134 -37
rect -44 -71 44 -37
rect 134 -71 222 -37
rect 312 -71 400 -37
rect -400 -581 -312 -547
rect -222 -581 -134 -547
rect -44 -581 44 -547
rect 134 -581 222 -547
rect 312 -581 400 -547
<< locali >>
rect -576 649 -480 683
rect 480 649 576 683
rect -576 587 -542 649
rect 542 587 576 649
rect -416 547 -400 581
rect -312 547 -296 581
rect -238 547 -222 581
rect -134 547 -118 581
rect -60 547 -44 581
rect 44 547 60 581
rect 118 547 134 581
rect 222 547 238 581
rect 296 547 312 581
rect 400 547 416 581
rect -462 497 -428 513
rect -462 105 -428 121
rect -284 497 -250 513
rect -284 105 -250 121
rect -106 497 -72 513
rect -106 105 -72 121
rect 72 497 106 513
rect 72 105 106 121
rect 250 497 284 513
rect 250 105 284 121
rect 428 497 462 513
rect 428 105 462 121
rect -416 37 -400 71
rect -312 37 -296 71
rect -238 37 -222 71
rect -134 37 -118 71
rect -60 37 -44 71
rect 44 37 60 71
rect 118 37 134 71
rect 222 37 238 71
rect 296 37 312 71
rect 400 37 416 71
rect -416 -71 -400 -37
rect -312 -71 -296 -37
rect -238 -71 -222 -37
rect -134 -71 -118 -37
rect -60 -71 -44 -37
rect 44 -71 60 -37
rect 118 -71 134 -37
rect 222 -71 238 -37
rect 296 -71 312 -37
rect 400 -71 416 -37
rect -462 -121 -428 -105
rect -462 -513 -428 -497
rect -284 -121 -250 -105
rect -284 -513 -250 -497
rect -106 -121 -72 -105
rect -106 -513 -72 -497
rect 72 -121 106 -105
rect 72 -513 106 -497
rect 250 -121 284 -105
rect 250 -513 284 -497
rect 428 -121 462 -105
rect 428 -513 462 -497
rect -416 -581 -400 -547
rect -312 -581 -296 -547
rect -238 -581 -222 -547
rect -134 -581 -118 -547
rect -60 -581 -44 -547
rect 44 -581 60 -547
rect 118 -581 134 -547
rect 222 -581 238 -547
rect 296 -581 312 -547
rect 400 -581 416 -547
rect -576 -649 -542 -587
rect 542 -649 576 -587
rect -576 -683 -480 -649
rect 480 -683 576 -649
<< viali >>
rect -400 547 -312 581
rect -222 547 -134 581
rect -44 547 44 581
rect 134 547 222 581
rect 312 547 400 581
rect -462 121 -428 497
rect -284 121 -250 497
rect -106 121 -72 497
rect 72 121 106 497
rect 250 121 284 497
rect 428 121 462 497
rect -400 37 -312 71
rect -222 37 -134 71
rect -44 37 44 71
rect 134 37 222 71
rect 312 37 400 71
rect -400 -71 -312 -37
rect -222 -71 -134 -37
rect -44 -71 44 -37
rect 134 -71 222 -37
rect 312 -71 400 -37
rect -462 -497 -428 -121
rect -284 -497 -250 -121
rect -106 -497 -72 -121
rect 72 -497 106 -121
rect 250 -497 284 -121
rect 428 -497 462 -121
rect -400 -581 -312 -547
rect -222 -581 -134 -547
rect -44 -581 44 -547
rect 134 -581 222 -547
rect 312 -581 400 -547
<< metal1 >>
rect -412 581 -300 587
rect -412 547 -400 581
rect -312 547 -300 581
rect -412 541 -300 547
rect -234 581 -122 587
rect -234 547 -222 581
rect -134 547 -122 581
rect -234 541 -122 547
rect -56 581 56 587
rect -56 547 -44 581
rect 44 547 56 581
rect -56 541 56 547
rect 122 581 234 587
rect 122 547 134 581
rect 222 547 234 581
rect 122 541 234 547
rect 300 581 412 587
rect 300 547 312 581
rect 400 547 412 581
rect 300 541 412 547
rect -468 497 -422 509
rect -468 121 -462 497
rect -428 121 -422 497
rect -468 109 -422 121
rect -290 497 -244 509
rect -290 121 -284 497
rect -250 121 -244 497
rect -290 109 -244 121
rect -112 497 -66 509
rect -112 121 -106 497
rect -72 121 -66 497
rect -112 109 -66 121
rect 66 497 112 509
rect 66 121 72 497
rect 106 121 112 497
rect 66 109 112 121
rect 244 497 290 509
rect 244 121 250 497
rect 284 121 290 497
rect 244 109 290 121
rect 422 497 468 509
rect 422 121 428 497
rect 462 121 468 497
rect 422 109 468 121
rect -412 71 -300 77
rect -412 37 -400 71
rect -312 37 -300 71
rect -412 31 -300 37
rect -234 71 -122 77
rect -234 37 -222 71
rect -134 37 -122 71
rect -234 31 -122 37
rect -56 71 56 77
rect -56 37 -44 71
rect 44 37 56 71
rect -56 31 56 37
rect 122 71 234 77
rect 122 37 134 71
rect 222 37 234 71
rect 122 31 234 37
rect 300 71 412 77
rect 300 37 312 71
rect 400 37 412 71
rect 300 31 412 37
rect -412 -37 -300 -31
rect -412 -71 -400 -37
rect -312 -71 -300 -37
rect -412 -77 -300 -71
rect -234 -37 -122 -31
rect -234 -71 -222 -37
rect -134 -71 -122 -37
rect -234 -77 -122 -71
rect -56 -37 56 -31
rect -56 -71 -44 -37
rect 44 -71 56 -37
rect -56 -77 56 -71
rect 122 -37 234 -31
rect 122 -71 134 -37
rect 222 -71 234 -37
rect 122 -77 234 -71
rect 300 -37 412 -31
rect 300 -71 312 -37
rect 400 -71 412 -37
rect 300 -77 412 -71
rect -468 -121 -422 -109
rect -468 -497 -462 -121
rect -428 -497 -422 -121
rect -468 -509 -422 -497
rect -290 -121 -244 -109
rect -290 -497 -284 -121
rect -250 -497 -244 -121
rect -290 -509 -244 -497
rect -112 -121 -66 -109
rect -112 -497 -106 -121
rect -72 -497 -66 -121
rect -112 -509 -66 -497
rect 66 -121 112 -109
rect 66 -497 72 -121
rect 106 -497 112 -121
rect 66 -509 112 -497
rect 244 -121 290 -109
rect 244 -497 250 -121
rect 284 -497 290 -121
rect 244 -509 290 -497
rect 422 -121 468 -109
rect 422 -497 428 -121
rect 462 -497 468 -121
rect 422 -509 468 -497
rect -412 -547 -300 -541
rect -412 -581 -400 -547
rect -312 -581 -300 -547
rect -412 -587 -300 -581
rect -234 -547 -122 -541
rect -234 -581 -222 -547
rect -134 -581 -122 -547
rect -234 -587 -122 -581
rect -56 -547 56 -541
rect -56 -581 -44 -547
rect 44 -581 56 -547
rect -56 -587 56 -581
rect 122 -547 234 -541
rect 122 -581 134 -547
rect 222 -581 234 -547
rect 122 -587 234 -581
rect 300 -547 412 -541
rect 300 -581 312 -547
rect 400 -581 412 -547
rect 300 -587 412 -581
<< properties >>
string FIXED_BBOX -559 -666 559 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.6 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
