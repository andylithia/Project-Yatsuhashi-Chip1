magic
tech sky130B
magscale 1 2
timestamp 1659903400
<< nwell >>
rect -140 -920 2560 2380
<< pmos >>
rect 94 1912 154 2112
rect 334 1912 394 2112
rect 574 1912 634 2112
rect 814 1912 874 2112
rect 1054 1912 1114 2112
rect 1294 1912 1354 2112
rect 1534 1912 1594 2112
rect 1774 1912 1834 2112
rect 2014 1912 2074 2112
rect 2254 1912 2314 2112
rect 94 1542 154 1742
rect 334 1542 394 1742
rect 574 1542 634 1742
rect 814 1542 874 1742
rect 1054 1542 1114 1742
rect 1294 1542 1354 1742
rect 1534 1542 1594 1742
rect 1774 1542 1834 1742
rect 2014 1542 2074 1742
rect 2254 1542 2314 1742
rect 94 1172 154 1372
rect 334 1172 394 1372
rect 574 1172 634 1372
rect 814 1172 874 1372
rect 1054 1172 1114 1372
rect 1294 1172 1354 1372
rect 1534 1172 1594 1372
rect 1774 1172 1834 1372
rect 2014 1172 2074 1372
rect 2254 1172 2314 1372
rect 94 802 154 1002
rect 334 802 394 1002
rect 574 802 634 1002
rect 814 802 874 1002
rect 1054 802 1114 1002
rect 1294 802 1354 1002
rect 1534 802 1594 1002
rect 1774 802 1834 1002
rect 2014 802 2074 1002
rect 2254 802 2314 1002
rect 94 478 154 678
rect 334 478 394 678
rect 574 478 634 678
rect 814 478 874 678
rect 1054 478 1114 678
rect 1294 478 1354 678
rect 1534 478 1594 678
rect 1774 478 1834 678
rect 2014 478 2074 678
rect 2254 478 2314 678
rect 94 108 154 308
rect 334 108 394 308
rect 574 108 634 308
rect 814 108 874 308
rect 1054 108 1114 308
rect 1294 108 1354 308
rect 1534 108 1594 308
rect 1774 108 1834 308
rect 2014 108 2074 308
rect 2254 108 2314 308
rect 94 -262 154 -62
rect 334 -262 394 -62
rect 574 -262 634 -62
rect 814 -262 874 -62
rect 1054 -262 1114 -62
rect 1294 -262 1354 -62
rect 1534 -262 1594 -62
rect 1774 -262 1834 -62
rect 2014 -262 2074 -62
rect 2254 -262 2314 -62
rect 94 -632 154 -432
rect 334 -632 394 -432
rect 574 -632 634 -432
rect 814 -632 874 -432
rect 1054 -632 1114 -432
rect 1294 -632 1354 -432
rect 1534 -632 1594 -432
rect 1774 -632 1834 -432
rect 2014 -632 2074 -432
rect 2254 -632 2314 -432
<< pdiff >>
rect 36 2100 94 2112
rect 36 1924 48 2100
rect 82 1924 94 2100
rect 36 1912 94 1924
rect 154 2100 212 2112
rect 154 1924 166 2100
rect 200 1924 212 2100
rect 154 1912 212 1924
rect 276 2100 334 2112
rect 276 1924 288 2100
rect 322 1924 334 2100
rect 276 1912 334 1924
rect 394 2100 452 2112
rect 394 1924 406 2100
rect 440 1924 452 2100
rect 394 1912 452 1924
rect 516 2100 574 2112
rect 516 1924 528 2100
rect 562 1924 574 2100
rect 516 1912 574 1924
rect 634 2100 692 2112
rect 634 1924 646 2100
rect 680 1924 692 2100
rect 634 1912 692 1924
rect 756 2100 814 2112
rect 756 1924 768 2100
rect 802 1924 814 2100
rect 756 1912 814 1924
rect 874 2100 932 2112
rect 874 1924 886 2100
rect 920 1924 932 2100
rect 874 1912 932 1924
rect 996 2100 1054 2112
rect 996 1924 1008 2100
rect 1042 1924 1054 2100
rect 996 1912 1054 1924
rect 1114 2100 1172 2112
rect 1114 1924 1126 2100
rect 1160 1924 1172 2100
rect 1114 1912 1172 1924
rect 1236 2100 1294 2112
rect 1236 1924 1248 2100
rect 1282 1924 1294 2100
rect 1236 1912 1294 1924
rect 1354 2100 1412 2112
rect 1354 1924 1366 2100
rect 1400 1924 1412 2100
rect 1354 1912 1412 1924
rect 1476 2100 1534 2112
rect 1476 1924 1488 2100
rect 1522 1924 1534 2100
rect 1476 1912 1534 1924
rect 1594 2100 1652 2112
rect 1594 1924 1606 2100
rect 1640 1924 1652 2100
rect 1594 1912 1652 1924
rect 1716 2100 1774 2112
rect 1716 1924 1728 2100
rect 1762 1924 1774 2100
rect 1716 1912 1774 1924
rect 1834 2100 1892 2112
rect 1834 1924 1846 2100
rect 1880 1924 1892 2100
rect 1834 1912 1892 1924
rect 1956 2100 2014 2112
rect 1956 1924 1968 2100
rect 2002 1924 2014 2100
rect 1956 1912 2014 1924
rect 2074 2100 2132 2112
rect 2074 1924 2086 2100
rect 2120 1924 2132 2100
rect 2074 1912 2132 1924
rect 2196 2100 2254 2112
rect 2196 1924 2208 2100
rect 2242 1924 2254 2100
rect 2196 1912 2254 1924
rect 2314 2100 2372 2112
rect 2314 1924 2326 2100
rect 2360 1924 2372 2100
rect 2314 1912 2372 1924
rect 36 1730 94 1742
rect 36 1554 48 1730
rect 82 1554 94 1730
rect 36 1542 94 1554
rect 154 1730 212 1742
rect 154 1554 166 1730
rect 200 1554 212 1730
rect 154 1542 212 1554
rect 276 1730 334 1742
rect 276 1554 288 1730
rect 322 1554 334 1730
rect 276 1542 334 1554
rect 394 1730 452 1742
rect 394 1554 406 1730
rect 440 1554 452 1730
rect 394 1542 452 1554
rect 516 1730 574 1742
rect 516 1554 528 1730
rect 562 1554 574 1730
rect 516 1542 574 1554
rect 634 1730 692 1742
rect 634 1554 646 1730
rect 680 1554 692 1730
rect 634 1542 692 1554
rect 756 1730 814 1742
rect 756 1554 768 1730
rect 802 1554 814 1730
rect 756 1542 814 1554
rect 874 1730 932 1742
rect 874 1554 886 1730
rect 920 1554 932 1730
rect 874 1542 932 1554
rect 996 1730 1054 1742
rect 996 1554 1008 1730
rect 1042 1554 1054 1730
rect 996 1542 1054 1554
rect 1114 1730 1172 1742
rect 1114 1554 1126 1730
rect 1160 1554 1172 1730
rect 1114 1542 1172 1554
rect 1236 1730 1294 1742
rect 1236 1554 1248 1730
rect 1282 1554 1294 1730
rect 1236 1542 1294 1554
rect 1354 1730 1412 1742
rect 1354 1554 1366 1730
rect 1400 1554 1412 1730
rect 1354 1542 1412 1554
rect 1476 1730 1534 1742
rect 1476 1554 1488 1730
rect 1522 1554 1534 1730
rect 1476 1542 1534 1554
rect 1594 1730 1652 1742
rect 1594 1554 1606 1730
rect 1640 1554 1652 1730
rect 1594 1542 1652 1554
rect 1716 1730 1774 1742
rect 1716 1554 1728 1730
rect 1762 1554 1774 1730
rect 1716 1542 1774 1554
rect 1834 1730 1892 1742
rect 1834 1554 1846 1730
rect 1880 1554 1892 1730
rect 1834 1542 1892 1554
rect 1956 1730 2014 1742
rect 1956 1554 1968 1730
rect 2002 1554 2014 1730
rect 1956 1542 2014 1554
rect 2074 1730 2132 1742
rect 2074 1554 2086 1730
rect 2120 1554 2132 1730
rect 2074 1542 2132 1554
rect 2196 1730 2254 1742
rect 2196 1554 2208 1730
rect 2242 1554 2254 1730
rect 2196 1542 2254 1554
rect 2314 1730 2372 1742
rect 2314 1554 2326 1730
rect 2360 1554 2372 1730
rect 2314 1542 2372 1554
rect 36 1360 94 1372
rect 36 1184 48 1360
rect 82 1184 94 1360
rect 36 1172 94 1184
rect 154 1360 212 1372
rect 154 1184 166 1360
rect 200 1184 212 1360
rect 154 1172 212 1184
rect 276 1360 334 1372
rect 276 1184 288 1360
rect 322 1184 334 1360
rect 276 1172 334 1184
rect 394 1360 452 1372
rect 394 1184 406 1360
rect 440 1184 452 1360
rect 394 1172 452 1184
rect 516 1360 574 1372
rect 516 1184 528 1360
rect 562 1184 574 1360
rect 516 1172 574 1184
rect 634 1360 692 1372
rect 634 1184 646 1360
rect 680 1184 692 1360
rect 634 1172 692 1184
rect 756 1360 814 1372
rect 756 1184 768 1360
rect 802 1184 814 1360
rect 756 1172 814 1184
rect 874 1360 932 1372
rect 874 1184 886 1360
rect 920 1184 932 1360
rect 874 1172 932 1184
rect 996 1360 1054 1372
rect 996 1184 1008 1360
rect 1042 1184 1054 1360
rect 996 1172 1054 1184
rect 1114 1360 1172 1372
rect 1114 1184 1126 1360
rect 1160 1184 1172 1360
rect 1114 1172 1172 1184
rect 1236 1360 1294 1372
rect 1236 1184 1248 1360
rect 1282 1184 1294 1360
rect 1236 1172 1294 1184
rect 1354 1360 1412 1372
rect 1354 1184 1366 1360
rect 1400 1184 1412 1360
rect 1354 1172 1412 1184
rect 1476 1360 1534 1372
rect 1476 1184 1488 1360
rect 1522 1184 1534 1360
rect 1476 1172 1534 1184
rect 1594 1360 1652 1372
rect 1594 1184 1606 1360
rect 1640 1184 1652 1360
rect 1594 1172 1652 1184
rect 1716 1360 1774 1372
rect 1716 1184 1728 1360
rect 1762 1184 1774 1360
rect 1716 1172 1774 1184
rect 1834 1360 1892 1372
rect 1834 1184 1846 1360
rect 1880 1184 1892 1360
rect 1834 1172 1892 1184
rect 1956 1360 2014 1372
rect 1956 1184 1968 1360
rect 2002 1184 2014 1360
rect 1956 1172 2014 1184
rect 2074 1360 2132 1372
rect 2074 1184 2086 1360
rect 2120 1184 2132 1360
rect 2074 1172 2132 1184
rect 2196 1360 2254 1372
rect 2196 1184 2208 1360
rect 2242 1184 2254 1360
rect 2196 1172 2254 1184
rect 2314 1360 2372 1372
rect 2314 1184 2326 1360
rect 2360 1184 2372 1360
rect 2314 1172 2372 1184
rect 36 990 94 1002
rect 36 814 48 990
rect 82 814 94 990
rect 36 802 94 814
rect 154 990 212 1002
rect 154 814 166 990
rect 200 814 212 990
rect 154 802 212 814
rect 276 990 334 1002
rect 276 814 288 990
rect 322 814 334 990
rect 276 802 334 814
rect 394 990 452 1002
rect 394 814 406 990
rect 440 814 452 990
rect 394 802 452 814
rect 516 990 574 1002
rect 516 814 528 990
rect 562 814 574 990
rect 516 802 574 814
rect 634 990 692 1002
rect 634 814 646 990
rect 680 814 692 990
rect 634 802 692 814
rect 756 990 814 1002
rect 756 814 768 990
rect 802 814 814 990
rect 756 802 814 814
rect 874 990 932 1002
rect 874 814 886 990
rect 920 814 932 990
rect 874 802 932 814
rect 996 990 1054 1002
rect 996 814 1008 990
rect 1042 814 1054 990
rect 996 802 1054 814
rect 1114 990 1172 1002
rect 1114 814 1126 990
rect 1160 814 1172 990
rect 1114 802 1172 814
rect 1236 990 1294 1002
rect 1236 814 1248 990
rect 1282 814 1294 990
rect 1236 802 1294 814
rect 1354 990 1412 1002
rect 1354 814 1366 990
rect 1400 814 1412 990
rect 1354 802 1412 814
rect 1476 990 1534 1002
rect 1476 814 1488 990
rect 1522 814 1534 990
rect 1476 802 1534 814
rect 1594 990 1652 1002
rect 1594 814 1606 990
rect 1640 814 1652 990
rect 1594 802 1652 814
rect 1716 990 1774 1002
rect 1716 814 1728 990
rect 1762 814 1774 990
rect 1716 802 1774 814
rect 1834 990 1892 1002
rect 1834 814 1846 990
rect 1880 814 1892 990
rect 1834 802 1892 814
rect 1956 990 2014 1002
rect 1956 814 1968 990
rect 2002 814 2014 990
rect 1956 802 2014 814
rect 2074 990 2132 1002
rect 2074 814 2086 990
rect 2120 814 2132 990
rect 2074 802 2132 814
rect 2196 990 2254 1002
rect 2196 814 2208 990
rect 2242 814 2254 990
rect 2196 802 2254 814
rect 2314 990 2372 1002
rect 2314 814 2326 990
rect 2360 814 2372 990
rect 2314 802 2372 814
rect 36 666 94 678
rect 36 490 48 666
rect 82 490 94 666
rect 36 478 94 490
rect 154 666 212 678
rect 154 490 166 666
rect 200 490 212 666
rect 154 478 212 490
rect 276 666 334 678
rect 276 490 288 666
rect 322 490 334 666
rect 276 478 334 490
rect 394 666 452 678
rect 394 490 406 666
rect 440 490 452 666
rect 394 478 452 490
rect 516 666 574 678
rect 516 490 528 666
rect 562 490 574 666
rect 516 478 574 490
rect 634 666 692 678
rect 634 490 646 666
rect 680 490 692 666
rect 634 478 692 490
rect 756 666 814 678
rect 756 490 768 666
rect 802 490 814 666
rect 756 478 814 490
rect 874 666 932 678
rect 874 490 886 666
rect 920 490 932 666
rect 874 478 932 490
rect 996 666 1054 678
rect 996 490 1008 666
rect 1042 490 1054 666
rect 996 478 1054 490
rect 1114 666 1172 678
rect 1114 490 1126 666
rect 1160 490 1172 666
rect 1114 478 1172 490
rect 1236 666 1294 678
rect 1236 490 1248 666
rect 1282 490 1294 666
rect 1236 478 1294 490
rect 1354 666 1412 678
rect 1354 490 1366 666
rect 1400 490 1412 666
rect 1354 478 1412 490
rect 1476 666 1534 678
rect 1476 490 1488 666
rect 1522 490 1534 666
rect 1476 478 1534 490
rect 1594 666 1652 678
rect 1594 490 1606 666
rect 1640 490 1652 666
rect 1594 478 1652 490
rect 1716 666 1774 678
rect 1716 490 1728 666
rect 1762 490 1774 666
rect 1716 478 1774 490
rect 1834 666 1892 678
rect 1834 490 1846 666
rect 1880 490 1892 666
rect 1834 478 1892 490
rect 1956 666 2014 678
rect 1956 490 1968 666
rect 2002 490 2014 666
rect 1956 478 2014 490
rect 2074 666 2132 678
rect 2074 490 2086 666
rect 2120 490 2132 666
rect 2074 478 2132 490
rect 2196 666 2254 678
rect 2196 490 2208 666
rect 2242 490 2254 666
rect 2196 478 2254 490
rect 2314 666 2372 678
rect 2314 490 2326 666
rect 2360 490 2372 666
rect 2314 478 2372 490
rect 36 296 94 308
rect 36 120 48 296
rect 82 120 94 296
rect 36 108 94 120
rect 154 296 212 308
rect 154 120 166 296
rect 200 120 212 296
rect 154 108 212 120
rect 276 296 334 308
rect 276 120 288 296
rect 322 120 334 296
rect 276 108 334 120
rect 394 296 452 308
rect 394 120 406 296
rect 440 120 452 296
rect 394 108 452 120
rect 516 296 574 308
rect 516 120 528 296
rect 562 120 574 296
rect 516 108 574 120
rect 634 296 692 308
rect 634 120 646 296
rect 680 120 692 296
rect 634 108 692 120
rect 756 296 814 308
rect 756 120 768 296
rect 802 120 814 296
rect 756 108 814 120
rect 874 296 932 308
rect 874 120 886 296
rect 920 120 932 296
rect 874 108 932 120
rect 996 296 1054 308
rect 996 120 1008 296
rect 1042 120 1054 296
rect 996 108 1054 120
rect 1114 296 1172 308
rect 1114 120 1126 296
rect 1160 120 1172 296
rect 1114 108 1172 120
rect 1236 296 1294 308
rect 1236 120 1248 296
rect 1282 120 1294 296
rect 1236 108 1294 120
rect 1354 296 1412 308
rect 1354 120 1366 296
rect 1400 120 1412 296
rect 1354 108 1412 120
rect 1476 296 1534 308
rect 1476 120 1488 296
rect 1522 120 1534 296
rect 1476 108 1534 120
rect 1594 296 1652 308
rect 1594 120 1606 296
rect 1640 120 1652 296
rect 1594 108 1652 120
rect 1716 296 1774 308
rect 1716 120 1728 296
rect 1762 120 1774 296
rect 1716 108 1774 120
rect 1834 296 1892 308
rect 1834 120 1846 296
rect 1880 120 1892 296
rect 1834 108 1892 120
rect 1956 296 2014 308
rect 1956 120 1968 296
rect 2002 120 2014 296
rect 1956 108 2014 120
rect 2074 296 2132 308
rect 2074 120 2086 296
rect 2120 120 2132 296
rect 2074 108 2132 120
rect 2196 296 2254 308
rect 2196 120 2208 296
rect 2242 120 2254 296
rect 2196 108 2254 120
rect 2314 296 2372 308
rect 2314 120 2326 296
rect 2360 120 2372 296
rect 2314 108 2372 120
rect 36 -74 94 -62
rect 36 -250 48 -74
rect 82 -250 94 -74
rect 36 -262 94 -250
rect 154 -74 212 -62
rect 154 -250 166 -74
rect 200 -250 212 -74
rect 154 -262 212 -250
rect 276 -74 334 -62
rect 276 -250 288 -74
rect 322 -250 334 -74
rect 276 -262 334 -250
rect 394 -74 452 -62
rect 394 -250 406 -74
rect 440 -250 452 -74
rect 394 -262 452 -250
rect 516 -74 574 -62
rect 516 -250 528 -74
rect 562 -250 574 -74
rect 516 -262 574 -250
rect 634 -74 692 -62
rect 634 -250 646 -74
rect 680 -250 692 -74
rect 634 -262 692 -250
rect 756 -74 814 -62
rect 756 -250 768 -74
rect 802 -250 814 -74
rect 756 -262 814 -250
rect 874 -74 932 -62
rect 874 -250 886 -74
rect 920 -250 932 -74
rect 874 -262 932 -250
rect 996 -74 1054 -62
rect 996 -250 1008 -74
rect 1042 -250 1054 -74
rect 996 -262 1054 -250
rect 1114 -74 1172 -62
rect 1114 -250 1126 -74
rect 1160 -250 1172 -74
rect 1114 -262 1172 -250
rect 1236 -74 1294 -62
rect 1236 -250 1248 -74
rect 1282 -250 1294 -74
rect 1236 -262 1294 -250
rect 1354 -74 1412 -62
rect 1354 -250 1366 -74
rect 1400 -250 1412 -74
rect 1354 -262 1412 -250
rect 1476 -74 1534 -62
rect 1476 -250 1488 -74
rect 1522 -250 1534 -74
rect 1476 -262 1534 -250
rect 1594 -74 1652 -62
rect 1594 -250 1606 -74
rect 1640 -250 1652 -74
rect 1594 -262 1652 -250
rect 1716 -74 1774 -62
rect 1716 -250 1728 -74
rect 1762 -250 1774 -74
rect 1716 -262 1774 -250
rect 1834 -74 1892 -62
rect 1834 -250 1846 -74
rect 1880 -250 1892 -74
rect 1834 -262 1892 -250
rect 1956 -74 2014 -62
rect 1956 -250 1968 -74
rect 2002 -250 2014 -74
rect 1956 -262 2014 -250
rect 2074 -74 2132 -62
rect 2074 -250 2086 -74
rect 2120 -250 2132 -74
rect 2074 -262 2132 -250
rect 2196 -74 2254 -62
rect 2196 -250 2208 -74
rect 2242 -250 2254 -74
rect 2196 -262 2254 -250
rect 2314 -74 2372 -62
rect 2314 -250 2326 -74
rect 2360 -250 2372 -74
rect 2314 -262 2372 -250
rect 36 -444 94 -432
rect 36 -620 48 -444
rect 82 -620 94 -444
rect 36 -632 94 -620
rect 154 -444 212 -432
rect 154 -620 166 -444
rect 200 -620 212 -444
rect 154 -632 212 -620
rect 276 -444 334 -432
rect 276 -620 288 -444
rect 322 -620 334 -444
rect 276 -632 334 -620
rect 394 -444 452 -432
rect 394 -620 406 -444
rect 440 -620 452 -444
rect 394 -632 452 -620
rect 516 -444 574 -432
rect 516 -620 528 -444
rect 562 -620 574 -444
rect 516 -632 574 -620
rect 634 -444 692 -432
rect 634 -620 646 -444
rect 680 -620 692 -444
rect 634 -632 692 -620
rect 756 -444 814 -432
rect 756 -620 768 -444
rect 802 -620 814 -444
rect 756 -632 814 -620
rect 874 -444 932 -432
rect 874 -620 886 -444
rect 920 -620 932 -444
rect 874 -632 932 -620
rect 996 -444 1054 -432
rect 996 -620 1008 -444
rect 1042 -620 1054 -444
rect 996 -632 1054 -620
rect 1114 -444 1172 -432
rect 1114 -620 1126 -444
rect 1160 -620 1172 -444
rect 1114 -632 1172 -620
rect 1236 -444 1294 -432
rect 1236 -620 1248 -444
rect 1282 -620 1294 -444
rect 1236 -632 1294 -620
rect 1354 -444 1412 -432
rect 1354 -620 1366 -444
rect 1400 -620 1412 -444
rect 1354 -632 1412 -620
rect 1476 -444 1534 -432
rect 1476 -620 1488 -444
rect 1522 -620 1534 -444
rect 1476 -632 1534 -620
rect 1594 -444 1652 -432
rect 1594 -620 1606 -444
rect 1640 -620 1652 -444
rect 1594 -632 1652 -620
rect 1716 -444 1774 -432
rect 1716 -620 1728 -444
rect 1762 -620 1774 -444
rect 1716 -632 1774 -620
rect 1834 -444 1892 -432
rect 1834 -620 1846 -444
rect 1880 -620 1892 -444
rect 1834 -632 1892 -620
rect 1956 -444 2014 -432
rect 1956 -620 1968 -444
rect 2002 -620 2014 -444
rect 1956 -632 2014 -620
rect 2074 -444 2132 -432
rect 2074 -620 2086 -444
rect 2120 -620 2132 -444
rect 2074 -632 2132 -620
rect 2196 -444 2254 -432
rect 2196 -620 2208 -444
rect 2242 -620 2254 -444
rect 2196 -632 2254 -620
rect 2314 -444 2372 -432
rect 2314 -620 2326 -444
rect 2360 -620 2372 -444
rect 2314 -632 2372 -620
<< pdiffc >>
rect 48 1924 82 2100
rect 166 1924 200 2100
rect 288 1924 322 2100
rect 406 1924 440 2100
rect 528 1924 562 2100
rect 646 1924 680 2100
rect 768 1924 802 2100
rect 886 1924 920 2100
rect 1008 1924 1042 2100
rect 1126 1924 1160 2100
rect 1248 1924 1282 2100
rect 1366 1924 1400 2100
rect 1488 1924 1522 2100
rect 1606 1924 1640 2100
rect 1728 1924 1762 2100
rect 1846 1924 1880 2100
rect 1968 1924 2002 2100
rect 2086 1924 2120 2100
rect 2208 1924 2242 2100
rect 2326 1924 2360 2100
rect 48 1554 82 1730
rect 166 1554 200 1730
rect 288 1554 322 1730
rect 406 1554 440 1730
rect 528 1554 562 1730
rect 646 1554 680 1730
rect 768 1554 802 1730
rect 886 1554 920 1730
rect 1008 1554 1042 1730
rect 1126 1554 1160 1730
rect 1248 1554 1282 1730
rect 1366 1554 1400 1730
rect 1488 1554 1522 1730
rect 1606 1554 1640 1730
rect 1728 1554 1762 1730
rect 1846 1554 1880 1730
rect 1968 1554 2002 1730
rect 2086 1554 2120 1730
rect 2208 1554 2242 1730
rect 2326 1554 2360 1730
rect 48 1184 82 1360
rect 166 1184 200 1360
rect 288 1184 322 1360
rect 406 1184 440 1360
rect 528 1184 562 1360
rect 646 1184 680 1360
rect 768 1184 802 1360
rect 886 1184 920 1360
rect 1008 1184 1042 1360
rect 1126 1184 1160 1360
rect 1248 1184 1282 1360
rect 1366 1184 1400 1360
rect 1488 1184 1522 1360
rect 1606 1184 1640 1360
rect 1728 1184 1762 1360
rect 1846 1184 1880 1360
rect 1968 1184 2002 1360
rect 2086 1184 2120 1360
rect 2208 1184 2242 1360
rect 2326 1184 2360 1360
rect 48 814 82 990
rect 166 814 200 990
rect 288 814 322 990
rect 406 814 440 990
rect 528 814 562 990
rect 646 814 680 990
rect 768 814 802 990
rect 886 814 920 990
rect 1008 814 1042 990
rect 1126 814 1160 990
rect 1248 814 1282 990
rect 1366 814 1400 990
rect 1488 814 1522 990
rect 1606 814 1640 990
rect 1728 814 1762 990
rect 1846 814 1880 990
rect 1968 814 2002 990
rect 2086 814 2120 990
rect 2208 814 2242 990
rect 2326 814 2360 990
rect 48 490 82 666
rect 166 490 200 666
rect 288 490 322 666
rect 406 490 440 666
rect 528 490 562 666
rect 646 490 680 666
rect 768 490 802 666
rect 886 490 920 666
rect 1008 490 1042 666
rect 1126 490 1160 666
rect 1248 490 1282 666
rect 1366 490 1400 666
rect 1488 490 1522 666
rect 1606 490 1640 666
rect 1728 490 1762 666
rect 1846 490 1880 666
rect 1968 490 2002 666
rect 2086 490 2120 666
rect 2208 490 2242 666
rect 2326 490 2360 666
rect 48 120 82 296
rect 166 120 200 296
rect 288 120 322 296
rect 406 120 440 296
rect 528 120 562 296
rect 646 120 680 296
rect 768 120 802 296
rect 886 120 920 296
rect 1008 120 1042 296
rect 1126 120 1160 296
rect 1248 120 1282 296
rect 1366 120 1400 296
rect 1488 120 1522 296
rect 1606 120 1640 296
rect 1728 120 1762 296
rect 1846 120 1880 296
rect 1968 120 2002 296
rect 2086 120 2120 296
rect 2208 120 2242 296
rect 2326 120 2360 296
rect 48 -250 82 -74
rect 166 -250 200 -74
rect 288 -250 322 -74
rect 406 -250 440 -74
rect 528 -250 562 -74
rect 646 -250 680 -74
rect 768 -250 802 -74
rect 886 -250 920 -74
rect 1008 -250 1042 -74
rect 1126 -250 1160 -74
rect 1248 -250 1282 -74
rect 1366 -250 1400 -74
rect 1488 -250 1522 -74
rect 1606 -250 1640 -74
rect 1728 -250 1762 -74
rect 1846 -250 1880 -74
rect 1968 -250 2002 -74
rect 2086 -250 2120 -74
rect 2208 -250 2242 -74
rect 2326 -250 2360 -74
rect 48 -620 82 -444
rect 166 -620 200 -444
rect 288 -620 322 -444
rect 406 -620 440 -444
rect 528 -620 562 -444
rect 646 -620 680 -444
rect 768 -620 802 -444
rect 886 -620 920 -444
rect 1008 -620 1042 -444
rect 1126 -620 1160 -444
rect 1248 -620 1282 -444
rect 1366 -620 1400 -444
rect 1488 -620 1522 -444
rect 1606 -620 1640 -444
rect 1728 -620 1762 -444
rect 1846 -620 1880 -444
rect 1968 -620 2002 -444
rect 2086 -620 2120 -444
rect 2208 -620 2242 -444
rect 2326 -620 2360 -444
<< nsubdiff >>
rect -100 2300 2520 2340
rect -100 -840 -80 2300
rect -40 2240 2460 2260
rect -40 -780 -20 2240
rect 2440 -780 2460 2240
rect -40 -800 2460 -780
rect 2500 -840 2520 2300
rect -100 -880 2520 -840
<< nsubdiffcont >>
rect -80 2260 2500 2300
rect -80 -800 -40 2260
rect 2460 -800 2500 2260
rect -80 -840 2500 -800
<< poly >>
rect 91 2193 157 2209
rect 91 2159 107 2193
rect 141 2159 157 2193
rect 91 2143 157 2159
rect 331 2193 397 2209
rect 331 2159 347 2193
rect 381 2159 397 2193
rect 331 2143 397 2159
rect 571 2193 637 2209
rect 571 2159 587 2193
rect 621 2159 637 2193
rect 571 2143 637 2159
rect 811 2193 877 2209
rect 811 2159 827 2193
rect 861 2159 877 2193
rect 811 2143 877 2159
rect 1051 2193 1117 2209
rect 1051 2159 1067 2193
rect 1101 2159 1117 2193
rect 1051 2143 1117 2159
rect 1291 2193 1357 2209
rect 1291 2159 1307 2193
rect 1341 2159 1357 2193
rect 1291 2143 1357 2159
rect 1531 2193 1597 2209
rect 1531 2159 1547 2193
rect 1581 2159 1597 2193
rect 1531 2143 1597 2159
rect 1771 2193 1837 2209
rect 1771 2159 1787 2193
rect 1821 2159 1837 2193
rect 1771 2143 1837 2159
rect 2011 2193 2077 2209
rect 2011 2159 2027 2193
rect 2061 2159 2077 2193
rect 2011 2143 2077 2159
rect 2251 2193 2317 2209
rect 2251 2159 2267 2193
rect 2301 2159 2317 2193
rect 2251 2143 2317 2159
rect 94 2112 154 2143
rect 334 2112 394 2143
rect 574 2112 634 2143
rect 814 2112 874 2143
rect 1054 2112 1114 2143
rect 1294 2112 1354 2143
rect 1534 2112 1594 2143
rect 1774 2112 1834 2143
rect 2014 2112 2074 2143
rect 2254 2112 2314 2143
rect 94 1886 154 1912
rect 334 1886 394 1912
rect 574 1886 634 1912
rect 814 1886 874 1912
rect 1054 1886 1114 1912
rect 1294 1886 1354 1912
rect 1534 1886 1594 1912
rect 1774 1886 1834 1912
rect 2014 1886 2074 1912
rect 2254 1886 2314 1912
rect 91 1823 157 1839
rect 91 1789 107 1823
rect 141 1789 157 1823
rect 91 1773 157 1789
rect 331 1823 397 1839
rect 331 1789 347 1823
rect 381 1789 397 1823
rect 331 1773 397 1789
rect 571 1823 637 1839
rect 571 1789 587 1823
rect 621 1789 637 1823
rect 571 1773 637 1789
rect 811 1823 877 1839
rect 811 1789 827 1823
rect 861 1789 877 1823
rect 811 1773 877 1789
rect 1051 1823 1117 1839
rect 1051 1789 1067 1823
rect 1101 1789 1117 1823
rect 1051 1773 1117 1789
rect 1291 1823 1357 1839
rect 1291 1789 1307 1823
rect 1341 1789 1357 1823
rect 1291 1773 1357 1789
rect 1531 1823 1597 1839
rect 1531 1789 1547 1823
rect 1581 1789 1597 1823
rect 1531 1773 1597 1789
rect 1771 1823 1837 1839
rect 1771 1789 1787 1823
rect 1821 1789 1837 1823
rect 1771 1773 1837 1789
rect 2011 1823 2077 1839
rect 2011 1789 2027 1823
rect 2061 1789 2077 1823
rect 2011 1773 2077 1789
rect 2251 1823 2317 1839
rect 2251 1789 2267 1823
rect 2301 1789 2317 1823
rect 2251 1773 2317 1789
rect 94 1742 154 1773
rect 334 1742 394 1773
rect 574 1742 634 1773
rect 814 1742 874 1773
rect 1054 1742 1114 1773
rect 1294 1742 1354 1773
rect 1534 1742 1594 1773
rect 1774 1742 1834 1773
rect 2014 1742 2074 1773
rect 2254 1742 2314 1773
rect 94 1516 154 1542
rect 334 1516 394 1542
rect 574 1516 634 1542
rect 814 1516 874 1542
rect 1054 1516 1114 1542
rect 1294 1516 1354 1542
rect 1534 1516 1594 1542
rect 1774 1516 1834 1542
rect 2014 1516 2074 1542
rect 2254 1516 2314 1542
rect 91 1453 157 1469
rect 91 1419 107 1453
rect 141 1419 157 1453
rect 91 1403 157 1419
rect 331 1453 397 1469
rect 331 1419 347 1453
rect 381 1419 397 1453
rect 331 1403 397 1419
rect 571 1453 637 1469
rect 571 1419 587 1453
rect 621 1419 637 1453
rect 571 1403 637 1419
rect 811 1453 877 1469
rect 811 1419 827 1453
rect 861 1419 877 1453
rect 811 1403 877 1419
rect 1051 1453 1117 1469
rect 1051 1419 1067 1453
rect 1101 1419 1117 1453
rect 1051 1403 1117 1419
rect 1291 1453 1357 1469
rect 1291 1419 1307 1453
rect 1341 1419 1357 1453
rect 1291 1403 1357 1419
rect 1531 1453 1597 1469
rect 1531 1419 1547 1453
rect 1581 1419 1597 1453
rect 1531 1403 1597 1419
rect 1771 1453 1837 1469
rect 1771 1419 1787 1453
rect 1821 1419 1837 1453
rect 1771 1403 1837 1419
rect 2011 1453 2077 1469
rect 2011 1419 2027 1453
rect 2061 1419 2077 1453
rect 2011 1403 2077 1419
rect 2251 1453 2317 1469
rect 2251 1419 2267 1453
rect 2301 1419 2317 1453
rect 2251 1403 2317 1419
rect 94 1372 154 1403
rect 334 1372 394 1403
rect 574 1372 634 1403
rect 814 1372 874 1403
rect 1054 1372 1114 1403
rect 1294 1372 1354 1403
rect 1534 1372 1594 1403
rect 1774 1372 1834 1403
rect 2014 1372 2074 1403
rect 2254 1372 2314 1403
rect 94 1146 154 1172
rect 334 1146 394 1172
rect 574 1146 634 1172
rect 814 1146 874 1172
rect 1054 1146 1114 1172
rect 1294 1146 1354 1172
rect 1534 1146 1594 1172
rect 1774 1146 1834 1172
rect 2014 1146 2074 1172
rect 2254 1146 2314 1172
rect 91 1083 157 1099
rect 91 1049 107 1083
rect 141 1049 157 1083
rect 91 1033 157 1049
rect 331 1083 397 1099
rect 331 1049 347 1083
rect 381 1049 397 1083
rect 331 1033 397 1049
rect 571 1083 637 1099
rect 571 1049 587 1083
rect 621 1049 637 1083
rect 571 1033 637 1049
rect 811 1083 877 1099
rect 811 1049 827 1083
rect 861 1049 877 1083
rect 811 1033 877 1049
rect 1051 1083 1117 1099
rect 1051 1049 1067 1083
rect 1101 1049 1117 1083
rect 1051 1033 1117 1049
rect 1291 1083 1357 1099
rect 1291 1049 1307 1083
rect 1341 1049 1357 1083
rect 1291 1033 1357 1049
rect 1531 1083 1597 1099
rect 1531 1049 1547 1083
rect 1581 1049 1597 1083
rect 1531 1033 1597 1049
rect 1771 1083 1837 1099
rect 1771 1049 1787 1083
rect 1821 1049 1837 1083
rect 1771 1033 1837 1049
rect 2011 1083 2077 1099
rect 2011 1049 2027 1083
rect 2061 1049 2077 1083
rect 2011 1033 2077 1049
rect 2251 1083 2317 1099
rect 2251 1049 2267 1083
rect 2301 1049 2317 1083
rect 2251 1033 2317 1049
rect 94 1002 154 1033
rect 334 1002 394 1033
rect 574 1002 634 1033
rect 814 1002 874 1033
rect 1054 1002 1114 1033
rect 1294 1002 1354 1033
rect 1534 1002 1594 1033
rect 1774 1002 1834 1033
rect 2014 1002 2074 1033
rect 2254 1002 2314 1033
rect 94 776 154 802
rect 334 776 394 802
rect 574 776 634 802
rect 814 776 874 802
rect 1054 776 1114 802
rect 1294 776 1354 802
rect 1534 776 1594 802
rect 1774 776 1834 802
rect 2014 776 2074 802
rect 2254 776 2314 802
rect 94 678 154 704
rect 334 678 394 704
rect 574 678 634 704
rect 814 678 874 704
rect 1054 678 1114 704
rect 1294 678 1354 704
rect 1534 678 1594 704
rect 1774 678 1834 704
rect 2014 678 2074 704
rect 2254 678 2314 704
rect 94 447 154 478
rect 334 447 394 478
rect 574 447 634 478
rect 814 447 874 478
rect 1054 447 1114 478
rect 1294 447 1354 478
rect 1534 447 1594 478
rect 1774 447 1834 478
rect 2014 447 2074 478
rect 2254 447 2314 478
rect 91 431 157 447
rect 91 397 107 431
rect 141 397 157 431
rect 91 381 157 397
rect 331 431 397 447
rect 331 397 347 431
rect 381 397 397 431
rect 331 381 397 397
rect 571 431 637 447
rect 571 397 587 431
rect 621 397 637 431
rect 571 381 637 397
rect 811 431 877 447
rect 811 397 827 431
rect 861 397 877 431
rect 811 381 877 397
rect 1051 431 1117 447
rect 1051 397 1067 431
rect 1101 397 1117 431
rect 1051 381 1117 397
rect 1291 431 1357 447
rect 1291 397 1307 431
rect 1341 397 1357 431
rect 1291 381 1357 397
rect 1531 431 1597 447
rect 1531 397 1547 431
rect 1581 397 1597 431
rect 1531 381 1597 397
rect 1771 431 1837 447
rect 1771 397 1787 431
rect 1821 397 1837 431
rect 1771 381 1837 397
rect 2011 431 2077 447
rect 2011 397 2027 431
rect 2061 397 2077 431
rect 2011 381 2077 397
rect 2251 431 2317 447
rect 2251 397 2267 431
rect 2301 397 2317 431
rect 2251 381 2317 397
rect 94 308 154 334
rect 334 308 394 334
rect 574 308 634 334
rect 814 308 874 334
rect 1054 308 1114 334
rect 1294 308 1354 334
rect 1534 308 1594 334
rect 1774 308 1834 334
rect 2014 308 2074 334
rect 2254 308 2314 334
rect 94 77 154 108
rect 334 77 394 108
rect 574 77 634 108
rect 814 77 874 108
rect 1054 77 1114 108
rect 1294 77 1354 108
rect 1534 77 1594 108
rect 1774 77 1834 108
rect 2014 77 2074 108
rect 2254 77 2314 108
rect 91 61 157 77
rect 91 27 107 61
rect 141 27 157 61
rect 91 11 157 27
rect 331 61 397 77
rect 331 27 347 61
rect 381 27 397 61
rect 331 11 397 27
rect 571 61 637 77
rect 571 27 587 61
rect 621 27 637 61
rect 571 11 637 27
rect 811 61 877 77
rect 811 27 827 61
rect 861 27 877 61
rect 811 11 877 27
rect 1051 61 1117 77
rect 1051 27 1067 61
rect 1101 27 1117 61
rect 1051 11 1117 27
rect 1291 61 1357 77
rect 1291 27 1307 61
rect 1341 27 1357 61
rect 1291 11 1357 27
rect 1531 61 1597 77
rect 1531 27 1547 61
rect 1581 27 1597 61
rect 1531 11 1597 27
rect 1771 61 1837 77
rect 1771 27 1787 61
rect 1821 27 1837 61
rect 1771 11 1837 27
rect 2011 61 2077 77
rect 2011 27 2027 61
rect 2061 27 2077 61
rect 2011 11 2077 27
rect 2251 61 2317 77
rect 2251 27 2267 61
rect 2301 27 2317 61
rect 2251 11 2317 27
rect 94 -62 154 -36
rect 334 -62 394 -36
rect 574 -62 634 -36
rect 814 -62 874 -36
rect 1054 -62 1114 -36
rect 1294 -62 1354 -36
rect 1534 -62 1594 -36
rect 1774 -62 1834 -36
rect 2014 -62 2074 -36
rect 2254 -62 2314 -36
rect 94 -293 154 -262
rect 334 -293 394 -262
rect 574 -293 634 -262
rect 814 -293 874 -262
rect 1054 -293 1114 -262
rect 1294 -293 1354 -262
rect 1534 -293 1594 -262
rect 1774 -293 1834 -262
rect 2014 -293 2074 -262
rect 2254 -293 2314 -262
rect 91 -309 157 -293
rect 91 -343 107 -309
rect 141 -343 157 -309
rect 91 -359 157 -343
rect 331 -309 397 -293
rect 331 -343 347 -309
rect 381 -343 397 -309
rect 331 -359 397 -343
rect 571 -309 637 -293
rect 571 -343 587 -309
rect 621 -343 637 -309
rect 571 -359 637 -343
rect 811 -309 877 -293
rect 811 -343 827 -309
rect 861 -343 877 -309
rect 811 -359 877 -343
rect 1051 -309 1117 -293
rect 1051 -343 1067 -309
rect 1101 -343 1117 -309
rect 1051 -359 1117 -343
rect 1291 -309 1357 -293
rect 1291 -343 1307 -309
rect 1341 -343 1357 -309
rect 1291 -359 1357 -343
rect 1531 -309 1597 -293
rect 1531 -343 1547 -309
rect 1581 -343 1597 -309
rect 1531 -359 1597 -343
rect 1771 -309 1837 -293
rect 1771 -343 1787 -309
rect 1821 -343 1837 -309
rect 1771 -359 1837 -343
rect 2011 -309 2077 -293
rect 2011 -343 2027 -309
rect 2061 -343 2077 -309
rect 2011 -359 2077 -343
rect 2251 -309 2317 -293
rect 2251 -343 2267 -309
rect 2301 -343 2317 -309
rect 2251 -359 2317 -343
rect 94 -432 154 -406
rect 334 -432 394 -406
rect 574 -432 634 -406
rect 814 -432 874 -406
rect 1054 -432 1114 -406
rect 1294 -432 1354 -406
rect 1534 -432 1594 -406
rect 1774 -432 1834 -406
rect 2014 -432 2074 -406
rect 2254 -432 2314 -406
rect 94 -663 154 -632
rect 334 -663 394 -632
rect 574 -663 634 -632
rect 814 -663 874 -632
rect 1054 -663 1114 -632
rect 1294 -663 1354 -632
rect 1534 -663 1594 -632
rect 1774 -663 1834 -632
rect 2014 -663 2074 -632
rect 2254 -663 2314 -632
rect 91 -679 157 -663
rect 91 -713 107 -679
rect 141 -713 157 -679
rect 91 -729 157 -713
rect 331 -679 397 -663
rect 331 -713 347 -679
rect 381 -713 397 -679
rect 331 -729 397 -713
rect 571 -679 637 -663
rect 571 -713 587 -679
rect 621 -713 637 -679
rect 571 -729 637 -713
rect 811 -679 877 -663
rect 811 -713 827 -679
rect 861 -713 877 -679
rect 811 -729 877 -713
rect 1051 -679 1117 -663
rect 1051 -713 1067 -679
rect 1101 -713 1117 -679
rect 1051 -729 1117 -713
rect 1291 -679 1357 -663
rect 1291 -713 1307 -679
rect 1341 -713 1357 -679
rect 1291 -729 1357 -713
rect 1531 -679 1597 -663
rect 1531 -713 1547 -679
rect 1581 -713 1597 -679
rect 1531 -729 1597 -713
rect 1771 -679 1837 -663
rect 1771 -713 1787 -679
rect 1821 -713 1837 -679
rect 1771 -729 1837 -713
rect 2011 -679 2077 -663
rect 2011 -713 2027 -679
rect 2061 -713 2077 -679
rect 2011 -729 2077 -713
rect 2251 -679 2317 -663
rect 2251 -713 2267 -679
rect 2301 -713 2317 -679
rect 2251 -729 2317 -713
<< polycont >>
rect 107 2159 141 2193
rect 347 2159 381 2193
rect 587 2159 621 2193
rect 827 2159 861 2193
rect 1067 2159 1101 2193
rect 1307 2159 1341 2193
rect 1547 2159 1581 2193
rect 1787 2159 1821 2193
rect 2027 2159 2061 2193
rect 2267 2159 2301 2193
rect 107 1789 141 1823
rect 347 1789 381 1823
rect 587 1789 621 1823
rect 827 1789 861 1823
rect 1067 1789 1101 1823
rect 1307 1789 1341 1823
rect 1547 1789 1581 1823
rect 1787 1789 1821 1823
rect 2027 1789 2061 1823
rect 2267 1789 2301 1823
rect 107 1419 141 1453
rect 347 1419 381 1453
rect 587 1419 621 1453
rect 827 1419 861 1453
rect 1067 1419 1101 1453
rect 1307 1419 1341 1453
rect 1547 1419 1581 1453
rect 1787 1419 1821 1453
rect 2027 1419 2061 1453
rect 2267 1419 2301 1453
rect 107 1049 141 1083
rect 347 1049 381 1083
rect 587 1049 621 1083
rect 827 1049 861 1083
rect 1067 1049 1101 1083
rect 1307 1049 1341 1083
rect 1547 1049 1581 1083
rect 1787 1049 1821 1083
rect 2027 1049 2061 1083
rect 2267 1049 2301 1083
rect 107 397 141 431
rect 347 397 381 431
rect 587 397 621 431
rect 827 397 861 431
rect 1067 397 1101 431
rect 1307 397 1341 431
rect 1547 397 1581 431
rect 1787 397 1821 431
rect 2027 397 2061 431
rect 2267 397 2301 431
rect 107 27 141 61
rect 347 27 381 61
rect 587 27 621 61
rect 827 27 861 61
rect 1067 27 1101 61
rect 1307 27 1341 61
rect 1547 27 1581 61
rect 1787 27 1821 61
rect 2027 27 2061 61
rect 2267 27 2301 61
rect 107 -343 141 -309
rect 347 -343 381 -309
rect 587 -343 621 -309
rect 827 -343 861 -309
rect 1067 -343 1101 -309
rect 1307 -343 1341 -309
rect 1547 -343 1581 -309
rect 1787 -343 1821 -309
rect 2027 -343 2061 -309
rect 2267 -343 2301 -309
rect 107 -713 141 -679
rect 347 -713 381 -679
rect 587 -713 621 -679
rect 827 -713 861 -679
rect 1067 -713 1101 -679
rect 1307 -713 1341 -679
rect 1547 -713 1581 -679
rect 1787 -713 1821 -679
rect 2027 -713 2061 -679
rect 2267 -713 2301 -679
<< locali >>
rect -100 2300 2520 2320
rect -100 -840 -80 2300
rect -40 2240 2460 2260
rect -40 -780 -20 2240
rect 91 2159 107 2193
rect 141 2159 157 2193
rect 331 2159 347 2193
rect 381 2159 397 2193
rect 571 2159 587 2193
rect 621 2159 637 2193
rect 811 2159 827 2193
rect 861 2159 877 2193
rect 1051 2159 1067 2193
rect 1101 2159 1117 2193
rect 1291 2159 1307 2193
rect 1341 2159 1357 2193
rect 1531 2159 1547 2193
rect 1581 2159 1597 2193
rect 1771 2159 1787 2193
rect 1821 2159 1837 2193
rect 2011 2159 2027 2193
rect 2061 2159 2077 2193
rect 2251 2159 2267 2193
rect 2301 2159 2317 2193
rect 48 2100 82 2116
rect 48 1908 82 1924
rect 166 2100 200 2116
rect 166 1908 200 1924
rect 288 2100 322 2116
rect 288 1908 322 1924
rect 406 2100 440 2116
rect 406 1908 440 1924
rect 528 2100 562 2116
rect 528 1908 562 1924
rect 646 2100 680 2116
rect 646 1908 680 1924
rect 768 2100 802 2116
rect 768 1908 802 1924
rect 886 2100 920 2116
rect 886 1908 920 1924
rect 1008 2100 1042 2116
rect 1008 1908 1042 1924
rect 1126 2100 1160 2116
rect 1126 1908 1160 1924
rect 1248 2100 1282 2116
rect 1248 1908 1282 1924
rect 1366 2100 1400 2116
rect 1366 1908 1400 1924
rect 1488 2100 1522 2116
rect 1488 1908 1522 1924
rect 1606 2100 1640 2116
rect 1606 1908 1640 1924
rect 1728 2100 1762 2116
rect 1728 1908 1762 1924
rect 1846 2100 1880 2116
rect 1846 1908 1880 1924
rect 1968 2100 2002 2116
rect 1968 1908 2002 1924
rect 2086 2100 2120 2116
rect 2086 1908 2120 1924
rect 2208 2100 2242 2116
rect 2208 1908 2242 1924
rect 2326 2100 2360 2116
rect 2326 1908 2360 1924
rect 91 1789 107 1823
rect 141 1789 157 1823
rect 331 1789 347 1823
rect 381 1789 397 1823
rect 571 1789 587 1823
rect 621 1789 637 1823
rect 811 1789 827 1823
rect 861 1789 877 1823
rect 1051 1789 1067 1823
rect 1101 1789 1117 1823
rect 1291 1789 1307 1823
rect 1341 1789 1357 1823
rect 1531 1789 1547 1823
rect 1581 1789 1597 1823
rect 1771 1789 1787 1823
rect 1821 1789 1837 1823
rect 2011 1789 2027 1823
rect 2061 1789 2077 1823
rect 2251 1789 2267 1823
rect 2301 1789 2317 1823
rect 48 1730 82 1746
rect 48 1538 82 1554
rect 166 1730 200 1746
rect 166 1538 200 1554
rect 288 1730 322 1746
rect 288 1538 322 1554
rect 406 1730 440 1746
rect 406 1538 440 1554
rect 528 1730 562 1746
rect 528 1538 562 1554
rect 646 1730 680 1746
rect 646 1538 680 1554
rect 768 1730 802 1746
rect 768 1538 802 1554
rect 886 1730 920 1746
rect 886 1538 920 1554
rect 1008 1730 1042 1746
rect 1008 1538 1042 1554
rect 1126 1730 1160 1746
rect 1126 1538 1160 1554
rect 1248 1730 1282 1746
rect 1248 1538 1282 1554
rect 1366 1730 1400 1746
rect 1366 1538 1400 1554
rect 1488 1730 1522 1746
rect 1488 1538 1522 1554
rect 1606 1730 1640 1746
rect 1606 1538 1640 1554
rect 1728 1730 1762 1746
rect 1728 1538 1762 1554
rect 1846 1730 1880 1746
rect 1846 1538 1880 1554
rect 1968 1730 2002 1746
rect 1968 1538 2002 1554
rect 2086 1730 2120 1746
rect 2086 1538 2120 1554
rect 2208 1730 2242 1746
rect 2208 1538 2242 1554
rect 2326 1730 2360 1746
rect 2326 1538 2360 1554
rect 91 1419 107 1453
rect 141 1419 157 1453
rect 331 1419 347 1453
rect 381 1419 397 1453
rect 571 1419 587 1453
rect 621 1419 637 1453
rect 811 1419 827 1453
rect 861 1419 877 1453
rect 1051 1419 1067 1453
rect 1101 1419 1117 1453
rect 1291 1419 1307 1453
rect 1341 1419 1357 1453
rect 1531 1419 1547 1453
rect 1581 1419 1597 1453
rect 1771 1419 1787 1453
rect 1821 1419 1837 1453
rect 2011 1419 2027 1453
rect 2061 1419 2077 1453
rect 2251 1419 2267 1453
rect 2301 1419 2317 1453
rect 48 1360 82 1376
rect 48 1168 82 1184
rect 166 1360 200 1376
rect 166 1168 200 1184
rect 288 1360 322 1376
rect 288 1168 322 1184
rect 406 1360 440 1376
rect 406 1168 440 1184
rect 528 1360 562 1376
rect 528 1168 562 1184
rect 646 1360 680 1376
rect 646 1168 680 1184
rect 768 1360 802 1376
rect 768 1168 802 1184
rect 886 1360 920 1376
rect 886 1168 920 1184
rect 1008 1360 1042 1376
rect 1008 1168 1042 1184
rect 1126 1360 1160 1376
rect 1126 1168 1160 1184
rect 1248 1360 1282 1376
rect 1248 1168 1282 1184
rect 1366 1360 1400 1376
rect 1366 1168 1400 1184
rect 1488 1360 1522 1376
rect 1488 1168 1522 1184
rect 1606 1360 1640 1376
rect 1606 1168 1640 1184
rect 1728 1360 1762 1376
rect 1728 1168 1762 1184
rect 1846 1360 1880 1376
rect 1846 1168 1880 1184
rect 1968 1360 2002 1376
rect 1968 1168 2002 1184
rect 2086 1360 2120 1376
rect 2086 1168 2120 1184
rect 2208 1360 2242 1376
rect 2208 1168 2242 1184
rect 2326 1360 2360 1376
rect 2326 1168 2360 1184
rect 91 1049 107 1083
rect 141 1049 157 1083
rect 331 1049 347 1083
rect 381 1049 397 1083
rect 571 1049 587 1083
rect 621 1049 637 1083
rect 811 1049 827 1083
rect 861 1049 877 1083
rect 1051 1049 1067 1083
rect 1101 1049 1117 1083
rect 1291 1049 1307 1083
rect 1341 1049 1357 1083
rect 1531 1049 1547 1083
rect 1581 1049 1597 1083
rect 1771 1049 1787 1083
rect 1821 1049 1837 1083
rect 2011 1049 2027 1083
rect 2061 1049 2077 1083
rect 2251 1049 2267 1083
rect 2301 1049 2317 1083
rect 48 990 82 1006
rect 48 798 82 814
rect 166 990 200 1006
rect 166 798 200 814
rect 288 990 322 1006
rect 288 798 322 814
rect 406 990 440 1006
rect 406 798 440 814
rect 528 990 562 1006
rect 528 798 562 814
rect 646 990 680 1006
rect 646 798 680 814
rect 768 990 802 1006
rect 768 798 802 814
rect 886 990 920 1006
rect 886 798 920 814
rect 1008 990 1042 1006
rect 1008 798 1042 814
rect 1126 990 1160 1006
rect 1126 798 1160 814
rect 1248 990 1282 1006
rect 1248 798 1282 814
rect 1366 990 1400 1006
rect 1366 798 1400 814
rect 1488 990 1522 1006
rect 1488 798 1522 814
rect 1606 990 1640 1006
rect 1606 798 1640 814
rect 1728 990 1762 1006
rect 1728 798 1762 814
rect 1846 990 1880 1006
rect 1846 798 1880 814
rect 1968 990 2002 1006
rect 1968 798 2002 814
rect 2086 990 2120 1006
rect 2086 798 2120 814
rect 2208 990 2242 1006
rect 2208 798 2242 814
rect 2326 990 2360 1006
rect 2326 798 2360 814
rect 48 666 82 682
rect 48 474 82 490
rect 166 666 200 682
rect 166 474 200 490
rect 288 666 322 682
rect 288 474 322 490
rect 406 666 440 682
rect 406 474 440 490
rect 528 666 562 682
rect 528 474 562 490
rect 646 666 680 682
rect 646 474 680 490
rect 768 666 802 682
rect 768 474 802 490
rect 886 666 920 682
rect 886 474 920 490
rect 1008 666 1042 682
rect 1008 474 1042 490
rect 1126 666 1160 682
rect 1126 474 1160 490
rect 1248 666 1282 682
rect 1248 474 1282 490
rect 1366 666 1400 682
rect 1366 474 1400 490
rect 1488 666 1522 682
rect 1488 474 1522 490
rect 1606 666 1640 682
rect 1606 474 1640 490
rect 1728 666 1762 682
rect 1728 474 1762 490
rect 1846 666 1880 682
rect 1846 474 1880 490
rect 1968 666 2002 682
rect 1968 474 2002 490
rect 2086 666 2120 682
rect 2086 474 2120 490
rect 2208 666 2242 682
rect 2208 474 2242 490
rect 2326 666 2360 682
rect 2326 474 2360 490
rect 91 397 107 431
rect 141 397 157 431
rect 331 397 347 431
rect 381 397 397 431
rect 571 397 587 431
rect 621 397 637 431
rect 811 397 827 431
rect 861 397 877 431
rect 1051 397 1067 431
rect 1101 397 1117 431
rect 1291 397 1307 431
rect 1341 397 1357 431
rect 1531 397 1547 431
rect 1581 397 1597 431
rect 1771 397 1787 431
rect 1821 397 1837 431
rect 2011 397 2027 431
rect 2061 397 2077 431
rect 2251 397 2267 431
rect 2301 397 2317 431
rect 48 296 82 312
rect 48 104 82 120
rect 166 296 200 312
rect 166 104 200 120
rect 288 296 322 312
rect 288 104 322 120
rect 406 296 440 312
rect 406 104 440 120
rect 528 296 562 312
rect 528 104 562 120
rect 646 296 680 312
rect 646 104 680 120
rect 768 296 802 312
rect 768 104 802 120
rect 886 296 920 312
rect 886 104 920 120
rect 1008 296 1042 312
rect 1008 104 1042 120
rect 1126 296 1160 312
rect 1126 104 1160 120
rect 1248 296 1282 312
rect 1248 104 1282 120
rect 1366 296 1400 312
rect 1366 104 1400 120
rect 1488 296 1522 312
rect 1488 104 1522 120
rect 1606 296 1640 312
rect 1606 104 1640 120
rect 1728 296 1762 312
rect 1728 104 1762 120
rect 1846 296 1880 312
rect 1846 104 1880 120
rect 1968 296 2002 312
rect 1968 104 2002 120
rect 2086 296 2120 312
rect 2086 104 2120 120
rect 2208 296 2242 312
rect 2208 104 2242 120
rect 2326 296 2360 312
rect 2326 104 2360 120
rect 91 27 107 61
rect 141 27 157 61
rect 331 27 347 61
rect 381 27 397 61
rect 571 27 587 61
rect 621 27 637 61
rect 811 27 827 61
rect 861 27 877 61
rect 1051 27 1067 61
rect 1101 27 1117 61
rect 1291 27 1307 61
rect 1341 27 1357 61
rect 1531 27 1547 61
rect 1581 27 1597 61
rect 1771 27 1787 61
rect 1821 27 1837 61
rect 2011 27 2027 61
rect 2061 27 2077 61
rect 2251 27 2267 61
rect 2301 27 2317 61
rect 48 -74 82 -58
rect 48 -266 82 -250
rect 166 -74 200 -58
rect 166 -266 200 -250
rect 288 -74 322 -58
rect 288 -266 322 -250
rect 406 -74 440 -58
rect 406 -266 440 -250
rect 528 -74 562 -58
rect 528 -266 562 -250
rect 646 -74 680 -58
rect 646 -266 680 -250
rect 768 -74 802 -58
rect 768 -266 802 -250
rect 886 -74 920 -58
rect 886 -266 920 -250
rect 1008 -74 1042 -58
rect 1008 -266 1042 -250
rect 1126 -74 1160 -58
rect 1126 -266 1160 -250
rect 1248 -74 1282 -58
rect 1248 -266 1282 -250
rect 1366 -74 1400 -58
rect 1366 -266 1400 -250
rect 1488 -74 1522 -58
rect 1488 -266 1522 -250
rect 1606 -74 1640 -58
rect 1606 -266 1640 -250
rect 1728 -74 1762 -58
rect 1728 -266 1762 -250
rect 1846 -74 1880 -58
rect 1846 -266 1880 -250
rect 1968 -74 2002 -58
rect 1968 -266 2002 -250
rect 2086 -74 2120 -58
rect 2086 -266 2120 -250
rect 2208 -74 2242 -58
rect 2208 -266 2242 -250
rect 2326 -74 2360 -58
rect 2326 -266 2360 -250
rect 91 -343 107 -309
rect 141 -343 157 -309
rect 331 -343 347 -309
rect 381 -343 397 -309
rect 571 -343 587 -309
rect 621 -343 637 -309
rect 811 -343 827 -309
rect 861 -343 877 -309
rect 1051 -343 1067 -309
rect 1101 -343 1117 -309
rect 1291 -343 1307 -309
rect 1341 -343 1357 -309
rect 1531 -343 1547 -309
rect 1581 -343 1597 -309
rect 1771 -343 1787 -309
rect 1821 -343 1837 -309
rect 2011 -343 2027 -309
rect 2061 -343 2077 -309
rect 2251 -343 2267 -309
rect 2301 -343 2317 -309
rect 48 -444 82 -428
rect 48 -636 82 -620
rect 166 -444 200 -428
rect 166 -636 200 -620
rect 288 -444 322 -428
rect 288 -636 322 -620
rect 406 -444 440 -428
rect 406 -636 440 -620
rect 528 -444 562 -428
rect 528 -636 562 -620
rect 646 -444 680 -428
rect 646 -636 680 -620
rect 768 -444 802 -428
rect 768 -636 802 -620
rect 886 -444 920 -428
rect 886 -636 920 -620
rect 1008 -444 1042 -428
rect 1008 -636 1042 -620
rect 1126 -444 1160 -428
rect 1126 -636 1160 -620
rect 1248 -444 1282 -428
rect 1248 -636 1282 -620
rect 1366 -444 1400 -428
rect 1366 -636 1400 -620
rect 1488 -444 1522 -428
rect 1488 -636 1522 -620
rect 1606 -444 1640 -428
rect 1606 -636 1640 -620
rect 1728 -444 1762 -428
rect 1728 -636 1762 -620
rect 1846 -444 1880 -428
rect 1846 -636 1880 -620
rect 1968 -444 2002 -428
rect 1968 -636 2002 -620
rect 2086 -444 2120 -428
rect 2086 -636 2120 -620
rect 2208 -444 2242 -428
rect 2208 -636 2242 -620
rect 2326 -444 2360 -428
rect 2326 -636 2360 -620
rect 91 -713 107 -679
rect 141 -713 157 -679
rect 331 -713 347 -679
rect 381 -713 397 -679
rect 571 -713 587 -679
rect 621 -713 637 -679
rect 811 -713 827 -679
rect 861 -713 877 -679
rect 1051 -713 1067 -679
rect 1101 -713 1117 -679
rect 1291 -713 1307 -679
rect 1341 -713 1357 -679
rect 1531 -713 1547 -679
rect 1581 -713 1597 -679
rect 1771 -713 1787 -679
rect 1821 -713 1837 -679
rect 2011 -713 2027 -679
rect 2061 -713 2077 -679
rect 2251 -713 2267 -679
rect 2301 -713 2317 -679
rect 2440 -780 2460 2240
rect -40 -800 2460 -780
rect 2500 -840 2520 2300
rect -100 -860 2520 -840
<< viali >>
rect 107 2159 141 2193
rect 347 2159 381 2193
rect 587 2159 621 2193
rect 827 2159 861 2193
rect 1067 2159 1101 2193
rect 1307 2159 1341 2193
rect 1547 2159 1581 2193
rect 1787 2159 1821 2193
rect 2027 2159 2061 2193
rect 2267 2159 2301 2193
rect 48 1924 82 2100
rect 166 1924 200 2100
rect 288 1924 322 2100
rect 406 1924 440 2100
rect 528 1924 562 2100
rect 646 1924 680 2100
rect 768 1924 802 2100
rect 886 1924 920 2100
rect 1008 1924 1042 2100
rect 1126 1924 1160 2100
rect 1248 1924 1282 2100
rect 1366 1924 1400 2100
rect 1488 1924 1522 2100
rect 1606 1924 1640 2100
rect 1728 1924 1762 2100
rect 1846 1924 1880 2100
rect 1968 1924 2002 2100
rect 2086 1924 2120 2100
rect 2208 1924 2242 2100
rect 2326 1924 2360 2100
rect 107 1789 141 1823
rect 347 1789 381 1823
rect 587 1789 621 1823
rect 827 1789 861 1823
rect 1067 1789 1101 1823
rect 1307 1789 1341 1823
rect 1547 1789 1581 1823
rect 1787 1789 1821 1823
rect 2027 1789 2061 1823
rect 2267 1789 2301 1823
rect 48 1554 82 1730
rect 166 1554 200 1730
rect 288 1554 322 1730
rect 406 1554 440 1730
rect 528 1554 562 1730
rect 646 1554 680 1730
rect 768 1554 802 1730
rect 886 1554 920 1730
rect 1008 1554 1042 1730
rect 1126 1554 1160 1730
rect 1248 1554 1282 1730
rect 1366 1554 1400 1730
rect 1488 1554 1522 1730
rect 1606 1554 1640 1730
rect 1728 1554 1762 1730
rect 1846 1554 1880 1730
rect 1968 1554 2002 1730
rect 2086 1554 2120 1730
rect 2208 1554 2242 1730
rect 2326 1554 2360 1730
rect 107 1419 141 1453
rect 347 1419 381 1453
rect 587 1419 621 1453
rect 827 1419 861 1453
rect 1067 1419 1101 1453
rect 1307 1419 1341 1453
rect 1547 1419 1581 1453
rect 1787 1419 1821 1453
rect 2027 1419 2061 1453
rect 2267 1419 2301 1453
rect 48 1184 82 1360
rect 166 1184 200 1360
rect 288 1184 322 1360
rect 406 1184 440 1360
rect 528 1184 562 1360
rect 646 1184 680 1360
rect 768 1184 802 1360
rect 886 1184 920 1360
rect 1008 1184 1042 1360
rect 1126 1184 1160 1360
rect 1248 1184 1282 1360
rect 1366 1184 1400 1360
rect 1488 1184 1522 1360
rect 1606 1184 1640 1360
rect 1728 1184 1762 1360
rect 1846 1184 1880 1360
rect 1968 1184 2002 1360
rect 2086 1184 2120 1360
rect 2208 1184 2242 1360
rect 2326 1184 2360 1360
rect 107 1049 141 1083
rect 347 1049 381 1083
rect 587 1049 621 1083
rect 827 1049 861 1083
rect 1067 1049 1101 1083
rect 1307 1049 1341 1083
rect 1547 1049 1581 1083
rect 1787 1049 1821 1083
rect 2027 1049 2061 1083
rect 2267 1049 2301 1083
rect 48 814 82 990
rect 166 814 200 990
rect 288 814 322 990
rect 406 814 440 990
rect 528 814 562 990
rect 646 814 680 990
rect 768 814 802 990
rect 886 814 920 990
rect 1008 814 1042 990
rect 1126 814 1160 990
rect 1248 814 1282 990
rect 1366 814 1400 990
rect 1488 814 1522 990
rect 1606 814 1640 990
rect 1728 814 1762 990
rect 1846 814 1880 990
rect 1968 814 2002 990
rect 2086 814 2120 990
rect 2208 814 2242 990
rect 2326 814 2360 990
rect 48 490 82 666
rect 166 490 200 666
rect 288 490 322 666
rect 406 490 440 666
rect 528 490 562 666
rect 646 490 680 666
rect 768 490 802 666
rect 886 490 920 666
rect 1008 490 1042 666
rect 1126 490 1160 666
rect 1248 490 1282 666
rect 1366 490 1400 666
rect 1488 490 1522 666
rect 1606 490 1640 666
rect 1728 490 1762 666
rect 1846 490 1880 666
rect 1968 490 2002 666
rect 2086 490 2120 666
rect 2208 490 2242 666
rect 2326 490 2360 666
rect 107 397 141 431
rect 347 397 381 431
rect 587 397 621 431
rect 827 397 861 431
rect 1067 397 1101 431
rect 1307 397 1341 431
rect 1547 397 1581 431
rect 1787 397 1821 431
rect 2027 397 2061 431
rect 2267 397 2301 431
rect 48 120 82 296
rect 166 120 200 296
rect 288 120 322 296
rect 406 120 440 296
rect 528 120 562 296
rect 646 120 680 296
rect 768 120 802 296
rect 886 120 920 296
rect 1008 120 1042 296
rect 1126 120 1160 296
rect 1248 120 1282 296
rect 1366 120 1400 296
rect 1488 120 1522 296
rect 1606 120 1640 296
rect 1728 120 1762 296
rect 1846 120 1880 296
rect 1968 120 2002 296
rect 2086 120 2120 296
rect 2208 120 2242 296
rect 2326 120 2360 296
rect 107 27 141 61
rect 347 27 381 61
rect 587 27 621 61
rect 827 27 861 61
rect 1067 27 1101 61
rect 1307 27 1341 61
rect 1547 27 1581 61
rect 1787 27 1821 61
rect 2027 27 2061 61
rect 2267 27 2301 61
rect 48 -250 82 -74
rect 166 -250 200 -74
rect 288 -250 322 -74
rect 406 -250 440 -74
rect 528 -250 562 -74
rect 646 -250 680 -74
rect 768 -250 802 -74
rect 886 -250 920 -74
rect 1008 -250 1042 -74
rect 1126 -250 1160 -74
rect 1248 -250 1282 -74
rect 1366 -250 1400 -74
rect 1488 -250 1522 -74
rect 1606 -250 1640 -74
rect 1728 -250 1762 -74
rect 1846 -250 1880 -74
rect 1968 -250 2002 -74
rect 2086 -250 2120 -74
rect 2208 -250 2242 -74
rect 2326 -250 2360 -74
rect 107 -343 141 -309
rect 347 -343 381 -309
rect 587 -343 621 -309
rect 827 -343 861 -309
rect 1067 -343 1101 -309
rect 1307 -343 1341 -309
rect 1547 -343 1581 -309
rect 1787 -343 1821 -309
rect 2027 -343 2061 -309
rect 2267 -343 2301 -309
rect 48 -620 82 -444
rect 166 -620 200 -444
rect 288 -620 322 -444
rect 406 -620 440 -444
rect 528 -620 562 -444
rect 646 -620 680 -444
rect 768 -620 802 -444
rect 886 -620 920 -444
rect 1008 -620 1042 -444
rect 1126 -620 1160 -444
rect 1248 -620 1282 -444
rect 1366 -620 1400 -444
rect 1488 -620 1522 -444
rect 1606 -620 1640 -444
rect 1728 -620 1762 -444
rect 1846 -620 1880 -444
rect 1968 -620 2002 -444
rect 2086 -620 2120 -444
rect 2208 -620 2242 -444
rect 2326 -620 2360 -444
rect 107 -713 141 -679
rect 347 -713 381 -679
rect 587 -713 621 -679
rect 827 -713 861 -679
rect 1067 -713 1101 -679
rect 1307 -713 1341 -679
rect 1547 -713 1581 -679
rect 1787 -713 1821 -679
rect 2027 -713 2061 -679
rect 2267 -713 2301 -679
rect 0 -840 2420 -800
<< metal1 >>
rect 30 2193 220 2220
rect 30 2159 107 2193
rect 141 2159 220 2193
rect 30 2120 220 2159
rect 320 2150 330 2220
rect 400 2150 410 2220
rect 560 2150 570 2220
rect 640 2150 650 2220
rect 800 2150 810 2220
rect 880 2150 890 2220
rect 1040 2150 1050 2220
rect 1120 2150 1130 2220
rect 1280 2150 1290 2220
rect 1360 2150 1370 2220
rect 1520 2150 1530 2220
rect 1600 2150 1610 2220
rect 1760 2150 1770 2220
rect 1840 2150 1850 2220
rect 2000 2150 2010 2220
rect 2080 2150 2090 2220
rect 2190 2193 2380 2220
rect 2190 2159 2267 2193
rect 2301 2159 2380 2193
rect 2190 2120 2380 2159
rect 30 2110 90 2120
rect 30 1920 38 2110
rect 30 1910 90 1920
rect 160 2110 220 2120
rect 212 1920 220 2110
rect 160 1910 220 1920
rect 270 2110 330 2120
rect 270 1920 278 2110
rect 270 1910 330 1920
rect 400 2110 460 2120
rect 452 1920 460 2110
rect 400 1910 460 1920
rect 510 2110 570 2120
rect 510 1920 518 2110
rect 510 1910 570 1920
rect 640 2110 700 2120
rect 692 1920 700 2110
rect 640 1910 700 1920
rect 750 2110 810 2120
rect 750 1920 758 2110
rect 750 1910 810 1920
rect 880 2110 940 2120
rect 932 1920 940 2110
rect 880 1910 940 1920
rect 990 2110 1050 2120
rect 990 1920 998 2110
rect 990 1910 1050 1920
rect 1120 2110 1180 2120
rect 1172 1920 1180 2110
rect 1120 1910 1180 1920
rect 1230 2110 1290 2120
rect 1230 1920 1238 2110
rect 1230 1910 1290 1920
rect 1360 2110 1420 2120
rect 1412 1920 1420 2110
rect 1360 1910 1420 1920
rect 1470 2110 1530 2120
rect 1470 1920 1478 2110
rect 1470 1910 1530 1920
rect 1600 2110 1660 2120
rect 1652 1920 1660 2110
rect 1600 1910 1660 1920
rect 1710 2110 1770 2120
rect 1710 1920 1718 2110
rect 1710 1910 1770 1920
rect 1840 2110 1900 2120
rect 1892 1920 1900 2110
rect 1840 1910 1900 1920
rect 1950 2110 2010 2120
rect 1950 1920 1958 2110
rect 1950 1910 2010 1920
rect 2080 2110 2140 2120
rect 2132 1920 2140 2110
rect 2080 1910 2140 1920
rect 2190 2110 2250 2120
rect 2190 1920 2198 2110
rect 2190 1910 2250 1920
rect 2320 2110 2380 2120
rect 2372 1920 2380 2110
rect 2320 1910 2380 1920
rect 30 1823 220 1850
rect 30 1789 107 1823
rect 141 1789 220 1823
rect 30 1750 220 1789
rect 320 1780 330 1850
rect 400 1780 410 1850
rect 560 1780 570 1850
rect 640 1780 650 1850
rect 800 1780 810 1850
rect 880 1780 890 1850
rect 1040 1780 1050 1850
rect 1120 1780 1130 1850
rect 1280 1780 1290 1850
rect 1360 1780 1370 1850
rect 1520 1780 1530 1850
rect 1600 1780 1610 1850
rect 1760 1780 1770 1850
rect 1840 1780 1850 1850
rect 2000 1780 2010 1850
rect 2080 1780 2090 1850
rect 2190 1823 2380 1850
rect 2190 1789 2267 1823
rect 2301 1789 2380 1823
rect 2190 1750 2380 1789
rect 30 1740 90 1750
rect 30 1550 38 1740
rect 30 1540 90 1550
rect 160 1740 220 1750
rect 212 1550 220 1740
rect 160 1540 220 1550
rect 270 1740 330 1750
rect 270 1550 278 1740
rect 270 1540 330 1550
rect 400 1740 460 1750
rect 452 1550 460 1740
rect 400 1540 460 1550
rect 510 1740 570 1750
rect 510 1550 518 1740
rect 510 1540 570 1550
rect 640 1740 700 1750
rect 692 1550 700 1740
rect 640 1540 700 1550
rect 750 1740 810 1750
rect 750 1550 758 1740
rect 750 1540 810 1550
rect 880 1740 940 1750
rect 932 1550 940 1740
rect 880 1540 940 1550
rect 990 1740 1050 1750
rect 990 1550 998 1740
rect 990 1540 1050 1550
rect 1120 1740 1180 1750
rect 1172 1550 1180 1740
rect 1120 1540 1180 1550
rect 1230 1740 1290 1750
rect 1230 1550 1238 1740
rect 1230 1540 1290 1550
rect 1360 1740 1420 1750
rect 1412 1550 1420 1740
rect 1360 1540 1420 1550
rect 1470 1740 1530 1750
rect 1470 1550 1478 1740
rect 1470 1540 1530 1550
rect 1600 1740 1660 1750
rect 1652 1550 1660 1740
rect 1600 1540 1660 1550
rect 1710 1740 1770 1750
rect 1710 1550 1718 1740
rect 1710 1540 1770 1550
rect 1840 1740 1900 1750
rect 1892 1550 1900 1740
rect 1840 1540 1900 1550
rect 1950 1740 2010 1750
rect 1950 1550 1958 1740
rect 1950 1540 2010 1550
rect 2080 1740 2140 1750
rect 2132 1550 2140 1740
rect 2080 1540 2140 1550
rect 2190 1740 2250 1750
rect 2190 1550 2198 1740
rect 2190 1540 2250 1550
rect 2320 1740 2380 1750
rect 2372 1550 2380 1740
rect 2320 1540 2380 1550
rect 30 1453 220 1480
rect 30 1419 107 1453
rect 141 1419 220 1453
rect 30 1380 220 1419
rect 320 1410 330 1480
rect 400 1410 410 1480
rect 560 1410 570 1480
rect 640 1410 650 1480
rect 800 1410 810 1480
rect 880 1410 890 1480
rect 1040 1410 1050 1480
rect 1120 1410 1130 1480
rect 1280 1410 1290 1480
rect 1360 1410 1370 1480
rect 1520 1410 1530 1480
rect 1600 1410 1610 1480
rect 1760 1410 1770 1480
rect 1840 1410 1850 1480
rect 2000 1410 2010 1480
rect 2080 1410 2090 1480
rect 2190 1453 2380 1480
rect 2190 1419 2267 1453
rect 2301 1419 2380 1453
rect 2190 1380 2380 1419
rect 30 1370 90 1380
rect 30 1180 38 1370
rect 30 1170 90 1180
rect 160 1370 220 1380
rect 212 1180 220 1370
rect 160 1170 220 1180
rect 270 1370 330 1380
rect 270 1180 278 1370
rect 270 1170 330 1180
rect 400 1370 460 1380
rect 452 1180 460 1370
rect 400 1170 460 1180
rect 510 1370 570 1380
rect 510 1180 518 1370
rect 510 1170 570 1180
rect 640 1370 700 1380
rect 692 1180 700 1370
rect 640 1170 700 1180
rect 750 1370 810 1380
rect 750 1180 758 1370
rect 750 1170 810 1180
rect 880 1370 940 1380
rect 932 1180 940 1370
rect 880 1170 940 1180
rect 990 1370 1050 1380
rect 990 1180 998 1370
rect 990 1170 1050 1180
rect 1120 1370 1180 1380
rect 1172 1180 1180 1370
rect 1120 1170 1180 1180
rect 1230 1370 1290 1380
rect 1230 1180 1238 1370
rect 1230 1170 1290 1180
rect 1360 1370 1420 1380
rect 1412 1180 1420 1370
rect 1360 1170 1420 1180
rect 1470 1370 1530 1380
rect 1470 1180 1478 1370
rect 1470 1170 1530 1180
rect 1600 1370 1660 1380
rect 1652 1180 1660 1370
rect 1600 1170 1660 1180
rect 1710 1370 1770 1380
rect 1710 1180 1718 1370
rect 1710 1170 1770 1180
rect 1840 1370 1900 1380
rect 1892 1180 1900 1370
rect 1840 1170 1900 1180
rect 1950 1370 2010 1380
rect 1950 1180 1958 1370
rect 1950 1170 2010 1180
rect 2080 1370 2140 1380
rect 2132 1180 2140 1370
rect 2080 1170 2140 1180
rect 2190 1370 2250 1380
rect 2190 1180 2198 1370
rect 2190 1170 2250 1180
rect 2320 1370 2380 1380
rect 2372 1180 2380 1370
rect 2320 1170 2380 1180
rect 30 1083 220 1110
rect 30 1049 107 1083
rect 141 1049 220 1083
rect 30 1010 220 1049
rect 320 1040 330 1110
rect 400 1040 410 1110
rect 560 1040 570 1110
rect 640 1040 650 1110
rect 800 1040 810 1110
rect 880 1040 890 1110
rect 1040 1040 1050 1110
rect 1120 1040 1130 1110
rect 1280 1040 1290 1110
rect 1360 1040 1370 1110
rect 1520 1040 1530 1110
rect 1600 1040 1610 1110
rect 1760 1040 1770 1110
rect 1840 1040 1850 1110
rect 2000 1040 2010 1110
rect 2080 1040 2090 1110
rect 2190 1083 2380 1110
rect 2190 1049 2267 1083
rect 2301 1049 2380 1083
rect 2190 1010 2380 1049
rect 30 1000 90 1010
rect 30 810 38 1000
rect 30 800 90 810
rect 160 1000 220 1010
rect 212 810 220 1000
rect 160 800 220 810
rect 270 1000 330 1010
rect 270 810 278 1000
rect 270 800 330 810
rect 400 1000 460 1010
rect 452 810 460 1000
rect 400 800 460 810
rect 510 1000 570 1010
rect 510 810 518 1000
rect 510 800 570 810
rect 640 1000 700 1010
rect 692 810 700 1000
rect 640 800 700 810
rect 750 1000 810 1010
rect 750 810 758 1000
rect 750 800 810 810
rect 880 1000 940 1010
rect 932 810 940 1000
rect 880 800 940 810
rect 990 1000 1050 1010
rect 990 810 998 1000
rect 990 800 1050 810
rect 1120 1000 1180 1010
rect 1172 810 1180 1000
rect 1120 800 1180 810
rect 1230 1000 1290 1010
rect 1230 810 1238 1000
rect 1230 800 1290 810
rect 1360 1000 1420 1010
rect 1412 810 1420 1000
rect 1360 800 1420 810
rect 1470 1000 1530 1010
rect 1470 810 1478 1000
rect 1470 800 1530 810
rect 1600 1000 1660 1010
rect 1652 810 1660 1000
rect 1600 800 1660 810
rect 1710 1000 1770 1010
rect 1710 810 1718 1000
rect 1710 800 1770 810
rect 1840 1000 1900 1010
rect 1892 810 1900 1000
rect 1840 800 1900 810
rect 1950 1000 2010 1010
rect 1950 810 1958 1000
rect 1950 800 2010 810
rect 2080 1000 2140 1010
rect 2132 810 2140 1000
rect 2080 800 2140 810
rect 2190 1000 2250 1010
rect 2190 810 2198 1000
rect 2190 800 2250 810
rect 2320 1000 2380 1010
rect 2372 810 2380 1000
rect 2320 800 2380 810
rect 30 670 90 680
rect 30 480 38 670
rect 30 470 90 480
rect 160 670 220 680
rect 212 480 220 670
rect 160 470 220 480
rect 270 670 330 680
rect 270 480 278 670
rect 270 470 330 480
rect 400 670 460 680
rect 452 480 460 670
rect 400 470 460 480
rect 510 670 570 680
rect 510 480 518 670
rect 510 470 570 480
rect 640 670 700 680
rect 692 480 700 670
rect 640 470 700 480
rect 750 670 810 680
rect 750 480 758 670
rect 750 470 810 480
rect 880 670 940 680
rect 932 480 940 670
rect 880 470 940 480
rect 990 670 1050 680
rect 990 480 998 670
rect 990 470 1050 480
rect 1120 670 1180 680
rect 1172 480 1180 670
rect 1120 470 1180 480
rect 1230 670 1290 680
rect 1230 480 1238 670
rect 1230 470 1290 480
rect 1360 666 1420 680
rect 1360 490 1366 666
rect 1400 490 1420 666
rect 30 431 220 470
rect 30 397 107 431
rect 141 397 220 431
rect 30 370 220 397
rect 320 370 330 440
rect 400 370 410 440
rect 560 370 570 440
rect 640 370 650 440
rect 800 370 810 440
rect 880 370 890 440
rect 1040 370 1050 440
rect 1120 370 1130 440
rect 1280 370 1290 440
rect 1360 360 1420 490
rect 1470 670 1530 680
rect 1470 480 1478 670
rect 1470 470 1530 480
rect 1600 670 1660 680
rect 1652 480 1660 670
rect 1600 470 1660 480
rect 1710 670 1770 680
rect 1710 480 1718 670
rect 1710 470 1770 480
rect 1840 670 1900 680
rect 1892 480 1900 670
rect 1840 470 1900 480
rect 1950 670 2010 680
rect 1950 480 1958 670
rect 1950 470 2010 480
rect 2080 670 2140 680
rect 2132 480 2140 670
rect 2080 470 2140 480
rect 2190 670 2250 680
rect 2190 480 2198 670
rect 2190 470 2250 480
rect 2320 670 2380 680
rect 2372 480 2380 670
rect 2320 470 2380 480
rect 1520 370 1530 440
rect 1600 370 1610 440
rect 1760 370 1770 440
rect 1840 370 1850 440
rect 2000 370 2010 440
rect 2080 370 2090 440
rect 2190 431 2380 470
rect 2190 397 2267 431
rect 2301 397 2380 431
rect 2190 370 2380 397
rect 30 300 90 310
rect 30 110 38 300
rect 30 100 90 110
rect 160 300 220 310
rect 212 110 220 300
rect 160 100 220 110
rect 270 300 330 310
rect 270 110 278 300
rect 270 100 330 110
rect 400 300 460 310
rect 452 110 460 300
rect 400 100 460 110
rect 510 300 570 310
rect 510 110 518 300
rect 510 100 570 110
rect 640 300 700 310
rect 692 110 700 300
rect 640 100 700 110
rect 750 300 810 310
rect 750 110 758 300
rect 750 100 810 110
rect 880 300 940 310
rect 932 110 940 300
rect 880 100 940 110
rect 990 300 1050 310
rect 990 110 998 300
rect 990 100 1050 110
rect 1120 300 1180 310
rect 1172 110 1180 300
rect 1120 100 1180 110
rect 1230 300 1290 310
rect 1230 110 1238 300
rect 1230 100 1290 110
rect 1360 300 1420 310
rect 1412 110 1420 300
rect 1360 100 1420 110
rect 1470 300 1530 310
rect 1470 110 1478 300
rect 1470 100 1530 110
rect 1600 300 1660 310
rect 1652 110 1660 300
rect 1600 100 1660 110
rect 1710 300 1770 310
rect 1710 110 1718 300
rect 1710 100 1770 110
rect 1840 300 1900 310
rect 1892 110 1900 300
rect 1840 100 1900 110
rect 1950 300 2010 310
rect 1950 110 1958 300
rect 1950 100 2010 110
rect 2080 300 2140 310
rect 2132 110 2140 300
rect 2080 100 2140 110
rect 2190 300 2250 310
rect 2190 110 2198 300
rect 2190 100 2250 110
rect 2320 300 2380 310
rect 2372 110 2380 300
rect 2320 100 2380 110
rect 30 61 220 100
rect 30 27 107 61
rect 141 27 220 61
rect 30 0 220 27
rect 320 0 330 70
rect 400 0 410 70
rect 560 0 570 70
rect 640 0 650 70
rect 800 0 810 70
rect 880 0 890 70
rect 1040 0 1050 70
rect 1120 0 1130 70
rect 1280 0 1290 70
rect 1360 0 1370 70
rect 1520 0 1530 70
rect 1600 0 1610 70
rect 1760 0 1770 70
rect 1840 0 1850 70
rect 2000 0 2010 70
rect 2080 0 2090 70
rect 2190 61 2380 100
rect 2190 27 2267 61
rect 2301 27 2380 61
rect 2190 0 2380 27
rect 30 -70 90 -60
rect 30 -260 38 -70
rect 30 -270 90 -260
rect 160 -70 220 -60
rect 212 -260 220 -70
rect 160 -270 220 -260
rect 270 -70 330 -60
rect 270 -260 278 -70
rect 270 -270 330 -260
rect 400 -70 460 -60
rect 452 -260 460 -70
rect 400 -270 460 -260
rect 510 -70 570 -60
rect 510 -260 518 -70
rect 510 -270 570 -260
rect 640 -70 700 -60
rect 692 -260 700 -70
rect 640 -270 700 -260
rect 750 -70 810 -60
rect 750 -260 758 -70
rect 750 -270 810 -260
rect 880 -70 940 -60
rect 932 -260 940 -70
rect 880 -270 940 -260
rect 990 -70 1050 -60
rect 990 -260 998 -70
rect 990 -270 1050 -260
rect 1120 -70 1180 -60
rect 1172 -260 1180 -70
rect 1120 -270 1180 -260
rect 1230 -70 1290 -60
rect 1230 -260 1238 -70
rect 1230 -270 1290 -260
rect 1360 -70 1420 -60
rect 1412 -260 1420 -70
rect 1360 -270 1420 -260
rect 1470 -70 1530 -60
rect 1470 -260 1478 -70
rect 1470 -270 1530 -260
rect 1600 -70 1660 -60
rect 1652 -260 1660 -70
rect 1600 -270 1660 -260
rect 1710 -70 1770 -60
rect 1710 -260 1718 -70
rect 1710 -270 1770 -260
rect 1840 -70 1900 -60
rect 1892 -260 1900 -70
rect 1840 -270 1900 -260
rect 1950 -70 2010 -60
rect 1950 -260 1958 -70
rect 1950 -270 2010 -260
rect 2080 -70 2140 -60
rect 2132 -260 2140 -70
rect 2080 -270 2140 -260
rect 2190 -70 2250 -60
rect 2190 -260 2198 -70
rect 2190 -270 2250 -260
rect 2320 -70 2380 -60
rect 2372 -260 2380 -70
rect 2320 -270 2380 -260
rect 30 -309 220 -270
rect 30 -343 107 -309
rect 141 -343 220 -309
rect 30 -370 220 -343
rect 320 -370 330 -300
rect 400 -370 410 -300
rect 560 -370 570 -300
rect 640 -370 650 -300
rect 800 -370 810 -300
rect 880 -370 890 -300
rect 1040 -370 1050 -300
rect 1120 -370 1130 -300
rect 1280 -370 1290 -300
rect 1360 -370 1370 -300
rect 1520 -370 1530 -300
rect 1600 -370 1610 -300
rect 1760 -370 1770 -300
rect 1840 -370 1850 -300
rect 2000 -370 2010 -300
rect 2080 -370 2090 -300
rect 2190 -309 2380 -270
rect 2190 -343 2267 -309
rect 2301 -343 2380 -309
rect 2190 -370 2380 -343
rect 30 -440 90 -430
rect 30 -630 38 -440
rect 30 -640 90 -630
rect 160 -440 220 -430
rect 212 -630 220 -440
rect 160 -640 220 -630
rect 270 -440 330 -430
rect 270 -630 278 -440
rect 270 -640 330 -630
rect 400 -440 460 -430
rect 452 -630 460 -440
rect 400 -640 460 -630
rect 510 -440 570 -430
rect 510 -630 518 -440
rect 510 -640 570 -630
rect 640 -440 700 -430
rect 692 -630 700 -440
rect 640 -640 700 -630
rect 750 -440 810 -430
rect 750 -630 758 -440
rect 750 -640 810 -630
rect 880 -440 940 -430
rect 932 -630 940 -440
rect 880 -640 940 -630
rect 990 -440 1050 -430
rect 990 -630 998 -440
rect 990 -640 1050 -630
rect 1120 -440 1180 -430
rect 1172 -630 1180 -440
rect 1120 -640 1180 -630
rect 1230 -440 1290 -430
rect 1230 -630 1238 -440
rect 1230 -640 1290 -630
rect 1360 -440 1420 -430
rect 1412 -630 1420 -440
rect 1360 -640 1420 -630
rect 1470 -440 1530 -430
rect 1470 -630 1478 -440
rect 1470 -640 1530 -630
rect 1600 -440 1660 -430
rect 1652 -630 1660 -440
rect 1600 -640 1660 -630
rect 1710 -440 1770 -430
rect 1710 -630 1718 -440
rect 1710 -640 1770 -630
rect 1840 -440 1900 -430
rect 1892 -630 1900 -440
rect 1840 -640 1900 -630
rect 1950 -440 2010 -430
rect 1950 -630 1958 -440
rect 1950 -640 2010 -630
rect 2080 -440 2140 -430
rect 2132 -630 2140 -440
rect 2080 -640 2140 -630
rect 2190 -440 2250 -430
rect 2190 -630 2198 -440
rect 2190 -640 2250 -630
rect 2320 -440 2380 -430
rect 2372 -630 2380 -440
rect 2320 -640 2380 -630
rect 30 -679 220 -640
rect 30 -713 107 -679
rect 141 -713 220 -679
rect 30 -740 220 -713
rect 320 -740 330 -670
rect 400 -740 410 -670
rect 560 -740 570 -670
rect 640 -740 650 -670
rect 800 -740 810 -670
rect 880 -740 890 -670
rect 1040 -740 1050 -670
rect 1120 -740 1130 -670
rect 1280 -740 1290 -670
rect 1360 -740 1370 -670
rect 1520 -740 1530 -670
rect 1600 -740 1610 -670
rect 1760 -740 1770 -670
rect 1840 -740 1850 -670
rect 2000 -740 2010 -670
rect 2080 -740 2090 -670
rect 2190 -679 2380 -640
rect 2190 -713 2267 -679
rect 2301 -713 2380 -679
rect 2190 -740 2380 -713
rect -20 -800 2440 -780
rect -20 -860 0 -800
rect 2420 -860 2440 -800
rect -20 -880 2440 -860
<< via1 >>
rect 330 2193 400 2220
rect 330 2159 347 2193
rect 347 2159 381 2193
rect 381 2159 400 2193
rect 330 2150 400 2159
rect 570 2193 640 2220
rect 570 2159 587 2193
rect 587 2159 621 2193
rect 621 2159 640 2193
rect 570 2150 640 2159
rect 810 2193 880 2220
rect 810 2159 827 2193
rect 827 2159 861 2193
rect 861 2159 880 2193
rect 810 2150 880 2159
rect 1050 2193 1120 2220
rect 1050 2159 1067 2193
rect 1067 2159 1101 2193
rect 1101 2159 1120 2193
rect 1050 2150 1120 2159
rect 1290 2193 1360 2220
rect 1290 2159 1307 2193
rect 1307 2159 1341 2193
rect 1341 2159 1360 2193
rect 1290 2150 1360 2159
rect 1530 2193 1600 2220
rect 1530 2159 1547 2193
rect 1547 2159 1581 2193
rect 1581 2159 1600 2193
rect 1530 2150 1600 2159
rect 1770 2193 1840 2220
rect 1770 2159 1787 2193
rect 1787 2159 1821 2193
rect 1821 2159 1840 2193
rect 1770 2150 1840 2159
rect 2010 2193 2080 2220
rect 2010 2159 2027 2193
rect 2027 2159 2061 2193
rect 2061 2159 2080 2193
rect 2010 2150 2080 2159
rect 38 2100 90 2110
rect 38 1924 48 2100
rect 48 1924 82 2100
rect 82 1924 90 2100
rect 38 1920 90 1924
rect 160 2100 212 2110
rect 160 1924 166 2100
rect 166 1924 200 2100
rect 200 1924 212 2100
rect 160 1920 212 1924
rect 278 2100 330 2110
rect 278 1924 288 2100
rect 288 1924 322 2100
rect 322 1924 330 2100
rect 278 1920 330 1924
rect 400 2100 452 2110
rect 400 1924 406 2100
rect 406 1924 440 2100
rect 440 1924 452 2100
rect 400 1920 452 1924
rect 518 2100 570 2110
rect 518 1924 528 2100
rect 528 1924 562 2100
rect 562 1924 570 2100
rect 518 1920 570 1924
rect 640 2100 692 2110
rect 640 1924 646 2100
rect 646 1924 680 2100
rect 680 1924 692 2100
rect 640 1920 692 1924
rect 758 2100 810 2110
rect 758 1924 768 2100
rect 768 1924 802 2100
rect 802 1924 810 2100
rect 758 1920 810 1924
rect 880 2100 932 2110
rect 880 1924 886 2100
rect 886 1924 920 2100
rect 920 1924 932 2100
rect 880 1920 932 1924
rect 998 2100 1050 2110
rect 998 1924 1008 2100
rect 1008 1924 1042 2100
rect 1042 1924 1050 2100
rect 998 1920 1050 1924
rect 1120 2100 1172 2110
rect 1120 1924 1126 2100
rect 1126 1924 1160 2100
rect 1160 1924 1172 2100
rect 1120 1920 1172 1924
rect 1238 2100 1290 2110
rect 1238 1924 1248 2100
rect 1248 1924 1282 2100
rect 1282 1924 1290 2100
rect 1238 1920 1290 1924
rect 1360 2100 1412 2110
rect 1360 1924 1366 2100
rect 1366 1924 1400 2100
rect 1400 1924 1412 2100
rect 1360 1920 1412 1924
rect 1478 2100 1530 2110
rect 1478 1924 1488 2100
rect 1488 1924 1522 2100
rect 1522 1924 1530 2100
rect 1478 1920 1530 1924
rect 1600 2100 1652 2110
rect 1600 1924 1606 2100
rect 1606 1924 1640 2100
rect 1640 1924 1652 2100
rect 1600 1920 1652 1924
rect 1718 2100 1770 2110
rect 1718 1924 1728 2100
rect 1728 1924 1762 2100
rect 1762 1924 1770 2100
rect 1718 1920 1770 1924
rect 1840 2100 1892 2110
rect 1840 1924 1846 2100
rect 1846 1924 1880 2100
rect 1880 1924 1892 2100
rect 1840 1920 1892 1924
rect 1958 2100 2010 2110
rect 1958 1924 1968 2100
rect 1968 1924 2002 2100
rect 2002 1924 2010 2100
rect 1958 1920 2010 1924
rect 2080 2100 2132 2110
rect 2080 1924 2086 2100
rect 2086 1924 2120 2100
rect 2120 1924 2132 2100
rect 2080 1920 2132 1924
rect 2198 2100 2250 2110
rect 2198 1924 2208 2100
rect 2208 1924 2242 2100
rect 2242 1924 2250 2100
rect 2198 1920 2250 1924
rect 2320 2100 2372 2110
rect 2320 1924 2326 2100
rect 2326 1924 2360 2100
rect 2360 1924 2372 2100
rect 2320 1920 2372 1924
rect 330 1823 400 1850
rect 330 1789 347 1823
rect 347 1789 381 1823
rect 381 1789 400 1823
rect 330 1780 400 1789
rect 570 1823 640 1850
rect 570 1789 587 1823
rect 587 1789 621 1823
rect 621 1789 640 1823
rect 570 1780 640 1789
rect 810 1823 880 1850
rect 810 1789 827 1823
rect 827 1789 861 1823
rect 861 1789 880 1823
rect 810 1780 880 1789
rect 1050 1823 1120 1850
rect 1050 1789 1067 1823
rect 1067 1789 1101 1823
rect 1101 1789 1120 1823
rect 1050 1780 1120 1789
rect 1290 1823 1360 1850
rect 1290 1789 1307 1823
rect 1307 1789 1341 1823
rect 1341 1789 1360 1823
rect 1290 1780 1360 1789
rect 1530 1823 1600 1850
rect 1530 1789 1547 1823
rect 1547 1789 1581 1823
rect 1581 1789 1600 1823
rect 1530 1780 1600 1789
rect 1770 1823 1840 1850
rect 1770 1789 1787 1823
rect 1787 1789 1821 1823
rect 1821 1789 1840 1823
rect 1770 1780 1840 1789
rect 2010 1823 2080 1850
rect 2010 1789 2027 1823
rect 2027 1789 2061 1823
rect 2061 1789 2080 1823
rect 2010 1780 2080 1789
rect 38 1730 90 1740
rect 38 1554 48 1730
rect 48 1554 82 1730
rect 82 1554 90 1730
rect 38 1550 90 1554
rect 160 1730 212 1740
rect 160 1554 166 1730
rect 166 1554 200 1730
rect 200 1554 212 1730
rect 160 1550 212 1554
rect 278 1730 330 1740
rect 278 1554 288 1730
rect 288 1554 322 1730
rect 322 1554 330 1730
rect 278 1550 330 1554
rect 400 1730 452 1740
rect 400 1554 406 1730
rect 406 1554 440 1730
rect 440 1554 452 1730
rect 400 1550 452 1554
rect 518 1730 570 1740
rect 518 1554 528 1730
rect 528 1554 562 1730
rect 562 1554 570 1730
rect 518 1550 570 1554
rect 640 1730 692 1740
rect 640 1554 646 1730
rect 646 1554 680 1730
rect 680 1554 692 1730
rect 640 1550 692 1554
rect 758 1730 810 1740
rect 758 1554 768 1730
rect 768 1554 802 1730
rect 802 1554 810 1730
rect 758 1550 810 1554
rect 880 1730 932 1740
rect 880 1554 886 1730
rect 886 1554 920 1730
rect 920 1554 932 1730
rect 880 1550 932 1554
rect 998 1730 1050 1740
rect 998 1554 1008 1730
rect 1008 1554 1042 1730
rect 1042 1554 1050 1730
rect 998 1550 1050 1554
rect 1120 1730 1172 1740
rect 1120 1554 1126 1730
rect 1126 1554 1160 1730
rect 1160 1554 1172 1730
rect 1120 1550 1172 1554
rect 1238 1730 1290 1740
rect 1238 1554 1248 1730
rect 1248 1554 1282 1730
rect 1282 1554 1290 1730
rect 1238 1550 1290 1554
rect 1360 1730 1412 1740
rect 1360 1554 1366 1730
rect 1366 1554 1400 1730
rect 1400 1554 1412 1730
rect 1360 1550 1412 1554
rect 1478 1730 1530 1740
rect 1478 1554 1488 1730
rect 1488 1554 1522 1730
rect 1522 1554 1530 1730
rect 1478 1550 1530 1554
rect 1600 1730 1652 1740
rect 1600 1554 1606 1730
rect 1606 1554 1640 1730
rect 1640 1554 1652 1730
rect 1600 1550 1652 1554
rect 1718 1730 1770 1740
rect 1718 1554 1728 1730
rect 1728 1554 1762 1730
rect 1762 1554 1770 1730
rect 1718 1550 1770 1554
rect 1840 1730 1892 1740
rect 1840 1554 1846 1730
rect 1846 1554 1880 1730
rect 1880 1554 1892 1730
rect 1840 1550 1892 1554
rect 1958 1730 2010 1740
rect 1958 1554 1968 1730
rect 1968 1554 2002 1730
rect 2002 1554 2010 1730
rect 1958 1550 2010 1554
rect 2080 1730 2132 1740
rect 2080 1554 2086 1730
rect 2086 1554 2120 1730
rect 2120 1554 2132 1730
rect 2080 1550 2132 1554
rect 2198 1730 2250 1740
rect 2198 1554 2208 1730
rect 2208 1554 2242 1730
rect 2242 1554 2250 1730
rect 2198 1550 2250 1554
rect 2320 1730 2372 1740
rect 2320 1554 2326 1730
rect 2326 1554 2360 1730
rect 2360 1554 2372 1730
rect 2320 1550 2372 1554
rect 330 1453 400 1480
rect 330 1419 347 1453
rect 347 1419 381 1453
rect 381 1419 400 1453
rect 330 1410 400 1419
rect 570 1453 640 1480
rect 570 1419 587 1453
rect 587 1419 621 1453
rect 621 1419 640 1453
rect 570 1410 640 1419
rect 810 1453 880 1480
rect 810 1419 827 1453
rect 827 1419 861 1453
rect 861 1419 880 1453
rect 810 1410 880 1419
rect 1050 1453 1120 1480
rect 1050 1419 1067 1453
rect 1067 1419 1101 1453
rect 1101 1419 1120 1453
rect 1050 1410 1120 1419
rect 1290 1453 1360 1480
rect 1290 1419 1307 1453
rect 1307 1419 1341 1453
rect 1341 1419 1360 1453
rect 1290 1410 1360 1419
rect 1530 1453 1600 1480
rect 1530 1419 1547 1453
rect 1547 1419 1581 1453
rect 1581 1419 1600 1453
rect 1530 1410 1600 1419
rect 1770 1453 1840 1480
rect 1770 1419 1787 1453
rect 1787 1419 1821 1453
rect 1821 1419 1840 1453
rect 1770 1410 1840 1419
rect 2010 1453 2080 1480
rect 2010 1419 2027 1453
rect 2027 1419 2061 1453
rect 2061 1419 2080 1453
rect 2010 1410 2080 1419
rect 38 1360 90 1370
rect 38 1184 48 1360
rect 48 1184 82 1360
rect 82 1184 90 1360
rect 38 1180 90 1184
rect 160 1360 212 1370
rect 160 1184 166 1360
rect 166 1184 200 1360
rect 200 1184 212 1360
rect 160 1180 212 1184
rect 278 1360 330 1370
rect 278 1184 288 1360
rect 288 1184 322 1360
rect 322 1184 330 1360
rect 278 1180 330 1184
rect 400 1360 452 1370
rect 400 1184 406 1360
rect 406 1184 440 1360
rect 440 1184 452 1360
rect 400 1180 452 1184
rect 518 1360 570 1370
rect 518 1184 528 1360
rect 528 1184 562 1360
rect 562 1184 570 1360
rect 518 1180 570 1184
rect 640 1360 692 1370
rect 640 1184 646 1360
rect 646 1184 680 1360
rect 680 1184 692 1360
rect 640 1180 692 1184
rect 758 1360 810 1370
rect 758 1184 768 1360
rect 768 1184 802 1360
rect 802 1184 810 1360
rect 758 1180 810 1184
rect 880 1360 932 1370
rect 880 1184 886 1360
rect 886 1184 920 1360
rect 920 1184 932 1360
rect 880 1180 932 1184
rect 998 1360 1050 1370
rect 998 1184 1008 1360
rect 1008 1184 1042 1360
rect 1042 1184 1050 1360
rect 998 1180 1050 1184
rect 1120 1360 1172 1370
rect 1120 1184 1126 1360
rect 1126 1184 1160 1360
rect 1160 1184 1172 1360
rect 1120 1180 1172 1184
rect 1238 1360 1290 1370
rect 1238 1184 1248 1360
rect 1248 1184 1282 1360
rect 1282 1184 1290 1360
rect 1238 1180 1290 1184
rect 1360 1360 1412 1370
rect 1360 1184 1366 1360
rect 1366 1184 1400 1360
rect 1400 1184 1412 1360
rect 1360 1180 1412 1184
rect 1478 1360 1530 1370
rect 1478 1184 1488 1360
rect 1488 1184 1522 1360
rect 1522 1184 1530 1360
rect 1478 1180 1530 1184
rect 1600 1360 1652 1370
rect 1600 1184 1606 1360
rect 1606 1184 1640 1360
rect 1640 1184 1652 1360
rect 1600 1180 1652 1184
rect 1718 1360 1770 1370
rect 1718 1184 1728 1360
rect 1728 1184 1762 1360
rect 1762 1184 1770 1360
rect 1718 1180 1770 1184
rect 1840 1360 1892 1370
rect 1840 1184 1846 1360
rect 1846 1184 1880 1360
rect 1880 1184 1892 1360
rect 1840 1180 1892 1184
rect 1958 1360 2010 1370
rect 1958 1184 1968 1360
rect 1968 1184 2002 1360
rect 2002 1184 2010 1360
rect 1958 1180 2010 1184
rect 2080 1360 2132 1370
rect 2080 1184 2086 1360
rect 2086 1184 2120 1360
rect 2120 1184 2132 1360
rect 2080 1180 2132 1184
rect 2198 1360 2250 1370
rect 2198 1184 2208 1360
rect 2208 1184 2242 1360
rect 2242 1184 2250 1360
rect 2198 1180 2250 1184
rect 2320 1360 2372 1370
rect 2320 1184 2326 1360
rect 2326 1184 2360 1360
rect 2360 1184 2372 1360
rect 2320 1180 2372 1184
rect 330 1083 400 1110
rect 330 1049 347 1083
rect 347 1049 381 1083
rect 381 1049 400 1083
rect 330 1040 400 1049
rect 570 1083 640 1110
rect 570 1049 587 1083
rect 587 1049 621 1083
rect 621 1049 640 1083
rect 570 1040 640 1049
rect 810 1083 880 1110
rect 810 1049 827 1083
rect 827 1049 861 1083
rect 861 1049 880 1083
rect 810 1040 880 1049
rect 1050 1083 1120 1110
rect 1050 1049 1067 1083
rect 1067 1049 1101 1083
rect 1101 1049 1120 1083
rect 1050 1040 1120 1049
rect 1290 1083 1360 1110
rect 1290 1049 1307 1083
rect 1307 1049 1341 1083
rect 1341 1049 1360 1083
rect 1290 1040 1360 1049
rect 1530 1083 1600 1110
rect 1530 1049 1547 1083
rect 1547 1049 1581 1083
rect 1581 1049 1600 1083
rect 1530 1040 1600 1049
rect 1770 1083 1840 1110
rect 1770 1049 1787 1083
rect 1787 1049 1821 1083
rect 1821 1049 1840 1083
rect 1770 1040 1840 1049
rect 2010 1083 2080 1110
rect 2010 1049 2027 1083
rect 2027 1049 2061 1083
rect 2061 1049 2080 1083
rect 2010 1040 2080 1049
rect 38 990 90 1000
rect 38 814 48 990
rect 48 814 82 990
rect 82 814 90 990
rect 38 810 90 814
rect 160 990 212 1000
rect 160 814 166 990
rect 166 814 200 990
rect 200 814 212 990
rect 160 810 212 814
rect 278 990 330 1000
rect 278 814 288 990
rect 288 814 322 990
rect 322 814 330 990
rect 278 810 330 814
rect 400 990 452 1000
rect 400 814 406 990
rect 406 814 440 990
rect 440 814 452 990
rect 400 810 452 814
rect 518 990 570 1000
rect 518 814 528 990
rect 528 814 562 990
rect 562 814 570 990
rect 518 810 570 814
rect 640 990 692 1000
rect 640 814 646 990
rect 646 814 680 990
rect 680 814 692 990
rect 640 810 692 814
rect 758 990 810 1000
rect 758 814 768 990
rect 768 814 802 990
rect 802 814 810 990
rect 758 810 810 814
rect 880 990 932 1000
rect 880 814 886 990
rect 886 814 920 990
rect 920 814 932 990
rect 880 810 932 814
rect 998 990 1050 1000
rect 998 814 1008 990
rect 1008 814 1042 990
rect 1042 814 1050 990
rect 998 810 1050 814
rect 1120 990 1172 1000
rect 1120 814 1126 990
rect 1126 814 1160 990
rect 1160 814 1172 990
rect 1120 810 1172 814
rect 1238 990 1290 1000
rect 1238 814 1248 990
rect 1248 814 1282 990
rect 1282 814 1290 990
rect 1238 810 1290 814
rect 1360 990 1412 1000
rect 1360 814 1366 990
rect 1366 814 1400 990
rect 1400 814 1412 990
rect 1360 810 1412 814
rect 1478 990 1530 1000
rect 1478 814 1488 990
rect 1488 814 1522 990
rect 1522 814 1530 990
rect 1478 810 1530 814
rect 1600 990 1652 1000
rect 1600 814 1606 990
rect 1606 814 1640 990
rect 1640 814 1652 990
rect 1600 810 1652 814
rect 1718 990 1770 1000
rect 1718 814 1728 990
rect 1728 814 1762 990
rect 1762 814 1770 990
rect 1718 810 1770 814
rect 1840 990 1892 1000
rect 1840 814 1846 990
rect 1846 814 1880 990
rect 1880 814 1892 990
rect 1840 810 1892 814
rect 1958 990 2010 1000
rect 1958 814 1968 990
rect 1968 814 2002 990
rect 2002 814 2010 990
rect 1958 810 2010 814
rect 2080 990 2132 1000
rect 2080 814 2086 990
rect 2086 814 2120 990
rect 2120 814 2132 990
rect 2080 810 2132 814
rect 2198 990 2250 1000
rect 2198 814 2208 990
rect 2208 814 2242 990
rect 2242 814 2250 990
rect 2198 810 2250 814
rect 2320 990 2372 1000
rect 2320 814 2326 990
rect 2326 814 2360 990
rect 2360 814 2372 990
rect 2320 810 2372 814
rect 38 666 90 670
rect 38 490 48 666
rect 48 490 82 666
rect 82 490 90 666
rect 38 480 90 490
rect 160 666 212 670
rect 160 490 166 666
rect 166 490 200 666
rect 200 490 212 666
rect 160 480 212 490
rect 278 666 330 670
rect 278 490 288 666
rect 288 490 322 666
rect 322 490 330 666
rect 278 480 330 490
rect 400 666 452 670
rect 400 490 406 666
rect 406 490 440 666
rect 440 490 452 666
rect 400 480 452 490
rect 518 666 570 670
rect 518 490 528 666
rect 528 490 562 666
rect 562 490 570 666
rect 518 480 570 490
rect 640 666 692 670
rect 640 490 646 666
rect 646 490 680 666
rect 680 490 692 666
rect 640 480 692 490
rect 758 666 810 670
rect 758 490 768 666
rect 768 490 802 666
rect 802 490 810 666
rect 758 480 810 490
rect 880 666 932 670
rect 880 490 886 666
rect 886 490 920 666
rect 920 490 932 666
rect 880 480 932 490
rect 998 666 1050 670
rect 998 490 1008 666
rect 1008 490 1042 666
rect 1042 490 1050 666
rect 998 480 1050 490
rect 1120 666 1172 670
rect 1120 490 1126 666
rect 1126 490 1160 666
rect 1160 490 1172 666
rect 1120 480 1172 490
rect 1238 666 1290 670
rect 1238 490 1248 666
rect 1248 490 1282 666
rect 1282 490 1290 666
rect 1238 480 1290 490
rect 330 431 400 440
rect 330 397 347 431
rect 347 397 381 431
rect 381 397 400 431
rect 330 370 400 397
rect 570 431 640 440
rect 570 397 587 431
rect 587 397 621 431
rect 621 397 640 431
rect 570 370 640 397
rect 810 431 880 440
rect 810 397 827 431
rect 827 397 861 431
rect 861 397 880 431
rect 810 370 880 397
rect 1050 431 1120 440
rect 1050 397 1067 431
rect 1067 397 1101 431
rect 1101 397 1120 431
rect 1050 370 1120 397
rect 1290 431 1360 440
rect 1290 397 1307 431
rect 1307 397 1341 431
rect 1341 397 1360 431
rect 1290 370 1360 397
rect 1478 666 1530 670
rect 1478 490 1488 666
rect 1488 490 1522 666
rect 1522 490 1530 666
rect 1478 480 1530 490
rect 1600 666 1652 670
rect 1600 490 1606 666
rect 1606 490 1640 666
rect 1640 490 1652 666
rect 1600 480 1652 490
rect 1718 666 1770 670
rect 1718 490 1728 666
rect 1728 490 1762 666
rect 1762 490 1770 666
rect 1718 480 1770 490
rect 1840 666 1892 670
rect 1840 490 1846 666
rect 1846 490 1880 666
rect 1880 490 1892 666
rect 1840 480 1892 490
rect 1958 666 2010 670
rect 1958 490 1968 666
rect 1968 490 2002 666
rect 2002 490 2010 666
rect 1958 480 2010 490
rect 2080 666 2132 670
rect 2080 490 2086 666
rect 2086 490 2120 666
rect 2120 490 2132 666
rect 2080 480 2132 490
rect 2198 666 2250 670
rect 2198 490 2208 666
rect 2208 490 2242 666
rect 2242 490 2250 666
rect 2198 480 2250 490
rect 2320 666 2372 670
rect 2320 490 2326 666
rect 2326 490 2360 666
rect 2360 490 2372 666
rect 2320 480 2372 490
rect 1530 431 1600 440
rect 1530 397 1547 431
rect 1547 397 1581 431
rect 1581 397 1600 431
rect 1530 370 1600 397
rect 1770 431 1840 440
rect 1770 397 1787 431
rect 1787 397 1821 431
rect 1821 397 1840 431
rect 1770 370 1840 397
rect 2010 431 2080 440
rect 2010 397 2027 431
rect 2027 397 2061 431
rect 2061 397 2080 431
rect 2010 370 2080 397
rect 38 296 90 300
rect 38 120 48 296
rect 48 120 82 296
rect 82 120 90 296
rect 38 110 90 120
rect 160 296 212 300
rect 160 120 166 296
rect 166 120 200 296
rect 200 120 212 296
rect 160 110 212 120
rect 278 296 330 300
rect 278 120 288 296
rect 288 120 322 296
rect 322 120 330 296
rect 278 110 330 120
rect 400 296 452 300
rect 400 120 406 296
rect 406 120 440 296
rect 440 120 452 296
rect 400 110 452 120
rect 518 296 570 300
rect 518 120 528 296
rect 528 120 562 296
rect 562 120 570 296
rect 518 110 570 120
rect 640 296 692 300
rect 640 120 646 296
rect 646 120 680 296
rect 680 120 692 296
rect 640 110 692 120
rect 758 296 810 300
rect 758 120 768 296
rect 768 120 802 296
rect 802 120 810 296
rect 758 110 810 120
rect 880 296 932 300
rect 880 120 886 296
rect 886 120 920 296
rect 920 120 932 296
rect 880 110 932 120
rect 998 296 1050 300
rect 998 120 1008 296
rect 1008 120 1042 296
rect 1042 120 1050 296
rect 998 110 1050 120
rect 1120 296 1172 300
rect 1120 120 1126 296
rect 1126 120 1160 296
rect 1160 120 1172 296
rect 1120 110 1172 120
rect 1238 296 1290 300
rect 1238 120 1248 296
rect 1248 120 1282 296
rect 1282 120 1290 296
rect 1238 110 1290 120
rect 1360 296 1412 300
rect 1360 120 1366 296
rect 1366 120 1400 296
rect 1400 120 1412 296
rect 1360 110 1412 120
rect 1478 296 1530 300
rect 1478 120 1488 296
rect 1488 120 1522 296
rect 1522 120 1530 296
rect 1478 110 1530 120
rect 1600 296 1652 300
rect 1600 120 1606 296
rect 1606 120 1640 296
rect 1640 120 1652 296
rect 1600 110 1652 120
rect 1718 296 1770 300
rect 1718 120 1728 296
rect 1728 120 1762 296
rect 1762 120 1770 296
rect 1718 110 1770 120
rect 1840 296 1892 300
rect 1840 120 1846 296
rect 1846 120 1880 296
rect 1880 120 1892 296
rect 1840 110 1892 120
rect 1958 296 2010 300
rect 1958 120 1968 296
rect 1968 120 2002 296
rect 2002 120 2010 296
rect 1958 110 2010 120
rect 2080 296 2132 300
rect 2080 120 2086 296
rect 2086 120 2120 296
rect 2120 120 2132 296
rect 2080 110 2132 120
rect 2198 296 2250 300
rect 2198 120 2208 296
rect 2208 120 2242 296
rect 2242 120 2250 296
rect 2198 110 2250 120
rect 2320 296 2372 300
rect 2320 120 2326 296
rect 2326 120 2360 296
rect 2360 120 2372 296
rect 2320 110 2372 120
rect 330 61 400 70
rect 330 27 347 61
rect 347 27 381 61
rect 381 27 400 61
rect 330 0 400 27
rect 570 61 640 70
rect 570 27 587 61
rect 587 27 621 61
rect 621 27 640 61
rect 570 0 640 27
rect 810 61 880 70
rect 810 27 827 61
rect 827 27 861 61
rect 861 27 880 61
rect 810 0 880 27
rect 1050 61 1120 70
rect 1050 27 1067 61
rect 1067 27 1101 61
rect 1101 27 1120 61
rect 1050 0 1120 27
rect 1290 61 1360 70
rect 1290 27 1307 61
rect 1307 27 1341 61
rect 1341 27 1360 61
rect 1290 0 1360 27
rect 1530 61 1600 70
rect 1530 27 1547 61
rect 1547 27 1581 61
rect 1581 27 1600 61
rect 1530 0 1600 27
rect 1770 61 1840 70
rect 1770 27 1787 61
rect 1787 27 1821 61
rect 1821 27 1840 61
rect 1770 0 1840 27
rect 2010 61 2080 70
rect 2010 27 2027 61
rect 2027 27 2061 61
rect 2061 27 2080 61
rect 2010 0 2080 27
rect 38 -74 90 -70
rect 38 -250 48 -74
rect 48 -250 82 -74
rect 82 -250 90 -74
rect 38 -260 90 -250
rect 160 -74 212 -70
rect 160 -250 166 -74
rect 166 -250 200 -74
rect 200 -250 212 -74
rect 160 -260 212 -250
rect 278 -74 330 -70
rect 278 -250 288 -74
rect 288 -250 322 -74
rect 322 -250 330 -74
rect 278 -260 330 -250
rect 400 -74 452 -70
rect 400 -250 406 -74
rect 406 -250 440 -74
rect 440 -250 452 -74
rect 400 -260 452 -250
rect 518 -74 570 -70
rect 518 -250 528 -74
rect 528 -250 562 -74
rect 562 -250 570 -74
rect 518 -260 570 -250
rect 640 -74 692 -70
rect 640 -250 646 -74
rect 646 -250 680 -74
rect 680 -250 692 -74
rect 640 -260 692 -250
rect 758 -74 810 -70
rect 758 -250 768 -74
rect 768 -250 802 -74
rect 802 -250 810 -74
rect 758 -260 810 -250
rect 880 -74 932 -70
rect 880 -250 886 -74
rect 886 -250 920 -74
rect 920 -250 932 -74
rect 880 -260 932 -250
rect 998 -74 1050 -70
rect 998 -250 1008 -74
rect 1008 -250 1042 -74
rect 1042 -250 1050 -74
rect 998 -260 1050 -250
rect 1120 -74 1172 -70
rect 1120 -250 1126 -74
rect 1126 -250 1160 -74
rect 1160 -250 1172 -74
rect 1120 -260 1172 -250
rect 1238 -74 1290 -70
rect 1238 -250 1248 -74
rect 1248 -250 1282 -74
rect 1282 -250 1290 -74
rect 1238 -260 1290 -250
rect 1360 -74 1412 -70
rect 1360 -250 1366 -74
rect 1366 -250 1400 -74
rect 1400 -250 1412 -74
rect 1360 -260 1412 -250
rect 1478 -74 1530 -70
rect 1478 -250 1488 -74
rect 1488 -250 1522 -74
rect 1522 -250 1530 -74
rect 1478 -260 1530 -250
rect 1600 -74 1652 -70
rect 1600 -250 1606 -74
rect 1606 -250 1640 -74
rect 1640 -250 1652 -74
rect 1600 -260 1652 -250
rect 1718 -74 1770 -70
rect 1718 -250 1728 -74
rect 1728 -250 1762 -74
rect 1762 -250 1770 -74
rect 1718 -260 1770 -250
rect 1840 -74 1892 -70
rect 1840 -250 1846 -74
rect 1846 -250 1880 -74
rect 1880 -250 1892 -74
rect 1840 -260 1892 -250
rect 1958 -74 2010 -70
rect 1958 -250 1968 -74
rect 1968 -250 2002 -74
rect 2002 -250 2010 -74
rect 1958 -260 2010 -250
rect 2080 -74 2132 -70
rect 2080 -250 2086 -74
rect 2086 -250 2120 -74
rect 2120 -250 2132 -74
rect 2080 -260 2132 -250
rect 2198 -74 2250 -70
rect 2198 -250 2208 -74
rect 2208 -250 2242 -74
rect 2242 -250 2250 -74
rect 2198 -260 2250 -250
rect 2320 -74 2372 -70
rect 2320 -250 2326 -74
rect 2326 -250 2360 -74
rect 2360 -250 2372 -74
rect 2320 -260 2372 -250
rect 330 -309 400 -300
rect 330 -343 347 -309
rect 347 -343 381 -309
rect 381 -343 400 -309
rect 330 -370 400 -343
rect 570 -309 640 -300
rect 570 -343 587 -309
rect 587 -343 621 -309
rect 621 -343 640 -309
rect 570 -370 640 -343
rect 810 -309 880 -300
rect 810 -343 827 -309
rect 827 -343 861 -309
rect 861 -343 880 -309
rect 810 -370 880 -343
rect 1050 -309 1120 -300
rect 1050 -343 1067 -309
rect 1067 -343 1101 -309
rect 1101 -343 1120 -309
rect 1050 -370 1120 -343
rect 1290 -309 1360 -300
rect 1290 -343 1307 -309
rect 1307 -343 1341 -309
rect 1341 -343 1360 -309
rect 1290 -370 1360 -343
rect 1530 -309 1600 -300
rect 1530 -343 1547 -309
rect 1547 -343 1581 -309
rect 1581 -343 1600 -309
rect 1530 -370 1600 -343
rect 1770 -309 1840 -300
rect 1770 -343 1787 -309
rect 1787 -343 1821 -309
rect 1821 -343 1840 -309
rect 1770 -370 1840 -343
rect 2010 -309 2080 -300
rect 2010 -343 2027 -309
rect 2027 -343 2061 -309
rect 2061 -343 2080 -309
rect 2010 -370 2080 -343
rect 38 -444 90 -440
rect 38 -620 48 -444
rect 48 -620 82 -444
rect 82 -620 90 -444
rect 38 -630 90 -620
rect 160 -444 212 -440
rect 160 -620 166 -444
rect 166 -620 200 -444
rect 200 -620 212 -444
rect 160 -630 212 -620
rect 278 -444 330 -440
rect 278 -620 288 -444
rect 288 -620 322 -444
rect 322 -620 330 -444
rect 278 -630 330 -620
rect 400 -444 452 -440
rect 400 -620 406 -444
rect 406 -620 440 -444
rect 440 -620 452 -444
rect 400 -630 452 -620
rect 518 -444 570 -440
rect 518 -620 528 -444
rect 528 -620 562 -444
rect 562 -620 570 -444
rect 518 -630 570 -620
rect 640 -444 692 -440
rect 640 -620 646 -444
rect 646 -620 680 -444
rect 680 -620 692 -444
rect 640 -630 692 -620
rect 758 -444 810 -440
rect 758 -620 768 -444
rect 768 -620 802 -444
rect 802 -620 810 -444
rect 758 -630 810 -620
rect 880 -444 932 -440
rect 880 -620 886 -444
rect 886 -620 920 -444
rect 920 -620 932 -444
rect 880 -630 932 -620
rect 998 -444 1050 -440
rect 998 -620 1008 -444
rect 1008 -620 1042 -444
rect 1042 -620 1050 -444
rect 998 -630 1050 -620
rect 1120 -444 1172 -440
rect 1120 -620 1126 -444
rect 1126 -620 1160 -444
rect 1160 -620 1172 -444
rect 1120 -630 1172 -620
rect 1238 -444 1290 -440
rect 1238 -620 1248 -444
rect 1248 -620 1282 -444
rect 1282 -620 1290 -444
rect 1238 -630 1290 -620
rect 1360 -444 1412 -440
rect 1360 -620 1366 -444
rect 1366 -620 1400 -444
rect 1400 -620 1412 -444
rect 1360 -630 1412 -620
rect 1478 -444 1530 -440
rect 1478 -620 1488 -444
rect 1488 -620 1522 -444
rect 1522 -620 1530 -444
rect 1478 -630 1530 -620
rect 1600 -444 1652 -440
rect 1600 -620 1606 -444
rect 1606 -620 1640 -444
rect 1640 -620 1652 -444
rect 1600 -630 1652 -620
rect 1718 -444 1770 -440
rect 1718 -620 1728 -444
rect 1728 -620 1762 -444
rect 1762 -620 1770 -444
rect 1718 -630 1770 -620
rect 1840 -444 1892 -440
rect 1840 -620 1846 -444
rect 1846 -620 1880 -444
rect 1880 -620 1892 -444
rect 1840 -630 1892 -620
rect 1958 -444 2010 -440
rect 1958 -620 1968 -444
rect 1968 -620 2002 -444
rect 2002 -620 2010 -444
rect 1958 -630 2010 -620
rect 2080 -444 2132 -440
rect 2080 -620 2086 -444
rect 2086 -620 2120 -444
rect 2120 -620 2132 -444
rect 2080 -630 2132 -620
rect 2198 -444 2250 -440
rect 2198 -620 2208 -444
rect 2208 -620 2242 -444
rect 2242 -620 2250 -444
rect 2198 -630 2250 -620
rect 2320 -444 2372 -440
rect 2320 -620 2326 -444
rect 2326 -620 2360 -444
rect 2360 -620 2372 -444
rect 2320 -630 2372 -620
rect 330 -679 400 -670
rect 330 -713 347 -679
rect 347 -713 381 -679
rect 381 -713 400 -679
rect 330 -740 400 -713
rect 570 -679 640 -670
rect 570 -713 587 -679
rect 587 -713 621 -679
rect 621 -713 640 -679
rect 570 -740 640 -713
rect 810 -679 880 -670
rect 810 -713 827 -679
rect 827 -713 861 -679
rect 861 -713 880 -679
rect 810 -740 880 -713
rect 1050 -679 1120 -670
rect 1050 -713 1067 -679
rect 1067 -713 1101 -679
rect 1101 -713 1120 -679
rect 1050 -740 1120 -713
rect 1290 -679 1360 -670
rect 1290 -713 1307 -679
rect 1307 -713 1341 -679
rect 1341 -713 1360 -679
rect 1290 -740 1360 -713
rect 1530 -679 1600 -670
rect 1530 -713 1547 -679
rect 1547 -713 1581 -679
rect 1581 -713 1600 -679
rect 1530 -740 1600 -713
rect 1770 -679 1840 -670
rect 1770 -713 1787 -679
rect 1787 -713 1821 -679
rect 1821 -713 1840 -679
rect 1770 -740 1840 -713
rect 2010 -679 2080 -670
rect 2010 -713 2027 -679
rect 2027 -713 2061 -679
rect 2061 -713 2080 -679
rect 2010 -740 2080 -713
rect 0 -840 2420 -800
rect 0 -860 2420 -840
<< metal2 >>
rect 450 2270 1960 2420
rect 320 2220 410 2230
rect 210 2120 280 2220
rect 320 2150 330 2220
rect 400 2150 410 2220
rect 450 2120 520 2270
rect 560 2220 650 2230
rect 800 2220 890 2230
rect 560 2150 570 2220
rect 640 2150 650 2220
rect 690 2120 760 2220
rect 800 2150 810 2220
rect 880 2150 890 2220
rect 930 2120 1000 2270
rect 1040 2220 1130 2230
rect 1280 2220 1370 2230
rect 1040 2150 1050 2220
rect 1120 2150 1130 2220
rect 1170 2120 1240 2220
rect 1280 2150 1290 2220
rect 1360 2150 1370 2220
rect 1410 2120 1480 2270
rect 1520 2220 1610 2230
rect 1760 2220 1850 2230
rect 1520 2150 1530 2220
rect 1600 2150 1610 2220
rect 1650 2120 1720 2220
rect 1760 2150 1770 2220
rect 1840 2150 1850 2220
rect 1890 2120 1960 2270
rect 2000 2220 2090 2230
rect 2000 2150 2010 2220
rect 2080 2150 2090 2220
rect 2130 2120 2200 2220
rect 30 2110 90 2120
rect 30 1920 38 2110
rect 30 1740 90 1920
rect 160 2110 330 2120
rect 212 1920 278 2110
rect 160 1910 330 1920
rect 400 2110 570 2120
rect 452 1920 518 2110
rect 400 1910 570 1920
rect 640 2110 810 2120
rect 692 1920 758 2110
rect 640 1910 810 1920
rect 880 2110 1050 2120
rect 932 1920 998 2110
rect 880 1910 1050 1920
rect 1120 2110 1290 2120
rect 1172 1920 1238 2110
rect 1120 1910 1290 1920
rect 1360 2110 1530 2120
rect 1412 1920 1478 2110
rect 1360 1910 1530 1920
rect 1600 2110 1770 2120
rect 1652 1920 1718 2110
rect 1600 1910 1770 1920
rect 1840 2110 2010 2120
rect 1892 1920 1958 2110
rect 1840 1910 2010 1920
rect 2080 2110 2250 2120
rect 2132 1920 2198 2110
rect 2080 1910 2250 1920
rect 2320 2110 2380 2120
rect 2372 1920 2380 2110
rect 210 1750 280 1910
rect 320 1850 410 1860
rect 320 1780 330 1850
rect 400 1780 410 1850
rect 450 1750 520 1910
rect 560 1850 650 1860
rect 560 1780 570 1850
rect 640 1780 650 1850
rect 690 1750 760 1910
rect 800 1850 890 1860
rect 800 1780 810 1850
rect 880 1780 890 1850
rect 930 1750 1000 1910
rect 1040 1850 1130 1860
rect 1040 1780 1050 1850
rect 1120 1780 1130 1850
rect 1170 1750 1240 1910
rect 1280 1850 1370 1860
rect 1280 1780 1290 1850
rect 1360 1780 1370 1850
rect 1410 1750 1480 1910
rect 1520 1850 1610 1860
rect 1520 1780 1530 1850
rect 1600 1780 1610 1850
rect 1650 1750 1720 1910
rect 1760 1850 1850 1860
rect 1760 1780 1770 1850
rect 1840 1780 1850 1850
rect 1890 1750 1960 1910
rect 2000 1850 2090 1860
rect 2000 1780 2010 1850
rect 2080 1780 2090 1850
rect 2130 1750 2200 1910
rect 30 1550 38 1740
rect 30 1370 90 1550
rect 160 1740 330 1750
rect 212 1550 278 1740
rect 160 1540 330 1550
rect 400 1740 570 1750
rect 452 1550 518 1740
rect 400 1540 570 1550
rect 640 1740 810 1750
rect 692 1550 758 1740
rect 640 1540 810 1550
rect 880 1740 1050 1750
rect 932 1550 998 1740
rect 880 1540 1050 1550
rect 1120 1740 1290 1750
rect 1172 1550 1238 1740
rect 1120 1540 1290 1550
rect 1360 1740 1530 1750
rect 1412 1550 1478 1740
rect 1360 1540 1530 1550
rect 1600 1740 1770 1750
rect 1652 1550 1718 1740
rect 1600 1540 1770 1550
rect 1840 1740 2010 1750
rect 1892 1550 1958 1740
rect 1840 1540 2010 1550
rect 2080 1740 2250 1750
rect 2132 1550 2198 1740
rect 2080 1540 2250 1550
rect 2320 1740 2380 1920
rect 2372 1550 2380 1740
rect 210 1380 280 1540
rect 320 1480 410 1490
rect 320 1410 330 1480
rect 400 1410 410 1480
rect 450 1380 520 1540
rect 560 1480 650 1490
rect 560 1410 570 1480
rect 640 1410 650 1480
rect 690 1380 760 1540
rect 800 1480 890 1490
rect 800 1410 810 1480
rect 880 1410 890 1480
rect 930 1380 1000 1540
rect 1040 1480 1130 1490
rect 1040 1410 1050 1480
rect 1120 1410 1130 1480
rect 1170 1380 1240 1540
rect 1280 1480 1370 1490
rect 1280 1410 1290 1480
rect 1360 1410 1370 1480
rect 1410 1380 1480 1540
rect 1520 1480 1610 1490
rect 1520 1410 1530 1480
rect 1600 1410 1610 1480
rect 1650 1380 1720 1540
rect 1760 1480 1850 1490
rect 1760 1410 1770 1480
rect 1840 1410 1850 1480
rect 1890 1380 1960 1540
rect 2000 1480 2090 1490
rect 2000 1410 2010 1480
rect 2080 1410 2090 1480
rect 2130 1380 2200 1540
rect 30 1180 38 1370
rect 30 1000 90 1180
rect 160 1370 330 1380
rect 212 1180 278 1370
rect 160 1170 330 1180
rect 400 1370 570 1380
rect 452 1180 518 1370
rect 400 1170 570 1180
rect 640 1370 810 1380
rect 692 1180 758 1370
rect 640 1170 810 1180
rect 880 1370 1050 1380
rect 932 1180 998 1370
rect 880 1170 1050 1180
rect 1120 1370 1290 1380
rect 1172 1180 1238 1370
rect 1120 1170 1290 1180
rect 1360 1370 1530 1380
rect 1412 1180 1478 1370
rect 1360 1170 1530 1180
rect 1600 1370 1770 1380
rect 1652 1180 1718 1370
rect 1600 1170 1770 1180
rect 1840 1370 2010 1380
rect 1892 1180 1958 1370
rect 1840 1170 2010 1180
rect 2080 1370 2250 1380
rect 2132 1180 2198 1370
rect 2080 1170 2250 1180
rect 2320 1370 2380 1550
rect 2372 1180 2380 1370
rect 210 1010 280 1170
rect 320 1110 410 1120
rect 320 1040 330 1110
rect 400 1040 410 1110
rect 450 1010 520 1170
rect 560 1110 650 1120
rect 560 1040 570 1110
rect 640 1040 650 1110
rect 690 1010 760 1170
rect 800 1110 890 1120
rect 800 1040 810 1110
rect 880 1040 890 1110
rect 930 1010 1000 1170
rect 1040 1110 1130 1120
rect 1040 1040 1050 1110
rect 1120 1040 1130 1110
rect 1170 1010 1240 1170
rect 1280 1110 1370 1120
rect 1280 1040 1290 1110
rect 1360 1040 1370 1110
rect 1410 1010 1480 1170
rect 1520 1110 1610 1120
rect 1520 1040 1530 1110
rect 1600 1040 1610 1110
rect 1650 1010 1720 1170
rect 1760 1110 1850 1120
rect 1760 1040 1770 1110
rect 1840 1040 1850 1110
rect 1890 1010 1960 1170
rect 2000 1110 2090 1120
rect 2000 1040 2010 1110
rect 2080 1040 2090 1110
rect 2130 1010 2200 1170
rect 30 810 38 1000
rect 30 670 90 810
rect 160 1000 330 1010
rect 212 810 278 1000
rect 160 800 330 810
rect 400 1000 570 1010
rect 452 810 518 1000
rect 400 800 570 810
rect 640 1000 810 1010
rect 692 810 758 1000
rect 640 800 810 810
rect 880 1000 1050 1010
rect 932 810 998 1000
rect 880 800 1050 810
rect 1120 1000 1290 1010
rect 1172 810 1238 1000
rect 1120 800 1290 810
rect 1360 1000 1530 1010
rect 1412 810 1478 1000
rect 1360 800 1530 810
rect 1600 1000 1770 1010
rect 1652 810 1718 1000
rect 1600 800 1770 810
rect 1840 1000 2010 1010
rect 1892 810 1958 1000
rect 1840 800 2010 810
rect 2080 1000 2250 1010
rect 2132 810 2198 1000
rect 2080 800 2250 810
rect 2320 1000 2380 1180
rect 2372 810 2380 1000
rect 210 680 280 800
rect 450 680 520 800
rect 690 680 760 800
rect 930 680 1000 800
rect 1170 680 1240 800
rect 1410 680 1480 800
rect 1650 680 1720 800
rect 1890 680 1960 800
rect 2130 680 2200 800
rect 30 480 38 670
rect 30 300 90 480
rect 160 670 330 680
rect 212 480 278 670
rect 160 470 330 480
rect 400 670 570 680
rect 452 480 518 670
rect 400 470 570 480
rect 640 670 810 680
rect 692 480 758 670
rect 640 470 810 480
rect 880 670 1050 680
rect 932 480 998 670
rect 880 470 1050 480
rect 1120 670 1290 680
rect 1172 480 1238 670
rect 1120 470 1290 480
rect 1410 670 1530 680
rect 1410 480 1478 670
rect 1410 470 1530 480
rect 1600 670 1770 680
rect 1652 480 1718 670
rect 1600 470 1770 480
rect 1840 670 2010 680
rect 1892 480 1958 670
rect 1840 470 2010 480
rect 2080 670 2250 680
rect 2132 480 2198 670
rect 2080 470 2250 480
rect 2320 670 2380 810
rect 2372 480 2380 670
rect 210 310 280 470
rect 320 370 330 440
rect 400 370 410 440
rect 320 360 410 370
rect 450 310 520 470
rect 560 370 570 440
rect 640 370 650 440
rect 560 360 650 370
rect 690 310 760 470
rect 800 370 810 440
rect 880 370 890 440
rect 800 360 890 370
rect 930 310 1000 470
rect 1040 370 1050 440
rect 1120 370 1130 440
rect 1040 360 1130 370
rect 1170 310 1240 470
rect 1280 370 1290 440
rect 1360 370 1370 440
rect 1280 360 1370 370
rect 1410 310 1480 470
rect 1520 370 1530 440
rect 1600 370 1610 440
rect 1520 360 1610 370
rect 1650 310 1720 470
rect 1760 370 1770 440
rect 1840 370 1850 440
rect 1760 360 1850 370
rect 1890 310 1960 470
rect 2000 370 2010 440
rect 2080 370 2090 440
rect 2000 360 2090 370
rect 2130 310 2200 470
rect 30 110 38 300
rect 30 -70 90 110
rect 160 300 330 310
rect 212 110 278 300
rect 160 100 330 110
rect 400 300 570 310
rect 452 110 518 300
rect 400 100 570 110
rect 640 300 810 310
rect 692 110 758 300
rect 640 100 810 110
rect 880 300 1050 310
rect 932 110 998 300
rect 880 100 1050 110
rect 1120 300 1290 310
rect 1172 110 1238 300
rect 1120 100 1290 110
rect 1360 300 1530 310
rect 1412 110 1478 300
rect 1360 100 1530 110
rect 1600 300 1770 310
rect 1652 110 1718 300
rect 1600 100 1770 110
rect 1840 300 2010 310
rect 1892 110 1958 300
rect 1840 100 2010 110
rect 2080 300 2250 310
rect 2132 110 2198 300
rect 2080 100 2250 110
rect 2320 300 2380 480
rect 2372 110 2380 300
rect 210 -60 280 100
rect 320 0 330 70
rect 400 0 410 70
rect 320 -10 410 0
rect 450 -60 520 100
rect 560 0 570 70
rect 640 0 650 70
rect 560 -10 650 0
rect 690 -60 760 100
rect 800 0 810 70
rect 880 0 890 70
rect 800 -10 890 0
rect 930 -60 1000 100
rect 1040 0 1050 70
rect 1120 0 1130 70
rect 1040 -10 1130 0
rect 1170 -60 1240 100
rect 1280 0 1290 70
rect 1360 0 1370 70
rect 1280 -10 1370 0
rect 1410 -60 1480 100
rect 1520 0 1530 70
rect 1600 0 1610 70
rect 1520 -10 1610 0
rect 1650 -60 1720 100
rect 1760 0 1770 70
rect 1840 0 1850 70
rect 1760 -10 1850 0
rect 1890 -60 1960 100
rect 2000 0 2010 70
rect 2080 0 2090 70
rect 2000 -10 2090 0
rect 2130 -60 2200 100
rect 30 -260 38 -70
rect 30 -440 90 -260
rect 160 -70 330 -60
rect 212 -260 278 -70
rect 160 -270 330 -260
rect 400 -70 570 -60
rect 452 -260 518 -70
rect 400 -270 570 -260
rect 640 -70 810 -60
rect 692 -260 758 -70
rect 640 -270 810 -260
rect 880 -70 1050 -60
rect 932 -260 998 -70
rect 880 -270 1050 -260
rect 1120 -70 1290 -60
rect 1172 -260 1238 -70
rect 1120 -270 1290 -260
rect 1360 -70 1530 -60
rect 1412 -260 1478 -70
rect 1360 -270 1530 -260
rect 1600 -70 1770 -60
rect 1652 -260 1718 -70
rect 1600 -270 1770 -260
rect 1840 -70 2010 -60
rect 1892 -260 1958 -70
rect 1840 -270 2010 -260
rect 2080 -70 2250 -60
rect 2132 -260 2198 -70
rect 2080 -270 2250 -260
rect 2320 -70 2380 110
rect 2372 -260 2380 -70
rect 210 -430 280 -270
rect 320 -370 330 -300
rect 400 -370 410 -300
rect 320 -380 410 -370
rect 450 -430 520 -270
rect 560 -370 570 -300
rect 640 -370 650 -300
rect 560 -380 650 -370
rect 690 -430 760 -270
rect 800 -370 810 -300
rect 880 -370 890 -300
rect 800 -380 890 -370
rect 930 -430 1000 -270
rect 1040 -370 1050 -300
rect 1120 -370 1130 -300
rect 1040 -380 1130 -370
rect 1170 -430 1240 -270
rect 1280 -370 1290 -300
rect 1360 -370 1370 -300
rect 1280 -380 1370 -370
rect 1410 -430 1480 -270
rect 1520 -370 1530 -300
rect 1600 -370 1610 -300
rect 1520 -380 1610 -370
rect 1650 -430 1720 -270
rect 1760 -370 1770 -300
rect 1840 -370 1850 -300
rect 1760 -380 1850 -370
rect 1890 -430 1960 -270
rect 2000 -370 2010 -300
rect 2080 -370 2090 -300
rect 2000 -380 2090 -370
rect 2130 -430 2200 -270
rect 30 -630 38 -440
rect 30 -780 90 -630
rect 160 -440 330 -430
rect 212 -630 278 -440
rect 160 -640 330 -630
rect 400 -440 570 -430
rect 452 -630 518 -440
rect 400 -640 570 -630
rect 640 -440 810 -430
rect 692 -630 758 -440
rect 640 -640 810 -630
rect 880 -440 1050 -430
rect 932 -630 998 -440
rect 880 -640 1050 -630
rect 1120 -440 1290 -430
rect 1172 -630 1238 -440
rect 1120 -640 1290 -630
rect 1360 -440 1530 -430
rect 1412 -630 1478 -440
rect 1360 -640 1530 -630
rect 1600 -440 1770 -430
rect 1652 -630 1718 -440
rect 1600 -640 1770 -630
rect 1840 -440 2010 -430
rect 1892 -630 1958 -440
rect 1840 -640 2010 -630
rect 2080 -440 2250 -430
rect 2132 -630 2198 -440
rect 2080 -640 2250 -630
rect 2320 -440 2380 -260
rect 2372 -630 2380 -440
rect 210 -780 280 -640
rect 320 -740 330 -670
rect 400 -740 410 -670
rect 450 -740 520 -640
rect 560 -740 570 -670
rect 640 -740 650 -670
rect 320 -750 410 -740
rect 560 -750 650 -740
rect 690 -780 760 -640
rect 800 -740 810 -670
rect 880 -740 890 -670
rect 930 -740 1000 -640
rect 1040 -740 1050 -670
rect 1120 -740 1130 -670
rect 800 -750 890 -740
rect 1040 -750 1130 -740
rect 1170 -780 1240 -640
rect 1280 -740 1290 -670
rect 1360 -740 1370 -670
rect 1410 -740 1480 -640
rect 1520 -740 1530 -670
rect 1600 -740 1610 -670
rect 1280 -750 1370 -740
rect 1520 -750 1610 -740
rect 1650 -780 1720 -640
rect 1760 -740 1770 -670
rect 1840 -740 1850 -670
rect 1890 -740 1960 -640
rect 2000 -740 2010 -670
rect 2080 -740 2090 -670
rect 1760 -750 1850 -740
rect 2000 -750 2090 -740
rect 2130 -780 2200 -640
rect 2320 -780 2380 -630
rect -20 -800 2440 -780
rect -20 -860 0 -800
rect 2420 -860 2440 -800
rect -20 -880 2440 -860
<< via2 >>
rect 330 2160 400 2220
rect 570 2160 640 2220
rect 810 2160 880 2220
rect 1050 2160 1120 2220
rect 1290 2160 1360 2220
rect 1530 2160 1600 2220
rect 1770 2160 1840 2220
rect 2010 2160 2080 2220
rect 330 1790 400 1850
rect 570 1790 640 1850
rect 810 1790 880 1850
rect 1050 1790 1120 1850
rect 1290 1790 1360 1850
rect 1530 1790 1600 1850
rect 1770 1790 1840 1850
rect 2010 1790 2080 1850
rect 330 1420 400 1480
rect 570 1420 640 1480
rect 810 1420 880 1480
rect 1050 1420 1120 1480
rect 1290 1420 1360 1480
rect 1530 1420 1600 1480
rect 1770 1420 1840 1480
rect 2010 1420 2080 1480
rect 330 1050 400 1110
rect 570 1050 640 1110
rect 810 1050 880 1110
rect 1050 1050 1120 1110
rect 1290 1050 1360 1110
rect 1530 1050 1600 1110
rect 1770 1050 1840 1110
rect 2010 1050 2080 1110
rect 330 370 400 430
rect 570 370 640 430
rect 810 370 880 430
rect 1050 370 1120 430
rect 1290 370 1360 430
rect 1530 370 1600 430
rect 1770 370 1840 430
rect 2010 370 2080 430
rect 330 0 400 60
rect 570 0 640 60
rect 810 0 880 60
rect 1050 0 1120 60
rect 1290 0 1360 60
rect 1530 0 1600 60
rect 1770 0 1840 60
rect 2010 0 2080 60
rect 330 -370 400 -310
rect 570 -370 640 -310
rect 810 -370 880 -310
rect 1050 -370 1120 -310
rect 1290 -370 1360 -310
rect 1530 -370 1600 -310
rect 1770 -370 1840 -310
rect 2010 -370 2080 -310
rect 330 -740 400 -680
rect 570 -740 640 -680
rect 810 -740 880 -680
rect 1050 -740 1120 -680
rect 1290 -740 1360 -680
rect 1530 -740 1600 -680
rect 1770 -740 1840 -680
rect 2010 -740 2080 -680
<< metal3 >>
rect 320 2220 2330 2230
rect 320 2160 330 2220
rect 400 2160 570 2220
rect 640 2160 810 2220
rect 880 2160 1050 2220
rect 1120 2160 1290 2220
rect 1360 2160 1530 2220
rect 1600 2160 1770 2220
rect 1840 2160 2010 2220
rect 2080 2160 2330 2220
rect 320 2150 2330 2160
rect 2240 1860 2330 2150
rect 2400 1880 2560 1890
rect 2400 1860 2420 1880
rect 320 1850 2420 1860
rect 320 1790 330 1850
rect 400 1790 570 1850
rect 640 1790 810 1850
rect 880 1790 1050 1850
rect 1120 1790 1290 1850
rect 1360 1790 1530 1850
rect 1600 1790 1770 1850
rect 1840 1790 2010 1850
rect 2080 1790 2420 1850
rect 320 1780 2420 1790
rect 2400 1760 2420 1780
rect 2550 1860 2560 1880
rect 2550 1780 2590 1860
rect 2550 1760 2560 1780
rect 2400 1750 2560 1760
rect 2200 1510 2350 1520
rect 2200 1490 2210 1510
rect 320 1480 2210 1490
rect 320 1420 330 1480
rect 400 1420 570 1480
rect 640 1420 810 1480
rect 880 1420 1050 1480
rect 1120 1420 1290 1480
rect 1360 1420 1530 1480
rect 1600 1420 1770 1480
rect 1840 1420 2010 1480
rect 2080 1420 2210 1480
rect 320 1410 2210 1420
rect 2200 1390 2210 1410
rect 2340 1490 2350 1510
rect 2340 1410 2590 1490
rect 2340 1390 2350 1410
rect 2200 1380 2350 1390
rect 560 1230 1850 1310
rect 560 1120 650 1230
rect 1760 1120 1850 1230
rect 1990 1250 2140 1260
rect 1990 1130 2000 1250
rect 2130 1130 2140 1250
rect 1990 1120 2140 1130
rect 320 1110 650 1120
rect 320 1050 330 1110
rect 400 1050 570 1110
rect 640 1050 650 1110
rect 320 1040 650 1050
rect 800 1110 1610 1120
rect 800 1050 810 1110
rect 880 1050 1050 1110
rect 1120 1050 1290 1110
rect 1360 1050 1530 1110
rect 1600 1050 1610 1110
rect 800 1040 1610 1050
rect 1760 1110 2590 1120
rect 1760 1050 1770 1110
rect 1840 1050 2010 1110
rect 2080 1050 2590 1110
rect 1760 1040 2590 1050
rect 1520 980 1610 1040
rect 1520 910 2590 980
rect 1040 780 2590 850
rect 1040 440 1130 780
rect 320 430 650 440
rect 320 370 330 430
rect 400 370 570 430
rect 640 370 650 430
rect 320 360 650 370
rect 800 430 1130 440
rect 800 370 810 430
rect 880 370 1050 430
rect 1120 370 1130 430
rect 800 360 1130 370
rect 1280 650 2590 720
rect 1280 430 1370 650
rect 1280 370 1290 430
rect 1360 370 1370 430
rect 1280 360 1370 370
rect 1520 510 2590 580
rect 1520 430 1610 510
rect 1520 370 1530 430
rect 1600 370 1610 430
rect 1520 360 1610 370
rect 1760 430 2140 440
rect 1760 370 1770 430
rect 1840 370 2010 430
rect 2080 370 2140 430
rect 1760 360 2140 370
rect 560 250 650 360
rect 1760 250 1850 360
rect 560 170 1850 250
rect 1990 350 2140 360
rect 1990 230 2000 350
rect 2130 230 2140 350
rect 1990 220 2140 230
rect 2200 90 2350 100
rect 2200 70 2210 90
rect 320 60 2210 70
rect 320 0 330 60
rect 400 0 570 60
rect 640 0 810 60
rect 880 0 1050 60
rect 1120 0 1290 60
rect 1360 0 1530 60
rect 1600 0 1770 60
rect 1840 0 2010 60
rect 2080 0 2210 60
rect 320 -10 2210 0
rect 2200 -30 2210 -10
rect 2340 -30 2350 90
rect 2200 -40 2350 -30
rect 2410 -280 2560 -270
rect 2410 -300 2420 -280
rect 320 -310 2420 -300
rect 320 -370 330 -310
rect 400 -370 570 -310
rect 640 -370 810 -310
rect 880 -370 1050 -310
rect 1120 -370 1290 -310
rect 1360 -370 1530 -310
rect 1600 -370 1770 -310
rect 1840 -370 2010 -310
rect 2080 -370 2420 -310
rect 320 -380 2420 -370
rect 2240 -670 2330 -380
rect 2410 -400 2420 -380
rect 2550 -400 2560 -280
rect 2410 -410 2560 -400
rect 320 -680 2330 -670
rect 320 -740 330 -680
rect 400 -740 570 -680
rect 640 -740 810 -680
rect 880 -740 1050 -680
rect 1120 -740 1290 -680
rect 1360 -740 1530 -680
rect 1600 -740 1770 -680
rect 1840 -740 2010 -680
rect 2080 -740 2330 -680
rect 320 -750 2330 -740
<< via3 >>
rect 2420 1760 2550 1880
rect 2210 1390 2340 1510
rect 2000 1130 2130 1250
rect 2000 230 2130 350
rect 2210 -30 2340 90
rect 2420 -400 2550 -280
<< metal4 >>
rect 2410 1880 2560 1890
rect 2410 1760 2420 1880
rect 2550 1760 2560 1880
rect 2200 1510 2350 1520
rect 2200 1390 2210 1510
rect 2340 1390 2350 1510
rect 1990 1250 2140 1260
rect 1990 1130 2000 1250
rect 2130 1130 2140 1250
rect 1990 350 2140 1130
rect 1990 230 2000 350
rect 2130 230 2140 350
rect 1990 220 2140 230
rect 2200 90 2350 1390
rect 2200 -30 2210 90
rect 2340 -30 2350 90
rect 2200 -40 2350 -30
rect 2410 -280 2560 1760
rect 2410 -400 2420 -280
rect 2550 -400 2560 -280
rect 2410 -410 2560 -400
<< labels >>
rlabel metal3 2570 1780 2590 1860 1 G32
rlabel metal3 2570 1410 2590 1490 1 G16
rlabel metal3 2570 1040 2590 1120 1 G8
rlabel metal3 2570 910 2590 980 1 G4
rlabel metal3 2570 780 2590 850 1 G2
rlabel metal3 2570 650 2590 720 1 IREF
rlabel metal3 2570 510 2590 580 1 G1
rlabel metal2 30 -880 2380 -780 1 VHI
rlabel metal2 450 2270 1960 2370 1 IOUT
<< end >>
