magic
tech sky130B
magscale 1 2
timestamp 1662001208
<< locali >>
rect -3600 8560 -2120 8580
rect -3600 8400 -3580 8560
rect -2140 8400 -2120 8560
rect -3600 8380 -2120 8400
rect -1400 7060 -1240 7080
rect -1400 5700 -1380 7060
rect -1260 5700 -1240 7060
rect -1400 5680 -1240 5700
rect -4560 -630 -4400 -620
rect -4560 -640 -4340 -630
rect -4560 -2220 -4540 -640
rect -4420 -2040 -4340 -640
rect -4420 -2060 -3720 -2040
rect -3740 -2220 -3720 -2060
rect -4560 -2240 -3720 -2220
<< viali >>
rect -3480 8820 -3320 8980
rect -2360 8660 -2260 8820
rect -3580 8400 -2140 8560
rect -1380 5700 -1260 7060
rect -960 6880 -840 7000
rect -1160 5780 -1040 5900
rect -4540 -2060 -4420 -640
rect -4260 -860 -4140 -720
rect -3940 -860 -3820 -720
rect -4540 -2220 -3740 -2060
<< metal1 >>
rect -3500 8980 -3300 9000
rect -3500 8820 -3480 8980
rect -3320 8820 -3300 8980
rect -3500 8800 -3300 8820
rect -2380 8820 -2240 8840
rect -4800 8600 -4000 8700
rect -2380 8660 -2360 8820
rect -2260 8660 -2240 8820
rect -2380 8640 -2240 8660
rect -1800 8780 3000 8800
rect -1800 8620 -1780 8780
rect -1620 8620 3000 8780
rect -1800 8600 3000 8620
rect -4800 7800 -4700 8600
rect -4500 8580 -4380 8600
rect -4120 8580 -4000 8600
rect -4500 8320 -4400 8580
rect -4100 8560 -2120 8580
rect -4100 8400 -3580 8560
rect -2140 8500 -2120 8560
rect -2140 8400 -150 8500
rect -4100 8320 -1400 8400
rect -4500 8300 -4380 8320
rect -4120 8300 -1400 8320
rect -700 8300 -150 8400
rect -4500 8200 -150 8300
rect -4500 8100 -1400 8200
rect -700 8100 -150 8200
rect -4500 8080 -4380 8100
rect -4120 8080 -3880 8100
rect -3620 8080 -3380 8100
rect -3120 8080 -2880 8100
rect -2620 8080 -2380 8100
rect -2120 8080 -1880 8100
rect -1620 8080 -150 8100
rect -4500 7820 -4400 8080
rect -4100 7820 -3900 8080
rect -3600 7820 -3400 8080
rect -3100 7820 -2900 8080
rect -2600 7820 -2400 8080
rect -2100 7820 -1900 8080
rect -1600 8000 -150 8080
rect -1600 7900 -1400 8000
rect -700 7900 -150 8000
rect -1600 7820 -150 7900
rect -4500 7800 -4380 7820
rect -4120 7800 -3880 7820
rect -3620 7800 -3380 7820
rect -3120 7800 -2880 7820
rect -2620 7800 -2380 7820
rect -2120 7800 -1880 7820
rect -1620 7800 -150 7820
rect -4800 7700 -1400 7800
rect -700 7700 -150 7800
rect -2500 7600 -150 7700
rect -2500 7580 -2380 7600
rect -2120 7580 -1880 7600
rect -1620 7580 -1400 7600
rect -2500 7320 -2400 7580
rect -2100 7320 -1900 7580
rect -1600 7500 -1400 7580
rect -700 7500 -150 7600
rect -1600 7400 -150 7500
rect 1100 8200 1860 8500
rect 1100 8180 1320 8200
rect 1580 8180 1860 8200
rect 1100 7920 1300 8180
rect 1600 7920 1860 8180
rect 1100 7900 1320 7920
rect 1580 7900 1860 7920
rect 1100 7700 1860 7900
rect 1100 7680 1320 7700
rect 1580 7680 1860 7700
rect 1100 7420 1300 7680
rect 1600 7420 1860 7680
rect 1100 7400 1320 7420
rect 1580 7400 1860 7420
rect -1600 7320 -1240 7400
rect -2500 7300 -2380 7320
rect -2120 7300 -1880 7320
rect -1620 7300 -1240 7320
rect -2500 7180 -1240 7300
rect -2500 7110 -2350 7180
rect -2150 7110 -1850 7180
rect -1650 7110 -1240 7180
rect -2500 7100 -1240 7110
rect -2500 7080 -2380 7100
rect -2120 7080 -1880 7100
rect -1620 7080 -1240 7100
rect -2500 7050 -2400 7080
rect -2500 6850 -2480 7050
rect -2410 6850 -2400 7050
rect -2500 6820 -2400 6850
rect -2100 7050 -1900 7080
rect -2100 6850 -2090 7050
rect -2020 6850 -1980 7050
rect -1910 6850 -1900 7050
rect -2100 6820 -1900 6850
rect -1600 7060 -1240 7080
rect -1600 7050 -1380 7060
rect -1600 6850 -1590 7050
rect -1520 6850 -1380 7050
rect -1600 6820 -1380 6850
rect -2500 6800 -2380 6820
rect -2120 6800 -1880 6820
rect -1620 6800 -1380 6820
rect -2500 6790 -1380 6800
rect -2500 6720 -2350 6790
rect -2150 6720 -1850 6790
rect -1650 6720 -1380 6790
rect -2500 6680 -1380 6720
rect -2500 6610 -2350 6680
rect -2150 6610 -1850 6680
rect -1650 6610 -1380 6680
rect -2500 6600 -1380 6610
rect -2500 6580 -2380 6600
rect -2120 6580 -1880 6600
rect -1620 6580 -1380 6600
rect -2500 6550 -2400 6580
rect -2500 6350 -2480 6550
rect -2410 6350 -2400 6550
rect -2500 6320 -2400 6350
rect -2100 6550 -1900 6580
rect -2100 6350 -2090 6550
rect -2020 6350 -1980 6550
rect -1910 6350 -1900 6550
rect -2100 6320 -1900 6350
rect -1600 6550 -1380 6580
rect -1600 6350 -1590 6550
rect -1520 6350 -1380 6550
rect -1600 6320 -1380 6350
rect -2500 6300 -2380 6320
rect -2120 6300 -1880 6320
rect -1620 6300 -1380 6320
rect -2500 6290 -1380 6300
rect -2500 6220 -2350 6290
rect -2150 6220 -1850 6290
rect -1650 6220 -1380 6290
rect -2500 6200 -1380 6220
rect -4000 6180 -1380 6200
rect -4000 6110 -3850 6180
rect -3650 6110 -3350 6180
rect -3150 6110 -2850 6180
rect -2650 6110 -2350 6180
rect -2150 6110 -1850 6180
rect -1650 6110 -1380 6180
rect -4000 6100 -1380 6110
rect -4000 6080 -3880 6100
rect -3620 6080 -3380 6100
rect -3120 6080 -2880 6100
rect -2620 6080 -2380 6100
rect -2120 6080 -1880 6100
rect -1620 6080 -1380 6100
rect -4000 6050 -3900 6080
rect -4000 5850 -3980 6050
rect -3910 5850 -3900 6050
rect -4000 5820 -3900 5850
rect -3600 6050 -3400 6080
rect -3600 5850 -3590 6050
rect -3520 5850 -3480 6050
rect -3410 5850 -3400 6050
rect -3600 5820 -3400 5850
rect -3100 6050 -2900 6080
rect -3100 5850 -3090 6050
rect -3020 5850 -2980 6050
rect -2910 5850 -2900 6050
rect -3100 5820 -2900 5850
rect -2600 6050 -2400 6080
rect -2600 5850 -2590 6050
rect -2520 5850 -2480 6050
rect -2410 5850 -2400 6050
rect -2600 5820 -2400 5850
rect -2100 6050 -1900 6080
rect -2100 5850 -2090 6050
rect -2020 5850 -1980 6050
rect -1910 5850 -1900 6050
rect -2100 5820 -1900 5850
rect -1600 6050 -1380 6080
rect -1600 5850 -1590 6050
rect -1520 5850 -1380 6050
rect -1600 5820 -1380 5850
rect -4000 5800 -3880 5820
rect -3620 5800 -3380 5820
rect -3120 5800 -2880 5820
rect -2620 5800 -2380 5820
rect -2120 5800 -1880 5820
rect -1620 5800 -1380 5820
rect -4000 5790 -1380 5800
rect -4000 5720 -3850 5790
rect -3650 5720 -3350 5790
rect -3150 5720 -2850 5790
rect -2650 5720 -2350 5790
rect -2150 5720 -1850 5790
rect -1650 5720 -1380 5790
rect -4000 5700 -1380 5720
rect -1260 5700 -1240 7060
rect 1100 7200 1860 7400
rect 1100 7180 1320 7200
rect 1580 7180 1860 7200
rect -1000 7020 -800 7040
rect -1000 6860 -980 7020
rect -820 6860 -800 7020
rect -1000 6840 -800 6860
rect 1100 6920 1300 7180
rect 1600 6920 1860 7180
rect 1100 6900 1320 6920
rect 1580 6900 1860 6920
rect 1100 6700 1860 6900
rect 1100 6680 1320 6700
rect 1580 6680 1860 6700
rect 1100 6420 1300 6680
rect 1600 6420 1860 6680
rect 1100 6400 1320 6420
rect 1580 6400 1860 6420
rect 1100 6200 1860 6400
rect 1100 6180 1320 6200
rect 1580 6180 1860 6200
rect -1200 5920 -1000 5940
rect -1200 5760 -1180 5920
rect -1020 5760 -1000 5920
rect 1100 5920 1300 6180
rect 1600 5920 1860 6180
rect 1100 5900 1320 5920
rect 1580 5900 1860 5920
rect 3100 8200 3800 8500
rect 3100 8180 3320 8200
rect 3580 8180 3800 8200
rect 3100 7920 3300 8180
rect 3600 7920 3800 8180
rect 3100 7900 3320 7920
rect 3580 7900 3800 7920
rect 3100 7700 3800 7900
rect 3100 7680 3320 7700
rect 3580 7680 3800 7700
rect 3100 7420 3300 7680
rect 3600 7420 3800 7680
rect 3100 7400 3320 7420
rect 3580 7400 3800 7420
rect 3100 7200 3800 7400
rect 3100 7180 3320 7200
rect 3580 7180 3800 7200
rect 3100 6920 3300 7180
rect 3600 6920 3800 7180
rect 3100 6900 3320 6920
rect 3580 6900 3800 6920
rect 3100 6700 3800 6900
rect 3100 6680 3320 6700
rect 3580 6680 3800 6700
rect 3100 6420 3300 6680
rect 3600 6420 3800 6680
rect 3100 6400 3320 6420
rect 3580 6400 3800 6420
rect 3100 6200 3800 6400
rect 3100 6180 3320 6200
rect 3580 6180 3800 6200
rect 3100 5920 3300 6180
rect 3600 5920 3800 6180
rect 3100 5900 3320 5920
rect 3580 5900 3800 5920
rect -1200 5740 -1000 5760
rect 500 5700 4000 5900
rect -4000 5680 -500 5700
rect -4000 5610 -3850 5680
rect -3650 5610 -3350 5680
rect -3150 5610 -2850 5680
rect -2650 5610 -2350 5680
rect -2150 5610 -500 5680
rect -4000 5600 -500 5610
rect -4000 5580 -3880 5600
rect -3620 5580 -3380 5600
rect -3120 5580 -2880 5600
rect -2620 5580 -2380 5600
rect -2120 5580 -1880 5600
rect -1620 5580 -1380 5600
rect -1120 5580 -880 5600
rect -620 5580 -500 5600
rect -4000 5550 -3900 5580
rect -4000 5350 -3980 5550
rect -3910 5350 -3900 5550
rect -4000 5320 -3900 5350
rect -3600 5550 -3400 5580
rect -3600 5350 -3590 5550
rect -3520 5350 -3480 5550
rect -3410 5350 -3400 5550
rect -3600 5320 -3400 5350
rect -3100 5550 -2900 5580
rect -3100 5350 -3090 5550
rect -3020 5350 -2980 5550
rect -2910 5350 -2900 5550
rect -3100 5320 -2900 5350
rect -2600 5550 -2400 5580
rect -2600 5350 -2590 5550
rect -2520 5350 -2480 5550
rect -2410 5350 -2400 5550
rect -2600 5320 -2400 5350
rect -2100 5550 -1900 5580
rect -2100 5350 -2090 5550
rect -2020 5350 -1900 5550
rect -2100 5320 -1900 5350
rect -1600 5320 -1400 5580
rect -1100 5320 -900 5580
rect -600 5320 -500 5580
rect -4000 5300 -3880 5320
rect -3620 5300 -3380 5320
rect -3120 5300 -2880 5320
rect -2620 5300 -2380 5320
rect -2120 5300 -1880 5320
rect -1620 5300 -1380 5320
rect -1120 5300 -880 5320
rect -620 5300 -500 5320
rect -4000 5290 -500 5300
rect -4000 5220 -3850 5290
rect -3650 5220 -3350 5290
rect -3150 5220 -2850 5290
rect -2650 5220 -2350 5290
rect -2150 5220 -500 5290
rect -4000 5200 -500 5220
rect 500 5680 620 5700
rect 880 5680 1120 5700
rect 1380 5680 1620 5700
rect 1880 5680 2120 5700
rect 2380 5680 2620 5700
rect 2880 5680 3120 5700
rect 3380 5680 3620 5700
rect 3880 5680 4000 5700
rect 500 5420 600 5680
rect 900 5420 1100 5680
rect 1400 5420 1600 5680
rect 1900 5420 2100 5680
rect 2400 5420 2600 5680
rect 2900 5420 3100 5680
rect 3400 5420 3600 5680
rect 3900 5420 4000 5680
rect 500 5400 620 5420
rect 880 5400 1120 5420
rect 1380 5400 1620 5420
rect 1880 5400 2120 5420
rect 2380 5400 2620 5420
rect 2880 5400 3120 5420
rect 3380 5400 3620 5420
rect 3880 5400 4000 5420
rect 500 5200 4000 5400
rect -5500 5100 -3500 5200
rect -5500 5080 -5380 5100
rect -5120 5080 -4880 5100
rect -4620 5080 -4380 5100
rect -4120 5080 -3880 5100
rect -3620 5080 -3500 5100
rect -5500 4820 -5400 5080
rect -5100 4820 -4900 5080
rect -4600 4820 -4400 5080
rect -4100 4820 -3900 5080
rect -3600 4820 -3500 5080
rect -5500 4800 -5380 4820
rect -5120 4800 -4880 4820
rect -4620 4800 -4380 4820
rect -4120 4800 -3880 4820
rect -3620 4800 -3500 4820
rect -5500 4600 -3500 4800
rect -5500 4580 -5380 4600
rect -5120 4580 -4880 4600
rect -4620 4580 -4380 4600
rect -4120 4580 -3880 4600
rect -3620 4580 -3500 4600
rect -5500 4320 -5400 4580
rect -5100 4320 -4900 4580
rect -4600 4320 -4400 4580
rect -4100 4320 -3900 4580
rect -3600 4320 -3500 4580
rect -5500 4300 -5380 4320
rect -5120 4300 -4880 4320
rect -4620 4300 -4380 4320
rect -4120 4300 -3880 4320
rect -3620 4300 -3500 4320
rect -5500 4100 -3500 4300
rect -5500 4080 -5380 4100
rect -5120 4080 -4880 4100
rect -4620 4080 -4380 4100
rect -4120 4080 -3880 4100
rect -3620 4080 -3500 4100
rect -5500 3820 -5400 4080
rect -5100 3820 -4900 4080
rect -4600 3820 -4400 4080
rect -4100 3820 -3900 4080
rect -3600 3820 -3500 4080
rect -5500 3800 -5380 3820
rect -5120 3800 -4880 3820
rect -4620 3800 -4380 3820
rect -4120 3800 -3880 3820
rect -3620 3800 -3500 3820
rect 500 5180 620 5200
rect 880 5180 1120 5200
rect 1380 5180 1620 5200
rect 1880 5180 2120 5200
rect 2380 5180 2620 5200
rect 2880 5180 3120 5200
rect 3380 5180 3620 5200
rect 3880 5180 4000 5200
rect 500 4920 600 5180
rect 900 4920 1100 5180
rect 1400 4920 1600 5180
rect 1900 4920 2100 5180
rect 2400 4920 2600 5180
rect 2900 4920 3100 5180
rect 3400 4920 3600 5180
rect 3900 4920 4000 5180
rect 500 4900 620 4920
rect 880 4900 1120 4920
rect 1380 4900 1620 4920
rect 1880 4900 2120 4920
rect 2380 4900 2620 4920
rect 2880 4900 3120 4920
rect 3380 4900 3620 4920
rect 3880 4900 4000 4920
rect 500 4700 4000 4900
rect 500 4680 620 4700
rect 880 4680 1120 4700
rect 1380 4680 1620 4700
rect 1880 4680 2120 4700
rect 2380 4680 2620 4700
rect 2880 4680 3120 4700
rect 3380 4680 3620 4700
rect 3880 4680 4000 4700
rect 500 4420 600 4680
rect 900 4420 1100 4680
rect 1400 4420 1600 4680
rect 1900 4420 2100 4680
rect 2400 4420 2600 4680
rect 2900 4420 3100 4680
rect 3400 4420 3600 4680
rect 3900 4420 4000 4680
rect 500 4400 620 4420
rect 880 4400 1120 4420
rect 1380 4400 1620 4420
rect 1880 4400 2120 4420
rect 2380 4400 2620 4420
rect 2880 4400 3120 4420
rect 3380 4400 3620 4420
rect 3880 4400 4000 4420
rect 500 4200 4000 4400
rect 500 4180 620 4200
rect 880 4180 1120 4200
rect 1380 4180 1620 4200
rect 1880 4180 2120 4200
rect 2380 4180 2620 4200
rect 2880 4180 3120 4200
rect 3380 4180 3620 4200
rect 3880 4180 4000 4200
rect 500 3920 600 4180
rect 900 3920 1100 4180
rect 1400 3920 1600 4180
rect 1900 3920 2100 4180
rect 2400 3920 2600 4180
rect 2900 3920 3100 4180
rect 3400 3920 3600 4180
rect 3900 3920 4000 4180
rect 500 3900 620 3920
rect 880 3900 1120 3920
rect 1380 3900 1620 3920
rect 1880 3900 2120 3920
rect 2380 3900 2620 3920
rect 2880 3900 3120 3920
rect 3380 3900 3620 3920
rect 3880 3900 4000 3920
rect 500 3800 4000 3900
rect -5500 3600 -3500 3800
rect -5500 3580 -5380 3600
rect -5120 3580 -4880 3600
rect -4620 3580 -4380 3600
rect -4120 3580 -3880 3600
rect -3620 3580 -3500 3600
rect -5500 3320 -5400 3580
rect -5100 3320 -4900 3580
rect -4600 3320 -4400 3580
rect -4100 3320 -3900 3580
rect -3600 3320 -3500 3580
rect -5500 3300 -5380 3320
rect -5120 3300 -4880 3320
rect -4620 3300 -4380 3320
rect -4120 3300 -3880 3320
rect -3620 3300 -3500 3320
rect -5500 3100 -3500 3300
rect -5500 3080 -5380 3100
rect -5120 3080 -4880 3100
rect -4620 3080 -4380 3100
rect -4120 3080 -3880 3100
rect -3620 3080 -3500 3100
rect -5500 2820 -5400 3080
rect -5100 2820 -4900 3080
rect -4600 2820 -4400 3080
rect -4100 2820 -3900 3080
rect -3600 2820 -3500 3080
rect -5500 2800 -5380 2820
rect -5120 2800 -4880 2820
rect -4620 2800 -4380 2820
rect -4120 2800 -3880 2820
rect -3620 2800 -3500 2820
rect -500 3700 4000 3800
rect -500 3680 -380 3700
rect -120 3680 120 3700
rect 380 3680 620 3700
rect 880 3680 1120 3700
rect 1380 3680 1620 3700
rect 1880 3680 2120 3700
rect 2380 3680 2620 3700
rect 2880 3680 3120 3700
rect 3380 3680 3620 3700
rect 3880 3680 4000 3700
rect -500 3420 -400 3680
rect -100 3420 100 3680
rect 400 3420 600 3680
rect 900 3420 1100 3680
rect 1400 3420 1600 3680
rect 1900 3420 2100 3680
rect 2400 3420 2600 3680
rect 2900 3420 3100 3680
rect 3400 3420 3600 3680
rect 3900 3420 4000 3680
rect -500 3400 -380 3420
rect -120 3400 120 3420
rect 380 3400 620 3420
rect 880 3400 1120 3420
rect 1380 3400 1620 3420
rect 1880 3400 2120 3420
rect 2380 3400 2620 3420
rect 2880 3400 3120 3420
rect 3380 3400 3620 3420
rect 3880 3400 4000 3420
rect -500 3200 4000 3400
rect -500 3180 -380 3200
rect -120 3180 120 3200
rect 380 3180 620 3200
rect 880 3180 1120 3200
rect 1380 3180 1620 3200
rect 1880 3180 2120 3200
rect 2380 3180 2620 3200
rect 2880 3180 3120 3200
rect 3380 3180 3620 3200
rect 3880 3180 4000 3200
rect -500 2920 -400 3180
rect -100 2920 100 3180
rect 400 2920 600 3180
rect 900 2920 1100 3180
rect 1400 2920 1600 3180
rect 1900 2920 2100 3180
rect 2400 2920 2600 3180
rect 2900 2920 3100 3180
rect 3400 2920 3600 3180
rect 3900 2920 4000 3180
rect -500 2900 -380 2920
rect -120 2900 120 2920
rect 380 2900 620 2920
rect 880 2900 1120 2920
rect 1380 2900 1620 2920
rect 1880 2900 2120 2920
rect 2380 2900 2620 2920
rect 2880 2900 3120 2920
rect 3380 2900 3620 2920
rect 3880 2900 4000 2920
rect -500 2800 4000 2900
rect -5500 2700 4000 2800
rect -5500 2680 -3380 2700
rect -3120 2680 -2880 2700
rect -2620 2680 -2380 2700
rect -2120 2680 -1880 2700
rect -1620 2680 -1380 2700
rect -1120 2680 -880 2700
rect -620 2680 -380 2700
rect -120 2680 120 2700
rect 380 2680 620 2700
rect 880 2680 1120 2700
rect 1380 2680 1620 2700
rect 1880 2680 2120 2700
rect 2380 2680 2620 2700
rect 2880 2680 3120 2700
rect 3380 2680 3620 2700
rect 3880 2680 4000 2700
rect -5500 2600 -3400 2680
rect -5500 2580 -5380 2600
rect -5120 2580 -4880 2600
rect -4620 2580 -4380 2600
rect -4120 2580 -3880 2600
rect -3620 2580 -3400 2600
rect -5500 2320 -5400 2580
rect -5100 2320 -4900 2580
rect -4600 2320 -4400 2580
rect -4100 2320 -3900 2580
rect -3600 2420 -3400 2580
rect -3100 2420 -2900 2680
rect -2600 2420 -2400 2680
rect -2100 2420 -1900 2680
rect -1600 2420 -1400 2680
rect -1100 2420 -900 2680
rect -600 2420 -400 2680
rect -100 2420 100 2680
rect 400 2420 600 2680
rect 900 2420 1100 2680
rect 1400 2420 1600 2680
rect 1900 2420 2100 2680
rect 2400 2420 2600 2680
rect 2900 2420 3100 2680
rect 3400 2420 3600 2680
rect 3900 2420 4000 2680
rect -3600 2400 -3380 2420
rect -3120 2400 -2880 2420
rect -2620 2400 -2380 2420
rect -2120 2400 -1880 2420
rect -1620 2400 -1380 2420
rect -1120 2400 -880 2420
rect -620 2400 -380 2420
rect -120 2400 120 2420
rect 380 2400 620 2420
rect 880 2400 1120 2420
rect 1380 2400 1620 2420
rect 1880 2400 2120 2420
rect 2380 2400 2620 2420
rect 2880 2400 3120 2420
rect 3380 2400 3620 2420
rect 3880 2400 4000 2420
rect -3600 2320 4000 2400
rect -5500 2300 -5380 2320
rect -5120 2300 -4880 2320
rect -4620 2300 -4380 2320
rect -4120 2300 -3880 2320
rect -3620 2300 4000 2320
rect -5500 2200 4000 2300
rect -5500 2180 -3380 2200
rect -3120 2180 -2880 2200
rect -2620 2180 -2380 2200
rect -2120 2180 -1880 2200
rect -1620 2180 -1380 2200
rect -1120 2180 -880 2200
rect -620 2180 -380 2200
rect -120 2180 120 2200
rect 380 2180 620 2200
rect 880 2180 1120 2200
rect 1380 2180 1620 2200
rect 1880 2180 2120 2200
rect 2380 2180 2620 2200
rect 2880 2180 3120 2200
rect 3380 2180 3620 2200
rect 3880 2180 4000 2200
rect -5500 2100 -3400 2180
rect -5500 2080 -5380 2100
rect -5120 2080 -4880 2100
rect -4620 2080 -4380 2100
rect -4120 2080 -3880 2100
rect -3620 2080 -3400 2100
rect -5500 1820 -5400 2080
rect -5100 1820 -4900 2080
rect -4600 1820 -4400 2080
rect -4100 1820 -3900 2080
rect -3600 1920 -3400 2080
rect -3100 1920 -2900 2180
rect -2600 1920 -2400 2180
rect -2100 1920 -1900 2180
rect -1600 1920 -1400 2180
rect -1100 1920 -900 2180
rect -600 1920 -400 2180
rect -100 1920 100 2180
rect 400 1920 600 2180
rect 900 1920 1100 2180
rect 1400 1920 1600 2180
rect 1900 1920 2100 2180
rect 2400 1920 2600 2180
rect 2900 1920 3100 2180
rect 3400 1920 3600 2180
rect 3900 1920 4000 2180
rect -3600 1900 -3380 1920
rect -3120 1900 -2880 1920
rect -2620 1900 -2380 1920
rect -2120 1900 -1880 1920
rect -1620 1900 -1380 1920
rect -1120 1900 -880 1920
rect -620 1900 -380 1920
rect -120 1900 120 1920
rect 380 1900 620 1920
rect 880 1900 1120 1920
rect 1380 1900 1620 1920
rect 1880 1900 2120 1920
rect 2380 1900 2620 1920
rect 2880 1900 3120 1920
rect 3380 1900 3620 1920
rect 3880 1900 4000 1920
rect -3600 1820 4000 1900
rect -5500 1800 -5380 1820
rect -5120 1800 -4880 1820
rect -4620 1800 -4380 1820
rect -4120 1800 -3880 1820
rect -3620 1800 4000 1820
rect -5500 1600 -3500 1800
rect -5500 1580 -5380 1600
rect -5120 1580 -4880 1600
rect -4620 1580 -4380 1600
rect -4120 1580 -3880 1600
rect -3620 1580 -3500 1600
rect -5500 1320 -5400 1580
rect -5100 1320 -4900 1580
rect -4600 1320 -4400 1580
rect -4100 1320 -3900 1580
rect -3600 1320 -3500 1580
rect -5500 1300 -5380 1320
rect -5120 1300 -4880 1320
rect -4620 1300 -4380 1320
rect -4120 1300 -3880 1320
rect -3620 1300 -3500 1320
rect -5500 1100 -3500 1300
rect -5500 1080 -5380 1100
rect -5120 1080 -4880 1100
rect -4620 1080 -4380 1100
rect -4120 1080 -3880 1100
rect -3620 1080 -3500 1100
rect -5500 820 -5400 1080
rect -5100 820 -4900 1080
rect -4600 820 -4400 1080
rect -4100 820 -3900 1080
rect -3600 820 -3500 1080
rect -5500 800 -5380 820
rect -5120 800 -4880 820
rect -4620 800 -4380 820
rect -4120 800 -3880 820
rect -3620 800 -3500 820
rect -5500 600 -3500 800
rect -5500 580 -5380 600
rect -5120 580 -4880 600
rect -4620 580 -4380 600
rect -4120 580 -3880 600
rect -3620 580 -3500 600
rect -5500 320 -5400 580
rect -5100 320 -4900 580
rect -4600 320 -4400 580
rect -4100 320 -3900 580
rect -3600 320 -3500 580
rect -5500 300 -5380 320
rect -5120 300 -4880 320
rect -4620 300 -4380 320
rect -4120 300 -3880 320
rect -3620 300 -3500 320
rect -700 1700 4000 1800
rect -700 1680 -580 1700
rect -320 1680 -200 1700
rect -700 1420 -600 1680
rect -300 1420 -200 1680
rect -700 1400 -580 1420
rect -320 1400 -200 1420
rect -700 1200 -200 1400
rect -700 1180 -580 1200
rect -320 1180 -200 1200
rect -700 920 -600 1180
rect -300 920 -200 1180
rect -700 900 -580 920
rect -320 900 -200 920
rect -700 700 -200 900
rect -700 680 -580 700
rect -320 680 -200 700
rect -700 420 -600 680
rect -300 420 -200 680
rect -700 400 -580 420
rect -320 400 -200 420
rect -700 300 -200 400
rect 1200 1680 1420 1700
rect 1680 1680 1900 1700
rect 1200 1420 1400 1680
rect 1700 1420 1900 1680
rect 1200 1400 1420 1420
rect 1680 1400 1900 1420
rect 1200 1200 1900 1400
rect 1200 1180 1420 1200
rect 1680 1180 1900 1200
rect 1200 920 1400 1180
rect 1700 920 1900 1180
rect 1200 900 1420 920
rect 1680 900 1900 920
rect 1200 700 1900 900
rect 1200 680 1420 700
rect 1680 680 1900 700
rect 1200 420 1400 680
rect 1700 420 1900 680
rect 1200 400 1420 420
rect 1680 400 1900 420
rect 1200 300 1900 400
rect -5500 100 -3500 300
rect -1000 200 50 300
rect -5500 80 -5380 100
rect -5120 80 -4880 100
rect -4620 80 -4380 100
rect -4120 80 -3880 100
rect -3620 80 -3500 100
rect -5500 -180 -5400 80
rect -5100 -180 -4900 80
rect -4600 -180 -4400 80
rect -4100 -180 -3900 80
rect -3600 -180 -3500 80
rect -5500 -200 -5380 -180
rect -5120 -200 -4880 -180
rect -4620 -200 -4380 -180
rect -4120 -200 -3880 -180
rect -3620 -200 -3500 -180
rect -5500 -300 -3500 -200
rect -1500 100 50 200
rect -1500 80 -1380 100
rect -1120 80 50 100
rect -1500 -180 -1400 80
rect -1100 -180 50 80
rect -1500 -200 -1380 -180
rect -1120 -200 50 -180
rect -5500 -400 -4500 -300
rect -5500 -420 -5380 -400
rect -5120 -420 -4880 -400
rect -4620 -420 -4500 -400
rect -5500 -680 -5400 -420
rect -5100 -680 -4900 -420
rect -4600 -600 -4500 -420
rect -1500 -400 50 -200
rect -1500 -420 -1380 -400
rect -1120 -420 50 -400
rect -4600 -640 -4400 -600
rect -4600 -680 -4540 -640
rect -5500 -700 -5380 -680
rect -5120 -700 -4880 -680
rect -4620 -700 -4540 -680
rect -5500 -900 -4540 -700
rect -5500 -920 -5380 -900
rect -5120 -920 -4880 -900
rect -4620 -920 -4540 -900
rect -5500 -1180 -5400 -920
rect -5100 -1180 -4900 -920
rect -4600 -1180 -4540 -920
rect -5500 -1200 -5380 -1180
rect -5120 -1200 -4880 -1180
rect -4620 -1200 -4540 -1180
rect -14500 -1400 -10000 -1300
rect -14500 -1420 -14380 -1400
rect -14120 -1420 -13880 -1400
rect -13620 -1420 -13380 -1400
rect -13120 -1420 -12880 -1400
rect -12620 -1420 -12380 -1400
rect -12120 -1420 -11880 -1400
rect -11620 -1420 -11380 -1400
rect -11120 -1420 -10880 -1400
rect -10620 -1420 -10380 -1400
rect -10120 -1420 -10000 -1400
rect -14500 -1680 -14400 -1420
rect -14100 -1680 -13900 -1420
rect -13600 -1680 -13400 -1420
rect -13100 -1680 -12900 -1420
rect -12600 -1680 -12400 -1420
rect -12100 -1680 -11900 -1420
rect -11600 -1680 -11400 -1420
rect -11100 -1680 -10900 -1420
rect -10600 -1680 -10400 -1420
rect -10100 -1680 -10000 -1420
rect -14500 -1700 -14380 -1680
rect -14120 -1700 -13880 -1680
rect -13620 -1700 -13380 -1680
rect -13120 -1700 -12880 -1680
rect -12620 -1700 -12380 -1680
rect -12120 -1700 -11880 -1680
rect -11620 -1700 -11380 -1680
rect -11120 -1700 -10880 -1680
rect -10620 -1700 -10380 -1680
rect -10120 -1700 -10000 -1680
rect -14500 -1900 -11600 -1700
rect -11400 -1900 -10000 -1700
rect -14500 -1920 -14380 -1900
rect -14120 -1920 -13880 -1900
rect -13620 -1920 -13380 -1900
rect -13120 -1920 -12880 -1900
rect -12620 -1920 -12380 -1900
rect -12120 -1920 -11880 -1900
rect -11620 -1920 -11380 -1900
rect -11120 -1920 -10880 -1900
rect -10620 -1920 -10380 -1900
rect -10120 -1920 -10000 -1900
rect -14500 -2180 -14400 -1920
rect -14100 -2180 -13900 -1920
rect -13600 -2180 -13400 -1920
rect -13100 -2180 -12900 -1920
rect -12600 -2180 -12400 -1920
rect -12100 -2180 -11900 -1920
rect -11600 -2180 -11400 -1920
rect -11100 -2180 -10900 -1920
rect -10600 -2180 -10400 -1920
rect -10100 -2180 -10000 -1920
rect -14500 -2200 -14380 -2180
rect -14120 -2200 -13880 -2180
rect -13620 -2200 -13380 -2180
rect -13120 -2200 -12880 -2180
rect -12620 -2200 -12380 -2180
rect -12120 -2200 -11880 -2180
rect -11620 -2200 -11380 -2180
rect -11120 -2200 -10880 -2180
rect -10620 -2200 -10380 -2180
rect -10120 -2200 -10000 -2180
rect -14500 -2400 -11600 -2200
rect -11400 -2300 -10000 -2200
rect -5500 -1400 -4540 -1200
rect -5500 -1420 -5380 -1400
rect -5120 -1420 -4880 -1400
rect -4620 -1420 -4540 -1400
rect -5500 -1680 -5400 -1420
rect -5100 -1680 -4900 -1420
rect -4600 -1680 -4540 -1420
rect -5500 -1700 -5380 -1680
rect -5120 -1700 -4880 -1680
rect -4620 -1700 -4540 -1680
rect -5500 -1900 -4540 -1700
rect -5500 -1920 -5380 -1900
rect -5120 -1920 -4880 -1900
rect -4620 -1920 -4540 -1900
rect -5500 -2180 -5400 -1920
rect -5100 -2180 -4900 -1920
rect -4600 -2180 -4540 -1920
rect -4420 -2000 -4400 -640
rect -4320 -690 -4120 -670
rect -4320 -890 -4300 -690
rect -4140 -890 -4120 -690
rect -4320 -910 -4120 -890
rect -3980 -690 -3780 -670
rect -3980 -890 -3960 -690
rect -3800 -890 -3780 -690
rect -3980 -910 -3780 -890
rect -1500 -680 -1400 -420
rect -1100 -680 50 -420
rect -1500 -700 -1380 -680
rect -1120 -700 50 -680
rect 950 200 2140 300
rect 950 180 1420 200
rect 1680 180 2140 200
rect 950 -80 1400 180
rect 1700 -80 2140 180
rect 950 -100 1420 -80
rect 1680 -100 2140 -80
rect 950 -300 2140 -100
rect 950 -320 1420 -300
rect 1680 -320 2140 -300
rect 950 -580 1400 -320
rect 1700 -580 2140 -320
rect 950 -600 1420 -580
rect 1680 -600 2140 -580
rect 950 -700 2140 -600
rect -1500 -800 -700 -700
rect -1500 -900 -1000 -800
rect -1500 -920 -1380 -900
rect -1120 -920 -1000 -900
rect -1500 -1180 -1400 -920
rect -1100 -1180 -1000 -920
rect 200 -1100 300 -900
rect 400 -1100 500 -900
rect 600 -1100 700 -900
rect 800 -1100 900 -900
rect 2300 -1100 2400 -900
rect 2500 -1100 2600 -900
rect 2700 -1100 2800 -900
rect 2900 -1100 3000 -900
rect -1500 -1200 -1380 -1180
rect -1120 -1200 -1000 -1180
rect -1500 -1400 -1000 -1200
rect -1500 -1420 -1380 -1400
rect -1120 -1420 -1000 -1400
rect -1500 -1680 -1400 -1420
rect -1100 -1680 -1000 -1420
rect -1500 -1700 -1380 -1680
rect -1120 -1700 -1000 -1680
rect -1500 -1900 -1000 -1700
rect -200 -1200 1000 -1100
rect -200 -1700 -100 -1200
rect 900 -1700 1000 -1200
rect -200 -1800 1000 -1700
rect 2200 -1200 3400 -1100
rect 2200 -1700 2300 -1200
rect 3300 -1700 3400 -1200
rect 2200 -1800 3400 -1700
rect -1500 -1920 -1380 -1900
rect -1120 -1920 -1000 -1900
rect -4420 -2060 -3600 -2000
rect -5500 -2200 -5380 -2180
rect -5120 -2200 -4880 -2180
rect -4620 -2200 -4540 -2180
rect -5500 -2220 -4540 -2200
rect -3740 -2220 -3600 -2060
rect -5500 -2300 -3600 -2220
rect -1500 -2180 -1400 -1920
rect -1100 -2180 -1000 -1920
rect -1500 -2200 -1380 -2180
rect -1120 -2200 -1000 -2180
rect -1500 -2300 -1000 -2200
rect -11400 -2400 -1000 -2300
rect -14500 -2420 -14380 -2400
rect -14120 -2420 -13880 -2400
rect -13620 -2420 -13380 -2400
rect -13120 -2420 -12880 -2400
rect -12620 -2420 -12380 -2400
rect -12120 -2420 -11880 -2400
rect -11620 -2420 -11380 -2400
rect -11120 -2420 -10880 -2400
rect -10620 -2420 -10380 -2400
rect -10120 -2420 -9880 -2400
rect -9620 -2420 -9380 -2400
rect -9120 -2420 -8880 -2400
rect -8620 -2420 -8380 -2400
rect -8120 -2420 -7880 -2400
rect -7620 -2420 -7380 -2400
rect -7120 -2420 -6880 -2400
rect -6620 -2420 -6380 -2400
rect -6120 -2420 -5880 -2400
rect -5620 -2420 -5380 -2400
rect -5120 -2420 -4880 -2400
rect -4620 -2420 -4380 -2400
rect -4120 -2420 -3880 -2400
rect -3620 -2420 -3380 -2400
rect -3120 -2420 -2880 -2400
rect -2620 -2420 -2380 -2400
rect -2120 -2420 -1880 -2400
rect -1620 -2420 -1380 -2400
rect -1120 -2420 -1000 -2400
rect -14500 -2680 -14400 -2420
rect -14100 -2680 -13900 -2420
rect -13600 -2680 -13400 -2420
rect -13100 -2680 -12900 -2420
rect -12600 -2680 -12400 -2420
rect -12100 -2680 -11900 -2420
rect -11600 -2680 -11400 -2420
rect -11100 -2680 -10900 -2420
rect -10600 -2680 -10400 -2420
rect -10100 -2680 -9900 -2420
rect -9600 -2680 -9400 -2420
rect -9100 -2680 -8900 -2420
rect -8600 -2680 -8400 -2420
rect -8100 -2680 -7900 -2420
rect -7600 -2680 -7400 -2420
rect -7100 -2680 -6900 -2420
rect -6600 -2680 -6400 -2420
rect -6100 -2680 -5900 -2420
rect -5600 -2680 -5400 -2420
rect -5100 -2680 -4900 -2420
rect -4600 -2680 -4400 -2420
rect -4100 -2680 -3900 -2420
rect -3600 -2680 -3400 -2420
rect -3100 -2680 -2900 -2420
rect -2600 -2680 -2400 -2420
rect -2100 -2680 -1900 -2420
rect -1600 -2680 -1400 -2420
rect -1100 -2680 -1000 -2420
rect -14500 -2700 -14380 -2680
rect -14120 -2700 -13880 -2680
rect -13620 -2700 -13380 -2680
rect -13120 -2700 -12880 -2680
rect -12620 -2700 -12380 -2680
rect -12120 -2700 -11880 -2680
rect -11620 -2700 -11380 -2680
rect -11120 -2700 -10880 -2680
rect -10620 -2700 -10380 -2680
rect -10120 -2700 -9880 -2680
rect -9620 -2700 -9380 -2680
rect -9120 -2700 -8880 -2680
rect -8620 -2700 -8380 -2680
rect -8120 -2700 -7880 -2680
rect -7620 -2700 -7380 -2680
rect -7120 -2700 -6880 -2680
rect -6620 -2700 -6380 -2680
rect -6120 -2700 -5880 -2680
rect -5620 -2700 -5380 -2680
rect -5120 -2700 -4880 -2680
rect -4620 -2700 -4380 -2680
rect -4120 -2700 -3880 -2680
rect -3620 -2700 -3380 -2680
rect -3120 -2700 -2880 -2680
rect -2620 -2700 -2380 -2680
rect -2120 -2700 -1880 -2680
rect -1620 -2700 -1380 -2680
rect -1120 -2700 -1000 -2680
rect -14500 -2900 -11600 -2700
rect -11400 -2900 -1000 -2700
rect -14500 -2920 -14380 -2900
rect -14120 -2920 -13880 -2900
rect -13620 -2920 -13380 -2900
rect -13120 -2920 -12880 -2900
rect -12620 -2920 -12380 -2900
rect -12120 -2920 -11880 -2900
rect -11620 -2920 -11380 -2900
rect -11120 -2920 -10880 -2900
rect -10620 -2920 -10380 -2900
rect -10120 -2920 -9880 -2900
rect -9620 -2920 -9380 -2900
rect -9120 -2920 -8880 -2900
rect -8620 -2920 -8380 -2900
rect -8120 -2920 -7880 -2900
rect -7620 -2920 -7380 -2900
rect -7120 -2920 -6880 -2900
rect -6620 -2920 -6380 -2900
rect -6120 -2920 -5880 -2900
rect -5620 -2920 -5380 -2900
rect -5120 -2920 -4880 -2900
rect -4620 -2920 -4380 -2900
rect -4120 -2920 -3880 -2900
rect -3620 -2920 -3380 -2900
rect -3120 -2920 -2880 -2900
rect -2620 -2920 -2380 -2900
rect -2120 -2920 -1880 -2900
rect -1620 -2920 -1380 -2900
rect -1120 -2920 -1000 -2900
rect -14500 -3180 -14400 -2920
rect -14100 -3180 -13900 -2920
rect -13600 -3180 -13400 -2920
rect -13100 -3180 -12900 -2920
rect -12600 -3180 -12400 -2920
rect -12100 -3180 -11900 -2920
rect -11600 -3180 -11400 -2920
rect -11100 -3180 -10900 -2920
rect -10600 -3180 -10400 -2920
rect -10100 -3180 -9900 -2920
rect -9600 -3180 -9400 -2920
rect -9100 -3180 -8900 -2920
rect -8600 -3180 -8400 -2920
rect -8100 -3180 -7900 -2920
rect -7600 -3180 -7400 -2920
rect -7100 -3180 -6900 -2920
rect -6600 -3180 -6400 -2920
rect -6100 -3180 -5900 -2920
rect -5600 -3180 -5400 -2920
rect -5100 -3180 -4900 -2920
rect -4600 -3180 -4400 -2920
rect -4100 -3180 -3900 -2920
rect -3600 -3180 -3400 -2920
rect -3100 -3180 -2900 -2920
rect -2600 -3180 -2400 -2920
rect -2100 -3180 -1900 -2920
rect -1600 -3180 -1400 -2920
rect -1100 -3180 -1000 -2920
rect -14500 -3200 -14380 -3180
rect -14120 -3200 -13880 -3180
rect -13620 -3200 -13380 -3180
rect -13120 -3200 -12880 -3180
rect -12620 -3200 -12380 -3180
rect -12120 -3200 -11880 -3180
rect -11620 -3200 -11380 -3180
rect -11120 -3200 -10880 -3180
rect -10620 -3200 -10380 -3180
rect -10120 -3200 -9880 -3180
rect -9620 -3200 -9380 -3180
rect -9120 -3200 -8880 -3180
rect -8620 -3200 -8380 -3180
rect -8120 -3200 -7880 -3180
rect -7620 -3200 -7380 -3180
rect -7120 -3200 -6880 -3180
rect -6620 -3200 -6380 -3180
rect -6120 -3200 -5880 -3180
rect -5620 -3200 -5380 -3180
rect -5120 -3200 -4880 -3180
rect -4620 -3200 -4380 -3180
rect -4120 -3200 -3880 -3180
rect -3620 -3200 -3380 -3180
rect -3120 -3200 -2880 -3180
rect -2620 -3200 -2380 -3180
rect -2120 -3200 -1880 -3180
rect -1620 -3200 -1380 -3180
rect -1120 -3200 -1000 -3180
rect -14500 -3300 -1000 -3200
<< via1 >>
rect -3480 8820 -3320 8980
rect -2360 8660 -2260 8820
rect -1780 8620 -1620 8780
rect -4700 7800 -4500 8600
rect -2350 7110 -2150 7180
rect -1850 7110 -1650 7180
rect -2480 6850 -2410 7050
rect -2090 6850 -2020 7050
rect -1980 6850 -1910 7050
rect -1590 6850 -1520 7050
rect -2350 6720 -2150 6790
rect -1850 6720 -1650 6790
rect -2350 6610 -2150 6680
rect -1850 6610 -1650 6680
rect -2480 6350 -2410 6550
rect -2090 6350 -2020 6550
rect -1980 6350 -1910 6550
rect -1590 6350 -1520 6550
rect -2350 6220 -2150 6290
rect -1850 6220 -1650 6290
rect -3850 6110 -3650 6180
rect -3350 6110 -3150 6180
rect -2850 6110 -2650 6180
rect -2350 6110 -2150 6180
rect -1850 6110 -1650 6180
rect -3980 5850 -3910 6050
rect -3590 5850 -3520 6050
rect -3480 5850 -3410 6050
rect -3090 5850 -3020 6050
rect -2980 5850 -2910 6050
rect -2590 5850 -2520 6050
rect -2480 5850 -2410 6050
rect -2090 5850 -2020 6050
rect -1980 5850 -1910 6050
rect -1590 5850 -1520 6050
rect -3850 5720 -3650 5790
rect -3350 5720 -3150 5790
rect -2850 5720 -2650 5790
rect -2350 5720 -2150 5790
rect -1850 5720 -1650 5790
rect -980 7000 -820 7020
rect -980 6880 -960 7000
rect -960 6880 -840 7000
rect -840 6880 -820 7000
rect -980 6860 -820 6880
rect -1180 5900 -1020 5920
rect -1180 5780 -1160 5900
rect -1160 5780 -1040 5900
rect -1040 5780 -1020 5900
rect -1180 5760 -1020 5780
rect -3850 5610 -3650 5680
rect -3350 5610 -3150 5680
rect -2850 5610 -2650 5680
rect -2350 5610 -2150 5680
rect -3980 5350 -3910 5550
rect -3590 5350 -3520 5550
rect -3480 5350 -3410 5550
rect -3090 5350 -3020 5550
rect -2980 5350 -2910 5550
rect -2590 5350 -2520 5550
rect -2480 5350 -2410 5550
rect -2090 5350 -2020 5550
rect -3850 5220 -3650 5290
rect -3350 5220 -3150 5290
rect -2850 5220 -2650 5290
rect -2350 5220 -2150 5290
rect -11600 -1900 -11400 -1700
rect -11600 -2400 -11400 -2200
rect -4300 -720 -4140 -690
rect -4300 -860 -4260 -720
rect -4260 -860 -4140 -720
rect -4300 -890 -4140 -860
rect -3960 -720 -3800 -690
rect -3960 -860 -3940 -720
rect -3940 -860 -3820 -720
rect -3820 -860 -3800 -720
rect -3960 -890 -3800 -860
rect -100 -1700 900 -1200
rect 2300 -1700 3300 -1200
rect -11600 -2900 -11400 -2700
<< metal2 >>
rect -6700 17200 -6600 18600
rect -6300 17200 -6200 18600
rect -5900 17200 -5800 18600
rect -5500 17200 -5400 18600
rect -4800 17100 -3300 17200
rect -5000 16600 -4700 17100
rect -3400 16600 -3300 17100
rect -4800 16500 -3300 16600
rect -6700 14800 -5300 15000
rect -6800 12600 -5200 14800
rect -4300 14180 -3760 14200
rect -4300 13620 -4280 14180
rect -3820 13620 -3760 14180
rect -4300 13600 -3760 13620
rect -15200 12400 -4400 12600
rect -15200 11600 -15000 12400
rect -4600 11600 -4400 12400
rect -15200 11400 -4400 11600
rect -15000 8000 -13200 11400
rect -12800 8000 -11800 11400
rect -11400 8000 -10600 11400
rect -10200 8000 -9400 11400
rect -9000 8000 -8200 11400
rect -7800 8000 -7000 11400
rect -6600 8000 -5800 11400
rect -5400 8600 -4400 11400
rect -3960 9000 -3760 13600
rect -800 12500 1000 12600
rect -800 9100 -700 12500
rect 900 10000 1000 12500
rect 900 9900 3100 10000
rect 3000 9100 3100 9900
rect -800 9000 3100 9100
rect -3960 8980 -3300 9000
rect -3960 8820 -3480 8980
rect -3320 8820 -3300 8980
rect -50 8930 1020 9000
rect 1960 8930 3100 9000
rect -50 8860 3100 8930
rect -3960 8800 -3300 8820
rect -2380 8820 -2080 8840
rect -2380 8620 -2360 8820
rect -2100 8620 -2080 8820
rect -2380 8600 -2080 8620
rect -1800 8780 -1600 8800
rect -1800 8620 -1780 8780
rect -1620 8620 -1600 8780
rect -1800 8600 -1600 8620
rect -5400 8000 -4700 8600
rect -15000 7800 -4700 8000
rect -4500 8000 -4400 8600
rect -50 8500 1020 8860
rect 1960 8500 3100 8860
rect -4500 7800 -4200 8000
rect -15000 3200 -14800 7800
rect -4400 6200 -4200 7800
rect 0 7210 1000 7400
rect 2000 7210 3000 7400
rect 0 7200 3000 7210
rect -2360 7180 -2140 7200
rect -2360 7110 -2350 7180
rect -2150 7110 -2140 7180
rect -2360 7060 -2140 7110
rect -1860 7180 -1640 7200
rect -1860 7110 -1850 7180
rect -1650 7110 -1640 7180
rect -1860 7060 -1640 7110
rect -2500 7050 -1500 7060
rect -2500 6850 -2480 7050
rect -2410 6850 -2090 7050
rect -2020 6850 -1980 7050
rect -1910 6850 -1590 7050
rect -1520 6850 -1500 7050
rect -2500 6840 -1500 6850
rect -1160 7020 -800 7040
rect -1160 6860 -1140 7020
rect -820 6860 -800 7020
rect -1160 6840 -800 6860
rect -2360 6790 -2140 6840
rect -2360 6720 -2350 6790
rect -2150 6720 -2140 6790
rect -2360 6680 -2140 6720
rect -2360 6610 -2350 6680
rect -2150 6610 -2140 6680
rect -2360 6560 -2140 6610
rect -1860 6790 -1640 6840
rect -1860 6720 -1850 6790
rect -1650 6720 -1640 6790
rect -1860 6680 -1640 6720
rect -1860 6610 -1850 6680
rect -1650 6610 -1640 6680
rect -1860 6560 -1640 6610
rect -2500 6550 -1500 6560
rect -2500 6350 -2480 6550
rect -2410 6350 -2090 6550
rect -2020 6350 -1980 6550
rect -1910 6350 -1590 6550
rect -1520 6350 -1500 6550
rect -2500 6340 -1500 6350
rect 0 6400 100 7200
rect 900 7170 2100 7200
rect 900 6400 1000 7170
rect -2360 6290 -2140 6340
rect -2360 6220 -2350 6290
rect -2150 6220 -2140 6290
rect -4400 6060 -4000 6200
rect -3860 6180 -3640 6200
rect -3860 6110 -3850 6180
rect -3650 6110 -3640 6180
rect -3860 6060 -3640 6110
rect -3360 6180 -3140 6200
rect -3360 6110 -3350 6180
rect -3150 6110 -3140 6180
rect -3360 6060 -3140 6110
rect -2860 6180 -2640 6200
rect -2860 6110 -2850 6180
rect -2650 6110 -2640 6180
rect -2860 6060 -2640 6110
rect -2360 6180 -2140 6220
rect -2360 6110 -2350 6180
rect -2150 6110 -2140 6180
rect -2360 6060 -2140 6110
rect -1860 6290 -1640 6340
rect 0 6300 1000 6400
rect 2000 6400 2100 7170
rect 2900 6400 3000 7200
rect 2000 6300 3000 6400
rect -1860 6220 -1850 6290
rect -1650 6220 -1640 6290
rect -1860 6180 -1640 6220
rect -1860 6110 -1850 6180
rect -1650 6110 -1640 6180
rect -1860 6060 -1640 6110
rect -4400 6050 -1500 6060
rect -4400 5850 -3980 6050
rect -3910 5850 -3590 6050
rect -3520 5850 -3480 6050
rect -3410 5850 -3090 6050
rect -3020 5850 -2980 6050
rect -2910 5850 -2590 6050
rect -2520 5850 -2480 6050
rect -2410 5850 -2090 6050
rect -2020 5850 -1980 6050
rect -1910 5850 -1590 6050
rect -1520 5850 -1500 6050
rect -4400 5840 -1500 5850
rect -1200 5920 -840 5940
rect -4400 5600 -4000 5840
rect -3860 5790 -3640 5840
rect -3860 5720 -3850 5790
rect -3650 5720 -3640 5790
rect -3860 5680 -3640 5720
rect -3860 5610 -3850 5680
rect -3650 5610 -3640 5680
rect -3860 5600 -3640 5610
rect -4400 5560 -3640 5600
rect -3360 5790 -3140 5840
rect -3360 5720 -3350 5790
rect -3150 5720 -3140 5790
rect -3360 5680 -3140 5720
rect -3360 5610 -3350 5680
rect -3150 5610 -3140 5680
rect -3360 5560 -3140 5610
rect -2860 5790 -2640 5840
rect -2860 5720 -2850 5790
rect -2650 5720 -2640 5790
rect -2860 5680 -2640 5720
rect -2860 5610 -2850 5680
rect -2650 5610 -2640 5680
rect -2860 5560 -2640 5610
rect -2360 5790 -2140 5840
rect -2360 5720 -2350 5790
rect -2150 5720 -2140 5790
rect -2360 5680 -2140 5720
rect -1860 5790 -1640 5840
rect -1860 5720 -1850 5790
rect -1650 5720 -1640 5790
rect -1200 5760 -1180 5920
rect -860 5760 -840 5920
rect -1200 5740 -840 5760
rect -1860 5700 -1640 5720
rect -2360 5610 -2350 5680
rect -2150 5610 -2140 5680
rect -2360 5560 -2140 5610
rect -4400 5550 -2000 5560
rect -4400 5400 -3980 5550
rect -4000 5350 -3980 5400
rect -3910 5350 -3590 5550
rect -3520 5350 -3480 5550
rect -3410 5350 -3090 5550
rect -3020 5350 -2980 5550
rect -2910 5350 -2590 5550
rect -2520 5350 -2480 5550
rect -2410 5350 -2090 5550
rect -2020 5350 -2000 5550
rect -4000 5340 -2000 5350
rect -4000 5290 -3640 5340
rect -4000 5220 -3850 5290
rect -3650 5220 -3640 5290
rect -4000 5200 -3640 5220
rect -3360 5290 -3140 5340
rect -3360 5220 -3350 5290
rect -3150 5220 -3140 5290
rect -3360 5200 -3140 5220
rect -2860 5290 -2640 5340
rect -2860 5220 -2850 5290
rect -2650 5220 -2640 5290
rect -2860 5200 -2640 5220
rect -2360 5290 -2140 5340
rect -2360 5220 -2350 5290
rect -2150 5220 -2140 5290
rect -2360 5200 -2140 5220
rect -4000 3200 -3800 5200
rect -15000 3000 -3800 3200
rect 0 1200 1000 1300
rect 0 500 100 1200
rect 900 500 1000 1200
rect 0 400 1000 500
rect 2100 1200 3100 1300
rect 2100 500 2200 1200
rect 3000 500 3100 1200
rect 2100 380 3100 500
rect -4320 -680 -4120 -660
rect -4320 -900 -4300 -680
rect -4140 -900 -4120 -680
rect -4320 -920 -4120 -900
rect -3980 -690 -3780 -670
rect -3980 -890 -3960 -690
rect -3800 -890 -3780 -690
rect -3980 -910 -3780 -890
rect -800 -1000 4200 -700
rect -12000 -1400 -11000 -1300
rect -12000 -3200 -11900 -1400
rect -11100 -3200 -11000 -1400
rect -12000 -3300 -11000 -3200
rect -800 -2100 -400 -1000
rect -200 -1200 1000 -1100
rect -200 -1700 -100 -1200
rect 900 -1700 1000 -1200
rect -200 -1800 1000 -1700
rect 1300 -2100 1900 -1000
rect 2200 -1200 3400 -1100
rect 2200 -1700 2300 -1200
rect 3300 -1700 3400 -1200
rect 2200 -1800 3400 -1700
rect 3800 -2100 4200 -1000
rect -800 -2300 4200 -2100
rect -800 -4700 -700 -2300
rect 1200 -2600 4200 -2300
rect 1200 -4700 1300 -2600
rect -800 -4800 1300 -4700
<< via2 >>
rect -4700 16600 -3400 17100
rect -4280 13620 -3820 14180
rect -15000 11600 -4600 12400
rect -700 9900 900 12500
rect -700 9100 3000 9900
rect -2360 8660 -2260 8820
rect -2260 8660 -2100 8820
rect -2360 8620 -2100 8660
rect -14800 5400 -4400 7800
rect -1140 6860 -980 7020
rect -980 6860 -820 7020
rect 100 6400 900 7200
rect 2100 6400 2900 7200
rect -1180 5760 -1020 5920
rect -1020 5760 -860 5920
rect -14800 3200 -4000 5400
rect 100 500 900 1200
rect 2200 500 3000 1200
rect -4300 -690 -4140 -680
rect -4300 -890 -4140 -690
rect -4300 -900 -4140 -890
rect -3960 -890 -3800 -690
rect -11900 -1700 -11100 -1400
rect -11900 -1900 -11600 -1700
rect -11600 -1900 -11400 -1700
rect -11400 -1900 -11100 -1700
rect -11900 -2200 -11100 -1900
rect -11900 -2400 -11600 -2200
rect -11600 -2400 -11400 -2200
rect -11400 -2400 -11100 -2200
rect -11900 -2700 -11100 -2400
rect -11900 -2900 -11600 -2700
rect -11600 -2900 -11400 -2700
rect -11400 -2900 -11100 -2700
rect -11900 -3200 -11100 -2900
rect -100 -1700 900 -1200
rect 2300 -1700 3300 -1200
rect -700 -4700 1200 -2300
<< metal3 >>
rect -18000 23700 -10400 23800
rect -18000 22400 -17900 23700
rect -10500 22400 -10400 23700
rect -18000 22000 -10400 22400
rect -20600 20000 -10400 22000
rect -20600 19800 -7600 20000
rect -20600 16600 -9000 19800
rect -7800 17600 -7600 19800
rect -4700 18400 1000 18500
rect -7800 16600 -7200 17600
rect -4700 17200 -4300 18400
rect -20600 16400 -7200 16600
rect -4800 17100 -4300 17200
rect -4800 16600 -4700 17100
rect 900 16600 1000 18400
rect -4800 16500 1000 16600
rect -20600 13000 -10400 16400
rect -8600 14200 -8000 16400
rect -8600 14180 -3800 14200
rect -8600 13620 -4280 14180
rect -3820 13620 -3800 14180
rect -8600 13600 -3800 13620
rect -18000 12400 -4400 12600
rect -18000 11600 -17800 12400
rect -4600 11600 -4400 12400
rect -18000 11400 -4400 11600
rect -1200 12500 1000 12600
rect -1200 9100 -700 12500
rect 900 10000 1000 12500
rect 900 9900 3100 10000
rect 3000 9100 3100 9900
rect -1200 9000 3100 9100
rect -2380 8820 -2080 8840
rect -2380 8620 -2360 8820
rect -2100 8620 -2080 8820
rect -2380 8200 -2080 8620
rect -3600 8150 -2080 8200
rect -15000 7800 -4200 8000
rect -15000 3200 -14800 7800
rect -4400 5600 -4200 7800
rect -3600 7850 -3550 8150
rect -2650 7850 -2080 8150
rect -3600 7820 -2080 7850
rect -3600 6000 -2600 7820
rect -1160 7020 -800 9000
rect 3500 8000 7700 8100
rect 3500 7300 3600 8000
rect -1160 6860 -1140 7020
rect -820 6860 -800 7020
rect -1160 6840 -800 6860
rect 0 7200 3600 7300
rect 0 6400 100 7200
rect 7600 6600 7700 8000
rect 3800 6400 7700 6600
rect 0 6300 7700 6400
rect -1200 5920 200 6000
rect -1200 5760 -1180 5920
rect -860 5900 200 5920
rect -860 5800 -300 5900
rect -860 5760 -840 5800
rect -1200 5740 -840 5760
rect -4400 5400 -3800 5600
rect -4000 3200 -3800 5400
rect -15000 3000 -3800 3200
rect -5600 -50 -3600 2600
rect -3200 600 -800 5200
rect -400 4400 -300 5800
rect 100 4400 200 5900
rect -400 4200 200 4400
rect 3700 1400 6400 1600
rect -3200 100 -3100 600
rect -900 100 -800 600
rect 0 1300 3900 1400
rect 0 500 100 1300
rect 0 400 3900 500
rect 2100 380 3100 400
rect -3200 0 -800 100
rect 3700 200 3900 400
rect 6300 200 6400 1400
rect 3700 0 6400 200
rect -5600 -350 -5550 -50
rect -3650 -350 -3600 -50
rect -5600 -400 -3600 -350
rect -4320 -680 -4120 -400
rect -4320 -900 -4300 -680
rect -4140 -900 -4120 -680
rect -4320 -920 -4120 -900
rect -3980 -680 -3780 -670
rect -3000 -680 -1000 0
rect -3980 -690 -1000 -680
rect -3980 -890 -3960 -690
rect -3800 -700 -1000 -690
rect -3800 -890 -2900 -700
rect -3980 -910 -2900 -890
rect -3660 -920 -2900 -910
rect -12000 -1400 -11000 -1300
rect -12000 -3200 -11900 -1400
rect -11100 -3200 -11000 -1400
rect -3000 -1700 -2900 -920
rect -1100 -1100 -1000 -700
rect -1100 -1200 3400 -1100
rect -3000 -1800 2300 -1700
rect -12000 -3300 -11000 -3200
rect -800 -2300 1300 -2200
rect -800 -4700 -700 -2300
rect 1200 -4700 1300 -2300
rect 2200 -3200 2300 -1800
rect 3300 -3200 3400 -1200
rect 2200 -3400 3400 -3200
rect -800 -4800 1300 -4700
<< via3 >>
rect -17900 22400 -10500 23700
rect -9000 16600 -7800 19800
rect -4300 17100 900 18400
rect -4300 16600 -3400 17100
rect -3400 16600 900 17100
rect -17800 11600 -15000 12400
rect -15000 11600 -4600 12400
rect -700 9900 900 12500
rect -700 9100 3000 9900
rect -14800 5400 -4400 7800
rect -3550 7850 -2650 8150
rect 3600 7200 7600 8000
rect 100 6400 900 7200
rect 900 6400 2100 7200
rect 2100 6400 2900 7200
rect 2900 6600 7600 7200
rect 2900 6400 3800 6600
rect -14800 3200 -4000 5400
rect -300 4400 100 5900
rect -3100 100 -900 600
rect 3900 1300 6300 1400
rect 100 1200 6300 1300
rect 100 500 900 1200
rect 900 500 2200 1200
rect 2200 500 3000 1200
rect 3000 500 6300 1200
rect 3900 200 6300 500
rect -5550 -350 -3650 -50
rect -11900 -3200 -11100 -1400
rect -2900 -1200 -1100 -700
rect -2900 -1700 -100 -1200
rect -100 -1700 900 -1200
rect 900 -1700 2300 -1200
rect 2300 -1700 3300 -1200
rect -700 -4700 1200 -2300
rect 2300 -3200 3300 -1700
<< mimcap >>
rect -20500 21800 -10500 21900
rect -20500 13200 -20400 21800
rect -10600 13200 -10500 21800
rect -20500 13100 -10500 13200
rect -3550 7500 -2650 7550
rect -3550 6100 -3500 7500
rect -2700 6100 -2650 7500
rect -3550 6050 -2650 6100
rect -3150 5100 -850 5150
rect -5550 2500 -3650 2550
rect -5550 300 -5500 2500
rect -3700 300 -3650 2500
rect -3150 1100 -3100 5100
rect -900 1100 -850 5100
rect -3150 1050 -850 1100
rect -5550 250 -3650 300
<< mimcapcontact >>
rect -20400 13200 -10600 21800
rect -3500 6100 -2700 7500
rect -5500 300 -3700 2500
rect -3100 1100 -900 5100
<< metal4 >>
rect -18000 23700 -10400 23800
rect -18000 22400 -17900 23700
rect -10500 22400 -10400 23700
rect -18000 22300 -10400 22400
rect -20600 21800 -10400 22200
rect -20600 13200 -20400 21800
rect -10600 15600 -10400 21800
rect -9200 19800 -7600 20000
rect -9200 16600 -9000 19800
rect -7800 17600 -7600 19800
rect -3600 18500 1000 23300
rect -4400 18400 1000 18500
rect -7800 16600 -7200 17600
rect -9200 16400 -7200 16600
rect -4400 16600 -4300 18400
rect 900 16600 1000 18400
rect -4400 16500 1000 16600
rect -10600 13200 -9400 15600
rect -20600 13000 -9400 13200
rect -20600 12400 -4400 13000
rect -20600 11600 -17800 12400
rect -4600 11600 -4400 12400
rect -20600 11400 -4400 11600
rect -3600 12500 1000 16500
rect -3600 10600 -700 12500
rect -21000 9100 -700 10600
rect 900 10000 1000 12500
rect 3500 10100 7700 10200
rect 900 9900 3100 10000
rect 3000 9100 3100 9900
rect -21000 9000 3100 9100
rect -3600 8150 -2600 8200
rect -15000 7800 -4200 8000
rect -3600 7850 -3550 8150
rect -2650 7850 -2600 8150
rect -3600 7800 -2600 7850
rect 3500 8000 3800 10100
rect -15000 3200 -14800 7800
rect -4400 7600 -4200 7800
rect -4400 7500 -2600 7600
rect -4400 7300 -3500 7500
rect -4400 7100 -4200 7300
rect -3600 7100 -3500 7300
rect -4400 6900 -3500 7100
rect -4400 6700 -4200 6900
rect -3600 6700 -3500 6900
rect -4400 6500 -3500 6700
rect -4400 6300 -4200 6500
rect -3600 6300 -3500 6500
rect -4400 6100 -3500 6300
rect -2700 6100 -2600 7500
rect 3500 7300 3600 8000
rect 0 7200 3600 7300
rect 0 6400 100 7200
rect 7600 6600 7700 10100
rect 3800 6500 7700 6600
rect 3800 6400 4000 6500
rect 0 6300 4000 6400
rect -4400 6000 -2600 6100
rect -4400 5600 -4200 6000
rect -400 5900 200 6000
rect -4400 5400 -3800 5600
rect -4000 3200 -3800 5400
rect -400 5200 -300 5900
rect -15000 3000 -3800 3200
rect -5600 2600 -5400 3000
rect -5200 2600 -5000 3000
rect -4800 2600 -4600 3000
rect -4400 2600 -4200 3000
rect -4000 2600 -3800 3000
rect -3200 5100 -300 5200
rect -5600 2500 -3600 2600
rect -5600 300 -5500 2500
rect -3700 300 -3600 2500
rect -3200 1100 -3100 5100
rect -900 4400 -300 5100
rect 100 4400 200 5900
rect -900 4200 200 4400
rect -900 1100 -800 4200
rect 3800 1500 6400 1600
rect 3800 1400 10900 1500
rect -3200 1000 -800 1100
rect 0 1300 3900 1400
rect -5600 200 -3600 300
rect -3200 600 -800 700
rect -3200 100 -3100 600
rect -900 100 -800 600
rect 0 500 100 1300
rect 0 400 3900 500
rect -3200 0 -800 100
rect 3800 200 3900 400
rect 6300 200 10900 1400
rect 3800 0 10900 200
rect -5600 -50 -3600 0
rect -5600 -350 -5550 -50
rect -3650 -350 -3600 -50
rect -5600 -400 -3600 -350
rect 6400 -400 10900 0
rect -3000 -700 -1000 -600
rect -12000 -1400 -11000 -1300
rect -12000 -3200 -11900 -1400
rect -11100 -3200 -11000 -1400
rect -3000 -1700 -2900 -700
rect -1100 -1100 -1000 -700
rect -1100 -1200 3400 -1100
rect -3000 -1800 2300 -1700
rect -12000 -3300 -11000 -3200
rect -800 -2300 1300 -2200
rect -800 -4700 -700 -2300
rect 1200 -4700 1300 -2300
rect 2200 -3200 2300 -1800
rect 3300 -3200 3400 -1200
rect 2200 -3400 3400 -3200
rect -800 -4800 1300 -4700
rect -800 -5000 1200 -4800
<< via4 >>
rect -17900 22400 -10500 23700
rect -3550 7850 -2650 8150
rect 3800 8000 7600 10100
rect -14800 3200 -6200 7800
rect 3800 6900 7600 8000
rect -3100 100 -900 600
rect -5550 -350 -3650 -50
rect -11900 -3200 -11100 -1400
<< mimcap2 >>
rect -20500 21800 -10500 21900
rect -20500 13200 -20400 21800
rect -10600 13200 -10500 21800
rect -20500 13100 -10500 13200
rect -3550 7500 -2650 7550
rect -3550 6100 -3500 7500
rect -2700 6100 -2650 7500
rect -3550 6050 -2650 6100
rect -3150 5100 -850 5150
rect -5550 2500 -3650 2550
rect -5550 300 -5500 2500
rect -3700 300 -3650 2500
rect -3150 1100 -3100 5100
rect -900 1100 -850 5100
rect -3150 1050 -850 1100
rect -5550 250 -3650 300
<< mimcap2contact >>
rect -20400 13200 -10600 21800
rect -3500 6100 -2700 7500
rect -5500 300 -3700 2500
rect -3100 1100 -900 5100
<< metal5 >>
rect -19000 23800 -18400 23900
rect -20600 23700 -10400 23800
rect -20600 22400 -17900 23700
rect -10500 22400 -10400 23700
rect -20600 21800 -10400 22400
rect -20600 13200 -20400 21800
rect -10600 13200 -10400 21800
rect -20600 13000 -10400 13200
rect 3700 10100 7700 10200
rect -3600 8150 -2600 8200
rect -19800 7800 -6000 8000
rect -19800 5800 -14800 7800
rect -19800 3000 -15800 5800
rect -15000 3200 -14800 5800
rect -6200 3200 -6000 7800
rect -3600 7850 -3550 8150
rect -2650 7850 -2600 8150
rect -3600 7500 -2600 7850
rect -3600 6100 -3500 7500
rect -2700 6100 -2600 7500
rect 3700 6900 3800 10100
rect 7600 6900 7700 10100
rect 3700 6800 7700 6900
rect -3600 6000 -2600 6100
rect -15000 3000 -6000 3200
rect -3200 5100 -800 5200
rect -19800 800 -11000 3000
rect -19800 -2000 -15800 800
rect -15000 -1400 -11000 800
rect -5600 2500 -3600 2600
rect -5600 300 -5500 2500
rect -3700 300 -3600 2500
rect -5600 -50 -3600 300
rect -3200 1100 -3100 5100
rect -900 1100 -800 5100
rect -3200 600 -800 1100
rect -3200 100 -3100 600
rect -900 100 -800 600
rect -3200 0 -800 100
rect -5600 -350 -5550 -50
rect -3650 -350 -3600 -50
rect -5600 -400 -3600 -350
rect -15000 -2000 -11900 -1400
rect -19800 -3200 -11900 -2000
rect -11100 -3200 -11000 -1400
rect -800 -3000 1300 -2200
rect -19800 -4200 -11000 -3200
rect -19800 -7000 -15800 -4200
rect -15000 -7000 -11000 -4200
rect -19800 -9200 -11000 -7000
rect -19800 -12000 -15800 -9200
rect -15000 -12000 -11000 -9200
rect -19800 -14200 -11000 -12000
use RF_nfet_8xW5p0L0p15_1  RF_nfet_8xW5p0L0p15_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1661277727
transform 1 0 510 0 -1 2680
box -510 2210 520 3580
use RF_nfet_8xW5p0L0p15_1  RF_nfet_8xW5p0L0p15_1_1
timestamp 1661277727
transform 1 0 2610 0 -1 2680
box -510 2210 520 3580
use RF_nfet_12xW5p0L0p15  RF_nfet_12xW5p0L0p15_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1661277727
transform 1 0 306 0 1 5100
box -506 2200 870 3580
use RF_nfet_12xW5p0L0p15  RF_nfet_12xW5p0L0p15_1
timestamp 1661277727
transform 1 0 2306 0 1 5100
box -506 2200 870 3580
use captuner_complete_1_r  captuner_complete_1_r_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1661915753
transform 1 0 -6860 0 1 16000
box -640 -1200 2480 2400
use sky130_fd_pr__res_generic_po_3AUR5J  sky130_fd_pr__res_generic_po_3AUR5J_0
timestamp 1661638576
transform 1 0 -4039 0 -1 -1345
box -361 -755 361 755
use sky130_fd_pr__res_generic_po_G5R3N7  sky130_fd_pr__res_generic_po_G5R3N7_0
timestamp 1661316842
transform 1 0 -993 0 1 6383
box -307 -743 307 743
use sky130_fd_pr__res_generic_po_G5R3N7  sky130_fd_pr__res_generic_po_G5R3N7_1
timestamp 1661316842
transform 0 1 -2857 -1 0 8807
box -307 -743 307 743
<< labels >>
rlabel metal5 -19800 6700 -15800 8000 1 VLO
rlabel metal5 -19000 23800 -18400 23900 1 VHI
rlabel metal4 -3600 22900 1000 23300 1 VOUT
rlabel metal3 -4300 -900 -4200 -700 1 BIAS_BOT
rlabel metal4 -400 4200 200 6000 1 RFB_MID
rlabel metal1 -1800 8600 -1600 8800 1 G_TOP
rlabel metal2 -5500 18500 -5400 18600 1 G4
rlabel metal2 -5900 18500 -5800 18600 1 G8
rlabel metal2 -6300 18500 -6200 18600 1 G1
rlabel metal2 -6700 18500 -6600 18600 1 G2
rlabel metal4 6400 -400 10900 1500 1 D1
rlabel space 3500 6500 7700 10200 1 S1
rlabel metal1 2200 -1800 2600 -1100 1 VIN
rlabel metal4 -800 -5000 1200 -4800 1 SS
rlabel metal3 -2380 8600 -2080 8840 1 BIAS_TOP
<< end >>
