magic
tech sky130A
magscale 1 2
timestamp 1663768690
<< pwell >>
rect 0 0 5138 6516
<< mvnmos >>
rect 228 258 328 6258
rect 386 258 486 6258
rect 544 258 644 6258
rect 702 258 802 6258
rect 860 258 960 6258
rect 1018 258 1118 6258
rect 1176 258 1276 6258
rect 1334 258 1434 6258
rect 1492 258 1592 6258
rect 1650 258 1750 6258
rect 1808 258 1908 6258
rect 1966 258 2066 6258
rect 2124 258 2224 6258
rect 2282 258 2382 6258
rect 2440 258 2540 6258
rect 2598 258 2698 6258
rect 2756 258 2856 6258
rect 2914 258 3014 6258
rect 3072 258 3172 6258
rect 3230 258 3330 6258
rect 3388 258 3488 6258
rect 3546 258 3646 6258
rect 3704 258 3804 6258
rect 3862 258 3962 6258
rect 4020 258 4120 6258
rect 4178 258 4278 6258
rect 4336 258 4436 6258
rect 4494 258 4594 6258
rect 4652 258 4752 6258
rect 4810 258 4910 6258
<< mvndiff >>
rect 170 6246 228 6258
rect 170 270 182 6246
rect 216 270 228 6246
rect 170 258 228 270
rect 328 6246 386 6258
rect 328 270 340 6246
rect 374 270 386 6246
rect 328 258 386 270
rect 486 6246 544 6258
rect 486 270 498 6246
rect 532 270 544 6246
rect 486 258 544 270
rect 644 6246 702 6258
rect 644 270 656 6246
rect 690 270 702 6246
rect 644 258 702 270
rect 802 6246 860 6258
rect 802 270 814 6246
rect 848 270 860 6246
rect 802 258 860 270
rect 960 6246 1018 6258
rect 960 270 972 6246
rect 1006 270 1018 6246
rect 960 258 1018 270
rect 1118 6246 1176 6258
rect 1118 270 1130 6246
rect 1164 270 1176 6246
rect 1118 258 1176 270
rect 1276 6246 1334 6258
rect 1276 270 1288 6246
rect 1322 270 1334 6246
rect 1276 258 1334 270
rect 1434 6246 1492 6258
rect 1434 270 1446 6246
rect 1480 270 1492 6246
rect 1434 258 1492 270
rect 1592 6246 1650 6258
rect 1592 270 1604 6246
rect 1638 270 1650 6246
rect 1592 258 1650 270
rect 1750 6246 1808 6258
rect 1750 270 1762 6246
rect 1796 270 1808 6246
rect 1750 258 1808 270
rect 1908 6246 1966 6258
rect 1908 270 1920 6246
rect 1954 270 1966 6246
rect 1908 258 1966 270
rect 2066 6246 2124 6258
rect 2066 270 2078 6246
rect 2112 270 2124 6246
rect 2066 258 2124 270
rect 2224 6246 2282 6258
rect 2224 270 2236 6246
rect 2270 270 2282 6246
rect 2224 258 2282 270
rect 2382 6246 2440 6258
rect 2382 270 2394 6246
rect 2428 270 2440 6246
rect 2382 258 2440 270
rect 2540 6246 2598 6258
rect 2540 270 2552 6246
rect 2586 270 2598 6246
rect 2540 258 2598 270
rect 2698 6246 2756 6258
rect 2698 270 2710 6246
rect 2744 270 2756 6246
rect 2698 258 2756 270
rect 2856 6246 2914 6258
rect 2856 270 2868 6246
rect 2902 270 2914 6246
rect 2856 258 2914 270
rect 3014 6246 3072 6258
rect 3014 270 3026 6246
rect 3060 270 3072 6246
rect 3014 258 3072 270
rect 3172 6246 3230 6258
rect 3172 270 3184 6246
rect 3218 270 3230 6246
rect 3172 258 3230 270
rect 3330 6246 3388 6258
rect 3330 270 3342 6246
rect 3376 270 3388 6246
rect 3330 258 3388 270
rect 3488 6246 3546 6258
rect 3488 270 3500 6246
rect 3534 270 3546 6246
rect 3488 258 3546 270
rect 3646 6246 3704 6258
rect 3646 270 3658 6246
rect 3692 270 3704 6246
rect 3646 258 3704 270
rect 3804 6246 3862 6258
rect 3804 270 3816 6246
rect 3850 270 3862 6246
rect 3804 258 3862 270
rect 3962 6246 4020 6258
rect 3962 270 3974 6246
rect 4008 270 4020 6246
rect 3962 258 4020 270
rect 4120 6246 4178 6258
rect 4120 270 4132 6246
rect 4166 270 4178 6246
rect 4120 258 4178 270
rect 4278 6246 4336 6258
rect 4278 270 4290 6246
rect 4324 270 4336 6246
rect 4278 258 4336 270
rect 4436 6246 4494 6258
rect 4436 270 4448 6246
rect 4482 270 4494 6246
rect 4436 258 4494 270
rect 4594 6246 4652 6258
rect 4594 270 4606 6246
rect 4640 270 4652 6246
rect 4594 258 4652 270
rect 4752 6246 4810 6258
rect 4752 270 4764 6246
rect 4798 270 4810 6246
rect 4752 258 4810 270
rect 4910 6246 4968 6258
rect 4910 270 4922 6246
rect 4956 270 4968 6246
rect 4910 258 4968 270
<< mvndiffc >>
rect 182 270 216 6246
rect 340 270 374 6246
rect 498 270 532 6246
rect 656 270 690 6246
rect 814 270 848 6246
rect 972 270 1006 6246
rect 1130 270 1164 6246
rect 1288 270 1322 6246
rect 1446 270 1480 6246
rect 1604 270 1638 6246
rect 1762 270 1796 6246
rect 1920 270 1954 6246
rect 2078 270 2112 6246
rect 2236 270 2270 6246
rect 2394 270 2428 6246
rect 2552 270 2586 6246
rect 2710 270 2744 6246
rect 2868 270 2902 6246
rect 3026 270 3060 6246
rect 3184 270 3218 6246
rect 3342 270 3376 6246
rect 3500 270 3534 6246
rect 3658 270 3692 6246
rect 3816 270 3850 6246
rect 3974 270 4008 6246
rect 4132 270 4166 6246
rect 4290 270 4324 6246
rect 4448 270 4482 6246
rect 4606 270 4640 6246
rect 4764 270 4798 6246
rect 4922 270 4956 6246
<< mvpsubdiff >>
rect 36 6468 5102 6480
rect 36 6434 144 6468
rect 4994 6434 5102 6468
rect 36 6422 5102 6434
rect 36 6372 94 6422
rect 36 144 48 6372
rect 82 144 94 6372
rect 5044 6372 5102 6422
rect 36 94 94 144
rect 5044 144 5056 6372
rect 5090 144 5102 6372
rect 5044 94 5102 144
rect 36 82 5102 94
rect 36 48 144 82
rect 4994 48 5102 82
rect 36 36 5102 48
<< mvpsubdiffcont >>
rect 144 6434 4994 6468
rect 48 144 82 6372
rect 5056 144 5090 6372
rect 144 48 4994 82
<< poly >>
rect 228 6330 328 6346
rect 228 6296 244 6330
rect 312 6296 328 6330
rect 228 6258 328 6296
rect 386 6330 486 6346
rect 386 6296 402 6330
rect 470 6296 486 6330
rect 386 6258 486 6296
rect 544 6330 644 6346
rect 544 6296 560 6330
rect 628 6296 644 6330
rect 544 6258 644 6296
rect 702 6330 802 6346
rect 702 6296 718 6330
rect 786 6296 802 6330
rect 702 6258 802 6296
rect 860 6330 960 6346
rect 860 6296 876 6330
rect 944 6296 960 6330
rect 860 6258 960 6296
rect 1018 6330 1118 6346
rect 1018 6296 1034 6330
rect 1102 6296 1118 6330
rect 1018 6258 1118 6296
rect 1176 6330 1276 6346
rect 1176 6296 1192 6330
rect 1260 6296 1276 6330
rect 1176 6258 1276 6296
rect 1334 6330 1434 6346
rect 1334 6296 1350 6330
rect 1418 6296 1434 6330
rect 1334 6258 1434 6296
rect 1492 6330 1592 6346
rect 1492 6296 1508 6330
rect 1576 6296 1592 6330
rect 1492 6258 1592 6296
rect 1650 6330 1750 6346
rect 1650 6296 1666 6330
rect 1734 6296 1750 6330
rect 1650 6258 1750 6296
rect 1808 6330 1908 6346
rect 1808 6296 1824 6330
rect 1892 6296 1908 6330
rect 1808 6258 1908 6296
rect 1966 6330 2066 6346
rect 1966 6296 1982 6330
rect 2050 6296 2066 6330
rect 1966 6258 2066 6296
rect 2124 6330 2224 6346
rect 2124 6296 2140 6330
rect 2208 6296 2224 6330
rect 2124 6258 2224 6296
rect 2282 6330 2382 6346
rect 2282 6296 2298 6330
rect 2366 6296 2382 6330
rect 2282 6258 2382 6296
rect 2440 6330 2540 6346
rect 2440 6296 2456 6330
rect 2524 6296 2540 6330
rect 2440 6258 2540 6296
rect 2598 6330 2698 6346
rect 2598 6296 2614 6330
rect 2682 6296 2698 6330
rect 2598 6258 2698 6296
rect 2756 6330 2856 6346
rect 2756 6296 2772 6330
rect 2840 6296 2856 6330
rect 2756 6258 2856 6296
rect 2914 6330 3014 6346
rect 2914 6296 2930 6330
rect 2998 6296 3014 6330
rect 2914 6258 3014 6296
rect 3072 6330 3172 6346
rect 3072 6296 3088 6330
rect 3156 6296 3172 6330
rect 3072 6258 3172 6296
rect 3230 6330 3330 6346
rect 3230 6296 3246 6330
rect 3314 6296 3330 6330
rect 3230 6258 3330 6296
rect 3388 6330 3488 6346
rect 3388 6296 3404 6330
rect 3472 6296 3488 6330
rect 3388 6258 3488 6296
rect 3546 6330 3646 6346
rect 3546 6296 3562 6330
rect 3630 6296 3646 6330
rect 3546 6258 3646 6296
rect 3704 6330 3804 6346
rect 3704 6296 3720 6330
rect 3788 6296 3804 6330
rect 3704 6258 3804 6296
rect 3862 6330 3962 6346
rect 3862 6296 3878 6330
rect 3946 6296 3962 6330
rect 3862 6258 3962 6296
rect 4020 6330 4120 6346
rect 4020 6296 4036 6330
rect 4104 6296 4120 6330
rect 4020 6258 4120 6296
rect 4178 6330 4278 6346
rect 4178 6296 4194 6330
rect 4262 6296 4278 6330
rect 4178 6258 4278 6296
rect 4336 6330 4436 6346
rect 4336 6296 4352 6330
rect 4420 6296 4436 6330
rect 4336 6258 4436 6296
rect 4494 6330 4594 6346
rect 4494 6296 4510 6330
rect 4578 6296 4594 6330
rect 4494 6258 4594 6296
rect 4652 6330 4752 6346
rect 4652 6296 4668 6330
rect 4736 6296 4752 6330
rect 4652 6258 4752 6296
rect 4810 6330 4910 6346
rect 4810 6296 4826 6330
rect 4894 6296 4910 6330
rect 4810 6258 4910 6296
rect 228 220 328 258
rect 228 186 244 220
rect 312 186 328 220
rect 228 170 328 186
rect 386 220 486 258
rect 386 186 402 220
rect 470 186 486 220
rect 386 170 486 186
rect 544 220 644 258
rect 544 186 560 220
rect 628 186 644 220
rect 544 170 644 186
rect 702 220 802 258
rect 702 186 718 220
rect 786 186 802 220
rect 702 170 802 186
rect 860 220 960 258
rect 860 186 876 220
rect 944 186 960 220
rect 860 170 960 186
rect 1018 220 1118 258
rect 1018 186 1034 220
rect 1102 186 1118 220
rect 1018 170 1118 186
rect 1176 220 1276 258
rect 1176 186 1192 220
rect 1260 186 1276 220
rect 1176 170 1276 186
rect 1334 220 1434 258
rect 1334 186 1350 220
rect 1418 186 1434 220
rect 1334 170 1434 186
rect 1492 220 1592 258
rect 1492 186 1508 220
rect 1576 186 1592 220
rect 1492 170 1592 186
rect 1650 220 1750 258
rect 1650 186 1666 220
rect 1734 186 1750 220
rect 1650 170 1750 186
rect 1808 220 1908 258
rect 1808 186 1824 220
rect 1892 186 1908 220
rect 1808 170 1908 186
rect 1966 220 2066 258
rect 1966 186 1982 220
rect 2050 186 2066 220
rect 1966 170 2066 186
rect 2124 220 2224 258
rect 2124 186 2140 220
rect 2208 186 2224 220
rect 2124 170 2224 186
rect 2282 220 2382 258
rect 2282 186 2298 220
rect 2366 186 2382 220
rect 2282 170 2382 186
rect 2440 220 2540 258
rect 2440 186 2456 220
rect 2524 186 2540 220
rect 2440 170 2540 186
rect 2598 220 2698 258
rect 2598 186 2614 220
rect 2682 186 2698 220
rect 2598 170 2698 186
rect 2756 220 2856 258
rect 2756 186 2772 220
rect 2840 186 2856 220
rect 2756 170 2856 186
rect 2914 220 3014 258
rect 2914 186 2930 220
rect 2998 186 3014 220
rect 2914 170 3014 186
rect 3072 220 3172 258
rect 3072 186 3088 220
rect 3156 186 3172 220
rect 3072 170 3172 186
rect 3230 220 3330 258
rect 3230 186 3246 220
rect 3314 186 3330 220
rect 3230 170 3330 186
rect 3388 220 3488 258
rect 3388 186 3404 220
rect 3472 186 3488 220
rect 3388 170 3488 186
rect 3546 220 3646 258
rect 3546 186 3562 220
rect 3630 186 3646 220
rect 3546 170 3646 186
rect 3704 220 3804 258
rect 3704 186 3720 220
rect 3788 186 3804 220
rect 3704 170 3804 186
rect 3862 220 3962 258
rect 3862 186 3878 220
rect 3946 186 3962 220
rect 3862 170 3962 186
rect 4020 220 4120 258
rect 4020 186 4036 220
rect 4104 186 4120 220
rect 4020 170 4120 186
rect 4178 220 4278 258
rect 4178 186 4194 220
rect 4262 186 4278 220
rect 4178 170 4278 186
rect 4336 220 4436 258
rect 4336 186 4352 220
rect 4420 186 4436 220
rect 4336 170 4436 186
rect 4494 220 4594 258
rect 4494 186 4510 220
rect 4578 186 4594 220
rect 4494 170 4594 186
rect 4652 220 4752 258
rect 4652 186 4668 220
rect 4736 186 4752 220
rect 4652 170 4752 186
rect 4810 220 4910 258
rect 4810 186 4826 220
rect 4894 186 4910 220
rect 4810 170 4910 186
<< polycont >>
rect 244 6296 312 6330
rect 402 6296 470 6330
rect 560 6296 628 6330
rect 718 6296 786 6330
rect 876 6296 944 6330
rect 1034 6296 1102 6330
rect 1192 6296 1260 6330
rect 1350 6296 1418 6330
rect 1508 6296 1576 6330
rect 1666 6296 1734 6330
rect 1824 6296 1892 6330
rect 1982 6296 2050 6330
rect 2140 6296 2208 6330
rect 2298 6296 2366 6330
rect 2456 6296 2524 6330
rect 2614 6296 2682 6330
rect 2772 6296 2840 6330
rect 2930 6296 2998 6330
rect 3088 6296 3156 6330
rect 3246 6296 3314 6330
rect 3404 6296 3472 6330
rect 3562 6296 3630 6330
rect 3720 6296 3788 6330
rect 3878 6296 3946 6330
rect 4036 6296 4104 6330
rect 4194 6296 4262 6330
rect 4352 6296 4420 6330
rect 4510 6296 4578 6330
rect 4668 6296 4736 6330
rect 4826 6296 4894 6330
rect 244 186 312 220
rect 402 186 470 220
rect 560 186 628 220
rect 718 186 786 220
rect 876 186 944 220
rect 1034 186 1102 220
rect 1192 186 1260 220
rect 1350 186 1418 220
rect 1508 186 1576 220
rect 1666 186 1734 220
rect 1824 186 1892 220
rect 1982 186 2050 220
rect 2140 186 2208 220
rect 2298 186 2366 220
rect 2456 186 2524 220
rect 2614 186 2682 220
rect 2772 186 2840 220
rect 2930 186 2998 220
rect 3088 186 3156 220
rect 3246 186 3314 220
rect 3404 186 3472 220
rect 3562 186 3630 220
rect 3720 186 3788 220
rect 3878 186 3946 220
rect 4036 186 4104 220
rect 4194 186 4262 220
rect 4352 186 4420 220
rect 4510 186 4578 220
rect 4668 186 4736 220
rect 4826 186 4894 220
<< locali >>
rect 48 6434 144 6468
rect 4994 6434 5090 6468
rect 48 6372 82 6434
rect 5056 6372 5090 6434
rect 228 6296 244 6330
rect 312 6296 328 6330
rect 386 6296 402 6330
rect 470 6296 486 6330
rect 544 6296 560 6330
rect 628 6296 644 6330
rect 702 6296 718 6330
rect 786 6296 802 6330
rect 860 6296 876 6330
rect 944 6296 960 6330
rect 1018 6296 1034 6330
rect 1102 6296 1118 6330
rect 1176 6296 1192 6330
rect 1260 6296 1276 6330
rect 1334 6296 1350 6330
rect 1418 6296 1434 6330
rect 1492 6296 1508 6330
rect 1576 6296 1592 6330
rect 1650 6296 1666 6330
rect 1734 6296 1750 6330
rect 1808 6296 1824 6330
rect 1892 6296 1908 6330
rect 1966 6296 1982 6330
rect 2050 6296 2066 6330
rect 2124 6296 2140 6330
rect 2208 6296 2224 6330
rect 2282 6296 2298 6330
rect 2366 6296 2382 6330
rect 2440 6296 2456 6330
rect 2524 6296 2540 6330
rect 2598 6296 2614 6330
rect 2682 6296 2698 6330
rect 2756 6296 2772 6330
rect 2840 6296 2856 6330
rect 2914 6296 2930 6330
rect 2998 6296 3014 6330
rect 3072 6296 3088 6330
rect 3156 6296 3172 6330
rect 3230 6296 3246 6330
rect 3314 6296 3330 6330
rect 3388 6296 3404 6330
rect 3472 6296 3488 6330
rect 3546 6296 3562 6330
rect 3630 6296 3646 6330
rect 3704 6296 3720 6330
rect 3788 6296 3804 6330
rect 3862 6296 3878 6330
rect 3946 6296 3962 6330
rect 4020 6296 4036 6330
rect 4104 6296 4120 6330
rect 4178 6296 4194 6330
rect 4262 6296 4278 6330
rect 4336 6296 4352 6330
rect 4420 6296 4436 6330
rect 4494 6296 4510 6330
rect 4578 6296 4594 6330
rect 4652 6296 4668 6330
rect 4736 6296 4752 6330
rect 4810 6296 4826 6330
rect 4894 6296 4910 6330
rect 182 6246 216 6262
rect 182 254 216 270
rect 340 6246 374 6262
rect 340 254 374 270
rect 498 6246 532 6262
rect 498 254 532 270
rect 656 6246 690 6262
rect 656 254 690 270
rect 814 6246 848 6262
rect 814 254 848 270
rect 972 6246 1006 6262
rect 972 254 1006 270
rect 1130 6246 1164 6262
rect 1130 254 1164 270
rect 1288 6246 1322 6262
rect 1288 254 1322 270
rect 1446 6246 1480 6262
rect 1446 254 1480 270
rect 1604 6246 1638 6262
rect 1604 254 1638 270
rect 1762 6246 1796 6262
rect 1762 254 1796 270
rect 1920 6246 1954 6262
rect 1920 254 1954 270
rect 2078 6246 2112 6262
rect 2078 254 2112 270
rect 2236 6246 2270 6262
rect 2236 254 2270 270
rect 2394 6246 2428 6262
rect 2394 254 2428 270
rect 2552 6246 2586 6262
rect 2552 254 2586 270
rect 2710 6246 2744 6262
rect 2710 254 2744 270
rect 2868 6246 2902 6262
rect 2868 254 2902 270
rect 3026 6246 3060 6262
rect 3026 254 3060 270
rect 3184 6246 3218 6262
rect 3184 254 3218 270
rect 3342 6246 3376 6262
rect 3342 254 3376 270
rect 3500 6246 3534 6262
rect 3500 254 3534 270
rect 3658 6246 3692 6262
rect 3658 254 3692 270
rect 3816 6246 3850 6262
rect 3816 254 3850 270
rect 3974 6246 4008 6262
rect 3974 254 4008 270
rect 4132 6246 4166 6262
rect 4132 254 4166 270
rect 4290 6246 4324 6262
rect 4290 254 4324 270
rect 4448 6246 4482 6262
rect 4448 254 4482 270
rect 4606 6246 4640 6262
rect 4606 254 4640 270
rect 4764 6246 4798 6262
rect 4764 254 4798 270
rect 4922 6246 4956 6262
rect 4922 254 4956 270
rect 228 186 244 220
rect 312 186 328 220
rect 386 186 402 220
rect 470 186 486 220
rect 544 186 560 220
rect 628 186 644 220
rect 702 186 718 220
rect 786 186 802 220
rect 860 186 876 220
rect 944 186 960 220
rect 1018 186 1034 220
rect 1102 186 1118 220
rect 1176 186 1192 220
rect 1260 186 1276 220
rect 1334 186 1350 220
rect 1418 186 1434 220
rect 1492 186 1508 220
rect 1576 186 1592 220
rect 1650 186 1666 220
rect 1734 186 1750 220
rect 1808 186 1824 220
rect 1892 186 1908 220
rect 1966 186 1982 220
rect 2050 186 2066 220
rect 2124 186 2140 220
rect 2208 186 2224 220
rect 2282 186 2298 220
rect 2366 186 2382 220
rect 2440 186 2456 220
rect 2524 186 2540 220
rect 2598 186 2614 220
rect 2682 186 2698 220
rect 2756 186 2772 220
rect 2840 186 2856 220
rect 2914 186 2930 220
rect 2998 186 3014 220
rect 3072 186 3088 220
rect 3156 186 3172 220
rect 3230 186 3246 220
rect 3314 186 3330 220
rect 3388 186 3404 220
rect 3472 186 3488 220
rect 3546 186 3562 220
rect 3630 186 3646 220
rect 3704 186 3720 220
rect 3788 186 3804 220
rect 3862 186 3878 220
rect 3946 186 3962 220
rect 4020 186 4036 220
rect 4104 186 4120 220
rect 4178 186 4194 220
rect 4262 186 4278 220
rect 4336 186 4352 220
rect 4420 186 4436 220
rect 4494 186 4510 220
rect 4578 186 4594 220
rect 4652 186 4668 220
rect 4736 186 4752 220
rect 4810 186 4826 220
rect 4894 186 4910 220
rect 48 82 82 144
rect 5056 82 5090 144
rect 48 48 144 82
rect 4994 48 5090 82
<< viali >>
rect 236 6468 4959 6470
rect 236 6434 4959 6468
rect 236 6432 4959 6434
rect 244 6296 312 6330
rect 402 6296 470 6330
rect 560 6296 628 6330
rect 718 6296 786 6330
rect 876 6296 944 6330
rect 1034 6296 1102 6330
rect 1192 6296 1260 6330
rect 1350 6296 1418 6330
rect 1508 6296 1576 6330
rect 1666 6296 1734 6330
rect 1824 6296 1892 6330
rect 1982 6296 2050 6330
rect 2140 6296 2208 6330
rect 2298 6296 2366 6330
rect 2456 6296 2524 6330
rect 2614 6296 2682 6330
rect 2772 6296 2840 6330
rect 2930 6296 2998 6330
rect 3088 6296 3156 6330
rect 3246 6296 3314 6330
rect 3404 6296 3472 6330
rect 3562 6296 3630 6330
rect 3720 6296 3788 6330
rect 3878 6296 3946 6330
rect 4036 6296 4104 6330
rect 4194 6296 4262 6330
rect 4352 6296 4420 6330
rect 4510 6296 4578 6330
rect 4668 6296 4736 6330
rect 4826 6296 4894 6330
rect 46 236 48 6280
rect 48 236 82 6280
rect 82 236 84 6280
rect 182 270 216 6246
rect 340 270 374 6246
rect 498 270 532 6246
rect 656 270 690 6246
rect 814 270 848 6246
rect 972 270 1006 6246
rect 1130 270 1164 6246
rect 1288 270 1322 6246
rect 1446 270 1480 6246
rect 1604 270 1638 6246
rect 1762 270 1796 6246
rect 1920 270 1954 6246
rect 2078 270 2112 6246
rect 2236 270 2270 6246
rect 2394 270 2428 6246
rect 2552 270 2586 6246
rect 2710 270 2744 6246
rect 2868 270 2902 6246
rect 3026 270 3060 6246
rect 3184 270 3218 6246
rect 3342 270 3376 6246
rect 3500 270 3534 6246
rect 3658 270 3692 6246
rect 3816 270 3850 6246
rect 3974 270 4008 6246
rect 4132 270 4166 6246
rect 4290 270 4324 6246
rect 4448 270 4482 6246
rect 4606 270 4640 6246
rect 4764 270 4798 6246
rect 4922 270 4956 6246
rect 5054 236 5056 6280
rect 5056 236 5090 6280
rect 5090 236 5092 6280
rect 244 186 312 220
rect 402 186 470 220
rect 560 186 628 220
rect 718 186 786 220
rect 876 186 944 220
rect 1034 186 1102 220
rect 1192 186 1260 220
rect 1350 186 1418 220
rect 1508 186 1576 220
rect 1666 186 1734 220
rect 1824 186 1892 220
rect 1982 186 2050 220
rect 2140 186 2208 220
rect 2298 186 2366 220
rect 2456 186 2524 220
rect 2614 186 2682 220
rect 2772 186 2840 220
rect 2930 186 2998 220
rect 3088 186 3156 220
rect 3246 186 3314 220
rect 3404 186 3472 220
rect 3562 186 3630 220
rect 3720 186 3788 220
rect 3878 186 3946 220
rect 4036 186 4104 220
rect 4194 186 4262 220
rect 4352 186 4420 220
rect 4510 186 4578 220
rect 4668 186 4736 220
rect 4826 186 4894 220
rect 236 82 4902 84
rect 236 48 4902 82
rect 236 46 4902 48
<< metal1 >>
rect 30 6470 5110 6480
rect 30 6432 236 6470
rect 4959 6432 5110 6470
rect 30 6422 5110 6432
rect 30 6420 100 6422
rect 5040 6420 5110 6422
rect 232 6330 252 6390
rect 4886 6330 4906 6390
rect 232 6296 244 6330
rect 4894 6296 4906 6330
rect 232 6290 252 6296
rect 4886 6290 4906 6296
rect 165 6246 231 6258
rect 165 6238 182 6246
rect 216 6238 231 6246
rect 165 270 182 278
rect 216 270 231 278
rect 165 258 231 270
rect 323 6246 389 6258
rect 323 6238 340 6246
rect 374 6238 389 6246
rect 323 270 340 278
rect 374 270 389 278
rect 323 258 389 270
rect 481 6246 547 6258
rect 481 6238 498 6246
rect 532 6238 547 6246
rect 481 270 498 278
rect 532 270 547 278
rect 481 258 547 270
rect 639 6246 705 6258
rect 639 6238 656 6246
rect 690 6238 705 6246
rect 639 270 656 278
rect 690 270 705 278
rect 639 258 705 270
rect 797 6246 863 6258
rect 797 6238 814 6246
rect 848 6238 863 6246
rect 797 270 814 278
rect 848 270 863 278
rect 797 258 863 270
rect 955 6246 1021 6258
rect 955 6238 972 6246
rect 1006 6238 1021 6246
rect 955 270 972 278
rect 1006 270 1021 278
rect 955 258 1021 270
rect 1113 6246 1179 6258
rect 1113 6238 1130 6246
rect 1164 6238 1179 6246
rect 1113 270 1130 278
rect 1164 270 1179 278
rect 1113 258 1179 270
rect 1271 6246 1337 6258
rect 1271 6238 1288 6246
rect 1322 6238 1337 6246
rect 1271 270 1288 278
rect 1322 270 1337 278
rect 1271 258 1337 270
rect 1429 6246 1495 6258
rect 1429 6238 1446 6246
rect 1480 6238 1495 6246
rect 1429 270 1446 278
rect 1480 270 1495 278
rect 1429 258 1495 270
rect 1587 6246 1653 6258
rect 1587 6238 1604 6246
rect 1638 6238 1653 6246
rect 1587 270 1604 278
rect 1638 270 1653 278
rect 1587 258 1653 270
rect 1745 6246 1811 6258
rect 1745 6238 1762 6246
rect 1796 6238 1811 6246
rect 1745 270 1762 278
rect 1796 270 1811 278
rect 1745 258 1811 270
rect 1903 6246 1969 6258
rect 1903 6238 1920 6246
rect 1954 6238 1969 6246
rect 1903 270 1920 278
rect 1954 270 1969 278
rect 1903 258 1969 270
rect 2061 6246 2127 6258
rect 2061 6238 2078 6246
rect 2112 6238 2127 6246
rect 2061 270 2078 278
rect 2112 270 2127 278
rect 2061 258 2127 270
rect 2219 6246 2285 6258
rect 2219 6238 2236 6246
rect 2270 6238 2285 6246
rect 2219 270 2236 278
rect 2270 270 2285 278
rect 2219 258 2285 270
rect 2377 6246 2443 6258
rect 2377 6238 2394 6246
rect 2428 6238 2443 6246
rect 2377 270 2394 278
rect 2428 270 2443 278
rect 2377 258 2443 270
rect 2535 6246 2601 6258
rect 2535 6238 2552 6246
rect 2586 6238 2601 6246
rect 2535 270 2552 278
rect 2586 270 2601 278
rect 2535 258 2601 270
rect 2693 6246 2759 6258
rect 2693 6238 2710 6246
rect 2744 6238 2759 6246
rect 2693 270 2710 278
rect 2744 270 2759 278
rect 2693 258 2759 270
rect 2851 6246 2917 6258
rect 2851 6238 2868 6246
rect 2902 6238 2917 6246
rect 2851 270 2868 278
rect 2902 270 2917 278
rect 2851 258 2917 270
rect 3009 6246 3075 6258
rect 3009 6238 3026 6246
rect 3060 6238 3075 6246
rect 3009 270 3026 278
rect 3060 270 3075 278
rect 3009 258 3075 270
rect 3167 6246 3233 6258
rect 3167 6238 3184 6246
rect 3218 6238 3233 6246
rect 3167 270 3184 278
rect 3218 270 3233 278
rect 3167 258 3233 270
rect 3325 6246 3391 6258
rect 3325 6238 3342 6246
rect 3376 6238 3391 6246
rect 3325 270 3342 278
rect 3376 270 3391 278
rect 3325 258 3391 270
rect 3483 6246 3549 6258
rect 3483 6238 3500 6246
rect 3534 6238 3549 6246
rect 3483 270 3500 278
rect 3534 270 3549 278
rect 3483 258 3549 270
rect 3641 6246 3707 6258
rect 3641 6238 3658 6246
rect 3692 6238 3707 6246
rect 3641 270 3658 278
rect 3692 270 3707 278
rect 3641 258 3707 270
rect 3799 6246 3865 6258
rect 3799 6238 3816 6246
rect 3850 6238 3865 6246
rect 3799 270 3816 278
rect 3850 270 3865 278
rect 3799 258 3865 270
rect 3957 6246 4023 6258
rect 3957 6238 3974 6246
rect 4008 6238 4023 6246
rect 3957 270 3974 278
rect 4008 270 4023 278
rect 3957 258 4023 270
rect 4115 6246 4181 6258
rect 4115 6238 4132 6246
rect 4166 6238 4181 6246
rect 4115 270 4132 278
rect 4166 270 4181 278
rect 4115 258 4181 270
rect 4273 6246 4339 6258
rect 4273 6238 4290 6246
rect 4324 6238 4339 6246
rect 4273 270 4290 278
rect 4324 270 4339 278
rect 4273 258 4339 270
rect 4431 6246 4497 6258
rect 4431 6238 4448 6246
rect 4482 6238 4497 6246
rect 4431 270 4448 278
rect 4482 270 4497 278
rect 4431 258 4497 270
rect 4589 6246 4655 6258
rect 4589 6238 4606 6246
rect 4640 6238 4655 6246
rect 4589 270 4606 278
rect 4640 270 4655 278
rect 4589 258 4655 270
rect 4747 6246 4813 6258
rect 4747 6238 4764 6246
rect 4798 6238 4813 6246
rect 4747 270 4764 278
rect 4798 270 4813 278
rect 4747 258 4813 270
rect 4905 6246 4971 6258
rect 4905 6238 4922 6246
rect 4956 6238 4971 6246
rect 4905 270 4922 278
rect 4956 270 4971 278
rect 4905 258 4971 270
rect 232 220 252 226
rect 4886 220 4906 226
rect 232 186 244 220
rect 4894 186 4906 220
rect 232 126 252 186
rect 4886 126 4906 186
rect 30 94 100 100
rect 5040 94 5110 100
rect 30 84 5110 94
rect 30 46 236 84
rect 4902 46 5110 84
rect 30 30 5110 46
<< via1 >>
rect 30 6280 100 6420
rect 252 6330 4886 6390
rect 252 6296 312 6330
rect 312 6296 402 6330
rect 402 6296 470 6330
rect 470 6296 560 6330
rect 560 6296 628 6330
rect 628 6296 718 6330
rect 718 6296 786 6330
rect 786 6296 876 6330
rect 876 6296 944 6330
rect 944 6296 1034 6330
rect 1034 6296 1102 6330
rect 1102 6296 1192 6330
rect 1192 6296 1260 6330
rect 1260 6296 1350 6330
rect 1350 6296 1418 6330
rect 1418 6296 1508 6330
rect 1508 6296 1576 6330
rect 1576 6296 1666 6330
rect 1666 6296 1734 6330
rect 1734 6296 1824 6330
rect 1824 6296 1892 6330
rect 1892 6296 1982 6330
rect 1982 6296 2050 6330
rect 2050 6296 2140 6330
rect 2140 6296 2208 6330
rect 2208 6296 2298 6330
rect 2298 6296 2366 6330
rect 2366 6296 2456 6330
rect 2456 6296 2524 6330
rect 2524 6296 2614 6330
rect 2614 6296 2682 6330
rect 2682 6296 2772 6330
rect 2772 6296 2840 6330
rect 2840 6296 2930 6330
rect 2930 6296 2998 6330
rect 2998 6296 3088 6330
rect 3088 6296 3156 6330
rect 3156 6296 3246 6330
rect 3246 6296 3314 6330
rect 3314 6296 3404 6330
rect 3404 6296 3472 6330
rect 3472 6296 3562 6330
rect 3562 6296 3630 6330
rect 3630 6296 3720 6330
rect 3720 6296 3788 6330
rect 3788 6296 3878 6330
rect 3878 6296 3946 6330
rect 3946 6296 4036 6330
rect 4036 6296 4104 6330
rect 4104 6296 4194 6330
rect 4194 6296 4262 6330
rect 4262 6296 4352 6330
rect 4352 6296 4420 6330
rect 4420 6296 4510 6330
rect 4510 6296 4578 6330
rect 4578 6296 4668 6330
rect 4668 6296 4736 6330
rect 4736 6296 4826 6330
rect 4826 6296 4886 6330
rect 252 6290 4886 6296
rect 30 236 46 6280
rect 46 236 84 6280
rect 84 236 100 6280
rect 5040 6280 5110 6420
rect 165 278 182 6238
rect 182 278 216 6238
rect 216 278 231 6238
rect 323 278 340 6238
rect 340 278 374 6238
rect 374 278 389 6238
rect 481 278 498 6238
rect 498 278 532 6238
rect 532 278 547 6238
rect 639 278 656 6238
rect 656 278 690 6238
rect 690 278 705 6238
rect 797 278 814 6238
rect 814 278 848 6238
rect 848 278 863 6238
rect 955 278 972 6238
rect 972 278 1006 6238
rect 1006 278 1021 6238
rect 1113 278 1130 6238
rect 1130 278 1164 6238
rect 1164 278 1179 6238
rect 1271 278 1288 6238
rect 1288 278 1322 6238
rect 1322 278 1337 6238
rect 1429 278 1446 6238
rect 1446 278 1480 6238
rect 1480 278 1495 6238
rect 1587 278 1604 6238
rect 1604 278 1638 6238
rect 1638 278 1653 6238
rect 1745 278 1762 6238
rect 1762 278 1796 6238
rect 1796 278 1811 6238
rect 1903 278 1920 6238
rect 1920 278 1954 6238
rect 1954 278 1969 6238
rect 2061 278 2078 6238
rect 2078 278 2112 6238
rect 2112 278 2127 6238
rect 2219 278 2236 6238
rect 2236 278 2270 6238
rect 2270 278 2285 6238
rect 2377 278 2394 6238
rect 2394 278 2428 6238
rect 2428 278 2443 6238
rect 2535 278 2552 6238
rect 2552 278 2586 6238
rect 2586 278 2601 6238
rect 2693 278 2710 6238
rect 2710 278 2744 6238
rect 2744 278 2759 6238
rect 2851 278 2868 6238
rect 2868 278 2902 6238
rect 2902 278 2917 6238
rect 3009 278 3026 6238
rect 3026 278 3060 6238
rect 3060 278 3075 6238
rect 3167 278 3184 6238
rect 3184 278 3218 6238
rect 3218 278 3233 6238
rect 3325 278 3342 6238
rect 3342 278 3376 6238
rect 3376 278 3391 6238
rect 3483 278 3500 6238
rect 3500 278 3534 6238
rect 3534 278 3549 6238
rect 3641 278 3658 6238
rect 3658 278 3692 6238
rect 3692 278 3707 6238
rect 3799 278 3816 6238
rect 3816 278 3850 6238
rect 3850 278 3865 6238
rect 3957 278 3974 6238
rect 3974 278 4008 6238
rect 4008 278 4023 6238
rect 4115 278 4132 6238
rect 4132 278 4166 6238
rect 4166 278 4181 6238
rect 4273 278 4290 6238
rect 4290 278 4324 6238
rect 4324 278 4339 6238
rect 4431 278 4448 6238
rect 4448 278 4482 6238
rect 4482 278 4497 6238
rect 4589 278 4606 6238
rect 4606 278 4640 6238
rect 4640 278 4655 6238
rect 4747 278 4764 6238
rect 4764 278 4798 6238
rect 4798 278 4813 6238
rect 4905 278 4922 6238
rect 4922 278 4956 6238
rect 4956 278 4971 6238
rect 30 100 100 236
rect 5040 236 5054 6280
rect 5054 236 5092 6280
rect 5092 236 5110 6280
rect 252 220 4886 226
rect 252 186 312 220
rect 312 186 402 220
rect 402 186 470 220
rect 470 186 560 220
rect 560 186 628 220
rect 628 186 718 220
rect 718 186 786 220
rect 786 186 876 220
rect 876 186 944 220
rect 944 186 1034 220
rect 1034 186 1102 220
rect 1102 186 1192 220
rect 1192 186 1260 220
rect 1260 186 1350 220
rect 1350 186 1418 220
rect 1418 186 1508 220
rect 1508 186 1576 220
rect 1576 186 1666 220
rect 1666 186 1734 220
rect 1734 186 1824 220
rect 1824 186 1892 220
rect 1892 186 1982 220
rect 1982 186 2050 220
rect 2050 186 2140 220
rect 2140 186 2208 220
rect 2208 186 2298 220
rect 2298 186 2366 220
rect 2366 186 2456 220
rect 2456 186 2524 220
rect 2524 186 2614 220
rect 2614 186 2682 220
rect 2682 186 2772 220
rect 2772 186 2840 220
rect 2840 186 2930 220
rect 2930 186 2998 220
rect 2998 186 3088 220
rect 3088 186 3156 220
rect 3156 186 3246 220
rect 3246 186 3314 220
rect 3314 186 3404 220
rect 3404 186 3472 220
rect 3472 186 3562 220
rect 3562 186 3630 220
rect 3630 186 3720 220
rect 3720 186 3788 220
rect 3788 186 3878 220
rect 3878 186 3946 220
rect 3946 186 4036 220
rect 4036 186 4104 220
rect 4104 186 4194 220
rect 4194 186 4262 220
rect 4262 186 4352 220
rect 4352 186 4420 220
rect 4420 186 4510 220
rect 4510 186 4578 220
rect 4578 186 4668 220
rect 4668 186 4736 220
rect 4736 186 4826 220
rect 4826 186 4886 220
rect 252 126 4886 186
rect 5040 100 5110 236
<< metal2 >>
rect 30 6420 100 6480
rect 5040 6420 5110 6480
rect 232 6380 252 6390
rect 4886 6380 4906 6390
rect 232 6310 240 6380
rect 4900 6310 4906 6380
rect 232 6290 252 6310
rect 4886 6290 4906 6310
rect 165 6238 231 6258
rect 165 258 231 278
rect 323 6238 389 6258
rect 323 258 389 278
rect 481 6238 547 6258
rect 481 258 547 278
rect 639 6238 705 6258
rect 639 258 705 278
rect 797 6238 863 6258
rect 797 258 863 278
rect 955 6238 1021 6258
rect 955 258 1021 278
rect 1113 6238 1179 6258
rect 1113 258 1179 278
rect 1271 6238 1337 6258
rect 1271 258 1337 278
rect 1429 6238 1495 6258
rect 1429 258 1495 278
rect 1587 6238 1653 6258
rect 1587 258 1653 278
rect 1745 6238 1811 6258
rect 1745 258 1811 278
rect 1903 6238 1969 6258
rect 1903 258 1969 278
rect 2061 6238 2127 6258
rect 2061 258 2127 278
rect 2219 6238 2285 6258
rect 2219 258 2285 278
rect 2377 6238 2443 6258
rect 2377 258 2443 278
rect 2535 6238 2601 6258
rect 2535 258 2601 278
rect 2693 6238 2759 6258
rect 2693 258 2759 278
rect 2851 6238 2917 6258
rect 2851 258 2917 278
rect 3009 6238 3075 6258
rect 3009 258 3075 278
rect 3167 6238 3233 6258
rect 3167 258 3233 278
rect 3325 6238 3391 6258
rect 3325 258 3391 278
rect 3483 6238 3549 6258
rect 3483 258 3549 278
rect 3641 6238 3707 6258
rect 3641 258 3707 278
rect 3799 6238 3865 6258
rect 3799 258 3865 278
rect 3957 6238 4023 6258
rect 3957 258 4023 278
rect 4115 6238 4181 6258
rect 4115 258 4181 278
rect 4273 6238 4339 6258
rect 4273 258 4339 278
rect 4431 6238 4497 6258
rect 4431 258 4497 278
rect 4589 6238 4655 6258
rect 4589 258 4655 278
rect 4747 6238 4813 6258
rect 4747 258 4813 278
rect 4905 6238 4971 6258
rect 4905 258 4971 278
rect 232 210 252 226
rect 4886 210 4906 226
rect 232 140 240 210
rect 4890 140 4906 210
rect 232 126 252 140
rect 4886 126 4906 140
rect 30 30 100 100
rect 5040 30 5110 100
<< via2 >>
rect 240 6310 252 6380
rect 252 6310 4886 6380
rect 4886 6310 4900 6380
rect 165 885 231 2645
rect 323 3885 389 5645
rect 481 885 547 2645
rect 639 3885 705 5645
rect 797 885 863 2645
rect 955 3885 1021 5645
rect 1113 885 1179 2645
rect 1271 3885 1337 5645
rect 1429 885 1495 2645
rect 1587 3885 1653 5645
rect 1745 885 1811 2645
rect 1903 3885 1969 5645
rect 2061 885 2127 2645
rect 2219 3885 2285 5645
rect 2377 885 2443 2645
rect 2535 3885 2601 5645
rect 2693 885 2759 2645
rect 2851 3885 2917 5645
rect 3009 885 3075 2645
rect 3167 3885 3233 5645
rect 3325 885 3391 2645
rect 3483 3885 3549 5645
rect 3641 885 3707 2645
rect 3799 3885 3865 5645
rect 3957 885 4023 2645
rect 4115 3885 4181 5645
rect 4273 885 4339 2645
rect 4431 3885 4497 5645
rect 4589 885 4655 2645
rect 4747 3885 4813 5645
rect 4905 885 4971 2645
rect 240 140 252 210
rect 252 140 4886 210
rect 4886 140 4890 210
<< metal3 >>
rect 100 6380 5100 6500
rect 100 6310 240 6380
rect 4900 6310 5100 6380
rect 100 6300 5100 6310
rect 30 5645 5110 5800
rect 30 3885 323 5645
rect 389 3885 639 5645
rect 705 3885 955 5645
rect 1021 3885 1271 5645
rect 1337 3885 1587 5645
rect 1653 3885 1903 5645
rect 1969 3885 2219 5645
rect 2285 3885 2535 5645
rect 2601 3885 2851 5645
rect 2917 3885 3167 5645
rect 3233 3885 3483 5645
rect 3549 3885 3799 5645
rect 3865 3885 4115 5645
rect 4181 3885 4431 5645
rect 4497 3885 4747 5645
rect 4813 3885 5110 5645
rect 30 3800 5110 3885
rect 30 2645 5110 2800
rect 30 885 165 2645
rect 231 885 481 2645
rect 547 885 797 2645
rect 863 885 1113 2645
rect 1179 885 1429 2645
rect 1495 885 1745 2645
rect 1811 885 2061 2645
rect 2127 885 2377 2645
rect 2443 885 2693 2645
rect 2759 885 3009 2645
rect 3075 885 3325 2645
rect 3391 885 3641 2645
rect 3707 885 3957 2645
rect 4023 885 4273 2645
rect 4339 885 4589 2645
rect 4655 885 4905 2645
rect 4971 885 5110 2645
rect 30 800 5110 885
rect 100 210 5100 230
rect 100 140 240 210
rect 4890 140 5100 210
rect 100 30 5100 140
<< labels >>
rlabel metal2 30 6420 100 6480 1 SUB
rlabel metal3 140 6300 200 6500 1 G
rlabel metal3 220 3810 260 5770 1 SD1
rlabel metal3 190 810 230 2770 1 SD2
<< end >>
