magic
tech sky130B
timestamp 1662171338
<< metal1 >>
rect 7000 60950 29000 61000
rect 7000 60940 7060 60950
rect 7190 60940 7310 60950
rect 7440 60940 7560 60950
rect 7690 60940 7810 60950
rect 7940 60940 8060 60950
rect 8190 60940 8310 60950
rect 8440 60940 8560 60950
rect 8690 60940 8810 60950
rect 8940 60940 9060 60950
rect 9190 60940 9310 60950
rect 9440 60940 9560 60950
rect 9690 60940 9810 60950
rect 9940 60940 10060 60950
rect 10190 60940 10310 60950
rect 10440 60940 10560 60950
rect 10690 60940 10810 60950
rect 10940 60940 11060 60950
rect 11190 60940 11310 60950
rect 11440 60940 11560 60950
rect 11690 60940 11810 60950
rect 11940 60940 12060 60950
rect 12190 60940 12310 60950
rect 12440 60940 12560 60950
rect 12690 60940 12810 60950
rect 12940 60940 13060 60950
rect 13190 60940 13310 60950
rect 13440 60940 13560 60950
rect 13690 60940 13810 60950
rect 13940 60940 14060 60950
rect 14190 60940 14310 60950
rect 14440 60940 14560 60950
rect 14690 60940 14810 60950
rect 14940 60940 15060 60950
rect 15190 60940 15310 60950
rect 15440 60940 15560 60950
rect 15690 60940 15810 60950
rect 15940 60940 16060 60950
rect 16190 60940 16310 60950
rect 16440 60940 16560 60950
rect 16690 60940 16810 60950
rect 16940 60940 17060 60950
rect 17190 60940 17310 60950
rect 17440 60940 17560 60950
rect 17690 60940 17810 60950
rect 17940 60940 18060 60950
rect 18190 60940 18310 60950
rect 18440 60940 18560 60950
rect 18690 60940 18810 60950
rect 18940 60940 19060 60950
rect 19190 60940 19310 60950
rect 19440 60940 19560 60950
rect 19690 60940 19810 60950
rect 19940 60940 20060 60950
rect 20190 60940 20310 60950
rect 20440 60940 20560 60950
rect 20690 60940 20810 60950
rect 20940 60940 21060 60950
rect 21190 60940 21310 60950
rect 21440 60940 21560 60950
rect 21690 60940 21810 60950
rect 21940 60940 22060 60950
rect 22190 60940 22310 60950
rect 22440 60940 22560 60950
rect 22690 60940 22810 60950
rect 22940 60940 23060 60950
rect 23190 60940 23310 60950
rect 23440 60940 23560 60950
rect 23690 60940 23810 60950
rect 23940 60940 24060 60950
rect 24190 60940 24310 60950
rect 24440 60940 24560 60950
rect 24690 60940 24810 60950
rect 24940 60940 25060 60950
rect 25190 60940 25310 60950
rect 25440 60940 25560 60950
rect 25690 60940 25810 60950
rect 25940 60940 26060 60950
rect 26190 60940 26310 60950
rect 26440 60940 26560 60950
rect 26690 60940 26810 60950
rect 26940 60940 27060 60950
rect 27190 60940 27310 60950
rect 27440 60940 27560 60950
rect 27690 60940 27810 60950
rect 27940 60940 28060 60950
rect 28190 60940 28310 60950
rect 28440 60940 28560 60950
rect 28690 60940 28810 60950
rect 28940 60940 29000 60950
rect 7000 60810 7050 60940
rect 7200 60810 7300 60940
rect 7450 60810 7550 60940
rect 7700 60810 7800 60940
rect 7950 60810 8050 60940
rect 8200 60810 8300 60940
rect 8450 60810 8550 60940
rect 8700 60810 8800 60940
rect 8950 60810 9050 60940
rect 9200 60810 9300 60940
rect 9450 60810 9550 60940
rect 9700 60810 9800 60940
rect 9950 60810 10050 60940
rect 10200 60810 10300 60940
rect 10450 60810 10550 60940
rect 10700 60810 10800 60940
rect 10950 60810 11050 60940
rect 11200 60810 11300 60940
rect 11450 60810 11550 60940
rect 11700 60810 11800 60940
rect 11950 60810 12050 60940
rect 12200 60810 12300 60940
rect 12450 60810 12550 60940
rect 12700 60810 12800 60940
rect 12950 60810 13050 60940
rect 13200 60810 13300 60940
rect 13450 60810 13550 60940
rect 13700 60810 13800 60940
rect 13950 60810 14050 60940
rect 14200 60810 14300 60940
rect 14450 60810 14550 60940
rect 14700 60810 14800 60940
rect 14950 60810 15050 60940
rect 15200 60810 15300 60940
rect 15450 60810 15550 60940
rect 15700 60810 15800 60940
rect 15950 60810 16050 60940
rect 16200 60810 16300 60940
rect 16450 60810 16550 60940
rect 16700 60810 16800 60940
rect 16950 60810 17050 60940
rect 17200 60810 17300 60940
rect 17450 60810 17550 60940
rect 17700 60810 17800 60940
rect 17950 60810 18050 60940
rect 18200 60810 18300 60940
rect 18450 60810 18550 60940
rect 18700 60810 18800 60940
rect 18950 60810 19050 60940
rect 19200 60810 19300 60940
rect 19450 60810 19550 60940
rect 19700 60810 19800 60940
rect 19950 60810 20050 60940
rect 20200 60810 20300 60940
rect 20450 60810 20550 60940
rect 20700 60810 20800 60940
rect 20950 60810 21050 60940
rect 21200 60810 21300 60940
rect 21450 60810 21550 60940
rect 21700 60810 21800 60940
rect 21950 60810 22050 60940
rect 22200 60810 22300 60940
rect 22450 60810 22550 60940
rect 22700 60810 22800 60940
rect 22950 60810 23050 60940
rect 23200 60810 23300 60940
rect 23450 60810 23550 60940
rect 23700 60810 23800 60940
rect 23950 60810 24050 60940
rect 24200 60810 24300 60940
rect 24450 60810 24550 60940
rect 24700 60810 24800 60940
rect 24950 60810 25050 60940
rect 25200 60810 25300 60940
rect 25450 60810 25550 60940
rect 25700 60810 25800 60940
rect 25950 60810 26050 60940
rect 26200 60810 26300 60940
rect 26450 60810 26550 60940
rect 26700 60810 26800 60940
rect 26950 60810 27050 60940
rect 27200 60810 27300 60940
rect 27450 60810 27550 60940
rect 27700 60810 27800 60940
rect 27950 60810 28050 60940
rect 28200 60810 28300 60940
rect 28450 60810 28550 60940
rect 28700 60810 28800 60940
rect 28950 60810 29000 60940
rect 7000 60800 7060 60810
rect 7190 60800 7310 60810
rect 7440 60800 7560 60810
rect 7690 60800 7810 60810
rect 7940 60800 8060 60810
rect 8190 60800 8310 60810
rect 8440 60800 8560 60810
rect 8690 60800 8810 60810
rect 8940 60800 9060 60810
rect 9190 60800 9310 60810
rect 9440 60800 9560 60810
rect 9690 60800 9810 60810
rect 9940 60800 10060 60810
rect 10190 60800 10310 60810
rect 10440 60800 10560 60810
rect 10690 60800 10810 60810
rect 10940 60800 11060 60810
rect 11190 60800 11310 60810
rect 11440 60800 11560 60810
rect 11690 60800 11810 60810
rect 11940 60800 12060 60810
rect 12190 60800 12310 60810
rect 12440 60800 12560 60810
rect 12690 60800 12810 60810
rect 12940 60800 13060 60810
rect 13190 60800 13310 60810
rect 13440 60800 13560 60810
rect 13690 60800 13810 60810
rect 13940 60800 14060 60810
rect 14190 60800 14310 60810
rect 14440 60800 14560 60810
rect 14690 60800 14810 60810
rect 14940 60800 15060 60810
rect 15190 60800 15310 60810
rect 15440 60800 15560 60810
rect 15690 60800 15810 60810
rect 15940 60800 16060 60810
rect 16190 60800 16310 60810
rect 16440 60800 16560 60810
rect 16690 60800 16810 60810
rect 16940 60800 17060 60810
rect 17190 60800 17310 60810
rect 17440 60800 17560 60810
rect 17690 60800 17810 60810
rect 17940 60800 18060 60810
rect 18190 60800 18310 60810
rect 18440 60800 18560 60810
rect 18690 60800 18810 60810
rect 18940 60800 19060 60810
rect 19190 60800 19310 60810
rect 19440 60800 19560 60810
rect 19690 60800 19810 60810
rect 19940 60800 20060 60810
rect 20190 60800 20310 60810
rect 20440 60800 20560 60810
rect 20690 60800 20810 60810
rect 20940 60800 21060 60810
rect 21190 60800 21310 60810
rect 21440 60800 21560 60810
rect 21690 60800 21810 60810
rect 21940 60800 22060 60810
rect 22190 60800 22310 60810
rect 22440 60800 22560 60810
rect 22690 60800 22810 60810
rect 22940 60800 23060 60810
rect 23190 60800 23310 60810
rect 23440 60800 23560 60810
rect 23690 60800 23810 60810
rect 23940 60800 24060 60810
rect 24190 60800 24310 60810
rect 24440 60800 24560 60810
rect 24690 60800 24810 60810
rect 24940 60800 25060 60810
rect 25190 60800 25310 60810
rect 25440 60800 25560 60810
rect 25690 60800 25810 60810
rect 25940 60800 26060 60810
rect 26190 60800 26310 60810
rect 26440 60800 26560 60810
rect 26690 60800 26810 60810
rect 26940 60800 27060 60810
rect 27190 60800 27310 60810
rect 27440 60800 27560 60810
rect 27690 60800 27810 60810
rect 27940 60800 28060 60810
rect 28190 60800 28310 60810
rect 28440 60800 28560 60810
rect 28690 60800 28810 60810
rect 28940 60800 29000 60810
rect 7000 60700 29000 60800
rect 7000 60690 7060 60700
rect 7190 60690 7310 60700
rect 7440 60690 7560 60700
rect 7690 60690 7810 60700
rect 7940 60690 8060 60700
rect 8190 60690 8310 60700
rect 8440 60690 8560 60700
rect 8690 60690 8810 60700
rect 8940 60690 9060 60700
rect 9190 60690 9310 60700
rect 9440 60690 9560 60700
rect 9690 60690 9810 60700
rect 9940 60690 10060 60700
rect 10190 60690 10310 60700
rect 10440 60690 10560 60700
rect 10690 60690 10810 60700
rect 10940 60690 11060 60700
rect 11190 60690 11310 60700
rect 11440 60690 11560 60700
rect 11690 60690 11810 60700
rect 11940 60690 12060 60700
rect 12190 60690 12310 60700
rect 12440 60690 12560 60700
rect 12690 60690 12810 60700
rect 12940 60690 13060 60700
rect 13190 60690 13310 60700
rect 13440 60690 13560 60700
rect 13690 60690 13810 60700
rect 13940 60690 14060 60700
rect 14190 60690 14310 60700
rect 14440 60690 14560 60700
rect 14690 60690 14810 60700
rect 14940 60690 15060 60700
rect 15190 60690 15310 60700
rect 15440 60690 15560 60700
rect 15690 60690 15810 60700
rect 15940 60690 16060 60700
rect 16190 60690 16310 60700
rect 16440 60690 16560 60700
rect 16690 60690 16810 60700
rect 16940 60690 17060 60700
rect 17190 60690 17310 60700
rect 17440 60690 17560 60700
rect 17690 60690 17810 60700
rect 17940 60690 18060 60700
rect 18190 60690 18310 60700
rect 18440 60690 18560 60700
rect 18690 60690 18810 60700
rect 18940 60690 19060 60700
rect 19190 60690 19310 60700
rect 19440 60690 19560 60700
rect 19690 60690 19810 60700
rect 19940 60690 20060 60700
rect 20190 60690 20310 60700
rect 20440 60690 20560 60700
rect 20690 60690 20810 60700
rect 20940 60690 21060 60700
rect 21190 60690 21310 60700
rect 21440 60690 21560 60700
rect 21690 60690 21810 60700
rect 21940 60690 22060 60700
rect 22190 60690 22310 60700
rect 22440 60690 22560 60700
rect 22690 60690 22810 60700
rect 22940 60690 23060 60700
rect 23190 60690 23310 60700
rect 23440 60690 23560 60700
rect 23690 60690 23810 60700
rect 23940 60690 24060 60700
rect 24190 60690 24310 60700
rect 24440 60690 24560 60700
rect 24690 60690 24810 60700
rect 24940 60690 25060 60700
rect 25190 60690 25310 60700
rect 25440 60690 25560 60700
rect 25690 60690 25810 60700
rect 25940 60690 26060 60700
rect 26190 60690 26310 60700
rect 26440 60690 26560 60700
rect 26690 60690 26810 60700
rect 26940 60690 27060 60700
rect 27190 60690 27310 60700
rect 27440 60690 27560 60700
rect 27690 60690 27810 60700
rect 27940 60690 28060 60700
rect 28190 60690 28310 60700
rect 28440 60690 28560 60700
rect 28690 60690 28810 60700
rect 28940 60690 29000 60700
rect 7000 60560 7050 60690
rect 7200 60560 7300 60690
rect 7450 60560 7550 60690
rect 7700 60560 7800 60690
rect 7950 60560 8050 60690
rect 8200 60560 8300 60690
rect 8450 60560 8550 60690
rect 8700 60560 8800 60690
rect 8950 60560 9050 60690
rect 9200 60560 9300 60690
rect 9450 60560 9550 60690
rect 9700 60560 9800 60690
rect 9950 60560 10050 60690
rect 10200 60560 10300 60690
rect 10450 60560 10550 60690
rect 10700 60560 10800 60690
rect 10950 60560 11050 60690
rect 11200 60560 11300 60690
rect 11450 60560 11550 60690
rect 11700 60560 11800 60690
rect 11950 60560 12050 60690
rect 12200 60560 12300 60690
rect 12450 60560 12550 60690
rect 12700 60560 12800 60690
rect 12950 60560 13050 60690
rect 13200 60560 13300 60690
rect 13450 60560 13550 60690
rect 13700 60560 13800 60690
rect 13950 60560 14050 60690
rect 14200 60560 14300 60690
rect 14450 60560 14550 60690
rect 14700 60560 14800 60690
rect 14950 60560 15050 60690
rect 15200 60560 15300 60690
rect 15450 60560 15550 60690
rect 15700 60560 15800 60690
rect 15950 60560 16050 60690
rect 16200 60560 16300 60690
rect 16450 60560 16550 60690
rect 16700 60560 16800 60690
rect 16950 60560 17050 60690
rect 17200 60560 17300 60690
rect 17450 60560 17550 60690
rect 17700 60560 17800 60690
rect 17950 60560 18050 60690
rect 18200 60560 18300 60690
rect 18450 60560 18550 60690
rect 18700 60560 18800 60690
rect 18950 60560 19050 60690
rect 19200 60560 19300 60690
rect 19450 60560 19550 60690
rect 19700 60560 19800 60690
rect 19950 60560 20050 60690
rect 20200 60560 20300 60690
rect 20450 60560 20550 60690
rect 20700 60560 20800 60690
rect 20950 60560 21050 60690
rect 21200 60560 21300 60690
rect 21450 60560 21550 60690
rect 21700 60560 21800 60690
rect 21950 60560 22050 60690
rect 22200 60560 22300 60690
rect 22450 60560 22550 60690
rect 22700 60560 22800 60690
rect 22950 60560 23050 60690
rect 23200 60560 23300 60690
rect 23450 60560 23550 60690
rect 23700 60560 23800 60690
rect 23950 60560 24050 60690
rect 24200 60560 24300 60690
rect 24450 60560 24550 60690
rect 24700 60560 24800 60690
rect 24950 60560 25050 60690
rect 25200 60560 25300 60690
rect 25450 60560 25550 60690
rect 25700 60560 25800 60690
rect 25950 60560 26050 60690
rect 26200 60560 26300 60690
rect 26450 60560 26550 60690
rect 26700 60560 26800 60690
rect 26950 60560 27050 60690
rect 27200 60560 27300 60690
rect 27450 60560 27550 60690
rect 27700 60560 27800 60690
rect 27950 60560 28050 60690
rect 28200 60560 28300 60690
rect 28450 60560 28550 60690
rect 28700 60560 28800 60690
rect 28950 60560 29000 60690
rect 7000 60550 7060 60560
rect 7190 60550 7310 60560
rect 7440 60550 7560 60560
rect 7690 60550 7810 60560
rect 7940 60550 8060 60560
rect 8190 60550 8310 60560
rect 8440 60550 8560 60560
rect 8690 60550 8810 60560
rect 8940 60550 9060 60560
rect 9190 60550 9310 60560
rect 9440 60550 9560 60560
rect 9690 60550 9810 60560
rect 9940 60550 10060 60560
rect 10190 60550 10310 60560
rect 10440 60550 10560 60560
rect 10690 60550 10810 60560
rect 10940 60550 11060 60560
rect 11190 60550 11310 60560
rect 11440 60550 11560 60560
rect 11690 60550 11810 60560
rect 11940 60550 12060 60560
rect 12190 60550 12310 60560
rect 12440 60550 12560 60560
rect 12690 60550 12810 60560
rect 12940 60550 13060 60560
rect 13190 60550 13310 60560
rect 13440 60550 13560 60560
rect 13690 60550 13810 60560
rect 13940 60550 14060 60560
rect 14190 60550 14310 60560
rect 14440 60550 14560 60560
rect 14690 60550 14810 60560
rect 14940 60550 15060 60560
rect 15190 60550 15310 60560
rect 15440 60550 15560 60560
rect 15690 60550 15810 60560
rect 15940 60550 16060 60560
rect 16190 60550 16310 60560
rect 16440 60550 16560 60560
rect 16690 60550 16810 60560
rect 16940 60550 17060 60560
rect 17190 60550 17310 60560
rect 17440 60550 17560 60560
rect 17690 60550 17810 60560
rect 17940 60550 18060 60560
rect 18190 60550 18310 60560
rect 18440 60550 18560 60560
rect 18690 60550 18810 60560
rect 18940 60550 19060 60560
rect 19190 60550 19310 60560
rect 19440 60550 19560 60560
rect 19690 60550 19810 60560
rect 19940 60550 20060 60560
rect 20190 60550 20310 60560
rect 20440 60550 20560 60560
rect 20690 60550 20810 60560
rect 20940 60550 21060 60560
rect 21190 60550 21310 60560
rect 21440 60550 21560 60560
rect 21690 60550 21810 60560
rect 21940 60550 22060 60560
rect 22190 60550 22310 60560
rect 22440 60550 22560 60560
rect 22690 60550 22810 60560
rect 22940 60550 23060 60560
rect 23190 60550 23310 60560
rect 23440 60550 23560 60560
rect 23690 60550 23810 60560
rect 23940 60550 24060 60560
rect 24190 60550 24310 60560
rect 24440 60550 24560 60560
rect 24690 60550 24810 60560
rect 24940 60550 25060 60560
rect 25190 60550 25310 60560
rect 25440 60550 25560 60560
rect 25690 60550 25810 60560
rect 25940 60550 26060 60560
rect 26190 60550 26310 60560
rect 26440 60550 26560 60560
rect 26690 60550 26810 60560
rect 26940 60550 27060 60560
rect 27190 60550 27310 60560
rect 27440 60550 27560 60560
rect 27690 60550 27810 60560
rect 27940 60550 28060 60560
rect 28190 60550 28310 60560
rect 28440 60550 28560 60560
rect 28690 60550 28810 60560
rect 28940 60550 29000 60560
rect 7000 60450 29000 60550
rect 7000 60440 7060 60450
rect 7190 60440 7310 60450
rect 7440 60440 7560 60450
rect 7690 60440 7810 60450
rect 7940 60440 8060 60450
rect 8190 60440 8310 60450
rect 8440 60440 8560 60450
rect 8690 60440 8810 60450
rect 8940 60440 9060 60450
rect 9190 60440 9310 60450
rect 9440 60440 9560 60450
rect 9690 60440 9810 60450
rect 9940 60440 10060 60450
rect 10190 60440 10310 60450
rect 10440 60440 10560 60450
rect 10690 60440 10810 60450
rect 10940 60440 11060 60450
rect 11190 60440 11310 60450
rect 11440 60440 11560 60450
rect 11690 60440 11810 60450
rect 11940 60440 12060 60450
rect 12190 60440 12310 60450
rect 12440 60440 12560 60450
rect 12690 60440 12810 60450
rect 12940 60440 13060 60450
rect 13190 60440 13310 60450
rect 13440 60440 13560 60450
rect 13690 60440 13810 60450
rect 13940 60440 14060 60450
rect 14190 60440 14310 60450
rect 14440 60440 14560 60450
rect 14690 60440 14810 60450
rect 14940 60440 15060 60450
rect 15190 60440 15310 60450
rect 15440 60440 15560 60450
rect 15690 60440 15810 60450
rect 15940 60440 16060 60450
rect 16190 60440 16310 60450
rect 16440 60440 16560 60450
rect 16690 60440 16810 60450
rect 16940 60440 17060 60450
rect 17190 60440 17310 60450
rect 17440 60440 17560 60450
rect 17690 60440 17810 60450
rect 17940 60440 18060 60450
rect 18190 60440 18310 60450
rect 18440 60440 18560 60450
rect 18690 60440 18810 60450
rect 18940 60440 19060 60450
rect 19190 60440 19310 60450
rect 19440 60440 19560 60450
rect 19690 60440 19810 60450
rect 19940 60440 20060 60450
rect 20190 60440 20310 60450
rect 20440 60440 20560 60450
rect 20690 60440 20810 60450
rect 20940 60440 21060 60450
rect 21190 60440 21310 60450
rect 21440 60440 21560 60450
rect 21690 60440 21810 60450
rect 21940 60440 22060 60450
rect 22190 60440 22310 60450
rect 22440 60440 22560 60450
rect 22690 60440 22810 60450
rect 22940 60440 23060 60450
rect 23190 60440 23310 60450
rect 23440 60440 23560 60450
rect 23690 60440 23810 60450
rect 23940 60440 24060 60450
rect 24190 60440 24310 60450
rect 24440 60440 24560 60450
rect 24690 60440 24810 60450
rect 24940 60440 25060 60450
rect 25190 60440 25310 60450
rect 25440 60440 25560 60450
rect 25690 60440 25810 60450
rect 25940 60440 26060 60450
rect 26190 60440 26310 60450
rect 26440 60440 26560 60450
rect 26690 60440 26810 60450
rect 26940 60440 27060 60450
rect 27190 60440 27310 60450
rect 27440 60440 27560 60450
rect 27690 60440 27810 60450
rect 27940 60440 28060 60450
rect 28190 60440 28310 60450
rect 28440 60440 28560 60450
rect 28690 60440 28810 60450
rect 28940 60440 29000 60450
rect 7000 60310 7050 60440
rect 7200 60310 7300 60440
rect 7450 60310 7550 60440
rect 7700 60310 7800 60440
rect 7950 60310 8050 60440
rect 8200 60310 8300 60440
rect 8450 60310 8550 60440
rect 8700 60310 8800 60440
rect 8950 60310 9050 60440
rect 9200 60310 9300 60440
rect 9450 60310 9550 60440
rect 9700 60310 9800 60440
rect 9950 60310 10050 60440
rect 10200 60310 10300 60440
rect 10450 60310 10550 60440
rect 10700 60310 10800 60440
rect 10950 60310 11050 60440
rect 11200 60310 11300 60440
rect 11450 60310 11550 60440
rect 11700 60310 11800 60440
rect 11950 60310 12050 60440
rect 12200 60310 12300 60440
rect 12450 60310 12550 60440
rect 12700 60310 12800 60440
rect 12950 60310 13050 60440
rect 13200 60310 13300 60440
rect 13450 60310 13550 60440
rect 13700 60310 13800 60440
rect 13950 60310 14050 60440
rect 14200 60310 14300 60440
rect 14450 60310 14550 60440
rect 14700 60310 14800 60440
rect 14950 60310 15050 60440
rect 15200 60310 15300 60440
rect 15450 60310 15550 60440
rect 15700 60310 15800 60440
rect 15950 60310 16050 60440
rect 16200 60310 16300 60440
rect 16450 60310 16550 60440
rect 16700 60310 16800 60440
rect 16950 60310 17050 60440
rect 17200 60310 17300 60440
rect 17450 60310 17550 60440
rect 17700 60310 17800 60440
rect 17950 60310 18050 60440
rect 18200 60310 18300 60440
rect 18450 60310 18550 60440
rect 18700 60310 18800 60440
rect 18950 60310 19050 60440
rect 19200 60310 19300 60440
rect 19450 60310 19550 60440
rect 19700 60310 19800 60440
rect 19950 60310 20050 60440
rect 20200 60310 20300 60440
rect 20450 60310 20550 60440
rect 20700 60310 20800 60440
rect 20950 60310 21050 60440
rect 21200 60310 21300 60440
rect 21450 60310 21550 60440
rect 21700 60310 21800 60440
rect 21950 60310 22050 60440
rect 22200 60310 22300 60440
rect 22450 60310 22550 60440
rect 22700 60310 22800 60440
rect 22950 60310 23050 60440
rect 23200 60310 23300 60440
rect 23450 60310 23550 60440
rect 23700 60310 23800 60440
rect 23950 60310 24050 60440
rect 24200 60310 24300 60440
rect 24450 60310 24550 60440
rect 24700 60310 24800 60440
rect 24950 60310 25050 60440
rect 25200 60310 25300 60440
rect 25450 60310 25550 60440
rect 25700 60310 25800 60440
rect 25950 60310 26050 60440
rect 26200 60310 26300 60440
rect 26450 60310 26550 60440
rect 26700 60310 26800 60440
rect 26950 60310 27050 60440
rect 27200 60310 27300 60440
rect 27450 60310 27550 60440
rect 27700 60310 27800 60440
rect 27950 60310 28050 60440
rect 28200 60310 28300 60440
rect 28450 60310 28550 60440
rect 28700 60310 28800 60440
rect 28950 60310 29000 60440
rect 7000 60300 7060 60310
rect 7190 60300 7310 60310
rect 7440 60300 7560 60310
rect 7690 60300 7810 60310
rect 7940 60300 8060 60310
rect 8190 60300 8310 60310
rect 8440 60300 8560 60310
rect 8690 60300 8810 60310
rect 8940 60300 9060 60310
rect 9190 60300 9310 60310
rect 9440 60300 9560 60310
rect 9690 60300 9810 60310
rect 9940 60300 10060 60310
rect 10190 60300 10310 60310
rect 10440 60300 10560 60310
rect 10690 60300 10810 60310
rect 10940 60300 11060 60310
rect 11190 60300 11310 60310
rect 11440 60300 11560 60310
rect 11690 60300 11810 60310
rect 11940 60300 12060 60310
rect 12190 60300 12310 60310
rect 12440 60300 12560 60310
rect 12690 60300 12810 60310
rect 12940 60300 13060 60310
rect 13190 60300 13310 60310
rect 13440 60300 13560 60310
rect 13690 60300 13810 60310
rect 13940 60300 14060 60310
rect 14190 60300 14310 60310
rect 14440 60300 14560 60310
rect 14690 60300 14810 60310
rect 14940 60300 15060 60310
rect 15190 60300 15310 60310
rect 15440 60300 15560 60310
rect 15690 60300 15810 60310
rect 15940 60300 16060 60310
rect 16190 60300 16310 60310
rect 16440 60300 16560 60310
rect 16690 60300 16810 60310
rect 16940 60300 17060 60310
rect 17190 60300 17310 60310
rect 17440 60300 17560 60310
rect 17690 60300 17810 60310
rect 17940 60300 18060 60310
rect 18190 60300 18310 60310
rect 18440 60300 18560 60310
rect 18690 60300 18810 60310
rect 18940 60300 19060 60310
rect 19190 60300 19310 60310
rect 19440 60300 19560 60310
rect 19690 60300 19810 60310
rect 19940 60300 20060 60310
rect 20190 60300 20310 60310
rect 20440 60300 20560 60310
rect 20690 60300 20810 60310
rect 20940 60300 21060 60310
rect 21190 60300 21310 60310
rect 21440 60300 21560 60310
rect 21690 60300 21810 60310
rect 21940 60300 22060 60310
rect 22190 60300 22310 60310
rect 22440 60300 22560 60310
rect 22690 60300 22810 60310
rect 22940 60300 23060 60310
rect 23190 60300 23310 60310
rect 23440 60300 23560 60310
rect 23690 60300 23810 60310
rect 23940 60300 24060 60310
rect 24190 60300 24310 60310
rect 24440 60300 24560 60310
rect 24690 60300 24810 60310
rect 24940 60300 25060 60310
rect 25190 60300 25310 60310
rect 25440 60300 25560 60310
rect 25690 60300 25810 60310
rect 25940 60300 26060 60310
rect 26190 60300 26310 60310
rect 26440 60300 26560 60310
rect 26690 60300 26810 60310
rect 26940 60300 27060 60310
rect 27190 60300 27310 60310
rect 27440 60300 27560 60310
rect 27690 60300 27810 60310
rect 27940 60300 28060 60310
rect 28190 60300 28310 60310
rect 28440 60300 28560 60310
rect 28690 60300 28810 60310
rect 28940 60300 29000 60310
rect 7000 60200 29000 60300
rect 7000 60190 7060 60200
rect 7190 60190 7310 60200
rect 7440 60190 7560 60200
rect 7690 60190 7810 60200
rect 7940 60190 8060 60200
rect 8190 60190 8310 60200
rect 8440 60190 8560 60200
rect 8690 60190 8810 60200
rect 8940 60190 9060 60200
rect 9190 60190 9310 60200
rect 9440 60190 9560 60200
rect 9690 60190 9810 60200
rect 9940 60190 10060 60200
rect 10190 60190 10310 60200
rect 10440 60190 10560 60200
rect 10690 60190 10810 60200
rect 10940 60190 11060 60200
rect 11190 60190 11310 60200
rect 11440 60190 11560 60200
rect 11690 60190 11810 60200
rect 11940 60190 12060 60200
rect 12190 60190 12310 60200
rect 12440 60190 12560 60200
rect 12690 60190 12810 60200
rect 12940 60190 13060 60200
rect 13190 60190 13310 60200
rect 13440 60190 13560 60200
rect 13690 60190 13810 60200
rect 13940 60190 14060 60200
rect 14190 60190 14310 60200
rect 14440 60190 14560 60200
rect 14690 60190 14810 60200
rect 14940 60190 15060 60200
rect 15190 60190 15310 60200
rect 15440 60190 15560 60200
rect 15690 60190 15810 60200
rect 15940 60190 16060 60200
rect 16190 60190 16310 60200
rect 16440 60190 16560 60200
rect 16690 60190 16810 60200
rect 16940 60190 17060 60200
rect 17190 60190 17310 60200
rect 17440 60190 17560 60200
rect 17690 60190 17810 60200
rect 17940 60190 18060 60200
rect 18190 60190 18310 60200
rect 18440 60190 18560 60200
rect 18690 60190 18810 60200
rect 18940 60190 19060 60200
rect 19190 60190 19310 60200
rect 19440 60190 19560 60200
rect 19690 60190 19810 60200
rect 19940 60190 20060 60200
rect 20190 60190 20310 60200
rect 20440 60190 20560 60200
rect 20690 60190 20810 60200
rect 20940 60190 21060 60200
rect 21190 60190 21310 60200
rect 21440 60190 21560 60200
rect 21690 60190 21810 60200
rect 21940 60190 22060 60200
rect 22190 60190 22310 60200
rect 22440 60190 22560 60200
rect 22690 60190 22810 60200
rect 22940 60190 23060 60200
rect 23190 60190 23310 60200
rect 23440 60190 23560 60200
rect 23690 60190 23810 60200
rect 23940 60190 24060 60200
rect 24190 60190 24310 60200
rect 24440 60190 24560 60200
rect 24690 60190 24810 60200
rect 24940 60190 25060 60200
rect 25190 60190 25310 60200
rect 25440 60190 25560 60200
rect 25690 60190 25810 60200
rect 25940 60190 26060 60200
rect 26190 60190 26310 60200
rect 26440 60190 26560 60200
rect 26690 60190 26810 60200
rect 26940 60190 27060 60200
rect 27190 60190 27310 60200
rect 27440 60190 27560 60200
rect 27690 60190 27810 60200
rect 27940 60190 28060 60200
rect 28190 60190 28310 60200
rect 28440 60190 28560 60200
rect 28690 60190 28810 60200
rect 28940 60190 29000 60200
rect 7000 60060 7050 60190
rect 7200 60060 7300 60190
rect 7450 60060 7550 60190
rect 7700 60060 7800 60190
rect 7950 60060 8050 60190
rect 8200 60060 8300 60190
rect 8450 60060 8550 60190
rect 8700 60060 8800 60190
rect 8950 60060 9050 60190
rect 9200 60060 9300 60190
rect 9450 60060 9550 60190
rect 9700 60060 9800 60190
rect 9950 60060 10050 60190
rect 10200 60060 10300 60190
rect 10450 60060 10550 60190
rect 10700 60060 10800 60190
rect 10950 60060 11050 60190
rect 11200 60060 11300 60190
rect 11450 60060 11550 60190
rect 11700 60060 11800 60190
rect 11950 60060 12050 60190
rect 12200 60060 12300 60190
rect 12450 60060 12550 60190
rect 12700 60060 12800 60190
rect 12950 60060 13050 60190
rect 13200 60060 13300 60190
rect 13450 60060 13550 60190
rect 13700 60060 13800 60190
rect 13950 60060 14050 60190
rect 14200 60060 14300 60190
rect 14450 60060 14550 60190
rect 14700 60060 14800 60190
rect 14950 60060 15050 60190
rect 15200 60060 15300 60190
rect 15450 60060 15550 60190
rect 15700 60060 15800 60190
rect 15950 60060 16050 60190
rect 16200 60060 16300 60190
rect 16450 60060 16550 60190
rect 16700 60060 16800 60190
rect 16950 60060 17050 60190
rect 17200 60060 17300 60190
rect 17450 60060 17550 60190
rect 17700 60060 17800 60190
rect 17950 60060 18050 60190
rect 18200 60060 18300 60190
rect 18450 60060 18550 60190
rect 18700 60060 18800 60190
rect 18950 60060 19050 60190
rect 19200 60060 19300 60190
rect 19450 60060 19550 60190
rect 19700 60060 19800 60190
rect 19950 60060 20050 60190
rect 20200 60060 20300 60190
rect 20450 60060 20550 60190
rect 20700 60060 20800 60190
rect 20950 60060 21050 60190
rect 21200 60060 21300 60190
rect 21450 60060 21550 60190
rect 21700 60060 21800 60190
rect 21950 60060 22050 60190
rect 22200 60060 22300 60190
rect 22450 60060 22550 60190
rect 22700 60060 22800 60190
rect 22950 60060 23050 60190
rect 23200 60060 23300 60190
rect 23450 60060 23550 60190
rect 23700 60060 23800 60190
rect 23950 60060 24050 60190
rect 24200 60060 24300 60190
rect 24450 60060 24550 60190
rect 24700 60060 24800 60190
rect 24950 60060 25050 60190
rect 25200 60060 25300 60190
rect 25450 60060 25550 60190
rect 25700 60060 25800 60190
rect 25950 60060 26050 60190
rect 26200 60060 26300 60190
rect 26450 60060 26550 60190
rect 26700 60060 26800 60190
rect 26950 60060 27050 60190
rect 27200 60060 27300 60190
rect 27450 60060 27550 60190
rect 27700 60060 27800 60190
rect 27950 60060 28050 60190
rect 28200 60060 28300 60190
rect 28450 60060 28550 60190
rect 28700 60060 28800 60190
rect 28950 60060 29000 60190
rect 7000 60050 7060 60060
rect 7190 60050 7310 60060
rect 7440 60050 7560 60060
rect 7690 60050 7810 60060
rect 7940 60050 8060 60060
rect 8190 60050 8310 60060
rect 8440 60050 8560 60060
rect 8690 60050 8810 60060
rect 8940 60050 9060 60060
rect 9190 60050 9310 60060
rect 9440 60050 9560 60060
rect 9690 60050 9810 60060
rect 9940 60050 10060 60060
rect 10190 60050 10310 60060
rect 10440 60050 10560 60060
rect 10690 60050 10810 60060
rect 10940 60050 11060 60060
rect 11190 60050 11310 60060
rect 11440 60050 11560 60060
rect 11690 60050 11810 60060
rect 11940 60050 12060 60060
rect 12190 60050 12310 60060
rect 12440 60050 12560 60060
rect 12690 60050 12810 60060
rect 12940 60050 13060 60060
rect 13190 60050 13310 60060
rect 13440 60050 13560 60060
rect 13690 60050 13810 60060
rect 13940 60050 14060 60060
rect 14190 60050 14310 60060
rect 14440 60050 14560 60060
rect 14690 60050 14810 60060
rect 14940 60050 15060 60060
rect 15190 60050 15310 60060
rect 15440 60050 15560 60060
rect 15690 60050 15810 60060
rect 15940 60050 16060 60060
rect 16190 60050 16310 60060
rect 16440 60050 16560 60060
rect 16690 60050 16810 60060
rect 16940 60050 17060 60060
rect 17190 60050 17310 60060
rect 17440 60050 17560 60060
rect 17690 60050 17810 60060
rect 17940 60050 18060 60060
rect 18190 60050 18310 60060
rect 18440 60050 18560 60060
rect 18690 60050 18810 60060
rect 18940 60050 19060 60060
rect 19190 60050 19310 60060
rect 19440 60050 19560 60060
rect 19690 60050 19810 60060
rect 19940 60050 20060 60060
rect 20190 60050 20310 60060
rect 20440 60050 20560 60060
rect 20690 60050 20810 60060
rect 20940 60050 21060 60060
rect 21190 60050 21310 60060
rect 21440 60050 21560 60060
rect 21690 60050 21810 60060
rect 21940 60050 22060 60060
rect 22190 60050 22310 60060
rect 22440 60050 22560 60060
rect 22690 60050 22810 60060
rect 22940 60050 23060 60060
rect 23190 60050 23310 60060
rect 23440 60050 23560 60060
rect 23690 60050 23810 60060
rect 23940 60050 24060 60060
rect 24190 60050 24310 60060
rect 24440 60050 24560 60060
rect 24690 60050 24810 60060
rect 24940 60050 25060 60060
rect 25190 60050 25310 60060
rect 25440 60050 25560 60060
rect 25690 60050 25810 60060
rect 25940 60050 26060 60060
rect 26190 60050 26310 60060
rect 26440 60050 26560 60060
rect 26690 60050 26810 60060
rect 26940 60050 27060 60060
rect 27190 60050 27310 60060
rect 27440 60050 27560 60060
rect 27690 60050 27810 60060
rect 27940 60050 28060 60060
rect 28190 60050 28310 60060
rect 28440 60050 28560 60060
rect 28690 60050 28810 60060
rect 28940 60050 29000 60060
rect 7000 59950 29000 60050
rect 7000 59940 7060 59950
rect 7190 59940 7310 59950
rect 7440 59940 7560 59950
rect 7690 59940 7810 59950
rect 7940 59940 8060 59950
rect 8190 59940 8310 59950
rect 8440 59940 8560 59950
rect 8690 59940 8810 59950
rect 8940 59940 9060 59950
rect 9190 59940 9310 59950
rect 9440 59940 9560 59950
rect 9690 59940 9810 59950
rect 9940 59940 10060 59950
rect 10190 59940 10310 59950
rect 10440 59940 10560 59950
rect 10690 59940 10810 59950
rect 10940 59940 11060 59950
rect 11190 59940 11310 59950
rect 11440 59940 11560 59950
rect 11690 59940 11810 59950
rect 11940 59940 12060 59950
rect 12190 59940 12310 59950
rect 12440 59940 12560 59950
rect 12690 59940 12810 59950
rect 12940 59940 13060 59950
rect 13190 59940 13310 59950
rect 13440 59940 13560 59950
rect 13690 59940 13810 59950
rect 13940 59940 14060 59950
rect 14190 59940 14310 59950
rect 14440 59940 14560 59950
rect 14690 59940 14810 59950
rect 14940 59940 15060 59950
rect 15190 59940 15310 59950
rect 15440 59940 15560 59950
rect 15690 59940 15810 59950
rect 15940 59940 16060 59950
rect 16190 59940 16310 59950
rect 16440 59940 16560 59950
rect 16690 59940 16810 59950
rect 16940 59940 17060 59950
rect 17190 59940 17310 59950
rect 17440 59940 17560 59950
rect 17690 59940 17810 59950
rect 17940 59940 18060 59950
rect 18190 59940 18310 59950
rect 18440 59940 18560 59950
rect 18690 59940 18810 59950
rect 18940 59940 19060 59950
rect 19190 59940 19310 59950
rect 19440 59940 19560 59950
rect 19690 59940 19810 59950
rect 19940 59940 20060 59950
rect 20190 59940 20310 59950
rect 20440 59940 20560 59950
rect 20690 59940 20810 59950
rect 20940 59940 21060 59950
rect 21190 59940 21310 59950
rect 21440 59940 21560 59950
rect 21690 59940 21810 59950
rect 21940 59940 22060 59950
rect 22190 59940 22310 59950
rect 22440 59940 22560 59950
rect 22690 59940 22810 59950
rect 22940 59940 23060 59950
rect 23190 59940 23310 59950
rect 23440 59940 23560 59950
rect 23690 59940 23810 59950
rect 23940 59940 24060 59950
rect 24190 59940 24310 59950
rect 24440 59940 24560 59950
rect 24690 59940 24810 59950
rect 24940 59940 25060 59950
rect 25190 59940 25310 59950
rect 25440 59940 25560 59950
rect 25690 59940 25810 59950
rect 25940 59940 26060 59950
rect 26190 59940 26310 59950
rect 26440 59940 26560 59950
rect 26690 59940 26810 59950
rect 26940 59940 27060 59950
rect 27190 59940 27310 59950
rect 27440 59940 27560 59950
rect 27690 59940 27810 59950
rect 27940 59940 28060 59950
rect 28190 59940 28310 59950
rect 28440 59940 28560 59950
rect 28690 59940 28810 59950
rect 28940 59940 29000 59950
rect 7000 59810 7050 59940
rect 7200 59810 7300 59940
rect 7450 59810 7550 59940
rect 7700 59810 7800 59940
rect 7950 59810 8050 59940
rect 8200 59810 8300 59940
rect 8450 59810 8550 59940
rect 8700 59810 8800 59940
rect 8950 59810 9050 59940
rect 9200 59810 9300 59940
rect 9450 59810 9550 59940
rect 9700 59810 9800 59940
rect 9950 59810 10050 59940
rect 10200 59810 10300 59940
rect 10450 59810 10550 59940
rect 10700 59810 10800 59940
rect 10950 59810 11050 59940
rect 11200 59810 11300 59940
rect 11450 59810 11550 59940
rect 11700 59810 11800 59940
rect 11950 59810 12050 59940
rect 12200 59810 12300 59940
rect 12450 59810 12550 59940
rect 12700 59810 12800 59940
rect 12950 59810 13050 59940
rect 13200 59810 13300 59940
rect 13450 59810 13550 59940
rect 13700 59810 13800 59940
rect 13950 59810 14050 59940
rect 14200 59810 14300 59940
rect 14450 59810 14550 59940
rect 14700 59810 14800 59940
rect 14950 59810 15050 59940
rect 15200 59810 15300 59940
rect 15450 59810 15550 59940
rect 15700 59810 15800 59940
rect 15950 59810 16050 59940
rect 16200 59810 16300 59940
rect 16450 59810 16550 59940
rect 16700 59810 16800 59940
rect 16950 59810 17050 59940
rect 17200 59810 17300 59940
rect 17450 59810 17550 59940
rect 17700 59810 17800 59940
rect 17950 59810 18050 59940
rect 18200 59810 18300 59940
rect 18450 59810 18550 59940
rect 18700 59810 18800 59940
rect 18950 59810 19050 59940
rect 19200 59810 19300 59940
rect 19450 59810 19550 59940
rect 19700 59810 19800 59940
rect 19950 59810 20050 59940
rect 20200 59810 20300 59940
rect 20450 59810 20550 59940
rect 20700 59810 20800 59940
rect 20950 59810 21050 59940
rect 21200 59810 21300 59940
rect 21450 59810 21550 59940
rect 21700 59810 21800 59940
rect 21950 59810 22050 59940
rect 22200 59810 22300 59940
rect 22450 59810 22550 59940
rect 22700 59810 22800 59940
rect 22950 59810 23050 59940
rect 23200 59810 23300 59940
rect 23450 59810 23550 59940
rect 23700 59810 23800 59940
rect 23950 59810 24050 59940
rect 24200 59810 24300 59940
rect 24450 59810 24550 59940
rect 24700 59810 24800 59940
rect 24950 59810 25050 59940
rect 25200 59810 25300 59940
rect 25450 59810 25550 59940
rect 25700 59810 25800 59940
rect 25950 59810 26050 59940
rect 26200 59810 26300 59940
rect 26450 59810 26550 59940
rect 26700 59810 26800 59940
rect 26950 59810 27050 59940
rect 27200 59810 27300 59940
rect 27450 59810 27550 59940
rect 27700 59810 27800 59940
rect 27950 59810 28050 59940
rect 28200 59810 28300 59940
rect 28450 59810 28550 59940
rect 28700 59810 28800 59940
rect 28950 59810 29000 59940
rect 7000 59800 7060 59810
rect 7190 59800 7310 59810
rect 7440 59800 7560 59810
rect 7690 59800 7810 59810
rect 7940 59800 8060 59810
rect 8190 59800 8310 59810
rect 8440 59800 8560 59810
rect 8690 59800 8810 59810
rect 8940 59800 9060 59810
rect 9190 59800 9310 59810
rect 9440 59800 9560 59810
rect 9690 59800 9810 59810
rect 9940 59800 10060 59810
rect 10190 59800 10310 59810
rect 10440 59800 10560 59810
rect 10690 59800 10810 59810
rect 10940 59800 11060 59810
rect 11190 59800 11310 59810
rect 11440 59800 11560 59810
rect 11690 59800 11810 59810
rect 11940 59800 12060 59810
rect 12190 59800 12310 59810
rect 12440 59800 12560 59810
rect 12690 59800 12810 59810
rect 12940 59800 13060 59810
rect 13190 59800 13310 59810
rect 13440 59800 13560 59810
rect 13690 59800 13810 59810
rect 13940 59800 14060 59810
rect 14190 59800 14310 59810
rect 14440 59800 14560 59810
rect 14690 59800 14810 59810
rect 14940 59800 15060 59810
rect 15190 59800 15310 59810
rect 15440 59800 15560 59810
rect 15690 59800 15810 59810
rect 15940 59800 16060 59810
rect 16190 59800 16310 59810
rect 16440 59800 16560 59810
rect 16690 59800 16810 59810
rect 16940 59800 17060 59810
rect 17190 59800 17310 59810
rect 17440 59800 17560 59810
rect 17690 59800 17810 59810
rect 17940 59800 18060 59810
rect 18190 59800 18310 59810
rect 18440 59800 18560 59810
rect 18690 59800 18810 59810
rect 18940 59800 19060 59810
rect 19190 59800 19310 59810
rect 19440 59800 19560 59810
rect 19690 59800 19810 59810
rect 19940 59800 20060 59810
rect 20190 59800 20310 59810
rect 20440 59800 20560 59810
rect 20690 59800 20810 59810
rect 20940 59800 21060 59810
rect 21190 59800 21310 59810
rect 21440 59800 21560 59810
rect 21690 59800 21810 59810
rect 21940 59800 22060 59810
rect 22190 59800 22310 59810
rect 22440 59800 22560 59810
rect 22690 59800 22810 59810
rect 22940 59800 23060 59810
rect 23190 59800 23310 59810
rect 23440 59800 23560 59810
rect 23690 59800 23810 59810
rect 23940 59800 24060 59810
rect 24190 59800 24310 59810
rect 24440 59800 24560 59810
rect 24690 59800 24810 59810
rect 24940 59800 25060 59810
rect 25190 59800 25310 59810
rect 25440 59800 25560 59810
rect 25690 59800 25810 59810
rect 25940 59800 26060 59810
rect 26190 59800 26310 59810
rect 26440 59800 26560 59810
rect 26690 59800 26810 59810
rect 26940 59800 27060 59810
rect 27190 59800 27310 59810
rect 27440 59800 27560 59810
rect 27690 59800 27810 59810
rect 27940 59800 28060 59810
rect 28190 59800 28310 59810
rect 28440 59800 28560 59810
rect 28690 59800 28810 59810
rect 28940 59800 29000 59810
rect 7000 59700 29000 59800
rect 7000 59690 7060 59700
rect 7190 59690 7310 59700
rect 7440 59690 7560 59700
rect 7690 59690 7810 59700
rect 7940 59690 8060 59700
rect 8190 59690 8310 59700
rect 8440 59690 8560 59700
rect 8690 59690 8810 59700
rect 8940 59690 9060 59700
rect 9190 59690 9310 59700
rect 9440 59690 9560 59700
rect 9690 59690 9810 59700
rect 9940 59690 10060 59700
rect 10190 59690 10310 59700
rect 10440 59690 10560 59700
rect 10690 59690 10810 59700
rect 10940 59690 11060 59700
rect 11190 59690 11310 59700
rect 11440 59690 11560 59700
rect 11690 59690 11810 59700
rect 11940 59690 12060 59700
rect 12190 59690 12310 59700
rect 12440 59690 12560 59700
rect 12690 59690 12810 59700
rect 12940 59690 13060 59700
rect 13190 59690 13310 59700
rect 13440 59690 13560 59700
rect 13690 59690 13810 59700
rect 13940 59690 14060 59700
rect 14190 59690 14310 59700
rect 14440 59690 14560 59700
rect 14690 59690 14810 59700
rect 14940 59690 15060 59700
rect 15190 59690 15310 59700
rect 15440 59690 15560 59700
rect 15690 59690 15810 59700
rect 15940 59690 16060 59700
rect 16190 59690 16310 59700
rect 16440 59690 16560 59700
rect 16690 59690 16810 59700
rect 16940 59690 17060 59700
rect 17190 59690 17310 59700
rect 17440 59690 17560 59700
rect 17690 59690 17810 59700
rect 17940 59690 18060 59700
rect 18190 59690 18310 59700
rect 18440 59690 18560 59700
rect 18690 59690 18810 59700
rect 18940 59690 19060 59700
rect 19190 59690 19310 59700
rect 19440 59690 19560 59700
rect 19690 59690 19810 59700
rect 19940 59690 20060 59700
rect 20190 59690 20310 59700
rect 20440 59690 20560 59700
rect 20690 59690 20810 59700
rect 20940 59690 21060 59700
rect 21190 59690 21310 59700
rect 21440 59690 21560 59700
rect 21690 59690 21810 59700
rect 21940 59690 22060 59700
rect 22190 59690 22310 59700
rect 22440 59690 22560 59700
rect 22690 59690 22810 59700
rect 22940 59690 23060 59700
rect 23190 59690 23310 59700
rect 23440 59690 23560 59700
rect 23690 59690 23810 59700
rect 23940 59690 24060 59700
rect 24190 59690 24310 59700
rect 24440 59690 24560 59700
rect 24690 59690 24810 59700
rect 24940 59690 25060 59700
rect 25190 59690 25310 59700
rect 25440 59690 25560 59700
rect 25690 59690 25810 59700
rect 25940 59690 26060 59700
rect 26190 59690 26310 59700
rect 26440 59690 26560 59700
rect 26690 59690 26810 59700
rect 26940 59690 27060 59700
rect 27190 59690 27310 59700
rect 27440 59690 27560 59700
rect 27690 59690 27810 59700
rect 27940 59690 28060 59700
rect 28190 59690 28310 59700
rect 28440 59690 28560 59700
rect 28690 59690 28810 59700
rect 28940 59690 29000 59700
rect 7000 59560 7050 59690
rect 7200 59560 7300 59690
rect 7450 59560 7550 59690
rect 7700 59560 7800 59690
rect 7950 59560 8050 59690
rect 8200 59560 8300 59690
rect 8450 59560 8550 59690
rect 8700 59560 8800 59690
rect 8950 59560 9050 59690
rect 9200 59560 9300 59690
rect 9450 59560 9550 59690
rect 9700 59560 9800 59690
rect 9950 59560 10050 59690
rect 10200 59560 10300 59690
rect 10450 59560 10550 59690
rect 10700 59560 10800 59690
rect 10950 59560 11050 59690
rect 11200 59560 11300 59690
rect 11450 59560 11550 59690
rect 11700 59560 11800 59690
rect 11950 59560 12050 59690
rect 12200 59560 12300 59690
rect 12450 59560 12550 59690
rect 12700 59560 12800 59690
rect 12950 59560 13050 59690
rect 13200 59560 13300 59690
rect 13450 59560 13550 59690
rect 13700 59560 13800 59690
rect 13950 59560 14050 59690
rect 14200 59560 14300 59690
rect 14450 59560 14550 59690
rect 14700 59560 14800 59690
rect 14950 59560 15050 59690
rect 15200 59560 15300 59690
rect 15450 59560 15550 59690
rect 15700 59560 15800 59690
rect 15950 59560 16050 59690
rect 16200 59560 16300 59690
rect 16450 59560 16550 59690
rect 16700 59560 16800 59690
rect 16950 59560 17050 59690
rect 17200 59560 17300 59690
rect 17450 59560 17550 59690
rect 17700 59560 17800 59690
rect 17950 59560 18050 59690
rect 18200 59560 18300 59690
rect 18450 59560 18550 59690
rect 18700 59560 18800 59690
rect 18950 59560 19050 59690
rect 19200 59560 19300 59690
rect 19450 59560 19550 59690
rect 19700 59560 19800 59690
rect 19950 59560 20050 59690
rect 20200 59560 20300 59690
rect 20450 59560 20550 59690
rect 20700 59560 20800 59690
rect 20950 59560 21050 59690
rect 21200 59560 21300 59690
rect 21450 59560 21550 59690
rect 21700 59560 21800 59690
rect 21950 59560 22050 59690
rect 22200 59560 22300 59690
rect 22450 59560 22550 59690
rect 22700 59560 22800 59690
rect 22950 59560 23050 59690
rect 23200 59560 23300 59690
rect 23450 59560 23550 59690
rect 23700 59560 23800 59690
rect 23950 59560 24050 59690
rect 24200 59560 24300 59690
rect 24450 59560 24550 59690
rect 24700 59560 24800 59690
rect 24950 59560 25050 59690
rect 25200 59560 25300 59690
rect 25450 59560 25550 59690
rect 25700 59560 25800 59690
rect 25950 59560 26050 59690
rect 26200 59560 26300 59690
rect 26450 59560 26550 59690
rect 26700 59560 26800 59690
rect 26950 59560 27050 59690
rect 27200 59560 27300 59690
rect 27450 59560 27550 59690
rect 27700 59560 27800 59690
rect 27950 59560 28050 59690
rect 28200 59560 28300 59690
rect 28450 59560 28550 59690
rect 28700 59560 28800 59690
rect 28950 59560 29000 59690
rect 7000 59550 7060 59560
rect 7190 59550 7310 59560
rect 7440 59550 7560 59560
rect 7690 59550 7810 59560
rect 7940 59550 8060 59560
rect 8190 59550 8310 59560
rect 8440 59550 8560 59560
rect 8690 59550 8810 59560
rect 8940 59550 9060 59560
rect 9190 59550 9310 59560
rect 9440 59550 9560 59560
rect 9690 59550 9810 59560
rect 9940 59550 10060 59560
rect 10190 59550 10310 59560
rect 10440 59550 10560 59560
rect 10690 59550 10810 59560
rect 10940 59550 11060 59560
rect 11190 59550 11310 59560
rect 11440 59550 11560 59560
rect 11690 59550 11810 59560
rect 11940 59550 12060 59560
rect 12190 59550 12310 59560
rect 12440 59550 12560 59560
rect 12690 59550 12810 59560
rect 12940 59550 13060 59560
rect 13190 59550 13310 59560
rect 13440 59550 13560 59560
rect 13690 59550 13810 59560
rect 13940 59550 14060 59560
rect 14190 59550 14310 59560
rect 14440 59550 14560 59560
rect 14690 59550 14810 59560
rect 14940 59550 15060 59560
rect 15190 59550 15310 59560
rect 15440 59550 15560 59560
rect 15690 59550 15810 59560
rect 15940 59550 16060 59560
rect 16190 59550 16310 59560
rect 16440 59550 16560 59560
rect 16690 59550 16810 59560
rect 16940 59550 17060 59560
rect 17190 59550 17310 59560
rect 17440 59550 17560 59560
rect 17690 59550 17810 59560
rect 17940 59550 18060 59560
rect 18190 59550 18310 59560
rect 18440 59550 18560 59560
rect 18690 59550 18810 59560
rect 18940 59550 19060 59560
rect 19190 59550 19310 59560
rect 19440 59550 19560 59560
rect 19690 59550 19810 59560
rect 19940 59550 20060 59560
rect 20190 59550 20310 59560
rect 20440 59550 20560 59560
rect 20690 59550 20810 59560
rect 20940 59550 21060 59560
rect 21190 59550 21310 59560
rect 21440 59550 21560 59560
rect 21690 59550 21810 59560
rect 21940 59550 22060 59560
rect 22190 59550 22310 59560
rect 22440 59550 22560 59560
rect 22690 59550 22810 59560
rect 22940 59550 23060 59560
rect 23190 59550 23310 59560
rect 23440 59550 23560 59560
rect 23690 59550 23810 59560
rect 23940 59550 24060 59560
rect 24190 59550 24310 59560
rect 24440 59550 24560 59560
rect 24690 59550 24810 59560
rect 24940 59550 25060 59560
rect 25190 59550 25310 59560
rect 25440 59550 25560 59560
rect 25690 59550 25810 59560
rect 25940 59550 26060 59560
rect 26190 59550 26310 59560
rect 26440 59550 26560 59560
rect 26690 59550 26810 59560
rect 26940 59550 27060 59560
rect 27190 59550 27310 59560
rect 27440 59550 27560 59560
rect 27690 59550 27810 59560
rect 27940 59550 28060 59560
rect 28190 59550 28310 59560
rect 28440 59550 28560 59560
rect 28690 59550 28810 59560
rect 28940 59550 29000 59560
rect 7000 59450 29000 59550
rect 7000 59440 7060 59450
rect 7190 59440 7310 59450
rect 7440 59440 7560 59450
rect 7690 59440 7810 59450
rect 7940 59440 8060 59450
rect 8190 59440 8310 59450
rect 8440 59440 8560 59450
rect 8690 59440 8810 59450
rect 8940 59440 9060 59450
rect 9190 59440 9310 59450
rect 9440 59440 9560 59450
rect 9690 59440 9810 59450
rect 9940 59440 10060 59450
rect 10190 59440 10310 59450
rect 10440 59440 10560 59450
rect 10690 59440 10810 59450
rect 10940 59440 11060 59450
rect 11190 59440 11310 59450
rect 11440 59440 11560 59450
rect 11690 59440 11810 59450
rect 11940 59440 12060 59450
rect 12190 59440 12310 59450
rect 12440 59440 12560 59450
rect 12690 59440 12810 59450
rect 12940 59440 13060 59450
rect 13190 59440 13310 59450
rect 13440 59440 13560 59450
rect 13690 59440 13810 59450
rect 13940 59440 14060 59450
rect 14190 59440 14310 59450
rect 14440 59440 14560 59450
rect 14690 59440 14810 59450
rect 14940 59440 15060 59450
rect 15190 59440 15310 59450
rect 15440 59440 15560 59450
rect 15690 59440 15810 59450
rect 15940 59440 16060 59450
rect 16190 59440 16310 59450
rect 16440 59440 16560 59450
rect 16690 59440 16810 59450
rect 16940 59440 17060 59450
rect 17190 59440 17310 59450
rect 17440 59440 17560 59450
rect 17690 59440 17810 59450
rect 17940 59440 18060 59450
rect 18190 59440 18310 59450
rect 18440 59440 18560 59450
rect 18690 59440 18810 59450
rect 18940 59440 19060 59450
rect 19190 59440 19310 59450
rect 19440 59440 19560 59450
rect 19690 59440 19810 59450
rect 19940 59440 20060 59450
rect 20190 59440 20310 59450
rect 20440 59440 20560 59450
rect 20690 59440 20810 59450
rect 20940 59440 21060 59450
rect 21190 59440 21310 59450
rect 21440 59440 21560 59450
rect 21690 59440 21810 59450
rect 21940 59440 22060 59450
rect 22190 59440 22310 59450
rect 22440 59440 22560 59450
rect 22690 59440 22810 59450
rect 22940 59440 23060 59450
rect 23190 59440 23310 59450
rect 23440 59440 23560 59450
rect 23690 59440 23810 59450
rect 23940 59440 24060 59450
rect 24190 59440 24310 59450
rect 24440 59440 24560 59450
rect 24690 59440 24810 59450
rect 24940 59440 25060 59450
rect 25190 59440 25310 59450
rect 25440 59440 25560 59450
rect 25690 59440 25810 59450
rect 25940 59440 26060 59450
rect 26190 59440 26310 59450
rect 26440 59440 26560 59450
rect 26690 59440 26810 59450
rect 26940 59440 27060 59450
rect 27190 59440 27310 59450
rect 27440 59440 27560 59450
rect 27690 59440 27810 59450
rect 27940 59440 28060 59450
rect 28190 59440 28310 59450
rect 28440 59440 28560 59450
rect 28690 59440 28810 59450
rect 28940 59440 29000 59450
rect 7000 59310 7050 59440
rect 7200 59310 7300 59440
rect 7450 59310 7550 59440
rect 7700 59310 7800 59440
rect 7950 59310 8050 59440
rect 8200 59310 8300 59440
rect 8450 59310 8550 59440
rect 8700 59310 8800 59440
rect 8950 59310 9050 59440
rect 9200 59310 9300 59440
rect 9450 59310 9550 59440
rect 9700 59310 9800 59440
rect 9950 59310 10050 59440
rect 10200 59310 10300 59440
rect 10450 59310 10550 59440
rect 10700 59310 10800 59440
rect 10950 59310 11050 59440
rect 11200 59310 11300 59440
rect 11450 59310 11550 59440
rect 11700 59310 11800 59440
rect 11950 59310 12050 59440
rect 12200 59310 12300 59440
rect 12450 59310 12550 59440
rect 12700 59310 12800 59440
rect 12950 59310 13050 59440
rect 13200 59310 13300 59440
rect 13450 59310 13550 59440
rect 13700 59310 13800 59440
rect 13950 59310 14050 59440
rect 14200 59310 14300 59440
rect 14450 59310 14550 59440
rect 14700 59310 14800 59440
rect 14950 59310 15050 59440
rect 15200 59310 15300 59440
rect 15450 59310 15550 59440
rect 15700 59310 15800 59440
rect 15950 59310 16050 59440
rect 16200 59310 16300 59440
rect 16450 59310 16550 59440
rect 16700 59310 16800 59440
rect 16950 59310 17050 59440
rect 17200 59310 17300 59440
rect 17450 59310 17550 59440
rect 17700 59310 17800 59440
rect 17950 59310 18050 59440
rect 18200 59310 18300 59440
rect 18450 59310 18550 59440
rect 18700 59310 18800 59440
rect 18950 59310 19050 59440
rect 19200 59310 19300 59440
rect 19450 59310 19550 59440
rect 19700 59310 19800 59440
rect 19950 59310 20050 59440
rect 20200 59310 20300 59440
rect 20450 59310 20550 59440
rect 20700 59310 20800 59440
rect 20950 59310 21050 59440
rect 21200 59310 21300 59440
rect 21450 59310 21550 59440
rect 21700 59310 21800 59440
rect 21950 59310 22050 59440
rect 22200 59310 22300 59440
rect 22450 59310 22550 59440
rect 22700 59310 22800 59440
rect 22950 59310 23050 59440
rect 23200 59310 23300 59440
rect 23450 59310 23550 59440
rect 23700 59310 23800 59440
rect 23950 59310 24050 59440
rect 24200 59310 24300 59440
rect 24450 59310 24550 59440
rect 24700 59310 24800 59440
rect 24950 59310 25050 59440
rect 25200 59310 25300 59440
rect 25450 59310 25550 59440
rect 25700 59310 25800 59440
rect 25950 59310 26050 59440
rect 26200 59310 26300 59440
rect 26450 59310 26550 59440
rect 26700 59310 26800 59440
rect 26950 59310 27050 59440
rect 27200 59310 27300 59440
rect 27450 59310 27550 59440
rect 27700 59310 27800 59440
rect 27950 59310 28050 59440
rect 28200 59310 28300 59440
rect 28450 59310 28550 59440
rect 28700 59310 28800 59440
rect 28950 59310 29000 59440
rect 7000 59300 7060 59310
rect 7190 59300 7310 59310
rect 7440 59300 7560 59310
rect 7690 59300 7810 59310
rect 7940 59300 8060 59310
rect 8190 59300 8310 59310
rect 8440 59300 8560 59310
rect 8690 59300 8810 59310
rect 8940 59300 9060 59310
rect 9190 59300 9310 59310
rect 9440 59300 9560 59310
rect 9690 59300 9810 59310
rect 9940 59300 10060 59310
rect 10190 59300 10310 59310
rect 10440 59300 10560 59310
rect 10690 59300 10810 59310
rect 10940 59300 11060 59310
rect 11190 59300 11310 59310
rect 11440 59300 11560 59310
rect 11690 59300 11810 59310
rect 11940 59300 12060 59310
rect 12190 59300 12310 59310
rect 12440 59300 12560 59310
rect 12690 59300 12810 59310
rect 12940 59300 13060 59310
rect 13190 59300 13310 59310
rect 13440 59300 13560 59310
rect 13690 59300 13810 59310
rect 13940 59300 14060 59310
rect 14190 59300 14310 59310
rect 14440 59300 14560 59310
rect 14690 59300 14810 59310
rect 14940 59300 15060 59310
rect 15190 59300 15310 59310
rect 15440 59300 15560 59310
rect 15690 59300 15810 59310
rect 15940 59300 16060 59310
rect 16190 59300 16310 59310
rect 16440 59300 16560 59310
rect 16690 59300 16810 59310
rect 16940 59300 17060 59310
rect 17190 59300 17310 59310
rect 17440 59300 17560 59310
rect 17690 59300 17810 59310
rect 17940 59300 18060 59310
rect 18190 59300 18310 59310
rect 18440 59300 18560 59310
rect 18690 59300 18810 59310
rect 18940 59300 19060 59310
rect 19190 59300 19310 59310
rect 19440 59300 19560 59310
rect 19690 59300 19810 59310
rect 19940 59300 20060 59310
rect 20190 59300 20310 59310
rect 20440 59300 20560 59310
rect 20690 59300 20810 59310
rect 20940 59300 21060 59310
rect 21190 59300 21310 59310
rect 21440 59300 21560 59310
rect 21690 59300 21810 59310
rect 21940 59300 22060 59310
rect 22190 59300 22310 59310
rect 22440 59300 22560 59310
rect 22690 59300 22810 59310
rect 22940 59300 23060 59310
rect 23190 59300 23310 59310
rect 23440 59300 23560 59310
rect 23690 59300 23810 59310
rect 23940 59300 24060 59310
rect 24190 59300 24310 59310
rect 24440 59300 24560 59310
rect 24690 59300 24810 59310
rect 24940 59300 25060 59310
rect 25190 59300 25310 59310
rect 25440 59300 25560 59310
rect 25690 59300 25810 59310
rect 25940 59300 26060 59310
rect 26190 59300 26310 59310
rect 26440 59300 26560 59310
rect 26690 59300 26810 59310
rect 26940 59300 27060 59310
rect 27190 59300 27310 59310
rect 27440 59300 27560 59310
rect 27690 59300 27810 59310
rect 27940 59300 28060 59310
rect 28190 59300 28310 59310
rect 28440 59300 28560 59310
rect 28690 59300 28810 59310
rect 28940 59300 29000 59310
rect 7000 59200 29000 59300
rect 7000 59190 7060 59200
rect 7190 59190 7310 59200
rect 7440 59190 7560 59200
rect 7690 59190 7810 59200
rect 7940 59190 8060 59200
rect 8190 59190 8310 59200
rect 8440 59190 8560 59200
rect 8690 59190 8810 59200
rect 8940 59190 9060 59200
rect 9190 59190 9310 59200
rect 9440 59190 9560 59200
rect 9690 59190 9810 59200
rect 9940 59190 10060 59200
rect 10190 59190 10310 59200
rect 10440 59190 10560 59200
rect 10690 59190 10810 59200
rect 10940 59190 11060 59200
rect 11190 59190 11310 59200
rect 11440 59190 11560 59200
rect 11690 59190 11810 59200
rect 11940 59190 12060 59200
rect 12190 59190 12310 59200
rect 12440 59190 12560 59200
rect 12690 59190 12810 59200
rect 12940 59190 13060 59200
rect 13190 59190 13310 59200
rect 13440 59190 13560 59200
rect 13690 59190 13810 59200
rect 13940 59190 14060 59200
rect 14190 59190 14310 59200
rect 14440 59190 14560 59200
rect 14690 59190 14810 59200
rect 14940 59190 15060 59200
rect 15190 59190 15310 59200
rect 15440 59190 15560 59200
rect 15690 59190 15810 59200
rect 15940 59190 16060 59200
rect 16190 59190 16310 59200
rect 16440 59190 16560 59200
rect 16690 59190 16810 59200
rect 16940 59190 17060 59200
rect 17190 59190 17310 59200
rect 17440 59190 17560 59200
rect 17690 59190 17810 59200
rect 17940 59190 18060 59200
rect 18190 59190 18310 59200
rect 18440 59190 18560 59200
rect 18690 59190 18810 59200
rect 18940 59190 19060 59200
rect 19190 59190 19310 59200
rect 19440 59190 19560 59200
rect 19690 59190 19810 59200
rect 19940 59190 20060 59200
rect 20190 59190 20310 59200
rect 20440 59190 20560 59200
rect 20690 59190 20810 59200
rect 20940 59190 21060 59200
rect 21190 59190 21310 59200
rect 21440 59190 21560 59200
rect 21690 59190 21810 59200
rect 21940 59190 22060 59200
rect 22190 59190 22310 59200
rect 22440 59190 22560 59200
rect 22690 59190 22810 59200
rect 22940 59190 23060 59200
rect 23190 59190 23310 59200
rect 23440 59190 23560 59200
rect 23690 59190 23810 59200
rect 23940 59190 24060 59200
rect 24190 59190 24310 59200
rect 24440 59190 24560 59200
rect 24690 59190 24810 59200
rect 24940 59190 25060 59200
rect 25190 59190 25310 59200
rect 25440 59190 25560 59200
rect 25690 59190 25810 59200
rect 25940 59190 26060 59200
rect 26190 59190 26310 59200
rect 26440 59190 26560 59200
rect 26690 59190 26810 59200
rect 26940 59190 27060 59200
rect 27190 59190 27310 59200
rect 27440 59190 27560 59200
rect 27690 59190 27810 59200
rect 27940 59190 28060 59200
rect 28190 59190 28310 59200
rect 28440 59190 28560 59200
rect 28690 59190 28810 59200
rect 28940 59190 29000 59200
rect 7000 59060 7050 59190
rect 7200 59060 7300 59190
rect 7450 59060 7550 59190
rect 7700 59060 7800 59190
rect 7950 59060 8050 59190
rect 8200 59060 8300 59190
rect 8450 59060 8550 59190
rect 8700 59060 8800 59190
rect 8950 59060 9050 59190
rect 9200 59060 9300 59190
rect 9450 59060 9550 59190
rect 9700 59060 9800 59190
rect 9950 59060 10050 59190
rect 10200 59060 10300 59190
rect 10450 59060 10550 59190
rect 10700 59060 10800 59190
rect 10950 59060 11050 59190
rect 11200 59060 11300 59190
rect 11450 59060 11550 59190
rect 11700 59060 11800 59190
rect 11950 59060 12050 59190
rect 12200 59060 12300 59190
rect 12450 59060 12550 59190
rect 12700 59060 12800 59190
rect 12950 59060 13050 59190
rect 13200 59060 13300 59190
rect 13450 59060 13550 59190
rect 13700 59060 13800 59190
rect 13950 59060 14050 59190
rect 14200 59060 14300 59190
rect 14450 59060 14550 59190
rect 14700 59060 14800 59190
rect 14950 59060 15050 59190
rect 15200 59060 15300 59190
rect 15450 59060 15550 59190
rect 15700 59060 15800 59190
rect 15950 59060 16050 59190
rect 16200 59060 16300 59190
rect 16450 59060 16550 59190
rect 16700 59060 16800 59190
rect 16950 59060 17050 59190
rect 17200 59060 17300 59190
rect 17450 59060 17550 59190
rect 17700 59060 17800 59190
rect 17950 59060 18050 59190
rect 18200 59060 18300 59190
rect 18450 59060 18550 59190
rect 18700 59060 18800 59190
rect 18950 59060 19050 59190
rect 19200 59060 19300 59190
rect 19450 59060 19550 59190
rect 19700 59060 19800 59190
rect 19950 59060 20050 59190
rect 20200 59060 20300 59190
rect 20450 59060 20550 59190
rect 20700 59060 20800 59190
rect 20950 59060 21050 59190
rect 21200 59060 21300 59190
rect 21450 59060 21550 59190
rect 21700 59060 21800 59190
rect 21950 59060 22050 59190
rect 22200 59060 22300 59190
rect 22450 59060 22550 59190
rect 22700 59060 22800 59190
rect 22950 59060 23050 59190
rect 23200 59060 23300 59190
rect 23450 59060 23550 59190
rect 23700 59060 23800 59190
rect 23950 59060 24050 59190
rect 24200 59060 24300 59190
rect 24450 59060 24550 59190
rect 24700 59060 24800 59190
rect 24950 59060 25050 59190
rect 25200 59060 25300 59190
rect 25450 59060 25550 59190
rect 25700 59060 25800 59190
rect 25950 59060 26050 59190
rect 26200 59060 26300 59190
rect 26450 59060 26550 59190
rect 26700 59060 26800 59190
rect 26950 59060 27050 59190
rect 27200 59060 27300 59190
rect 27450 59060 27550 59190
rect 27700 59060 27800 59190
rect 27950 59060 28050 59190
rect 28200 59060 28300 59190
rect 28450 59060 28550 59190
rect 28700 59060 28800 59190
rect 28950 59060 29000 59190
rect 7000 59050 7060 59060
rect 7190 59050 7310 59060
rect 7440 59050 7560 59060
rect 7690 59050 7810 59060
rect 7940 59050 8060 59060
rect 8190 59050 8310 59060
rect 8440 59050 8560 59060
rect 8690 59050 8810 59060
rect 8940 59050 9060 59060
rect 9190 59050 9310 59060
rect 9440 59050 9560 59060
rect 9690 59050 9810 59060
rect 9940 59050 10060 59060
rect 10190 59050 10310 59060
rect 10440 59050 10560 59060
rect 10690 59050 10810 59060
rect 10940 59050 11060 59060
rect 11190 59050 11310 59060
rect 11440 59050 11560 59060
rect 11690 59050 11810 59060
rect 11940 59050 12060 59060
rect 12190 59050 12310 59060
rect 12440 59050 12560 59060
rect 12690 59050 12810 59060
rect 12940 59050 13060 59060
rect 13190 59050 13310 59060
rect 13440 59050 13560 59060
rect 13690 59050 13810 59060
rect 13940 59050 14060 59060
rect 14190 59050 14310 59060
rect 14440 59050 14560 59060
rect 14690 59050 14810 59060
rect 14940 59050 15060 59060
rect 15190 59050 15310 59060
rect 15440 59050 15560 59060
rect 15690 59050 15810 59060
rect 15940 59050 16060 59060
rect 16190 59050 16310 59060
rect 16440 59050 16560 59060
rect 16690 59050 16810 59060
rect 16940 59050 17060 59060
rect 17190 59050 17310 59060
rect 17440 59050 17560 59060
rect 17690 59050 17810 59060
rect 17940 59050 18060 59060
rect 18190 59050 18310 59060
rect 18440 59050 18560 59060
rect 18690 59050 18810 59060
rect 18940 59050 19060 59060
rect 19190 59050 19310 59060
rect 19440 59050 19560 59060
rect 19690 59050 19810 59060
rect 19940 59050 20060 59060
rect 20190 59050 20310 59060
rect 20440 59050 20560 59060
rect 20690 59050 20810 59060
rect 20940 59050 21060 59060
rect 21190 59050 21310 59060
rect 21440 59050 21560 59060
rect 21690 59050 21810 59060
rect 21940 59050 22060 59060
rect 22190 59050 22310 59060
rect 22440 59050 22560 59060
rect 22690 59050 22810 59060
rect 22940 59050 23060 59060
rect 23190 59050 23310 59060
rect 23440 59050 23560 59060
rect 23690 59050 23810 59060
rect 23940 59050 24060 59060
rect 24190 59050 24310 59060
rect 24440 59050 24560 59060
rect 24690 59050 24810 59060
rect 24940 59050 25060 59060
rect 25190 59050 25310 59060
rect 25440 59050 25560 59060
rect 25690 59050 25810 59060
rect 25940 59050 26060 59060
rect 26190 59050 26310 59060
rect 26440 59050 26560 59060
rect 26690 59050 26810 59060
rect 26940 59050 27060 59060
rect 27190 59050 27310 59060
rect 27440 59050 27560 59060
rect 27690 59050 27810 59060
rect 27940 59050 28060 59060
rect 28190 59050 28310 59060
rect 28440 59050 28560 59060
rect 28690 59050 28810 59060
rect 28940 59050 29000 59060
rect 7000 58950 29000 59050
rect 7000 58940 7060 58950
rect 7190 58940 7310 58950
rect 7440 58940 7560 58950
rect 7690 58940 7810 58950
rect 7940 58940 8060 58950
rect 8190 58940 8310 58950
rect 8440 58940 8560 58950
rect 8690 58940 8810 58950
rect 8940 58940 9060 58950
rect 9190 58940 9310 58950
rect 9440 58940 9560 58950
rect 9690 58940 9810 58950
rect 9940 58940 10060 58950
rect 10190 58940 10310 58950
rect 10440 58940 10560 58950
rect 10690 58940 10810 58950
rect 10940 58940 11060 58950
rect 11190 58940 11310 58950
rect 11440 58940 11560 58950
rect 11690 58940 11810 58950
rect 11940 58940 12060 58950
rect 12190 58940 12310 58950
rect 12440 58940 12560 58950
rect 12690 58940 12810 58950
rect 12940 58940 13060 58950
rect 13190 58940 13310 58950
rect 13440 58940 13560 58950
rect 13690 58940 13810 58950
rect 13940 58940 14060 58950
rect 14190 58940 14310 58950
rect 14440 58940 14560 58950
rect 14690 58940 14810 58950
rect 14940 58940 15060 58950
rect 15190 58940 15310 58950
rect 15440 58940 15560 58950
rect 15690 58940 15810 58950
rect 15940 58940 16060 58950
rect 16190 58940 16310 58950
rect 16440 58940 16560 58950
rect 16690 58940 16810 58950
rect 16940 58940 17060 58950
rect 17190 58940 17310 58950
rect 17440 58940 17560 58950
rect 17690 58940 17810 58950
rect 17940 58940 18060 58950
rect 18190 58940 18310 58950
rect 18440 58940 18560 58950
rect 18690 58940 18810 58950
rect 18940 58940 19060 58950
rect 19190 58940 19310 58950
rect 19440 58940 19560 58950
rect 19690 58940 19810 58950
rect 19940 58940 20060 58950
rect 20190 58940 20310 58950
rect 20440 58940 20560 58950
rect 20690 58940 20810 58950
rect 20940 58940 21060 58950
rect 21190 58940 21310 58950
rect 21440 58940 21560 58950
rect 21690 58940 21810 58950
rect 21940 58940 22060 58950
rect 22190 58940 22310 58950
rect 22440 58940 22560 58950
rect 22690 58940 22810 58950
rect 22940 58940 23060 58950
rect 23190 58940 23310 58950
rect 23440 58940 23560 58950
rect 23690 58940 23810 58950
rect 23940 58940 24060 58950
rect 24190 58940 24310 58950
rect 24440 58940 24560 58950
rect 24690 58940 24810 58950
rect 24940 58940 25060 58950
rect 25190 58940 25310 58950
rect 25440 58940 25560 58950
rect 25690 58940 25810 58950
rect 25940 58940 26060 58950
rect 26190 58940 26310 58950
rect 26440 58940 26560 58950
rect 26690 58940 26810 58950
rect 26940 58940 27060 58950
rect 27190 58940 27310 58950
rect 27440 58940 27560 58950
rect 27690 58940 27810 58950
rect 27940 58940 28060 58950
rect 28190 58940 28310 58950
rect 28440 58940 28560 58950
rect 28690 58940 28810 58950
rect 28940 58940 29000 58950
rect 7000 58810 7050 58940
rect 7200 58810 7300 58940
rect 7450 58810 7550 58940
rect 7700 58810 7800 58940
rect 7950 58810 8050 58940
rect 8200 58810 8300 58940
rect 8450 58810 8550 58940
rect 8700 58810 8800 58940
rect 8950 58810 9050 58940
rect 9200 58810 9300 58940
rect 9450 58810 9550 58940
rect 9700 58810 9800 58940
rect 9950 58810 10050 58940
rect 10200 58810 10300 58940
rect 10450 58810 10550 58940
rect 10700 58810 10800 58940
rect 10950 58810 11050 58940
rect 11200 58810 11300 58940
rect 11450 58810 11550 58940
rect 11700 58810 11800 58940
rect 11950 58810 12050 58940
rect 12200 58810 12300 58940
rect 12450 58810 12550 58940
rect 12700 58810 12800 58940
rect 12950 58810 13050 58940
rect 13200 58810 13300 58940
rect 13450 58810 13550 58940
rect 13700 58810 13800 58940
rect 13950 58810 14050 58940
rect 14200 58810 14300 58940
rect 14450 58810 14550 58940
rect 14700 58810 14800 58940
rect 14950 58810 15050 58940
rect 15200 58810 15300 58940
rect 15450 58810 15550 58940
rect 15700 58810 15800 58940
rect 15950 58810 16050 58940
rect 16200 58810 16300 58940
rect 16450 58810 16550 58940
rect 16700 58810 16800 58940
rect 16950 58810 17050 58940
rect 17200 58810 17300 58940
rect 17450 58810 17550 58940
rect 17700 58810 17800 58940
rect 17950 58810 18050 58940
rect 18200 58810 18300 58940
rect 18450 58810 18550 58940
rect 18700 58810 18800 58940
rect 18950 58810 19050 58940
rect 19200 58810 19300 58940
rect 19450 58810 19550 58940
rect 19700 58810 19800 58940
rect 19950 58810 20050 58940
rect 20200 58810 20300 58940
rect 20450 58810 20550 58940
rect 20700 58810 20800 58940
rect 20950 58810 21050 58940
rect 21200 58810 21300 58940
rect 21450 58810 21550 58940
rect 21700 58810 21800 58940
rect 21950 58810 22050 58940
rect 22200 58810 22300 58940
rect 22450 58810 22550 58940
rect 22700 58810 22800 58940
rect 22950 58810 23050 58940
rect 23200 58810 23300 58940
rect 23450 58810 23550 58940
rect 23700 58810 23800 58940
rect 23950 58810 24050 58940
rect 24200 58810 24300 58940
rect 24450 58810 24550 58940
rect 24700 58810 24800 58940
rect 24950 58810 25050 58940
rect 25200 58810 25300 58940
rect 25450 58810 25550 58940
rect 25700 58810 25800 58940
rect 25950 58810 26050 58940
rect 26200 58810 26300 58940
rect 26450 58810 26550 58940
rect 26700 58810 26800 58940
rect 26950 58810 27050 58940
rect 27200 58810 27300 58940
rect 27450 58810 27550 58940
rect 27700 58810 27800 58940
rect 27950 58810 28050 58940
rect 28200 58810 28300 58940
rect 28450 58810 28550 58940
rect 28700 58810 28800 58940
rect 28950 58810 29000 58940
rect 7000 58800 7060 58810
rect 7190 58800 7310 58810
rect 7440 58800 7560 58810
rect 7690 58800 7810 58810
rect 7940 58800 8060 58810
rect 8190 58800 8310 58810
rect 8440 58800 8560 58810
rect 8690 58800 8810 58810
rect 8940 58800 9060 58810
rect 9190 58800 9310 58810
rect 9440 58800 9560 58810
rect 9690 58800 9810 58810
rect 9940 58800 10060 58810
rect 10190 58800 10310 58810
rect 10440 58800 10560 58810
rect 10690 58800 10810 58810
rect 10940 58800 11060 58810
rect 11190 58800 11310 58810
rect 11440 58800 11560 58810
rect 11690 58800 11810 58810
rect 11940 58800 12060 58810
rect 12190 58800 12310 58810
rect 12440 58800 12560 58810
rect 12690 58800 12810 58810
rect 12940 58800 13060 58810
rect 13190 58800 13310 58810
rect 13440 58800 13560 58810
rect 13690 58800 13810 58810
rect 13940 58800 14060 58810
rect 14190 58800 14310 58810
rect 14440 58800 14560 58810
rect 14690 58800 14810 58810
rect 14940 58800 15060 58810
rect 15190 58800 15310 58810
rect 15440 58800 15560 58810
rect 15690 58800 15810 58810
rect 15940 58800 16060 58810
rect 16190 58800 16310 58810
rect 16440 58800 16560 58810
rect 16690 58800 16810 58810
rect 16940 58800 17060 58810
rect 17190 58800 17310 58810
rect 17440 58800 17560 58810
rect 17690 58800 17810 58810
rect 17940 58800 18060 58810
rect 18190 58800 18310 58810
rect 18440 58800 18560 58810
rect 18690 58800 18810 58810
rect 18940 58800 19060 58810
rect 19190 58800 19310 58810
rect 19440 58800 19560 58810
rect 19690 58800 19810 58810
rect 19940 58800 20060 58810
rect 20190 58800 20310 58810
rect 20440 58800 20560 58810
rect 20690 58800 20810 58810
rect 20940 58800 21060 58810
rect 21190 58800 21310 58810
rect 21440 58800 21560 58810
rect 21690 58800 21810 58810
rect 21940 58800 22060 58810
rect 22190 58800 22310 58810
rect 22440 58800 22560 58810
rect 22690 58800 22810 58810
rect 22940 58800 23060 58810
rect 23190 58800 23310 58810
rect 23440 58800 23560 58810
rect 23690 58800 23810 58810
rect 23940 58800 24060 58810
rect 24190 58800 24310 58810
rect 24440 58800 24560 58810
rect 24690 58800 24810 58810
rect 24940 58800 25060 58810
rect 25190 58800 25310 58810
rect 25440 58800 25560 58810
rect 25690 58800 25810 58810
rect 25940 58800 26060 58810
rect 26190 58800 26310 58810
rect 26440 58800 26560 58810
rect 26690 58800 26810 58810
rect 26940 58800 27060 58810
rect 27190 58800 27310 58810
rect 27440 58800 27560 58810
rect 27690 58800 27810 58810
rect 27940 58800 28060 58810
rect 28190 58800 28310 58810
rect 28440 58800 28560 58810
rect 28690 58800 28810 58810
rect 28940 58800 29000 58810
rect 7000 58700 29000 58800
rect 7000 58690 7060 58700
rect 7190 58690 7310 58700
rect 7440 58690 7560 58700
rect 7690 58690 7810 58700
rect 7940 58690 8060 58700
rect 8190 58690 8310 58700
rect 8440 58690 8560 58700
rect 8690 58690 8810 58700
rect 8940 58690 9060 58700
rect 9190 58690 9310 58700
rect 9440 58690 9560 58700
rect 9690 58690 9810 58700
rect 9940 58690 10060 58700
rect 10190 58690 10310 58700
rect 10440 58690 10560 58700
rect 10690 58690 10810 58700
rect 10940 58690 11060 58700
rect 11190 58690 11310 58700
rect 11440 58690 11560 58700
rect 11690 58690 11810 58700
rect 11940 58690 12060 58700
rect 12190 58690 12310 58700
rect 12440 58690 12560 58700
rect 12690 58690 12810 58700
rect 12940 58690 13060 58700
rect 13190 58690 13310 58700
rect 13440 58690 13560 58700
rect 13690 58690 13810 58700
rect 13940 58690 14060 58700
rect 14190 58690 14310 58700
rect 14440 58690 14560 58700
rect 14690 58690 14810 58700
rect 14940 58690 15060 58700
rect 15190 58690 15310 58700
rect 15440 58690 15560 58700
rect 15690 58690 15810 58700
rect 15940 58690 16060 58700
rect 16190 58690 16310 58700
rect 16440 58690 16560 58700
rect 16690 58690 16810 58700
rect 16940 58690 17060 58700
rect 17190 58690 17310 58700
rect 17440 58690 17560 58700
rect 17690 58690 17810 58700
rect 17940 58690 18060 58700
rect 18190 58690 18310 58700
rect 18440 58690 18560 58700
rect 18690 58690 18810 58700
rect 18940 58690 19060 58700
rect 19190 58690 19310 58700
rect 19440 58690 19560 58700
rect 19690 58690 19810 58700
rect 19940 58690 20060 58700
rect 20190 58690 20310 58700
rect 20440 58690 20560 58700
rect 20690 58690 20810 58700
rect 20940 58690 21060 58700
rect 21190 58690 21310 58700
rect 21440 58690 21560 58700
rect 21690 58690 21810 58700
rect 21940 58690 22060 58700
rect 22190 58690 22310 58700
rect 22440 58690 22560 58700
rect 22690 58690 22810 58700
rect 22940 58690 23060 58700
rect 23190 58690 23310 58700
rect 23440 58690 23560 58700
rect 23690 58690 23810 58700
rect 23940 58690 24060 58700
rect 24190 58690 24310 58700
rect 24440 58690 24560 58700
rect 24690 58690 24810 58700
rect 24940 58690 25060 58700
rect 25190 58690 25310 58700
rect 25440 58690 25560 58700
rect 25690 58690 25810 58700
rect 25940 58690 26060 58700
rect 26190 58690 26310 58700
rect 26440 58690 26560 58700
rect 26690 58690 26810 58700
rect 26940 58690 27060 58700
rect 27190 58690 27310 58700
rect 27440 58690 27560 58700
rect 27690 58690 27810 58700
rect 27940 58690 28060 58700
rect 28190 58690 28310 58700
rect 28440 58690 28560 58700
rect 28690 58690 28810 58700
rect 28940 58690 29000 58700
rect 7000 58560 7050 58690
rect 7200 58560 7300 58690
rect 7450 58560 7550 58690
rect 7700 58560 7800 58690
rect 7950 58560 8050 58690
rect 8200 58560 8300 58690
rect 8450 58560 8550 58690
rect 8700 58560 8800 58690
rect 8950 58560 9050 58690
rect 9200 58560 9300 58690
rect 9450 58560 9550 58690
rect 9700 58560 9800 58690
rect 9950 58560 10050 58690
rect 10200 58560 10300 58690
rect 10450 58560 10550 58690
rect 10700 58560 10800 58690
rect 10950 58560 11050 58690
rect 11200 58560 11300 58690
rect 11450 58560 11550 58690
rect 11700 58560 11800 58690
rect 11950 58560 12050 58690
rect 12200 58560 12300 58690
rect 12450 58560 12550 58690
rect 12700 58560 12800 58690
rect 12950 58560 13050 58690
rect 13200 58560 13300 58690
rect 13450 58560 13550 58690
rect 13700 58560 13800 58690
rect 13950 58560 14050 58690
rect 14200 58560 14300 58690
rect 14450 58560 14550 58690
rect 14700 58560 14800 58690
rect 14950 58560 15050 58690
rect 15200 58560 15300 58690
rect 15450 58560 15550 58690
rect 15700 58560 15800 58690
rect 15950 58560 16050 58690
rect 16200 58560 16300 58690
rect 16450 58560 16550 58690
rect 16700 58560 16800 58690
rect 16950 58560 17050 58690
rect 17200 58560 17300 58690
rect 17450 58560 17550 58690
rect 17700 58560 17800 58690
rect 17950 58560 18050 58690
rect 18200 58560 18300 58690
rect 18450 58560 18550 58690
rect 18700 58560 18800 58690
rect 18950 58560 19050 58690
rect 19200 58560 19300 58690
rect 19450 58560 19550 58690
rect 19700 58560 19800 58690
rect 19950 58560 20050 58690
rect 20200 58560 20300 58690
rect 20450 58560 20550 58690
rect 20700 58560 20800 58690
rect 20950 58560 21050 58690
rect 21200 58560 21300 58690
rect 21450 58560 21550 58690
rect 21700 58560 21800 58690
rect 21950 58560 22050 58690
rect 22200 58560 22300 58690
rect 22450 58560 22550 58690
rect 22700 58560 22800 58690
rect 22950 58560 23050 58690
rect 23200 58560 23300 58690
rect 23450 58560 23550 58690
rect 23700 58560 23800 58690
rect 23950 58560 24050 58690
rect 24200 58560 24300 58690
rect 24450 58560 24550 58690
rect 24700 58560 24800 58690
rect 24950 58560 25050 58690
rect 25200 58560 25300 58690
rect 25450 58560 25550 58690
rect 25700 58560 25800 58690
rect 25950 58560 26050 58690
rect 26200 58560 26300 58690
rect 26450 58560 26550 58690
rect 26700 58560 26800 58690
rect 26950 58560 27050 58690
rect 27200 58560 27300 58690
rect 27450 58560 27550 58690
rect 27700 58560 27800 58690
rect 27950 58560 28050 58690
rect 28200 58560 28300 58690
rect 28450 58560 28550 58690
rect 28700 58560 28800 58690
rect 28950 58560 29000 58690
rect 7000 58550 7060 58560
rect 7190 58550 7310 58560
rect 7440 58550 7560 58560
rect 7690 58550 7810 58560
rect 7940 58550 8060 58560
rect 8190 58550 8310 58560
rect 8440 58550 8560 58560
rect 8690 58550 8810 58560
rect 8940 58550 9060 58560
rect 9190 58550 9310 58560
rect 9440 58550 9560 58560
rect 9690 58550 9810 58560
rect 9940 58550 10060 58560
rect 10190 58550 10310 58560
rect 10440 58550 10560 58560
rect 10690 58550 10810 58560
rect 10940 58550 11060 58560
rect 11190 58550 11310 58560
rect 11440 58550 11560 58560
rect 11690 58550 11810 58560
rect 11940 58550 12060 58560
rect 12190 58550 12310 58560
rect 12440 58550 12560 58560
rect 12690 58550 12810 58560
rect 12940 58550 13060 58560
rect 13190 58550 13310 58560
rect 13440 58550 13560 58560
rect 13690 58550 13810 58560
rect 13940 58550 14060 58560
rect 14190 58550 14310 58560
rect 14440 58550 14560 58560
rect 14690 58550 14810 58560
rect 14940 58550 15060 58560
rect 15190 58550 15310 58560
rect 15440 58550 15560 58560
rect 15690 58550 15810 58560
rect 15940 58550 16060 58560
rect 16190 58550 16310 58560
rect 16440 58550 16560 58560
rect 16690 58550 16810 58560
rect 16940 58550 17060 58560
rect 17190 58550 17310 58560
rect 17440 58550 17560 58560
rect 17690 58550 17810 58560
rect 17940 58550 18060 58560
rect 18190 58550 18310 58560
rect 18440 58550 18560 58560
rect 18690 58550 18810 58560
rect 18940 58550 19060 58560
rect 19190 58550 19310 58560
rect 19440 58550 19560 58560
rect 19690 58550 19810 58560
rect 19940 58550 20060 58560
rect 20190 58550 20310 58560
rect 20440 58550 20560 58560
rect 20690 58550 20810 58560
rect 20940 58550 21060 58560
rect 21190 58550 21310 58560
rect 21440 58550 21560 58560
rect 21690 58550 21810 58560
rect 21940 58550 22060 58560
rect 22190 58550 22310 58560
rect 22440 58550 22560 58560
rect 22690 58550 22810 58560
rect 22940 58550 23060 58560
rect 23190 58550 23310 58560
rect 23440 58550 23560 58560
rect 23690 58550 23810 58560
rect 23940 58550 24060 58560
rect 24190 58550 24310 58560
rect 24440 58550 24560 58560
rect 24690 58550 24810 58560
rect 24940 58550 25060 58560
rect 25190 58550 25310 58560
rect 25440 58550 25560 58560
rect 25690 58550 25810 58560
rect 25940 58550 26060 58560
rect 26190 58550 26310 58560
rect 26440 58550 26560 58560
rect 26690 58550 26810 58560
rect 26940 58550 27060 58560
rect 27190 58550 27310 58560
rect 27440 58550 27560 58560
rect 27690 58550 27810 58560
rect 27940 58550 28060 58560
rect 28190 58550 28310 58560
rect 28440 58550 28560 58560
rect 28690 58550 28810 58560
rect 28940 58550 29000 58560
rect 7000 58450 29000 58550
rect 7000 58440 7060 58450
rect 7190 58440 7310 58450
rect 7440 58440 7560 58450
rect 7690 58440 7810 58450
rect 7940 58440 8060 58450
rect 8190 58440 8310 58450
rect 8440 58440 8560 58450
rect 8690 58440 8810 58450
rect 8940 58440 9060 58450
rect 9190 58440 9310 58450
rect 9440 58440 9560 58450
rect 9690 58440 9810 58450
rect 9940 58440 10060 58450
rect 10190 58440 10310 58450
rect 10440 58440 10560 58450
rect 10690 58440 10810 58450
rect 10940 58440 11060 58450
rect 11190 58440 11310 58450
rect 11440 58440 11560 58450
rect 11690 58440 11810 58450
rect 11940 58440 12060 58450
rect 12190 58440 12310 58450
rect 12440 58440 12560 58450
rect 12690 58440 12810 58450
rect 12940 58440 13060 58450
rect 13190 58440 13310 58450
rect 13440 58440 13560 58450
rect 13690 58440 13810 58450
rect 13940 58440 14060 58450
rect 14190 58440 14310 58450
rect 14440 58440 14560 58450
rect 14690 58440 14810 58450
rect 14940 58440 15060 58450
rect 15190 58440 15310 58450
rect 15440 58440 15560 58450
rect 15690 58440 15810 58450
rect 15940 58440 16060 58450
rect 16190 58440 16310 58450
rect 16440 58440 16560 58450
rect 16690 58440 16810 58450
rect 16940 58440 17060 58450
rect 17190 58440 17310 58450
rect 17440 58440 17560 58450
rect 17690 58440 17810 58450
rect 17940 58440 18060 58450
rect 18190 58440 18310 58450
rect 18440 58440 18560 58450
rect 18690 58440 18810 58450
rect 18940 58440 19060 58450
rect 19190 58440 19310 58450
rect 19440 58440 19560 58450
rect 19690 58440 19810 58450
rect 19940 58440 20060 58450
rect 20190 58440 20310 58450
rect 20440 58440 20560 58450
rect 20690 58440 20810 58450
rect 20940 58440 21060 58450
rect 21190 58440 21310 58450
rect 21440 58440 21560 58450
rect 21690 58440 21810 58450
rect 21940 58440 22060 58450
rect 22190 58440 22310 58450
rect 22440 58440 22560 58450
rect 22690 58440 22810 58450
rect 22940 58440 23060 58450
rect 23190 58440 23310 58450
rect 23440 58440 23560 58450
rect 23690 58440 23810 58450
rect 23940 58440 24060 58450
rect 24190 58440 24310 58450
rect 24440 58440 24560 58450
rect 24690 58440 24810 58450
rect 24940 58440 25060 58450
rect 25190 58440 25310 58450
rect 25440 58440 25560 58450
rect 25690 58440 25810 58450
rect 25940 58440 26060 58450
rect 26190 58440 26310 58450
rect 26440 58440 26560 58450
rect 26690 58440 26810 58450
rect 26940 58440 27060 58450
rect 27190 58440 27310 58450
rect 27440 58440 27560 58450
rect 27690 58440 27810 58450
rect 27940 58440 28060 58450
rect 28190 58440 28310 58450
rect 28440 58440 28560 58450
rect 28690 58440 28810 58450
rect 28940 58440 29000 58450
rect 7000 58310 7050 58440
rect 7200 58310 7300 58440
rect 7450 58310 7550 58440
rect 7700 58310 7800 58440
rect 7950 58310 8050 58440
rect 8200 58310 8300 58440
rect 8450 58310 8550 58440
rect 8700 58310 8800 58440
rect 8950 58310 9050 58440
rect 9200 58310 9300 58440
rect 9450 58310 9550 58440
rect 9700 58310 9800 58440
rect 9950 58310 10050 58440
rect 10200 58310 10300 58440
rect 10450 58310 10550 58440
rect 10700 58310 10800 58440
rect 10950 58310 11050 58440
rect 11200 58310 11300 58440
rect 11450 58310 11550 58440
rect 11700 58310 11800 58440
rect 11950 58310 12050 58440
rect 12200 58310 12300 58440
rect 12450 58310 12550 58440
rect 12700 58310 12800 58440
rect 12950 58310 13050 58440
rect 13200 58310 13300 58440
rect 13450 58310 13550 58440
rect 13700 58310 13800 58440
rect 13950 58310 14050 58440
rect 14200 58310 14300 58440
rect 14450 58310 14550 58440
rect 14700 58310 14800 58440
rect 14950 58310 15050 58440
rect 15200 58310 15300 58440
rect 15450 58310 15550 58440
rect 15700 58310 15800 58440
rect 15950 58310 16050 58440
rect 16200 58310 16300 58440
rect 16450 58310 16550 58440
rect 16700 58310 16800 58440
rect 16950 58310 17050 58440
rect 17200 58310 17300 58440
rect 17450 58310 17550 58440
rect 17700 58310 17800 58440
rect 17950 58310 18050 58440
rect 18200 58310 18300 58440
rect 18450 58310 18550 58440
rect 18700 58310 18800 58440
rect 18950 58310 19050 58440
rect 19200 58310 19300 58440
rect 19450 58310 19550 58440
rect 19700 58310 19800 58440
rect 19950 58310 20050 58440
rect 20200 58310 20300 58440
rect 20450 58310 20550 58440
rect 20700 58310 20800 58440
rect 20950 58310 21050 58440
rect 21200 58310 21300 58440
rect 21450 58310 21550 58440
rect 21700 58310 21800 58440
rect 21950 58310 22050 58440
rect 22200 58310 22300 58440
rect 22450 58310 22550 58440
rect 22700 58310 22800 58440
rect 22950 58310 23050 58440
rect 23200 58310 23300 58440
rect 23450 58310 23550 58440
rect 23700 58310 23800 58440
rect 23950 58310 24050 58440
rect 24200 58310 24300 58440
rect 24450 58310 24550 58440
rect 24700 58310 24800 58440
rect 24950 58310 25050 58440
rect 25200 58310 25300 58440
rect 25450 58310 25550 58440
rect 25700 58310 25800 58440
rect 25950 58310 26050 58440
rect 26200 58310 26300 58440
rect 26450 58310 26550 58440
rect 26700 58310 26800 58440
rect 26950 58310 27050 58440
rect 27200 58310 27300 58440
rect 27450 58310 27550 58440
rect 27700 58310 27800 58440
rect 27950 58310 28050 58440
rect 28200 58310 28300 58440
rect 28450 58310 28550 58440
rect 28700 58310 28800 58440
rect 28950 58310 29000 58440
rect 7000 58300 7060 58310
rect 7190 58300 7310 58310
rect 7440 58300 7560 58310
rect 7690 58300 7810 58310
rect 7940 58300 8060 58310
rect 8190 58300 8310 58310
rect 8440 58300 8560 58310
rect 8690 58300 8810 58310
rect 8940 58300 9060 58310
rect 9190 58300 9310 58310
rect 9440 58300 9560 58310
rect 9690 58300 9810 58310
rect 9940 58300 10060 58310
rect 10190 58300 10310 58310
rect 10440 58300 10560 58310
rect 10690 58300 10810 58310
rect 10940 58300 11060 58310
rect 11190 58300 11310 58310
rect 11440 58300 11560 58310
rect 11690 58300 11810 58310
rect 11940 58300 12060 58310
rect 12190 58300 12310 58310
rect 12440 58300 12560 58310
rect 12690 58300 12810 58310
rect 12940 58300 13060 58310
rect 13190 58300 13310 58310
rect 13440 58300 13560 58310
rect 13690 58300 13810 58310
rect 13940 58300 14060 58310
rect 14190 58300 14310 58310
rect 14440 58300 14560 58310
rect 14690 58300 14810 58310
rect 14940 58300 15060 58310
rect 15190 58300 15310 58310
rect 15440 58300 15560 58310
rect 15690 58300 15810 58310
rect 15940 58300 16060 58310
rect 16190 58300 16310 58310
rect 16440 58300 16560 58310
rect 16690 58300 16810 58310
rect 16940 58300 17060 58310
rect 17190 58300 17310 58310
rect 17440 58300 17560 58310
rect 17690 58300 17810 58310
rect 17940 58300 18060 58310
rect 18190 58300 18310 58310
rect 18440 58300 18560 58310
rect 18690 58300 18810 58310
rect 18940 58300 19060 58310
rect 19190 58300 19310 58310
rect 19440 58300 19560 58310
rect 19690 58300 19810 58310
rect 19940 58300 20060 58310
rect 20190 58300 20310 58310
rect 20440 58300 20560 58310
rect 20690 58300 20810 58310
rect 20940 58300 21060 58310
rect 21190 58300 21310 58310
rect 21440 58300 21560 58310
rect 21690 58300 21810 58310
rect 21940 58300 22060 58310
rect 22190 58300 22310 58310
rect 22440 58300 22560 58310
rect 22690 58300 22810 58310
rect 22940 58300 23060 58310
rect 23190 58300 23310 58310
rect 23440 58300 23560 58310
rect 23690 58300 23810 58310
rect 23940 58300 24060 58310
rect 24190 58300 24310 58310
rect 24440 58300 24560 58310
rect 24690 58300 24810 58310
rect 24940 58300 25060 58310
rect 25190 58300 25310 58310
rect 25440 58300 25560 58310
rect 25690 58300 25810 58310
rect 25940 58300 26060 58310
rect 26190 58300 26310 58310
rect 26440 58300 26560 58310
rect 26690 58300 26810 58310
rect 26940 58300 27060 58310
rect 27190 58300 27310 58310
rect 27440 58300 27560 58310
rect 27690 58300 27810 58310
rect 27940 58300 28060 58310
rect 28190 58300 28310 58310
rect 28440 58300 28560 58310
rect 28690 58300 28810 58310
rect 28940 58300 29000 58310
rect 7000 58200 29000 58300
rect 7000 58190 7060 58200
rect 7190 58190 7310 58200
rect 7440 58190 7560 58200
rect 7690 58190 7810 58200
rect 7940 58190 8060 58200
rect 8190 58190 8310 58200
rect 8440 58190 8560 58200
rect 8690 58190 8810 58200
rect 8940 58190 9060 58200
rect 9190 58190 9310 58200
rect 9440 58190 9560 58200
rect 9690 58190 9810 58200
rect 9940 58190 10060 58200
rect 10190 58190 10310 58200
rect 10440 58190 10560 58200
rect 10690 58190 10810 58200
rect 10940 58190 11060 58200
rect 11190 58190 11310 58200
rect 11440 58190 11560 58200
rect 11690 58190 11810 58200
rect 11940 58190 12060 58200
rect 12190 58190 12310 58200
rect 12440 58190 12560 58200
rect 12690 58190 12810 58200
rect 12940 58190 13060 58200
rect 13190 58190 13310 58200
rect 13440 58190 13560 58200
rect 13690 58190 13810 58200
rect 13940 58190 14060 58200
rect 14190 58190 14310 58200
rect 14440 58190 14560 58200
rect 14690 58190 14810 58200
rect 14940 58190 15060 58200
rect 15190 58190 15310 58200
rect 15440 58190 15560 58200
rect 15690 58190 15810 58200
rect 15940 58190 16060 58200
rect 16190 58190 16310 58200
rect 16440 58190 16560 58200
rect 16690 58190 16810 58200
rect 16940 58190 17060 58200
rect 17190 58190 17310 58200
rect 17440 58190 17560 58200
rect 17690 58190 17810 58200
rect 17940 58190 18060 58200
rect 18190 58190 18310 58200
rect 18440 58190 18560 58200
rect 18690 58190 18810 58200
rect 18940 58190 19060 58200
rect 19190 58190 19310 58200
rect 19440 58190 19560 58200
rect 19690 58190 19810 58200
rect 19940 58190 20060 58200
rect 20190 58190 20310 58200
rect 20440 58190 20560 58200
rect 20690 58190 20810 58200
rect 20940 58190 21060 58200
rect 21190 58190 21310 58200
rect 21440 58190 21560 58200
rect 21690 58190 21810 58200
rect 21940 58190 22060 58200
rect 22190 58190 22310 58200
rect 22440 58190 22560 58200
rect 22690 58190 22810 58200
rect 22940 58190 23060 58200
rect 23190 58190 23310 58200
rect 23440 58190 23560 58200
rect 23690 58190 23810 58200
rect 23940 58190 24060 58200
rect 24190 58190 24310 58200
rect 24440 58190 24560 58200
rect 24690 58190 24810 58200
rect 24940 58190 25060 58200
rect 25190 58190 25310 58200
rect 25440 58190 25560 58200
rect 25690 58190 25810 58200
rect 25940 58190 26060 58200
rect 26190 58190 26310 58200
rect 26440 58190 26560 58200
rect 26690 58190 26810 58200
rect 26940 58190 27060 58200
rect 27190 58190 27310 58200
rect 27440 58190 27560 58200
rect 27690 58190 27810 58200
rect 27940 58190 28060 58200
rect 28190 58190 28310 58200
rect 28440 58190 28560 58200
rect 28690 58190 28810 58200
rect 28940 58190 29000 58200
rect 7000 58060 7050 58190
rect 7200 58060 7300 58190
rect 7450 58060 7550 58190
rect 7700 58060 7800 58190
rect 7950 58060 8050 58190
rect 8200 58060 8300 58190
rect 8450 58060 8550 58190
rect 8700 58060 8800 58190
rect 8950 58060 9050 58190
rect 9200 58060 9300 58190
rect 9450 58060 9550 58190
rect 9700 58060 9800 58190
rect 9950 58060 10050 58190
rect 10200 58060 10300 58190
rect 10450 58060 10550 58190
rect 10700 58060 10800 58190
rect 10950 58060 11050 58190
rect 11200 58060 11300 58190
rect 11450 58060 11550 58190
rect 11700 58060 11800 58190
rect 11950 58060 12050 58190
rect 12200 58060 12300 58190
rect 12450 58060 12550 58190
rect 12700 58060 12800 58190
rect 12950 58060 13050 58190
rect 13200 58060 13300 58190
rect 13450 58060 13550 58190
rect 13700 58060 13800 58190
rect 13950 58060 14050 58190
rect 14200 58060 14300 58190
rect 14450 58060 14550 58190
rect 14700 58060 14800 58190
rect 14950 58060 15050 58190
rect 15200 58060 15300 58190
rect 15450 58060 15550 58190
rect 15700 58060 15800 58190
rect 15950 58060 16050 58190
rect 16200 58060 16300 58190
rect 16450 58060 16550 58190
rect 16700 58060 16800 58190
rect 16950 58060 17050 58190
rect 17200 58060 17300 58190
rect 17450 58060 17550 58190
rect 17700 58060 17800 58190
rect 17950 58060 18050 58190
rect 18200 58060 18300 58190
rect 18450 58060 18550 58190
rect 18700 58060 18800 58190
rect 18950 58060 19050 58190
rect 19200 58060 19300 58190
rect 19450 58060 19550 58190
rect 19700 58060 19800 58190
rect 19950 58060 20050 58190
rect 20200 58060 20300 58190
rect 20450 58060 20550 58190
rect 20700 58060 20800 58190
rect 20950 58060 21050 58190
rect 21200 58060 21300 58190
rect 21450 58060 21550 58190
rect 21700 58060 21800 58190
rect 21950 58060 22050 58190
rect 22200 58060 22300 58190
rect 22450 58060 22550 58190
rect 22700 58060 22800 58190
rect 22950 58060 23050 58190
rect 23200 58060 23300 58190
rect 23450 58060 23550 58190
rect 23700 58060 23800 58190
rect 23950 58060 24050 58190
rect 24200 58060 24300 58190
rect 24450 58060 24550 58190
rect 24700 58060 24800 58190
rect 24950 58060 25050 58190
rect 25200 58060 25300 58190
rect 25450 58060 25550 58190
rect 25700 58060 25800 58190
rect 25950 58060 26050 58190
rect 26200 58060 26300 58190
rect 26450 58060 26550 58190
rect 26700 58060 26800 58190
rect 26950 58060 27050 58190
rect 27200 58060 27300 58190
rect 27450 58060 27550 58190
rect 27700 58060 27800 58190
rect 27950 58060 28050 58190
rect 28200 58060 28300 58190
rect 28450 58060 28550 58190
rect 28700 58060 28800 58190
rect 28950 58060 29000 58190
rect 7000 58050 7060 58060
rect 7190 58050 7310 58060
rect 7440 58050 7560 58060
rect 7690 58050 7810 58060
rect 7940 58050 8060 58060
rect 8190 58050 8310 58060
rect 8440 58050 8560 58060
rect 8690 58050 8810 58060
rect 8940 58050 9060 58060
rect 9190 58050 9310 58060
rect 9440 58050 9560 58060
rect 9690 58050 9810 58060
rect 9940 58050 10060 58060
rect 10190 58050 10310 58060
rect 10440 58050 10560 58060
rect 10690 58050 10810 58060
rect 10940 58050 11060 58060
rect 11190 58050 11310 58060
rect 11440 58050 11560 58060
rect 11690 58050 11810 58060
rect 11940 58050 12060 58060
rect 12190 58050 12310 58060
rect 12440 58050 12560 58060
rect 12690 58050 12810 58060
rect 12940 58050 13060 58060
rect 13190 58050 13310 58060
rect 13440 58050 13560 58060
rect 13690 58050 13810 58060
rect 13940 58050 14060 58060
rect 14190 58050 14310 58060
rect 14440 58050 14560 58060
rect 14690 58050 14810 58060
rect 14940 58050 15060 58060
rect 15190 58050 15310 58060
rect 15440 58050 15560 58060
rect 15690 58050 15810 58060
rect 15940 58050 16060 58060
rect 16190 58050 16310 58060
rect 16440 58050 16560 58060
rect 16690 58050 16810 58060
rect 16940 58050 17060 58060
rect 17190 58050 17310 58060
rect 17440 58050 17560 58060
rect 17690 58050 17810 58060
rect 17940 58050 18060 58060
rect 18190 58050 18310 58060
rect 18440 58050 18560 58060
rect 18690 58050 18810 58060
rect 18940 58050 19060 58060
rect 19190 58050 19310 58060
rect 19440 58050 19560 58060
rect 19690 58050 19810 58060
rect 19940 58050 20060 58060
rect 20190 58050 20310 58060
rect 20440 58050 20560 58060
rect 20690 58050 20810 58060
rect 20940 58050 21060 58060
rect 21190 58050 21310 58060
rect 21440 58050 21560 58060
rect 21690 58050 21810 58060
rect 21940 58050 22060 58060
rect 22190 58050 22310 58060
rect 22440 58050 22560 58060
rect 22690 58050 22810 58060
rect 22940 58050 23060 58060
rect 23190 58050 23310 58060
rect 23440 58050 23560 58060
rect 23690 58050 23810 58060
rect 23940 58050 24060 58060
rect 24190 58050 24310 58060
rect 24440 58050 24560 58060
rect 24690 58050 24810 58060
rect 24940 58050 25060 58060
rect 25190 58050 25310 58060
rect 25440 58050 25560 58060
rect 25690 58050 25810 58060
rect 25940 58050 26060 58060
rect 26190 58050 26310 58060
rect 26440 58050 26560 58060
rect 26690 58050 26810 58060
rect 26940 58050 27060 58060
rect 27190 58050 27310 58060
rect 27440 58050 27560 58060
rect 27690 58050 27810 58060
rect 27940 58050 28060 58060
rect 28190 58050 28310 58060
rect 28440 58050 28560 58060
rect 28690 58050 28810 58060
rect 28940 58050 29000 58060
rect 7000 57950 29000 58050
rect 7000 57940 7060 57950
rect 7190 57940 7310 57950
rect 7440 57940 7560 57950
rect 7690 57940 7810 57950
rect 7940 57940 8060 57950
rect 8190 57940 8310 57950
rect 8440 57940 8560 57950
rect 8690 57940 8810 57950
rect 8940 57940 9060 57950
rect 9190 57940 9310 57950
rect 9440 57940 9560 57950
rect 9690 57940 9810 57950
rect 9940 57940 10060 57950
rect 10190 57940 10310 57950
rect 10440 57940 10560 57950
rect 10690 57940 10810 57950
rect 10940 57940 11060 57950
rect 11190 57940 11310 57950
rect 11440 57940 11560 57950
rect 11690 57940 11810 57950
rect 11940 57940 12060 57950
rect 12190 57940 12310 57950
rect 12440 57940 12560 57950
rect 12690 57940 12810 57950
rect 12940 57940 13060 57950
rect 13190 57940 13310 57950
rect 13440 57940 13560 57950
rect 13690 57940 13810 57950
rect 13940 57940 14060 57950
rect 14190 57940 14310 57950
rect 14440 57940 14560 57950
rect 14690 57940 14810 57950
rect 14940 57940 15060 57950
rect 15190 57940 15310 57950
rect 15440 57940 15560 57950
rect 15690 57940 15810 57950
rect 15940 57940 16060 57950
rect 16190 57940 16310 57950
rect 16440 57940 16560 57950
rect 16690 57940 16810 57950
rect 16940 57940 17060 57950
rect 17190 57940 17310 57950
rect 17440 57940 17560 57950
rect 17690 57940 17810 57950
rect 17940 57940 18060 57950
rect 18190 57940 18310 57950
rect 18440 57940 18560 57950
rect 18690 57940 18810 57950
rect 18940 57940 19060 57950
rect 19190 57940 19310 57950
rect 19440 57940 19560 57950
rect 19690 57940 19810 57950
rect 19940 57940 20060 57950
rect 20190 57940 20310 57950
rect 20440 57940 20560 57950
rect 20690 57940 20810 57950
rect 20940 57940 21060 57950
rect 21190 57940 21310 57950
rect 21440 57940 21560 57950
rect 21690 57940 21810 57950
rect 21940 57940 22060 57950
rect 22190 57940 22310 57950
rect 22440 57940 22560 57950
rect 22690 57940 22810 57950
rect 22940 57940 23060 57950
rect 23190 57940 23310 57950
rect 23440 57940 23560 57950
rect 23690 57940 23810 57950
rect 23940 57940 24060 57950
rect 24190 57940 24310 57950
rect 24440 57940 24560 57950
rect 24690 57940 24810 57950
rect 24940 57940 25060 57950
rect 25190 57940 25310 57950
rect 25440 57940 25560 57950
rect 25690 57940 25810 57950
rect 25940 57940 26060 57950
rect 26190 57940 26310 57950
rect 26440 57940 26560 57950
rect 26690 57940 26810 57950
rect 26940 57940 27060 57950
rect 27190 57940 27310 57950
rect 27440 57940 27560 57950
rect 27690 57940 27810 57950
rect 27940 57940 28060 57950
rect 28190 57940 28310 57950
rect 28440 57940 28560 57950
rect 28690 57940 28810 57950
rect 28940 57940 29000 57950
rect 7000 57810 7050 57940
rect 7200 57810 7300 57940
rect 7450 57810 7550 57940
rect 7700 57810 7800 57940
rect 7950 57810 8050 57940
rect 8200 57810 8300 57940
rect 8450 57810 8550 57940
rect 8700 57810 8800 57940
rect 8950 57810 9050 57940
rect 9200 57810 9300 57940
rect 9450 57810 9550 57940
rect 9700 57810 9800 57940
rect 9950 57810 10050 57940
rect 10200 57810 10300 57940
rect 10450 57810 10550 57940
rect 10700 57810 10800 57940
rect 10950 57810 11050 57940
rect 11200 57810 11300 57940
rect 11450 57810 11550 57940
rect 11700 57810 11800 57940
rect 11950 57810 12050 57940
rect 12200 57810 12300 57940
rect 12450 57810 12550 57940
rect 12700 57810 12800 57940
rect 12950 57810 13050 57940
rect 13200 57810 13300 57940
rect 13450 57810 13550 57940
rect 13700 57810 13800 57940
rect 13950 57810 14050 57940
rect 14200 57810 14300 57940
rect 14450 57810 14550 57940
rect 14700 57810 14800 57940
rect 14950 57810 15050 57940
rect 15200 57810 15300 57940
rect 15450 57810 15550 57940
rect 15700 57810 15800 57940
rect 15950 57810 16050 57940
rect 16200 57810 16300 57940
rect 16450 57810 16550 57940
rect 16700 57810 16800 57940
rect 16950 57810 17050 57940
rect 17200 57810 17300 57940
rect 17450 57810 17550 57940
rect 17700 57810 17800 57940
rect 17950 57810 18050 57940
rect 18200 57810 18300 57940
rect 18450 57810 18550 57940
rect 18700 57810 18800 57940
rect 18950 57810 19050 57940
rect 19200 57810 19300 57940
rect 19450 57810 19550 57940
rect 19700 57810 19800 57940
rect 19950 57810 20050 57940
rect 20200 57810 20300 57940
rect 20450 57810 20550 57940
rect 20700 57810 20800 57940
rect 20950 57810 21050 57940
rect 21200 57810 21300 57940
rect 21450 57810 21550 57940
rect 21700 57810 21800 57940
rect 21950 57810 22050 57940
rect 22200 57810 22300 57940
rect 22450 57810 22550 57940
rect 22700 57810 22800 57940
rect 22950 57810 23050 57940
rect 23200 57810 23300 57940
rect 23450 57810 23550 57940
rect 23700 57810 23800 57940
rect 23950 57810 24050 57940
rect 24200 57810 24300 57940
rect 24450 57810 24550 57940
rect 24700 57810 24800 57940
rect 24950 57810 25050 57940
rect 25200 57810 25300 57940
rect 25450 57810 25550 57940
rect 25700 57810 25800 57940
rect 25950 57810 26050 57940
rect 26200 57810 26300 57940
rect 26450 57810 26550 57940
rect 26700 57810 26800 57940
rect 26950 57810 27050 57940
rect 27200 57810 27300 57940
rect 27450 57810 27550 57940
rect 27700 57810 27800 57940
rect 27950 57810 28050 57940
rect 28200 57810 28300 57940
rect 28450 57810 28550 57940
rect 28700 57810 28800 57940
rect 28950 57810 29000 57940
rect 7000 57800 7060 57810
rect 7190 57800 7310 57810
rect 7440 57800 7560 57810
rect 7690 57800 7810 57810
rect 7940 57800 8060 57810
rect 8190 57800 8310 57810
rect 8440 57800 8560 57810
rect 8690 57800 8810 57810
rect 8940 57800 9060 57810
rect 9190 57800 9310 57810
rect 9440 57800 9560 57810
rect 9690 57800 9810 57810
rect 9940 57800 10060 57810
rect 10190 57800 10310 57810
rect 10440 57800 10560 57810
rect 10690 57800 10810 57810
rect 10940 57800 11060 57810
rect 11190 57800 11310 57810
rect 11440 57800 11560 57810
rect 11690 57800 11810 57810
rect 11940 57800 12060 57810
rect 12190 57800 12310 57810
rect 12440 57800 12560 57810
rect 12690 57800 12810 57810
rect 12940 57800 13060 57810
rect 13190 57800 13310 57810
rect 13440 57800 13560 57810
rect 13690 57800 13810 57810
rect 13940 57800 14060 57810
rect 14190 57800 14310 57810
rect 14440 57800 14560 57810
rect 14690 57800 14810 57810
rect 14940 57800 15060 57810
rect 15190 57800 15310 57810
rect 15440 57800 15560 57810
rect 15690 57800 15810 57810
rect 15940 57800 16060 57810
rect 16190 57800 16310 57810
rect 16440 57800 16560 57810
rect 16690 57800 16810 57810
rect 16940 57800 17060 57810
rect 17190 57800 17310 57810
rect 17440 57800 17560 57810
rect 17690 57800 17810 57810
rect 17940 57800 18060 57810
rect 18190 57800 18310 57810
rect 18440 57800 18560 57810
rect 18690 57800 18810 57810
rect 18940 57800 19060 57810
rect 19190 57800 19310 57810
rect 19440 57800 19560 57810
rect 19690 57800 19810 57810
rect 19940 57800 20060 57810
rect 20190 57800 20310 57810
rect 20440 57800 20560 57810
rect 20690 57800 20810 57810
rect 20940 57800 21060 57810
rect 21190 57800 21310 57810
rect 21440 57800 21560 57810
rect 21690 57800 21810 57810
rect 21940 57800 22060 57810
rect 22190 57800 22310 57810
rect 22440 57800 22560 57810
rect 22690 57800 22810 57810
rect 22940 57800 23060 57810
rect 23190 57800 23310 57810
rect 23440 57800 23560 57810
rect 23690 57800 23810 57810
rect 23940 57800 24060 57810
rect 24190 57800 24310 57810
rect 24440 57800 24560 57810
rect 24690 57800 24810 57810
rect 24940 57800 25060 57810
rect 25190 57800 25310 57810
rect 25440 57800 25560 57810
rect 25690 57800 25810 57810
rect 25940 57800 26060 57810
rect 26190 57800 26310 57810
rect 26440 57800 26560 57810
rect 26690 57800 26810 57810
rect 26940 57800 27060 57810
rect 27190 57800 27310 57810
rect 27440 57800 27560 57810
rect 27690 57800 27810 57810
rect 27940 57800 28060 57810
rect 28190 57800 28310 57810
rect 28440 57800 28560 57810
rect 28690 57800 28810 57810
rect 28940 57800 29000 57810
rect 7000 57700 29000 57800
rect 7000 57690 7060 57700
rect 7190 57690 7310 57700
rect 7440 57690 7560 57700
rect 7690 57690 7810 57700
rect 7940 57690 8060 57700
rect 8190 57690 8310 57700
rect 8440 57690 8560 57700
rect 8690 57690 8810 57700
rect 8940 57690 9060 57700
rect 9190 57690 9310 57700
rect 9440 57690 9560 57700
rect 9690 57690 9810 57700
rect 9940 57690 10060 57700
rect 10190 57690 10310 57700
rect 10440 57690 10560 57700
rect 10690 57690 10810 57700
rect 10940 57690 11060 57700
rect 11190 57690 11310 57700
rect 11440 57690 11560 57700
rect 11690 57690 11810 57700
rect 11940 57690 12060 57700
rect 12190 57690 12310 57700
rect 12440 57690 12560 57700
rect 12690 57690 12810 57700
rect 12940 57690 13060 57700
rect 13190 57690 13310 57700
rect 13440 57690 13560 57700
rect 13690 57690 13810 57700
rect 13940 57690 14060 57700
rect 14190 57690 14310 57700
rect 14440 57690 14560 57700
rect 14690 57690 14810 57700
rect 14940 57690 15060 57700
rect 15190 57690 15310 57700
rect 15440 57690 15560 57700
rect 15690 57690 15810 57700
rect 15940 57690 16060 57700
rect 16190 57690 16310 57700
rect 16440 57690 16560 57700
rect 16690 57690 16810 57700
rect 16940 57690 17060 57700
rect 17190 57690 17310 57700
rect 17440 57690 17560 57700
rect 17690 57690 17810 57700
rect 17940 57690 18060 57700
rect 18190 57690 18310 57700
rect 18440 57690 18560 57700
rect 18690 57690 18810 57700
rect 18940 57690 19060 57700
rect 19190 57690 19310 57700
rect 19440 57690 19560 57700
rect 19690 57690 19810 57700
rect 19940 57690 20060 57700
rect 20190 57690 20310 57700
rect 20440 57690 20560 57700
rect 20690 57690 20810 57700
rect 20940 57690 21060 57700
rect 21190 57690 21310 57700
rect 21440 57690 21560 57700
rect 21690 57690 21810 57700
rect 21940 57690 22060 57700
rect 22190 57690 22310 57700
rect 22440 57690 22560 57700
rect 22690 57690 22810 57700
rect 22940 57690 23060 57700
rect 23190 57690 23310 57700
rect 23440 57690 23560 57700
rect 23690 57690 23810 57700
rect 23940 57690 24060 57700
rect 24190 57690 24310 57700
rect 24440 57690 24560 57700
rect 24690 57690 24810 57700
rect 24940 57690 25060 57700
rect 25190 57690 25310 57700
rect 25440 57690 25560 57700
rect 25690 57690 25810 57700
rect 25940 57690 26060 57700
rect 26190 57690 26310 57700
rect 26440 57690 26560 57700
rect 26690 57690 26810 57700
rect 26940 57690 27060 57700
rect 27190 57690 27310 57700
rect 27440 57690 27560 57700
rect 27690 57690 27810 57700
rect 27940 57690 28060 57700
rect 28190 57690 28310 57700
rect 28440 57690 28560 57700
rect 28690 57690 28810 57700
rect 28940 57690 29000 57700
rect 7000 57560 7050 57690
rect 7200 57560 7300 57690
rect 7450 57560 7550 57690
rect 7700 57560 7800 57690
rect 7950 57560 8050 57690
rect 8200 57560 8300 57690
rect 8450 57560 8550 57690
rect 8700 57560 8800 57690
rect 8950 57560 9050 57690
rect 9200 57560 9300 57690
rect 9450 57560 9550 57690
rect 9700 57560 9800 57690
rect 9950 57560 10050 57690
rect 10200 57560 10300 57690
rect 10450 57560 10550 57690
rect 10700 57560 10800 57690
rect 10950 57560 11050 57690
rect 11200 57560 11300 57690
rect 11450 57560 11550 57690
rect 11700 57560 11800 57690
rect 11950 57560 12050 57690
rect 12200 57560 12300 57690
rect 12450 57560 12550 57690
rect 12700 57560 12800 57690
rect 12950 57560 13050 57690
rect 13200 57560 13300 57690
rect 13450 57560 13550 57690
rect 13700 57560 13800 57690
rect 13950 57560 14050 57690
rect 14200 57560 14300 57690
rect 14450 57560 14550 57690
rect 14700 57560 14800 57690
rect 14950 57560 15050 57690
rect 15200 57560 15300 57690
rect 15450 57560 15550 57690
rect 15700 57560 15800 57690
rect 15950 57560 16050 57690
rect 16200 57560 16300 57690
rect 16450 57560 16550 57690
rect 16700 57560 16800 57690
rect 16950 57560 17050 57690
rect 17200 57560 17300 57690
rect 17450 57560 17550 57690
rect 17700 57560 17800 57690
rect 17950 57560 18050 57690
rect 18200 57560 18300 57690
rect 18450 57560 18550 57690
rect 18700 57560 18800 57690
rect 18950 57560 19050 57690
rect 19200 57560 19300 57690
rect 19450 57560 19550 57690
rect 19700 57560 19800 57690
rect 19950 57560 20050 57690
rect 20200 57560 20300 57690
rect 20450 57560 20550 57690
rect 20700 57560 20800 57690
rect 20950 57560 21050 57690
rect 21200 57560 21300 57690
rect 21450 57560 21550 57690
rect 21700 57560 21800 57690
rect 21950 57560 22050 57690
rect 22200 57560 22300 57690
rect 22450 57560 22550 57690
rect 22700 57560 22800 57690
rect 22950 57560 23050 57690
rect 23200 57560 23300 57690
rect 23450 57560 23550 57690
rect 23700 57560 23800 57690
rect 23950 57560 24050 57690
rect 24200 57560 24300 57690
rect 24450 57560 24550 57690
rect 24700 57560 24800 57690
rect 24950 57560 25050 57690
rect 25200 57560 25300 57690
rect 25450 57560 25550 57690
rect 25700 57560 25800 57690
rect 25950 57560 26050 57690
rect 26200 57560 26300 57690
rect 26450 57560 26550 57690
rect 26700 57560 26800 57690
rect 26950 57560 27050 57690
rect 27200 57560 27300 57690
rect 27450 57560 27550 57690
rect 27700 57560 27800 57690
rect 27950 57560 28050 57690
rect 28200 57560 28300 57690
rect 28450 57560 28550 57690
rect 28700 57560 28800 57690
rect 28950 57560 29000 57690
rect 7000 57550 7060 57560
rect 7190 57550 7310 57560
rect 7440 57550 7560 57560
rect 7690 57550 7810 57560
rect 7940 57550 8060 57560
rect 8190 57550 8310 57560
rect 8440 57550 8560 57560
rect 8690 57550 8810 57560
rect 8940 57550 9060 57560
rect 9190 57550 9310 57560
rect 9440 57550 9560 57560
rect 9690 57550 9810 57560
rect 9940 57550 10060 57560
rect 10190 57550 10310 57560
rect 10440 57550 10560 57560
rect 10690 57550 10810 57560
rect 10940 57550 11060 57560
rect 11190 57550 11310 57560
rect 11440 57550 11560 57560
rect 11690 57550 11810 57560
rect 11940 57550 12060 57560
rect 12190 57550 12310 57560
rect 12440 57550 12560 57560
rect 12690 57550 12810 57560
rect 12940 57550 13060 57560
rect 13190 57550 13310 57560
rect 13440 57550 13560 57560
rect 13690 57550 13810 57560
rect 13940 57550 14060 57560
rect 14190 57550 14310 57560
rect 14440 57550 14560 57560
rect 14690 57550 14810 57560
rect 14940 57550 15060 57560
rect 15190 57550 15310 57560
rect 15440 57550 15560 57560
rect 15690 57550 15810 57560
rect 15940 57550 16060 57560
rect 16190 57550 16310 57560
rect 16440 57550 16560 57560
rect 16690 57550 16810 57560
rect 16940 57550 17060 57560
rect 17190 57550 17310 57560
rect 17440 57550 17560 57560
rect 17690 57550 17810 57560
rect 17940 57550 18060 57560
rect 18190 57550 18310 57560
rect 18440 57550 18560 57560
rect 18690 57550 18810 57560
rect 18940 57550 19060 57560
rect 19190 57550 19310 57560
rect 19440 57550 19560 57560
rect 19690 57550 19810 57560
rect 19940 57550 20060 57560
rect 20190 57550 20310 57560
rect 20440 57550 20560 57560
rect 20690 57550 20810 57560
rect 20940 57550 21060 57560
rect 21190 57550 21310 57560
rect 21440 57550 21560 57560
rect 21690 57550 21810 57560
rect 21940 57550 22060 57560
rect 22190 57550 22310 57560
rect 22440 57550 22560 57560
rect 22690 57550 22810 57560
rect 22940 57550 23060 57560
rect 23190 57550 23310 57560
rect 23440 57550 23560 57560
rect 23690 57550 23810 57560
rect 23940 57550 24060 57560
rect 24190 57550 24310 57560
rect 24440 57550 24560 57560
rect 24690 57550 24810 57560
rect 24940 57550 25060 57560
rect 25190 57550 25310 57560
rect 25440 57550 25560 57560
rect 25690 57550 25810 57560
rect 25940 57550 26060 57560
rect 26190 57550 26310 57560
rect 26440 57550 26560 57560
rect 26690 57550 26810 57560
rect 26940 57550 27060 57560
rect 27190 57550 27310 57560
rect 27440 57550 27560 57560
rect 27690 57550 27810 57560
rect 27940 57550 28060 57560
rect 28190 57550 28310 57560
rect 28440 57550 28560 57560
rect 28690 57550 28810 57560
rect 28940 57550 29000 57560
rect 7000 57450 29000 57550
rect 7000 57440 7060 57450
rect 7190 57440 7310 57450
rect 7440 57440 7560 57450
rect 7690 57440 7810 57450
rect 7940 57440 8060 57450
rect 8190 57440 8310 57450
rect 8440 57440 8560 57450
rect 8690 57440 8810 57450
rect 8940 57440 9060 57450
rect 9190 57440 9310 57450
rect 9440 57440 9560 57450
rect 9690 57440 9810 57450
rect 9940 57440 10060 57450
rect 10190 57440 10310 57450
rect 10440 57440 10560 57450
rect 10690 57440 10810 57450
rect 10940 57440 11060 57450
rect 11190 57440 11310 57450
rect 11440 57440 11560 57450
rect 11690 57440 11810 57450
rect 11940 57440 12060 57450
rect 12190 57440 12310 57450
rect 12440 57440 12560 57450
rect 12690 57440 12810 57450
rect 12940 57440 13060 57450
rect 13190 57440 13310 57450
rect 13440 57440 13560 57450
rect 13690 57440 13810 57450
rect 13940 57440 14060 57450
rect 14190 57440 14310 57450
rect 14440 57440 14560 57450
rect 14690 57440 14810 57450
rect 14940 57440 15060 57450
rect 15190 57440 15310 57450
rect 15440 57440 15560 57450
rect 15690 57440 15810 57450
rect 15940 57440 16060 57450
rect 16190 57440 16310 57450
rect 16440 57440 16560 57450
rect 16690 57440 16810 57450
rect 16940 57440 17060 57450
rect 17190 57440 17310 57450
rect 17440 57440 17560 57450
rect 17690 57440 17810 57450
rect 17940 57440 18060 57450
rect 18190 57440 18310 57450
rect 18440 57440 18560 57450
rect 18690 57440 18810 57450
rect 18940 57440 19060 57450
rect 19190 57440 19310 57450
rect 19440 57440 19560 57450
rect 19690 57440 19810 57450
rect 19940 57440 20060 57450
rect 20190 57440 20310 57450
rect 20440 57440 20560 57450
rect 20690 57440 20810 57450
rect 20940 57440 21060 57450
rect 21190 57440 21310 57450
rect 21440 57440 21560 57450
rect 21690 57440 21810 57450
rect 21940 57440 22060 57450
rect 22190 57440 22310 57450
rect 22440 57440 22560 57450
rect 22690 57440 22810 57450
rect 22940 57440 23060 57450
rect 23190 57440 23310 57450
rect 23440 57440 23560 57450
rect 23690 57440 23810 57450
rect 23940 57440 24060 57450
rect 24190 57440 24310 57450
rect 24440 57440 24560 57450
rect 24690 57440 24810 57450
rect 24940 57440 25060 57450
rect 25190 57440 25310 57450
rect 25440 57440 25560 57450
rect 25690 57440 25810 57450
rect 25940 57440 26060 57450
rect 26190 57440 26310 57450
rect 26440 57440 26560 57450
rect 26690 57440 26810 57450
rect 26940 57440 27060 57450
rect 27190 57440 27310 57450
rect 27440 57440 27560 57450
rect 27690 57440 27810 57450
rect 27940 57440 28060 57450
rect 28190 57440 28310 57450
rect 28440 57440 28560 57450
rect 28690 57440 28810 57450
rect 28940 57440 29000 57450
rect 7000 57310 7050 57440
rect 7200 57310 7300 57440
rect 7450 57310 7550 57440
rect 7700 57310 7800 57440
rect 7950 57310 8050 57440
rect 8200 57310 8300 57440
rect 8450 57310 8550 57440
rect 8700 57310 8800 57440
rect 8950 57310 9050 57440
rect 9200 57310 9300 57440
rect 9450 57310 9550 57440
rect 9700 57310 9800 57440
rect 9950 57310 10050 57440
rect 10200 57310 10300 57440
rect 10450 57310 10550 57440
rect 10700 57310 10800 57440
rect 10950 57310 11050 57440
rect 11200 57310 11300 57440
rect 11450 57310 11550 57440
rect 11700 57310 11800 57440
rect 11950 57310 12050 57440
rect 12200 57310 12300 57440
rect 12450 57310 12550 57440
rect 12700 57310 12800 57440
rect 12950 57310 13050 57440
rect 13200 57310 13300 57440
rect 13450 57310 13550 57440
rect 13700 57310 13800 57440
rect 13950 57310 14050 57440
rect 14200 57310 14300 57440
rect 14450 57310 14550 57440
rect 14700 57310 14800 57440
rect 14950 57310 15050 57440
rect 15200 57310 15300 57440
rect 15450 57310 15550 57440
rect 15700 57310 15800 57440
rect 15950 57310 16050 57440
rect 16200 57310 16300 57440
rect 16450 57310 16550 57440
rect 16700 57310 16800 57440
rect 16950 57310 17050 57440
rect 17200 57310 17300 57440
rect 17450 57310 17550 57440
rect 17700 57310 17800 57440
rect 17950 57310 18050 57440
rect 18200 57310 18300 57440
rect 18450 57310 18550 57440
rect 18700 57310 18800 57440
rect 18950 57310 19050 57440
rect 19200 57310 19300 57440
rect 19450 57310 19550 57440
rect 19700 57310 19800 57440
rect 19950 57310 20050 57440
rect 20200 57310 20300 57440
rect 20450 57310 20550 57440
rect 20700 57310 20800 57440
rect 20950 57310 21050 57440
rect 21200 57310 21300 57440
rect 21450 57310 21550 57440
rect 21700 57310 21800 57440
rect 21950 57310 22050 57440
rect 22200 57310 22300 57440
rect 22450 57310 22550 57440
rect 22700 57310 22800 57440
rect 22950 57310 23050 57440
rect 23200 57310 23300 57440
rect 23450 57310 23550 57440
rect 23700 57310 23800 57440
rect 23950 57310 24050 57440
rect 24200 57310 24300 57440
rect 24450 57310 24550 57440
rect 24700 57310 24800 57440
rect 24950 57310 25050 57440
rect 25200 57310 25300 57440
rect 25450 57310 25550 57440
rect 25700 57310 25800 57440
rect 25950 57310 26050 57440
rect 26200 57310 26300 57440
rect 26450 57310 26550 57440
rect 26700 57310 26800 57440
rect 26950 57310 27050 57440
rect 27200 57310 27300 57440
rect 27450 57310 27550 57440
rect 27700 57310 27800 57440
rect 27950 57310 28050 57440
rect 28200 57310 28300 57440
rect 28450 57310 28550 57440
rect 28700 57310 28800 57440
rect 28950 57310 29000 57440
rect 7000 57300 7060 57310
rect 7190 57300 7310 57310
rect 7440 57300 7560 57310
rect 7690 57300 7810 57310
rect 7940 57300 8060 57310
rect 8190 57300 8310 57310
rect 8440 57300 8560 57310
rect 8690 57300 8810 57310
rect 8940 57300 9060 57310
rect 9190 57300 9310 57310
rect 9440 57300 9560 57310
rect 9690 57300 9810 57310
rect 9940 57300 10060 57310
rect 10190 57300 10310 57310
rect 10440 57300 10560 57310
rect 10690 57300 10810 57310
rect 10940 57300 11060 57310
rect 11190 57300 11310 57310
rect 11440 57300 11560 57310
rect 11690 57300 11810 57310
rect 11940 57300 12060 57310
rect 12190 57300 12310 57310
rect 12440 57300 12560 57310
rect 12690 57300 12810 57310
rect 12940 57300 13060 57310
rect 13190 57300 13310 57310
rect 13440 57300 13560 57310
rect 13690 57300 13810 57310
rect 13940 57300 14060 57310
rect 14190 57300 14310 57310
rect 14440 57300 14560 57310
rect 14690 57300 14810 57310
rect 14940 57300 15060 57310
rect 15190 57300 15310 57310
rect 15440 57300 15560 57310
rect 15690 57300 15810 57310
rect 15940 57300 16060 57310
rect 16190 57300 16310 57310
rect 16440 57300 16560 57310
rect 16690 57300 16810 57310
rect 16940 57300 17060 57310
rect 17190 57300 17310 57310
rect 17440 57300 17560 57310
rect 17690 57300 17810 57310
rect 17940 57300 18060 57310
rect 18190 57300 18310 57310
rect 18440 57300 18560 57310
rect 18690 57300 18810 57310
rect 18940 57300 19060 57310
rect 19190 57300 19310 57310
rect 19440 57300 19560 57310
rect 19690 57300 19810 57310
rect 19940 57300 20060 57310
rect 20190 57300 20310 57310
rect 20440 57300 20560 57310
rect 20690 57300 20810 57310
rect 20940 57300 21060 57310
rect 21190 57300 21310 57310
rect 21440 57300 21560 57310
rect 21690 57300 21810 57310
rect 21940 57300 22060 57310
rect 22190 57300 22310 57310
rect 22440 57300 22560 57310
rect 22690 57300 22810 57310
rect 22940 57300 23060 57310
rect 23190 57300 23310 57310
rect 23440 57300 23560 57310
rect 23690 57300 23810 57310
rect 23940 57300 24060 57310
rect 24190 57300 24310 57310
rect 24440 57300 24560 57310
rect 24690 57300 24810 57310
rect 24940 57300 25060 57310
rect 25190 57300 25310 57310
rect 25440 57300 25560 57310
rect 25690 57300 25810 57310
rect 25940 57300 26060 57310
rect 26190 57300 26310 57310
rect 26440 57300 26560 57310
rect 26690 57300 26810 57310
rect 26940 57300 27060 57310
rect 27190 57300 27310 57310
rect 27440 57300 27560 57310
rect 27690 57300 27810 57310
rect 27940 57300 28060 57310
rect 28190 57300 28310 57310
rect 28440 57300 28560 57310
rect 28690 57300 28810 57310
rect 28940 57300 29000 57310
rect 7000 57200 29000 57300
rect 7000 57190 7060 57200
rect 7190 57190 7310 57200
rect 7440 57190 7560 57200
rect 7690 57190 7810 57200
rect 7940 57190 8060 57200
rect 8190 57190 8310 57200
rect 8440 57190 8560 57200
rect 8690 57190 8810 57200
rect 8940 57190 9060 57200
rect 9190 57190 9310 57200
rect 9440 57190 9560 57200
rect 9690 57190 9810 57200
rect 9940 57190 10060 57200
rect 10190 57190 10310 57200
rect 10440 57190 10560 57200
rect 10690 57190 10810 57200
rect 10940 57190 11060 57200
rect 11190 57190 11310 57200
rect 11440 57190 11560 57200
rect 11690 57190 11810 57200
rect 11940 57190 12060 57200
rect 12190 57190 12310 57200
rect 12440 57190 12560 57200
rect 12690 57190 12810 57200
rect 12940 57190 13060 57200
rect 13190 57190 13310 57200
rect 13440 57190 13560 57200
rect 13690 57190 13810 57200
rect 13940 57190 14060 57200
rect 14190 57190 14310 57200
rect 14440 57190 14560 57200
rect 14690 57190 14810 57200
rect 14940 57190 15060 57200
rect 15190 57190 15310 57200
rect 15440 57190 15560 57200
rect 15690 57190 15810 57200
rect 15940 57190 16060 57200
rect 16190 57190 16310 57200
rect 16440 57190 16560 57200
rect 16690 57190 16810 57200
rect 16940 57190 17060 57200
rect 17190 57190 17310 57200
rect 17440 57190 17560 57200
rect 17690 57190 17810 57200
rect 17940 57190 18060 57200
rect 18190 57190 18310 57200
rect 18440 57190 18560 57200
rect 18690 57190 18810 57200
rect 18940 57190 19060 57200
rect 19190 57190 19310 57200
rect 19440 57190 19560 57200
rect 19690 57190 19810 57200
rect 19940 57190 20060 57200
rect 20190 57190 20310 57200
rect 20440 57190 20560 57200
rect 20690 57190 20810 57200
rect 20940 57190 21060 57200
rect 21190 57190 21310 57200
rect 21440 57190 21560 57200
rect 21690 57190 21810 57200
rect 21940 57190 22060 57200
rect 22190 57190 22310 57200
rect 22440 57190 22560 57200
rect 22690 57190 22810 57200
rect 22940 57190 23060 57200
rect 23190 57190 23310 57200
rect 23440 57190 23560 57200
rect 23690 57190 23810 57200
rect 23940 57190 24060 57200
rect 24190 57190 24310 57200
rect 24440 57190 24560 57200
rect 24690 57190 24810 57200
rect 24940 57190 25060 57200
rect 25190 57190 25310 57200
rect 25440 57190 25560 57200
rect 25690 57190 25810 57200
rect 25940 57190 26060 57200
rect 26190 57190 26310 57200
rect 26440 57190 26560 57200
rect 26690 57190 26810 57200
rect 26940 57190 27060 57200
rect 27190 57190 27310 57200
rect 27440 57190 27560 57200
rect 27690 57190 27810 57200
rect 27940 57190 28060 57200
rect 28190 57190 28310 57200
rect 28440 57190 28560 57200
rect 28690 57190 28810 57200
rect 28940 57190 29000 57200
rect 7000 57060 7050 57190
rect 7200 57060 7300 57190
rect 7450 57060 7550 57190
rect 7700 57060 7800 57190
rect 7950 57060 8050 57190
rect 8200 57060 8300 57190
rect 8450 57060 8550 57190
rect 8700 57060 8800 57190
rect 8950 57060 9050 57190
rect 9200 57060 9300 57190
rect 9450 57060 9550 57190
rect 9700 57060 9800 57190
rect 9950 57060 10050 57190
rect 10200 57060 10300 57190
rect 10450 57060 10550 57190
rect 10700 57060 10800 57190
rect 10950 57060 11050 57190
rect 11200 57060 11300 57190
rect 11450 57060 11550 57190
rect 11700 57060 11800 57190
rect 11950 57060 12050 57190
rect 12200 57060 12300 57190
rect 12450 57060 12550 57190
rect 12700 57060 12800 57190
rect 12950 57060 13050 57190
rect 13200 57060 13300 57190
rect 13450 57060 13550 57190
rect 13700 57060 13800 57190
rect 13950 57060 14050 57190
rect 14200 57060 14300 57190
rect 14450 57060 14550 57190
rect 14700 57060 14800 57190
rect 14950 57060 15050 57190
rect 15200 57060 15300 57190
rect 15450 57060 15550 57190
rect 15700 57060 15800 57190
rect 15950 57060 16050 57190
rect 16200 57060 16300 57190
rect 16450 57060 16550 57190
rect 16700 57060 16800 57190
rect 16950 57060 17050 57190
rect 17200 57060 17300 57190
rect 17450 57060 17550 57190
rect 17700 57060 17800 57190
rect 17950 57060 18050 57190
rect 18200 57060 18300 57190
rect 18450 57060 18550 57190
rect 18700 57060 18800 57190
rect 18950 57060 19050 57190
rect 19200 57060 19300 57190
rect 19450 57060 19550 57190
rect 19700 57060 19800 57190
rect 19950 57060 20050 57190
rect 20200 57060 20300 57190
rect 20450 57060 20550 57190
rect 20700 57060 20800 57190
rect 20950 57060 21050 57190
rect 21200 57060 21300 57190
rect 21450 57060 21550 57190
rect 21700 57060 21800 57190
rect 21950 57060 22050 57190
rect 22200 57060 22300 57190
rect 22450 57060 22550 57190
rect 22700 57060 22800 57190
rect 22950 57060 23050 57190
rect 23200 57060 23300 57190
rect 23450 57060 23550 57190
rect 23700 57060 23800 57190
rect 23950 57060 24050 57190
rect 24200 57060 24300 57190
rect 24450 57060 24550 57190
rect 24700 57060 24800 57190
rect 24950 57060 25050 57190
rect 25200 57060 25300 57190
rect 25450 57060 25550 57190
rect 25700 57060 25800 57190
rect 25950 57060 26050 57190
rect 26200 57060 26300 57190
rect 26450 57060 26550 57190
rect 26700 57060 26800 57190
rect 26950 57060 27050 57190
rect 27200 57060 27300 57190
rect 27450 57060 27550 57190
rect 27700 57060 27800 57190
rect 27950 57060 28050 57190
rect 28200 57060 28300 57190
rect 28450 57060 28550 57190
rect 28700 57060 28800 57190
rect 28950 57060 29000 57190
rect 7000 57050 7060 57060
rect 7190 57050 7310 57060
rect 7440 57050 7560 57060
rect 7690 57050 7810 57060
rect 7940 57050 8060 57060
rect 8190 57050 8310 57060
rect 8440 57050 8560 57060
rect 8690 57050 8810 57060
rect 8940 57050 9060 57060
rect 9190 57050 9310 57060
rect 9440 57050 9560 57060
rect 9690 57050 9810 57060
rect 9940 57050 10060 57060
rect 10190 57050 10310 57060
rect 10440 57050 10560 57060
rect 10690 57050 10810 57060
rect 10940 57050 11060 57060
rect 11190 57050 11310 57060
rect 11440 57050 11560 57060
rect 11690 57050 11810 57060
rect 11940 57050 12060 57060
rect 12190 57050 12310 57060
rect 12440 57050 12560 57060
rect 12690 57050 12810 57060
rect 12940 57050 13060 57060
rect 13190 57050 13310 57060
rect 13440 57050 13560 57060
rect 13690 57050 13810 57060
rect 13940 57050 14060 57060
rect 14190 57050 14310 57060
rect 14440 57050 14560 57060
rect 14690 57050 14810 57060
rect 14940 57050 15060 57060
rect 15190 57050 15310 57060
rect 15440 57050 15560 57060
rect 15690 57050 15810 57060
rect 15940 57050 16060 57060
rect 16190 57050 16310 57060
rect 16440 57050 16560 57060
rect 16690 57050 16810 57060
rect 16940 57050 17060 57060
rect 17190 57050 17310 57060
rect 17440 57050 17560 57060
rect 17690 57050 17810 57060
rect 17940 57050 18060 57060
rect 18190 57050 18310 57060
rect 18440 57050 18560 57060
rect 18690 57050 18810 57060
rect 18940 57050 19060 57060
rect 19190 57050 19310 57060
rect 19440 57050 19560 57060
rect 19690 57050 19810 57060
rect 19940 57050 20060 57060
rect 20190 57050 20310 57060
rect 20440 57050 20560 57060
rect 20690 57050 20810 57060
rect 20940 57050 21060 57060
rect 21190 57050 21310 57060
rect 21440 57050 21560 57060
rect 21690 57050 21810 57060
rect 21940 57050 22060 57060
rect 22190 57050 22310 57060
rect 22440 57050 22560 57060
rect 22690 57050 22810 57060
rect 22940 57050 23060 57060
rect 23190 57050 23310 57060
rect 23440 57050 23560 57060
rect 23690 57050 23810 57060
rect 23940 57050 24060 57060
rect 24190 57050 24310 57060
rect 24440 57050 24560 57060
rect 24690 57050 24810 57060
rect 24940 57050 25060 57060
rect 25190 57050 25310 57060
rect 25440 57050 25560 57060
rect 25690 57050 25810 57060
rect 25940 57050 26060 57060
rect 26190 57050 26310 57060
rect 26440 57050 26560 57060
rect 26690 57050 26810 57060
rect 26940 57050 27060 57060
rect 27190 57050 27310 57060
rect 27440 57050 27560 57060
rect 27690 57050 27810 57060
rect 27940 57050 28060 57060
rect 28190 57050 28310 57060
rect 28440 57050 28560 57060
rect 28690 57050 28810 57060
rect 28940 57050 29000 57060
rect 7000 57000 29000 57050
rect 59000 60950 71000 61000
rect 59000 60940 59060 60950
rect 59190 60940 59310 60950
rect 59440 60940 59560 60950
rect 59690 60940 59810 60950
rect 59940 60940 60060 60950
rect 60190 60940 60310 60950
rect 60440 60940 60560 60950
rect 60690 60940 60810 60950
rect 60940 60940 61060 60950
rect 61190 60940 61310 60950
rect 61440 60940 61560 60950
rect 61690 60940 61810 60950
rect 61940 60940 62060 60950
rect 62190 60940 62310 60950
rect 62440 60940 62560 60950
rect 62690 60940 62810 60950
rect 62940 60940 63060 60950
rect 63190 60940 63310 60950
rect 63440 60940 63560 60950
rect 63690 60940 63810 60950
rect 63940 60940 64060 60950
rect 64190 60940 64310 60950
rect 64440 60940 64560 60950
rect 64690 60940 64810 60950
rect 64940 60940 65060 60950
rect 65190 60940 65310 60950
rect 65440 60940 65560 60950
rect 65690 60940 65810 60950
rect 65940 60940 66060 60950
rect 66190 60940 66310 60950
rect 66440 60940 66560 60950
rect 66690 60940 66810 60950
rect 66940 60940 67060 60950
rect 67190 60940 67310 60950
rect 67440 60940 67560 60950
rect 67690 60940 67810 60950
rect 67940 60940 68060 60950
rect 68190 60940 68310 60950
rect 68440 60940 68560 60950
rect 68690 60940 68810 60950
rect 68940 60940 69060 60950
rect 69190 60940 69310 60950
rect 69440 60940 69560 60950
rect 69690 60940 69810 60950
rect 69940 60940 70060 60950
rect 70190 60940 70310 60950
rect 70440 60940 70560 60950
rect 70690 60940 70810 60950
rect 70940 60940 71000 60950
rect 59000 60810 59050 60940
rect 59200 60810 59300 60940
rect 59450 60810 59550 60940
rect 59700 60810 59800 60940
rect 59950 60810 60050 60940
rect 60200 60810 60300 60940
rect 60450 60810 60550 60940
rect 60700 60810 60800 60940
rect 60950 60810 61050 60940
rect 61200 60810 61300 60940
rect 61450 60810 61550 60940
rect 61700 60810 61800 60940
rect 61950 60810 62050 60940
rect 62200 60810 62300 60940
rect 62450 60810 62550 60940
rect 62700 60810 62800 60940
rect 62950 60810 63050 60940
rect 63200 60810 63300 60940
rect 63450 60810 63550 60940
rect 63700 60810 63800 60940
rect 63950 60810 64050 60940
rect 64200 60810 64300 60940
rect 64450 60810 64550 60940
rect 64700 60810 64800 60940
rect 64950 60810 65050 60940
rect 65200 60810 65300 60940
rect 65450 60810 65550 60940
rect 65700 60810 65800 60940
rect 65950 60810 66050 60940
rect 66200 60810 66300 60940
rect 66450 60810 66550 60940
rect 66700 60810 66800 60940
rect 66950 60810 67050 60940
rect 67200 60810 67300 60940
rect 67450 60810 67550 60940
rect 67700 60810 67800 60940
rect 67950 60810 68050 60940
rect 68200 60810 68300 60940
rect 68450 60810 68550 60940
rect 68700 60810 68800 60940
rect 68950 60810 69050 60940
rect 69200 60810 69300 60940
rect 69450 60810 69550 60940
rect 69700 60810 69800 60940
rect 69950 60810 70050 60940
rect 70200 60810 70300 60940
rect 70450 60810 70550 60940
rect 70700 60810 70800 60940
rect 70950 60810 71000 60940
rect 59000 60800 59060 60810
rect 59190 60800 59310 60810
rect 59440 60800 59560 60810
rect 59690 60800 59810 60810
rect 59940 60800 60060 60810
rect 60190 60800 60310 60810
rect 60440 60800 60560 60810
rect 60690 60800 60810 60810
rect 60940 60800 61060 60810
rect 61190 60800 61310 60810
rect 61440 60800 61560 60810
rect 61690 60800 61810 60810
rect 61940 60800 62060 60810
rect 62190 60800 62310 60810
rect 62440 60800 62560 60810
rect 62690 60800 62810 60810
rect 62940 60800 63060 60810
rect 63190 60800 63310 60810
rect 63440 60800 63560 60810
rect 63690 60800 63810 60810
rect 63940 60800 64060 60810
rect 64190 60800 64310 60810
rect 64440 60800 64560 60810
rect 64690 60800 64810 60810
rect 64940 60800 65060 60810
rect 65190 60800 65310 60810
rect 65440 60800 65560 60810
rect 65690 60800 65810 60810
rect 65940 60800 66060 60810
rect 66190 60800 66310 60810
rect 66440 60800 66560 60810
rect 66690 60800 66810 60810
rect 66940 60800 67060 60810
rect 67190 60800 67310 60810
rect 67440 60800 67560 60810
rect 67690 60800 67810 60810
rect 67940 60800 68060 60810
rect 68190 60800 68310 60810
rect 68440 60800 68560 60810
rect 68690 60800 68810 60810
rect 68940 60800 69060 60810
rect 69190 60800 69310 60810
rect 69440 60800 69560 60810
rect 69690 60800 69810 60810
rect 69940 60800 70060 60810
rect 70190 60800 70310 60810
rect 70440 60800 70560 60810
rect 70690 60800 70810 60810
rect 70940 60800 71000 60810
rect 59000 60700 71000 60800
rect 59000 60690 59060 60700
rect 59190 60690 59310 60700
rect 59440 60690 59560 60700
rect 59690 60690 59810 60700
rect 59940 60690 60060 60700
rect 60190 60690 60310 60700
rect 60440 60690 60560 60700
rect 60690 60690 60810 60700
rect 60940 60690 61060 60700
rect 61190 60690 61310 60700
rect 61440 60690 61560 60700
rect 61690 60690 61810 60700
rect 61940 60690 62060 60700
rect 62190 60690 62310 60700
rect 62440 60690 62560 60700
rect 62690 60690 62810 60700
rect 62940 60690 63060 60700
rect 63190 60690 63310 60700
rect 63440 60690 63560 60700
rect 63690 60690 63810 60700
rect 63940 60690 64060 60700
rect 64190 60690 64310 60700
rect 64440 60690 64560 60700
rect 64690 60690 64810 60700
rect 64940 60690 65060 60700
rect 65190 60690 65310 60700
rect 65440 60690 65560 60700
rect 65690 60690 65810 60700
rect 65940 60690 66060 60700
rect 66190 60690 66310 60700
rect 66440 60690 66560 60700
rect 66690 60690 66810 60700
rect 66940 60690 67060 60700
rect 67190 60690 67310 60700
rect 67440 60690 67560 60700
rect 67690 60690 67810 60700
rect 67940 60690 68060 60700
rect 68190 60690 68310 60700
rect 68440 60690 68560 60700
rect 68690 60690 68810 60700
rect 68940 60690 69060 60700
rect 69190 60690 69310 60700
rect 69440 60690 69560 60700
rect 69690 60690 69810 60700
rect 69940 60690 70060 60700
rect 70190 60690 70310 60700
rect 70440 60690 70560 60700
rect 70690 60690 70810 60700
rect 70940 60690 71000 60700
rect 59000 60560 59050 60690
rect 59200 60560 59300 60690
rect 59450 60560 59550 60690
rect 59700 60560 59800 60690
rect 59950 60560 60050 60690
rect 60200 60560 60300 60690
rect 60450 60560 60550 60690
rect 60700 60560 60800 60690
rect 60950 60560 61050 60690
rect 61200 60560 61300 60690
rect 61450 60560 61550 60690
rect 61700 60560 61800 60690
rect 61950 60560 62050 60690
rect 62200 60560 62300 60690
rect 62450 60560 62550 60690
rect 62700 60560 62800 60690
rect 62950 60560 63050 60690
rect 63200 60560 63300 60690
rect 63450 60560 63550 60690
rect 63700 60560 63800 60690
rect 63950 60560 64050 60690
rect 64200 60560 64300 60690
rect 64450 60560 64550 60690
rect 64700 60560 64800 60690
rect 64950 60560 65050 60690
rect 65200 60560 65300 60690
rect 65450 60560 65550 60690
rect 65700 60560 65800 60690
rect 65950 60560 66050 60690
rect 66200 60560 66300 60690
rect 66450 60560 66550 60690
rect 66700 60560 66800 60690
rect 66950 60560 67050 60690
rect 67200 60560 67300 60690
rect 67450 60560 67550 60690
rect 67700 60560 67800 60690
rect 67950 60560 68050 60690
rect 68200 60560 68300 60690
rect 68450 60560 68550 60690
rect 68700 60560 68800 60690
rect 68950 60560 69050 60690
rect 69200 60560 69300 60690
rect 69450 60560 69550 60690
rect 69700 60560 69800 60690
rect 69950 60560 70050 60690
rect 70200 60560 70300 60690
rect 70450 60560 70550 60690
rect 70700 60560 70800 60690
rect 70950 60560 71000 60690
rect 59000 60550 59060 60560
rect 59190 60550 59310 60560
rect 59440 60550 59560 60560
rect 59690 60550 59810 60560
rect 59940 60550 60060 60560
rect 60190 60550 60310 60560
rect 60440 60550 60560 60560
rect 60690 60550 60810 60560
rect 60940 60550 61060 60560
rect 61190 60550 61310 60560
rect 61440 60550 61560 60560
rect 61690 60550 61810 60560
rect 61940 60550 62060 60560
rect 62190 60550 62310 60560
rect 62440 60550 62560 60560
rect 62690 60550 62810 60560
rect 62940 60550 63060 60560
rect 63190 60550 63310 60560
rect 63440 60550 63560 60560
rect 63690 60550 63810 60560
rect 63940 60550 64060 60560
rect 64190 60550 64310 60560
rect 64440 60550 64560 60560
rect 64690 60550 64810 60560
rect 64940 60550 65060 60560
rect 65190 60550 65310 60560
rect 65440 60550 65560 60560
rect 65690 60550 65810 60560
rect 65940 60550 66060 60560
rect 66190 60550 66310 60560
rect 66440 60550 66560 60560
rect 66690 60550 66810 60560
rect 66940 60550 67060 60560
rect 67190 60550 67310 60560
rect 67440 60550 67560 60560
rect 67690 60550 67810 60560
rect 67940 60550 68060 60560
rect 68190 60550 68310 60560
rect 68440 60550 68560 60560
rect 68690 60550 68810 60560
rect 68940 60550 69060 60560
rect 69190 60550 69310 60560
rect 69440 60550 69560 60560
rect 69690 60550 69810 60560
rect 69940 60550 70060 60560
rect 70190 60550 70310 60560
rect 70440 60550 70560 60560
rect 70690 60550 70810 60560
rect 70940 60550 71000 60560
rect 59000 60450 71000 60550
rect 59000 60440 59060 60450
rect 59190 60440 59310 60450
rect 59440 60440 59560 60450
rect 59690 60440 59810 60450
rect 59940 60440 60060 60450
rect 60190 60440 60310 60450
rect 60440 60440 60560 60450
rect 60690 60440 60810 60450
rect 60940 60440 61060 60450
rect 61190 60440 61310 60450
rect 61440 60440 61560 60450
rect 61690 60440 61810 60450
rect 61940 60440 62060 60450
rect 62190 60440 62310 60450
rect 62440 60440 62560 60450
rect 62690 60440 62810 60450
rect 62940 60440 63060 60450
rect 63190 60440 63310 60450
rect 63440 60440 63560 60450
rect 63690 60440 63810 60450
rect 63940 60440 64060 60450
rect 64190 60440 64310 60450
rect 64440 60440 64560 60450
rect 64690 60440 64810 60450
rect 64940 60440 65060 60450
rect 65190 60440 65310 60450
rect 65440 60440 65560 60450
rect 65690 60440 65810 60450
rect 65940 60440 66060 60450
rect 66190 60440 66310 60450
rect 66440 60440 66560 60450
rect 66690 60440 66810 60450
rect 66940 60440 67060 60450
rect 67190 60440 67310 60450
rect 67440 60440 67560 60450
rect 67690 60440 67810 60450
rect 67940 60440 68060 60450
rect 68190 60440 68310 60450
rect 68440 60440 68560 60450
rect 68690 60440 68810 60450
rect 68940 60440 69060 60450
rect 69190 60440 69310 60450
rect 69440 60440 69560 60450
rect 69690 60440 69810 60450
rect 69940 60440 70060 60450
rect 70190 60440 70310 60450
rect 70440 60440 70560 60450
rect 70690 60440 70810 60450
rect 70940 60440 71000 60450
rect 59000 60310 59050 60440
rect 59200 60310 59300 60440
rect 59450 60310 59550 60440
rect 59700 60310 59800 60440
rect 59950 60310 60050 60440
rect 60200 60310 60300 60440
rect 60450 60310 60550 60440
rect 60700 60310 60800 60440
rect 60950 60310 61050 60440
rect 61200 60310 61300 60440
rect 61450 60310 61550 60440
rect 61700 60310 61800 60440
rect 61950 60310 62050 60440
rect 62200 60310 62300 60440
rect 62450 60310 62550 60440
rect 62700 60310 62800 60440
rect 62950 60310 63050 60440
rect 63200 60310 63300 60440
rect 63450 60310 63550 60440
rect 63700 60310 63800 60440
rect 63950 60310 64050 60440
rect 64200 60310 64300 60440
rect 64450 60310 64550 60440
rect 64700 60310 64800 60440
rect 64950 60310 65050 60440
rect 65200 60310 65300 60440
rect 65450 60310 65550 60440
rect 65700 60310 65800 60440
rect 65950 60310 66050 60440
rect 66200 60310 66300 60440
rect 66450 60310 66550 60440
rect 66700 60310 66800 60440
rect 66950 60310 67050 60440
rect 67200 60310 67300 60440
rect 67450 60310 67550 60440
rect 67700 60310 67800 60440
rect 67950 60310 68050 60440
rect 68200 60310 68300 60440
rect 68450 60310 68550 60440
rect 68700 60310 68800 60440
rect 68950 60310 69050 60440
rect 69200 60310 69300 60440
rect 69450 60310 69550 60440
rect 69700 60310 69800 60440
rect 69950 60310 70050 60440
rect 70200 60310 70300 60440
rect 70450 60310 70550 60440
rect 70700 60310 70800 60440
rect 70950 60310 71000 60440
rect 59000 60300 59060 60310
rect 59190 60300 59310 60310
rect 59440 60300 59560 60310
rect 59690 60300 59810 60310
rect 59940 60300 60060 60310
rect 60190 60300 60310 60310
rect 60440 60300 60560 60310
rect 60690 60300 60810 60310
rect 60940 60300 61060 60310
rect 61190 60300 61310 60310
rect 61440 60300 61560 60310
rect 61690 60300 61810 60310
rect 61940 60300 62060 60310
rect 62190 60300 62310 60310
rect 62440 60300 62560 60310
rect 62690 60300 62810 60310
rect 62940 60300 63060 60310
rect 63190 60300 63310 60310
rect 63440 60300 63560 60310
rect 63690 60300 63810 60310
rect 63940 60300 64060 60310
rect 64190 60300 64310 60310
rect 64440 60300 64560 60310
rect 64690 60300 64810 60310
rect 64940 60300 65060 60310
rect 65190 60300 65310 60310
rect 65440 60300 65560 60310
rect 65690 60300 65810 60310
rect 65940 60300 66060 60310
rect 66190 60300 66310 60310
rect 66440 60300 66560 60310
rect 66690 60300 66810 60310
rect 66940 60300 67060 60310
rect 67190 60300 67310 60310
rect 67440 60300 67560 60310
rect 67690 60300 67810 60310
rect 67940 60300 68060 60310
rect 68190 60300 68310 60310
rect 68440 60300 68560 60310
rect 68690 60300 68810 60310
rect 68940 60300 69060 60310
rect 69190 60300 69310 60310
rect 69440 60300 69560 60310
rect 69690 60300 69810 60310
rect 69940 60300 70060 60310
rect 70190 60300 70310 60310
rect 70440 60300 70560 60310
rect 70690 60300 70810 60310
rect 70940 60300 71000 60310
rect 59000 60200 71000 60300
rect 59000 60190 59060 60200
rect 59190 60190 59310 60200
rect 59440 60190 59560 60200
rect 59690 60190 59810 60200
rect 59940 60190 60060 60200
rect 60190 60190 60310 60200
rect 60440 60190 60560 60200
rect 60690 60190 60810 60200
rect 60940 60190 61060 60200
rect 61190 60190 61310 60200
rect 61440 60190 61560 60200
rect 61690 60190 61810 60200
rect 61940 60190 62060 60200
rect 62190 60190 62310 60200
rect 62440 60190 62560 60200
rect 62690 60190 62810 60200
rect 62940 60190 63060 60200
rect 63190 60190 63310 60200
rect 63440 60190 63560 60200
rect 63690 60190 63810 60200
rect 63940 60190 64060 60200
rect 64190 60190 64310 60200
rect 64440 60190 64560 60200
rect 64690 60190 64810 60200
rect 64940 60190 65060 60200
rect 65190 60190 65310 60200
rect 65440 60190 65560 60200
rect 65690 60190 65810 60200
rect 65940 60190 66060 60200
rect 66190 60190 66310 60200
rect 66440 60190 66560 60200
rect 66690 60190 66810 60200
rect 66940 60190 67060 60200
rect 67190 60190 67310 60200
rect 67440 60190 67560 60200
rect 67690 60190 67810 60200
rect 67940 60190 68060 60200
rect 68190 60190 68310 60200
rect 68440 60190 68560 60200
rect 68690 60190 68810 60200
rect 68940 60190 69060 60200
rect 69190 60190 69310 60200
rect 69440 60190 69560 60200
rect 69690 60190 69810 60200
rect 69940 60190 70060 60200
rect 70190 60190 70310 60200
rect 70440 60190 70560 60200
rect 70690 60190 70810 60200
rect 70940 60190 71000 60200
rect 59000 60060 59050 60190
rect 59200 60060 59300 60190
rect 59450 60060 59550 60190
rect 59700 60060 59800 60190
rect 59950 60060 60050 60190
rect 60200 60060 60300 60190
rect 60450 60060 60550 60190
rect 60700 60060 60800 60190
rect 60950 60060 61050 60190
rect 61200 60060 61300 60190
rect 61450 60060 61550 60190
rect 61700 60060 61800 60190
rect 61950 60060 62050 60190
rect 62200 60060 62300 60190
rect 62450 60060 62550 60190
rect 62700 60060 62800 60190
rect 62950 60060 63050 60190
rect 63200 60060 63300 60190
rect 63450 60060 63550 60190
rect 63700 60060 63800 60190
rect 63950 60060 64050 60190
rect 64200 60060 64300 60190
rect 64450 60060 64550 60190
rect 64700 60060 64800 60190
rect 64950 60060 65050 60190
rect 65200 60060 65300 60190
rect 65450 60060 65550 60190
rect 65700 60060 65800 60190
rect 65950 60060 66050 60190
rect 66200 60060 66300 60190
rect 66450 60060 66550 60190
rect 66700 60060 66800 60190
rect 66950 60060 67050 60190
rect 67200 60060 67300 60190
rect 67450 60060 67550 60190
rect 67700 60060 67800 60190
rect 67950 60060 68050 60190
rect 68200 60060 68300 60190
rect 68450 60060 68550 60190
rect 68700 60060 68800 60190
rect 68950 60060 69050 60190
rect 69200 60060 69300 60190
rect 69450 60060 69550 60190
rect 69700 60060 69800 60190
rect 69950 60060 70050 60190
rect 70200 60060 70300 60190
rect 70450 60060 70550 60190
rect 70700 60060 70800 60190
rect 70950 60060 71000 60190
rect 59000 60050 59060 60060
rect 59190 60050 59310 60060
rect 59440 60050 59560 60060
rect 59690 60050 59810 60060
rect 59940 60050 60060 60060
rect 60190 60050 60310 60060
rect 60440 60050 60560 60060
rect 60690 60050 60810 60060
rect 60940 60050 61060 60060
rect 61190 60050 61310 60060
rect 61440 60050 61560 60060
rect 61690 60050 61810 60060
rect 61940 60050 62060 60060
rect 62190 60050 62310 60060
rect 62440 60050 62560 60060
rect 62690 60050 62810 60060
rect 62940 60050 63060 60060
rect 63190 60050 63310 60060
rect 63440 60050 63560 60060
rect 63690 60050 63810 60060
rect 63940 60050 64060 60060
rect 64190 60050 64310 60060
rect 64440 60050 64560 60060
rect 64690 60050 64810 60060
rect 64940 60050 65060 60060
rect 65190 60050 65310 60060
rect 65440 60050 65560 60060
rect 65690 60050 65810 60060
rect 65940 60050 66060 60060
rect 66190 60050 66310 60060
rect 66440 60050 66560 60060
rect 66690 60050 66810 60060
rect 66940 60050 67060 60060
rect 67190 60050 67310 60060
rect 67440 60050 67560 60060
rect 67690 60050 67810 60060
rect 67940 60050 68060 60060
rect 68190 60050 68310 60060
rect 68440 60050 68560 60060
rect 68690 60050 68810 60060
rect 68940 60050 69060 60060
rect 69190 60050 69310 60060
rect 69440 60050 69560 60060
rect 69690 60050 69810 60060
rect 69940 60050 70060 60060
rect 70190 60050 70310 60060
rect 70440 60050 70560 60060
rect 70690 60050 70810 60060
rect 70940 60050 71000 60060
rect 59000 59950 71000 60050
rect 59000 59940 59060 59950
rect 59190 59940 59310 59950
rect 59440 59940 59560 59950
rect 59690 59940 59810 59950
rect 59940 59940 60060 59950
rect 60190 59940 60310 59950
rect 60440 59940 60560 59950
rect 60690 59940 60810 59950
rect 60940 59940 61060 59950
rect 61190 59940 61310 59950
rect 61440 59940 61560 59950
rect 61690 59940 61810 59950
rect 61940 59940 62060 59950
rect 62190 59940 62310 59950
rect 62440 59940 62560 59950
rect 62690 59940 62810 59950
rect 62940 59940 63060 59950
rect 63190 59940 63310 59950
rect 63440 59940 63560 59950
rect 63690 59940 63810 59950
rect 63940 59940 64060 59950
rect 64190 59940 64310 59950
rect 64440 59940 64560 59950
rect 64690 59940 64810 59950
rect 64940 59940 65060 59950
rect 65190 59940 65310 59950
rect 65440 59940 65560 59950
rect 65690 59940 65810 59950
rect 65940 59940 66060 59950
rect 66190 59940 66310 59950
rect 66440 59940 66560 59950
rect 66690 59940 66810 59950
rect 66940 59940 67060 59950
rect 67190 59940 67310 59950
rect 67440 59940 67560 59950
rect 67690 59940 67810 59950
rect 67940 59940 68060 59950
rect 68190 59940 68310 59950
rect 68440 59940 68560 59950
rect 68690 59940 68810 59950
rect 68940 59940 69060 59950
rect 69190 59940 69310 59950
rect 69440 59940 69560 59950
rect 69690 59940 69810 59950
rect 69940 59940 70060 59950
rect 70190 59940 70310 59950
rect 70440 59940 70560 59950
rect 70690 59940 70810 59950
rect 70940 59940 71000 59950
rect 59000 59810 59050 59940
rect 59200 59810 59300 59940
rect 59450 59810 59550 59940
rect 59700 59810 59800 59940
rect 59950 59810 60050 59940
rect 60200 59810 60300 59940
rect 60450 59810 60550 59940
rect 60700 59810 60800 59940
rect 60950 59810 61050 59940
rect 61200 59810 61300 59940
rect 61450 59810 61550 59940
rect 61700 59810 61800 59940
rect 61950 59810 62050 59940
rect 62200 59810 62300 59940
rect 62450 59810 62550 59940
rect 62700 59810 62800 59940
rect 62950 59810 63050 59940
rect 63200 59810 63300 59940
rect 63450 59810 63550 59940
rect 63700 59810 63800 59940
rect 63950 59810 64050 59940
rect 64200 59810 64300 59940
rect 64450 59810 64550 59940
rect 64700 59810 64800 59940
rect 64950 59810 65050 59940
rect 65200 59810 65300 59940
rect 65450 59810 65550 59940
rect 65700 59810 65800 59940
rect 65950 59810 66050 59940
rect 66200 59810 66300 59940
rect 66450 59810 66550 59940
rect 66700 59810 66800 59940
rect 66950 59810 67050 59940
rect 67200 59810 67300 59940
rect 67450 59810 67550 59940
rect 67700 59810 67800 59940
rect 67950 59810 68050 59940
rect 68200 59810 68300 59940
rect 68450 59810 68550 59940
rect 68700 59810 68800 59940
rect 68950 59810 69050 59940
rect 69200 59810 69300 59940
rect 69450 59810 69550 59940
rect 69700 59810 69800 59940
rect 69950 59810 70050 59940
rect 70200 59810 70300 59940
rect 70450 59810 70550 59940
rect 70700 59810 70800 59940
rect 70950 59810 71000 59940
rect 59000 59800 59060 59810
rect 59190 59800 59310 59810
rect 59440 59800 59560 59810
rect 59690 59800 59810 59810
rect 59940 59800 60060 59810
rect 60190 59800 60310 59810
rect 60440 59800 60560 59810
rect 60690 59800 60810 59810
rect 60940 59800 61060 59810
rect 61190 59800 61310 59810
rect 61440 59800 61560 59810
rect 61690 59800 61810 59810
rect 61940 59800 62060 59810
rect 62190 59800 62310 59810
rect 62440 59800 62560 59810
rect 62690 59800 62810 59810
rect 62940 59800 63060 59810
rect 63190 59800 63310 59810
rect 63440 59800 63560 59810
rect 63690 59800 63810 59810
rect 63940 59800 64060 59810
rect 64190 59800 64310 59810
rect 64440 59800 64560 59810
rect 64690 59800 64810 59810
rect 64940 59800 65060 59810
rect 65190 59800 65310 59810
rect 65440 59800 65560 59810
rect 65690 59800 65810 59810
rect 65940 59800 66060 59810
rect 66190 59800 66310 59810
rect 66440 59800 66560 59810
rect 66690 59800 66810 59810
rect 66940 59800 67060 59810
rect 67190 59800 67310 59810
rect 67440 59800 67560 59810
rect 67690 59800 67810 59810
rect 67940 59800 68060 59810
rect 68190 59800 68310 59810
rect 68440 59800 68560 59810
rect 68690 59800 68810 59810
rect 68940 59800 69060 59810
rect 69190 59800 69310 59810
rect 69440 59800 69560 59810
rect 69690 59800 69810 59810
rect 69940 59800 70060 59810
rect 70190 59800 70310 59810
rect 70440 59800 70560 59810
rect 70690 59800 70810 59810
rect 70940 59800 71000 59810
rect 59000 59700 71000 59800
rect 59000 59690 59060 59700
rect 59190 59690 59310 59700
rect 59440 59690 59560 59700
rect 59690 59690 59810 59700
rect 59940 59690 60060 59700
rect 60190 59690 60310 59700
rect 60440 59690 60560 59700
rect 60690 59690 60810 59700
rect 60940 59690 61060 59700
rect 61190 59690 61310 59700
rect 61440 59690 61560 59700
rect 61690 59690 61810 59700
rect 61940 59690 62060 59700
rect 62190 59690 62310 59700
rect 62440 59690 62560 59700
rect 62690 59690 62810 59700
rect 62940 59690 63060 59700
rect 63190 59690 63310 59700
rect 63440 59690 63560 59700
rect 63690 59690 63810 59700
rect 63940 59690 64060 59700
rect 64190 59690 64310 59700
rect 64440 59690 64560 59700
rect 64690 59690 64810 59700
rect 64940 59690 65060 59700
rect 65190 59690 65310 59700
rect 65440 59690 65560 59700
rect 65690 59690 65810 59700
rect 65940 59690 66060 59700
rect 66190 59690 66310 59700
rect 66440 59690 66560 59700
rect 66690 59690 66810 59700
rect 66940 59690 67060 59700
rect 67190 59690 67310 59700
rect 67440 59690 67560 59700
rect 67690 59690 67810 59700
rect 67940 59690 68060 59700
rect 68190 59690 68310 59700
rect 68440 59690 68560 59700
rect 68690 59690 68810 59700
rect 68940 59690 69060 59700
rect 69190 59690 69310 59700
rect 69440 59690 69560 59700
rect 69690 59690 69810 59700
rect 69940 59690 70060 59700
rect 70190 59690 70310 59700
rect 70440 59690 70560 59700
rect 70690 59690 70810 59700
rect 70940 59690 71000 59700
rect 59000 59560 59050 59690
rect 59200 59560 59300 59690
rect 59450 59560 59550 59690
rect 59700 59560 59800 59690
rect 59950 59560 60050 59690
rect 60200 59560 60300 59690
rect 60450 59560 60550 59690
rect 60700 59560 60800 59690
rect 60950 59560 61050 59690
rect 61200 59560 61300 59690
rect 61450 59560 61550 59690
rect 61700 59560 61800 59690
rect 61950 59560 62050 59690
rect 62200 59560 62300 59690
rect 62450 59560 62550 59690
rect 62700 59560 62800 59690
rect 62950 59560 63050 59690
rect 63200 59560 63300 59690
rect 63450 59560 63550 59690
rect 63700 59560 63800 59690
rect 63950 59560 64050 59690
rect 64200 59560 64300 59690
rect 64450 59560 64550 59690
rect 64700 59560 64800 59690
rect 64950 59560 65050 59690
rect 65200 59560 65300 59690
rect 65450 59560 65550 59690
rect 65700 59560 65800 59690
rect 65950 59560 66050 59690
rect 66200 59560 66300 59690
rect 66450 59560 66550 59690
rect 66700 59560 66800 59690
rect 66950 59560 67050 59690
rect 67200 59560 67300 59690
rect 67450 59560 67550 59690
rect 67700 59560 67800 59690
rect 67950 59560 68050 59690
rect 68200 59560 68300 59690
rect 68450 59560 68550 59690
rect 68700 59560 68800 59690
rect 68950 59560 69050 59690
rect 69200 59560 69300 59690
rect 69450 59560 69550 59690
rect 69700 59560 69800 59690
rect 69950 59560 70050 59690
rect 70200 59560 70300 59690
rect 70450 59560 70550 59690
rect 70700 59560 70800 59690
rect 70950 59560 71000 59690
rect 59000 59550 59060 59560
rect 59190 59550 59310 59560
rect 59440 59550 59560 59560
rect 59690 59550 59810 59560
rect 59940 59550 60060 59560
rect 60190 59550 60310 59560
rect 60440 59550 60560 59560
rect 60690 59550 60810 59560
rect 60940 59550 61060 59560
rect 61190 59550 61310 59560
rect 61440 59550 61560 59560
rect 61690 59550 61810 59560
rect 61940 59550 62060 59560
rect 62190 59550 62310 59560
rect 62440 59550 62560 59560
rect 62690 59550 62810 59560
rect 62940 59550 63060 59560
rect 63190 59550 63310 59560
rect 63440 59550 63560 59560
rect 63690 59550 63810 59560
rect 63940 59550 64060 59560
rect 64190 59550 64310 59560
rect 64440 59550 64560 59560
rect 64690 59550 64810 59560
rect 64940 59550 65060 59560
rect 65190 59550 65310 59560
rect 65440 59550 65560 59560
rect 65690 59550 65810 59560
rect 65940 59550 66060 59560
rect 66190 59550 66310 59560
rect 66440 59550 66560 59560
rect 66690 59550 66810 59560
rect 66940 59550 67060 59560
rect 67190 59550 67310 59560
rect 67440 59550 67560 59560
rect 67690 59550 67810 59560
rect 67940 59550 68060 59560
rect 68190 59550 68310 59560
rect 68440 59550 68560 59560
rect 68690 59550 68810 59560
rect 68940 59550 69060 59560
rect 69190 59550 69310 59560
rect 69440 59550 69560 59560
rect 69690 59550 69810 59560
rect 69940 59550 70060 59560
rect 70190 59550 70310 59560
rect 70440 59550 70560 59560
rect 70690 59550 70810 59560
rect 70940 59550 71000 59560
rect 59000 59450 71000 59550
rect 59000 59440 59060 59450
rect 59190 59440 59310 59450
rect 59440 59440 59560 59450
rect 59690 59440 59810 59450
rect 59940 59440 60060 59450
rect 60190 59440 60310 59450
rect 60440 59440 60560 59450
rect 60690 59440 60810 59450
rect 60940 59440 61060 59450
rect 61190 59440 61310 59450
rect 61440 59440 61560 59450
rect 61690 59440 61810 59450
rect 61940 59440 62060 59450
rect 62190 59440 62310 59450
rect 62440 59440 62560 59450
rect 62690 59440 62810 59450
rect 62940 59440 63060 59450
rect 63190 59440 63310 59450
rect 63440 59440 63560 59450
rect 63690 59440 63810 59450
rect 63940 59440 64060 59450
rect 64190 59440 64310 59450
rect 64440 59440 64560 59450
rect 64690 59440 64810 59450
rect 64940 59440 65060 59450
rect 65190 59440 65310 59450
rect 65440 59440 65560 59450
rect 65690 59440 65810 59450
rect 65940 59440 66060 59450
rect 66190 59440 66310 59450
rect 66440 59440 66560 59450
rect 66690 59440 66810 59450
rect 66940 59440 67060 59450
rect 67190 59440 67310 59450
rect 67440 59440 67560 59450
rect 67690 59440 67810 59450
rect 67940 59440 68060 59450
rect 68190 59440 68310 59450
rect 68440 59440 68560 59450
rect 68690 59440 68810 59450
rect 68940 59440 69060 59450
rect 69190 59440 69310 59450
rect 69440 59440 69560 59450
rect 69690 59440 69810 59450
rect 69940 59440 70060 59450
rect 70190 59440 70310 59450
rect 70440 59440 70560 59450
rect 70690 59440 70810 59450
rect 70940 59440 71000 59450
rect 59000 59310 59050 59440
rect 59200 59310 59300 59440
rect 59450 59310 59550 59440
rect 59700 59310 59800 59440
rect 59950 59310 60050 59440
rect 60200 59310 60300 59440
rect 60450 59310 60550 59440
rect 60700 59310 60800 59440
rect 60950 59310 61050 59440
rect 61200 59310 61300 59440
rect 61450 59310 61550 59440
rect 61700 59310 61800 59440
rect 61950 59310 62050 59440
rect 62200 59310 62300 59440
rect 62450 59310 62550 59440
rect 62700 59310 62800 59440
rect 62950 59310 63050 59440
rect 63200 59310 63300 59440
rect 63450 59310 63550 59440
rect 63700 59310 63800 59440
rect 63950 59310 64050 59440
rect 64200 59310 64300 59440
rect 64450 59310 64550 59440
rect 64700 59310 64800 59440
rect 64950 59310 65050 59440
rect 65200 59310 65300 59440
rect 65450 59310 65550 59440
rect 65700 59310 65800 59440
rect 65950 59310 66050 59440
rect 66200 59310 66300 59440
rect 66450 59310 66550 59440
rect 66700 59310 66800 59440
rect 66950 59310 67050 59440
rect 67200 59310 67300 59440
rect 67450 59310 67550 59440
rect 67700 59310 67800 59440
rect 67950 59310 68050 59440
rect 68200 59310 68300 59440
rect 68450 59310 68550 59440
rect 68700 59310 68800 59440
rect 68950 59310 69050 59440
rect 69200 59310 69300 59440
rect 69450 59310 69550 59440
rect 69700 59310 69800 59440
rect 69950 59310 70050 59440
rect 70200 59310 70300 59440
rect 70450 59310 70550 59440
rect 70700 59310 70800 59440
rect 70950 59310 71000 59440
rect 59000 59300 59060 59310
rect 59190 59300 59310 59310
rect 59440 59300 59560 59310
rect 59690 59300 59810 59310
rect 59940 59300 60060 59310
rect 60190 59300 60310 59310
rect 60440 59300 60560 59310
rect 60690 59300 60810 59310
rect 60940 59300 61060 59310
rect 61190 59300 61310 59310
rect 61440 59300 61560 59310
rect 61690 59300 61810 59310
rect 61940 59300 62060 59310
rect 62190 59300 62310 59310
rect 62440 59300 62560 59310
rect 62690 59300 62810 59310
rect 62940 59300 63060 59310
rect 63190 59300 63310 59310
rect 63440 59300 63560 59310
rect 63690 59300 63810 59310
rect 63940 59300 64060 59310
rect 64190 59300 64310 59310
rect 64440 59300 64560 59310
rect 64690 59300 64810 59310
rect 64940 59300 65060 59310
rect 65190 59300 65310 59310
rect 65440 59300 65560 59310
rect 65690 59300 65810 59310
rect 65940 59300 66060 59310
rect 66190 59300 66310 59310
rect 66440 59300 66560 59310
rect 66690 59300 66810 59310
rect 66940 59300 67060 59310
rect 67190 59300 67310 59310
rect 67440 59300 67560 59310
rect 67690 59300 67810 59310
rect 67940 59300 68060 59310
rect 68190 59300 68310 59310
rect 68440 59300 68560 59310
rect 68690 59300 68810 59310
rect 68940 59300 69060 59310
rect 69190 59300 69310 59310
rect 69440 59300 69560 59310
rect 69690 59300 69810 59310
rect 69940 59300 70060 59310
rect 70190 59300 70310 59310
rect 70440 59300 70560 59310
rect 70690 59300 70810 59310
rect 70940 59300 71000 59310
rect 59000 59200 71000 59300
rect 59000 59190 59060 59200
rect 59190 59190 59310 59200
rect 59440 59190 59560 59200
rect 59690 59190 59810 59200
rect 59940 59190 60060 59200
rect 60190 59190 60310 59200
rect 60440 59190 60560 59200
rect 60690 59190 60810 59200
rect 60940 59190 61060 59200
rect 61190 59190 61310 59200
rect 61440 59190 61560 59200
rect 61690 59190 61810 59200
rect 61940 59190 62060 59200
rect 62190 59190 62310 59200
rect 62440 59190 62560 59200
rect 62690 59190 62810 59200
rect 62940 59190 63060 59200
rect 63190 59190 63310 59200
rect 63440 59190 63560 59200
rect 63690 59190 63810 59200
rect 63940 59190 64060 59200
rect 64190 59190 64310 59200
rect 64440 59190 64560 59200
rect 64690 59190 64810 59200
rect 64940 59190 65060 59200
rect 65190 59190 65310 59200
rect 65440 59190 65560 59200
rect 65690 59190 65810 59200
rect 65940 59190 66060 59200
rect 66190 59190 66310 59200
rect 66440 59190 66560 59200
rect 66690 59190 66810 59200
rect 66940 59190 67060 59200
rect 67190 59190 67310 59200
rect 67440 59190 67560 59200
rect 67690 59190 67810 59200
rect 67940 59190 68060 59200
rect 68190 59190 68310 59200
rect 68440 59190 68560 59200
rect 68690 59190 68810 59200
rect 68940 59190 69060 59200
rect 69190 59190 69310 59200
rect 69440 59190 69560 59200
rect 69690 59190 69810 59200
rect 69940 59190 70060 59200
rect 70190 59190 70310 59200
rect 70440 59190 70560 59200
rect 70690 59190 70810 59200
rect 70940 59190 71000 59200
rect 59000 59060 59050 59190
rect 59200 59060 59300 59190
rect 59450 59060 59550 59190
rect 59700 59060 59800 59190
rect 59950 59060 60050 59190
rect 60200 59060 60300 59190
rect 60450 59060 60550 59190
rect 60700 59060 60800 59190
rect 60950 59060 61050 59190
rect 61200 59060 61300 59190
rect 61450 59060 61550 59190
rect 61700 59060 61800 59190
rect 61950 59060 62050 59190
rect 62200 59060 62300 59190
rect 62450 59060 62550 59190
rect 62700 59060 62800 59190
rect 62950 59060 63050 59190
rect 63200 59060 63300 59190
rect 63450 59060 63550 59190
rect 63700 59060 63800 59190
rect 63950 59060 64050 59190
rect 64200 59060 64300 59190
rect 64450 59060 64550 59190
rect 64700 59060 64800 59190
rect 64950 59060 65050 59190
rect 65200 59060 65300 59190
rect 65450 59060 65550 59190
rect 65700 59060 65800 59190
rect 65950 59060 66050 59190
rect 66200 59060 66300 59190
rect 66450 59060 66550 59190
rect 66700 59060 66800 59190
rect 66950 59060 67050 59190
rect 67200 59060 67300 59190
rect 67450 59060 67550 59190
rect 67700 59060 67800 59190
rect 67950 59060 68050 59190
rect 68200 59060 68300 59190
rect 68450 59060 68550 59190
rect 68700 59060 68800 59190
rect 68950 59060 69050 59190
rect 69200 59060 69300 59190
rect 69450 59060 69550 59190
rect 69700 59060 69800 59190
rect 69950 59060 70050 59190
rect 70200 59060 70300 59190
rect 70450 59060 70550 59190
rect 70700 59060 70800 59190
rect 70950 59060 71000 59190
rect 59000 59050 59060 59060
rect 59190 59050 59310 59060
rect 59440 59050 59560 59060
rect 59690 59050 59810 59060
rect 59940 59050 60060 59060
rect 60190 59050 60310 59060
rect 60440 59050 60560 59060
rect 60690 59050 60810 59060
rect 60940 59050 61060 59060
rect 61190 59050 61310 59060
rect 61440 59050 61560 59060
rect 61690 59050 61810 59060
rect 61940 59050 62060 59060
rect 62190 59050 62310 59060
rect 62440 59050 62560 59060
rect 62690 59050 62810 59060
rect 62940 59050 63060 59060
rect 63190 59050 63310 59060
rect 63440 59050 63560 59060
rect 63690 59050 63810 59060
rect 63940 59050 64060 59060
rect 64190 59050 64310 59060
rect 64440 59050 64560 59060
rect 64690 59050 64810 59060
rect 64940 59050 65060 59060
rect 65190 59050 65310 59060
rect 65440 59050 65560 59060
rect 65690 59050 65810 59060
rect 65940 59050 66060 59060
rect 66190 59050 66310 59060
rect 66440 59050 66560 59060
rect 66690 59050 66810 59060
rect 66940 59050 67060 59060
rect 67190 59050 67310 59060
rect 67440 59050 67560 59060
rect 67690 59050 67810 59060
rect 67940 59050 68060 59060
rect 68190 59050 68310 59060
rect 68440 59050 68560 59060
rect 68690 59050 68810 59060
rect 68940 59050 69060 59060
rect 69190 59050 69310 59060
rect 69440 59050 69560 59060
rect 69690 59050 69810 59060
rect 69940 59050 70060 59060
rect 70190 59050 70310 59060
rect 70440 59050 70560 59060
rect 70690 59050 70810 59060
rect 70940 59050 71000 59060
rect 59000 58950 71000 59050
rect 59000 58940 59060 58950
rect 59190 58940 59310 58950
rect 59440 58940 59560 58950
rect 59690 58940 59810 58950
rect 59940 58940 60060 58950
rect 60190 58940 60310 58950
rect 60440 58940 60560 58950
rect 60690 58940 60810 58950
rect 60940 58940 61060 58950
rect 61190 58940 61310 58950
rect 61440 58940 61560 58950
rect 61690 58940 61810 58950
rect 61940 58940 62060 58950
rect 62190 58940 62310 58950
rect 62440 58940 62560 58950
rect 62690 58940 62810 58950
rect 62940 58940 63060 58950
rect 63190 58940 63310 58950
rect 63440 58940 63560 58950
rect 63690 58940 63810 58950
rect 63940 58940 64060 58950
rect 64190 58940 64310 58950
rect 64440 58940 64560 58950
rect 64690 58940 64810 58950
rect 64940 58940 65060 58950
rect 65190 58940 65310 58950
rect 65440 58940 65560 58950
rect 65690 58940 65810 58950
rect 65940 58940 66060 58950
rect 66190 58940 66310 58950
rect 66440 58940 66560 58950
rect 66690 58940 66810 58950
rect 66940 58940 67060 58950
rect 67190 58940 67310 58950
rect 67440 58940 67560 58950
rect 67690 58940 67810 58950
rect 67940 58940 68060 58950
rect 68190 58940 68310 58950
rect 68440 58940 68560 58950
rect 68690 58940 68810 58950
rect 68940 58940 69060 58950
rect 69190 58940 69310 58950
rect 69440 58940 69560 58950
rect 69690 58940 69810 58950
rect 69940 58940 70060 58950
rect 70190 58940 70310 58950
rect 70440 58940 70560 58950
rect 70690 58940 70810 58950
rect 70940 58940 71000 58950
rect 59000 58810 59050 58940
rect 59200 58810 59300 58940
rect 59450 58810 59550 58940
rect 59700 58810 59800 58940
rect 59950 58810 60050 58940
rect 60200 58810 60300 58940
rect 60450 58810 60550 58940
rect 60700 58810 60800 58940
rect 60950 58810 61050 58940
rect 61200 58810 61300 58940
rect 61450 58810 61550 58940
rect 61700 58810 61800 58940
rect 61950 58810 62050 58940
rect 62200 58810 62300 58940
rect 62450 58810 62550 58940
rect 62700 58810 62800 58940
rect 62950 58810 63050 58940
rect 63200 58810 63300 58940
rect 63450 58810 63550 58940
rect 63700 58810 63800 58940
rect 63950 58810 64050 58940
rect 64200 58810 64300 58940
rect 64450 58810 64550 58940
rect 64700 58810 64800 58940
rect 64950 58810 65050 58940
rect 65200 58810 65300 58940
rect 65450 58810 65550 58940
rect 65700 58810 65800 58940
rect 65950 58810 66050 58940
rect 66200 58810 66300 58940
rect 66450 58810 66550 58940
rect 66700 58810 66800 58940
rect 66950 58810 67050 58940
rect 67200 58810 67300 58940
rect 67450 58810 67550 58940
rect 67700 58810 67800 58940
rect 67950 58810 68050 58940
rect 68200 58810 68300 58940
rect 68450 58810 68550 58940
rect 68700 58810 68800 58940
rect 68950 58810 69050 58940
rect 69200 58810 69300 58940
rect 69450 58810 69550 58940
rect 69700 58810 69800 58940
rect 69950 58810 70050 58940
rect 70200 58810 70300 58940
rect 70450 58810 70550 58940
rect 70700 58810 70800 58940
rect 70950 58810 71000 58940
rect 59000 58800 59060 58810
rect 59190 58800 59310 58810
rect 59440 58800 59560 58810
rect 59690 58800 59810 58810
rect 59940 58800 60060 58810
rect 60190 58800 60310 58810
rect 60440 58800 60560 58810
rect 60690 58800 60810 58810
rect 60940 58800 61060 58810
rect 61190 58800 61310 58810
rect 61440 58800 61560 58810
rect 61690 58800 61810 58810
rect 61940 58800 62060 58810
rect 62190 58800 62310 58810
rect 62440 58800 62560 58810
rect 62690 58800 62810 58810
rect 62940 58800 63060 58810
rect 63190 58800 63310 58810
rect 63440 58800 63560 58810
rect 63690 58800 63810 58810
rect 63940 58800 64060 58810
rect 64190 58800 64310 58810
rect 64440 58800 64560 58810
rect 64690 58800 64810 58810
rect 64940 58800 65060 58810
rect 65190 58800 65310 58810
rect 65440 58800 65560 58810
rect 65690 58800 65810 58810
rect 65940 58800 66060 58810
rect 66190 58800 66310 58810
rect 66440 58800 66560 58810
rect 66690 58800 66810 58810
rect 66940 58800 67060 58810
rect 67190 58800 67310 58810
rect 67440 58800 67560 58810
rect 67690 58800 67810 58810
rect 67940 58800 68060 58810
rect 68190 58800 68310 58810
rect 68440 58800 68560 58810
rect 68690 58800 68810 58810
rect 68940 58800 69060 58810
rect 69190 58800 69310 58810
rect 69440 58800 69560 58810
rect 69690 58800 69810 58810
rect 69940 58800 70060 58810
rect 70190 58800 70310 58810
rect 70440 58800 70560 58810
rect 70690 58800 70810 58810
rect 70940 58800 71000 58810
rect 59000 58700 71000 58800
rect 59000 58690 59060 58700
rect 59190 58690 59310 58700
rect 59440 58690 59560 58700
rect 59690 58690 59810 58700
rect 59940 58690 60060 58700
rect 60190 58690 60310 58700
rect 60440 58690 60560 58700
rect 60690 58690 60810 58700
rect 60940 58690 61060 58700
rect 61190 58690 61310 58700
rect 61440 58690 61560 58700
rect 61690 58690 61810 58700
rect 61940 58690 62060 58700
rect 62190 58690 62310 58700
rect 62440 58690 62560 58700
rect 62690 58690 62810 58700
rect 62940 58690 63060 58700
rect 63190 58690 63310 58700
rect 63440 58690 63560 58700
rect 63690 58690 63810 58700
rect 63940 58690 64060 58700
rect 64190 58690 64310 58700
rect 64440 58690 64560 58700
rect 64690 58690 64810 58700
rect 64940 58690 65060 58700
rect 65190 58690 65310 58700
rect 65440 58690 65560 58700
rect 65690 58690 65810 58700
rect 65940 58690 66060 58700
rect 66190 58690 66310 58700
rect 66440 58690 66560 58700
rect 66690 58690 66810 58700
rect 66940 58690 67060 58700
rect 67190 58690 67310 58700
rect 67440 58690 67560 58700
rect 67690 58690 67810 58700
rect 67940 58690 68060 58700
rect 68190 58690 68310 58700
rect 68440 58690 68560 58700
rect 68690 58690 68810 58700
rect 68940 58690 69060 58700
rect 69190 58690 69310 58700
rect 69440 58690 69560 58700
rect 69690 58690 69810 58700
rect 69940 58690 70060 58700
rect 70190 58690 70310 58700
rect 70440 58690 70560 58700
rect 70690 58690 70810 58700
rect 70940 58690 71000 58700
rect 59000 58560 59050 58690
rect 59200 58560 59300 58690
rect 59450 58560 59550 58690
rect 59700 58560 59800 58690
rect 59950 58560 60050 58690
rect 60200 58560 60300 58690
rect 60450 58560 60550 58690
rect 60700 58560 60800 58690
rect 60950 58560 61050 58690
rect 61200 58560 61300 58690
rect 61450 58560 61550 58690
rect 61700 58560 61800 58690
rect 61950 58560 62050 58690
rect 62200 58560 62300 58690
rect 62450 58560 62550 58690
rect 62700 58560 62800 58690
rect 62950 58560 63050 58690
rect 63200 58560 63300 58690
rect 63450 58560 63550 58690
rect 63700 58560 63800 58690
rect 63950 58560 64050 58690
rect 64200 58560 64300 58690
rect 64450 58560 64550 58690
rect 64700 58560 64800 58690
rect 64950 58560 65050 58690
rect 65200 58560 65300 58690
rect 65450 58560 65550 58690
rect 65700 58560 65800 58690
rect 65950 58560 66050 58690
rect 66200 58560 66300 58690
rect 66450 58560 66550 58690
rect 66700 58560 66800 58690
rect 66950 58560 67050 58690
rect 67200 58560 67300 58690
rect 67450 58560 67550 58690
rect 67700 58560 67800 58690
rect 67950 58560 68050 58690
rect 68200 58560 68300 58690
rect 68450 58560 68550 58690
rect 68700 58560 68800 58690
rect 68950 58560 69050 58690
rect 69200 58560 69300 58690
rect 69450 58560 69550 58690
rect 69700 58560 69800 58690
rect 69950 58560 70050 58690
rect 70200 58560 70300 58690
rect 70450 58560 70550 58690
rect 70700 58560 70800 58690
rect 70950 58560 71000 58690
rect 59000 58550 59060 58560
rect 59190 58550 59310 58560
rect 59440 58550 59560 58560
rect 59690 58550 59810 58560
rect 59940 58550 60060 58560
rect 60190 58550 60310 58560
rect 60440 58550 60560 58560
rect 60690 58550 60810 58560
rect 60940 58550 61060 58560
rect 61190 58550 61310 58560
rect 61440 58550 61560 58560
rect 61690 58550 61810 58560
rect 61940 58550 62060 58560
rect 62190 58550 62310 58560
rect 62440 58550 62560 58560
rect 62690 58550 62810 58560
rect 62940 58550 63060 58560
rect 63190 58550 63310 58560
rect 63440 58550 63560 58560
rect 63690 58550 63810 58560
rect 63940 58550 64060 58560
rect 64190 58550 64310 58560
rect 64440 58550 64560 58560
rect 64690 58550 64810 58560
rect 64940 58550 65060 58560
rect 65190 58550 65310 58560
rect 65440 58550 65560 58560
rect 65690 58550 65810 58560
rect 65940 58550 66060 58560
rect 66190 58550 66310 58560
rect 66440 58550 66560 58560
rect 66690 58550 66810 58560
rect 66940 58550 67060 58560
rect 67190 58550 67310 58560
rect 67440 58550 67560 58560
rect 67690 58550 67810 58560
rect 67940 58550 68060 58560
rect 68190 58550 68310 58560
rect 68440 58550 68560 58560
rect 68690 58550 68810 58560
rect 68940 58550 69060 58560
rect 69190 58550 69310 58560
rect 69440 58550 69560 58560
rect 69690 58550 69810 58560
rect 69940 58550 70060 58560
rect 70190 58550 70310 58560
rect 70440 58550 70560 58560
rect 70690 58550 70810 58560
rect 70940 58550 71000 58560
rect 59000 58450 71000 58550
rect 59000 58440 59060 58450
rect 59190 58440 59310 58450
rect 59440 58440 59560 58450
rect 59690 58440 59810 58450
rect 59940 58440 60060 58450
rect 60190 58440 60310 58450
rect 60440 58440 60560 58450
rect 60690 58440 60810 58450
rect 60940 58440 61060 58450
rect 61190 58440 61310 58450
rect 61440 58440 61560 58450
rect 61690 58440 61810 58450
rect 61940 58440 62060 58450
rect 62190 58440 62310 58450
rect 62440 58440 62560 58450
rect 62690 58440 62810 58450
rect 62940 58440 63060 58450
rect 63190 58440 63310 58450
rect 63440 58440 63560 58450
rect 63690 58440 63810 58450
rect 63940 58440 64060 58450
rect 64190 58440 64310 58450
rect 64440 58440 64560 58450
rect 64690 58440 64810 58450
rect 64940 58440 65060 58450
rect 65190 58440 65310 58450
rect 65440 58440 65560 58450
rect 65690 58440 65810 58450
rect 65940 58440 66060 58450
rect 66190 58440 66310 58450
rect 66440 58440 66560 58450
rect 66690 58440 66810 58450
rect 66940 58440 67060 58450
rect 67190 58440 67310 58450
rect 67440 58440 67560 58450
rect 67690 58440 67810 58450
rect 67940 58440 68060 58450
rect 68190 58440 68310 58450
rect 68440 58440 68560 58450
rect 68690 58440 68810 58450
rect 68940 58440 69060 58450
rect 69190 58440 69310 58450
rect 69440 58440 69560 58450
rect 69690 58440 69810 58450
rect 69940 58440 70060 58450
rect 70190 58440 70310 58450
rect 70440 58440 70560 58450
rect 70690 58440 70810 58450
rect 70940 58440 71000 58450
rect 59000 58310 59050 58440
rect 59200 58310 59300 58440
rect 59450 58310 59550 58440
rect 59700 58310 59800 58440
rect 59950 58310 60050 58440
rect 60200 58310 60300 58440
rect 60450 58310 60550 58440
rect 60700 58310 60800 58440
rect 60950 58310 61050 58440
rect 61200 58310 61300 58440
rect 61450 58310 61550 58440
rect 61700 58310 61800 58440
rect 61950 58310 62050 58440
rect 62200 58310 62300 58440
rect 62450 58310 62550 58440
rect 62700 58310 62800 58440
rect 62950 58310 63050 58440
rect 63200 58310 63300 58440
rect 63450 58310 63550 58440
rect 63700 58310 63800 58440
rect 63950 58310 64050 58440
rect 64200 58310 64300 58440
rect 64450 58310 64550 58440
rect 64700 58310 64800 58440
rect 64950 58310 65050 58440
rect 65200 58310 65300 58440
rect 65450 58310 65550 58440
rect 65700 58310 65800 58440
rect 65950 58310 66050 58440
rect 66200 58310 66300 58440
rect 66450 58310 66550 58440
rect 66700 58310 66800 58440
rect 66950 58310 67050 58440
rect 67200 58310 67300 58440
rect 67450 58310 67550 58440
rect 67700 58310 67800 58440
rect 67950 58310 68050 58440
rect 68200 58310 68300 58440
rect 68450 58310 68550 58440
rect 68700 58310 68800 58440
rect 68950 58310 69050 58440
rect 69200 58310 69300 58440
rect 69450 58310 69550 58440
rect 69700 58310 69800 58440
rect 69950 58310 70050 58440
rect 70200 58310 70300 58440
rect 70450 58310 70550 58440
rect 70700 58310 70800 58440
rect 70950 58310 71000 58440
rect 59000 58300 59060 58310
rect 59190 58300 59310 58310
rect 59440 58300 59560 58310
rect 59690 58300 59810 58310
rect 59940 58300 60060 58310
rect 60190 58300 60310 58310
rect 60440 58300 60560 58310
rect 60690 58300 60810 58310
rect 60940 58300 61060 58310
rect 61190 58300 61310 58310
rect 61440 58300 61560 58310
rect 61690 58300 61810 58310
rect 61940 58300 62060 58310
rect 62190 58300 62310 58310
rect 62440 58300 62560 58310
rect 62690 58300 62810 58310
rect 62940 58300 63060 58310
rect 63190 58300 63310 58310
rect 63440 58300 63560 58310
rect 63690 58300 63810 58310
rect 63940 58300 64060 58310
rect 64190 58300 64310 58310
rect 64440 58300 64560 58310
rect 64690 58300 64810 58310
rect 64940 58300 65060 58310
rect 65190 58300 65310 58310
rect 65440 58300 65560 58310
rect 65690 58300 65810 58310
rect 65940 58300 66060 58310
rect 66190 58300 66310 58310
rect 66440 58300 66560 58310
rect 66690 58300 66810 58310
rect 66940 58300 67060 58310
rect 67190 58300 67310 58310
rect 67440 58300 67560 58310
rect 67690 58300 67810 58310
rect 67940 58300 68060 58310
rect 68190 58300 68310 58310
rect 68440 58300 68560 58310
rect 68690 58300 68810 58310
rect 68940 58300 69060 58310
rect 69190 58300 69310 58310
rect 69440 58300 69560 58310
rect 69690 58300 69810 58310
rect 69940 58300 70060 58310
rect 70190 58300 70310 58310
rect 70440 58300 70560 58310
rect 70690 58300 70810 58310
rect 70940 58300 71000 58310
rect 59000 58200 71000 58300
rect 59000 58190 59060 58200
rect 59190 58190 59310 58200
rect 59440 58190 59560 58200
rect 59690 58190 59810 58200
rect 59940 58190 60060 58200
rect 60190 58190 60310 58200
rect 60440 58190 60560 58200
rect 60690 58190 60810 58200
rect 60940 58190 61060 58200
rect 61190 58190 61310 58200
rect 61440 58190 61560 58200
rect 61690 58190 61810 58200
rect 61940 58190 62060 58200
rect 62190 58190 62310 58200
rect 62440 58190 62560 58200
rect 62690 58190 62810 58200
rect 62940 58190 63060 58200
rect 63190 58190 63310 58200
rect 63440 58190 63560 58200
rect 63690 58190 63810 58200
rect 63940 58190 64060 58200
rect 64190 58190 64310 58200
rect 64440 58190 64560 58200
rect 64690 58190 64810 58200
rect 64940 58190 65060 58200
rect 65190 58190 65310 58200
rect 65440 58190 65560 58200
rect 65690 58190 65810 58200
rect 65940 58190 66060 58200
rect 66190 58190 66310 58200
rect 66440 58190 66560 58200
rect 66690 58190 66810 58200
rect 66940 58190 67060 58200
rect 67190 58190 67310 58200
rect 67440 58190 67560 58200
rect 67690 58190 67810 58200
rect 67940 58190 68060 58200
rect 68190 58190 68310 58200
rect 68440 58190 68560 58200
rect 68690 58190 68810 58200
rect 68940 58190 69060 58200
rect 69190 58190 69310 58200
rect 69440 58190 69560 58200
rect 69690 58190 69810 58200
rect 69940 58190 70060 58200
rect 70190 58190 70310 58200
rect 70440 58190 70560 58200
rect 70690 58190 70810 58200
rect 70940 58190 71000 58200
rect 59000 58060 59050 58190
rect 59200 58060 59300 58190
rect 59450 58060 59550 58190
rect 59700 58060 59800 58190
rect 59950 58060 60050 58190
rect 60200 58060 60300 58190
rect 60450 58060 60550 58190
rect 60700 58060 60800 58190
rect 60950 58060 61050 58190
rect 61200 58060 61300 58190
rect 61450 58060 61550 58190
rect 61700 58060 61800 58190
rect 61950 58060 62050 58190
rect 62200 58060 62300 58190
rect 62450 58060 62550 58190
rect 62700 58060 62800 58190
rect 62950 58060 63050 58190
rect 63200 58060 63300 58190
rect 63450 58060 63550 58190
rect 63700 58060 63800 58190
rect 63950 58060 64050 58190
rect 64200 58060 64300 58190
rect 64450 58060 64550 58190
rect 64700 58060 64800 58190
rect 64950 58060 65050 58190
rect 65200 58060 65300 58190
rect 65450 58060 65550 58190
rect 65700 58060 65800 58190
rect 65950 58060 66050 58190
rect 66200 58060 66300 58190
rect 66450 58060 66550 58190
rect 66700 58060 66800 58190
rect 66950 58060 67050 58190
rect 67200 58060 67300 58190
rect 67450 58060 67550 58190
rect 67700 58060 67800 58190
rect 67950 58060 68050 58190
rect 68200 58060 68300 58190
rect 68450 58060 68550 58190
rect 68700 58060 68800 58190
rect 68950 58060 69050 58190
rect 69200 58060 69300 58190
rect 69450 58060 69550 58190
rect 69700 58060 69800 58190
rect 69950 58060 70050 58190
rect 70200 58060 70300 58190
rect 70450 58060 70550 58190
rect 70700 58060 70800 58190
rect 70950 58060 71000 58190
rect 59000 58050 59060 58060
rect 59190 58050 59310 58060
rect 59440 58050 59560 58060
rect 59690 58050 59810 58060
rect 59940 58050 60060 58060
rect 60190 58050 60310 58060
rect 60440 58050 60560 58060
rect 60690 58050 60810 58060
rect 60940 58050 61060 58060
rect 61190 58050 61310 58060
rect 61440 58050 61560 58060
rect 61690 58050 61810 58060
rect 61940 58050 62060 58060
rect 62190 58050 62310 58060
rect 62440 58050 62560 58060
rect 62690 58050 62810 58060
rect 62940 58050 63060 58060
rect 63190 58050 63310 58060
rect 63440 58050 63560 58060
rect 63690 58050 63810 58060
rect 63940 58050 64060 58060
rect 64190 58050 64310 58060
rect 64440 58050 64560 58060
rect 64690 58050 64810 58060
rect 64940 58050 65060 58060
rect 65190 58050 65310 58060
rect 65440 58050 65560 58060
rect 65690 58050 65810 58060
rect 65940 58050 66060 58060
rect 66190 58050 66310 58060
rect 66440 58050 66560 58060
rect 66690 58050 66810 58060
rect 66940 58050 67060 58060
rect 67190 58050 67310 58060
rect 67440 58050 67560 58060
rect 67690 58050 67810 58060
rect 67940 58050 68060 58060
rect 68190 58050 68310 58060
rect 68440 58050 68560 58060
rect 68690 58050 68810 58060
rect 68940 58050 69060 58060
rect 69190 58050 69310 58060
rect 69440 58050 69560 58060
rect 69690 58050 69810 58060
rect 69940 58050 70060 58060
rect 70190 58050 70310 58060
rect 70440 58050 70560 58060
rect 70690 58050 70810 58060
rect 70940 58050 71000 58060
rect 59000 57950 71000 58050
rect 59000 57940 59060 57950
rect 59190 57940 59310 57950
rect 59440 57940 59560 57950
rect 59690 57940 59810 57950
rect 59940 57940 60060 57950
rect 60190 57940 60310 57950
rect 60440 57940 60560 57950
rect 60690 57940 60810 57950
rect 60940 57940 61060 57950
rect 61190 57940 61310 57950
rect 61440 57940 61560 57950
rect 61690 57940 61810 57950
rect 61940 57940 62060 57950
rect 62190 57940 62310 57950
rect 62440 57940 62560 57950
rect 62690 57940 62810 57950
rect 62940 57940 63060 57950
rect 63190 57940 63310 57950
rect 63440 57940 63560 57950
rect 63690 57940 63810 57950
rect 63940 57940 64060 57950
rect 64190 57940 64310 57950
rect 64440 57940 64560 57950
rect 64690 57940 64810 57950
rect 64940 57940 65060 57950
rect 65190 57940 65310 57950
rect 65440 57940 65560 57950
rect 65690 57940 65810 57950
rect 65940 57940 66060 57950
rect 66190 57940 66310 57950
rect 66440 57940 66560 57950
rect 66690 57940 66810 57950
rect 66940 57940 67060 57950
rect 67190 57940 67310 57950
rect 67440 57940 67560 57950
rect 67690 57940 67810 57950
rect 67940 57940 68060 57950
rect 68190 57940 68310 57950
rect 68440 57940 68560 57950
rect 68690 57940 68810 57950
rect 68940 57940 69060 57950
rect 69190 57940 69310 57950
rect 69440 57940 69560 57950
rect 69690 57940 69810 57950
rect 69940 57940 70060 57950
rect 70190 57940 70310 57950
rect 70440 57940 70560 57950
rect 70690 57940 70810 57950
rect 70940 57940 71000 57950
rect 59000 57810 59050 57940
rect 59200 57810 59300 57940
rect 59450 57810 59550 57940
rect 59700 57810 59800 57940
rect 59950 57810 60050 57940
rect 60200 57810 60300 57940
rect 60450 57810 60550 57940
rect 60700 57810 60800 57940
rect 60950 57810 61050 57940
rect 61200 57810 61300 57940
rect 61450 57810 61550 57940
rect 61700 57810 61800 57940
rect 61950 57810 62050 57940
rect 62200 57810 62300 57940
rect 62450 57810 62550 57940
rect 62700 57810 62800 57940
rect 62950 57810 63050 57940
rect 63200 57810 63300 57940
rect 63450 57810 63550 57940
rect 63700 57810 63800 57940
rect 63950 57810 64050 57940
rect 64200 57810 64300 57940
rect 64450 57810 64550 57940
rect 64700 57810 64800 57940
rect 64950 57810 65050 57940
rect 65200 57810 65300 57940
rect 65450 57810 65550 57940
rect 65700 57810 65800 57940
rect 65950 57810 66050 57940
rect 66200 57810 66300 57940
rect 66450 57810 66550 57940
rect 66700 57810 66800 57940
rect 66950 57810 67050 57940
rect 67200 57810 67300 57940
rect 67450 57810 67550 57940
rect 67700 57810 67800 57940
rect 67950 57810 68050 57940
rect 68200 57810 68300 57940
rect 68450 57810 68550 57940
rect 68700 57810 68800 57940
rect 68950 57810 69050 57940
rect 69200 57810 69300 57940
rect 69450 57810 69550 57940
rect 69700 57810 69800 57940
rect 69950 57810 70050 57940
rect 70200 57810 70300 57940
rect 70450 57810 70550 57940
rect 70700 57810 70800 57940
rect 70950 57810 71000 57940
rect 59000 57800 59060 57810
rect 59190 57800 59310 57810
rect 59440 57800 59560 57810
rect 59690 57800 59810 57810
rect 59940 57800 60060 57810
rect 60190 57800 60310 57810
rect 60440 57800 60560 57810
rect 60690 57800 60810 57810
rect 60940 57800 61060 57810
rect 61190 57800 61310 57810
rect 61440 57800 61560 57810
rect 61690 57800 61810 57810
rect 61940 57800 62060 57810
rect 62190 57800 62310 57810
rect 62440 57800 62560 57810
rect 62690 57800 62810 57810
rect 62940 57800 63060 57810
rect 63190 57800 63310 57810
rect 63440 57800 63560 57810
rect 63690 57800 63810 57810
rect 63940 57800 64060 57810
rect 64190 57800 64310 57810
rect 64440 57800 64560 57810
rect 64690 57800 64810 57810
rect 64940 57800 65060 57810
rect 65190 57800 65310 57810
rect 65440 57800 65560 57810
rect 65690 57800 65810 57810
rect 65940 57800 66060 57810
rect 66190 57800 66310 57810
rect 66440 57800 66560 57810
rect 66690 57800 66810 57810
rect 66940 57800 67060 57810
rect 67190 57800 67310 57810
rect 67440 57800 67560 57810
rect 67690 57800 67810 57810
rect 67940 57800 68060 57810
rect 68190 57800 68310 57810
rect 68440 57800 68560 57810
rect 68690 57800 68810 57810
rect 68940 57800 69060 57810
rect 69190 57800 69310 57810
rect 69440 57800 69560 57810
rect 69690 57800 69810 57810
rect 69940 57800 70060 57810
rect 70190 57800 70310 57810
rect 70440 57800 70560 57810
rect 70690 57800 70810 57810
rect 70940 57800 71000 57810
rect 59000 57700 71000 57800
rect 59000 57690 59060 57700
rect 59190 57690 59310 57700
rect 59440 57690 59560 57700
rect 59690 57690 59810 57700
rect 59940 57690 60060 57700
rect 60190 57690 60310 57700
rect 60440 57690 60560 57700
rect 60690 57690 60810 57700
rect 60940 57690 61060 57700
rect 61190 57690 61310 57700
rect 61440 57690 61560 57700
rect 61690 57690 61810 57700
rect 61940 57690 62060 57700
rect 62190 57690 62310 57700
rect 62440 57690 62560 57700
rect 62690 57690 62810 57700
rect 62940 57690 63060 57700
rect 63190 57690 63310 57700
rect 63440 57690 63560 57700
rect 63690 57690 63810 57700
rect 63940 57690 64060 57700
rect 64190 57690 64310 57700
rect 64440 57690 64560 57700
rect 64690 57690 64810 57700
rect 64940 57690 65060 57700
rect 65190 57690 65310 57700
rect 65440 57690 65560 57700
rect 65690 57690 65810 57700
rect 65940 57690 66060 57700
rect 66190 57690 66310 57700
rect 66440 57690 66560 57700
rect 66690 57690 66810 57700
rect 66940 57690 67060 57700
rect 67190 57690 67310 57700
rect 67440 57690 67560 57700
rect 67690 57690 67810 57700
rect 67940 57690 68060 57700
rect 68190 57690 68310 57700
rect 68440 57690 68560 57700
rect 68690 57690 68810 57700
rect 68940 57690 69060 57700
rect 69190 57690 69310 57700
rect 69440 57690 69560 57700
rect 69690 57690 69810 57700
rect 69940 57690 70060 57700
rect 70190 57690 70310 57700
rect 70440 57690 70560 57700
rect 70690 57690 70810 57700
rect 70940 57690 71000 57700
rect 59000 57560 59050 57690
rect 59200 57560 59300 57690
rect 59450 57560 59550 57690
rect 59700 57560 59800 57690
rect 59950 57560 60050 57690
rect 60200 57560 60300 57690
rect 60450 57560 60550 57690
rect 60700 57560 60800 57690
rect 60950 57560 61050 57690
rect 61200 57560 61300 57690
rect 61450 57560 61550 57690
rect 61700 57560 61800 57690
rect 61950 57560 62050 57690
rect 62200 57560 62300 57690
rect 62450 57560 62550 57690
rect 62700 57560 62800 57690
rect 62950 57560 63050 57690
rect 63200 57560 63300 57690
rect 63450 57560 63550 57690
rect 63700 57560 63800 57690
rect 63950 57560 64050 57690
rect 64200 57560 64300 57690
rect 64450 57560 64550 57690
rect 64700 57560 64800 57690
rect 64950 57560 65050 57690
rect 65200 57560 65300 57690
rect 65450 57560 65550 57690
rect 65700 57560 65800 57690
rect 65950 57560 66050 57690
rect 66200 57560 66300 57690
rect 66450 57560 66550 57690
rect 66700 57560 66800 57690
rect 66950 57560 67050 57690
rect 67200 57560 67300 57690
rect 67450 57560 67550 57690
rect 67700 57560 67800 57690
rect 67950 57560 68050 57690
rect 68200 57560 68300 57690
rect 68450 57560 68550 57690
rect 68700 57560 68800 57690
rect 68950 57560 69050 57690
rect 69200 57560 69300 57690
rect 69450 57560 69550 57690
rect 69700 57560 69800 57690
rect 69950 57560 70050 57690
rect 70200 57560 70300 57690
rect 70450 57560 70550 57690
rect 70700 57560 70800 57690
rect 70950 57560 71000 57690
rect 59000 57550 59060 57560
rect 59190 57550 59310 57560
rect 59440 57550 59560 57560
rect 59690 57550 59810 57560
rect 59940 57550 60060 57560
rect 60190 57550 60310 57560
rect 60440 57550 60560 57560
rect 60690 57550 60810 57560
rect 60940 57550 61060 57560
rect 61190 57550 61310 57560
rect 61440 57550 61560 57560
rect 61690 57550 61810 57560
rect 61940 57550 62060 57560
rect 62190 57550 62310 57560
rect 62440 57550 62560 57560
rect 62690 57550 62810 57560
rect 62940 57550 63060 57560
rect 63190 57550 63310 57560
rect 63440 57550 63560 57560
rect 63690 57550 63810 57560
rect 63940 57550 64060 57560
rect 64190 57550 64310 57560
rect 64440 57550 64560 57560
rect 64690 57550 64810 57560
rect 64940 57550 65060 57560
rect 65190 57550 65310 57560
rect 65440 57550 65560 57560
rect 65690 57550 65810 57560
rect 65940 57550 66060 57560
rect 66190 57550 66310 57560
rect 66440 57550 66560 57560
rect 66690 57550 66810 57560
rect 66940 57550 67060 57560
rect 67190 57550 67310 57560
rect 67440 57550 67560 57560
rect 67690 57550 67810 57560
rect 67940 57550 68060 57560
rect 68190 57550 68310 57560
rect 68440 57550 68560 57560
rect 68690 57550 68810 57560
rect 68940 57550 69060 57560
rect 69190 57550 69310 57560
rect 69440 57550 69560 57560
rect 69690 57550 69810 57560
rect 69940 57550 70060 57560
rect 70190 57550 70310 57560
rect 70440 57550 70560 57560
rect 70690 57550 70810 57560
rect 70940 57550 71000 57560
rect 59000 57450 71000 57550
rect 59000 57440 59060 57450
rect 59190 57440 59310 57450
rect 59440 57440 59560 57450
rect 59690 57440 59810 57450
rect 59940 57440 60060 57450
rect 60190 57440 60310 57450
rect 60440 57440 60560 57450
rect 60690 57440 60810 57450
rect 60940 57440 61060 57450
rect 61190 57440 61310 57450
rect 61440 57440 61560 57450
rect 61690 57440 61810 57450
rect 61940 57440 62060 57450
rect 62190 57440 62310 57450
rect 62440 57440 62560 57450
rect 62690 57440 62810 57450
rect 62940 57440 63060 57450
rect 63190 57440 63310 57450
rect 63440 57440 63560 57450
rect 63690 57440 63810 57450
rect 63940 57440 64060 57450
rect 64190 57440 64310 57450
rect 64440 57440 64560 57450
rect 64690 57440 64810 57450
rect 64940 57440 65060 57450
rect 65190 57440 65310 57450
rect 65440 57440 65560 57450
rect 65690 57440 65810 57450
rect 65940 57440 66060 57450
rect 66190 57440 66310 57450
rect 66440 57440 66560 57450
rect 66690 57440 66810 57450
rect 66940 57440 67060 57450
rect 67190 57440 67310 57450
rect 67440 57440 67560 57450
rect 67690 57440 67810 57450
rect 67940 57440 68060 57450
rect 68190 57440 68310 57450
rect 68440 57440 68560 57450
rect 68690 57440 68810 57450
rect 68940 57440 69060 57450
rect 69190 57440 69310 57450
rect 69440 57440 69560 57450
rect 69690 57440 69810 57450
rect 69940 57440 70060 57450
rect 70190 57440 70310 57450
rect 70440 57440 70560 57450
rect 70690 57440 70810 57450
rect 70940 57440 71000 57450
rect 59000 57310 59050 57440
rect 59200 57310 59300 57440
rect 59450 57310 59550 57440
rect 59700 57310 59800 57440
rect 59950 57310 60050 57440
rect 60200 57310 60300 57440
rect 60450 57310 60550 57440
rect 60700 57310 60800 57440
rect 60950 57310 61050 57440
rect 61200 57310 61300 57440
rect 61450 57310 61550 57440
rect 61700 57310 61800 57440
rect 61950 57310 62050 57440
rect 62200 57310 62300 57440
rect 62450 57310 62550 57440
rect 62700 57310 62800 57440
rect 62950 57310 63050 57440
rect 63200 57310 63300 57440
rect 63450 57310 63550 57440
rect 63700 57310 63800 57440
rect 63950 57310 64050 57440
rect 64200 57310 64300 57440
rect 64450 57310 64550 57440
rect 64700 57310 64800 57440
rect 64950 57310 65050 57440
rect 65200 57310 65300 57440
rect 65450 57310 65550 57440
rect 65700 57310 65800 57440
rect 65950 57310 66050 57440
rect 66200 57310 66300 57440
rect 66450 57310 66550 57440
rect 66700 57310 66800 57440
rect 66950 57310 67050 57440
rect 67200 57310 67300 57440
rect 67450 57310 67550 57440
rect 67700 57310 67800 57440
rect 67950 57310 68050 57440
rect 68200 57310 68300 57440
rect 68450 57310 68550 57440
rect 68700 57310 68800 57440
rect 68950 57310 69050 57440
rect 69200 57310 69300 57440
rect 69450 57310 69550 57440
rect 69700 57310 69800 57440
rect 69950 57310 70050 57440
rect 70200 57310 70300 57440
rect 70450 57310 70550 57440
rect 70700 57310 70800 57440
rect 70950 57310 71000 57440
rect 59000 57300 59060 57310
rect 59190 57300 59310 57310
rect 59440 57300 59560 57310
rect 59690 57300 59810 57310
rect 59940 57300 60060 57310
rect 60190 57300 60310 57310
rect 60440 57300 60560 57310
rect 60690 57300 60810 57310
rect 60940 57300 61060 57310
rect 61190 57300 61310 57310
rect 61440 57300 61560 57310
rect 61690 57300 61810 57310
rect 61940 57300 62060 57310
rect 62190 57300 62310 57310
rect 62440 57300 62560 57310
rect 62690 57300 62810 57310
rect 62940 57300 63060 57310
rect 63190 57300 63310 57310
rect 63440 57300 63560 57310
rect 63690 57300 63810 57310
rect 63940 57300 64060 57310
rect 64190 57300 64310 57310
rect 64440 57300 64560 57310
rect 64690 57300 64810 57310
rect 64940 57300 65060 57310
rect 65190 57300 65310 57310
rect 65440 57300 65560 57310
rect 65690 57300 65810 57310
rect 65940 57300 66060 57310
rect 66190 57300 66310 57310
rect 66440 57300 66560 57310
rect 66690 57300 66810 57310
rect 66940 57300 67060 57310
rect 67190 57300 67310 57310
rect 67440 57300 67560 57310
rect 67690 57300 67810 57310
rect 67940 57300 68060 57310
rect 68190 57300 68310 57310
rect 68440 57300 68560 57310
rect 68690 57300 68810 57310
rect 68940 57300 69060 57310
rect 69190 57300 69310 57310
rect 69440 57300 69560 57310
rect 69690 57300 69810 57310
rect 69940 57300 70060 57310
rect 70190 57300 70310 57310
rect 70440 57300 70560 57310
rect 70690 57300 70810 57310
rect 70940 57300 71000 57310
rect 59000 57200 71000 57300
rect 59000 57190 59060 57200
rect 59190 57190 59310 57200
rect 59440 57190 59560 57200
rect 59690 57190 59810 57200
rect 59940 57190 60060 57200
rect 60190 57190 60310 57200
rect 60440 57190 60560 57200
rect 60690 57190 60810 57200
rect 60940 57190 61060 57200
rect 61190 57190 61310 57200
rect 61440 57190 61560 57200
rect 61690 57190 61810 57200
rect 61940 57190 62060 57200
rect 62190 57190 62310 57200
rect 62440 57190 62560 57200
rect 62690 57190 62810 57200
rect 62940 57190 63060 57200
rect 63190 57190 63310 57200
rect 63440 57190 63560 57200
rect 63690 57190 63810 57200
rect 63940 57190 64060 57200
rect 64190 57190 64310 57200
rect 64440 57190 64560 57200
rect 64690 57190 64810 57200
rect 64940 57190 65060 57200
rect 65190 57190 65310 57200
rect 65440 57190 65560 57200
rect 65690 57190 65810 57200
rect 65940 57190 66060 57200
rect 66190 57190 66310 57200
rect 66440 57190 66560 57200
rect 66690 57190 66810 57200
rect 66940 57190 67060 57200
rect 67190 57190 67310 57200
rect 67440 57190 67560 57200
rect 67690 57190 67810 57200
rect 67940 57190 68060 57200
rect 68190 57190 68310 57200
rect 68440 57190 68560 57200
rect 68690 57190 68810 57200
rect 68940 57190 69060 57200
rect 69190 57190 69310 57200
rect 69440 57190 69560 57200
rect 69690 57190 69810 57200
rect 69940 57190 70060 57200
rect 70190 57190 70310 57200
rect 70440 57190 70560 57200
rect 70690 57190 70810 57200
rect 70940 57190 71000 57200
rect 59000 57060 59050 57190
rect 59200 57060 59300 57190
rect 59450 57060 59550 57190
rect 59700 57060 59800 57190
rect 59950 57060 60050 57190
rect 60200 57060 60300 57190
rect 60450 57060 60550 57190
rect 60700 57060 60800 57190
rect 60950 57060 61050 57190
rect 61200 57060 61300 57190
rect 61450 57060 61550 57190
rect 61700 57060 61800 57190
rect 61950 57060 62050 57190
rect 62200 57060 62300 57190
rect 62450 57060 62550 57190
rect 62700 57060 62800 57190
rect 62950 57060 63050 57190
rect 63200 57060 63300 57190
rect 63450 57060 63550 57190
rect 63700 57060 63800 57190
rect 63950 57060 64050 57190
rect 64200 57060 64300 57190
rect 64450 57060 64550 57190
rect 64700 57060 64800 57190
rect 64950 57060 65050 57190
rect 65200 57060 65300 57190
rect 65450 57060 65550 57190
rect 65700 57060 65800 57190
rect 65950 57060 66050 57190
rect 66200 57060 66300 57190
rect 66450 57060 66550 57190
rect 66700 57060 66800 57190
rect 66950 57060 67050 57190
rect 67200 57060 67300 57190
rect 67450 57060 67550 57190
rect 67700 57060 67800 57190
rect 67950 57060 68050 57190
rect 68200 57060 68300 57190
rect 68450 57060 68550 57190
rect 68700 57060 68800 57190
rect 68950 57060 69050 57190
rect 69200 57060 69300 57190
rect 69450 57060 69550 57190
rect 69700 57060 69800 57190
rect 69950 57060 70050 57190
rect 70200 57060 70300 57190
rect 70450 57060 70550 57190
rect 70700 57060 70800 57190
rect 70950 57060 71000 57190
rect 59000 57050 59060 57060
rect 59190 57050 59310 57060
rect 59440 57050 59560 57060
rect 59690 57050 59810 57060
rect 59940 57050 60060 57060
rect 60190 57050 60310 57060
rect 60440 57050 60560 57060
rect 60690 57050 60810 57060
rect 60940 57050 61060 57060
rect 61190 57050 61310 57060
rect 61440 57050 61560 57060
rect 61690 57050 61810 57060
rect 61940 57050 62060 57060
rect 62190 57050 62310 57060
rect 62440 57050 62560 57060
rect 62690 57050 62810 57060
rect 62940 57050 63060 57060
rect 63190 57050 63310 57060
rect 63440 57050 63560 57060
rect 63690 57050 63810 57060
rect 63940 57050 64060 57060
rect 64190 57050 64310 57060
rect 64440 57050 64560 57060
rect 64690 57050 64810 57060
rect 64940 57050 65060 57060
rect 65190 57050 65310 57060
rect 65440 57050 65560 57060
rect 65690 57050 65810 57060
rect 65940 57050 66060 57060
rect 66190 57050 66310 57060
rect 66440 57050 66560 57060
rect 66690 57050 66810 57060
rect 66940 57050 67060 57060
rect 67190 57050 67310 57060
rect 67440 57050 67560 57060
rect 67690 57050 67810 57060
rect 67940 57050 68060 57060
rect 68190 57050 68310 57060
rect 68440 57050 68560 57060
rect 68690 57050 68810 57060
rect 68940 57050 69060 57060
rect 69190 57050 69310 57060
rect 69440 57050 69560 57060
rect 69690 57050 69810 57060
rect 69940 57050 70060 57060
rect 70190 57050 70310 57060
rect 70440 57050 70560 57060
rect 70690 57050 70810 57060
rect 70940 57050 71000 57060
rect 59000 57000 71000 57050
rect 81000 60950 92000 61000
rect 81000 60940 81060 60950
rect 81190 60940 81310 60950
rect 81440 60940 81560 60950
rect 81690 60940 81810 60950
rect 81940 60940 82060 60950
rect 82190 60940 82310 60950
rect 82440 60940 82560 60950
rect 82690 60940 82810 60950
rect 82940 60940 83060 60950
rect 83190 60940 83310 60950
rect 83440 60940 83560 60950
rect 83690 60940 83810 60950
rect 83940 60940 84060 60950
rect 84190 60940 84310 60950
rect 84440 60940 84560 60950
rect 84690 60940 84810 60950
rect 84940 60940 85060 60950
rect 85190 60940 85310 60950
rect 85440 60940 85560 60950
rect 85690 60940 85810 60950
rect 85940 60940 86060 60950
rect 86190 60940 86310 60950
rect 86440 60940 86560 60950
rect 86690 60940 86810 60950
rect 86940 60940 87060 60950
rect 87190 60940 87310 60950
rect 87440 60940 87560 60950
rect 87690 60940 87810 60950
rect 87940 60940 88060 60950
rect 88190 60940 88310 60950
rect 88440 60940 88560 60950
rect 88690 60940 88810 60950
rect 88940 60940 89060 60950
rect 89190 60940 89310 60950
rect 89440 60940 89560 60950
rect 89690 60940 89810 60950
rect 89940 60940 90060 60950
rect 90190 60940 90310 60950
rect 90440 60940 90560 60950
rect 90690 60940 90810 60950
rect 90940 60940 91060 60950
rect 91190 60940 91310 60950
rect 91440 60940 91560 60950
rect 91690 60940 91810 60950
rect 91940 60940 92000 60950
rect 81000 60810 81050 60940
rect 81200 60810 81300 60940
rect 81450 60810 81550 60940
rect 81700 60810 81800 60940
rect 81950 60810 82050 60940
rect 82200 60810 82300 60940
rect 82450 60810 82550 60940
rect 82700 60810 82800 60940
rect 82950 60810 83050 60940
rect 83200 60810 83300 60940
rect 83450 60810 83550 60940
rect 83700 60810 83800 60940
rect 83950 60810 84050 60940
rect 84200 60810 84300 60940
rect 84450 60810 84550 60940
rect 84700 60810 84800 60940
rect 84950 60810 85050 60940
rect 85200 60810 85300 60940
rect 85450 60810 85550 60940
rect 85700 60810 85800 60940
rect 85950 60810 86050 60940
rect 86200 60810 86300 60940
rect 86450 60810 86550 60940
rect 86700 60810 86800 60940
rect 86950 60810 87050 60940
rect 87200 60810 87300 60940
rect 87450 60810 87550 60940
rect 87700 60810 87800 60940
rect 87950 60810 88050 60940
rect 88200 60810 88300 60940
rect 88450 60810 88550 60940
rect 88700 60810 88800 60940
rect 88950 60810 89050 60940
rect 89200 60810 89300 60940
rect 89450 60810 89550 60940
rect 89700 60810 89800 60940
rect 89950 60810 90050 60940
rect 90200 60810 90300 60940
rect 90450 60810 90550 60940
rect 90700 60810 90800 60940
rect 90950 60810 91050 60940
rect 91200 60810 91300 60940
rect 91450 60810 91550 60940
rect 91700 60810 91800 60940
rect 91950 60810 92000 60940
rect 81000 60800 81060 60810
rect 81190 60800 81310 60810
rect 81440 60800 81560 60810
rect 81690 60800 81810 60810
rect 81940 60800 82060 60810
rect 82190 60800 82310 60810
rect 82440 60800 82560 60810
rect 82690 60800 82810 60810
rect 82940 60800 83060 60810
rect 83190 60800 83310 60810
rect 83440 60800 83560 60810
rect 83690 60800 83810 60810
rect 83940 60800 84060 60810
rect 84190 60800 84310 60810
rect 84440 60800 84560 60810
rect 84690 60800 84810 60810
rect 84940 60800 85060 60810
rect 85190 60800 85310 60810
rect 85440 60800 85560 60810
rect 85690 60800 85810 60810
rect 85940 60800 86060 60810
rect 86190 60800 86310 60810
rect 86440 60800 86560 60810
rect 86690 60800 86810 60810
rect 86940 60800 87060 60810
rect 87190 60800 87310 60810
rect 87440 60800 87560 60810
rect 87690 60800 87810 60810
rect 87940 60800 88060 60810
rect 88190 60800 88310 60810
rect 88440 60800 88560 60810
rect 88690 60800 88810 60810
rect 88940 60800 89060 60810
rect 89190 60800 89310 60810
rect 89440 60800 89560 60810
rect 89690 60800 89810 60810
rect 89940 60800 90060 60810
rect 90190 60800 90310 60810
rect 90440 60800 90560 60810
rect 90690 60800 90810 60810
rect 90940 60800 91060 60810
rect 91190 60800 91310 60810
rect 91440 60800 91560 60810
rect 91690 60800 91810 60810
rect 91940 60800 92000 60810
rect 81000 60700 92000 60800
rect 81000 60690 81060 60700
rect 81190 60690 81310 60700
rect 81440 60690 81560 60700
rect 81690 60690 81810 60700
rect 81940 60690 82060 60700
rect 82190 60690 82310 60700
rect 82440 60690 82560 60700
rect 82690 60690 82810 60700
rect 82940 60690 83060 60700
rect 83190 60690 83310 60700
rect 83440 60690 83560 60700
rect 83690 60690 83810 60700
rect 83940 60690 84060 60700
rect 84190 60690 84310 60700
rect 84440 60690 84560 60700
rect 84690 60690 84810 60700
rect 84940 60690 85060 60700
rect 85190 60690 85310 60700
rect 85440 60690 85560 60700
rect 85690 60690 85810 60700
rect 85940 60690 86060 60700
rect 86190 60690 86310 60700
rect 86440 60690 86560 60700
rect 86690 60690 86810 60700
rect 86940 60690 87060 60700
rect 87190 60690 87310 60700
rect 87440 60690 87560 60700
rect 87690 60690 87810 60700
rect 87940 60690 88060 60700
rect 88190 60690 88310 60700
rect 88440 60690 88560 60700
rect 88690 60690 88810 60700
rect 88940 60690 89060 60700
rect 89190 60690 89310 60700
rect 89440 60690 89560 60700
rect 89690 60690 89810 60700
rect 89940 60690 90060 60700
rect 90190 60690 90310 60700
rect 90440 60690 90560 60700
rect 90690 60690 90810 60700
rect 90940 60690 91060 60700
rect 91190 60690 91310 60700
rect 91440 60690 91560 60700
rect 91690 60690 91810 60700
rect 91940 60690 92000 60700
rect 81000 60560 81050 60690
rect 81200 60560 81300 60690
rect 81450 60560 81550 60690
rect 81700 60560 81800 60690
rect 81950 60560 82050 60690
rect 82200 60560 82300 60690
rect 82450 60560 82550 60690
rect 82700 60560 82800 60690
rect 82950 60560 83050 60690
rect 83200 60560 83300 60690
rect 83450 60560 83550 60690
rect 83700 60560 83800 60690
rect 83950 60560 84050 60690
rect 84200 60560 84300 60690
rect 84450 60560 84550 60690
rect 84700 60560 84800 60690
rect 84950 60560 85050 60690
rect 85200 60560 85300 60690
rect 85450 60560 85550 60690
rect 85700 60560 85800 60690
rect 85950 60560 86050 60690
rect 86200 60560 86300 60690
rect 86450 60560 86550 60690
rect 86700 60560 86800 60690
rect 86950 60560 87050 60690
rect 87200 60560 87300 60690
rect 87450 60560 87550 60690
rect 87700 60560 87800 60690
rect 87950 60560 88050 60690
rect 88200 60560 88300 60690
rect 88450 60560 88550 60690
rect 88700 60560 88800 60690
rect 88950 60560 89050 60690
rect 89200 60560 89300 60690
rect 89450 60560 89550 60690
rect 89700 60560 89800 60690
rect 89950 60560 90050 60690
rect 90200 60560 90300 60690
rect 90450 60560 90550 60690
rect 90700 60560 90800 60690
rect 90950 60560 91050 60690
rect 91200 60560 91300 60690
rect 91450 60560 91550 60690
rect 91700 60560 91800 60690
rect 91950 60560 92000 60690
rect 81000 60550 81060 60560
rect 81190 60550 81310 60560
rect 81440 60550 81560 60560
rect 81690 60550 81810 60560
rect 81940 60550 82060 60560
rect 82190 60550 82310 60560
rect 82440 60550 82560 60560
rect 82690 60550 82810 60560
rect 82940 60550 83060 60560
rect 83190 60550 83310 60560
rect 83440 60550 83560 60560
rect 83690 60550 83810 60560
rect 83940 60550 84060 60560
rect 84190 60550 84310 60560
rect 84440 60550 84560 60560
rect 84690 60550 84810 60560
rect 84940 60550 85060 60560
rect 85190 60550 85310 60560
rect 85440 60550 85560 60560
rect 85690 60550 85810 60560
rect 85940 60550 86060 60560
rect 86190 60550 86310 60560
rect 86440 60550 86560 60560
rect 86690 60550 86810 60560
rect 86940 60550 87060 60560
rect 87190 60550 87310 60560
rect 87440 60550 87560 60560
rect 87690 60550 87810 60560
rect 87940 60550 88060 60560
rect 88190 60550 88310 60560
rect 88440 60550 88560 60560
rect 88690 60550 88810 60560
rect 88940 60550 89060 60560
rect 89190 60550 89310 60560
rect 89440 60550 89560 60560
rect 89690 60550 89810 60560
rect 89940 60550 90060 60560
rect 90190 60550 90310 60560
rect 90440 60550 90560 60560
rect 90690 60550 90810 60560
rect 90940 60550 91060 60560
rect 91190 60550 91310 60560
rect 91440 60550 91560 60560
rect 91690 60550 91810 60560
rect 91940 60550 92000 60560
rect 81000 60450 92000 60550
rect 81000 60440 81060 60450
rect 81190 60440 81310 60450
rect 81440 60440 81560 60450
rect 81690 60440 81810 60450
rect 81940 60440 82060 60450
rect 82190 60440 82310 60450
rect 82440 60440 82560 60450
rect 82690 60440 82810 60450
rect 82940 60440 83060 60450
rect 83190 60440 83310 60450
rect 83440 60440 83560 60450
rect 83690 60440 83810 60450
rect 83940 60440 84060 60450
rect 84190 60440 84310 60450
rect 84440 60440 84560 60450
rect 84690 60440 84810 60450
rect 84940 60440 85060 60450
rect 85190 60440 85310 60450
rect 85440 60440 85560 60450
rect 85690 60440 85810 60450
rect 85940 60440 86060 60450
rect 86190 60440 86310 60450
rect 86440 60440 86560 60450
rect 86690 60440 86810 60450
rect 86940 60440 87060 60450
rect 87190 60440 87310 60450
rect 87440 60440 87560 60450
rect 87690 60440 87810 60450
rect 87940 60440 88060 60450
rect 88190 60440 88310 60450
rect 88440 60440 88560 60450
rect 88690 60440 88810 60450
rect 88940 60440 89060 60450
rect 89190 60440 89310 60450
rect 89440 60440 89560 60450
rect 89690 60440 89810 60450
rect 89940 60440 90060 60450
rect 90190 60440 90310 60450
rect 90440 60440 90560 60450
rect 90690 60440 90810 60450
rect 90940 60440 91060 60450
rect 91190 60440 91310 60450
rect 91440 60440 91560 60450
rect 91690 60440 91810 60450
rect 91940 60440 92000 60450
rect 81000 60310 81050 60440
rect 81200 60310 81300 60440
rect 81450 60310 81550 60440
rect 81700 60310 81800 60440
rect 81950 60310 82050 60440
rect 82200 60310 82300 60440
rect 82450 60310 82550 60440
rect 82700 60310 82800 60440
rect 82950 60310 83050 60440
rect 83200 60310 83300 60440
rect 83450 60310 83550 60440
rect 83700 60310 83800 60440
rect 83950 60310 84050 60440
rect 84200 60310 84300 60440
rect 84450 60310 84550 60440
rect 84700 60310 84800 60440
rect 84950 60310 85050 60440
rect 85200 60310 85300 60440
rect 85450 60310 85550 60440
rect 85700 60310 85800 60440
rect 85950 60310 86050 60440
rect 86200 60310 86300 60440
rect 86450 60310 86550 60440
rect 86700 60310 86800 60440
rect 86950 60310 87050 60440
rect 87200 60310 87300 60440
rect 87450 60310 87550 60440
rect 87700 60310 87800 60440
rect 87950 60310 88050 60440
rect 88200 60310 88300 60440
rect 88450 60310 88550 60440
rect 88700 60310 88800 60440
rect 88950 60310 89050 60440
rect 89200 60310 89300 60440
rect 89450 60310 89550 60440
rect 89700 60310 89800 60440
rect 89950 60310 90050 60440
rect 90200 60310 90300 60440
rect 90450 60310 90550 60440
rect 90700 60310 90800 60440
rect 90950 60310 91050 60440
rect 91200 60310 91300 60440
rect 91450 60310 91550 60440
rect 91700 60310 91800 60440
rect 91950 60310 92000 60440
rect 81000 60300 81060 60310
rect 81190 60300 81310 60310
rect 81440 60300 81560 60310
rect 81690 60300 81810 60310
rect 81940 60300 82060 60310
rect 82190 60300 82310 60310
rect 82440 60300 82560 60310
rect 82690 60300 82810 60310
rect 82940 60300 83060 60310
rect 83190 60300 83310 60310
rect 83440 60300 83560 60310
rect 83690 60300 83810 60310
rect 83940 60300 84060 60310
rect 84190 60300 84310 60310
rect 84440 60300 84560 60310
rect 84690 60300 84810 60310
rect 84940 60300 85060 60310
rect 85190 60300 85310 60310
rect 85440 60300 85560 60310
rect 85690 60300 85810 60310
rect 85940 60300 86060 60310
rect 86190 60300 86310 60310
rect 86440 60300 86560 60310
rect 86690 60300 86810 60310
rect 86940 60300 87060 60310
rect 87190 60300 87310 60310
rect 87440 60300 87560 60310
rect 87690 60300 87810 60310
rect 87940 60300 88060 60310
rect 88190 60300 88310 60310
rect 88440 60300 88560 60310
rect 88690 60300 88810 60310
rect 88940 60300 89060 60310
rect 89190 60300 89310 60310
rect 89440 60300 89560 60310
rect 89690 60300 89810 60310
rect 89940 60300 90060 60310
rect 90190 60300 90310 60310
rect 90440 60300 90560 60310
rect 90690 60300 90810 60310
rect 90940 60300 91060 60310
rect 91190 60300 91310 60310
rect 91440 60300 91560 60310
rect 91690 60300 91810 60310
rect 91940 60300 92000 60310
rect 81000 60200 92000 60300
rect 81000 60190 81060 60200
rect 81190 60190 81310 60200
rect 81440 60190 81560 60200
rect 81690 60190 81810 60200
rect 81940 60190 82060 60200
rect 82190 60190 82310 60200
rect 82440 60190 82560 60200
rect 82690 60190 82810 60200
rect 82940 60190 83060 60200
rect 83190 60190 83310 60200
rect 83440 60190 83560 60200
rect 83690 60190 83810 60200
rect 83940 60190 84060 60200
rect 84190 60190 84310 60200
rect 84440 60190 84560 60200
rect 84690 60190 84810 60200
rect 84940 60190 85060 60200
rect 85190 60190 85310 60200
rect 85440 60190 85560 60200
rect 85690 60190 85810 60200
rect 85940 60190 86060 60200
rect 86190 60190 86310 60200
rect 86440 60190 86560 60200
rect 86690 60190 86810 60200
rect 86940 60190 87060 60200
rect 87190 60190 87310 60200
rect 87440 60190 87560 60200
rect 87690 60190 87810 60200
rect 87940 60190 88060 60200
rect 88190 60190 88310 60200
rect 88440 60190 88560 60200
rect 88690 60190 88810 60200
rect 88940 60190 89060 60200
rect 89190 60190 89310 60200
rect 89440 60190 89560 60200
rect 89690 60190 89810 60200
rect 89940 60190 90060 60200
rect 90190 60190 90310 60200
rect 90440 60190 90560 60200
rect 90690 60190 90810 60200
rect 90940 60190 91060 60200
rect 91190 60190 91310 60200
rect 91440 60190 91560 60200
rect 91690 60190 91810 60200
rect 91940 60190 92000 60200
rect 81000 60060 81050 60190
rect 81200 60060 81300 60190
rect 81450 60060 81550 60190
rect 81700 60060 81800 60190
rect 81950 60060 82050 60190
rect 82200 60060 82300 60190
rect 82450 60060 82550 60190
rect 82700 60060 82800 60190
rect 82950 60060 83050 60190
rect 83200 60060 83300 60190
rect 83450 60060 83550 60190
rect 83700 60060 83800 60190
rect 83950 60060 84050 60190
rect 84200 60060 84300 60190
rect 84450 60060 84550 60190
rect 84700 60060 84800 60190
rect 84950 60060 85050 60190
rect 85200 60060 85300 60190
rect 85450 60060 85550 60190
rect 85700 60060 85800 60190
rect 85950 60060 86050 60190
rect 86200 60060 86300 60190
rect 86450 60060 86550 60190
rect 86700 60060 86800 60190
rect 86950 60060 87050 60190
rect 87200 60060 87300 60190
rect 87450 60060 87550 60190
rect 87700 60060 87800 60190
rect 87950 60060 88050 60190
rect 88200 60060 88300 60190
rect 88450 60060 88550 60190
rect 88700 60060 88800 60190
rect 88950 60060 89050 60190
rect 89200 60060 89300 60190
rect 89450 60060 89550 60190
rect 89700 60060 89800 60190
rect 89950 60060 90050 60190
rect 90200 60060 90300 60190
rect 90450 60060 90550 60190
rect 90700 60060 90800 60190
rect 90950 60060 91050 60190
rect 91200 60060 91300 60190
rect 91450 60060 91550 60190
rect 91700 60060 91800 60190
rect 91950 60060 92000 60190
rect 81000 60050 81060 60060
rect 81190 60050 81310 60060
rect 81440 60050 81560 60060
rect 81690 60050 81810 60060
rect 81940 60050 82060 60060
rect 82190 60050 82310 60060
rect 82440 60050 82560 60060
rect 82690 60050 82810 60060
rect 82940 60050 83060 60060
rect 83190 60050 83310 60060
rect 83440 60050 83560 60060
rect 83690 60050 83810 60060
rect 83940 60050 84060 60060
rect 84190 60050 84310 60060
rect 84440 60050 84560 60060
rect 84690 60050 84810 60060
rect 84940 60050 85060 60060
rect 85190 60050 85310 60060
rect 85440 60050 85560 60060
rect 85690 60050 85810 60060
rect 85940 60050 86060 60060
rect 86190 60050 86310 60060
rect 86440 60050 86560 60060
rect 86690 60050 86810 60060
rect 86940 60050 87060 60060
rect 87190 60050 87310 60060
rect 87440 60050 87560 60060
rect 87690 60050 87810 60060
rect 87940 60050 88060 60060
rect 88190 60050 88310 60060
rect 88440 60050 88560 60060
rect 88690 60050 88810 60060
rect 88940 60050 89060 60060
rect 89190 60050 89310 60060
rect 89440 60050 89560 60060
rect 89690 60050 89810 60060
rect 89940 60050 90060 60060
rect 90190 60050 90310 60060
rect 90440 60050 90560 60060
rect 90690 60050 90810 60060
rect 90940 60050 91060 60060
rect 91190 60050 91310 60060
rect 91440 60050 91560 60060
rect 91690 60050 91810 60060
rect 91940 60050 92000 60060
rect 81000 59950 92000 60050
rect 81000 59940 81060 59950
rect 81190 59940 81310 59950
rect 81440 59940 81560 59950
rect 81690 59940 81810 59950
rect 81940 59940 82060 59950
rect 82190 59940 82310 59950
rect 82440 59940 82560 59950
rect 82690 59940 82810 59950
rect 82940 59940 83060 59950
rect 83190 59940 83310 59950
rect 83440 59940 83560 59950
rect 83690 59940 83810 59950
rect 83940 59940 84060 59950
rect 84190 59940 84310 59950
rect 84440 59940 84560 59950
rect 84690 59940 84810 59950
rect 84940 59940 85060 59950
rect 85190 59940 85310 59950
rect 85440 59940 85560 59950
rect 85690 59940 85810 59950
rect 85940 59940 86060 59950
rect 86190 59940 86310 59950
rect 86440 59940 86560 59950
rect 86690 59940 86810 59950
rect 86940 59940 87060 59950
rect 87190 59940 87310 59950
rect 87440 59940 87560 59950
rect 87690 59940 87810 59950
rect 87940 59940 88060 59950
rect 88190 59940 88310 59950
rect 88440 59940 88560 59950
rect 88690 59940 88810 59950
rect 88940 59940 89060 59950
rect 89190 59940 89310 59950
rect 89440 59940 89560 59950
rect 89690 59940 89810 59950
rect 89940 59940 90060 59950
rect 90190 59940 90310 59950
rect 90440 59940 90560 59950
rect 90690 59940 90810 59950
rect 90940 59940 91060 59950
rect 91190 59940 91310 59950
rect 91440 59940 91560 59950
rect 91690 59940 91810 59950
rect 91940 59940 92000 59950
rect 81000 59810 81050 59940
rect 81200 59810 81300 59940
rect 81450 59810 81550 59940
rect 81700 59810 81800 59940
rect 81950 59810 82050 59940
rect 82200 59810 82300 59940
rect 82450 59810 82550 59940
rect 82700 59810 82800 59940
rect 82950 59810 83050 59940
rect 83200 59810 83300 59940
rect 83450 59810 83550 59940
rect 83700 59810 83800 59940
rect 83950 59810 84050 59940
rect 84200 59810 84300 59940
rect 84450 59810 84550 59940
rect 84700 59810 84800 59940
rect 84950 59810 85050 59940
rect 85200 59810 85300 59940
rect 85450 59810 85550 59940
rect 85700 59810 85800 59940
rect 85950 59810 86050 59940
rect 86200 59810 86300 59940
rect 86450 59810 86550 59940
rect 86700 59810 86800 59940
rect 86950 59810 87050 59940
rect 87200 59810 87300 59940
rect 87450 59810 87550 59940
rect 87700 59810 87800 59940
rect 87950 59810 88050 59940
rect 88200 59810 88300 59940
rect 88450 59810 88550 59940
rect 88700 59810 88800 59940
rect 88950 59810 89050 59940
rect 89200 59810 89300 59940
rect 89450 59810 89550 59940
rect 89700 59810 89800 59940
rect 89950 59810 90050 59940
rect 90200 59810 90300 59940
rect 90450 59810 90550 59940
rect 90700 59810 90800 59940
rect 90950 59810 91050 59940
rect 91200 59810 91300 59940
rect 91450 59810 91550 59940
rect 91700 59810 91800 59940
rect 91950 59810 92000 59940
rect 81000 59800 81060 59810
rect 81190 59800 81310 59810
rect 81440 59800 81560 59810
rect 81690 59800 81810 59810
rect 81940 59800 82060 59810
rect 82190 59800 82310 59810
rect 82440 59800 82560 59810
rect 82690 59800 82810 59810
rect 82940 59800 83060 59810
rect 83190 59800 83310 59810
rect 83440 59800 83560 59810
rect 83690 59800 83810 59810
rect 83940 59800 84060 59810
rect 84190 59800 84310 59810
rect 84440 59800 84560 59810
rect 84690 59800 84810 59810
rect 84940 59800 85060 59810
rect 85190 59800 85310 59810
rect 85440 59800 85560 59810
rect 85690 59800 85810 59810
rect 85940 59800 86060 59810
rect 86190 59800 86310 59810
rect 86440 59800 86560 59810
rect 86690 59800 86810 59810
rect 86940 59800 87060 59810
rect 87190 59800 87310 59810
rect 87440 59800 87560 59810
rect 87690 59800 87810 59810
rect 87940 59800 88060 59810
rect 88190 59800 88310 59810
rect 88440 59800 88560 59810
rect 88690 59800 88810 59810
rect 88940 59800 89060 59810
rect 89190 59800 89310 59810
rect 89440 59800 89560 59810
rect 89690 59800 89810 59810
rect 89940 59800 90060 59810
rect 90190 59800 90310 59810
rect 90440 59800 90560 59810
rect 90690 59800 90810 59810
rect 90940 59800 91060 59810
rect 91190 59800 91310 59810
rect 91440 59800 91560 59810
rect 91690 59800 91810 59810
rect 91940 59800 92000 59810
rect 81000 59700 92000 59800
rect 81000 59690 81060 59700
rect 81190 59690 81310 59700
rect 81440 59690 81560 59700
rect 81690 59690 81810 59700
rect 81940 59690 82060 59700
rect 82190 59690 82310 59700
rect 82440 59690 82560 59700
rect 82690 59690 82810 59700
rect 82940 59690 83060 59700
rect 83190 59690 83310 59700
rect 83440 59690 83560 59700
rect 83690 59690 83810 59700
rect 83940 59690 84060 59700
rect 84190 59690 84310 59700
rect 84440 59690 84560 59700
rect 84690 59690 84810 59700
rect 84940 59690 85060 59700
rect 85190 59690 85310 59700
rect 85440 59690 85560 59700
rect 85690 59690 85810 59700
rect 85940 59690 86060 59700
rect 86190 59690 86310 59700
rect 86440 59690 86560 59700
rect 86690 59690 86810 59700
rect 86940 59690 87060 59700
rect 87190 59690 87310 59700
rect 87440 59690 87560 59700
rect 87690 59690 87810 59700
rect 87940 59690 88060 59700
rect 88190 59690 88310 59700
rect 88440 59690 88560 59700
rect 88690 59690 88810 59700
rect 88940 59690 89060 59700
rect 89190 59690 89310 59700
rect 89440 59690 89560 59700
rect 89690 59690 89810 59700
rect 89940 59690 90060 59700
rect 90190 59690 90310 59700
rect 90440 59690 90560 59700
rect 90690 59690 90810 59700
rect 90940 59690 91060 59700
rect 91190 59690 91310 59700
rect 91440 59690 91560 59700
rect 91690 59690 91810 59700
rect 91940 59690 92000 59700
rect 81000 59560 81050 59690
rect 81200 59560 81300 59690
rect 81450 59560 81550 59690
rect 81700 59560 81800 59690
rect 81950 59560 82050 59690
rect 82200 59560 82300 59690
rect 82450 59560 82550 59690
rect 82700 59560 82800 59690
rect 82950 59560 83050 59690
rect 83200 59560 83300 59690
rect 83450 59560 83550 59690
rect 83700 59560 83800 59690
rect 83950 59560 84050 59690
rect 84200 59560 84300 59690
rect 84450 59560 84550 59690
rect 84700 59560 84800 59690
rect 84950 59560 85050 59690
rect 85200 59560 85300 59690
rect 85450 59560 85550 59690
rect 85700 59560 85800 59690
rect 85950 59560 86050 59690
rect 86200 59560 86300 59690
rect 86450 59560 86550 59690
rect 86700 59560 86800 59690
rect 86950 59560 87050 59690
rect 87200 59560 87300 59690
rect 87450 59560 87550 59690
rect 87700 59560 87800 59690
rect 87950 59560 88050 59690
rect 88200 59560 88300 59690
rect 88450 59560 88550 59690
rect 88700 59560 88800 59690
rect 88950 59560 89050 59690
rect 89200 59560 89300 59690
rect 89450 59560 89550 59690
rect 89700 59560 89800 59690
rect 89950 59560 90050 59690
rect 90200 59560 90300 59690
rect 90450 59560 90550 59690
rect 90700 59560 90800 59690
rect 90950 59560 91050 59690
rect 91200 59560 91300 59690
rect 91450 59560 91550 59690
rect 91700 59560 91800 59690
rect 91950 59560 92000 59690
rect 81000 59550 81060 59560
rect 81190 59550 81310 59560
rect 81440 59550 81560 59560
rect 81690 59550 81810 59560
rect 81940 59550 82060 59560
rect 82190 59550 82310 59560
rect 82440 59550 82560 59560
rect 82690 59550 82810 59560
rect 82940 59550 83060 59560
rect 83190 59550 83310 59560
rect 83440 59550 83560 59560
rect 83690 59550 83810 59560
rect 83940 59550 84060 59560
rect 84190 59550 84310 59560
rect 84440 59550 84560 59560
rect 84690 59550 84810 59560
rect 84940 59550 85060 59560
rect 85190 59550 85310 59560
rect 85440 59550 85560 59560
rect 85690 59550 85810 59560
rect 85940 59550 86060 59560
rect 86190 59550 86310 59560
rect 86440 59550 86560 59560
rect 86690 59550 86810 59560
rect 86940 59550 87060 59560
rect 87190 59550 87310 59560
rect 87440 59550 87560 59560
rect 87690 59550 87810 59560
rect 87940 59550 88060 59560
rect 88190 59550 88310 59560
rect 88440 59550 88560 59560
rect 88690 59550 88810 59560
rect 88940 59550 89060 59560
rect 89190 59550 89310 59560
rect 89440 59550 89560 59560
rect 89690 59550 89810 59560
rect 89940 59550 90060 59560
rect 90190 59550 90310 59560
rect 90440 59550 90560 59560
rect 90690 59550 90810 59560
rect 90940 59550 91060 59560
rect 91190 59550 91310 59560
rect 91440 59550 91560 59560
rect 91690 59550 91810 59560
rect 91940 59550 92000 59560
rect 81000 59450 92000 59550
rect 81000 59440 81060 59450
rect 81190 59440 81310 59450
rect 81440 59440 81560 59450
rect 81690 59440 81810 59450
rect 81940 59440 82060 59450
rect 82190 59440 82310 59450
rect 82440 59440 82560 59450
rect 82690 59440 82810 59450
rect 82940 59440 83060 59450
rect 83190 59440 83310 59450
rect 83440 59440 83560 59450
rect 83690 59440 83810 59450
rect 83940 59440 84060 59450
rect 84190 59440 84310 59450
rect 84440 59440 84560 59450
rect 84690 59440 84810 59450
rect 84940 59440 85060 59450
rect 85190 59440 85310 59450
rect 85440 59440 85560 59450
rect 85690 59440 85810 59450
rect 85940 59440 86060 59450
rect 86190 59440 86310 59450
rect 86440 59440 86560 59450
rect 86690 59440 86810 59450
rect 86940 59440 87060 59450
rect 87190 59440 87310 59450
rect 87440 59440 87560 59450
rect 87690 59440 87810 59450
rect 87940 59440 88060 59450
rect 88190 59440 88310 59450
rect 88440 59440 88560 59450
rect 88690 59440 88810 59450
rect 88940 59440 89060 59450
rect 89190 59440 89310 59450
rect 89440 59440 89560 59450
rect 89690 59440 89810 59450
rect 89940 59440 90060 59450
rect 90190 59440 90310 59450
rect 90440 59440 90560 59450
rect 90690 59440 90810 59450
rect 90940 59440 91060 59450
rect 91190 59440 91310 59450
rect 91440 59440 91560 59450
rect 91690 59440 91810 59450
rect 91940 59440 92000 59450
rect 81000 59310 81050 59440
rect 81200 59310 81300 59440
rect 81450 59310 81550 59440
rect 81700 59310 81800 59440
rect 81950 59310 82050 59440
rect 82200 59310 82300 59440
rect 82450 59310 82550 59440
rect 82700 59310 82800 59440
rect 82950 59310 83050 59440
rect 83200 59310 83300 59440
rect 83450 59310 83550 59440
rect 83700 59310 83800 59440
rect 83950 59310 84050 59440
rect 84200 59310 84300 59440
rect 84450 59310 84550 59440
rect 84700 59310 84800 59440
rect 84950 59310 85050 59440
rect 85200 59310 85300 59440
rect 85450 59310 85550 59440
rect 85700 59310 85800 59440
rect 85950 59310 86050 59440
rect 86200 59310 86300 59440
rect 86450 59310 86550 59440
rect 86700 59310 86800 59440
rect 86950 59310 87050 59440
rect 87200 59310 87300 59440
rect 87450 59310 87550 59440
rect 87700 59310 87800 59440
rect 87950 59310 88050 59440
rect 88200 59310 88300 59440
rect 88450 59310 88550 59440
rect 88700 59310 88800 59440
rect 88950 59310 89050 59440
rect 89200 59310 89300 59440
rect 89450 59310 89550 59440
rect 89700 59310 89800 59440
rect 89950 59310 90050 59440
rect 90200 59310 90300 59440
rect 90450 59310 90550 59440
rect 90700 59310 90800 59440
rect 90950 59310 91050 59440
rect 91200 59310 91300 59440
rect 91450 59310 91550 59440
rect 91700 59310 91800 59440
rect 91950 59310 92000 59440
rect 81000 59300 81060 59310
rect 81190 59300 81310 59310
rect 81440 59300 81560 59310
rect 81690 59300 81810 59310
rect 81940 59300 82060 59310
rect 82190 59300 82310 59310
rect 82440 59300 82560 59310
rect 82690 59300 82810 59310
rect 82940 59300 83060 59310
rect 83190 59300 83310 59310
rect 83440 59300 83560 59310
rect 83690 59300 83810 59310
rect 83940 59300 84060 59310
rect 84190 59300 84310 59310
rect 84440 59300 84560 59310
rect 84690 59300 84810 59310
rect 84940 59300 85060 59310
rect 85190 59300 85310 59310
rect 85440 59300 85560 59310
rect 85690 59300 85810 59310
rect 85940 59300 86060 59310
rect 86190 59300 86310 59310
rect 86440 59300 86560 59310
rect 86690 59300 86810 59310
rect 86940 59300 87060 59310
rect 87190 59300 87310 59310
rect 87440 59300 87560 59310
rect 87690 59300 87810 59310
rect 87940 59300 88060 59310
rect 88190 59300 88310 59310
rect 88440 59300 88560 59310
rect 88690 59300 88810 59310
rect 88940 59300 89060 59310
rect 89190 59300 89310 59310
rect 89440 59300 89560 59310
rect 89690 59300 89810 59310
rect 89940 59300 90060 59310
rect 90190 59300 90310 59310
rect 90440 59300 90560 59310
rect 90690 59300 90810 59310
rect 90940 59300 91060 59310
rect 91190 59300 91310 59310
rect 91440 59300 91560 59310
rect 91690 59300 91810 59310
rect 91940 59300 92000 59310
rect 81000 59200 92000 59300
rect 81000 59190 81060 59200
rect 81190 59190 81310 59200
rect 81440 59190 81560 59200
rect 81690 59190 81810 59200
rect 81940 59190 82060 59200
rect 82190 59190 82310 59200
rect 82440 59190 82560 59200
rect 82690 59190 82810 59200
rect 82940 59190 83060 59200
rect 83190 59190 83310 59200
rect 83440 59190 83560 59200
rect 83690 59190 83810 59200
rect 83940 59190 84060 59200
rect 84190 59190 84310 59200
rect 84440 59190 84560 59200
rect 84690 59190 84810 59200
rect 84940 59190 85060 59200
rect 85190 59190 85310 59200
rect 85440 59190 85560 59200
rect 85690 59190 85810 59200
rect 85940 59190 86060 59200
rect 86190 59190 86310 59200
rect 86440 59190 86560 59200
rect 86690 59190 86810 59200
rect 86940 59190 87060 59200
rect 87190 59190 87310 59200
rect 87440 59190 87560 59200
rect 87690 59190 87810 59200
rect 87940 59190 88060 59200
rect 88190 59190 88310 59200
rect 88440 59190 88560 59200
rect 88690 59190 88810 59200
rect 88940 59190 89060 59200
rect 89190 59190 89310 59200
rect 89440 59190 89560 59200
rect 89690 59190 89810 59200
rect 89940 59190 90060 59200
rect 90190 59190 90310 59200
rect 90440 59190 90560 59200
rect 90690 59190 90810 59200
rect 90940 59190 91060 59200
rect 91190 59190 91310 59200
rect 91440 59190 91560 59200
rect 91690 59190 91810 59200
rect 91940 59190 92000 59200
rect 81000 59060 81050 59190
rect 81200 59060 81300 59190
rect 81450 59060 81550 59190
rect 81700 59060 81800 59190
rect 81950 59060 82050 59190
rect 82200 59060 82300 59190
rect 82450 59060 82550 59190
rect 82700 59060 82800 59190
rect 82950 59060 83050 59190
rect 83200 59060 83300 59190
rect 83450 59060 83550 59190
rect 83700 59060 83800 59190
rect 83950 59060 84050 59190
rect 84200 59060 84300 59190
rect 84450 59060 84550 59190
rect 84700 59060 84800 59190
rect 84950 59060 85050 59190
rect 85200 59060 85300 59190
rect 85450 59060 85550 59190
rect 85700 59060 85800 59190
rect 85950 59060 86050 59190
rect 86200 59060 86300 59190
rect 86450 59060 86550 59190
rect 86700 59060 86800 59190
rect 86950 59060 87050 59190
rect 87200 59060 87300 59190
rect 87450 59060 87550 59190
rect 87700 59060 87800 59190
rect 87950 59060 88050 59190
rect 88200 59060 88300 59190
rect 88450 59060 88550 59190
rect 88700 59060 88800 59190
rect 88950 59060 89050 59190
rect 89200 59060 89300 59190
rect 89450 59060 89550 59190
rect 89700 59060 89800 59190
rect 89950 59060 90050 59190
rect 90200 59060 90300 59190
rect 90450 59060 90550 59190
rect 90700 59060 90800 59190
rect 90950 59060 91050 59190
rect 91200 59060 91300 59190
rect 91450 59060 91550 59190
rect 91700 59060 91800 59190
rect 91950 59060 92000 59190
rect 81000 59050 81060 59060
rect 81190 59050 81310 59060
rect 81440 59050 81560 59060
rect 81690 59050 81810 59060
rect 81940 59050 82060 59060
rect 82190 59050 82310 59060
rect 82440 59050 82560 59060
rect 82690 59050 82810 59060
rect 82940 59050 83060 59060
rect 83190 59050 83310 59060
rect 83440 59050 83560 59060
rect 83690 59050 83810 59060
rect 83940 59050 84060 59060
rect 84190 59050 84310 59060
rect 84440 59050 84560 59060
rect 84690 59050 84810 59060
rect 84940 59050 85060 59060
rect 85190 59050 85310 59060
rect 85440 59050 85560 59060
rect 85690 59050 85810 59060
rect 85940 59050 86060 59060
rect 86190 59050 86310 59060
rect 86440 59050 86560 59060
rect 86690 59050 86810 59060
rect 86940 59050 87060 59060
rect 87190 59050 87310 59060
rect 87440 59050 87560 59060
rect 87690 59050 87810 59060
rect 87940 59050 88060 59060
rect 88190 59050 88310 59060
rect 88440 59050 88560 59060
rect 88690 59050 88810 59060
rect 88940 59050 89060 59060
rect 89190 59050 89310 59060
rect 89440 59050 89560 59060
rect 89690 59050 89810 59060
rect 89940 59050 90060 59060
rect 90190 59050 90310 59060
rect 90440 59050 90560 59060
rect 90690 59050 90810 59060
rect 90940 59050 91060 59060
rect 91190 59050 91310 59060
rect 91440 59050 91560 59060
rect 91690 59050 91810 59060
rect 91940 59050 92000 59060
rect 81000 58950 92000 59050
rect 81000 58940 81060 58950
rect 81190 58940 81310 58950
rect 81440 58940 81560 58950
rect 81690 58940 81810 58950
rect 81940 58940 82060 58950
rect 82190 58940 82310 58950
rect 82440 58940 82560 58950
rect 82690 58940 82810 58950
rect 82940 58940 83060 58950
rect 83190 58940 83310 58950
rect 83440 58940 83560 58950
rect 83690 58940 83810 58950
rect 83940 58940 84060 58950
rect 84190 58940 84310 58950
rect 84440 58940 84560 58950
rect 84690 58940 84810 58950
rect 84940 58940 85060 58950
rect 85190 58940 85310 58950
rect 85440 58940 85560 58950
rect 85690 58940 85810 58950
rect 85940 58940 86060 58950
rect 86190 58940 86310 58950
rect 86440 58940 86560 58950
rect 86690 58940 86810 58950
rect 86940 58940 87060 58950
rect 87190 58940 87310 58950
rect 87440 58940 87560 58950
rect 87690 58940 87810 58950
rect 87940 58940 88060 58950
rect 88190 58940 88310 58950
rect 88440 58940 88560 58950
rect 88690 58940 88810 58950
rect 88940 58940 89060 58950
rect 89190 58940 89310 58950
rect 89440 58940 89560 58950
rect 89690 58940 89810 58950
rect 89940 58940 90060 58950
rect 90190 58940 90310 58950
rect 90440 58940 90560 58950
rect 90690 58940 90810 58950
rect 90940 58940 91060 58950
rect 91190 58940 91310 58950
rect 91440 58940 91560 58950
rect 91690 58940 91810 58950
rect 91940 58940 92000 58950
rect 81000 58810 81050 58940
rect 81200 58810 81300 58940
rect 81450 58810 81550 58940
rect 81700 58810 81800 58940
rect 81950 58810 82050 58940
rect 82200 58810 82300 58940
rect 82450 58810 82550 58940
rect 82700 58810 82800 58940
rect 82950 58810 83050 58940
rect 83200 58810 83300 58940
rect 83450 58810 83550 58940
rect 83700 58810 83800 58940
rect 83950 58810 84050 58940
rect 84200 58810 84300 58940
rect 84450 58810 84550 58940
rect 84700 58810 84800 58940
rect 84950 58810 85050 58940
rect 85200 58810 85300 58940
rect 85450 58810 85550 58940
rect 85700 58810 85800 58940
rect 85950 58810 86050 58940
rect 86200 58810 86300 58940
rect 86450 58810 86550 58940
rect 86700 58810 86800 58940
rect 86950 58810 87050 58940
rect 87200 58810 87300 58940
rect 87450 58810 87550 58940
rect 87700 58810 87800 58940
rect 87950 58810 88050 58940
rect 88200 58810 88300 58940
rect 88450 58810 88550 58940
rect 88700 58810 88800 58940
rect 88950 58810 89050 58940
rect 89200 58810 89300 58940
rect 89450 58810 89550 58940
rect 89700 58810 89800 58940
rect 89950 58810 90050 58940
rect 90200 58810 90300 58940
rect 90450 58810 90550 58940
rect 90700 58810 90800 58940
rect 90950 58810 91050 58940
rect 91200 58810 91300 58940
rect 91450 58810 91550 58940
rect 91700 58810 91800 58940
rect 91950 58810 92000 58940
rect 81000 58800 81060 58810
rect 81190 58800 81310 58810
rect 81440 58800 81560 58810
rect 81690 58800 81810 58810
rect 81940 58800 82060 58810
rect 82190 58800 82310 58810
rect 82440 58800 82560 58810
rect 82690 58800 82810 58810
rect 82940 58800 83060 58810
rect 83190 58800 83310 58810
rect 83440 58800 83560 58810
rect 83690 58800 83810 58810
rect 83940 58800 84060 58810
rect 84190 58800 84310 58810
rect 84440 58800 84560 58810
rect 84690 58800 84810 58810
rect 84940 58800 85060 58810
rect 85190 58800 85310 58810
rect 85440 58800 85560 58810
rect 85690 58800 85810 58810
rect 85940 58800 86060 58810
rect 86190 58800 86310 58810
rect 86440 58800 86560 58810
rect 86690 58800 86810 58810
rect 86940 58800 87060 58810
rect 87190 58800 87310 58810
rect 87440 58800 87560 58810
rect 87690 58800 87810 58810
rect 87940 58800 88060 58810
rect 88190 58800 88310 58810
rect 88440 58800 88560 58810
rect 88690 58800 88810 58810
rect 88940 58800 89060 58810
rect 89190 58800 89310 58810
rect 89440 58800 89560 58810
rect 89690 58800 89810 58810
rect 89940 58800 90060 58810
rect 90190 58800 90310 58810
rect 90440 58800 90560 58810
rect 90690 58800 90810 58810
rect 90940 58800 91060 58810
rect 91190 58800 91310 58810
rect 91440 58800 91560 58810
rect 91690 58800 91810 58810
rect 91940 58800 92000 58810
rect 81000 58700 92000 58800
rect 81000 58690 81060 58700
rect 81190 58690 81310 58700
rect 81440 58690 81560 58700
rect 81690 58690 81810 58700
rect 81940 58690 82060 58700
rect 82190 58690 82310 58700
rect 82440 58690 82560 58700
rect 82690 58690 82810 58700
rect 82940 58690 83060 58700
rect 83190 58690 83310 58700
rect 83440 58690 83560 58700
rect 83690 58690 83810 58700
rect 83940 58690 84060 58700
rect 84190 58690 84310 58700
rect 84440 58690 84560 58700
rect 84690 58690 84810 58700
rect 84940 58690 85060 58700
rect 85190 58690 85310 58700
rect 85440 58690 85560 58700
rect 85690 58690 85810 58700
rect 85940 58690 86060 58700
rect 86190 58690 86310 58700
rect 86440 58690 86560 58700
rect 86690 58690 86810 58700
rect 86940 58690 87060 58700
rect 87190 58690 87310 58700
rect 87440 58690 87560 58700
rect 87690 58690 87810 58700
rect 87940 58690 88060 58700
rect 88190 58690 88310 58700
rect 88440 58690 88560 58700
rect 88690 58690 88810 58700
rect 88940 58690 89060 58700
rect 89190 58690 89310 58700
rect 89440 58690 89560 58700
rect 89690 58690 89810 58700
rect 89940 58690 90060 58700
rect 90190 58690 90310 58700
rect 90440 58690 90560 58700
rect 90690 58690 90810 58700
rect 90940 58690 91060 58700
rect 91190 58690 91310 58700
rect 91440 58690 91560 58700
rect 91690 58690 91810 58700
rect 91940 58690 92000 58700
rect 81000 58560 81050 58690
rect 81200 58560 81300 58690
rect 81450 58560 81550 58690
rect 81700 58560 81800 58690
rect 81950 58560 82050 58690
rect 82200 58560 82300 58690
rect 82450 58560 82550 58690
rect 82700 58560 82800 58690
rect 82950 58560 83050 58690
rect 83200 58560 83300 58690
rect 83450 58560 83550 58690
rect 83700 58560 83800 58690
rect 83950 58560 84050 58690
rect 84200 58560 84300 58690
rect 84450 58560 84550 58690
rect 84700 58560 84800 58690
rect 84950 58560 85050 58690
rect 85200 58560 85300 58690
rect 85450 58560 85550 58690
rect 85700 58560 85800 58690
rect 85950 58560 86050 58690
rect 86200 58560 86300 58690
rect 86450 58560 86550 58690
rect 86700 58560 86800 58690
rect 86950 58560 87050 58690
rect 87200 58560 87300 58690
rect 87450 58560 87550 58690
rect 87700 58560 87800 58690
rect 87950 58560 88050 58690
rect 88200 58560 88300 58690
rect 88450 58560 88550 58690
rect 88700 58560 88800 58690
rect 88950 58560 89050 58690
rect 89200 58560 89300 58690
rect 89450 58560 89550 58690
rect 89700 58560 89800 58690
rect 89950 58560 90050 58690
rect 90200 58560 90300 58690
rect 90450 58560 90550 58690
rect 90700 58560 90800 58690
rect 90950 58560 91050 58690
rect 91200 58560 91300 58690
rect 91450 58560 91550 58690
rect 91700 58560 91800 58690
rect 91950 58560 92000 58690
rect 81000 58550 81060 58560
rect 81190 58550 81310 58560
rect 81440 58550 81560 58560
rect 81690 58550 81810 58560
rect 81940 58550 82060 58560
rect 82190 58550 82310 58560
rect 82440 58550 82560 58560
rect 82690 58550 82810 58560
rect 82940 58550 83060 58560
rect 83190 58550 83310 58560
rect 83440 58550 83560 58560
rect 83690 58550 83810 58560
rect 83940 58550 84060 58560
rect 84190 58550 84310 58560
rect 84440 58550 84560 58560
rect 84690 58550 84810 58560
rect 84940 58550 85060 58560
rect 85190 58550 85310 58560
rect 85440 58550 85560 58560
rect 85690 58550 85810 58560
rect 85940 58550 86060 58560
rect 86190 58550 86310 58560
rect 86440 58550 86560 58560
rect 86690 58550 86810 58560
rect 86940 58550 87060 58560
rect 87190 58550 87310 58560
rect 87440 58550 87560 58560
rect 87690 58550 87810 58560
rect 87940 58550 88060 58560
rect 88190 58550 88310 58560
rect 88440 58550 88560 58560
rect 88690 58550 88810 58560
rect 88940 58550 89060 58560
rect 89190 58550 89310 58560
rect 89440 58550 89560 58560
rect 89690 58550 89810 58560
rect 89940 58550 90060 58560
rect 90190 58550 90310 58560
rect 90440 58550 90560 58560
rect 90690 58550 90810 58560
rect 90940 58550 91060 58560
rect 91190 58550 91310 58560
rect 91440 58550 91560 58560
rect 91690 58550 91810 58560
rect 91940 58550 92000 58560
rect 81000 58450 92000 58550
rect 81000 58440 81060 58450
rect 81190 58440 81310 58450
rect 81440 58440 81560 58450
rect 81690 58440 81810 58450
rect 81940 58440 82060 58450
rect 82190 58440 82310 58450
rect 82440 58440 82560 58450
rect 82690 58440 82810 58450
rect 82940 58440 83060 58450
rect 83190 58440 83310 58450
rect 83440 58440 83560 58450
rect 83690 58440 83810 58450
rect 83940 58440 84060 58450
rect 84190 58440 84310 58450
rect 84440 58440 84560 58450
rect 84690 58440 84810 58450
rect 84940 58440 85060 58450
rect 85190 58440 85310 58450
rect 85440 58440 85560 58450
rect 85690 58440 85810 58450
rect 85940 58440 86060 58450
rect 86190 58440 86310 58450
rect 86440 58440 86560 58450
rect 86690 58440 86810 58450
rect 86940 58440 87060 58450
rect 87190 58440 87310 58450
rect 87440 58440 87560 58450
rect 87690 58440 87810 58450
rect 87940 58440 88060 58450
rect 88190 58440 88310 58450
rect 88440 58440 88560 58450
rect 88690 58440 88810 58450
rect 88940 58440 89060 58450
rect 89190 58440 89310 58450
rect 89440 58440 89560 58450
rect 89690 58440 89810 58450
rect 89940 58440 90060 58450
rect 90190 58440 90310 58450
rect 90440 58440 90560 58450
rect 90690 58440 90810 58450
rect 90940 58440 91060 58450
rect 91190 58440 91310 58450
rect 91440 58440 91560 58450
rect 91690 58440 91810 58450
rect 91940 58440 92000 58450
rect 81000 58310 81050 58440
rect 81200 58310 81300 58440
rect 81450 58310 81550 58440
rect 81700 58310 81800 58440
rect 81950 58310 82050 58440
rect 82200 58310 82300 58440
rect 82450 58310 82550 58440
rect 82700 58310 82800 58440
rect 82950 58310 83050 58440
rect 83200 58310 83300 58440
rect 83450 58310 83550 58440
rect 83700 58310 83800 58440
rect 83950 58310 84050 58440
rect 84200 58310 84300 58440
rect 84450 58310 84550 58440
rect 84700 58310 84800 58440
rect 84950 58310 85050 58440
rect 85200 58310 85300 58440
rect 85450 58310 85550 58440
rect 85700 58310 85800 58440
rect 85950 58310 86050 58440
rect 86200 58310 86300 58440
rect 86450 58310 86550 58440
rect 86700 58310 86800 58440
rect 86950 58310 87050 58440
rect 87200 58310 87300 58440
rect 87450 58310 87550 58440
rect 87700 58310 87800 58440
rect 87950 58310 88050 58440
rect 88200 58310 88300 58440
rect 88450 58310 88550 58440
rect 88700 58310 88800 58440
rect 88950 58310 89050 58440
rect 89200 58310 89300 58440
rect 89450 58310 89550 58440
rect 89700 58310 89800 58440
rect 89950 58310 90050 58440
rect 90200 58310 90300 58440
rect 90450 58310 90550 58440
rect 90700 58310 90800 58440
rect 90950 58310 91050 58440
rect 91200 58310 91300 58440
rect 91450 58310 91550 58440
rect 91700 58310 91800 58440
rect 91950 58310 92000 58440
rect 81000 58300 81060 58310
rect 81190 58300 81310 58310
rect 81440 58300 81560 58310
rect 81690 58300 81810 58310
rect 81940 58300 82060 58310
rect 82190 58300 82310 58310
rect 82440 58300 82560 58310
rect 82690 58300 82810 58310
rect 82940 58300 83060 58310
rect 83190 58300 83310 58310
rect 83440 58300 83560 58310
rect 83690 58300 83810 58310
rect 83940 58300 84060 58310
rect 84190 58300 84310 58310
rect 84440 58300 84560 58310
rect 84690 58300 84810 58310
rect 84940 58300 85060 58310
rect 85190 58300 85310 58310
rect 85440 58300 85560 58310
rect 85690 58300 85810 58310
rect 85940 58300 86060 58310
rect 86190 58300 86310 58310
rect 86440 58300 86560 58310
rect 86690 58300 86810 58310
rect 86940 58300 87060 58310
rect 87190 58300 87310 58310
rect 87440 58300 87560 58310
rect 87690 58300 87810 58310
rect 87940 58300 88060 58310
rect 88190 58300 88310 58310
rect 88440 58300 88560 58310
rect 88690 58300 88810 58310
rect 88940 58300 89060 58310
rect 89190 58300 89310 58310
rect 89440 58300 89560 58310
rect 89690 58300 89810 58310
rect 89940 58300 90060 58310
rect 90190 58300 90310 58310
rect 90440 58300 90560 58310
rect 90690 58300 90810 58310
rect 90940 58300 91060 58310
rect 91190 58300 91310 58310
rect 91440 58300 91560 58310
rect 91690 58300 91810 58310
rect 91940 58300 92000 58310
rect 81000 58200 92000 58300
rect 81000 58190 81060 58200
rect 81190 58190 81310 58200
rect 81440 58190 81560 58200
rect 81690 58190 81810 58200
rect 81940 58190 82060 58200
rect 82190 58190 82310 58200
rect 82440 58190 82560 58200
rect 82690 58190 82810 58200
rect 82940 58190 83060 58200
rect 83190 58190 83310 58200
rect 83440 58190 83560 58200
rect 83690 58190 83810 58200
rect 83940 58190 84060 58200
rect 84190 58190 84310 58200
rect 84440 58190 84560 58200
rect 84690 58190 84810 58200
rect 84940 58190 85060 58200
rect 85190 58190 85310 58200
rect 85440 58190 85560 58200
rect 85690 58190 85810 58200
rect 85940 58190 86060 58200
rect 86190 58190 86310 58200
rect 86440 58190 86560 58200
rect 86690 58190 86810 58200
rect 86940 58190 87060 58200
rect 87190 58190 87310 58200
rect 87440 58190 87560 58200
rect 87690 58190 87810 58200
rect 87940 58190 88060 58200
rect 88190 58190 88310 58200
rect 88440 58190 88560 58200
rect 88690 58190 88810 58200
rect 88940 58190 89060 58200
rect 89190 58190 89310 58200
rect 89440 58190 89560 58200
rect 89690 58190 89810 58200
rect 89940 58190 90060 58200
rect 90190 58190 90310 58200
rect 90440 58190 90560 58200
rect 90690 58190 90810 58200
rect 90940 58190 91060 58200
rect 91190 58190 91310 58200
rect 91440 58190 91560 58200
rect 91690 58190 91810 58200
rect 91940 58190 92000 58200
rect 81000 58060 81050 58190
rect 81200 58060 81300 58190
rect 81450 58060 81550 58190
rect 81700 58060 81800 58190
rect 81950 58060 82050 58190
rect 82200 58060 82300 58190
rect 82450 58060 82550 58190
rect 82700 58060 82800 58190
rect 82950 58060 83050 58190
rect 83200 58060 83300 58190
rect 83450 58060 83550 58190
rect 83700 58060 83800 58190
rect 83950 58060 84050 58190
rect 84200 58060 84300 58190
rect 84450 58060 84550 58190
rect 84700 58060 84800 58190
rect 84950 58060 85050 58190
rect 85200 58060 85300 58190
rect 85450 58060 85550 58190
rect 85700 58060 85800 58190
rect 85950 58060 86050 58190
rect 86200 58060 86300 58190
rect 86450 58060 86550 58190
rect 86700 58060 86800 58190
rect 86950 58060 87050 58190
rect 87200 58060 87300 58190
rect 87450 58060 87550 58190
rect 87700 58060 87800 58190
rect 87950 58060 88050 58190
rect 88200 58060 88300 58190
rect 88450 58060 88550 58190
rect 88700 58060 88800 58190
rect 88950 58060 89050 58190
rect 89200 58060 89300 58190
rect 89450 58060 89550 58190
rect 89700 58060 89800 58190
rect 89950 58060 90050 58190
rect 90200 58060 90300 58190
rect 90450 58060 90550 58190
rect 90700 58060 90800 58190
rect 90950 58060 91050 58190
rect 91200 58060 91300 58190
rect 91450 58060 91550 58190
rect 91700 58060 91800 58190
rect 91950 58060 92000 58190
rect 81000 58050 81060 58060
rect 81190 58050 81310 58060
rect 81440 58050 81560 58060
rect 81690 58050 81810 58060
rect 81940 58050 82060 58060
rect 82190 58050 82310 58060
rect 82440 58050 82560 58060
rect 82690 58050 82810 58060
rect 82940 58050 83060 58060
rect 83190 58050 83310 58060
rect 83440 58050 83560 58060
rect 83690 58050 83810 58060
rect 83940 58050 84060 58060
rect 84190 58050 84310 58060
rect 84440 58050 84560 58060
rect 84690 58050 84810 58060
rect 84940 58050 85060 58060
rect 85190 58050 85310 58060
rect 85440 58050 85560 58060
rect 85690 58050 85810 58060
rect 85940 58050 86060 58060
rect 86190 58050 86310 58060
rect 86440 58050 86560 58060
rect 86690 58050 86810 58060
rect 86940 58050 87060 58060
rect 87190 58050 87310 58060
rect 87440 58050 87560 58060
rect 87690 58050 87810 58060
rect 87940 58050 88060 58060
rect 88190 58050 88310 58060
rect 88440 58050 88560 58060
rect 88690 58050 88810 58060
rect 88940 58050 89060 58060
rect 89190 58050 89310 58060
rect 89440 58050 89560 58060
rect 89690 58050 89810 58060
rect 89940 58050 90060 58060
rect 90190 58050 90310 58060
rect 90440 58050 90560 58060
rect 90690 58050 90810 58060
rect 90940 58050 91060 58060
rect 91190 58050 91310 58060
rect 91440 58050 91560 58060
rect 91690 58050 91810 58060
rect 91940 58050 92000 58060
rect 81000 57950 92000 58050
rect 81000 57940 81060 57950
rect 81190 57940 81310 57950
rect 81440 57940 81560 57950
rect 81690 57940 81810 57950
rect 81940 57940 82060 57950
rect 82190 57940 82310 57950
rect 82440 57940 82560 57950
rect 82690 57940 82810 57950
rect 82940 57940 83060 57950
rect 83190 57940 83310 57950
rect 83440 57940 83560 57950
rect 83690 57940 83810 57950
rect 83940 57940 84060 57950
rect 84190 57940 84310 57950
rect 84440 57940 84560 57950
rect 84690 57940 84810 57950
rect 84940 57940 85060 57950
rect 85190 57940 85310 57950
rect 85440 57940 85560 57950
rect 85690 57940 85810 57950
rect 85940 57940 86060 57950
rect 86190 57940 86310 57950
rect 86440 57940 86560 57950
rect 86690 57940 86810 57950
rect 86940 57940 87060 57950
rect 87190 57940 87310 57950
rect 87440 57940 87560 57950
rect 87690 57940 87810 57950
rect 87940 57940 88060 57950
rect 88190 57940 88310 57950
rect 88440 57940 88560 57950
rect 88690 57940 88810 57950
rect 88940 57940 89060 57950
rect 89190 57940 89310 57950
rect 89440 57940 89560 57950
rect 89690 57940 89810 57950
rect 89940 57940 90060 57950
rect 90190 57940 90310 57950
rect 90440 57940 90560 57950
rect 90690 57940 90810 57950
rect 90940 57940 91060 57950
rect 91190 57940 91310 57950
rect 91440 57940 91560 57950
rect 91690 57940 91810 57950
rect 91940 57940 92000 57950
rect 81000 57810 81050 57940
rect 81200 57810 81300 57940
rect 81450 57810 81550 57940
rect 81700 57810 81800 57940
rect 81950 57810 82050 57940
rect 82200 57810 82300 57940
rect 82450 57810 82550 57940
rect 82700 57810 82800 57940
rect 82950 57810 83050 57940
rect 83200 57810 83300 57940
rect 83450 57810 83550 57940
rect 83700 57810 83800 57940
rect 83950 57810 84050 57940
rect 84200 57810 84300 57940
rect 84450 57810 84550 57940
rect 84700 57810 84800 57940
rect 84950 57810 85050 57940
rect 85200 57810 85300 57940
rect 85450 57810 85550 57940
rect 85700 57810 85800 57940
rect 85950 57810 86050 57940
rect 86200 57810 86300 57940
rect 86450 57810 86550 57940
rect 86700 57810 86800 57940
rect 86950 57810 87050 57940
rect 87200 57810 87300 57940
rect 87450 57810 87550 57940
rect 87700 57810 87800 57940
rect 87950 57810 88050 57940
rect 88200 57810 88300 57940
rect 88450 57810 88550 57940
rect 88700 57810 88800 57940
rect 88950 57810 89050 57940
rect 89200 57810 89300 57940
rect 89450 57810 89550 57940
rect 89700 57810 89800 57940
rect 89950 57810 90050 57940
rect 90200 57810 90300 57940
rect 90450 57810 90550 57940
rect 90700 57810 90800 57940
rect 90950 57810 91050 57940
rect 91200 57810 91300 57940
rect 91450 57810 91550 57940
rect 91700 57810 91800 57940
rect 91950 57810 92000 57940
rect 81000 57800 81060 57810
rect 81190 57800 81310 57810
rect 81440 57800 81560 57810
rect 81690 57800 81810 57810
rect 81940 57800 82060 57810
rect 82190 57800 82310 57810
rect 82440 57800 82560 57810
rect 82690 57800 82810 57810
rect 82940 57800 83060 57810
rect 83190 57800 83310 57810
rect 83440 57800 83560 57810
rect 83690 57800 83810 57810
rect 83940 57800 84060 57810
rect 84190 57800 84310 57810
rect 84440 57800 84560 57810
rect 84690 57800 84810 57810
rect 84940 57800 85060 57810
rect 85190 57800 85310 57810
rect 85440 57800 85560 57810
rect 85690 57800 85810 57810
rect 85940 57800 86060 57810
rect 86190 57800 86310 57810
rect 86440 57800 86560 57810
rect 86690 57800 86810 57810
rect 86940 57800 87060 57810
rect 87190 57800 87310 57810
rect 87440 57800 87560 57810
rect 87690 57800 87810 57810
rect 87940 57800 88060 57810
rect 88190 57800 88310 57810
rect 88440 57800 88560 57810
rect 88690 57800 88810 57810
rect 88940 57800 89060 57810
rect 89190 57800 89310 57810
rect 89440 57800 89560 57810
rect 89690 57800 89810 57810
rect 89940 57800 90060 57810
rect 90190 57800 90310 57810
rect 90440 57800 90560 57810
rect 90690 57800 90810 57810
rect 90940 57800 91060 57810
rect 91190 57800 91310 57810
rect 91440 57800 91560 57810
rect 91690 57800 91810 57810
rect 91940 57800 92000 57810
rect 81000 57700 92000 57800
rect 81000 57690 81060 57700
rect 81190 57690 81310 57700
rect 81440 57690 81560 57700
rect 81690 57690 81810 57700
rect 81940 57690 82060 57700
rect 82190 57690 82310 57700
rect 82440 57690 82560 57700
rect 82690 57690 82810 57700
rect 82940 57690 83060 57700
rect 83190 57690 83310 57700
rect 83440 57690 83560 57700
rect 83690 57690 83810 57700
rect 83940 57690 84060 57700
rect 84190 57690 84310 57700
rect 84440 57690 84560 57700
rect 84690 57690 84810 57700
rect 84940 57690 85060 57700
rect 85190 57690 85310 57700
rect 85440 57690 85560 57700
rect 85690 57690 85810 57700
rect 85940 57690 86060 57700
rect 86190 57690 86310 57700
rect 86440 57690 86560 57700
rect 86690 57690 86810 57700
rect 86940 57690 87060 57700
rect 87190 57690 87310 57700
rect 87440 57690 87560 57700
rect 87690 57690 87810 57700
rect 87940 57690 88060 57700
rect 88190 57690 88310 57700
rect 88440 57690 88560 57700
rect 88690 57690 88810 57700
rect 88940 57690 89060 57700
rect 89190 57690 89310 57700
rect 89440 57690 89560 57700
rect 89690 57690 89810 57700
rect 89940 57690 90060 57700
rect 90190 57690 90310 57700
rect 90440 57690 90560 57700
rect 90690 57690 90810 57700
rect 90940 57690 91060 57700
rect 91190 57690 91310 57700
rect 91440 57690 91560 57700
rect 91690 57690 91810 57700
rect 91940 57690 92000 57700
rect 81000 57560 81050 57690
rect 81200 57560 81300 57690
rect 81450 57560 81550 57690
rect 81700 57560 81800 57690
rect 81950 57560 82050 57690
rect 82200 57560 82300 57690
rect 82450 57560 82550 57690
rect 82700 57560 82800 57690
rect 82950 57560 83050 57690
rect 83200 57560 83300 57690
rect 83450 57560 83550 57690
rect 83700 57560 83800 57690
rect 83950 57560 84050 57690
rect 84200 57560 84300 57690
rect 84450 57560 84550 57690
rect 84700 57560 84800 57690
rect 84950 57560 85050 57690
rect 85200 57560 85300 57690
rect 85450 57560 85550 57690
rect 85700 57560 85800 57690
rect 85950 57560 86050 57690
rect 86200 57560 86300 57690
rect 86450 57560 86550 57690
rect 86700 57560 86800 57690
rect 86950 57560 87050 57690
rect 87200 57560 87300 57690
rect 87450 57560 87550 57690
rect 87700 57560 87800 57690
rect 87950 57560 88050 57690
rect 88200 57560 88300 57690
rect 88450 57560 88550 57690
rect 88700 57560 88800 57690
rect 88950 57560 89050 57690
rect 89200 57560 89300 57690
rect 89450 57560 89550 57690
rect 89700 57560 89800 57690
rect 89950 57560 90050 57690
rect 90200 57560 90300 57690
rect 90450 57560 90550 57690
rect 90700 57560 90800 57690
rect 90950 57560 91050 57690
rect 91200 57560 91300 57690
rect 91450 57560 91550 57690
rect 91700 57560 91800 57690
rect 91950 57560 92000 57690
rect 81000 57550 81060 57560
rect 81190 57550 81310 57560
rect 81440 57550 81560 57560
rect 81690 57550 81810 57560
rect 81940 57550 82060 57560
rect 82190 57550 82310 57560
rect 82440 57550 82560 57560
rect 82690 57550 82810 57560
rect 82940 57550 83060 57560
rect 83190 57550 83310 57560
rect 83440 57550 83560 57560
rect 83690 57550 83810 57560
rect 83940 57550 84060 57560
rect 84190 57550 84310 57560
rect 84440 57550 84560 57560
rect 84690 57550 84810 57560
rect 84940 57550 85060 57560
rect 85190 57550 85310 57560
rect 85440 57550 85560 57560
rect 85690 57550 85810 57560
rect 85940 57550 86060 57560
rect 86190 57550 86310 57560
rect 86440 57550 86560 57560
rect 86690 57550 86810 57560
rect 86940 57550 87060 57560
rect 87190 57550 87310 57560
rect 87440 57550 87560 57560
rect 87690 57550 87810 57560
rect 87940 57550 88060 57560
rect 88190 57550 88310 57560
rect 88440 57550 88560 57560
rect 88690 57550 88810 57560
rect 88940 57550 89060 57560
rect 89190 57550 89310 57560
rect 89440 57550 89560 57560
rect 89690 57550 89810 57560
rect 89940 57550 90060 57560
rect 90190 57550 90310 57560
rect 90440 57550 90560 57560
rect 90690 57550 90810 57560
rect 90940 57550 91060 57560
rect 91190 57550 91310 57560
rect 91440 57550 91560 57560
rect 91690 57550 91810 57560
rect 91940 57550 92000 57560
rect 81000 57450 92000 57550
rect 81000 57440 81060 57450
rect 81190 57440 81310 57450
rect 81440 57440 81560 57450
rect 81690 57440 81810 57450
rect 81940 57440 82060 57450
rect 82190 57440 82310 57450
rect 82440 57440 82560 57450
rect 82690 57440 82810 57450
rect 82940 57440 83060 57450
rect 83190 57440 83310 57450
rect 83440 57440 83560 57450
rect 83690 57440 83810 57450
rect 83940 57440 84060 57450
rect 84190 57440 84310 57450
rect 84440 57440 84560 57450
rect 84690 57440 84810 57450
rect 84940 57440 85060 57450
rect 85190 57440 85310 57450
rect 85440 57440 85560 57450
rect 85690 57440 85810 57450
rect 85940 57440 86060 57450
rect 86190 57440 86310 57450
rect 86440 57440 86560 57450
rect 86690 57440 86810 57450
rect 86940 57440 87060 57450
rect 87190 57440 87310 57450
rect 87440 57440 87560 57450
rect 87690 57440 87810 57450
rect 87940 57440 88060 57450
rect 88190 57440 88310 57450
rect 88440 57440 88560 57450
rect 88690 57440 88810 57450
rect 88940 57440 89060 57450
rect 89190 57440 89310 57450
rect 89440 57440 89560 57450
rect 89690 57440 89810 57450
rect 89940 57440 90060 57450
rect 90190 57440 90310 57450
rect 90440 57440 90560 57450
rect 90690 57440 90810 57450
rect 90940 57440 91060 57450
rect 91190 57440 91310 57450
rect 91440 57440 91560 57450
rect 91690 57440 91810 57450
rect 91940 57440 92000 57450
rect 81000 57310 81050 57440
rect 81200 57310 81300 57440
rect 81450 57310 81550 57440
rect 81700 57310 81800 57440
rect 81950 57310 82050 57440
rect 82200 57310 82300 57440
rect 82450 57310 82550 57440
rect 82700 57310 82800 57440
rect 82950 57310 83050 57440
rect 83200 57310 83300 57440
rect 83450 57310 83550 57440
rect 83700 57310 83800 57440
rect 83950 57310 84050 57440
rect 84200 57310 84300 57440
rect 84450 57310 84550 57440
rect 84700 57310 84800 57440
rect 84950 57310 85050 57440
rect 85200 57310 85300 57440
rect 85450 57310 85550 57440
rect 85700 57310 85800 57440
rect 85950 57310 86050 57440
rect 86200 57310 86300 57440
rect 86450 57310 86550 57440
rect 86700 57310 86800 57440
rect 86950 57310 87050 57440
rect 87200 57310 87300 57440
rect 87450 57310 87550 57440
rect 87700 57310 87800 57440
rect 87950 57310 88050 57440
rect 88200 57310 88300 57440
rect 88450 57310 88550 57440
rect 88700 57310 88800 57440
rect 88950 57310 89050 57440
rect 89200 57310 89300 57440
rect 89450 57310 89550 57440
rect 89700 57310 89800 57440
rect 89950 57310 90050 57440
rect 90200 57310 90300 57440
rect 90450 57310 90550 57440
rect 90700 57310 90800 57440
rect 90950 57310 91050 57440
rect 91200 57310 91300 57440
rect 91450 57310 91550 57440
rect 91700 57310 91800 57440
rect 91950 57310 92000 57440
rect 81000 57300 81060 57310
rect 81190 57300 81310 57310
rect 81440 57300 81560 57310
rect 81690 57300 81810 57310
rect 81940 57300 82060 57310
rect 82190 57300 82310 57310
rect 82440 57300 82560 57310
rect 82690 57300 82810 57310
rect 82940 57300 83060 57310
rect 83190 57300 83310 57310
rect 83440 57300 83560 57310
rect 83690 57300 83810 57310
rect 83940 57300 84060 57310
rect 84190 57300 84310 57310
rect 84440 57300 84560 57310
rect 84690 57300 84810 57310
rect 84940 57300 85060 57310
rect 85190 57300 85310 57310
rect 85440 57300 85560 57310
rect 85690 57300 85810 57310
rect 85940 57300 86060 57310
rect 86190 57300 86310 57310
rect 86440 57300 86560 57310
rect 86690 57300 86810 57310
rect 86940 57300 87060 57310
rect 87190 57300 87310 57310
rect 87440 57300 87560 57310
rect 87690 57300 87810 57310
rect 87940 57300 88060 57310
rect 88190 57300 88310 57310
rect 88440 57300 88560 57310
rect 88690 57300 88810 57310
rect 88940 57300 89060 57310
rect 89190 57300 89310 57310
rect 89440 57300 89560 57310
rect 89690 57300 89810 57310
rect 89940 57300 90060 57310
rect 90190 57300 90310 57310
rect 90440 57300 90560 57310
rect 90690 57300 90810 57310
rect 90940 57300 91060 57310
rect 91190 57300 91310 57310
rect 91440 57300 91560 57310
rect 91690 57300 91810 57310
rect 91940 57300 92000 57310
rect 81000 57200 92000 57300
rect 81000 57190 81060 57200
rect 81190 57190 81310 57200
rect 81440 57190 81560 57200
rect 81690 57190 81810 57200
rect 81940 57190 82060 57200
rect 82190 57190 82310 57200
rect 82440 57190 82560 57200
rect 82690 57190 82810 57200
rect 82940 57190 83060 57200
rect 83190 57190 83310 57200
rect 83440 57190 83560 57200
rect 83690 57190 83810 57200
rect 83940 57190 84060 57200
rect 84190 57190 84310 57200
rect 84440 57190 84560 57200
rect 84690 57190 84810 57200
rect 84940 57190 85060 57200
rect 85190 57190 85310 57200
rect 85440 57190 85560 57200
rect 85690 57190 85810 57200
rect 85940 57190 86060 57200
rect 86190 57190 86310 57200
rect 86440 57190 86560 57200
rect 86690 57190 86810 57200
rect 86940 57190 87060 57200
rect 87190 57190 87310 57200
rect 87440 57190 87560 57200
rect 87690 57190 87810 57200
rect 87940 57190 88060 57200
rect 88190 57190 88310 57200
rect 88440 57190 88560 57200
rect 88690 57190 88810 57200
rect 88940 57190 89060 57200
rect 89190 57190 89310 57200
rect 89440 57190 89560 57200
rect 89690 57190 89810 57200
rect 89940 57190 90060 57200
rect 90190 57190 90310 57200
rect 90440 57190 90560 57200
rect 90690 57190 90810 57200
rect 90940 57190 91060 57200
rect 91190 57190 91310 57200
rect 91440 57190 91560 57200
rect 91690 57190 91810 57200
rect 91940 57190 92000 57200
rect 81000 57060 81050 57190
rect 81200 57060 81300 57190
rect 81450 57060 81550 57190
rect 81700 57060 81800 57190
rect 81950 57060 82050 57190
rect 82200 57060 82300 57190
rect 82450 57060 82550 57190
rect 82700 57060 82800 57190
rect 82950 57060 83050 57190
rect 83200 57060 83300 57190
rect 83450 57060 83550 57190
rect 83700 57060 83800 57190
rect 83950 57060 84050 57190
rect 84200 57060 84300 57190
rect 84450 57060 84550 57190
rect 84700 57060 84800 57190
rect 84950 57060 85050 57190
rect 85200 57060 85300 57190
rect 85450 57060 85550 57190
rect 85700 57060 85800 57190
rect 85950 57060 86050 57190
rect 86200 57060 86300 57190
rect 86450 57060 86550 57190
rect 86700 57060 86800 57190
rect 86950 57060 87050 57190
rect 87200 57060 87300 57190
rect 87450 57060 87550 57190
rect 87700 57060 87800 57190
rect 87950 57060 88050 57190
rect 88200 57060 88300 57190
rect 88450 57060 88550 57190
rect 88700 57060 88800 57190
rect 88950 57060 89050 57190
rect 89200 57060 89300 57190
rect 89450 57060 89550 57190
rect 89700 57060 89800 57190
rect 89950 57060 90050 57190
rect 90200 57060 90300 57190
rect 90450 57060 90550 57190
rect 90700 57060 90800 57190
rect 90950 57060 91050 57190
rect 91200 57060 91300 57190
rect 91450 57060 91550 57190
rect 91700 57060 91800 57190
rect 91950 57060 92000 57190
rect 81000 57050 81060 57060
rect 81190 57050 81310 57060
rect 81440 57050 81560 57060
rect 81690 57050 81810 57060
rect 81940 57050 82060 57060
rect 82190 57050 82310 57060
rect 82440 57050 82560 57060
rect 82690 57050 82810 57060
rect 82940 57050 83060 57060
rect 83190 57050 83310 57060
rect 83440 57050 83560 57060
rect 83690 57050 83810 57060
rect 83940 57050 84060 57060
rect 84190 57050 84310 57060
rect 84440 57050 84560 57060
rect 84690 57050 84810 57060
rect 84940 57050 85060 57060
rect 85190 57050 85310 57060
rect 85440 57050 85560 57060
rect 85690 57050 85810 57060
rect 85940 57050 86060 57060
rect 86190 57050 86310 57060
rect 86440 57050 86560 57060
rect 86690 57050 86810 57060
rect 86940 57050 87060 57060
rect 87190 57050 87310 57060
rect 87440 57050 87560 57060
rect 87690 57050 87810 57060
rect 87940 57050 88060 57060
rect 88190 57050 88310 57060
rect 88440 57050 88560 57060
rect 88690 57050 88810 57060
rect 88940 57050 89060 57060
rect 89190 57050 89310 57060
rect 89440 57050 89560 57060
rect 89690 57050 89810 57060
rect 89940 57050 90060 57060
rect 90190 57050 90310 57060
rect 90440 57050 90560 57060
rect 90690 57050 90810 57060
rect 90940 57050 91060 57060
rect 91190 57050 91310 57060
rect 91440 57050 91560 57060
rect 91690 57050 91810 57060
rect 91940 57050 92000 57060
rect 81000 57000 92000 57050
rect 107000 60950 116000 61000
rect 107000 60940 107060 60950
rect 107190 60940 107310 60950
rect 107440 60940 107560 60950
rect 107690 60940 107810 60950
rect 107940 60940 108060 60950
rect 108190 60940 108310 60950
rect 108440 60940 108560 60950
rect 108690 60940 108810 60950
rect 108940 60940 109060 60950
rect 109190 60940 109310 60950
rect 109440 60940 109560 60950
rect 109690 60940 109810 60950
rect 109940 60940 110060 60950
rect 110190 60940 110310 60950
rect 110440 60940 110560 60950
rect 110690 60940 110810 60950
rect 110940 60940 111060 60950
rect 111190 60940 111310 60950
rect 111440 60940 111560 60950
rect 111690 60940 111810 60950
rect 111940 60940 112060 60950
rect 112190 60940 112310 60950
rect 112440 60940 112560 60950
rect 112690 60940 112810 60950
rect 112940 60940 113060 60950
rect 113190 60940 113310 60950
rect 113440 60940 113560 60950
rect 113690 60940 113810 60950
rect 113940 60940 114060 60950
rect 114190 60940 114310 60950
rect 114440 60940 114560 60950
rect 114690 60940 114810 60950
rect 114940 60940 115060 60950
rect 115190 60940 115310 60950
rect 115440 60940 115560 60950
rect 115690 60940 115810 60950
rect 115940 60940 116000 60950
rect 107000 60810 107050 60940
rect 107200 60810 107300 60940
rect 107450 60810 107550 60940
rect 107700 60810 107800 60940
rect 107950 60810 108050 60940
rect 108200 60810 108300 60940
rect 108450 60810 108550 60940
rect 108700 60810 108800 60940
rect 108950 60810 109050 60940
rect 109200 60810 109300 60940
rect 109450 60810 109550 60940
rect 109700 60810 109800 60940
rect 109950 60810 110050 60940
rect 110200 60810 110300 60940
rect 110450 60810 110550 60940
rect 110700 60810 110800 60940
rect 110950 60810 111050 60940
rect 111200 60810 111300 60940
rect 111450 60810 111550 60940
rect 111700 60810 111800 60940
rect 111950 60810 112050 60940
rect 112200 60810 112300 60940
rect 112450 60810 112550 60940
rect 112700 60810 112800 60940
rect 112950 60810 113050 60940
rect 113200 60810 113300 60940
rect 113450 60810 113550 60940
rect 113700 60810 113800 60940
rect 113950 60810 114050 60940
rect 114200 60810 114300 60940
rect 114450 60810 114550 60940
rect 114700 60810 114800 60940
rect 114950 60810 115050 60940
rect 115200 60810 115300 60940
rect 115450 60810 115550 60940
rect 115700 60810 115800 60940
rect 115950 60810 116000 60940
rect 107000 60800 107060 60810
rect 107190 60800 107310 60810
rect 107440 60800 107560 60810
rect 107690 60800 107810 60810
rect 107940 60800 108060 60810
rect 108190 60800 108310 60810
rect 108440 60800 108560 60810
rect 108690 60800 108810 60810
rect 108940 60800 109060 60810
rect 109190 60800 109310 60810
rect 109440 60800 109560 60810
rect 109690 60800 109810 60810
rect 109940 60800 110060 60810
rect 110190 60800 110310 60810
rect 110440 60800 110560 60810
rect 110690 60800 110810 60810
rect 110940 60800 111060 60810
rect 111190 60800 111310 60810
rect 111440 60800 111560 60810
rect 111690 60800 111810 60810
rect 111940 60800 112060 60810
rect 112190 60800 112310 60810
rect 112440 60800 112560 60810
rect 112690 60800 112810 60810
rect 112940 60800 113060 60810
rect 113190 60800 113310 60810
rect 113440 60800 113560 60810
rect 113690 60800 113810 60810
rect 113940 60800 114060 60810
rect 114190 60800 114310 60810
rect 114440 60800 114560 60810
rect 114690 60800 114810 60810
rect 114940 60800 115060 60810
rect 115190 60800 115310 60810
rect 115440 60800 115560 60810
rect 115690 60800 115810 60810
rect 115940 60800 116000 60810
rect 107000 60700 116000 60800
rect 107000 60690 107060 60700
rect 107190 60690 107310 60700
rect 107440 60690 107560 60700
rect 107690 60690 107810 60700
rect 107940 60690 108060 60700
rect 108190 60690 108310 60700
rect 108440 60690 108560 60700
rect 108690 60690 108810 60700
rect 108940 60690 109060 60700
rect 109190 60690 109310 60700
rect 109440 60690 109560 60700
rect 109690 60690 109810 60700
rect 109940 60690 110060 60700
rect 110190 60690 110310 60700
rect 110440 60690 110560 60700
rect 110690 60690 110810 60700
rect 110940 60690 111060 60700
rect 111190 60690 111310 60700
rect 111440 60690 111560 60700
rect 111690 60690 111810 60700
rect 111940 60690 112060 60700
rect 112190 60690 112310 60700
rect 112440 60690 112560 60700
rect 112690 60690 112810 60700
rect 112940 60690 113060 60700
rect 113190 60690 113310 60700
rect 113440 60690 113560 60700
rect 113690 60690 113810 60700
rect 113940 60690 114060 60700
rect 114190 60690 114310 60700
rect 114440 60690 114560 60700
rect 114690 60690 114810 60700
rect 114940 60690 115060 60700
rect 115190 60690 115310 60700
rect 115440 60690 115560 60700
rect 115690 60690 115810 60700
rect 115940 60690 116000 60700
rect 107000 60560 107050 60690
rect 107200 60560 107300 60690
rect 107450 60560 107550 60690
rect 107700 60560 107800 60690
rect 107950 60560 108050 60690
rect 108200 60560 108300 60690
rect 108450 60560 108550 60690
rect 108700 60560 108800 60690
rect 108950 60560 109050 60690
rect 109200 60560 109300 60690
rect 109450 60560 109550 60690
rect 109700 60560 109800 60690
rect 109950 60560 110050 60690
rect 110200 60560 110300 60690
rect 110450 60560 110550 60690
rect 110700 60560 110800 60690
rect 110950 60560 111050 60690
rect 111200 60560 111300 60690
rect 111450 60560 111550 60690
rect 111700 60560 111800 60690
rect 111950 60560 112050 60690
rect 112200 60560 112300 60690
rect 112450 60560 112550 60690
rect 112700 60560 112800 60690
rect 112950 60560 113050 60690
rect 113200 60560 113300 60690
rect 113450 60560 113550 60690
rect 113700 60560 113800 60690
rect 113950 60560 114050 60690
rect 114200 60560 114300 60690
rect 114450 60560 114550 60690
rect 114700 60560 114800 60690
rect 114950 60560 115050 60690
rect 115200 60560 115300 60690
rect 115450 60560 115550 60690
rect 115700 60560 115800 60690
rect 115950 60560 116000 60690
rect 107000 60550 107060 60560
rect 107190 60550 107310 60560
rect 107440 60550 107560 60560
rect 107690 60550 107810 60560
rect 107940 60550 108060 60560
rect 108190 60550 108310 60560
rect 108440 60550 108560 60560
rect 108690 60550 108810 60560
rect 108940 60550 109060 60560
rect 109190 60550 109310 60560
rect 109440 60550 109560 60560
rect 109690 60550 109810 60560
rect 109940 60550 110060 60560
rect 110190 60550 110310 60560
rect 110440 60550 110560 60560
rect 110690 60550 110810 60560
rect 110940 60550 111060 60560
rect 111190 60550 111310 60560
rect 111440 60550 111560 60560
rect 111690 60550 111810 60560
rect 111940 60550 112060 60560
rect 112190 60550 112310 60560
rect 112440 60550 112560 60560
rect 112690 60550 112810 60560
rect 112940 60550 113060 60560
rect 113190 60550 113310 60560
rect 113440 60550 113560 60560
rect 113690 60550 113810 60560
rect 113940 60550 114060 60560
rect 114190 60550 114310 60560
rect 114440 60550 114560 60560
rect 114690 60550 114810 60560
rect 114940 60550 115060 60560
rect 115190 60550 115310 60560
rect 115440 60550 115560 60560
rect 115690 60550 115810 60560
rect 115940 60550 116000 60560
rect 107000 60450 116000 60550
rect 107000 60440 107060 60450
rect 107190 60440 107310 60450
rect 107440 60440 107560 60450
rect 107690 60440 107810 60450
rect 107940 60440 108060 60450
rect 108190 60440 108310 60450
rect 108440 60440 108560 60450
rect 108690 60440 108810 60450
rect 108940 60440 109060 60450
rect 109190 60440 109310 60450
rect 109440 60440 109560 60450
rect 109690 60440 109810 60450
rect 109940 60440 110060 60450
rect 110190 60440 110310 60450
rect 110440 60440 110560 60450
rect 110690 60440 110810 60450
rect 110940 60440 111060 60450
rect 111190 60440 111310 60450
rect 111440 60440 111560 60450
rect 111690 60440 111810 60450
rect 111940 60440 112060 60450
rect 112190 60440 112310 60450
rect 112440 60440 112560 60450
rect 112690 60440 112810 60450
rect 112940 60440 113060 60450
rect 113190 60440 113310 60450
rect 113440 60440 113560 60450
rect 113690 60440 113810 60450
rect 113940 60440 114060 60450
rect 114190 60440 114310 60450
rect 114440 60440 114560 60450
rect 114690 60440 114810 60450
rect 114940 60440 115060 60450
rect 115190 60440 115310 60450
rect 115440 60440 115560 60450
rect 115690 60440 115810 60450
rect 115940 60440 116000 60450
rect 107000 60310 107050 60440
rect 107200 60310 107300 60440
rect 107450 60310 107550 60440
rect 107700 60310 107800 60440
rect 107950 60310 108050 60440
rect 108200 60310 108300 60440
rect 108450 60310 108550 60440
rect 108700 60310 108800 60440
rect 108950 60310 109050 60440
rect 109200 60310 109300 60440
rect 109450 60310 109550 60440
rect 109700 60310 109800 60440
rect 109950 60310 110050 60440
rect 110200 60310 110300 60440
rect 110450 60310 110550 60440
rect 110700 60310 110800 60440
rect 110950 60310 111050 60440
rect 111200 60310 111300 60440
rect 111450 60310 111550 60440
rect 111700 60310 111800 60440
rect 111950 60310 112050 60440
rect 112200 60310 112300 60440
rect 112450 60310 112550 60440
rect 112700 60310 112800 60440
rect 112950 60310 113050 60440
rect 113200 60310 113300 60440
rect 113450 60310 113550 60440
rect 113700 60310 113800 60440
rect 113950 60310 114050 60440
rect 114200 60310 114300 60440
rect 114450 60310 114550 60440
rect 114700 60310 114800 60440
rect 114950 60310 115050 60440
rect 115200 60310 115300 60440
rect 115450 60310 115550 60440
rect 115700 60310 115800 60440
rect 115950 60310 116000 60440
rect 107000 60300 107060 60310
rect 107190 60300 107310 60310
rect 107440 60300 107560 60310
rect 107690 60300 107810 60310
rect 107940 60300 108060 60310
rect 108190 60300 108310 60310
rect 108440 60300 108560 60310
rect 108690 60300 108810 60310
rect 108940 60300 109060 60310
rect 109190 60300 109310 60310
rect 109440 60300 109560 60310
rect 109690 60300 109810 60310
rect 109940 60300 110060 60310
rect 110190 60300 110310 60310
rect 110440 60300 110560 60310
rect 110690 60300 110810 60310
rect 110940 60300 111060 60310
rect 111190 60300 111310 60310
rect 111440 60300 111560 60310
rect 111690 60300 111810 60310
rect 111940 60300 112060 60310
rect 112190 60300 112310 60310
rect 112440 60300 112560 60310
rect 112690 60300 112810 60310
rect 112940 60300 113060 60310
rect 113190 60300 113310 60310
rect 113440 60300 113560 60310
rect 113690 60300 113810 60310
rect 113940 60300 114060 60310
rect 114190 60300 114310 60310
rect 114440 60300 114560 60310
rect 114690 60300 114810 60310
rect 114940 60300 115060 60310
rect 115190 60300 115310 60310
rect 115440 60300 115560 60310
rect 115690 60300 115810 60310
rect 115940 60300 116000 60310
rect 107000 60200 116000 60300
rect 107000 60190 107060 60200
rect 107190 60190 107310 60200
rect 107440 60190 107560 60200
rect 107690 60190 107810 60200
rect 107940 60190 108060 60200
rect 108190 60190 108310 60200
rect 108440 60190 108560 60200
rect 108690 60190 108810 60200
rect 108940 60190 109060 60200
rect 109190 60190 109310 60200
rect 109440 60190 109560 60200
rect 109690 60190 109810 60200
rect 109940 60190 110060 60200
rect 110190 60190 110310 60200
rect 110440 60190 110560 60200
rect 110690 60190 110810 60200
rect 110940 60190 111060 60200
rect 111190 60190 111310 60200
rect 111440 60190 111560 60200
rect 111690 60190 111810 60200
rect 111940 60190 112060 60200
rect 112190 60190 112310 60200
rect 112440 60190 112560 60200
rect 112690 60190 112810 60200
rect 112940 60190 113060 60200
rect 113190 60190 113310 60200
rect 113440 60190 113560 60200
rect 113690 60190 113810 60200
rect 113940 60190 114060 60200
rect 114190 60190 114310 60200
rect 114440 60190 114560 60200
rect 114690 60190 114810 60200
rect 114940 60190 115060 60200
rect 115190 60190 115310 60200
rect 115440 60190 115560 60200
rect 115690 60190 115810 60200
rect 115940 60190 116000 60200
rect 107000 60060 107050 60190
rect 107200 60060 107300 60190
rect 107450 60060 107550 60190
rect 107700 60060 107800 60190
rect 107950 60060 108050 60190
rect 108200 60060 108300 60190
rect 108450 60060 108550 60190
rect 108700 60060 108800 60190
rect 108950 60060 109050 60190
rect 109200 60060 109300 60190
rect 109450 60060 109550 60190
rect 109700 60060 109800 60190
rect 109950 60060 110050 60190
rect 110200 60060 110300 60190
rect 110450 60060 110550 60190
rect 110700 60060 110800 60190
rect 110950 60060 111050 60190
rect 111200 60060 111300 60190
rect 111450 60060 111550 60190
rect 111700 60060 111800 60190
rect 111950 60060 112050 60190
rect 112200 60060 112300 60190
rect 112450 60060 112550 60190
rect 112700 60060 112800 60190
rect 112950 60060 113050 60190
rect 113200 60060 113300 60190
rect 113450 60060 113550 60190
rect 113700 60060 113800 60190
rect 113950 60060 114050 60190
rect 114200 60060 114300 60190
rect 114450 60060 114550 60190
rect 114700 60060 114800 60190
rect 114950 60060 115050 60190
rect 115200 60060 115300 60190
rect 115450 60060 115550 60190
rect 115700 60060 115800 60190
rect 115950 60060 116000 60190
rect 107000 60050 107060 60060
rect 107190 60050 107310 60060
rect 107440 60050 107560 60060
rect 107690 60050 107810 60060
rect 107940 60050 108060 60060
rect 108190 60050 108310 60060
rect 108440 60050 108560 60060
rect 108690 60050 108810 60060
rect 108940 60050 109060 60060
rect 109190 60050 109310 60060
rect 109440 60050 109560 60060
rect 109690 60050 109810 60060
rect 109940 60050 110060 60060
rect 110190 60050 110310 60060
rect 110440 60050 110560 60060
rect 110690 60050 110810 60060
rect 110940 60050 111060 60060
rect 111190 60050 111310 60060
rect 111440 60050 111560 60060
rect 111690 60050 111810 60060
rect 111940 60050 112060 60060
rect 112190 60050 112310 60060
rect 112440 60050 112560 60060
rect 112690 60050 112810 60060
rect 112940 60050 113060 60060
rect 113190 60050 113310 60060
rect 113440 60050 113560 60060
rect 113690 60050 113810 60060
rect 113940 60050 114060 60060
rect 114190 60050 114310 60060
rect 114440 60050 114560 60060
rect 114690 60050 114810 60060
rect 114940 60050 115060 60060
rect 115190 60050 115310 60060
rect 115440 60050 115560 60060
rect 115690 60050 115810 60060
rect 115940 60050 116000 60060
rect 107000 59950 116000 60050
rect 107000 59940 107060 59950
rect 107190 59940 107310 59950
rect 107440 59940 107560 59950
rect 107690 59940 107810 59950
rect 107940 59940 108060 59950
rect 108190 59940 108310 59950
rect 108440 59940 108560 59950
rect 108690 59940 108810 59950
rect 108940 59940 109060 59950
rect 109190 59940 109310 59950
rect 109440 59940 109560 59950
rect 109690 59940 109810 59950
rect 109940 59940 110060 59950
rect 110190 59940 110310 59950
rect 110440 59940 110560 59950
rect 110690 59940 110810 59950
rect 110940 59940 111060 59950
rect 111190 59940 111310 59950
rect 111440 59940 111560 59950
rect 111690 59940 111810 59950
rect 111940 59940 112060 59950
rect 112190 59940 112310 59950
rect 112440 59940 112560 59950
rect 112690 59940 112810 59950
rect 112940 59940 113060 59950
rect 113190 59940 113310 59950
rect 113440 59940 113560 59950
rect 113690 59940 113810 59950
rect 113940 59940 114060 59950
rect 114190 59940 114310 59950
rect 114440 59940 114560 59950
rect 114690 59940 114810 59950
rect 114940 59940 115060 59950
rect 115190 59940 115310 59950
rect 115440 59940 115560 59950
rect 115690 59940 115810 59950
rect 115940 59940 116000 59950
rect 107000 59810 107050 59940
rect 107200 59810 107300 59940
rect 107450 59810 107550 59940
rect 107700 59810 107800 59940
rect 107950 59810 108050 59940
rect 108200 59810 108300 59940
rect 108450 59810 108550 59940
rect 108700 59810 108800 59940
rect 108950 59810 109050 59940
rect 109200 59810 109300 59940
rect 109450 59810 109550 59940
rect 109700 59810 109800 59940
rect 109950 59810 110050 59940
rect 110200 59810 110300 59940
rect 110450 59810 110550 59940
rect 110700 59810 110800 59940
rect 110950 59810 111050 59940
rect 111200 59810 111300 59940
rect 111450 59810 111550 59940
rect 111700 59810 111800 59940
rect 111950 59810 112050 59940
rect 112200 59810 112300 59940
rect 112450 59810 112550 59940
rect 112700 59810 112800 59940
rect 112950 59810 113050 59940
rect 113200 59810 113300 59940
rect 113450 59810 113550 59940
rect 113700 59810 113800 59940
rect 113950 59810 114050 59940
rect 114200 59810 114300 59940
rect 114450 59810 114550 59940
rect 114700 59810 114800 59940
rect 114950 59810 115050 59940
rect 115200 59810 115300 59940
rect 115450 59810 115550 59940
rect 115700 59810 115800 59940
rect 115950 59810 116000 59940
rect 107000 59800 107060 59810
rect 107190 59800 107310 59810
rect 107440 59800 107560 59810
rect 107690 59800 107810 59810
rect 107940 59800 108060 59810
rect 108190 59800 108310 59810
rect 108440 59800 108560 59810
rect 108690 59800 108810 59810
rect 108940 59800 109060 59810
rect 109190 59800 109310 59810
rect 109440 59800 109560 59810
rect 109690 59800 109810 59810
rect 109940 59800 110060 59810
rect 110190 59800 110310 59810
rect 110440 59800 110560 59810
rect 110690 59800 110810 59810
rect 110940 59800 111060 59810
rect 111190 59800 111310 59810
rect 111440 59800 111560 59810
rect 111690 59800 111810 59810
rect 111940 59800 112060 59810
rect 112190 59800 112310 59810
rect 112440 59800 112560 59810
rect 112690 59800 112810 59810
rect 112940 59800 113060 59810
rect 113190 59800 113310 59810
rect 113440 59800 113560 59810
rect 113690 59800 113810 59810
rect 113940 59800 114060 59810
rect 114190 59800 114310 59810
rect 114440 59800 114560 59810
rect 114690 59800 114810 59810
rect 114940 59800 115060 59810
rect 115190 59800 115310 59810
rect 115440 59800 115560 59810
rect 115690 59800 115810 59810
rect 115940 59800 116000 59810
rect 107000 59700 116000 59800
rect 107000 59690 107060 59700
rect 107190 59690 107310 59700
rect 107440 59690 107560 59700
rect 107690 59690 107810 59700
rect 107940 59690 108060 59700
rect 108190 59690 108310 59700
rect 108440 59690 108560 59700
rect 108690 59690 108810 59700
rect 108940 59690 109060 59700
rect 109190 59690 109310 59700
rect 109440 59690 109560 59700
rect 109690 59690 109810 59700
rect 109940 59690 110060 59700
rect 110190 59690 110310 59700
rect 110440 59690 110560 59700
rect 110690 59690 110810 59700
rect 110940 59690 111060 59700
rect 111190 59690 111310 59700
rect 111440 59690 111560 59700
rect 111690 59690 111810 59700
rect 111940 59690 112060 59700
rect 112190 59690 112310 59700
rect 112440 59690 112560 59700
rect 112690 59690 112810 59700
rect 112940 59690 113060 59700
rect 113190 59690 113310 59700
rect 113440 59690 113560 59700
rect 113690 59690 113810 59700
rect 113940 59690 114060 59700
rect 114190 59690 114310 59700
rect 114440 59690 114560 59700
rect 114690 59690 114810 59700
rect 114940 59690 115060 59700
rect 115190 59690 115310 59700
rect 115440 59690 115560 59700
rect 115690 59690 115810 59700
rect 115940 59690 116000 59700
rect 107000 59560 107050 59690
rect 107200 59560 107300 59690
rect 107450 59560 107550 59690
rect 107700 59560 107800 59690
rect 107950 59560 108050 59690
rect 108200 59560 108300 59690
rect 108450 59560 108550 59690
rect 108700 59560 108800 59690
rect 108950 59560 109050 59690
rect 109200 59560 109300 59690
rect 109450 59560 109550 59690
rect 109700 59560 109800 59690
rect 109950 59560 110050 59690
rect 110200 59560 110300 59690
rect 110450 59560 110550 59690
rect 110700 59560 110800 59690
rect 110950 59560 111050 59690
rect 111200 59560 111300 59690
rect 111450 59560 111550 59690
rect 111700 59560 111800 59690
rect 111950 59560 112050 59690
rect 112200 59560 112300 59690
rect 112450 59560 112550 59690
rect 112700 59560 112800 59690
rect 112950 59560 113050 59690
rect 113200 59560 113300 59690
rect 113450 59560 113550 59690
rect 113700 59560 113800 59690
rect 113950 59560 114050 59690
rect 114200 59560 114300 59690
rect 114450 59560 114550 59690
rect 114700 59560 114800 59690
rect 114950 59560 115050 59690
rect 115200 59560 115300 59690
rect 115450 59560 115550 59690
rect 115700 59560 115800 59690
rect 115950 59560 116000 59690
rect 107000 59550 107060 59560
rect 107190 59550 107310 59560
rect 107440 59550 107560 59560
rect 107690 59550 107810 59560
rect 107940 59550 108060 59560
rect 108190 59550 108310 59560
rect 108440 59550 108560 59560
rect 108690 59550 108810 59560
rect 108940 59550 109060 59560
rect 109190 59550 109310 59560
rect 109440 59550 109560 59560
rect 109690 59550 109810 59560
rect 109940 59550 110060 59560
rect 110190 59550 110310 59560
rect 110440 59550 110560 59560
rect 110690 59550 110810 59560
rect 110940 59550 111060 59560
rect 111190 59550 111310 59560
rect 111440 59550 111560 59560
rect 111690 59550 111810 59560
rect 111940 59550 112060 59560
rect 112190 59550 112310 59560
rect 112440 59550 112560 59560
rect 112690 59550 112810 59560
rect 112940 59550 113060 59560
rect 113190 59550 113310 59560
rect 113440 59550 113560 59560
rect 113690 59550 113810 59560
rect 113940 59550 114060 59560
rect 114190 59550 114310 59560
rect 114440 59550 114560 59560
rect 114690 59550 114810 59560
rect 114940 59550 115060 59560
rect 115190 59550 115310 59560
rect 115440 59550 115560 59560
rect 115690 59550 115810 59560
rect 115940 59550 116000 59560
rect 107000 59450 116000 59550
rect 107000 59440 107060 59450
rect 107190 59440 107310 59450
rect 107440 59440 107560 59450
rect 107690 59440 107810 59450
rect 107940 59440 108060 59450
rect 108190 59440 108310 59450
rect 108440 59440 108560 59450
rect 108690 59440 108810 59450
rect 108940 59440 109060 59450
rect 109190 59440 109310 59450
rect 109440 59440 109560 59450
rect 109690 59440 109810 59450
rect 109940 59440 110060 59450
rect 110190 59440 110310 59450
rect 110440 59440 110560 59450
rect 110690 59440 110810 59450
rect 110940 59440 111060 59450
rect 111190 59440 111310 59450
rect 111440 59440 111560 59450
rect 111690 59440 111810 59450
rect 111940 59440 112060 59450
rect 112190 59440 112310 59450
rect 112440 59440 112560 59450
rect 112690 59440 112810 59450
rect 112940 59440 113060 59450
rect 113190 59440 113310 59450
rect 113440 59440 113560 59450
rect 113690 59440 113810 59450
rect 113940 59440 114060 59450
rect 114190 59440 114310 59450
rect 114440 59440 114560 59450
rect 114690 59440 114810 59450
rect 114940 59440 115060 59450
rect 115190 59440 115310 59450
rect 115440 59440 115560 59450
rect 115690 59440 115810 59450
rect 115940 59440 116000 59450
rect 107000 59310 107050 59440
rect 107200 59310 107300 59440
rect 107450 59310 107550 59440
rect 107700 59310 107800 59440
rect 107950 59310 108050 59440
rect 108200 59310 108300 59440
rect 108450 59310 108550 59440
rect 108700 59310 108800 59440
rect 108950 59310 109050 59440
rect 109200 59310 109300 59440
rect 109450 59310 109550 59440
rect 109700 59310 109800 59440
rect 109950 59310 110050 59440
rect 110200 59310 110300 59440
rect 110450 59310 110550 59440
rect 110700 59310 110800 59440
rect 110950 59310 111050 59440
rect 111200 59310 111300 59440
rect 111450 59310 111550 59440
rect 111700 59310 111800 59440
rect 111950 59310 112050 59440
rect 112200 59310 112300 59440
rect 112450 59310 112550 59440
rect 112700 59310 112800 59440
rect 112950 59310 113050 59440
rect 113200 59310 113300 59440
rect 113450 59310 113550 59440
rect 113700 59310 113800 59440
rect 113950 59310 114050 59440
rect 114200 59310 114300 59440
rect 114450 59310 114550 59440
rect 114700 59310 114800 59440
rect 114950 59310 115050 59440
rect 115200 59310 115300 59440
rect 115450 59310 115550 59440
rect 115700 59310 115800 59440
rect 115950 59310 116000 59440
rect 107000 59300 107060 59310
rect 107190 59300 107310 59310
rect 107440 59300 107560 59310
rect 107690 59300 107810 59310
rect 107940 59300 108060 59310
rect 108190 59300 108310 59310
rect 108440 59300 108560 59310
rect 108690 59300 108810 59310
rect 108940 59300 109060 59310
rect 109190 59300 109310 59310
rect 109440 59300 109560 59310
rect 109690 59300 109810 59310
rect 109940 59300 110060 59310
rect 110190 59300 110310 59310
rect 110440 59300 110560 59310
rect 110690 59300 110810 59310
rect 110940 59300 111060 59310
rect 111190 59300 111310 59310
rect 111440 59300 111560 59310
rect 111690 59300 111810 59310
rect 111940 59300 112060 59310
rect 112190 59300 112310 59310
rect 112440 59300 112560 59310
rect 112690 59300 112810 59310
rect 112940 59300 113060 59310
rect 113190 59300 113310 59310
rect 113440 59300 113560 59310
rect 113690 59300 113810 59310
rect 113940 59300 114060 59310
rect 114190 59300 114310 59310
rect 114440 59300 114560 59310
rect 114690 59300 114810 59310
rect 114940 59300 115060 59310
rect 115190 59300 115310 59310
rect 115440 59300 115560 59310
rect 115690 59300 115810 59310
rect 115940 59300 116000 59310
rect 107000 59200 116000 59300
rect 107000 59190 107060 59200
rect 107190 59190 107310 59200
rect 107440 59190 107560 59200
rect 107690 59190 107810 59200
rect 107940 59190 108060 59200
rect 108190 59190 108310 59200
rect 108440 59190 108560 59200
rect 108690 59190 108810 59200
rect 108940 59190 109060 59200
rect 109190 59190 109310 59200
rect 109440 59190 109560 59200
rect 109690 59190 109810 59200
rect 109940 59190 110060 59200
rect 110190 59190 110310 59200
rect 110440 59190 110560 59200
rect 110690 59190 110810 59200
rect 110940 59190 111060 59200
rect 111190 59190 111310 59200
rect 111440 59190 111560 59200
rect 111690 59190 111810 59200
rect 111940 59190 112060 59200
rect 112190 59190 112310 59200
rect 112440 59190 112560 59200
rect 112690 59190 112810 59200
rect 112940 59190 113060 59200
rect 113190 59190 113310 59200
rect 113440 59190 113560 59200
rect 113690 59190 113810 59200
rect 113940 59190 114060 59200
rect 114190 59190 114310 59200
rect 114440 59190 114560 59200
rect 114690 59190 114810 59200
rect 114940 59190 115060 59200
rect 115190 59190 115310 59200
rect 115440 59190 115560 59200
rect 115690 59190 115810 59200
rect 115940 59190 116000 59200
rect 107000 59060 107050 59190
rect 107200 59060 107300 59190
rect 107450 59060 107550 59190
rect 107700 59060 107800 59190
rect 107950 59060 108050 59190
rect 108200 59060 108300 59190
rect 108450 59060 108550 59190
rect 108700 59060 108800 59190
rect 108950 59060 109050 59190
rect 109200 59060 109300 59190
rect 109450 59060 109550 59190
rect 109700 59060 109800 59190
rect 109950 59060 110050 59190
rect 110200 59060 110300 59190
rect 110450 59060 110550 59190
rect 110700 59060 110800 59190
rect 110950 59060 111050 59190
rect 111200 59060 111300 59190
rect 111450 59060 111550 59190
rect 111700 59060 111800 59190
rect 111950 59060 112050 59190
rect 112200 59060 112300 59190
rect 112450 59060 112550 59190
rect 112700 59060 112800 59190
rect 112950 59060 113050 59190
rect 113200 59060 113300 59190
rect 113450 59060 113550 59190
rect 113700 59060 113800 59190
rect 113950 59060 114050 59190
rect 114200 59060 114300 59190
rect 114450 59060 114550 59190
rect 114700 59060 114800 59190
rect 114950 59060 115050 59190
rect 115200 59060 115300 59190
rect 115450 59060 115550 59190
rect 115700 59060 115800 59190
rect 115950 59060 116000 59190
rect 107000 59050 107060 59060
rect 107190 59050 107310 59060
rect 107440 59050 107560 59060
rect 107690 59050 107810 59060
rect 107940 59050 108060 59060
rect 108190 59050 108310 59060
rect 108440 59050 108560 59060
rect 108690 59050 108810 59060
rect 108940 59050 109060 59060
rect 109190 59050 109310 59060
rect 109440 59050 109560 59060
rect 109690 59050 109810 59060
rect 109940 59050 110060 59060
rect 110190 59050 110310 59060
rect 110440 59050 110560 59060
rect 110690 59050 110810 59060
rect 110940 59050 111060 59060
rect 111190 59050 111310 59060
rect 111440 59050 111560 59060
rect 111690 59050 111810 59060
rect 111940 59050 112060 59060
rect 112190 59050 112310 59060
rect 112440 59050 112560 59060
rect 112690 59050 112810 59060
rect 112940 59050 113060 59060
rect 113190 59050 113310 59060
rect 113440 59050 113560 59060
rect 113690 59050 113810 59060
rect 113940 59050 114060 59060
rect 114190 59050 114310 59060
rect 114440 59050 114560 59060
rect 114690 59050 114810 59060
rect 114940 59050 115060 59060
rect 115190 59050 115310 59060
rect 115440 59050 115560 59060
rect 115690 59050 115810 59060
rect 115940 59050 116000 59060
rect 107000 58950 116000 59050
rect 107000 58940 107060 58950
rect 107190 58940 107310 58950
rect 107440 58940 107560 58950
rect 107690 58940 107810 58950
rect 107940 58940 108060 58950
rect 108190 58940 108310 58950
rect 108440 58940 108560 58950
rect 108690 58940 108810 58950
rect 108940 58940 109060 58950
rect 109190 58940 109310 58950
rect 109440 58940 109560 58950
rect 109690 58940 109810 58950
rect 109940 58940 110060 58950
rect 110190 58940 110310 58950
rect 110440 58940 110560 58950
rect 110690 58940 110810 58950
rect 110940 58940 111060 58950
rect 111190 58940 111310 58950
rect 111440 58940 111560 58950
rect 111690 58940 111810 58950
rect 111940 58940 112060 58950
rect 112190 58940 112310 58950
rect 112440 58940 112560 58950
rect 112690 58940 112810 58950
rect 112940 58940 113060 58950
rect 113190 58940 113310 58950
rect 113440 58940 113560 58950
rect 113690 58940 113810 58950
rect 113940 58940 114060 58950
rect 114190 58940 114310 58950
rect 114440 58940 114560 58950
rect 114690 58940 114810 58950
rect 114940 58940 115060 58950
rect 115190 58940 115310 58950
rect 115440 58940 115560 58950
rect 115690 58940 115810 58950
rect 115940 58940 116000 58950
rect 107000 58810 107050 58940
rect 107200 58810 107300 58940
rect 107450 58810 107550 58940
rect 107700 58810 107800 58940
rect 107950 58810 108050 58940
rect 108200 58810 108300 58940
rect 108450 58810 108550 58940
rect 108700 58810 108800 58940
rect 108950 58810 109050 58940
rect 109200 58810 109300 58940
rect 109450 58810 109550 58940
rect 109700 58810 109800 58940
rect 109950 58810 110050 58940
rect 110200 58810 110300 58940
rect 110450 58810 110550 58940
rect 110700 58810 110800 58940
rect 110950 58810 111050 58940
rect 111200 58810 111300 58940
rect 111450 58810 111550 58940
rect 111700 58810 111800 58940
rect 111950 58810 112050 58940
rect 112200 58810 112300 58940
rect 112450 58810 112550 58940
rect 112700 58810 112800 58940
rect 112950 58810 113050 58940
rect 113200 58810 113300 58940
rect 113450 58810 113550 58940
rect 113700 58810 113800 58940
rect 113950 58810 114050 58940
rect 114200 58810 114300 58940
rect 114450 58810 114550 58940
rect 114700 58810 114800 58940
rect 114950 58810 115050 58940
rect 115200 58810 115300 58940
rect 115450 58810 115550 58940
rect 115700 58810 115800 58940
rect 115950 58810 116000 58940
rect 107000 58800 107060 58810
rect 107190 58800 107310 58810
rect 107440 58800 107560 58810
rect 107690 58800 107810 58810
rect 107940 58800 108060 58810
rect 108190 58800 108310 58810
rect 108440 58800 108560 58810
rect 108690 58800 108810 58810
rect 108940 58800 109060 58810
rect 109190 58800 109310 58810
rect 109440 58800 109560 58810
rect 109690 58800 109810 58810
rect 109940 58800 110060 58810
rect 110190 58800 110310 58810
rect 110440 58800 110560 58810
rect 110690 58800 110810 58810
rect 110940 58800 111060 58810
rect 111190 58800 111310 58810
rect 111440 58800 111560 58810
rect 111690 58800 111810 58810
rect 111940 58800 112060 58810
rect 112190 58800 112310 58810
rect 112440 58800 112560 58810
rect 112690 58800 112810 58810
rect 112940 58800 113060 58810
rect 113190 58800 113310 58810
rect 113440 58800 113560 58810
rect 113690 58800 113810 58810
rect 113940 58800 114060 58810
rect 114190 58800 114310 58810
rect 114440 58800 114560 58810
rect 114690 58800 114810 58810
rect 114940 58800 115060 58810
rect 115190 58800 115310 58810
rect 115440 58800 115560 58810
rect 115690 58800 115810 58810
rect 115940 58800 116000 58810
rect 107000 58700 116000 58800
rect 107000 58690 107060 58700
rect 107190 58690 107310 58700
rect 107440 58690 107560 58700
rect 107690 58690 107810 58700
rect 107940 58690 108060 58700
rect 108190 58690 108310 58700
rect 108440 58690 108560 58700
rect 108690 58690 108810 58700
rect 108940 58690 109060 58700
rect 109190 58690 109310 58700
rect 109440 58690 109560 58700
rect 109690 58690 109810 58700
rect 109940 58690 110060 58700
rect 110190 58690 110310 58700
rect 110440 58690 110560 58700
rect 110690 58690 110810 58700
rect 110940 58690 111060 58700
rect 111190 58690 111310 58700
rect 111440 58690 111560 58700
rect 111690 58690 111810 58700
rect 111940 58690 112060 58700
rect 112190 58690 112310 58700
rect 112440 58690 112560 58700
rect 112690 58690 112810 58700
rect 112940 58690 113060 58700
rect 113190 58690 113310 58700
rect 113440 58690 113560 58700
rect 113690 58690 113810 58700
rect 113940 58690 114060 58700
rect 114190 58690 114310 58700
rect 114440 58690 114560 58700
rect 114690 58690 114810 58700
rect 114940 58690 115060 58700
rect 115190 58690 115310 58700
rect 115440 58690 115560 58700
rect 115690 58690 115810 58700
rect 115940 58690 116000 58700
rect 107000 58560 107050 58690
rect 107200 58560 107300 58690
rect 107450 58560 107550 58690
rect 107700 58560 107800 58690
rect 107950 58560 108050 58690
rect 108200 58560 108300 58690
rect 108450 58560 108550 58690
rect 108700 58560 108800 58690
rect 108950 58560 109050 58690
rect 109200 58560 109300 58690
rect 109450 58560 109550 58690
rect 109700 58560 109800 58690
rect 109950 58560 110050 58690
rect 110200 58560 110300 58690
rect 110450 58560 110550 58690
rect 110700 58560 110800 58690
rect 110950 58560 111050 58690
rect 111200 58560 111300 58690
rect 111450 58560 111550 58690
rect 111700 58560 111800 58690
rect 111950 58560 112050 58690
rect 112200 58560 112300 58690
rect 112450 58560 112550 58690
rect 112700 58560 112800 58690
rect 112950 58560 113050 58690
rect 113200 58560 113300 58690
rect 113450 58560 113550 58690
rect 113700 58560 113800 58690
rect 113950 58560 114050 58690
rect 114200 58560 114300 58690
rect 114450 58560 114550 58690
rect 114700 58560 114800 58690
rect 114950 58560 115050 58690
rect 115200 58560 115300 58690
rect 115450 58560 115550 58690
rect 115700 58560 115800 58690
rect 115950 58560 116000 58690
rect 107000 58550 107060 58560
rect 107190 58550 107310 58560
rect 107440 58550 107560 58560
rect 107690 58550 107810 58560
rect 107940 58550 108060 58560
rect 108190 58550 108310 58560
rect 108440 58550 108560 58560
rect 108690 58550 108810 58560
rect 108940 58550 109060 58560
rect 109190 58550 109310 58560
rect 109440 58550 109560 58560
rect 109690 58550 109810 58560
rect 109940 58550 110060 58560
rect 110190 58550 110310 58560
rect 110440 58550 110560 58560
rect 110690 58550 110810 58560
rect 110940 58550 111060 58560
rect 111190 58550 111310 58560
rect 111440 58550 111560 58560
rect 111690 58550 111810 58560
rect 111940 58550 112060 58560
rect 112190 58550 112310 58560
rect 112440 58550 112560 58560
rect 112690 58550 112810 58560
rect 112940 58550 113060 58560
rect 113190 58550 113310 58560
rect 113440 58550 113560 58560
rect 113690 58550 113810 58560
rect 113940 58550 114060 58560
rect 114190 58550 114310 58560
rect 114440 58550 114560 58560
rect 114690 58550 114810 58560
rect 114940 58550 115060 58560
rect 115190 58550 115310 58560
rect 115440 58550 115560 58560
rect 115690 58550 115810 58560
rect 115940 58550 116000 58560
rect 107000 58450 116000 58550
rect 107000 58440 107060 58450
rect 107190 58440 107310 58450
rect 107440 58440 107560 58450
rect 107690 58440 107810 58450
rect 107940 58440 108060 58450
rect 108190 58440 108310 58450
rect 108440 58440 108560 58450
rect 108690 58440 108810 58450
rect 108940 58440 109060 58450
rect 109190 58440 109310 58450
rect 109440 58440 109560 58450
rect 109690 58440 109810 58450
rect 109940 58440 110060 58450
rect 110190 58440 110310 58450
rect 110440 58440 110560 58450
rect 110690 58440 110810 58450
rect 110940 58440 111060 58450
rect 111190 58440 111310 58450
rect 111440 58440 111560 58450
rect 111690 58440 111810 58450
rect 111940 58440 112060 58450
rect 112190 58440 112310 58450
rect 112440 58440 112560 58450
rect 112690 58440 112810 58450
rect 112940 58440 113060 58450
rect 113190 58440 113310 58450
rect 113440 58440 113560 58450
rect 113690 58440 113810 58450
rect 113940 58440 114060 58450
rect 114190 58440 114310 58450
rect 114440 58440 114560 58450
rect 114690 58440 114810 58450
rect 114940 58440 115060 58450
rect 115190 58440 115310 58450
rect 115440 58440 115560 58450
rect 115690 58440 115810 58450
rect 115940 58440 116000 58450
rect 107000 58310 107050 58440
rect 107200 58310 107300 58440
rect 107450 58310 107550 58440
rect 107700 58310 107800 58440
rect 107950 58310 108050 58440
rect 108200 58310 108300 58440
rect 108450 58310 108550 58440
rect 108700 58310 108800 58440
rect 108950 58310 109050 58440
rect 109200 58310 109300 58440
rect 109450 58310 109550 58440
rect 109700 58310 109800 58440
rect 109950 58310 110050 58440
rect 110200 58310 110300 58440
rect 110450 58310 110550 58440
rect 110700 58310 110800 58440
rect 110950 58310 111050 58440
rect 111200 58310 111300 58440
rect 111450 58310 111550 58440
rect 111700 58310 111800 58440
rect 111950 58310 112050 58440
rect 112200 58310 112300 58440
rect 112450 58310 112550 58440
rect 112700 58310 112800 58440
rect 112950 58310 113050 58440
rect 113200 58310 113300 58440
rect 113450 58310 113550 58440
rect 113700 58310 113800 58440
rect 113950 58310 114050 58440
rect 114200 58310 114300 58440
rect 114450 58310 114550 58440
rect 114700 58310 114800 58440
rect 114950 58310 115050 58440
rect 115200 58310 115300 58440
rect 115450 58310 115550 58440
rect 115700 58310 115800 58440
rect 115950 58310 116000 58440
rect 107000 58300 107060 58310
rect 107190 58300 107310 58310
rect 107440 58300 107560 58310
rect 107690 58300 107810 58310
rect 107940 58300 108060 58310
rect 108190 58300 108310 58310
rect 108440 58300 108560 58310
rect 108690 58300 108810 58310
rect 108940 58300 109060 58310
rect 109190 58300 109310 58310
rect 109440 58300 109560 58310
rect 109690 58300 109810 58310
rect 109940 58300 110060 58310
rect 110190 58300 110310 58310
rect 110440 58300 110560 58310
rect 110690 58300 110810 58310
rect 110940 58300 111060 58310
rect 111190 58300 111310 58310
rect 111440 58300 111560 58310
rect 111690 58300 111810 58310
rect 111940 58300 112060 58310
rect 112190 58300 112310 58310
rect 112440 58300 112560 58310
rect 112690 58300 112810 58310
rect 112940 58300 113060 58310
rect 113190 58300 113310 58310
rect 113440 58300 113560 58310
rect 113690 58300 113810 58310
rect 113940 58300 114060 58310
rect 114190 58300 114310 58310
rect 114440 58300 114560 58310
rect 114690 58300 114810 58310
rect 114940 58300 115060 58310
rect 115190 58300 115310 58310
rect 115440 58300 115560 58310
rect 115690 58300 115810 58310
rect 115940 58300 116000 58310
rect 107000 58200 116000 58300
rect 107000 58190 107060 58200
rect 107190 58190 107310 58200
rect 107440 58190 107560 58200
rect 107690 58190 107810 58200
rect 107940 58190 108060 58200
rect 108190 58190 108310 58200
rect 108440 58190 108560 58200
rect 108690 58190 108810 58200
rect 108940 58190 109060 58200
rect 109190 58190 109310 58200
rect 109440 58190 109560 58200
rect 109690 58190 109810 58200
rect 109940 58190 110060 58200
rect 110190 58190 110310 58200
rect 110440 58190 110560 58200
rect 110690 58190 110810 58200
rect 110940 58190 111060 58200
rect 111190 58190 111310 58200
rect 111440 58190 111560 58200
rect 111690 58190 111810 58200
rect 111940 58190 112060 58200
rect 112190 58190 112310 58200
rect 112440 58190 112560 58200
rect 112690 58190 112810 58200
rect 112940 58190 113060 58200
rect 113190 58190 113310 58200
rect 113440 58190 113560 58200
rect 113690 58190 113810 58200
rect 113940 58190 114060 58200
rect 114190 58190 114310 58200
rect 114440 58190 114560 58200
rect 114690 58190 114810 58200
rect 114940 58190 115060 58200
rect 115190 58190 115310 58200
rect 115440 58190 115560 58200
rect 115690 58190 115810 58200
rect 115940 58190 116000 58200
rect 107000 58060 107050 58190
rect 107200 58060 107300 58190
rect 107450 58060 107550 58190
rect 107700 58060 107800 58190
rect 107950 58060 108050 58190
rect 108200 58060 108300 58190
rect 108450 58060 108550 58190
rect 108700 58060 108800 58190
rect 108950 58060 109050 58190
rect 109200 58060 109300 58190
rect 109450 58060 109550 58190
rect 109700 58060 109800 58190
rect 109950 58060 110050 58190
rect 110200 58060 110300 58190
rect 110450 58060 110550 58190
rect 110700 58060 110800 58190
rect 110950 58060 111050 58190
rect 111200 58060 111300 58190
rect 111450 58060 111550 58190
rect 111700 58060 111800 58190
rect 111950 58060 112050 58190
rect 112200 58060 112300 58190
rect 112450 58060 112550 58190
rect 112700 58060 112800 58190
rect 112950 58060 113050 58190
rect 113200 58060 113300 58190
rect 113450 58060 113550 58190
rect 113700 58060 113800 58190
rect 113950 58060 114050 58190
rect 114200 58060 114300 58190
rect 114450 58060 114550 58190
rect 114700 58060 114800 58190
rect 114950 58060 115050 58190
rect 115200 58060 115300 58190
rect 115450 58060 115550 58190
rect 115700 58060 115800 58190
rect 115950 58060 116000 58190
rect 107000 58050 107060 58060
rect 107190 58050 107310 58060
rect 107440 58050 107560 58060
rect 107690 58050 107810 58060
rect 107940 58050 108060 58060
rect 108190 58050 108310 58060
rect 108440 58050 108560 58060
rect 108690 58050 108810 58060
rect 108940 58050 109060 58060
rect 109190 58050 109310 58060
rect 109440 58050 109560 58060
rect 109690 58050 109810 58060
rect 109940 58050 110060 58060
rect 110190 58050 110310 58060
rect 110440 58050 110560 58060
rect 110690 58050 110810 58060
rect 110940 58050 111060 58060
rect 111190 58050 111310 58060
rect 111440 58050 111560 58060
rect 111690 58050 111810 58060
rect 111940 58050 112060 58060
rect 112190 58050 112310 58060
rect 112440 58050 112560 58060
rect 112690 58050 112810 58060
rect 112940 58050 113060 58060
rect 113190 58050 113310 58060
rect 113440 58050 113560 58060
rect 113690 58050 113810 58060
rect 113940 58050 114060 58060
rect 114190 58050 114310 58060
rect 114440 58050 114560 58060
rect 114690 58050 114810 58060
rect 114940 58050 115060 58060
rect 115190 58050 115310 58060
rect 115440 58050 115560 58060
rect 115690 58050 115810 58060
rect 115940 58050 116000 58060
rect 107000 57950 116000 58050
rect 107000 57940 107060 57950
rect 107190 57940 107310 57950
rect 107440 57940 107560 57950
rect 107690 57940 107810 57950
rect 107940 57940 108060 57950
rect 108190 57940 108310 57950
rect 108440 57940 108560 57950
rect 108690 57940 108810 57950
rect 108940 57940 109060 57950
rect 109190 57940 109310 57950
rect 109440 57940 109560 57950
rect 109690 57940 109810 57950
rect 109940 57940 110060 57950
rect 110190 57940 110310 57950
rect 110440 57940 110560 57950
rect 110690 57940 110810 57950
rect 110940 57940 111060 57950
rect 111190 57940 111310 57950
rect 111440 57940 111560 57950
rect 111690 57940 111810 57950
rect 111940 57940 112060 57950
rect 112190 57940 112310 57950
rect 112440 57940 112560 57950
rect 112690 57940 112810 57950
rect 112940 57940 113060 57950
rect 113190 57940 113310 57950
rect 113440 57940 113560 57950
rect 113690 57940 113810 57950
rect 113940 57940 114060 57950
rect 114190 57940 114310 57950
rect 114440 57940 114560 57950
rect 114690 57940 114810 57950
rect 114940 57940 115060 57950
rect 115190 57940 115310 57950
rect 115440 57940 115560 57950
rect 115690 57940 115810 57950
rect 115940 57940 116000 57950
rect 107000 57810 107050 57940
rect 107200 57810 107300 57940
rect 107450 57810 107550 57940
rect 107700 57810 107800 57940
rect 107950 57810 108050 57940
rect 108200 57810 108300 57940
rect 108450 57810 108550 57940
rect 108700 57810 108800 57940
rect 108950 57810 109050 57940
rect 109200 57810 109300 57940
rect 109450 57810 109550 57940
rect 109700 57810 109800 57940
rect 109950 57810 110050 57940
rect 110200 57810 110300 57940
rect 110450 57810 110550 57940
rect 110700 57810 110800 57940
rect 110950 57810 111050 57940
rect 111200 57810 111300 57940
rect 111450 57810 111550 57940
rect 111700 57810 111800 57940
rect 111950 57810 112050 57940
rect 112200 57810 112300 57940
rect 112450 57810 112550 57940
rect 112700 57810 112800 57940
rect 112950 57810 113050 57940
rect 113200 57810 113300 57940
rect 113450 57810 113550 57940
rect 113700 57810 113800 57940
rect 113950 57810 114050 57940
rect 114200 57810 114300 57940
rect 114450 57810 114550 57940
rect 114700 57810 114800 57940
rect 114950 57810 115050 57940
rect 115200 57810 115300 57940
rect 115450 57810 115550 57940
rect 115700 57810 115800 57940
rect 115950 57810 116000 57940
rect 107000 57800 107060 57810
rect 107190 57800 107310 57810
rect 107440 57800 107560 57810
rect 107690 57800 107810 57810
rect 107940 57800 108060 57810
rect 108190 57800 108310 57810
rect 108440 57800 108560 57810
rect 108690 57800 108810 57810
rect 108940 57800 109060 57810
rect 109190 57800 109310 57810
rect 109440 57800 109560 57810
rect 109690 57800 109810 57810
rect 109940 57800 110060 57810
rect 110190 57800 110310 57810
rect 110440 57800 110560 57810
rect 110690 57800 110810 57810
rect 110940 57800 111060 57810
rect 111190 57800 111310 57810
rect 111440 57800 111560 57810
rect 111690 57800 111810 57810
rect 111940 57800 112060 57810
rect 112190 57800 112310 57810
rect 112440 57800 112560 57810
rect 112690 57800 112810 57810
rect 112940 57800 113060 57810
rect 113190 57800 113310 57810
rect 113440 57800 113560 57810
rect 113690 57800 113810 57810
rect 113940 57800 114060 57810
rect 114190 57800 114310 57810
rect 114440 57800 114560 57810
rect 114690 57800 114810 57810
rect 114940 57800 115060 57810
rect 115190 57800 115310 57810
rect 115440 57800 115560 57810
rect 115690 57800 115810 57810
rect 115940 57800 116000 57810
rect 107000 57700 116000 57800
rect 107000 57690 107060 57700
rect 107190 57690 107310 57700
rect 107440 57690 107560 57700
rect 107690 57690 107810 57700
rect 107940 57690 108060 57700
rect 108190 57690 108310 57700
rect 108440 57690 108560 57700
rect 108690 57690 108810 57700
rect 108940 57690 109060 57700
rect 109190 57690 109310 57700
rect 109440 57690 109560 57700
rect 109690 57690 109810 57700
rect 109940 57690 110060 57700
rect 110190 57690 110310 57700
rect 110440 57690 110560 57700
rect 110690 57690 110810 57700
rect 110940 57690 111060 57700
rect 111190 57690 111310 57700
rect 111440 57690 111560 57700
rect 111690 57690 111810 57700
rect 111940 57690 112060 57700
rect 112190 57690 112310 57700
rect 112440 57690 112560 57700
rect 112690 57690 112810 57700
rect 112940 57690 113060 57700
rect 113190 57690 113310 57700
rect 113440 57690 113560 57700
rect 113690 57690 113810 57700
rect 113940 57690 114060 57700
rect 114190 57690 114310 57700
rect 114440 57690 114560 57700
rect 114690 57690 114810 57700
rect 114940 57690 115060 57700
rect 115190 57690 115310 57700
rect 115440 57690 115560 57700
rect 115690 57690 115810 57700
rect 115940 57690 116000 57700
rect 107000 57560 107050 57690
rect 107200 57560 107300 57690
rect 107450 57560 107550 57690
rect 107700 57560 107800 57690
rect 107950 57560 108050 57690
rect 108200 57560 108300 57690
rect 108450 57560 108550 57690
rect 108700 57560 108800 57690
rect 108950 57560 109050 57690
rect 109200 57560 109300 57690
rect 109450 57560 109550 57690
rect 109700 57560 109800 57690
rect 109950 57560 110050 57690
rect 110200 57560 110300 57690
rect 110450 57560 110550 57690
rect 110700 57560 110800 57690
rect 110950 57560 111050 57690
rect 111200 57560 111300 57690
rect 111450 57560 111550 57690
rect 111700 57560 111800 57690
rect 111950 57560 112050 57690
rect 112200 57560 112300 57690
rect 112450 57560 112550 57690
rect 112700 57560 112800 57690
rect 112950 57560 113050 57690
rect 113200 57560 113300 57690
rect 113450 57560 113550 57690
rect 113700 57560 113800 57690
rect 113950 57560 114050 57690
rect 114200 57560 114300 57690
rect 114450 57560 114550 57690
rect 114700 57560 114800 57690
rect 114950 57560 115050 57690
rect 115200 57560 115300 57690
rect 115450 57560 115550 57690
rect 115700 57560 115800 57690
rect 115950 57560 116000 57690
rect 107000 57550 107060 57560
rect 107190 57550 107310 57560
rect 107440 57550 107560 57560
rect 107690 57550 107810 57560
rect 107940 57550 108060 57560
rect 108190 57550 108310 57560
rect 108440 57550 108560 57560
rect 108690 57550 108810 57560
rect 108940 57550 109060 57560
rect 109190 57550 109310 57560
rect 109440 57550 109560 57560
rect 109690 57550 109810 57560
rect 109940 57550 110060 57560
rect 110190 57550 110310 57560
rect 110440 57550 110560 57560
rect 110690 57550 110810 57560
rect 110940 57550 111060 57560
rect 111190 57550 111310 57560
rect 111440 57550 111560 57560
rect 111690 57550 111810 57560
rect 111940 57550 112060 57560
rect 112190 57550 112310 57560
rect 112440 57550 112560 57560
rect 112690 57550 112810 57560
rect 112940 57550 113060 57560
rect 113190 57550 113310 57560
rect 113440 57550 113560 57560
rect 113690 57550 113810 57560
rect 113940 57550 114060 57560
rect 114190 57550 114310 57560
rect 114440 57550 114560 57560
rect 114690 57550 114810 57560
rect 114940 57550 115060 57560
rect 115190 57550 115310 57560
rect 115440 57550 115560 57560
rect 115690 57550 115810 57560
rect 115940 57550 116000 57560
rect 107000 57450 116000 57550
rect 107000 57440 107060 57450
rect 107190 57440 107310 57450
rect 107440 57440 107560 57450
rect 107690 57440 107810 57450
rect 107940 57440 108060 57450
rect 108190 57440 108310 57450
rect 108440 57440 108560 57450
rect 108690 57440 108810 57450
rect 108940 57440 109060 57450
rect 109190 57440 109310 57450
rect 109440 57440 109560 57450
rect 109690 57440 109810 57450
rect 109940 57440 110060 57450
rect 110190 57440 110310 57450
rect 110440 57440 110560 57450
rect 110690 57440 110810 57450
rect 110940 57440 111060 57450
rect 111190 57440 111310 57450
rect 111440 57440 111560 57450
rect 111690 57440 111810 57450
rect 111940 57440 112060 57450
rect 112190 57440 112310 57450
rect 112440 57440 112560 57450
rect 112690 57440 112810 57450
rect 112940 57440 113060 57450
rect 113190 57440 113310 57450
rect 113440 57440 113560 57450
rect 113690 57440 113810 57450
rect 113940 57440 114060 57450
rect 114190 57440 114310 57450
rect 114440 57440 114560 57450
rect 114690 57440 114810 57450
rect 114940 57440 115060 57450
rect 115190 57440 115310 57450
rect 115440 57440 115560 57450
rect 115690 57440 115810 57450
rect 115940 57440 116000 57450
rect 107000 57310 107050 57440
rect 107200 57310 107300 57440
rect 107450 57310 107550 57440
rect 107700 57310 107800 57440
rect 107950 57310 108050 57440
rect 108200 57310 108300 57440
rect 108450 57310 108550 57440
rect 108700 57310 108800 57440
rect 108950 57310 109050 57440
rect 109200 57310 109300 57440
rect 109450 57310 109550 57440
rect 109700 57310 109800 57440
rect 109950 57310 110050 57440
rect 110200 57310 110300 57440
rect 110450 57310 110550 57440
rect 110700 57310 110800 57440
rect 110950 57310 111050 57440
rect 111200 57310 111300 57440
rect 111450 57310 111550 57440
rect 111700 57310 111800 57440
rect 111950 57310 112050 57440
rect 112200 57310 112300 57440
rect 112450 57310 112550 57440
rect 112700 57310 112800 57440
rect 112950 57310 113050 57440
rect 113200 57310 113300 57440
rect 113450 57310 113550 57440
rect 113700 57310 113800 57440
rect 113950 57310 114050 57440
rect 114200 57310 114300 57440
rect 114450 57310 114550 57440
rect 114700 57310 114800 57440
rect 114950 57310 115050 57440
rect 115200 57310 115300 57440
rect 115450 57310 115550 57440
rect 115700 57310 115800 57440
rect 115950 57310 116000 57440
rect 107000 57300 107060 57310
rect 107190 57300 107310 57310
rect 107440 57300 107560 57310
rect 107690 57300 107810 57310
rect 107940 57300 108060 57310
rect 108190 57300 108310 57310
rect 108440 57300 108560 57310
rect 108690 57300 108810 57310
rect 108940 57300 109060 57310
rect 109190 57300 109310 57310
rect 109440 57300 109560 57310
rect 109690 57300 109810 57310
rect 109940 57300 110060 57310
rect 110190 57300 110310 57310
rect 110440 57300 110560 57310
rect 110690 57300 110810 57310
rect 110940 57300 111060 57310
rect 111190 57300 111310 57310
rect 111440 57300 111560 57310
rect 111690 57300 111810 57310
rect 111940 57300 112060 57310
rect 112190 57300 112310 57310
rect 112440 57300 112560 57310
rect 112690 57300 112810 57310
rect 112940 57300 113060 57310
rect 113190 57300 113310 57310
rect 113440 57300 113560 57310
rect 113690 57300 113810 57310
rect 113940 57300 114060 57310
rect 114190 57300 114310 57310
rect 114440 57300 114560 57310
rect 114690 57300 114810 57310
rect 114940 57300 115060 57310
rect 115190 57300 115310 57310
rect 115440 57300 115560 57310
rect 115690 57300 115810 57310
rect 115940 57300 116000 57310
rect 107000 57200 116000 57300
rect 107000 57190 107060 57200
rect 107190 57190 107310 57200
rect 107440 57190 107560 57200
rect 107690 57190 107810 57200
rect 107940 57190 108060 57200
rect 108190 57190 108310 57200
rect 108440 57190 108560 57200
rect 108690 57190 108810 57200
rect 108940 57190 109060 57200
rect 109190 57190 109310 57200
rect 109440 57190 109560 57200
rect 109690 57190 109810 57200
rect 109940 57190 110060 57200
rect 110190 57190 110310 57200
rect 110440 57190 110560 57200
rect 110690 57190 110810 57200
rect 110940 57190 111060 57200
rect 111190 57190 111310 57200
rect 111440 57190 111560 57200
rect 111690 57190 111810 57200
rect 111940 57190 112060 57200
rect 112190 57190 112310 57200
rect 112440 57190 112560 57200
rect 112690 57190 112810 57200
rect 112940 57190 113060 57200
rect 113190 57190 113310 57200
rect 113440 57190 113560 57200
rect 113690 57190 113810 57200
rect 113940 57190 114060 57200
rect 114190 57190 114310 57200
rect 114440 57190 114560 57200
rect 114690 57190 114810 57200
rect 114940 57190 115060 57200
rect 115190 57190 115310 57200
rect 115440 57190 115560 57200
rect 115690 57190 115810 57200
rect 115940 57190 116000 57200
rect 107000 57060 107050 57190
rect 107200 57060 107300 57190
rect 107450 57060 107550 57190
rect 107700 57060 107800 57190
rect 107950 57060 108050 57190
rect 108200 57060 108300 57190
rect 108450 57060 108550 57190
rect 108700 57060 108800 57190
rect 108950 57060 109050 57190
rect 109200 57060 109300 57190
rect 109450 57060 109550 57190
rect 109700 57060 109800 57190
rect 109950 57060 110050 57190
rect 110200 57060 110300 57190
rect 110450 57060 110550 57190
rect 110700 57060 110800 57190
rect 110950 57060 111050 57190
rect 111200 57060 111300 57190
rect 111450 57060 111550 57190
rect 111700 57060 111800 57190
rect 111950 57060 112050 57190
rect 112200 57060 112300 57190
rect 112450 57060 112550 57190
rect 112700 57060 112800 57190
rect 112950 57060 113050 57190
rect 113200 57060 113300 57190
rect 113450 57060 113550 57190
rect 113700 57060 113800 57190
rect 113950 57060 114050 57190
rect 114200 57060 114300 57190
rect 114450 57060 114550 57190
rect 114700 57060 114800 57190
rect 114950 57060 115050 57190
rect 115200 57060 115300 57190
rect 115450 57060 115550 57190
rect 115700 57060 115800 57190
rect 115950 57060 116000 57190
rect 107000 57050 107060 57060
rect 107190 57050 107310 57060
rect 107440 57050 107560 57060
rect 107690 57050 107810 57060
rect 107940 57050 108060 57060
rect 108190 57050 108310 57060
rect 108440 57050 108560 57060
rect 108690 57050 108810 57060
rect 108940 57050 109060 57060
rect 109190 57050 109310 57060
rect 109440 57050 109560 57060
rect 109690 57050 109810 57060
rect 109940 57050 110060 57060
rect 110190 57050 110310 57060
rect 110440 57050 110560 57060
rect 110690 57050 110810 57060
rect 110940 57050 111060 57060
rect 111190 57050 111310 57060
rect 111440 57050 111560 57060
rect 111690 57050 111810 57060
rect 111940 57050 112060 57060
rect 112190 57050 112310 57060
rect 112440 57050 112560 57060
rect 112690 57050 112810 57060
rect 112940 57050 113060 57060
rect 113190 57050 113310 57060
rect 113440 57050 113560 57060
rect 113690 57050 113810 57060
rect 113940 57050 114060 57060
rect 114190 57050 114310 57060
rect 114440 57050 114560 57060
rect 114690 57050 114810 57060
rect 114940 57050 115060 57060
rect 115190 57050 115310 57060
rect 115440 57050 115560 57060
rect 115690 57050 115810 57060
rect 115940 57050 116000 57060
rect 107000 57000 116000 57050
rect 89000 56950 116000 57000
rect 89000 56940 89060 56950
rect 89190 56940 89310 56950
rect 89440 56940 89560 56950
rect 89690 56940 89810 56950
rect 89940 56940 90060 56950
rect 90190 56940 90310 56950
rect 90440 56940 90560 56950
rect 90690 56940 90810 56950
rect 90940 56940 91060 56950
rect 91190 56940 91310 56950
rect 91440 56940 91560 56950
rect 91690 56940 91810 56950
rect 91940 56940 92060 56950
rect 92190 56940 92310 56950
rect 92440 56940 92560 56950
rect 92690 56940 92810 56950
rect 92940 56940 93060 56950
rect 93190 56940 93310 56950
rect 93440 56940 93560 56950
rect 93690 56940 93810 56950
rect 93940 56940 94060 56950
rect 94190 56940 94310 56950
rect 94440 56940 94560 56950
rect 94690 56940 94810 56950
rect 94940 56940 95060 56950
rect 95190 56940 95310 56950
rect 95440 56940 95560 56950
rect 95690 56940 95810 56950
rect 95940 56940 96060 56950
rect 96190 56940 96310 56950
rect 96440 56940 96560 56950
rect 96690 56940 96810 56950
rect 96940 56940 97060 56950
rect 97190 56940 97310 56950
rect 97440 56940 97560 56950
rect 97690 56940 97810 56950
rect 97940 56940 98060 56950
rect 98190 56940 98310 56950
rect 98440 56940 98560 56950
rect 98690 56940 98810 56950
rect 98940 56940 99060 56950
rect 99190 56940 99310 56950
rect 99440 56940 99560 56950
rect 99690 56940 99810 56950
rect 99940 56940 100060 56950
rect 100190 56940 100310 56950
rect 100440 56940 100560 56950
rect 100690 56940 100810 56950
rect 100940 56940 101060 56950
rect 101190 56940 101310 56950
rect 101440 56940 101560 56950
rect 101690 56940 101810 56950
rect 101940 56940 102060 56950
rect 102190 56940 102310 56950
rect 102440 56940 102560 56950
rect 102690 56940 102810 56950
rect 102940 56940 103060 56950
rect 103190 56940 103310 56950
rect 103440 56940 103560 56950
rect 103690 56940 103810 56950
rect 103940 56940 104060 56950
rect 104190 56940 104310 56950
rect 104440 56940 104560 56950
rect 104690 56940 104810 56950
rect 104940 56940 105060 56950
rect 105190 56940 105310 56950
rect 105440 56940 105560 56950
rect 105690 56940 105810 56950
rect 105940 56940 106060 56950
rect 106190 56940 106310 56950
rect 106440 56940 106560 56950
rect 106690 56940 106810 56950
rect 106940 56940 107060 56950
rect 107190 56940 107310 56950
rect 107440 56940 107560 56950
rect 107690 56940 107810 56950
rect 107940 56940 108060 56950
rect 108190 56940 108310 56950
rect 108440 56940 108560 56950
rect 108690 56940 108810 56950
rect 108940 56940 109060 56950
rect 109190 56940 109310 56950
rect 109440 56940 109560 56950
rect 109690 56940 109810 56950
rect 109940 56940 110060 56950
rect 110190 56940 110310 56950
rect 110440 56940 110560 56950
rect 110690 56940 110810 56950
rect 110940 56940 111060 56950
rect 111190 56940 111310 56950
rect 111440 56940 111560 56950
rect 111690 56940 111810 56950
rect 111940 56940 112060 56950
rect 112190 56940 112310 56950
rect 112440 56940 112560 56950
rect 112690 56940 112810 56950
rect 112940 56940 113060 56950
rect 113190 56940 113310 56950
rect 113440 56940 113560 56950
rect 113690 56940 113810 56950
rect 113940 56940 114060 56950
rect 114190 56940 114310 56950
rect 114440 56940 114560 56950
rect 114690 56940 114810 56950
rect 114940 56940 115060 56950
rect 115190 56940 115310 56950
rect 115440 56940 115560 56950
rect 115690 56940 115810 56950
rect 115940 56940 116000 56950
rect 89000 56810 89050 56940
rect 89200 56810 89300 56940
rect 89450 56810 89550 56940
rect 89700 56810 89800 56940
rect 89950 56810 90050 56940
rect 90200 56810 90300 56940
rect 90450 56810 90550 56940
rect 90700 56810 90800 56940
rect 90950 56810 91050 56940
rect 91200 56810 91300 56940
rect 91450 56810 91550 56940
rect 91700 56810 91800 56940
rect 91950 56810 92050 56940
rect 92200 56810 92300 56940
rect 92450 56810 92550 56940
rect 92700 56810 92800 56940
rect 92950 56810 93050 56940
rect 93200 56810 93300 56940
rect 93450 56810 93550 56940
rect 93700 56810 93800 56940
rect 93950 56810 94050 56940
rect 94200 56810 94300 56940
rect 94450 56810 94550 56940
rect 94700 56810 94800 56940
rect 94950 56810 95050 56940
rect 95200 56810 95300 56940
rect 95450 56810 95550 56940
rect 95700 56810 95800 56940
rect 95950 56810 96050 56940
rect 96200 56810 96300 56940
rect 96450 56810 96550 56940
rect 96700 56810 96800 56940
rect 96950 56810 97050 56940
rect 97200 56810 97300 56940
rect 97450 56810 97550 56940
rect 97700 56810 97800 56940
rect 97950 56810 98050 56940
rect 98200 56810 98300 56940
rect 98450 56810 98550 56940
rect 98700 56810 98800 56940
rect 98950 56810 99050 56940
rect 99200 56810 99300 56940
rect 99450 56810 99550 56940
rect 99700 56810 99800 56940
rect 99950 56810 100050 56940
rect 100200 56810 100300 56940
rect 100450 56810 100550 56940
rect 100700 56810 100800 56940
rect 100950 56810 101050 56940
rect 101200 56810 101300 56940
rect 101450 56810 101550 56940
rect 101700 56810 101800 56940
rect 101950 56810 102050 56940
rect 102200 56810 102300 56940
rect 102450 56810 102550 56940
rect 102700 56810 102800 56940
rect 102950 56810 103050 56940
rect 103200 56810 103300 56940
rect 103450 56810 103550 56940
rect 103700 56810 103800 56940
rect 103950 56810 104050 56940
rect 104200 56810 104300 56940
rect 104450 56810 104550 56940
rect 104700 56810 104800 56940
rect 104950 56810 105050 56940
rect 105200 56810 105300 56940
rect 105450 56810 105550 56940
rect 105700 56810 105800 56940
rect 105950 56810 106050 56940
rect 106200 56810 106300 56940
rect 106450 56810 106550 56940
rect 106700 56810 106800 56940
rect 106950 56810 107050 56940
rect 107200 56810 107300 56940
rect 107450 56810 107550 56940
rect 107700 56810 107800 56940
rect 107950 56810 108050 56940
rect 108200 56810 108300 56940
rect 108450 56810 108550 56940
rect 108700 56810 108800 56940
rect 108950 56810 109050 56940
rect 109200 56810 109300 56940
rect 109450 56810 109550 56940
rect 109700 56810 109800 56940
rect 109950 56810 110050 56940
rect 110200 56810 110300 56940
rect 110450 56810 110550 56940
rect 110700 56810 110800 56940
rect 110950 56810 111050 56940
rect 111200 56810 111300 56940
rect 111450 56810 111550 56940
rect 111700 56810 111800 56940
rect 111950 56810 112050 56940
rect 112200 56810 112300 56940
rect 112450 56810 112550 56940
rect 112700 56810 112800 56940
rect 112950 56810 113050 56940
rect 113200 56810 113300 56940
rect 113450 56810 113550 56940
rect 113700 56810 113800 56940
rect 113950 56810 114050 56940
rect 114200 56810 114300 56940
rect 114450 56810 114550 56940
rect 114700 56810 114800 56940
rect 114950 56810 115050 56940
rect 115200 56810 115300 56940
rect 115450 56810 115550 56940
rect 115700 56810 115800 56940
rect 115950 56810 116000 56940
rect 89000 56800 89060 56810
rect 89190 56800 89310 56810
rect 89440 56800 89560 56810
rect 89690 56800 89810 56810
rect 89940 56800 90060 56810
rect 90190 56800 90310 56810
rect 90440 56800 90560 56810
rect 90690 56800 90810 56810
rect 90940 56800 91060 56810
rect 91190 56800 91310 56810
rect 91440 56800 91560 56810
rect 91690 56800 91810 56810
rect 91940 56800 92060 56810
rect 92190 56800 92310 56810
rect 92440 56800 92560 56810
rect 92690 56800 92810 56810
rect 92940 56800 93060 56810
rect 93190 56800 93310 56810
rect 93440 56800 93560 56810
rect 93690 56800 93810 56810
rect 93940 56800 94060 56810
rect 94190 56800 94310 56810
rect 94440 56800 94560 56810
rect 94690 56800 94810 56810
rect 94940 56800 95060 56810
rect 95190 56800 95310 56810
rect 95440 56800 95560 56810
rect 95690 56800 95810 56810
rect 95940 56800 96060 56810
rect 96190 56800 96310 56810
rect 96440 56800 96560 56810
rect 96690 56800 96810 56810
rect 96940 56800 97060 56810
rect 97190 56800 97310 56810
rect 97440 56800 97560 56810
rect 97690 56800 97810 56810
rect 97940 56800 98060 56810
rect 98190 56800 98310 56810
rect 98440 56800 98560 56810
rect 98690 56800 98810 56810
rect 98940 56800 99060 56810
rect 99190 56800 99310 56810
rect 99440 56800 99560 56810
rect 99690 56800 99810 56810
rect 99940 56800 100060 56810
rect 100190 56800 100310 56810
rect 100440 56800 100560 56810
rect 100690 56800 100810 56810
rect 100940 56800 101060 56810
rect 101190 56800 101310 56810
rect 101440 56800 101560 56810
rect 101690 56800 101810 56810
rect 101940 56800 102060 56810
rect 102190 56800 102310 56810
rect 102440 56800 102560 56810
rect 102690 56800 102810 56810
rect 102940 56800 103060 56810
rect 103190 56800 103310 56810
rect 103440 56800 103560 56810
rect 103690 56800 103810 56810
rect 103940 56800 104060 56810
rect 104190 56800 104310 56810
rect 104440 56800 104560 56810
rect 104690 56800 104810 56810
rect 104940 56800 105060 56810
rect 105190 56800 105310 56810
rect 105440 56800 105560 56810
rect 105690 56800 105810 56810
rect 105940 56800 106060 56810
rect 106190 56800 106310 56810
rect 106440 56800 106560 56810
rect 106690 56800 106810 56810
rect 106940 56800 107060 56810
rect 107190 56800 107310 56810
rect 107440 56800 107560 56810
rect 107690 56800 107810 56810
rect 107940 56800 108060 56810
rect 108190 56800 108310 56810
rect 108440 56800 108560 56810
rect 108690 56800 108810 56810
rect 108940 56800 109060 56810
rect 109190 56800 109310 56810
rect 109440 56800 109560 56810
rect 109690 56800 109810 56810
rect 109940 56800 110060 56810
rect 110190 56800 110310 56810
rect 110440 56800 110560 56810
rect 110690 56800 110810 56810
rect 110940 56800 111060 56810
rect 111190 56800 111310 56810
rect 111440 56800 111560 56810
rect 111690 56800 111810 56810
rect 111940 56800 112060 56810
rect 112190 56800 112310 56810
rect 112440 56800 112560 56810
rect 112690 56800 112810 56810
rect 112940 56800 113060 56810
rect 113190 56800 113310 56810
rect 113440 56800 113560 56810
rect 113690 56800 113810 56810
rect 113940 56800 114060 56810
rect 114190 56800 114310 56810
rect 114440 56800 114560 56810
rect 114690 56800 114810 56810
rect 114940 56800 115060 56810
rect 115190 56800 115310 56810
rect 115440 56800 115560 56810
rect 115690 56800 115810 56810
rect 115940 56800 116000 56810
rect 89000 56700 116000 56800
rect 89000 56690 89060 56700
rect 89190 56690 89310 56700
rect 89440 56690 89560 56700
rect 89690 56690 89810 56700
rect 89940 56690 90060 56700
rect 90190 56690 90310 56700
rect 90440 56690 90560 56700
rect 90690 56690 90810 56700
rect 90940 56690 91060 56700
rect 91190 56690 91310 56700
rect 91440 56690 91560 56700
rect 91690 56690 91810 56700
rect 91940 56690 92060 56700
rect 92190 56690 92310 56700
rect 92440 56690 92560 56700
rect 92690 56690 92810 56700
rect 92940 56690 93060 56700
rect 93190 56690 93310 56700
rect 93440 56690 93560 56700
rect 93690 56690 93810 56700
rect 93940 56690 94060 56700
rect 94190 56690 94310 56700
rect 94440 56690 94560 56700
rect 94690 56690 94810 56700
rect 94940 56690 95060 56700
rect 95190 56690 95310 56700
rect 95440 56690 95560 56700
rect 95690 56690 95810 56700
rect 95940 56690 96060 56700
rect 96190 56690 96310 56700
rect 96440 56690 96560 56700
rect 96690 56690 96810 56700
rect 96940 56690 97060 56700
rect 97190 56690 97310 56700
rect 97440 56690 97560 56700
rect 97690 56690 97810 56700
rect 97940 56690 98060 56700
rect 98190 56690 98310 56700
rect 98440 56690 98560 56700
rect 98690 56690 98810 56700
rect 98940 56690 99060 56700
rect 99190 56690 99310 56700
rect 99440 56690 99560 56700
rect 99690 56690 99810 56700
rect 99940 56690 100060 56700
rect 100190 56690 100310 56700
rect 100440 56690 100560 56700
rect 100690 56690 100810 56700
rect 100940 56690 101060 56700
rect 101190 56690 101310 56700
rect 101440 56690 101560 56700
rect 101690 56690 101810 56700
rect 101940 56690 102060 56700
rect 102190 56690 102310 56700
rect 102440 56690 102560 56700
rect 102690 56690 102810 56700
rect 102940 56690 103060 56700
rect 103190 56690 103310 56700
rect 103440 56690 103560 56700
rect 103690 56690 103810 56700
rect 103940 56690 104060 56700
rect 104190 56690 104310 56700
rect 104440 56690 104560 56700
rect 104690 56690 104810 56700
rect 104940 56690 105060 56700
rect 105190 56690 105310 56700
rect 105440 56690 105560 56700
rect 105690 56690 105810 56700
rect 105940 56690 106060 56700
rect 106190 56690 106310 56700
rect 106440 56690 106560 56700
rect 106690 56690 106810 56700
rect 106940 56690 107060 56700
rect 107190 56690 107310 56700
rect 107440 56690 107560 56700
rect 107690 56690 107810 56700
rect 107940 56690 108060 56700
rect 108190 56690 108310 56700
rect 108440 56690 108560 56700
rect 108690 56690 108810 56700
rect 108940 56690 109060 56700
rect 109190 56690 109310 56700
rect 109440 56690 109560 56700
rect 109690 56690 109810 56700
rect 109940 56690 110060 56700
rect 110190 56690 110310 56700
rect 110440 56690 110560 56700
rect 110690 56690 110810 56700
rect 110940 56690 111060 56700
rect 111190 56690 111310 56700
rect 111440 56690 111560 56700
rect 111690 56690 111810 56700
rect 111940 56690 112060 56700
rect 112190 56690 112310 56700
rect 112440 56690 112560 56700
rect 112690 56690 112810 56700
rect 112940 56690 113060 56700
rect 113190 56690 113310 56700
rect 113440 56690 113560 56700
rect 113690 56690 113810 56700
rect 113940 56690 114060 56700
rect 114190 56690 114310 56700
rect 114440 56690 114560 56700
rect 114690 56690 114810 56700
rect 114940 56690 115060 56700
rect 115190 56690 115310 56700
rect 115440 56690 115560 56700
rect 115690 56690 115810 56700
rect 115940 56690 116000 56700
rect 89000 56560 89050 56690
rect 89200 56560 89300 56690
rect 89450 56560 89550 56690
rect 89700 56560 89800 56690
rect 89950 56560 90050 56690
rect 90200 56560 90300 56690
rect 90450 56560 90550 56690
rect 90700 56560 90800 56690
rect 90950 56560 91050 56690
rect 91200 56560 91300 56690
rect 91450 56560 91550 56690
rect 91700 56560 91800 56690
rect 91950 56560 92050 56690
rect 92200 56560 92300 56690
rect 92450 56560 92550 56690
rect 92700 56560 92800 56690
rect 92950 56560 93050 56690
rect 93200 56560 93300 56690
rect 93450 56560 93550 56690
rect 93700 56560 93800 56690
rect 93950 56560 94050 56690
rect 94200 56560 94300 56690
rect 94450 56560 94550 56690
rect 94700 56560 94800 56690
rect 94950 56560 95050 56690
rect 95200 56560 95300 56690
rect 95450 56560 95550 56690
rect 95700 56560 95800 56690
rect 95950 56560 96050 56690
rect 96200 56560 96300 56690
rect 96450 56560 96550 56690
rect 96700 56560 96800 56690
rect 96950 56560 97050 56690
rect 97200 56560 97300 56690
rect 97450 56560 97550 56690
rect 97700 56560 97800 56690
rect 97950 56560 98050 56690
rect 98200 56560 98300 56690
rect 98450 56560 98550 56690
rect 98700 56560 98800 56690
rect 98950 56560 99050 56690
rect 99200 56560 99300 56690
rect 99450 56560 99550 56690
rect 99700 56560 99800 56690
rect 99950 56560 100050 56690
rect 100200 56560 100300 56690
rect 100450 56560 100550 56690
rect 100700 56560 100800 56690
rect 100950 56560 101050 56690
rect 101200 56560 101300 56690
rect 101450 56560 101550 56690
rect 101700 56560 101800 56690
rect 101950 56560 102050 56690
rect 102200 56560 102300 56690
rect 102450 56560 102550 56690
rect 102700 56560 102800 56690
rect 102950 56560 103050 56690
rect 103200 56560 103300 56690
rect 103450 56560 103550 56690
rect 103700 56560 103800 56690
rect 103950 56560 104050 56690
rect 104200 56560 104300 56690
rect 104450 56560 104550 56690
rect 104700 56560 104800 56690
rect 104950 56560 105050 56690
rect 105200 56560 105300 56690
rect 105450 56560 105550 56690
rect 105700 56560 105800 56690
rect 105950 56560 106050 56690
rect 106200 56560 106300 56690
rect 106450 56560 106550 56690
rect 106700 56560 106800 56690
rect 106950 56560 107050 56690
rect 107200 56560 107300 56690
rect 107450 56560 107550 56690
rect 107700 56560 107800 56690
rect 107950 56560 108050 56690
rect 108200 56560 108300 56690
rect 108450 56560 108550 56690
rect 108700 56560 108800 56690
rect 108950 56560 109050 56690
rect 109200 56560 109300 56690
rect 109450 56560 109550 56690
rect 109700 56560 109800 56690
rect 109950 56560 110050 56690
rect 110200 56560 110300 56690
rect 110450 56560 110550 56690
rect 110700 56560 110800 56690
rect 110950 56560 111050 56690
rect 111200 56560 111300 56690
rect 111450 56560 111550 56690
rect 111700 56560 111800 56690
rect 111950 56560 112050 56690
rect 112200 56560 112300 56690
rect 112450 56560 112550 56690
rect 112700 56560 112800 56690
rect 112950 56560 113050 56690
rect 113200 56560 113300 56690
rect 113450 56560 113550 56690
rect 113700 56560 113800 56690
rect 113950 56560 114050 56690
rect 114200 56560 114300 56690
rect 114450 56560 114550 56690
rect 114700 56560 114800 56690
rect 114950 56560 115050 56690
rect 115200 56560 115300 56690
rect 115450 56560 115550 56690
rect 115700 56560 115800 56690
rect 115950 56560 116000 56690
rect 89000 56550 89060 56560
rect 89190 56550 89310 56560
rect 89440 56550 89560 56560
rect 89690 56550 89810 56560
rect 89940 56550 90060 56560
rect 90190 56550 90310 56560
rect 90440 56550 90560 56560
rect 90690 56550 90810 56560
rect 90940 56550 91060 56560
rect 91190 56550 91310 56560
rect 91440 56550 91560 56560
rect 91690 56550 91810 56560
rect 91940 56550 92060 56560
rect 92190 56550 92310 56560
rect 92440 56550 92560 56560
rect 92690 56550 92810 56560
rect 92940 56550 93060 56560
rect 93190 56550 93310 56560
rect 93440 56550 93560 56560
rect 93690 56550 93810 56560
rect 93940 56550 94060 56560
rect 94190 56550 94310 56560
rect 94440 56550 94560 56560
rect 94690 56550 94810 56560
rect 94940 56550 95060 56560
rect 95190 56550 95310 56560
rect 95440 56550 95560 56560
rect 95690 56550 95810 56560
rect 95940 56550 96060 56560
rect 96190 56550 96310 56560
rect 96440 56550 96560 56560
rect 96690 56550 96810 56560
rect 96940 56550 97060 56560
rect 97190 56550 97310 56560
rect 97440 56550 97560 56560
rect 97690 56550 97810 56560
rect 97940 56550 98060 56560
rect 98190 56550 98310 56560
rect 98440 56550 98560 56560
rect 98690 56550 98810 56560
rect 98940 56550 99060 56560
rect 99190 56550 99310 56560
rect 99440 56550 99560 56560
rect 99690 56550 99810 56560
rect 99940 56550 100060 56560
rect 100190 56550 100310 56560
rect 100440 56550 100560 56560
rect 100690 56550 100810 56560
rect 100940 56550 101060 56560
rect 101190 56550 101310 56560
rect 101440 56550 101560 56560
rect 101690 56550 101810 56560
rect 101940 56550 102060 56560
rect 102190 56550 102310 56560
rect 102440 56550 102560 56560
rect 102690 56550 102810 56560
rect 102940 56550 103060 56560
rect 103190 56550 103310 56560
rect 103440 56550 103560 56560
rect 103690 56550 103810 56560
rect 103940 56550 104060 56560
rect 104190 56550 104310 56560
rect 104440 56550 104560 56560
rect 104690 56550 104810 56560
rect 104940 56550 105060 56560
rect 105190 56550 105310 56560
rect 105440 56550 105560 56560
rect 105690 56550 105810 56560
rect 105940 56550 106060 56560
rect 106190 56550 106310 56560
rect 106440 56550 106560 56560
rect 106690 56550 106810 56560
rect 106940 56550 107060 56560
rect 107190 56550 107310 56560
rect 107440 56550 107560 56560
rect 107690 56550 107810 56560
rect 107940 56550 108060 56560
rect 108190 56550 108310 56560
rect 108440 56550 108560 56560
rect 108690 56550 108810 56560
rect 108940 56550 109060 56560
rect 109190 56550 109310 56560
rect 109440 56550 109560 56560
rect 109690 56550 109810 56560
rect 109940 56550 110060 56560
rect 110190 56550 110310 56560
rect 110440 56550 110560 56560
rect 110690 56550 110810 56560
rect 110940 56550 111060 56560
rect 111190 56550 111310 56560
rect 111440 56550 111560 56560
rect 111690 56550 111810 56560
rect 111940 56550 112060 56560
rect 112190 56550 112310 56560
rect 112440 56550 112560 56560
rect 112690 56550 112810 56560
rect 112940 56550 113060 56560
rect 113190 56550 113310 56560
rect 113440 56550 113560 56560
rect 113690 56550 113810 56560
rect 113940 56550 114060 56560
rect 114190 56550 114310 56560
rect 114440 56550 114560 56560
rect 114690 56550 114810 56560
rect 114940 56550 115060 56560
rect 115190 56550 115310 56560
rect 115440 56550 115560 56560
rect 115690 56550 115810 56560
rect 115940 56550 116000 56560
rect 89000 56450 116000 56550
rect 89000 56440 89060 56450
rect 89190 56440 89310 56450
rect 89440 56440 89560 56450
rect 89690 56440 89810 56450
rect 89940 56440 90060 56450
rect 90190 56440 90310 56450
rect 90440 56440 90560 56450
rect 90690 56440 90810 56450
rect 90940 56440 91060 56450
rect 91190 56440 91310 56450
rect 91440 56440 91560 56450
rect 91690 56440 91810 56450
rect 91940 56440 92060 56450
rect 92190 56440 92310 56450
rect 92440 56440 92560 56450
rect 92690 56440 92810 56450
rect 92940 56440 93060 56450
rect 93190 56440 93310 56450
rect 93440 56440 93560 56450
rect 93690 56440 93810 56450
rect 93940 56440 94060 56450
rect 94190 56440 94310 56450
rect 94440 56440 94560 56450
rect 94690 56440 94810 56450
rect 94940 56440 95060 56450
rect 95190 56440 95310 56450
rect 95440 56440 95560 56450
rect 95690 56440 95810 56450
rect 95940 56440 96060 56450
rect 96190 56440 96310 56450
rect 96440 56440 96560 56450
rect 96690 56440 96810 56450
rect 96940 56440 97060 56450
rect 97190 56440 97310 56450
rect 97440 56440 97560 56450
rect 97690 56440 97810 56450
rect 97940 56440 98060 56450
rect 98190 56440 98310 56450
rect 98440 56440 98560 56450
rect 98690 56440 98810 56450
rect 98940 56440 99060 56450
rect 99190 56440 99310 56450
rect 99440 56440 99560 56450
rect 99690 56440 99810 56450
rect 99940 56440 100060 56450
rect 100190 56440 100310 56450
rect 100440 56440 100560 56450
rect 100690 56440 100810 56450
rect 100940 56440 101060 56450
rect 101190 56440 101310 56450
rect 101440 56440 101560 56450
rect 101690 56440 101810 56450
rect 101940 56440 102060 56450
rect 102190 56440 102310 56450
rect 102440 56440 102560 56450
rect 102690 56440 102810 56450
rect 102940 56440 103060 56450
rect 103190 56440 103310 56450
rect 103440 56440 103560 56450
rect 103690 56440 103810 56450
rect 103940 56440 104060 56450
rect 104190 56440 104310 56450
rect 104440 56440 104560 56450
rect 104690 56440 104810 56450
rect 104940 56440 105060 56450
rect 105190 56440 105310 56450
rect 105440 56440 105560 56450
rect 105690 56440 105810 56450
rect 105940 56440 106060 56450
rect 106190 56440 106310 56450
rect 106440 56440 106560 56450
rect 106690 56440 106810 56450
rect 106940 56440 107060 56450
rect 107190 56440 107310 56450
rect 107440 56440 107560 56450
rect 107690 56440 107810 56450
rect 107940 56440 108060 56450
rect 108190 56440 108310 56450
rect 108440 56440 108560 56450
rect 108690 56440 108810 56450
rect 108940 56440 109060 56450
rect 109190 56440 109310 56450
rect 109440 56440 109560 56450
rect 109690 56440 109810 56450
rect 109940 56440 110060 56450
rect 110190 56440 110310 56450
rect 110440 56440 110560 56450
rect 110690 56440 110810 56450
rect 110940 56440 111060 56450
rect 111190 56440 111310 56450
rect 111440 56440 111560 56450
rect 111690 56440 111810 56450
rect 111940 56440 112060 56450
rect 112190 56440 112310 56450
rect 112440 56440 112560 56450
rect 112690 56440 112810 56450
rect 112940 56440 113060 56450
rect 113190 56440 113310 56450
rect 113440 56440 113560 56450
rect 113690 56440 113810 56450
rect 113940 56440 114060 56450
rect 114190 56440 114310 56450
rect 114440 56440 114560 56450
rect 114690 56440 114810 56450
rect 114940 56440 115060 56450
rect 115190 56440 115310 56450
rect 115440 56440 115560 56450
rect 115690 56440 115810 56450
rect 115940 56440 116000 56450
rect 89000 56310 89050 56440
rect 89200 56310 89300 56440
rect 89450 56310 89550 56440
rect 89700 56310 89800 56440
rect 89950 56310 90050 56440
rect 90200 56310 90300 56440
rect 90450 56310 90550 56440
rect 90700 56310 90800 56440
rect 90950 56310 91050 56440
rect 91200 56310 91300 56440
rect 91450 56310 91550 56440
rect 91700 56310 91800 56440
rect 91950 56310 92050 56440
rect 92200 56310 92300 56440
rect 92450 56310 92550 56440
rect 92700 56310 92800 56440
rect 92950 56310 93050 56440
rect 93200 56310 93300 56440
rect 93450 56310 93550 56440
rect 93700 56310 93800 56440
rect 93950 56310 94050 56440
rect 94200 56310 94300 56440
rect 94450 56310 94550 56440
rect 94700 56310 94800 56440
rect 94950 56310 95050 56440
rect 95200 56310 95300 56440
rect 95450 56310 95550 56440
rect 95700 56310 95800 56440
rect 95950 56310 96050 56440
rect 96200 56310 96300 56440
rect 96450 56310 96550 56440
rect 96700 56310 96800 56440
rect 96950 56310 97050 56440
rect 97200 56310 97300 56440
rect 97450 56310 97550 56440
rect 97700 56310 97800 56440
rect 97950 56310 98050 56440
rect 98200 56310 98300 56440
rect 98450 56310 98550 56440
rect 98700 56310 98800 56440
rect 98950 56310 99050 56440
rect 99200 56310 99300 56440
rect 99450 56310 99550 56440
rect 99700 56310 99800 56440
rect 99950 56310 100050 56440
rect 100200 56310 100300 56440
rect 100450 56310 100550 56440
rect 100700 56310 100800 56440
rect 100950 56310 101050 56440
rect 101200 56310 101300 56440
rect 101450 56310 101550 56440
rect 101700 56310 101800 56440
rect 101950 56310 102050 56440
rect 102200 56310 102300 56440
rect 102450 56310 102550 56440
rect 102700 56310 102800 56440
rect 102950 56310 103050 56440
rect 103200 56310 103300 56440
rect 103450 56310 103550 56440
rect 103700 56310 103800 56440
rect 103950 56310 104050 56440
rect 104200 56310 104300 56440
rect 104450 56310 104550 56440
rect 104700 56310 104800 56440
rect 104950 56310 105050 56440
rect 105200 56310 105300 56440
rect 105450 56310 105550 56440
rect 105700 56310 105800 56440
rect 105950 56310 106050 56440
rect 106200 56310 106300 56440
rect 106450 56310 106550 56440
rect 106700 56310 106800 56440
rect 106950 56310 107050 56440
rect 107200 56310 107300 56440
rect 107450 56310 107550 56440
rect 107700 56310 107800 56440
rect 107950 56310 108050 56440
rect 108200 56310 108300 56440
rect 108450 56310 108550 56440
rect 108700 56310 108800 56440
rect 108950 56310 109050 56440
rect 109200 56310 109300 56440
rect 109450 56310 109550 56440
rect 109700 56310 109800 56440
rect 109950 56310 110050 56440
rect 110200 56310 110300 56440
rect 110450 56310 110550 56440
rect 110700 56310 110800 56440
rect 110950 56310 111050 56440
rect 111200 56310 111300 56440
rect 111450 56310 111550 56440
rect 111700 56310 111800 56440
rect 111950 56310 112050 56440
rect 112200 56310 112300 56440
rect 112450 56310 112550 56440
rect 112700 56310 112800 56440
rect 112950 56310 113050 56440
rect 113200 56310 113300 56440
rect 113450 56310 113550 56440
rect 113700 56310 113800 56440
rect 113950 56310 114050 56440
rect 114200 56310 114300 56440
rect 114450 56310 114550 56440
rect 114700 56310 114800 56440
rect 114950 56310 115050 56440
rect 115200 56310 115300 56440
rect 115450 56310 115550 56440
rect 115700 56310 115800 56440
rect 115950 56310 116000 56440
rect 89000 56300 89060 56310
rect 89190 56300 89310 56310
rect 89440 56300 89560 56310
rect 89690 56300 89810 56310
rect 89940 56300 90060 56310
rect 90190 56300 90310 56310
rect 90440 56300 90560 56310
rect 90690 56300 90810 56310
rect 90940 56300 91060 56310
rect 91190 56300 91310 56310
rect 91440 56300 91560 56310
rect 91690 56300 91810 56310
rect 91940 56300 92060 56310
rect 92190 56300 92310 56310
rect 92440 56300 92560 56310
rect 92690 56300 92810 56310
rect 92940 56300 93060 56310
rect 93190 56300 93310 56310
rect 93440 56300 93560 56310
rect 93690 56300 93810 56310
rect 93940 56300 94060 56310
rect 94190 56300 94310 56310
rect 94440 56300 94560 56310
rect 94690 56300 94810 56310
rect 94940 56300 95060 56310
rect 95190 56300 95310 56310
rect 95440 56300 95560 56310
rect 95690 56300 95810 56310
rect 95940 56300 96060 56310
rect 96190 56300 96310 56310
rect 96440 56300 96560 56310
rect 96690 56300 96810 56310
rect 96940 56300 97060 56310
rect 97190 56300 97310 56310
rect 97440 56300 97560 56310
rect 97690 56300 97810 56310
rect 97940 56300 98060 56310
rect 98190 56300 98310 56310
rect 98440 56300 98560 56310
rect 98690 56300 98810 56310
rect 98940 56300 99060 56310
rect 99190 56300 99310 56310
rect 99440 56300 99560 56310
rect 99690 56300 99810 56310
rect 99940 56300 100060 56310
rect 100190 56300 100310 56310
rect 100440 56300 100560 56310
rect 100690 56300 100810 56310
rect 100940 56300 101060 56310
rect 101190 56300 101310 56310
rect 101440 56300 101560 56310
rect 101690 56300 101810 56310
rect 101940 56300 102060 56310
rect 102190 56300 102310 56310
rect 102440 56300 102560 56310
rect 102690 56300 102810 56310
rect 102940 56300 103060 56310
rect 103190 56300 103310 56310
rect 103440 56300 103560 56310
rect 103690 56300 103810 56310
rect 103940 56300 104060 56310
rect 104190 56300 104310 56310
rect 104440 56300 104560 56310
rect 104690 56300 104810 56310
rect 104940 56300 105060 56310
rect 105190 56300 105310 56310
rect 105440 56300 105560 56310
rect 105690 56300 105810 56310
rect 105940 56300 106060 56310
rect 106190 56300 106310 56310
rect 106440 56300 106560 56310
rect 106690 56300 106810 56310
rect 106940 56300 107060 56310
rect 107190 56300 107310 56310
rect 107440 56300 107560 56310
rect 107690 56300 107810 56310
rect 107940 56300 108060 56310
rect 108190 56300 108310 56310
rect 108440 56300 108560 56310
rect 108690 56300 108810 56310
rect 108940 56300 109060 56310
rect 109190 56300 109310 56310
rect 109440 56300 109560 56310
rect 109690 56300 109810 56310
rect 109940 56300 110060 56310
rect 110190 56300 110310 56310
rect 110440 56300 110560 56310
rect 110690 56300 110810 56310
rect 110940 56300 111060 56310
rect 111190 56300 111310 56310
rect 111440 56300 111560 56310
rect 111690 56300 111810 56310
rect 111940 56300 112060 56310
rect 112190 56300 112310 56310
rect 112440 56300 112560 56310
rect 112690 56300 112810 56310
rect 112940 56300 113060 56310
rect 113190 56300 113310 56310
rect 113440 56300 113560 56310
rect 113690 56300 113810 56310
rect 113940 56300 114060 56310
rect 114190 56300 114310 56310
rect 114440 56300 114560 56310
rect 114690 56300 114810 56310
rect 114940 56300 115060 56310
rect 115190 56300 115310 56310
rect 115440 56300 115560 56310
rect 115690 56300 115810 56310
rect 115940 56300 116000 56310
rect 89000 56200 116000 56300
rect 89000 56190 89060 56200
rect 89190 56190 89310 56200
rect 89440 56190 89560 56200
rect 89690 56190 89810 56200
rect 89940 56190 90060 56200
rect 90190 56190 90310 56200
rect 90440 56190 90560 56200
rect 90690 56190 90810 56200
rect 90940 56190 91060 56200
rect 91190 56190 91310 56200
rect 91440 56190 91560 56200
rect 91690 56190 91810 56200
rect 91940 56190 92060 56200
rect 92190 56190 92310 56200
rect 92440 56190 92560 56200
rect 92690 56190 92810 56200
rect 92940 56190 93060 56200
rect 93190 56190 93310 56200
rect 93440 56190 93560 56200
rect 93690 56190 93810 56200
rect 93940 56190 94060 56200
rect 94190 56190 94310 56200
rect 94440 56190 94560 56200
rect 94690 56190 94810 56200
rect 94940 56190 95060 56200
rect 95190 56190 95310 56200
rect 95440 56190 95560 56200
rect 95690 56190 95810 56200
rect 95940 56190 96060 56200
rect 96190 56190 96310 56200
rect 96440 56190 96560 56200
rect 96690 56190 96810 56200
rect 96940 56190 97060 56200
rect 97190 56190 97310 56200
rect 97440 56190 97560 56200
rect 97690 56190 97810 56200
rect 97940 56190 98060 56200
rect 98190 56190 98310 56200
rect 98440 56190 98560 56200
rect 98690 56190 98810 56200
rect 98940 56190 99060 56200
rect 99190 56190 99310 56200
rect 99440 56190 99560 56200
rect 99690 56190 99810 56200
rect 99940 56190 100060 56200
rect 100190 56190 100310 56200
rect 100440 56190 100560 56200
rect 100690 56190 100810 56200
rect 100940 56190 101060 56200
rect 101190 56190 101310 56200
rect 101440 56190 101560 56200
rect 101690 56190 101810 56200
rect 101940 56190 102060 56200
rect 102190 56190 102310 56200
rect 102440 56190 102560 56200
rect 102690 56190 102810 56200
rect 102940 56190 103060 56200
rect 103190 56190 103310 56200
rect 103440 56190 103560 56200
rect 103690 56190 103810 56200
rect 103940 56190 104060 56200
rect 104190 56190 104310 56200
rect 104440 56190 104560 56200
rect 104690 56190 104810 56200
rect 104940 56190 105060 56200
rect 105190 56190 105310 56200
rect 105440 56190 105560 56200
rect 105690 56190 105810 56200
rect 105940 56190 106060 56200
rect 106190 56190 106310 56200
rect 106440 56190 106560 56200
rect 106690 56190 106810 56200
rect 106940 56190 107060 56200
rect 107190 56190 107310 56200
rect 107440 56190 107560 56200
rect 107690 56190 107810 56200
rect 107940 56190 108060 56200
rect 108190 56190 108310 56200
rect 108440 56190 108560 56200
rect 108690 56190 108810 56200
rect 108940 56190 109060 56200
rect 109190 56190 109310 56200
rect 109440 56190 109560 56200
rect 109690 56190 109810 56200
rect 109940 56190 110060 56200
rect 110190 56190 110310 56200
rect 110440 56190 110560 56200
rect 110690 56190 110810 56200
rect 110940 56190 111060 56200
rect 111190 56190 111310 56200
rect 111440 56190 111560 56200
rect 111690 56190 111810 56200
rect 111940 56190 112060 56200
rect 112190 56190 112310 56200
rect 112440 56190 112560 56200
rect 112690 56190 112810 56200
rect 112940 56190 113060 56200
rect 113190 56190 113310 56200
rect 113440 56190 113560 56200
rect 113690 56190 113810 56200
rect 113940 56190 114060 56200
rect 114190 56190 114310 56200
rect 114440 56190 114560 56200
rect 114690 56190 114810 56200
rect 114940 56190 115060 56200
rect 115190 56190 115310 56200
rect 115440 56190 115560 56200
rect 115690 56190 115810 56200
rect 115940 56190 116000 56200
rect 89000 56060 89050 56190
rect 89200 56060 89300 56190
rect 89450 56060 89550 56190
rect 89700 56060 89800 56190
rect 89950 56060 90050 56190
rect 90200 56060 90300 56190
rect 90450 56060 90550 56190
rect 90700 56060 90800 56190
rect 90950 56060 91050 56190
rect 91200 56060 91300 56190
rect 91450 56060 91550 56190
rect 91700 56060 91800 56190
rect 91950 56060 92050 56190
rect 92200 56060 92300 56190
rect 92450 56060 92550 56190
rect 92700 56060 92800 56190
rect 92950 56060 93050 56190
rect 93200 56060 93300 56190
rect 93450 56060 93550 56190
rect 93700 56060 93800 56190
rect 93950 56060 94050 56190
rect 94200 56060 94300 56190
rect 94450 56060 94550 56190
rect 94700 56060 94800 56190
rect 94950 56060 95050 56190
rect 95200 56060 95300 56190
rect 95450 56060 95550 56190
rect 95700 56060 95800 56190
rect 95950 56060 96050 56190
rect 96200 56060 96300 56190
rect 96450 56060 96550 56190
rect 96700 56060 96800 56190
rect 96950 56060 97050 56190
rect 97200 56060 97300 56190
rect 97450 56060 97550 56190
rect 97700 56060 97800 56190
rect 97950 56060 98050 56190
rect 98200 56060 98300 56190
rect 98450 56060 98550 56190
rect 98700 56060 98800 56190
rect 98950 56060 99050 56190
rect 99200 56060 99300 56190
rect 99450 56060 99550 56190
rect 99700 56060 99800 56190
rect 99950 56060 100050 56190
rect 100200 56060 100300 56190
rect 100450 56060 100550 56190
rect 100700 56060 100800 56190
rect 100950 56060 101050 56190
rect 101200 56060 101300 56190
rect 101450 56060 101550 56190
rect 101700 56060 101800 56190
rect 101950 56060 102050 56190
rect 102200 56060 102300 56190
rect 102450 56060 102550 56190
rect 102700 56060 102800 56190
rect 102950 56060 103050 56190
rect 103200 56060 103300 56190
rect 103450 56060 103550 56190
rect 103700 56060 103800 56190
rect 103950 56060 104050 56190
rect 104200 56060 104300 56190
rect 104450 56060 104550 56190
rect 104700 56060 104800 56190
rect 104950 56060 105050 56190
rect 105200 56060 105300 56190
rect 105450 56060 105550 56190
rect 105700 56060 105800 56190
rect 105950 56060 106050 56190
rect 106200 56060 106300 56190
rect 106450 56060 106550 56190
rect 106700 56060 106800 56190
rect 106950 56060 107050 56190
rect 107200 56060 107300 56190
rect 107450 56060 107550 56190
rect 107700 56060 107800 56190
rect 107950 56060 108050 56190
rect 108200 56060 108300 56190
rect 108450 56060 108550 56190
rect 108700 56060 108800 56190
rect 108950 56060 109050 56190
rect 109200 56060 109300 56190
rect 109450 56060 109550 56190
rect 109700 56060 109800 56190
rect 109950 56060 110050 56190
rect 110200 56060 110300 56190
rect 110450 56060 110550 56190
rect 110700 56060 110800 56190
rect 110950 56060 111050 56190
rect 111200 56060 111300 56190
rect 111450 56060 111550 56190
rect 111700 56060 111800 56190
rect 111950 56060 112050 56190
rect 112200 56060 112300 56190
rect 112450 56060 112550 56190
rect 112700 56060 112800 56190
rect 112950 56060 113050 56190
rect 113200 56060 113300 56190
rect 113450 56060 113550 56190
rect 113700 56060 113800 56190
rect 113950 56060 114050 56190
rect 114200 56060 114300 56190
rect 114450 56060 114550 56190
rect 114700 56060 114800 56190
rect 114950 56060 115050 56190
rect 115200 56060 115300 56190
rect 115450 56060 115550 56190
rect 115700 56060 115800 56190
rect 115950 56060 116000 56190
rect 89000 56050 89060 56060
rect 89190 56050 89310 56060
rect 89440 56050 89560 56060
rect 89690 56050 89810 56060
rect 89940 56050 90060 56060
rect 90190 56050 90310 56060
rect 90440 56050 90560 56060
rect 90690 56050 90810 56060
rect 90940 56050 91060 56060
rect 91190 56050 91310 56060
rect 91440 56050 91560 56060
rect 91690 56050 91810 56060
rect 91940 56050 92060 56060
rect 92190 56050 92310 56060
rect 92440 56050 92560 56060
rect 92690 56050 92810 56060
rect 92940 56050 93060 56060
rect 93190 56050 93310 56060
rect 93440 56050 93560 56060
rect 93690 56050 93810 56060
rect 93940 56050 94060 56060
rect 94190 56050 94310 56060
rect 94440 56050 94560 56060
rect 94690 56050 94810 56060
rect 94940 56050 95060 56060
rect 95190 56050 95310 56060
rect 95440 56050 95560 56060
rect 95690 56050 95810 56060
rect 95940 56050 96060 56060
rect 96190 56050 96310 56060
rect 96440 56050 96560 56060
rect 96690 56050 96810 56060
rect 96940 56050 97060 56060
rect 97190 56050 97310 56060
rect 97440 56050 97560 56060
rect 97690 56050 97810 56060
rect 97940 56050 98060 56060
rect 98190 56050 98310 56060
rect 98440 56050 98560 56060
rect 98690 56050 98810 56060
rect 98940 56050 99060 56060
rect 99190 56050 99310 56060
rect 99440 56050 99560 56060
rect 99690 56050 99810 56060
rect 99940 56050 100060 56060
rect 100190 56050 100310 56060
rect 100440 56050 100560 56060
rect 100690 56050 100810 56060
rect 100940 56050 101060 56060
rect 101190 56050 101310 56060
rect 101440 56050 101560 56060
rect 101690 56050 101810 56060
rect 101940 56050 102060 56060
rect 102190 56050 102310 56060
rect 102440 56050 102560 56060
rect 102690 56050 102810 56060
rect 102940 56050 103060 56060
rect 103190 56050 103310 56060
rect 103440 56050 103560 56060
rect 103690 56050 103810 56060
rect 103940 56050 104060 56060
rect 104190 56050 104310 56060
rect 104440 56050 104560 56060
rect 104690 56050 104810 56060
rect 104940 56050 105060 56060
rect 105190 56050 105310 56060
rect 105440 56050 105560 56060
rect 105690 56050 105810 56060
rect 105940 56050 106060 56060
rect 106190 56050 106310 56060
rect 106440 56050 106560 56060
rect 106690 56050 106810 56060
rect 106940 56050 107060 56060
rect 107190 56050 107310 56060
rect 107440 56050 107560 56060
rect 107690 56050 107810 56060
rect 107940 56050 108060 56060
rect 108190 56050 108310 56060
rect 108440 56050 108560 56060
rect 108690 56050 108810 56060
rect 108940 56050 109060 56060
rect 109190 56050 109310 56060
rect 109440 56050 109560 56060
rect 109690 56050 109810 56060
rect 109940 56050 110060 56060
rect 110190 56050 110310 56060
rect 110440 56050 110560 56060
rect 110690 56050 110810 56060
rect 110940 56050 111060 56060
rect 111190 56050 111310 56060
rect 111440 56050 111560 56060
rect 111690 56050 111810 56060
rect 111940 56050 112060 56060
rect 112190 56050 112310 56060
rect 112440 56050 112560 56060
rect 112690 56050 112810 56060
rect 112940 56050 113060 56060
rect 113190 56050 113310 56060
rect 113440 56050 113560 56060
rect 113690 56050 113810 56060
rect 113940 56050 114060 56060
rect 114190 56050 114310 56060
rect 114440 56050 114560 56060
rect 114690 56050 114810 56060
rect 114940 56050 115060 56060
rect 115190 56050 115310 56060
rect 115440 56050 115560 56060
rect 115690 56050 115810 56060
rect 115940 56050 116000 56060
rect 89000 55950 116000 56050
rect 89000 55940 89060 55950
rect 89190 55940 89310 55950
rect 89440 55940 89560 55950
rect 89690 55940 89810 55950
rect 89940 55940 90060 55950
rect 90190 55940 90310 55950
rect 90440 55940 90560 55950
rect 90690 55940 90810 55950
rect 90940 55940 91060 55950
rect 91190 55940 91310 55950
rect 91440 55940 91560 55950
rect 91690 55940 91810 55950
rect 91940 55940 92060 55950
rect 92190 55940 92310 55950
rect 92440 55940 92560 55950
rect 92690 55940 92810 55950
rect 92940 55940 93060 55950
rect 93190 55940 93310 55950
rect 93440 55940 93560 55950
rect 93690 55940 93810 55950
rect 93940 55940 94060 55950
rect 94190 55940 94310 55950
rect 94440 55940 94560 55950
rect 94690 55940 94810 55950
rect 94940 55940 95060 55950
rect 95190 55940 95310 55950
rect 95440 55940 95560 55950
rect 95690 55940 95810 55950
rect 95940 55940 96060 55950
rect 96190 55940 96310 55950
rect 96440 55940 96560 55950
rect 96690 55940 96810 55950
rect 96940 55940 97060 55950
rect 97190 55940 97310 55950
rect 97440 55940 97560 55950
rect 97690 55940 97810 55950
rect 97940 55940 98060 55950
rect 98190 55940 98310 55950
rect 98440 55940 98560 55950
rect 98690 55940 98810 55950
rect 98940 55940 99060 55950
rect 99190 55940 99310 55950
rect 99440 55940 99560 55950
rect 99690 55940 99810 55950
rect 99940 55940 100060 55950
rect 100190 55940 100310 55950
rect 100440 55940 100560 55950
rect 100690 55940 100810 55950
rect 100940 55940 101060 55950
rect 101190 55940 101310 55950
rect 101440 55940 101560 55950
rect 101690 55940 101810 55950
rect 101940 55940 102060 55950
rect 102190 55940 102310 55950
rect 102440 55940 102560 55950
rect 102690 55940 102810 55950
rect 102940 55940 103060 55950
rect 103190 55940 103310 55950
rect 103440 55940 103560 55950
rect 103690 55940 103810 55950
rect 103940 55940 104060 55950
rect 104190 55940 104310 55950
rect 104440 55940 104560 55950
rect 104690 55940 104810 55950
rect 104940 55940 105060 55950
rect 105190 55940 105310 55950
rect 105440 55940 105560 55950
rect 105690 55940 105810 55950
rect 105940 55940 106060 55950
rect 106190 55940 106310 55950
rect 106440 55940 106560 55950
rect 106690 55940 106810 55950
rect 106940 55940 107060 55950
rect 107190 55940 107310 55950
rect 107440 55940 107560 55950
rect 107690 55940 107810 55950
rect 107940 55940 108060 55950
rect 108190 55940 108310 55950
rect 108440 55940 108560 55950
rect 108690 55940 108810 55950
rect 108940 55940 109060 55950
rect 109190 55940 109310 55950
rect 109440 55940 109560 55950
rect 109690 55940 109810 55950
rect 109940 55940 110060 55950
rect 110190 55940 110310 55950
rect 110440 55940 110560 55950
rect 110690 55940 110810 55950
rect 110940 55940 111060 55950
rect 111190 55940 111310 55950
rect 111440 55940 111560 55950
rect 111690 55940 111810 55950
rect 111940 55940 112060 55950
rect 112190 55940 112310 55950
rect 112440 55940 112560 55950
rect 112690 55940 112810 55950
rect 112940 55940 113060 55950
rect 113190 55940 113310 55950
rect 113440 55940 113560 55950
rect 113690 55940 113810 55950
rect 113940 55940 114060 55950
rect 114190 55940 114310 55950
rect 114440 55940 114560 55950
rect 114690 55940 114810 55950
rect 114940 55940 115060 55950
rect 115190 55940 115310 55950
rect 115440 55940 115560 55950
rect 115690 55940 115810 55950
rect 115940 55940 116000 55950
rect 89000 55810 89050 55940
rect 89200 55810 89300 55940
rect 89450 55810 89550 55940
rect 89700 55810 89800 55940
rect 89950 55810 90050 55940
rect 90200 55810 90300 55940
rect 90450 55810 90550 55940
rect 90700 55810 90800 55940
rect 90950 55810 91050 55940
rect 91200 55810 91300 55940
rect 91450 55810 91550 55940
rect 91700 55810 91800 55940
rect 91950 55810 92050 55940
rect 92200 55810 92300 55940
rect 92450 55810 92550 55940
rect 92700 55810 92800 55940
rect 92950 55810 93050 55940
rect 93200 55810 93300 55940
rect 93450 55810 93550 55940
rect 93700 55810 93800 55940
rect 93950 55810 94050 55940
rect 94200 55810 94300 55940
rect 94450 55810 94550 55940
rect 94700 55810 94800 55940
rect 94950 55810 95050 55940
rect 95200 55810 95300 55940
rect 95450 55810 95550 55940
rect 95700 55810 95800 55940
rect 95950 55810 96050 55940
rect 96200 55810 96300 55940
rect 96450 55810 96550 55940
rect 96700 55810 96800 55940
rect 96950 55810 97050 55940
rect 97200 55810 97300 55940
rect 97450 55810 97550 55940
rect 97700 55810 97800 55940
rect 97950 55810 98050 55940
rect 98200 55810 98300 55940
rect 98450 55810 98550 55940
rect 98700 55810 98800 55940
rect 98950 55810 99050 55940
rect 99200 55810 99300 55940
rect 99450 55810 99550 55940
rect 99700 55810 99800 55940
rect 99950 55810 100050 55940
rect 100200 55810 100300 55940
rect 100450 55810 100550 55940
rect 100700 55810 100800 55940
rect 100950 55810 101050 55940
rect 101200 55810 101300 55940
rect 101450 55810 101550 55940
rect 101700 55810 101800 55940
rect 101950 55810 102050 55940
rect 102200 55810 102300 55940
rect 102450 55810 102550 55940
rect 102700 55810 102800 55940
rect 102950 55810 103050 55940
rect 103200 55810 103300 55940
rect 103450 55810 103550 55940
rect 103700 55810 103800 55940
rect 103950 55810 104050 55940
rect 104200 55810 104300 55940
rect 104450 55810 104550 55940
rect 104700 55810 104800 55940
rect 104950 55810 105050 55940
rect 105200 55810 105300 55940
rect 105450 55810 105550 55940
rect 105700 55810 105800 55940
rect 105950 55810 106050 55940
rect 106200 55810 106300 55940
rect 106450 55810 106550 55940
rect 106700 55810 106800 55940
rect 106950 55810 107050 55940
rect 107200 55810 107300 55940
rect 107450 55810 107550 55940
rect 107700 55810 107800 55940
rect 107950 55810 108050 55940
rect 108200 55810 108300 55940
rect 108450 55810 108550 55940
rect 108700 55810 108800 55940
rect 108950 55810 109050 55940
rect 109200 55810 109300 55940
rect 109450 55810 109550 55940
rect 109700 55810 109800 55940
rect 109950 55810 110050 55940
rect 110200 55810 110300 55940
rect 110450 55810 110550 55940
rect 110700 55810 110800 55940
rect 110950 55810 111050 55940
rect 111200 55810 111300 55940
rect 111450 55810 111550 55940
rect 111700 55810 111800 55940
rect 111950 55810 112050 55940
rect 112200 55810 112300 55940
rect 112450 55810 112550 55940
rect 112700 55810 112800 55940
rect 112950 55810 113050 55940
rect 113200 55810 113300 55940
rect 113450 55810 113550 55940
rect 113700 55810 113800 55940
rect 113950 55810 114050 55940
rect 114200 55810 114300 55940
rect 114450 55810 114550 55940
rect 114700 55810 114800 55940
rect 114950 55810 115050 55940
rect 115200 55810 115300 55940
rect 115450 55810 115550 55940
rect 115700 55810 115800 55940
rect 115950 55810 116000 55940
rect 89000 55800 89060 55810
rect 89190 55800 89310 55810
rect 89440 55800 89560 55810
rect 89690 55800 89810 55810
rect 89940 55800 90060 55810
rect 90190 55800 90310 55810
rect 90440 55800 90560 55810
rect 90690 55800 90810 55810
rect 90940 55800 91060 55810
rect 91190 55800 91310 55810
rect 91440 55800 91560 55810
rect 91690 55800 91810 55810
rect 91940 55800 92060 55810
rect 92190 55800 92310 55810
rect 92440 55800 92560 55810
rect 92690 55800 92810 55810
rect 92940 55800 93060 55810
rect 93190 55800 93310 55810
rect 93440 55800 93560 55810
rect 93690 55800 93810 55810
rect 93940 55800 94060 55810
rect 94190 55800 94310 55810
rect 94440 55800 94560 55810
rect 94690 55800 94810 55810
rect 94940 55800 95060 55810
rect 95190 55800 95310 55810
rect 95440 55800 95560 55810
rect 95690 55800 95810 55810
rect 95940 55800 96060 55810
rect 96190 55800 96310 55810
rect 96440 55800 96560 55810
rect 96690 55800 96810 55810
rect 96940 55800 97060 55810
rect 97190 55800 97310 55810
rect 97440 55800 97560 55810
rect 97690 55800 97810 55810
rect 97940 55800 98060 55810
rect 98190 55800 98310 55810
rect 98440 55800 98560 55810
rect 98690 55800 98810 55810
rect 98940 55800 99060 55810
rect 99190 55800 99310 55810
rect 99440 55800 99560 55810
rect 99690 55800 99810 55810
rect 99940 55800 100060 55810
rect 100190 55800 100310 55810
rect 100440 55800 100560 55810
rect 100690 55800 100810 55810
rect 100940 55800 101060 55810
rect 101190 55800 101310 55810
rect 101440 55800 101560 55810
rect 101690 55800 101810 55810
rect 101940 55800 102060 55810
rect 102190 55800 102310 55810
rect 102440 55800 102560 55810
rect 102690 55800 102810 55810
rect 102940 55800 103060 55810
rect 103190 55800 103310 55810
rect 103440 55800 103560 55810
rect 103690 55800 103810 55810
rect 103940 55800 104060 55810
rect 104190 55800 104310 55810
rect 104440 55800 104560 55810
rect 104690 55800 104810 55810
rect 104940 55800 105060 55810
rect 105190 55800 105310 55810
rect 105440 55800 105560 55810
rect 105690 55800 105810 55810
rect 105940 55800 106060 55810
rect 106190 55800 106310 55810
rect 106440 55800 106560 55810
rect 106690 55800 106810 55810
rect 106940 55800 107060 55810
rect 107190 55800 107310 55810
rect 107440 55800 107560 55810
rect 107690 55800 107810 55810
rect 107940 55800 108060 55810
rect 108190 55800 108310 55810
rect 108440 55800 108560 55810
rect 108690 55800 108810 55810
rect 108940 55800 109060 55810
rect 109190 55800 109310 55810
rect 109440 55800 109560 55810
rect 109690 55800 109810 55810
rect 109940 55800 110060 55810
rect 110190 55800 110310 55810
rect 110440 55800 110560 55810
rect 110690 55800 110810 55810
rect 110940 55800 111060 55810
rect 111190 55800 111310 55810
rect 111440 55800 111560 55810
rect 111690 55800 111810 55810
rect 111940 55800 112060 55810
rect 112190 55800 112310 55810
rect 112440 55800 112560 55810
rect 112690 55800 112810 55810
rect 112940 55800 113060 55810
rect 113190 55800 113310 55810
rect 113440 55800 113560 55810
rect 113690 55800 113810 55810
rect 113940 55800 114060 55810
rect 114190 55800 114310 55810
rect 114440 55800 114560 55810
rect 114690 55800 114810 55810
rect 114940 55800 115060 55810
rect 115190 55800 115310 55810
rect 115440 55800 115560 55810
rect 115690 55800 115810 55810
rect 115940 55800 116000 55810
rect 89000 55700 116000 55800
rect 89000 55690 89060 55700
rect 89190 55690 89310 55700
rect 89440 55690 89560 55700
rect 89690 55690 89810 55700
rect 89940 55690 90060 55700
rect 90190 55690 90310 55700
rect 90440 55690 90560 55700
rect 90690 55690 90810 55700
rect 90940 55690 91060 55700
rect 91190 55690 91310 55700
rect 91440 55690 91560 55700
rect 91690 55690 91810 55700
rect 91940 55690 92060 55700
rect 92190 55690 92310 55700
rect 92440 55690 92560 55700
rect 92690 55690 92810 55700
rect 92940 55690 93060 55700
rect 93190 55690 93310 55700
rect 93440 55690 93560 55700
rect 93690 55690 93810 55700
rect 93940 55690 94060 55700
rect 94190 55690 94310 55700
rect 94440 55690 94560 55700
rect 94690 55690 94810 55700
rect 94940 55690 95060 55700
rect 95190 55690 95310 55700
rect 95440 55690 95560 55700
rect 95690 55690 95810 55700
rect 95940 55690 96060 55700
rect 96190 55690 96310 55700
rect 96440 55690 96560 55700
rect 96690 55690 96810 55700
rect 96940 55690 97060 55700
rect 97190 55690 97310 55700
rect 97440 55690 97560 55700
rect 97690 55690 97810 55700
rect 97940 55690 98060 55700
rect 98190 55690 98310 55700
rect 98440 55690 98560 55700
rect 98690 55690 98810 55700
rect 98940 55690 99060 55700
rect 99190 55690 99310 55700
rect 99440 55690 99560 55700
rect 99690 55690 99810 55700
rect 99940 55690 100060 55700
rect 100190 55690 100310 55700
rect 100440 55690 100560 55700
rect 100690 55690 100810 55700
rect 100940 55690 101060 55700
rect 101190 55690 101310 55700
rect 101440 55690 101560 55700
rect 101690 55690 101810 55700
rect 101940 55690 102060 55700
rect 102190 55690 102310 55700
rect 102440 55690 102560 55700
rect 102690 55690 102810 55700
rect 102940 55690 103060 55700
rect 103190 55690 103310 55700
rect 103440 55690 103560 55700
rect 103690 55690 103810 55700
rect 103940 55690 104060 55700
rect 104190 55690 104310 55700
rect 104440 55690 104560 55700
rect 104690 55690 104810 55700
rect 104940 55690 105060 55700
rect 105190 55690 105310 55700
rect 105440 55690 105560 55700
rect 105690 55690 105810 55700
rect 105940 55690 106060 55700
rect 106190 55690 106310 55700
rect 106440 55690 106560 55700
rect 106690 55690 106810 55700
rect 106940 55690 107060 55700
rect 107190 55690 107310 55700
rect 107440 55690 107560 55700
rect 107690 55690 107810 55700
rect 107940 55690 108060 55700
rect 108190 55690 108310 55700
rect 108440 55690 108560 55700
rect 108690 55690 108810 55700
rect 108940 55690 109060 55700
rect 109190 55690 109310 55700
rect 109440 55690 109560 55700
rect 109690 55690 109810 55700
rect 109940 55690 110060 55700
rect 110190 55690 110310 55700
rect 110440 55690 110560 55700
rect 110690 55690 110810 55700
rect 110940 55690 111060 55700
rect 111190 55690 111310 55700
rect 111440 55690 111560 55700
rect 111690 55690 111810 55700
rect 111940 55690 112060 55700
rect 112190 55690 112310 55700
rect 112440 55690 112560 55700
rect 112690 55690 112810 55700
rect 112940 55690 113060 55700
rect 113190 55690 113310 55700
rect 113440 55690 113560 55700
rect 113690 55690 113810 55700
rect 113940 55690 114060 55700
rect 114190 55690 114310 55700
rect 114440 55690 114560 55700
rect 114690 55690 114810 55700
rect 114940 55690 115060 55700
rect 115190 55690 115310 55700
rect 115440 55690 115560 55700
rect 115690 55690 115810 55700
rect 115940 55690 116000 55700
rect 89000 55560 89050 55690
rect 89200 55560 89300 55690
rect 89450 55560 89550 55690
rect 89700 55560 89800 55690
rect 89950 55560 90050 55690
rect 90200 55560 90300 55690
rect 90450 55560 90550 55690
rect 90700 55560 90800 55690
rect 90950 55560 91050 55690
rect 91200 55560 91300 55690
rect 91450 55560 91550 55690
rect 91700 55560 91800 55690
rect 91950 55560 92050 55690
rect 92200 55560 92300 55690
rect 92450 55560 92550 55690
rect 92700 55560 92800 55690
rect 92950 55560 93050 55690
rect 93200 55560 93300 55690
rect 93450 55560 93550 55690
rect 93700 55560 93800 55690
rect 93950 55560 94050 55690
rect 94200 55560 94300 55690
rect 94450 55560 94550 55690
rect 94700 55560 94800 55690
rect 94950 55560 95050 55690
rect 95200 55560 95300 55690
rect 95450 55560 95550 55690
rect 95700 55560 95800 55690
rect 95950 55560 96050 55690
rect 96200 55560 96300 55690
rect 96450 55560 96550 55690
rect 96700 55560 96800 55690
rect 96950 55560 97050 55690
rect 97200 55560 97300 55690
rect 97450 55560 97550 55690
rect 97700 55560 97800 55690
rect 97950 55560 98050 55690
rect 98200 55560 98300 55690
rect 98450 55560 98550 55690
rect 98700 55560 98800 55690
rect 98950 55560 99050 55690
rect 99200 55560 99300 55690
rect 99450 55560 99550 55690
rect 99700 55560 99800 55690
rect 99950 55560 100050 55690
rect 100200 55560 100300 55690
rect 100450 55560 100550 55690
rect 100700 55560 100800 55690
rect 100950 55560 101050 55690
rect 101200 55560 101300 55690
rect 101450 55560 101550 55690
rect 101700 55560 101800 55690
rect 101950 55560 102050 55690
rect 102200 55560 102300 55690
rect 102450 55560 102550 55690
rect 102700 55560 102800 55690
rect 102950 55560 103050 55690
rect 103200 55560 103300 55690
rect 103450 55560 103550 55690
rect 103700 55560 103800 55690
rect 103950 55560 104050 55690
rect 104200 55560 104300 55690
rect 104450 55560 104550 55690
rect 104700 55560 104800 55690
rect 104950 55560 105050 55690
rect 105200 55560 105300 55690
rect 105450 55560 105550 55690
rect 105700 55560 105800 55690
rect 105950 55560 106050 55690
rect 106200 55560 106300 55690
rect 106450 55560 106550 55690
rect 106700 55560 106800 55690
rect 106950 55560 107050 55690
rect 107200 55560 107300 55690
rect 107450 55560 107550 55690
rect 107700 55560 107800 55690
rect 107950 55560 108050 55690
rect 108200 55560 108300 55690
rect 108450 55560 108550 55690
rect 108700 55560 108800 55690
rect 108950 55560 109050 55690
rect 109200 55560 109300 55690
rect 109450 55560 109550 55690
rect 109700 55560 109800 55690
rect 109950 55560 110050 55690
rect 110200 55560 110300 55690
rect 110450 55560 110550 55690
rect 110700 55560 110800 55690
rect 110950 55560 111050 55690
rect 111200 55560 111300 55690
rect 111450 55560 111550 55690
rect 111700 55560 111800 55690
rect 111950 55560 112050 55690
rect 112200 55560 112300 55690
rect 112450 55560 112550 55690
rect 112700 55560 112800 55690
rect 112950 55560 113050 55690
rect 113200 55560 113300 55690
rect 113450 55560 113550 55690
rect 113700 55560 113800 55690
rect 113950 55560 114050 55690
rect 114200 55560 114300 55690
rect 114450 55560 114550 55690
rect 114700 55560 114800 55690
rect 114950 55560 115050 55690
rect 115200 55560 115300 55690
rect 115450 55560 115550 55690
rect 115700 55560 115800 55690
rect 115950 55560 116000 55690
rect 89000 55550 89060 55560
rect 89190 55550 89310 55560
rect 89440 55550 89560 55560
rect 89690 55550 89810 55560
rect 89940 55550 90060 55560
rect 90190 55550 90310 55560
rect 90440 55550 90560 55560
rect 90690 55550 90810 55560
rect 90940 55550 91060 55560
rect 91190 55550 91310 55560
rect 91440 55550 91560 55560
rect 91690 55550 91810 55560
rect 91940 55550 92060 55560
rect 92190 55550 92310 55560
rect 92440 55550 92560 55560
rect 92690 55550 92810 55560
rect 92940 55550 93060 55560
rect 93190 55550 93310 55560
rect 93440 55550 93560 55560
rect 93690 55550 93810 55560
rect 93940 55550 94060 55560
rect 94190 55550 94310 55560
rect 94440 55550 94560 55560
rect 94690 55550 94810 55560
rect 94940 55550 95060 55560
rect 95190 55550 95310 55560
rect 95440 55550 95560 55560
rect 95690 55550 95810 55560
rect 95940 55550 96060 55560
rect 96190 55550 96310 55560
rect 96440 55550 96560 55560
rect 96690 55550 96810 55560
rect 96940 55550 97060 55560
rect 97190 55550 97310 55560
rect 97440 55550 97560 55560
rect 97690 55550 97810 55560
rect 97940 55550 98060 55560
rect 98190 55550 98310 55560
rect 98440 55550 98560 55560
rect 98690 55550 98810 55560
rect 98940 55550 99060 55560
rect 99190 55550 99310 55560
rect 99440 55550 99560 55560
rect 99690 55550 99810 55560
rect 99940 55550 100060 55560
rect 100190 55550 100310 55560
rect 100440 55550 100560 55560
rect 100690 55550 100810 55560
rect 100940 55550 101060 55560
rect 101190 55550 101310 55560
rect 101440 55550 101560 55560
rect 101690 55550 101810 55560
rect 101940 55550 102060 55560
rect 102190 55550 102310 55560
rect 102440 55550 102560 55560
rect 102690 55550 102810 55560
rect 102940 55550 103060 55560
rect 103190 55550 103310 55560
rect 103440 55550 103560 55560
rect 103690 55550 103810 55560
rect 103940 55550 104060 55560
rect 104190 55550 104310 55560
rect 104440 55550 104560 55560
rect 104690 55550 104810 55560
rect 104940 55550 105060 55560
rect 105190 55550 105310 55560
rect 105440 55550 105560 55560
rect 105690 55550 105810 55560
rect 105940 55550 106060 55560
rect 106190 55550 106310 55560
rect 106440 55550 106560 55560
rect 106690 55550 106810 55560
rect 106940 55550 107060 55560
rect 107190 55550 107310 55560
rect 107440 55550 107560 55560
rect 107690 55550 107810 55560
rect 107940 55550 108060 55560
rect 108190 55550 108310 55560
rect 108440 55550 108560 55560
rect 108690 55550 108810 55560
rect 108940 55550 109060 55560
rect 109190 55550 109310 55560
rect 109440 55550 109560 55560
rect 109690 55550 109810 55560
rect 109940 55550 110060 55560
rect 110190 55550 110310 55560
rect 110440 55550 110560 55560
rect 110690 55550 110810 55560
rect 110940 55550 111060 55560
rect 111190 55550 111310 55560
rect 111440 55550 111560 55560
rect 111690 55550 111810 55560
rect 111940 55550 112060 55560
rect 112190 55550 112310 55560
rect 112440 55550 112560 55560
rect 112690 55550 112810 55560
rect 112940 55550 113060 55560
rect 113190 55550 113310 55560
rect 113440 55550 113560 55560
rect 113690 55550 113810 55560
rect 113940 55550 114060 55560
rect 114190 55550 114310 55560
rect 114440 55550 114560 55560
rect 114690 55550 114810 55560
rect 114940 55550 115060 55560
rect 115190 55550 115310 55560
rect 115440 55550 115560 55560
rect 115690 55550 115810 55560
rect 115940 55550 116000 55560
rect 89000 55450 116000 55550
rect 89000 55440 89060 55450
rect 89190 55440 89310 55450
rect 89440 55440 89560 55450
rect 89690 55440 89810 55450
rect 89940 55440 90060 55450
rect 90190 55440 90310 55450
rect 90440 55440 90560 55450
rect 90690 55440 90810 55450
rect 90940 55440 91060 55450
rect 91190 55440 91310 55450
rect 91440 55440 91560 55450
rect 91690 55440 91810 55450
rect 91940 55440 92060 55450
rect 92190 55440 92310 55450
rect 92440 55440 92560 55450
rect 92690 55440 92810 55450
rect 92940 55440 93060 55450
rect 93190 55440 93310 55450
rect 93440 55440 93560 55450
rect 93690 55440 93810 55450
rect 93940 55440 94060 55450
rect 94190 55440 94310 55450
rect 94440 55440 94560 55450
rect 94690 55440 94810 55450
rect 94940 55440 95060 55450
rect 95190 55440 95310 55450
rect 95440 55440 95560 55450
rect 95690 55440 95810 55450
rect 95940 55440 96060 55450
rect 96190 55440 96310 55450
rect 96440 55440 96560 55450
rect 96690 55440 96810 55450
rect 96940 55440 97060 55450
rect 97190 55440 97310 55450
rect 97440 55440 97560 55450
rect 97690 55440 97810 55450
rect 97940 55440 98060 55450
rect 98190 55440 98310 55450
rect 98440 55440 98560 55450
rect 98690 55440 98810 55450
rect 98940 55440 99060 55450
rect 99190 55440 99310 55450
rect 99440 55440 99560 55450
rect 99690 55440 99810 55450
rect 99940 55440 100060 55450
rect 100190 55440 100310 55450
rect 100440 55440 100560 55450
rect 100690 55440 100810 55450
rect 100940 55440 101060 55450
rect 101190 55440 101310 55450
rect 101440 55440 101560 55450
rect 101690 55440 101810 55450
rect 101940 55440 102060 55450
rect 102190 55440 102310 55450
rect 102440 55440 102560 55450
rect 102690 55440 102810 55450
rect 102940 55440 103060 55450
rect 103190 55440 103310 55450
rect 103440 55440 103560 55450
rect 103690 55440 103810 55450
rect 103940 55440 104060 55450
rect 104190 55440 104310 55450
rect 104440 55440 104560 55450
rect 104690 55440 104810 55450
rect 104940 55440 105060 55450
rect 105190 55440 105310 55450
rect 105440 55440 105560 55450
rect 105690 55440 105810 55450
rect 105940 55440 106060 55450
rect 106190 55440 106310 55450
rect 106440 55440 106560 55450
rect 106690 55440 106810 55450
rect 106940 55440 107060 55450
rect 107190 55440 107310 55450
rect 107440 55440 107560 55450
rect 107690 55440 107810 55450
rect 107940 55440 108060 55450
rect 108190 55440 108310 55450
rect 108440 55440 108560 55450
rect 108690 55440 108810 55450
rect 108940 55440 109060 55450
rect 109190 55440 109310 55450
rect 109440 55440 109560 55450
rect 109690 55440 109810 55450
rect 109940 55440 110060 55450
rect 110190 55440 110310 55450
rect 110440 55440 110560 55450
rect 110690 55440 110810 55450
rect 110940 55440 111060 55450
rect 111190 55440 111310 55450
rect 111440 55440 111560 55450
rect 111690 55440 111810 55450
rect 111940 55440 112060 55450
rect 112190 55440 112310 55450
rect 112440 55440 112560 55450
rect 112690 55440 112810 55450
rect 112940 55440 113060 55450
rect 113190 55440 113310 55450
rect 113440 55440 113560 55450
rect 113690 55440 113810 55450
rect 113940 55440 114060 55450
rect 114190 55440 114310 55450
rect 114440 55440 114560 55450
rect 114690 55440 114810 55450
rect 114940 55440 115060 55450
rect 115190 55440 115310 55450
rect 115440 55440 115560 55450
rect 115690 55440 115810 55450
rect 115940 55440 116000 55450
rect 89000 55310 89050 55440
rect 89200 55310 89300 55440
rect 89450 55310 89550 55440
rect 89700 55310 89800 55440
rect 89950 55310 90050 55440
rect 90200 55310 90300 55440
rect 90450 55310 90550 55440
rect 90700 55310 90800 55440
rect 90950 55310 91050 55440
rect 91200 55310 91300 55440
rect 91450 55310 91550 55440
rect 91700 55310 91800 55440
rect 91950 55310 92050 55440
rect 92200 55310 92300 55440
rect 92450 55310 92550 55440
rect 92700 55310 92800 55440
rect 92950 55310 93050 55440
rect 93200 55310 93300 55440
rect 93450 55310 93550 55440
rect 93700 55310 93800 55440
rect 93950 55310 94050 55440
rect 94200 55310 94300 55440
rect 94450 55310 94550 55440
rect 94700 55310 94800 55440
rect 94950 55310 95050 55440
rect 95200 55310 95300 55440
rect 95450 55310 95550 55440
rect 95700 55310 95800 55440
rect 95950 55310 96050 55440
rect 96200 55310 96300 55440
rect 96450 55310 96550 55440
rect 96700 55310 96800 55440
rect 96950 55310 97050 55440
rect 97200 55310 97300 55440
rect 97450 55310 97550 55440
rect 97700 55310 97800 55440
rect 97950 55310 98050 55440
rect 98200 55310 98300 55440
rect 98450 55310 98550 55440
rect 98700 55310 98800 55440
rect 98950 55310 99050 55440
rect 99200 55310 99300 55440
rect 99450 55310 99550 55440
rect 99700 55310 99800 55440
rect 99950 55310 100050 55440
rect 100200 55310 100300 55440
rect 100450 55310 100550 55440
rect 100700 55310 100800 55440
rect 100950 55310 101050 55440
rect 101200 55310 101300 55440
rect 101450 55310 101550 55440
rect 101700 55310 101800 55440
rect 101950 55310 102050 55440
rect 102200 55310 102300 55440
rect 102450 55310 102550 55440
rect 102700 55310 102800 55440
rect 102950 55310 103050 55440
rect 103200 55310 103300 55440
rect 103450 55310 103550 55440
rect 103700 55310 103800 55440
rect 103950 55310 104050 55440
rect 104200 55310 104300 55440
rect 104450 55310 104550 55440
rect 104700 55310 104800 55440
rect 104950 55310 105050 55440
rect 105200 55310 105300 55440
rect 105450 55310 105550 55440
rect 105700 55310 105800 55440
rect 105950 55310 106050 55440
rect 106200 55310 106300 55440
rect 106450 55310 106550 55440
rect 106700 55310 106800 55440
rect 106950 55310 107050 55440
rect 107200 55310 107300 55440
rect 107450 55310 107550 55440
rect 107700 55310 107800 55440
rect 107950 55310 108050 55440
rect 108200 55310 108300 55440
rect 108450 55310 108550 55440
rect 108700 55310 108800 55440
rect 108950 55310 109050 55440
rect 109200 55310 109300 55440
rect 109450 55310 109550 55440
rect 109700 55310 109800 55440
rect 109950 55310 110050 55440
rect 110200 55310 110300 55440
rect 110450 55310 110550 55440
rect 110700 55310 110800 55440
rect 110950 55310 111050 55440
rect 111200 55310 111300 55440
rect 111450 55310 111550 55440
rect 111700 55310 111800 55440
rect 111950 55310 112050 55440
rect 112200 55310 112300 55440
rect 112450 55310 112550 55440
rect 112700 55310 112800 55440
rect 112950 55310 113050 55440
rect 113200 55310 113300 55440
rect 113450 55310 113550 55440
rect 113700 55310 113800 55440
rect 113950 55310 114050 55440
rect 114200 55310 114300 55440
rect 114450 55310 114550 55440
rect 114700 55310 114800 55440
rect 114950 55310 115050 55440
rect 115200 55310 115300 55440
rect 115450 55310 115550 55440
rect 115700 55310 115800 55440
rect 115950 55310 116000 55440
rect 89000 55300 89060 55310
rect 89190 55300 89310 55310
rect 89440 55300 89560 55310
rect 89690 55300 89810 55310
rect 89940 55300 90060 55310
rect 90190 55300 90310 55310
rect 90440 55300 90560 55310
rect 90690 55300 90810 55310
rect 90940 55300 91060 55310
rect 91190 55300 91310 55310
rect 91440 55300 91560 55310
rect 91690 55300 91810 55310
rect 91940 55300 92060 55310
rect 92190 55300 92310 55310
rect 92440 55300 92560 55310
rect 92690 55300 92810 55310
rect 92940 55300 93060 55310
rect 93190 55300 93310 55310
rect 93440 55300 93560 55310
rect 93690 55300 93810 55310
rect 93940 55300 94060 55310
rect 94190 55300 94310 55310
rect 94440 55300 94560 55310
rect 94690 55300 94810 55310
rect 94940 55300 95060 55310
rect 95190 55300 95310 55310
rect 95440 55300 95560 55310
rect 95690 55300 95810 55310
rect 95940 55300 96060 55310
rect 96190 55300 96310 55310
rect 96440 55300 96560 55310
rect 96690 55300 96810 55310
rect 96940 55300 97060 55310
rect 97190 55300 97310 55310
rect 97440 55300 97560 55310
rect 97690 55300 97810 55310
rect 97940 55300 98060 55310
rect 98190 55300 98310 55310
rect 98440 55300 98560 55310
rect 98690 55300 98810 55310
rect 98940 55300 99060 55310
rect 99190 55300 99310 55310
rect 99440 55300 99560 55310
rect 99690 55300 99810 55310
rect 99940 55300 100060 55310
rect 100190 55300 100310 55310
rect 100440 55300 100560 55310
rect 100690 55300 100810 55310
rect 100940 55300 101060 55310
rect 101190 55300 101310 55310
rect 101440 55300 101560 55310
rect 101690 55300 101810 55310
rect 101940 55300 102060 55310
rect 102190 55300 102310 55310
rect 102440 55300 102560 55310
rect 102690 55300 102810 55310
rect 102940 55300 103060 55310
rect 103190 55300 103310 55310
rect 103440 55300 103560 55310
rect 103690 55300 103810 55310
rect 103940 55300 104060 55310
rect 104190 55300 104310 55310
rect 104440 55300 104560 55310
rect 104690 55300 104810 55310
rect 104940 55300 105060 55310
rect 105190 55300 105310 55310
rect 105440 55300 105560 55310
rect 105690 55300 105810 55310
rect 105940 55300 106060 55310
rect 106190 55300 106310 55310
rect 106440 55300 106560 55310
rect 106690 55300 106810 55310
rect 106940 55300 107060 55310
rect 107190 55300 107310 55310
rect 107440 55300 107560 55310
rect 107690 55300 107810 55310
rect 107940 55300 108060 55310
rect 108190 55300 108310 55310
rect 108440 55300 108560 55310
rect 108690 55300 108810 55310
rect 108940 55300 109060 55310
rect 109190 55300 109310 55310
rect 109440 55300 109560 55310
rect 109690 55300 109810 55310
rect 109940 55300 110060 55310
rect 110190 55300 110310 55310
rect 110440 55300 110560 55310
rect 110690 55300 110810 55310
rect 110940 55300 111060 55310
rect 111190 55300 111310 55310
rect 111440 55300 111560 55310
rect 111690 55300 111810 55310
rect 111940 55300 112060 55310
rect 112190 55300 112310 55310
rect 112440 55300 112560 55310
rect 112690 55300 112810 55310
rect 112940 55300 113060 55310
rect 113190 55300 113310 55310
rect 113440 55300 113560 55310
rect 113690 55300 113810 55310
rect 113940 55300 114060 55310
rect 114190 55300 114310 55310
rect 114440 55300 114560 55310
rect 114690 55300 114810 55310
rect 114940 55300 115060 55310
rect 115190 55300 115310 55310
rect 115440 55300 115560 55310
rect 115690 55300 115810 55310
rect 115940 55300 116000 55310
rect 89000 55200 116000 55300
rect 89000 55190 89060 55200
rect 89190 55190 89310 55200
rect 89440 55190 89560 55200
rect 89690 55190 89810 55200
rect 89940 55190 90060 55200
rect 90190 55190 90310 55200
rect 90440 55190 90560 55200
rect 90690 55190 90810 55200
rect 90940 55190 91060 55200
rect 91190 55190 91310 55200
rect 91440 55190 91560 55200
rect 91690 55190 91810 55200
rect 91940 55190 92060 55200
rect 92190 55190 92310 55200
rect 92440 55190 92560 55200
rect 92690 55190 92810 55200
rect 92940 55190 93060 55200
rect 93190 55190 93310 55200
rect 93440 55190 93560 55200
rect 93690 55190 93810 55200
rect 93940 55190 94060 55200
rect 94190 55190 94310 55200
rect 94440 55190 94560 55200
rect 94690 55190 94810 55200
rect 94940 55190 95060 55200
rect 95190 55190 95310 55200
rect 95440 55190 95560 55200
rect 95690 55190 95810 55200
rect 95940 55190 96060 55200
rect 96190 55190 96310 55200
rect 96440 55190 96560 55200
rect 96690 55190 96810 55200
rect 96940 55190 97060 55200
rect 97190 55190 97310 55200
rect 97440 55190 97560 55200
rect 97690 55190 97810 55200
rect 97940 55190 98060 55200
rect 98190 55190 98310 55200
rect 98440 55190 98560 55200
rect 98690 55190 98810 55200
rect 98940 55190 99060 55200
rect 99190 55190 99310 55200
rect 99440 55190 99560 55200
rect 99690 55190 99810 55200
rect 99940 55190 100060 55200
rect 100190 55190 100310 55200
rect 100440 55190 100560 55200
rect 100690 55190 100810 55200
rect 100940 55190 101060 55200
rect 101190 55190 101310 55200
rect 101440 55190 101560 55200
rect 101690 55190 101810 55200
rect 101940 55190 102060 55200
rect 102190 55190 102310 55200
rect 102440 55190 102560 55200
rect 102690 55190 102810 55200
rect 102940 55190 103060 55200
rect 103190 55190 103310 55200
rect 103440 55190 103560 55200
rect 103690 55190 103810 55200
rect 103940 55190 104060 55200
rect 104190 55190 104310 55200
rect 104440 55190 104560 55200
rect 104690 55190 104810 55200
rect 104940 55190 105060 55200
rect 105190 55190 105310 55200
rect 105440 55190 105560 55200
rect 105690 55190 105810 55200
rect 105940 55190 106060 55200
rect 106190 55190 106310 55200
rect 106440 55190 106560 55200
rect 106690 55190 106810 55200
rect 106940 55190 107060 55200
rect 107190 55190 107310 55200
rect 107440 55190 107560 55200
rect 107690 55190 107810 55200
rect 107940 55190 108060 55200
rect 108190 55190 108310 55200
rect 108440 55190 108560 55200
rect 108690 55190 108810 55200
rect 108940 55190 109060 55200
rect 109190 55190 109310 55200
rect 109440 55190 109560 55200
rect 109690 55190 109810 55200
rect 109940 55190 110060 55200
rect 110190 55190 110310 55200
rect 110440 55190 110560 55200
rect 110690 55190 110810 55200
rect 110940 55190 111060 55200
rect 111190 55190 111310 55200
rect 111440 55190 111560 55200
rect 111690 55190 111810 55200
rect 111940 55190 112060 55200
rect 112190 55190 112310 55200
rect 112440 55190 112560 55200
rect 112690 55190 112810 55200
rect 112940 55190 113060 55200
rect 113190 55190 113310 55200
rect 113440 55190 113560 55200
rect 113690 55190 113810 55200
rect 113940 55190 114060 55200
rect 114190 55190 114310 55200
rect 114440 55190 114560 55200
rect 114690 55190 114810 55200
rect 114940 55190 115060 55200
rect 115190 55190 115310 55200
rect 115440 55190 115560 55200
rect 115690 55190 115810 55200
rect 115940 55190 116000 55200
rect 89000 55060 89050 55190
rect 89200 55060 89300 55190
rect 89450 55060 89550 55190
rect 89700 55060 89800 55190
rect 89950 55060 90050 55190
rect 90200 55060 90300 55190
rect 90450 55060 90550 55190
rect 90700 55060 90800 55190
rect 90950 55060 91050 55190
rect 91200 55060 91300 55190
rect 91450 55060 91550 55190
rect 91700 55060 91800 55190
rect 91950 55060 92050 55190
rect 92200 55060 92300 55190
rect 92450 55060 92550 55190
rect 92700 55060 92800 55190
rect 92950 55060 93050 55190
rect 93200 55060 93300 55190
rect 93450 55060 93550 55190
rect 93700 55060 93800 55190
rect 93950 55060 94050 55190
rect 94200 55060 94300 55190
rect 94450 55060 94550 55190
rect 94700 55060 94800 55190
rect 94950 55060 95050 55190
rect 95200 55060 95300 55190
rect 95450 55060 95550 55190
rect 95700 55060 95800 55190
rect 95950 55060 96050 55190
rect 96200 55060 96300 55190
rect 96450 55060 96550 55190
rect 96700 55060 96800 55190
rect 96950 55060 97050 55190
rect 97200 55060 97300 55190
rect 97450 55060 97550 55190
rect 97700 55060 97800 55190
rect 97950 55060 98050 55190
rect 98200 55060 98300 55190
rect 98450 55060 98550 55190
rect 98700 55060 98800 55190
rect 98950 55060 99050 55190
rect 99200 55060 99300 55190
rect 99450 55060 99550 55190
rect 99700 55060 99800 55190
rect 99950 55060 100050 55190
rect 100200 55060 100300 55190
rect 100450 55060 100550 55190
rect 100700 55060 100800 55190
rect 100950 55060 101050 55190
rect 101200 55060 101300 55190
rect 101450 55060 101550 55190
rect 101700 55060 101800 55190
rect 101950 55060 102050 55190
rect 102200 55060 102300 55190
rect 102450 55060 102550 55190
rect 102700 55060 102800 55190
rect 102950 55060 103050 55190
rect 103200 55060 103300 55190
rect 103450 55060 103550 55190
rect 103700 55060 103800 55190
rect 103950 55060 104050 55190
rect 104200 55060 104300 55190
rect 104450 55060 104550 55190
rect 104700 55060 104800 55190
rect 104950 55060 105050 55190
rect 105200 55060 105300 55190
rect 105450 55060 105550 55190
rect 105700 55060 105800 55190
rect 105950 55060 106050 55190
rect 106200 55060 106300 55190
rect 106450 55060 106550 55190
rect 106700 55060 106800 55190
rect 106950 55060 107050 55190
rect 107200 55060 107300 55190
rect 107450 55060 107550 55190
rect 107700 55060 107800 55190
rect 107950 55060 108050 55190
rect 108200 55060 108300 55190
rect 108450 55060 108550 55190
rect 108700 55060 108800 55190
rect 108950 55060 109050 55190
rect 109200 55060 109300 55190
rect 109450 55060 109550 55190
rect 109700 55060 109800 55190
rect 109950 55060 110050 55190
rect 110200 55060 110300 55190
rect 110450 55060 110550 55190
rect 110700 55060 110800 55190
rect 110950 55060 111050 55190
rect 111200 55060 111300 55190
rect 111450 55060 111550 55190
rect 111700 55060 111800 55190
rect 111950 55060 112050 55190
rect 112200 55060 112300 55190
rect 112450 55060 112550 55190
rect 112700 55060 112800 55190
rect 112950 55060 113050 55190
rect 113200 55060 113300 55190
rect 113450 55060 113550 55190
rect 113700 55060 113800 55190
rect 113950 55060 114050 55190
rect 114200 55060 114300 55190
rect 114450 55060 114550 55190
rect 114700 55060 114800 55190
rect 114950 55060 115050 55190
rect 115200 55060 115300 55190
rect 115450 55060 115550 55190
rect 115700 55060 115800 55190
rect 115950 55060 116000 55190
rect 89000 55050 89060 55060
rect 89190 55050 89310 55060
rect 89440 55050 89560 55060
rect 89690 55050 89810 55060
rect 89940 55050 90060 55060
rect 90190 55050 90310 55060
rect 90440 55050 90560 55060
rect 90690 55050 90810 55060
rect 90940 55050 91060 55060
rect 91190 55050 91310 55060
rect 91440 55050 91560 55060
rect 91690 55050 91810 55060
rect 91940 55050 92060 55060
rect 92190 55050 92310 55060
rect 92440 55050 92560 55060
rect 92690 55050 92810 55060
rect 92940 55050 93060 55060
rect 93190 55050 93310 55060
rect 93440 55050 93560 55060
rect 93690 55050 93810 55060
rect 93940 55050 94060 55060
rect 94190 55050 94310 55060
rect 94440 55050 94560 55060
rect 94690 55050 94810 55060
rect 94940 55050 95060 55060
rect 95190 55050 95310 55060
rect 95440 55050 95560 55060
rect 95690 55050 95810 55060
rect 95940 55050 96060 55060
rect 96190 55050 96310 55060
rect 96440 55050 96560 55060
rect 96690 55050 96810 55060
rect 96940 55050 97060 55060
rect 97190 55050 97310 55060
rect 97440 55050 97560 55060
rect 97690 55050 97810 55060
rect 97940 55050 98060 55060
rect 98190 55050 98310 55060
rect 98440 55050 98560 55060
rect 98690 55050 98810 55060
rect 98940 55050 99060 55060
rect 99190 55050 99310 55060
rect 99440 55050 99560 55060
rect 99690 55050 99810 55060
rect 99940 55050 100060 55060
rect 100190 55050 100310 55060
rect 100440 55050 100560 55060
rect 100690 55050 100810 55060
rect 100940 55050 101060 55060
rect 101190 55050 101310 55060
rect 101440 55050 101560 55060
rect 101690 55050 101810 55060
rect 101940 55050 102060 55060
rect 102190 55050 102310 55060
rect 102440 55050 102560 55060
rect 102690 55050 102810 55060
rect 102940 55050 103060 55060
rect 103190 55050 103310 55060
rect 103440 55050 103560 55060
rect 103690 55050 103810 55060
rect 103940 55050 104060 55060
rect 104190 55050 104310 55060
rect 104440 55050 104560 55060
rect 104690 55050 104810 55060
rect 104940 55050 105060 55060
rect 105190 55050 105310 55060
rect 105440 55050 105560 55060
rect 105690 55050 105810 55060
rect 105940 55050 106060 55060
rect 106190 55050 106310 55060
rect 106440 55050 106560 55060
rect 106690 55050 106810 55060
rect 106940 55050 107060 55060
rect 107190 55050 107310 55060
rect 107440 55050 107560 55060
rect 107690 55050 107810 55060
rect 107940 55050 108060 55060
rect 108190 55050 108310 55060
rect 108440 55050 108560 55060
rect 108690 55050 108810 55060
rect 108940 55050 109060 55060
rect 109190 55050 109310 55060
rect 109440 55050 109560 55060
rect 109690 55050 109810 55060
rect 109940 55050 110060 55060
rect 110190 55050 110310 55060
rect 110440 55050 110560 55060
rect 110690 55050 110810 55060
rect 110940 55050 111060 55060
rect 111190 55050 111310 55060
rect 111440 55050 111560 55060
rect 111690 55050 111810 55060
rect 111940 55050 112060 55060
rect 112190 55050 112310 55060
rect 112440 55050 112560 55060
rect 112690 55050 112810 55060
rect 112940 55050 113060 55060
rect 113190 55050 113310 55060
rect 113440 55050 113560 55060
rect 113690 55050 113810 55060
rect 113940 55050 114060 55060
rect 114190 55050 114310 55060
rect 114440 55050 114560 55060
rect 114690 55050 114810 55060
rect 114940 55050 115060 55060
rect 115190 55050 115310 55060
rect 115440 55050 115560 55060
rect 115690 55050 115810 55060
rect 115940 55050 116000 55060
rect 89000 54950 116000 55050
rect 89000 54940 89060 54950
rect 89190 54940 89310 54950
rect 89440 54940 89560 54950
rect 89690 54940 89810 54950
rect 89940 54940 90060 54950
rect 90190 54940 90310 54950
rect 90440 54940 90560 54950
rect 90690 54940 90810 54950
rect 90940 54940 91060 54950
rect 91190 54940 91310 54950
rect 91440 54940 91560 54950
rect 91690 54940 91810 54950
rect 91940 54940 92060 54950
rect 92190 54940 92310 54950
rect 92440 54940 92560 54950
rect 92690 54940 92810 54950
rect 92940 54940 93060 54950
rect 93190 54940 93310 54950
rect 93440 54940 93560 54950
rect 93690 54940 93810 54950
rect 93940 54940 94060 54950
rect 94190 54940 94310 54950
rect 94440 54940 94560 54950
rect 94690 54940 94810 54950
rect 94940 54940 95060 54950
rect 95190 54940 95310 54950
rect 95440 54940 95560 54950
rect 95690 54940 95810 54950
rect 95940 54940 96060 54950
rect 96190 54940 96310 54950
rect 96440 54940 96560 54950
rect 96690 54940 96810 54950
rect 96940 54940 97060 54950
rect 97190 54940 97310 54950
rect 97440 54940 97560 54950
rect 97690 54940 97810 54950
rect 97940 54940 98060 54950
rect 98190 54940 98310 54950
rect 98440 54940 98560 54950
rect 98690 54940 98810 54950
rect 98940 54940 99060 54950
rect 99190 54940 99310 54950
rect 99440 54940 99560 54950
rect 99690 54940 99810 54950
rect 99940 54940 100060 54950
rect 100190 54940 100310 54950
rect 100440 54940 100560 54950
rect 100690 54940 100810 54950
rect 100940 54940 101060 54950
rect 101190 54940 101310 54950
rect 101440 54940 101560 54950
rect 101690 54940 101810 54950
rect 101940 54940 102060 54950
rect 102190 54940 102310 54950
rect 102440 54940 102560 54950
rect 102690 54940 102810 54950
rect 102940 54940 103060 54950
rect 103190 54940 103310 54950
rect 103440 54940 103560 54950
rect 103690 54940 103810 54950
rect 103940 54940 104060 54950
rect 104190 54940 104310 54950
rect 104440 54940 104560 54950
rect 104690 54940 104810 54950
rect 104940 54940 105060 54950
rect 105190 54940 105310 54950
rect 105440 54940 105560 54950
rect 105690 54940 105810 54950
rect 105940 54940 106060 54950
rect 106190 54940 106310 54950
rect 106440 54940 106560 54950
rect 106690 54940 106810 54950
rect 106940 54940 107060 54950
rect 107190 54940 107310 54950
rect 107440 54940 107560 54950
rect 107690 54940 107810 54950
rect 107940 54940 108060 54950
rect 108190 54940 108310 54950
rect 108440 54940 108560 54950
rect 108690 54940 108810 54950
rect 108940 54940 109060 54950
rect 109190 54940 109310 54950
rect 109440 54940 109560 54950
rect 109690 54940 109810 54950
rect 109940 54940 110060 54950
rect 110190 54940 110310 54950
rect 110440 54940 110560 54950
rect 110690 54940 110810 54950
rect 110940 54940 111060 54950
rect 111190 54940 111310 54950
rect 111440 54940 111560 54950
rect 111690 54940 111810 54950
rect 111940 54940 112060 54950
rect 112190 54940 112310 54950
rect 112440 54940 112560 54950
rect 112690 54940 112810 54950
rect 112940 54940 113060 54950
rect 113190 54940 113310 54950
rect 113440 54940 113560 54950
rect 113690 54940 113810 54950
rect 113940 54940 114060 54950
rect 114190 54940 114310 54950
rect 114440 54940 114560 54950
rect 114690 54940 114810 54950
rect 114940 54940 115060 54950
rect 115190 54940 115310 54950
rect 115440 54940 115560 54950
rect 115690 54940 115810 54950
rect 115940 54940 116000 54950
rect 89000 54810 89050 54940
rect 89200 54810 89300 54940
rect 89450 54810 89550 54940
rect 89700 54810 89800 54940
rect 89950 54810 90050 54940
rect 90200 54810 90300 54940
rect 90450 54810 90550 54940
rect 90700 54810 90800 54940
rect 90950 54810 91050 54940
rect 91200 54810 91300 54940
rect 91450 54810 91550 54940
rect 91700 54810 91800 54940
rect 91950 54810 92050 54940
rect 92200 54810 92300 54940
rect 92450 54810 92550 54940
rect 92700 54810 92800 54940
rect 92950 54810 93050 54940
rect 93200 54810 93300 54940
rect 93450 54810 93550 54940
rect 93700 54810 93800 54940
rect 93950 54810 94050 54940
rect 94200 54810 94300 54940
rect 94450 54810 94550 54940
rect 94700 54810 94800 54940
rect 94950 54810 95050 54940
rect 95200 54810 95300 54940
rect 95450 54810 95550 54940
rect 95700 54810 95800 54940
rect 95950 54810 96050 54940
rect 96200 54810 96300 54940
rect 96450 54810 96550 54940
rect 96700 54810 96800 54940
rect 96950 54810 97050 54940
rect 97200 54810 97300 54940
rect 97450 54810 97550 54940
rect 97700 54810 97800 54940
rect 97950 54810 98050 54940
rect 98200 54810 98300 54940
rect 98450 54810 98550 54940
rect 98700 54810 98800 54940
rect 98950 54810 99050 54940
rect 99200 54810 99300 54940
rect 99450 54810 99550 54940
rect 99700 54810 99800 54940
rect 99950 54810 100050 54940
rect 100200 54810 100300 54940
rect 100450 54810 100550 54940
rect 100700 54810 100800 54940
rect 100950 54810 101050 54940
rect 101200 54810 101300 54940
rect 101450 54810 101550 54940
rect 101700 54810 101800 54940
rect 101950 54810 102050 54940
rect 102200 54810 102300 54940
rect 102450 54810 102550 54940
rect 102700 54810 102800 54940
rect 102950 54810 103050 54940
rect 103200 54810 103300 54940
rect 103450 54810 103550 54940
rect 103700 54810 103800 54940
rect 103950 54810 104050 54940
rect 104200 54810 104300 54940
rect 104450 54810 104550 54940
rect 104700 54810 104800 54940
rect 104950 54810 105050 54940
rect 105200 54810 105300 54940
rect 105450 54810 105550 54940
rect 105700 54810 105800 54940
rect 105950 54810 106050 54940
rect 106200 54810 106300 54940
rect 106450 54810 106550 54940
rect 106700 54810 106800 54940
rect 106950 54810 107050 54940
rect 107200 54810 107300 54940
rect 107450 54810 107550 54940
rect 107700 54810 107800 54940
rect 107950 54810 108050 54940
rect 108200 54810 108300 54940
rect 108450 54810 108550 54940
rect 108700 54810 108800 54940
rect 108950 54810 109050 54940
rect 109200 54810 109300 54940
rect 109450 54810 109550 54940
rect 109700 54810 109800 54940
rect 109950 54810 110050 54940
rect 110200 54810 110300 54940
rect 110450 54810 110550 54940
rect 110700 54810 110800 54940
rect 110950 54810 111050 54940
rect 111200 54810 111300 54940
rect 111450 54810 111550 54940
rect 111700 54810 111800 54940
rect 111950 54810 112050 54940
rect 112200 54810 112300 54940
rect 112450 54810 112550 54940
rect 112700 54810 112800 54940
rect 112950 54810 113050 54940
rect 113200 54810 113300 54940
rect 113450 54810 113550 54940
rect 113700 54810 113800 54940
rect 113950 54810 114050 54940
rect 114200 54810 114300 54940
rect 114450 54810 114550 54940
rect 114700 54810 114800 54940
rect 114950 54810 115050 54940
rect 115200 54810 115300 54940
rect 115450 54810 115550 54940
rect 115700 54810 115800 54940
rect 115950 54810 116000 54940
rect 89000 54800 89060 54810
rect 89190 54800 89310 54810
rect 89440 54800 89560 54810
rect 89690 54800 89810 54810
rect 89940 54800 90060 54810
rect 90190 54800 90310 54810
rect 90440 54800 90560 54810
rect 90690 54800 90810 54810
rect 90940 54800 91060 54810
rect 91190 54800 91310 54810
rect 91440 54800 91560 54810
rect 91690 54800 91810 54810
rect 91940 54800 92060 54810
rect 92190 54800 92310 54810
rect 92440 54800 92560 54810
rect 92690 54800 92810 54810
rect 92940 54800 93060 54810
rect 93190 54800 93310 54810
rect 93440 54800 93560 54810
rect 93690 54800 93810 54810
rect 93940 54800 94060 54810
rect 94190 54800 94310 54810
rect 94440 54800 94560 54810
rect 94690 54800 94810 54810
rect 94940 54800 95060 54810
rect 95190 54800 95310 54810
rect 95440 54800 95560 54810
rect 95690 54800 95810 54810
rect 95940 54800 96060 54810
rect 96190 54800 96310 54810
rect 96440 54800 96560 54810
rect 96690 54800 96810 54810
rect 96940 54800 97060 54810
rect 97190 54800 97310 54810
rect 97440 54800 97560 54810
rect 97690 54800 97810 54810
rect 97940 54800 98060 54810
rect 98190 54800 98310 54810
rect 98440 54800 98560 54810
rect 98690 54800 98810 54810
rect 98940 54800 99060 54810
rect 99190 54800 99310 54810
rect 99440 54800 99560 54810
rect 99690 54800 99810 54810
rect 99940 54800 100060 54810
rect 100190 54800 100310 54810
rect 100440 54800 100560 54810
rect 100690 54800 100810 54810
rect 100940 54800 101060 54810
rect 101190 54800 101310 54810
rect 101440 54800 101560 54810
rect 101690 54800 101810 54810
rect 101940 54800 102060 54810
rect 102190 54800 102310 54810
rect 102440 54800 102560 54810
rect 102690 54800 102810 54810
rect 102940 54800 103060 54810
rect 103190 54800 103310 54810
rect 103440 54800 103560 54810
rect 103690 54800 103810 54810
rect 103940 54800 104060 54810
rect 104190 54800 104310 54810
rect 104440 54800 104560 54810
rect 104690 54800 104810 54810
rect 104940 54800 105060 54810
rect 105190 54800 105310 54810
rect 105440 54800 105560 54810
rect 105690 54800 105810 54810
rect 105940 54800 106060 54810
rect 106190 54800 106310 54810
rect 106440 54800 106560 54810
rect 106690 54800 106810 54810
rect 106940 54800 107060 54810
rect 107190 54800 107310 54810
rect 107440 54800 107560 54810
rect 107690 54800 107810 54810
rect 107940 54800 108060 54810
rect 108190 54800 108310 54810
rect 108440 54800 108560 54810
rect 108690 54800 108810 54810
rect 108940 54800 109060 54810
rect 109190 54800 109310 54810
rect 109440 54800 109560 54810
rect 109690 54800 109810 54810
rect 109940 54800 110060 54810
rect 110190 54800 110310 54810
rect 110440 54800 110560 54810
rect 110690 54800 110810 54810
rect 110940 54800 111060 54810
rect 111190 54800 111310 54810
rect 111440 54800 111560 54810
rect 111690 54800 111810 54810
rect 111940 54800 112060 54810
rect 112190 54800 112310 54810
rect 112440 54800 112560 54810
rect 112690 54800 112810 54810
rect 112940 54800 113060 54810
rect 113190 54800 113310 54810
rect 113440 54800 113560 54810
rect 113690 54800 113810 54810
rect 113940 54800 114060 54810
rect 114190 54800 114310 54810
rect 114440 54800 114560 54810
rect 114690 54800 114810 54810
rect 114940 54800 115060 54810
rect 115190 54800 115310 54810
rect 115440 54800 115560 54810
rect 115690 54800 115810 54810
rect 115940 54800 116000 54810
rect 89000 54700 116000 54800
rect 89000 54690 89060 54700
rect 89190 54690 89310 54700
rect 89440 54690 89560 54700
rect 89690 54690 89810 54700
rect 89940 54690 90060 54700
rect 90190 54690 90310 54700
rect 90440 54690 90560 54700
rect 90690 54690 90810 54700
rect 90940 54690 91060 54700
rect 91190 54690 91310 54700
rect 91440 54690 91560 54700
rect 91690 54690 91810 54700
rect 91940 54690 92060 54700
rect 92190 54690 92310 54700
rect 92440 54690 92560 54700
rect 92690 54690 92810 54700
rect 92940 54690 93060 54700
rect 93190 54690 93310 54700
rect 93440 54690 93560 54700
rect 93690 54690 93810 54700
rect 93940 54690 94060 54700
rect 94190 54690 94310 54700
rect 94440 54690 94560 54700
rect 94690 54690 94810 54700
rect 94940 54690 95060 54700
rect 95190 54690 95310 54700
rect 95440 54690 95560 54700
rect 95690 54690 95810 54700
rect 95940 54690 96060 54700
rect 96190 54690 96310 54700
rect 96440 54690 96560 54700
rect 96690 54690 96810 54700
rect 96940 54690 97060 54700
rect 97190 54690 97310 54700
rect 97440 54690 97560 54700
rect 97690 54690 97810 54700
rect 97940 54690 98060 54700
rect 98190 54690 98310 54700
rect 98440 54690 98560 54700
rect 98690 54690 98810 54700
rect 98940 54690 99060 54700
rect 99190 54690 99310 54700
rect 99440 54690 99560 54700
rect 99690 54690 99810 54700
rect 99940 54690 100060 54700
rect 100190 54690 100310 54700
rect 100440 54690 100560 54700
rect 100690 54690 100810 54700
rect 100940 54690 101060 54700
rect 101190 54690 101310 54700
rect 101440 54690 101560 54700
rect 101690 54690 101810 54700
rect 101940 54690 102060 54700
rect 102190 54690 102310 54700
rect 102440 54690 102560 54700
rect 102690 54690 102810 54700
rect 102940 54690 103060 54700
rect 103190 54690 103310 54700
rect 103440 54690 103560 54700
rect 103690 54690 103810 54700
rect 103940 54690 104060 54700
rect 104190 54690 104310 54700
rect 104440 54690 104560 54700
rect 104690 54690 104810 54700
rect 104940 54690 105060 54700
rect 105190 54690 105310 54700
rect 105440 54690 105560 54700
rect 105690 54690 105810 54700
rect 105940 54690 106060 54700
rect 106190 54690 106310 54700
rect 106440 54690 106560 54700
rect 106690 54690 106810 54700
rect 106940 54690 107060 54700
rect 107190 54690 107310 54700
rect 107440 54690 107560 54700
rect 107690 54690 107810 54700
rect 107940 54690 108060 54700
rect 108190 54690 108310 54700
rect 108440 54690 108560 54700
rect 108690 54690 108810 54700
rect 108940 54690 109060 54700
rect 109190 54690 109310 54700
rect 109440 54690 109560 54700
rect 109690 54690 109810 54700
rect 109940 54690 110060 54700
rect 110190 54690 110310 54700
rect 110440 54690 110560 54700
rect 110690 54690 110810 54700
rect 110940 54690 111060 54700
rect 111190 54690 111310 54700
rect 111440 54690 111560 54700
rect 111690 54690 111810 54700
rect 111940 54690 112060 54700
rect 112190 54690 112310 54700
rect 112440 54690 112560 54700
rect 112690 54690 112810 54700
rect 112940 54690 113060 54700
rect 113190 54690 113310 54700
rect 113440 54690 113560 54700
rect 113690 54690 113810 54700
rect 113940 54690 114060 54700
rect 114190 54690 114310 54700
rect 114440 54690 114560 54700
rect 114690 54690 114810 54700
rect 114940 54690 115060 54700
rect 115190 54690 115310 54700
rect 115440 54690 115560 54700
rect 115690 54690 115810 54700
rect 115940 54690 116000 54700
rect 89000 54560 89050 54690
rect 89200 54560 89300 54690
rect 89450 54560 89550 54690
rect 89700 54560 89800 54690
rect 89950 54560 90050 54690
rect 90200 54560 90300 54690
rect 90450 54560 90550 54690
rect 90700 54560 90800 54690
rect 90950 54560 91050 54690
rect 91200 54560 91300 54690
rect 91450 54560 91550 54690
rect 91700 54560 91800 54690
rect 91950 54560 92050 54690
rect 92200 54560 92300 54690
rect 92450 54560 92550 54690
rect 92700 54560 92800 54690
rect 92950 54560 93050 54690
rect 93200 54560 93300 54690
rect 93450 54560 93550 54690
rect 93700 54560 93800 54690
rect 93950 54560 94050 54690
rect 94200 54560 94300 54690
rect 94450 54560 94550 54690
rect 94700 54560 94800 54690
rect 94950 54560 95050 54690
rect 95200 54560 95300 54690
rect 95450 54560 95550 54690
rect 95700 54560 95800 54690
rect 95950 54560 96050 54690
rect 96200 54560 96300 54690
rect 96450 54560 96550 54690
rect 96700 54560 96800 54690
rect 96950 54560 97050 54690
rect 97200 54560 97300 54690
rect 97450 54560 97550 54690
rect 97700 54560 97800 54690
rect 97950 54560 98050 54690
rect 98200 54560 98300 54690
rect 98450 54560 98550 54690
rect 98700 54560 98800 54690
rect 98950 54560 99050 54690
rect 99200 54560 99300 54690
rect 99450 54560 99550 54690
rect 99700 54560 99800 54690
rect 99950 54560 100050 54690
rect 100200 54560 100300 54690
rect 100450 54560 100550 54690
rect 100700 54560 100800 54690
rect 100950 54560 101050 54690
rect 101200 54560 101300 54690
rect 101450 54560 101550 54690
rect 101700 54560 101800 54690
rect 101950 54560 102050 54690
rect 102200 54560 102300 54690
rect 102450 54560 102550 54690
rect 102700 54560 102800 54690
rect 102950 54560 103050 54690
rect 103200 54560 103300 54690
rect 103450 54560 103550 54690
rect 103700 54560 103800 54690
rect 103950 54560 104050 54690
rect 104200 54560 104300 54690
rect 104450 54560 104550 54690
rect 104700 54560 104800 54690
rect 104950 54560 105050 54690
rect 105200 54560 105300 54690
rect 105450 54560 105550 54690
rect 105700 54560 105800 54690
rect 105950 54560 106050 54690
rect 106200 54560 106300 54690
rect 106450 54560 106550 54690
rect 106700 54560 106800 54690
rect 106950 54560 107050 54690
rect 107200 54560 107300 54690
rect 107450 54560 107550 54690
rect 107700 54560 107800 54690
rect 107950 54560 108050 54690
rect 108200 54560 108300 54690
rect 108450 54560 108550 54690
rect 108700 54560 108800 54690
rect 108950 54560 109050 54690
rect 109200 54560 109300 54690
rect 109450 54560 109550 54690
rect 109700 54560 109800 54690
rect 109950 54560 110050 54690
rect 110200 54560 110300 54690
rect 110450 54560 110550 54690
rect 110700 54560 110800 54690
rect 110950 54560 111050 54690
rect 111200 54560 111300 54690
rect 111450 54560 111550 54690
rect 111700 54560 111800 54690
rect 111950 54560 112050 54690
rect 112200 54560 112300 54690
rect 112450 54560 112550 54690
rect 112700 54560 112800 54690
rect 112950 54560 113050 54690
rect 113200 54560 113300 54690
rect 113450 54560 113550 54690
rect 113700 54560 113800 54690
rect 113950 54560 114050 54690
rect 114200 54560 114300 54690
rect 114450 54560 114550 54690
rect 114700 54560 114800 54690
rect 114950 54560 115050 54690
rect 115200 54560 115300 54690
rect 115450 54560 115550 54690
rect 115700 54560 115800 54690
rect 115950 54560 116000 54690
rect 89000 54550 89060 54560
rect 89190 54550 89310 54560
rect 89440 54550 89560 54560
rect 89690 54550 89810 54560
rect 89940 54550 90060 54560
rect 90190 54550 90310 54560
rect 90440 54550 90560 54560
rect 90690 54550 90810 54560
rect 90940 54550 91060 54560
rect 91190 54550 91310 54560
rect 91440 54550 91560 54560
rect 91690 54550 91810 54560
rect 91940 54550 92060 54560
rect 92190 54550 92310 54560
rect 92440 54550 92560 54560
rect 92690 54550 92810 54560
rect 92940 54550 93060 54560
rect 93190 54550 93310 54560
rect 93440 54550 93560 54560
rect 93690 54550 93810 54560
rect 93940 54550 94060 54560
rect 94190 54550 94310 54560
rect 94440 54550 94560 54560
rect 94690 54550 94810 54560
rect 94940 54550 95060 54560
rect 95190 54550 95310 54560
rect 95440 54550 95560 54560
rect 95690 54550 95810 54560
rect 95940 54550 96060 54560
rect 96190 54550 96310 54560
rect 96440 54550 96560 54560
rect 96690 54550 96810 54560
rect 96940 54550 97060 54560
rect 97190 54550 97310 54560
rect 97440 54550 97560 54560
rect 97690 54550 97810 54560
rect 97940 54550 98060 54560
rect 98190 54550 98310 54560
rect 98440 54550 98560 54560
rect 98690 54550 98810 54560
rect 98940 54550 99060 54560
rect 99190 54550 99310 54560
rect 99440 54550 99560 54560
rect 99690 54550 99810 54560
rect 99940 54550 100060 54560
rect 100190 54550 100310 54560
rect 100440 54550 100560 54560
rect 100690 54550 100810 54560
rect 100940 54550 101060 54560
rect 101190 54550 101310 54560
rect 101440 54550 101560 54560
rect 101690 54550 101810 54560
rect 101940 54550 102060 54560
rect 102190 54550 102310 54560
rect 102440 54550 102560 54560
rect 102690 54550 102810 54560
rect 102940 54550 103060 54560
rect 103190 54550 103310 54560
rect 103440 54550 103560 54560
rect 103690 54550 103810 54560
rect 103940 54550 104060 54560
rect 104190 54550 104310 54560
rect 104440 54550 104560 54560
rect 104690 54550 104810 54560
rect 104940 54550 105060 54560
rect 105190 54550 105310 54560
rect 105440 54550 105560 54560
rect 105690 54550 105810 54560
rect 105940 54550 106060 54560
rect 106190 54550 106310 54560
rect 106440 54550 106560 54560
rect 106690 54550 106810 54560
rect 106940 54550 107060 54560
rect 107190 54550 107310 54560
rect 107440 54550 107560 54560
rect 107690 54550 107810 54560
rect 107940 54550 108060 54560
rect 108190 54550 108310 54560
rect 108440 54550 108560 54560
rect 108690 54550 108810 54560
rect 108940 54550 109060 54560
rect 109190 54550 109310 54560
rect 109440 54550 109560 54560
rect 109690 54550 109810 54560
rect 109940 54550 110060 54560
rect 110190 54550 110310 54560
rect 110440 54550 110560 54560
rect 110690 54550 110810 54560
rect 110940 54550 111060 54560
rect 111190 54550 111310 54560
rect 111440 54550 111560 54560
rect 111690 54550 111810 54560
rect 111940 54550 112060 54560
rect 112190 54550 112310 54560
rect 112440 54550 112560 54560
rect 112690 54550 112810 54560
rect 112940 54550 113060 54560
rect 113190 54550 113310 54560
rect 113440 54550 113560 54560
rect 113690 54550 113810 54560
rect 113940 54550 114060 54560
rect 114190 54550 114310 54560
rect 114440 54550 114560 54560
rect 114690 54550 114810 54560
rect 114940 54550 115060 54560
rect 115190 54550 115310 54560
rect 115440 54550 115560 54560
rect 115690 54550 115810 54560
rect 115940 54550 116000 54560
rect 89000 54450 116000 54550
rect 89000 54440 89060 54450
rect 89190 54440 89310 54450
rect 89440 54440 89560 54450
rect 89690 54440 89810 54450
rect 89940 54440 90060 54450
rect 90190 54440 90310 54450
rect 90440 54440 90560 54450
rect 90690 54440 90810 54450
rect 90940 54440 91060 54450
rect 91190 54440 91310 54450
rect 91440 54440 91560 54450
rect 91690 54440 91810 54450
rect 91940 54440 92060 54450
rect 92190 54440 92310 54450
rect 92440 54440 92560 54450
rect 92690 54440 92810 54450
rect 92940 54440 93060 54450
rect 93190 54440 93310 54450
rect 93440 54440 93560 54450
rect 93690 54440 93810 54450
rect 93940 54440 94060 54450
rect 94190 54440 94310 54450
rect 94440 54440 94560 54450
rect 94690 54440 94810 54450
rect 94940 54440 95060 54450
rect 95190 54440 95310 54450
rect 95440 54440 95560 54450
rect 95690 54440 95810 54450
rect 95940 54440 96060 54450
rect 96190 54440 96310 54450
rect 96440 54440 96560 54450
rect 96690 54440 96810 54450
rect 96940 54440 97060 54450
rect 97190 54440 97310 54450
rect 97440 54440 97560 54450
rect 97690 54440 97810 54450
rect 97940 54440 98060 54450
rect 98190 54440 98310 54450
rect 98440 54440 98560 54450
rect 98690 54440 98810 54450
rect 98940 54440 99060 54450
rect 99190 54440 99310 54450
rect 99440 54440 99560 54450
rect 99690 54440 99810 54450
rect 99940 54440 100060 54450
rect 100190 54440 100310 54450
rect 100440 54440 100560 54450
rect 100690 54440 100810 54450
rect 100940 54440 101060 54450
rect 101190 54440 101310 54450
rect 101440 54440 101560 54450
rect 101690 54440 101810 54450
rect 101940 54440 102060 54450
rect 102190 54440 102310 54450
rect 102440 54440 102560 54450
rect 102690 54440 102810 54450
rect 102940 54440 103060 54450
rect 103190 54440 103310 54450
rect 103440 54440 103560 54450
rect 103690 54440 103810 54450
rect 103940 54440 104060 54450
rect 104190 54440 104310 54450
rect 104440 54440 104560 54450
rect 104690 54440 104810 54450
rect 104940 54440 105060 54450
rect 105190 54440 105310 54450
rect 105440 54440 105560 54450
rect 105690 54440 105810 54450
rect 105940 54440 106060 54450
rect 106190 54440 106310 54450
rect 106440 54440 106560 54450
rect 106690 54440 106810 54450
rect 106940 54440 107060 54450
rect 107190 54440 107310 54450
rect 107440 54440 107560 54450
rect 107690 54440 107810 54450
rect 107940 54440 108060 54450
rect 108190 54440 108310 54450
rect 108440 54440 108560 54450
rect 108690 54440 108810 54450
rect 108940 54440 109060 54450
rect 109190 54440 109310 54450
rect 109440 54440 109560 54450
rect 109690 54440 109810 54450
rect 109940 54440 110060 54450
rect 110190 54440 110310 54450
rect 110440 54440 110560 54450
rect 110690 54440 110810 54450
rect 110940 54440 111060 54450
rect 111190 54440 111310 54450
rect 111440 54440 111560 54450
rect 111690 54440 111810 54450
rect 111940 54440 112060 54450
rect 112190 54440 112310 54450
rect 112440 54440 112560 54450
rect 112690 54440 112810 54450
rect 112940 54440 113060 54450
rect 113190 54440 113310 54450
rect 113440 54440 113560 54450
rect 113690 54440 113810 54450
rect 113940 54440 114060 54450
rect 114190 54440 114310 54450
rect 114440 54440 114560 54450
rect 114690 54440 114810 54450
rect 114940 54440 115060 54450
rect 115190 54440 115310 54450
rect 115440 54440 115560 54450
rect 115690 54440 115810 54450
rect 115940 54440 116000 54450
rect 89000 54310 89050 54440
rect 89200 54310 89300 54440
rect 89450 54310 89550 54440
rect 89700 54310 89800 54440
rect 89950 54310 90050 54440
rect 90200 54310 90300 54440
rect 90450 54310 90550 54440
rect 90700 54310 90800 54440
rect 90950 54310 91050 54440
rect 91200 54310 91300 54440
rect 91450 54310 91550 54440
rect 91700 54310 91800 54440
rect 91950 54310 92050 54440
rect 92200 54310 92300 54440
rect 92450 54310 92550 54440
rect 92700 54310 92800 54440
rect 92950 54310 93050 54440
rect 93200 54310 93300 54440
rect 93450 54310 93550 54440
rect 93700 54310 93800 54440
rect 93950 54310 94050 54440
rect 94200 54310 94300 54440
rect 94450 54310 94550 54440
rect 94700 54310 94800 54440
rect 94950 54310 95050 54440
rect 95200 54310 95300 54440
rect 95450 54310 95550 54440
rect 95700 54310 95800 54440
rect 95950 54310 96050 54440
rect 96200 54310 96300 54440
rect 96450 54310 96550 54440
rect 96700 54310 96800 54440
rect 96950 54310 97050 54440
rect 97200 54310 97300 54440
rect 97450 54310 97550 54440
rect 97700 54310 97800 54440
rect 97950 54310 98050 54440
rect 98200 54310 98300 54440
rect 98450 54310 98550 54440
rect 98700 54310 98800 54440
rect 98950 54310 99050 54440
rect 99200 54310 99300 54440
rect 99450 54310 99550 54440
rect 99700 54310 99800 54440
rect 99950 54310 100050 54440
rect 100200 54310 100300 54440
rect 100450 54310 100550 54440
rect 100700 54310 100800 54440
rect 100950 54310 101050 54440
rect 101200 54310 101300 54440
rect 101450 54310 101550 54440
rect 101700 54310 101800 54440
rect 101950 54310 102050 54440
rect 102200 54310 102300 54440
rect 102450 54310 102550 54440
rect 102700 54310 102800 54440
rect 102950 54310 103050 54440
rect 103200 54310 103300 54440
rect 103450 54310 103550 54440
rect 103700 54310 103800 54440
rect 103950 54310 104050 54440
rect 104200 54310 104300 54440
rect 104450 54310 104550 54440
rect 104700 54310 104800 54440
rect 104950 54310 105050 54440
rect 105200 54310 105300 54440
rect 105450 54310 105550 54440
rect 105700 54310 105800 54440
rect 105950 54310 106050 54440
rect 106200 54310 106300 54440
rect 106450 54310 106550 54440
rect 106700 54310 106800 54440
rect 106950 54310 107050 54440
rect 107200 54310 107300 54440
rect 107450 54310 107550 54440
rect 107700 54310 107800 54440
rect 107950 54310 108050 54440
rect 108200 54310 108300 54440
rect 108450 54310 108550 54440
rect 108700 54310 108800 54440
rect 108950 54310 109050 54440
rect 109200 54310 109300 54440
rect 109450 54310 109550 54440
rect 109700 54310 109800 54440
rect 109950 54310 110050 54440
rect 110200 54310 110300 54440
rect 110450 54310 110550 54440
rect 110700 54310 110800 54440
rect 110950 54310 111050 54440
rect 111200 54310 111300 54440
rect 111450 54310 111550 54440
rect 111700 54310 111800 54440
rect 111950 54310 112050 54440
rect 112200 54310 112300 54440
rect 112450 54310 112550 54440
rect 112700 54310 112800 54440
rect 112950 54310 113050 54440
rect 113200 54310 113300 54440
rect 113450 54310 113550 54440
rect 113700 54310 113800 54440
rect 113950 54310 114050 54440
rect 114200 54310 114300 54440
rect 114450 54310 114550 54440
rect 114700 54310 114800 54440
rect 114950 54310 115050 54440
rect 115200 54310 115300 54440
rect 115450 54310 115550 54440
rect 115700 54310 115800 54440
rect 115950 54310 116000 54440
rect 89000 54300 89060 54310
rect 89190 54300 89310 54310
rect 89440 54300 89560 54310
rect 89690 54300 89810 54310
rect 89940 54300 90060 54310
rect 90190 54300 90310 54310
rect 90440 54300 90560 54310
rect 90690 54300 90810 54310
rect 90940 54300 91060 54310
rect 91190 54300 91310 54310
rect 91440 54300 91560 54310
rect 91690 54300 91810 54310
rect 91940 54300 92060 54310
rect 92190 54300 92310 54310
rect 92440 54300 92560 54310
rect 92690 54300 92810 54310
rect 92940 54300 93060 54310
rect 93190 54300 93310 54310
rect 93440 54300 93560 54310
rect 93690 54300 93810 54310
rect 93940 54300 94060 54310
rect 94190 54300 94310 54310
rect 94440 54300 94560 54310
rect 94690 54300 94810 54310
rect 94940 54300 95060 54310
rect 95190 54300 95310 54310
rect 95440 54300 95560 54310
rect 95690 54300 95810 54310
rect 95940 54300 96060 54310
rect 96190 54300 96310 54310
rect 96440 54300 96560 54310
rect 96690 54300 96810 54310
rect 96940 54300 97060 54310
rect 97190 54300 97310 54310
rect 97440 54300 97560 54310
rect 97690 54300 97810 54310
rect 97940 54300 98060 54310
rect 98190 54300 98310 54310
rect 98440 54300 98560 54310
rect 98690 54300 98810 54310
rect 98940 54300 99060 54310
rect 99190 54300 99310 54310
rect 99440 54300 99560 54310
rect 99690 54300 99810 54310
rect 99940 54300 100060 54310
rect 100190 54300 100310 54310
rect 100440 54300 100560 54310
rect 100690 54300 100810 54310
rect 100940 54300 101060 54310
rect 101190 54300 101310 54310
rect 101440 54300 101560 54310
rect 101690 54300 101810 54310
rect 101940 54300 102060 54310
rect 102190 54300 102310 54310
rect 102440 54300 102560 54310
rect 102690 54300 102810 54310
rect 102940 54300 103060 54310
rect 103190 54300 103310 54310
rect 103440 54300 103560 54310
rect 103690 54300 103810 54310
rect 103940 54300 104060 54310
rect 104190 54300 104310 54310
rect 104440 54300 104560 54310
rect 104690 54300 104810 54310
rect 104940 54300 105060 54310
rect 105190 54300 105310 54310
rect 105440 54300 105560 54310
rect 105690 54300 105810 54310
rect 105940 54300 106060 54310
rect 106190 54300 106310 54310
rect 106440 54300 106560 54310
rect 106690 54300 106810 54310
rect 106940 54300 107060 54310
rect 107190 54300 107310 54310
rect 107440 54300 107560 54310
rect 107690 54300 107810 54310
rect 107940 54300 108060 54310
rect 108190 54300 108310 54310
rect 108440 54300 108560 54310
rect 108690 54300 108810 54310
rect 108940 54300 109060 54310
rect 109190 54300 109310 54310
rect 109440 54300 109560 54310
rect 109690 54300 109810 54310
rect 109940 54300 110060 54310
rect 110190 54300 110310 54310
rect 110440 54300 110560 54310
rect 110690 54300 110810 54310
rect 110940 54300 111060 54310
rect 111190 54300 111310 54310
rect 111440 54300 111560 54310
rect 111690 54300 111810 54310
rect 111940 54300 112060 54310
rect 112190 54300 112310 54310
rect 112440 54300 112560 54310
rect 112690 54300 112810 54310
rect 112940 54300 113060 54310
rect 113190 54300 113310 54310
rect 113440 54300 113560 54310
rect 113690 54300 113810 54310
rect 113940 54300 114060 54310
rect 114190 54300 114310 54310
rect 114440 54300 114560 54310
rect 114690 54300 114810 54310
rect 114940 54300 115060 54310
rect 115190 54300 115310 54310
rect 115440 54300 115560 54310
rect 115690 54300 115810 54310
rect 115940 54300 116000 54310
rect 89000 54200 116000 54300
rect 89000 54190 89060 54200
rect 89190 54190 89310 54200
rect 89440 54190 89560 54200
rect 89690 54190 89810 54200
rect 89940 54190 90060 54200
rect 90190 54190 90310 54200
rect 90440 54190 90560 54200
rect 90690 54190 90810 54200
rect 90940 54190 91060 54200
rect 91190 54190 91310 54200
rect 91440 54190 91560 54200
rect 91690 54190 91810 54200
rect 91940 54190 92060 54200
rect 92190 54190 92310 54200
rect 92440 54190 92560 54200
rect 92690 54190 92810 54200
rect 92940 54190 93060 54200
rect 93190 54190 93310 54200
rect 93440 54190 93560 54200
rect 93690 54190 93810 54200
rect 93940 54190 94060 54200
rect 94190 54190 94310 54200
rect 94440 54190 94560 54200
rect 94690 54190 94810 54200
rect 94940 54190 95060 54200
rect 95190 54190 95310 54200
rect 95440 54190 95560 54200
rect 95690 54190 95810 54200
rect 95940 54190 96060 54200
rect 96190 54190 96310 54200
rect 96440 54190 96560 54200
rect 96690 54190 96810 54200
rect 96940 54190 97060 54200
rect 97190 54190 97310 54200
rect 97440 54190 97560 54200
rect 97690 54190 97810 54200
rect 97940 54190 98060 54200
rect 98190 54190 98310 54200
rect 98440 54190 98560 54200
rect 98690 54190 98810 54200
rect 98940 54190 99060 54200
rect 99190 54190 99310 54200
rect 99440 54190 99560 54200
rect 99690 54190 99810 54200
rect 99940 54190 100060 54200
rect 100190 54190 100310 54200
rect 100440 54190 100560 54200
rect 100690 54190 100810 54200
rect 100940 54190 101060 54200
rect 101190 54190 101310 54200
rect 101440 54190 101560 54200
rect 101690 54190 101810 54200
rect 101940 54190 102060 54200
rect 102190 54190 102310 54200
rect 102440 54190 102560 54200
rect 102690 54190 102810 54200
rect 102940 54190 103060 54200
rect 103190 54190 103310 54200
rect 103440 54190 103560 54200
rect 103690 54190 103810 54200
rect 103940 54190 104060 54200
rect 104190 54190 104310 54200
rect 104440 54190 104560 54200
rect 104690 54190 104810 54200
rect 104940 54190 105060 54200
rect 105190 54190 105310 54200
rect 105440 54190 105560 54200
rect 105690 54190 105810 54200
rect 105940 54190 106060 54200
rect 106190 54190 106310 54200
rect 106440 54190 106560 54200
rect 106690 54190 106810 54200
rect 106940 54190 107060 54200
rect 107190 54190 107310 54200
rect 107440 54190 107560 54200
rect 107690 54190 107810 54200
rect 107940 54190 108060 54200
rect 108190 54190 108310 54200
rect 108440 54190 108560 54200
rect 108690 54190 108810 54200
rect 108940 54190 109060 54200
rect 109190 54190 109310 54200
rect 109440 54190 109560 54200
rect 109690 54190 109810 54200
rect 109940 54190 110060 54200
rect 110190 54190 110310 54200
rect 110440 54190 110560 54200
rect 110690 54190 110810 54200
rect 110940 54190 111060 54200
rect 111190 54190 111310 54200
rect 111440 54190 111560 54200
rect 111690 54190 111810 54200
rect 111940 54190 112060 54200
rect 112190 54190 112310 54200
rect 112440 54190 112560 54200
rect 112690 54190 112810 54200
rect 112940 54190 113060 54200
rect 113190 54190 113310 54200
rect 113440 54190 113560 54200
rect 113690 54190 113810 54200
rect 113940 54190 114060 54200
rect 114190 54190 114310 54200
rect 114440 54190 114560 54200
rect 114690 54190 114810 54200
rect 114940 54190 115060 54200
rect 115190 54190 115310 54200
rect 115440 54190 115560 54200
rect 115690 54190 115810 54200
rect 115940 54190 116000 54200
rect 89000 54060 89050 54190
rect 89200 54060 89300 54190
rect 89450 54060 89550 54190
rect 89700 54060 89800 54190
rect 89950 54060 90050 54190
rect 90200 54060 90300 54190
rect 90450 54060 90550 54190
rect 90700 54060 90800 54190
rect 90950 54060 91050 54190
rect 91200 54060 91300 54190
rect 91450 54060 91550 54190
rect 91700 54060 91800 54190
rect 91950 54060 92050 54190
rect 92200 54060 92300 54190
rect 92450 54060 92550 54190
rect 92700 54060 92800 54190
rect 92950 54060 93050 54190
rect 93200 54060 93300 54190
rect 93450 54060 93550 54190
rect 93700 54060 93800 54190
rect 93950 54060 94050 54190
rect 94200 54060 94300 54190
rect 94450 54060 94550 54190
rect 94700 54060 94800 54190
rect 94950 54060 95050 54190
rect 95200 54060 95300 54190
rect 95450 54060 95550 54190
rect 95700 54060 95800 54190
rect 95950 54060 96050 54190
rect 96200 54060 96300 54190
rect 96450 54060 96550 54190
rect 96700 54060 96800 54190
rect 96950 54060 97050 54190
rect 97200 54060 97300 54190
rect 97450 54060 97550 54190
rect 97700 54060 97800 54190
rect 97950 54060 98050 54190
rect 98200 54060 98300 54190
rect 98450 54060 98550 54190
rect 98700 54060 98800 54190
rect 98950 54060 99050 54190
rect 99200 54060 99300 54190
rect 99450 54060 99550 54190
rect 99700 54060 99800 54190
rect 99950 54060 100050 54190
rect 100200 54060 100300 54190
rect 100450 54060 100550 54190
rect 100700 54060 100800 54190
rect 100950 54060 101050 54190
rect 101200 54060 101300 54190
rect 101450 54060 101550 54190
rect 101700 54060 101800 54190
rect 101950 54060 102050 54190
rect 102200 54060 102300 54190
rect 102450 54060 102550 54190
rect 102700 54060 102800 54190
rect 102950 54060 103050 54190
rect 103200 54060 103300 54190
rect 103450 54060 103550 54190
rect 103700 54060 103800 54190
rect 103950 54060 104050 54190
rect 104200 54060 104300 54190
rect 104450 54060 104550 54190
rect 104700 54060 104800 54190
rect 104950 54060 105050 54190
rect 105200 54060 105300 54190
rect 105450 54060 105550 54190
rect 105700 54060 105800 54190
rect 105950 54060 106050 54190
rect 106200 54060 106300 54190
rect 106450 54060 106550 54190
rect 106700 54060 106800 54190
rect 106950 54060 107050 54190
rect 107200 54060 107300 54190
rect 107450 54060 107550 54190
rect 107700 54060 107800 54190
rect 107950 54060 108050 54190
rect 108200 54060 108300 54190
rect 108450 54060 108550 54190
rect 108700 54060 108800 54190
rect 108950 54060 109050 54190
rect 109200 54060 109300 54190
rect 109450 54060 109550 54190
rect 109700 54060 109800 54190
rect 109950 54060 110050 54190
rect 110200 54060 110300 54190
rect 110450 54060 110550 54190
rect 110700 54060 110800 54190
rect 110950 54060 111050 54190
rect 111200 54060 111300 54190
rect 111450 54060 111550 54190
rect 111700 54060 111800 54190
rect 111950 54060 112050 54190
rect 112200 54060 112300 54190
rect 112450 54060 112550 54190
rect 112700 54060 112800 54190
rect 112950 54060 113050 54190
rect 113200 54060 113300 54190
rect 113450 54060 113550 54190
rect 113700 54060 113800 54190
rect 113950 54060 114050 54190
rect 114200 54060 114300 54190
rect 114450 54060 114550 54190
rect 114700 54060 114800 54190
rect 114950 54060 115050 54190
rect 115200 54060 115300 54190
rect 115450 54060 115550 54190
rect 115700 54060 115800 54190
rect 115950 54060 116000 54190
rect 89000 54050 89060 54060
rect 89190 54050 89310 54060
rect 89440 54050 89560 54060
rect 89690 54050 89810 54060
rect 89940 54050 90060 54060
rect 90190 54050 90310 54060
rect 90440 54050 90560 54060
rect 90690 54050 90810 54060
rect 90940 54050 91060 54060
rect 91190 54050 91310 54060
rect 91440 54050 91560 54060
rect 91690 54050 91810 54060
rect 91940 54050 92060 54060
rect 92190 54050 92310 54060
rect 92440 54050 92560 54060
rect 92690 54050 92810 54060
rect 92940 54050 93060 54060
rect 93190 54050 93310 54060
rect 93440 54050 93560 54060
rect 93690 54050 93810 54060
rect 93940 54050 94060 54060
rect 94190 54050 94310 54060
rect 94440 54050 94560 54060
rect 94690 54050 94810 54060
rect 94940 54050 95060 54060
rect 95190 54050 95310 54060
rect 95440 54050 95560 54060
rect 95690 54050 95810 54060
rect 95940 54050 96060 54060
rect 96190 54050 96310 54060
rect 96440 54050 96560 54060
rect 96690 54050 96810 54060
rect 96940 54050 97060 54060
rect 97190 54050 97310 54060
rect 97440 54050 97560 54060
rect 97690 54050 97810 54060
rect 97940 54050 98060 54060
rect 98190 54050 98310 54060
rect 98440 54050 98560 54060
rect 98690 54050 98810 54060
rect 98940 54050 99060 54060
rect 99190 54050 99310 54060
rect 99440 54050 99560 54060
rect 99690 54050 99810 54060
rect 99940 54050 100060 54060
rect 100190 54050 100310 54060
rect 100440 54050 100560 54060
rect 100690 54050 100810 54060
rect 100940 54050 101060 54060
rect 101190 54050 101310 54060
rect 101440 54050 101560 54060
rect 101690 54050 101810 54060
rect 101940 54050 102060 54060
rect 102190 54050 102310 54060
rect 102440 54050 102560 54060
rect 102690 54050 102810 54060
rect 102940 54050 103060 54060
rect 103190 54050 103310 54060
rect 103440 54050 103560 54060
rect 103690 54050 103810 54060
rect 103940 54050 104060 54060
rect 104190 54050 104310 54060
rect 104440 54050 104560 54060
rect 104690 54050 104810 54060
rect 104940 54050 105060 54060
rect 105190 54050 105310 54060
rect 105440 54050 105560 54060
rect 105690 54050 105810 54060
rect 105940 54050 106060 54060
rect 106190 54050 106310 54060
rect 106440 54050 106560 54060
rect 106690 54050 106810 54060
rect 106940 54050 107060 54060
rect 107190 54050 107310 54060
rect 107440 54050 107560 54060
rect 107690 54050 107810 54060
rect 107940 54050 108060 54060
rect 108190 54050 108310 54060
rect 108440 54050 108560 54060
rect 108690 54050 108810 54060
rect 108940 54050 109060 54060
rect 109190 54050 109310 54060
rect 109440 54050 109560 54060
rect 109690 54050 109810 54060
rect 109940 54050 110060 54060
rect 110190 54050 110310 54060
rect 110440 54050 110560 54060
rect 110690 54050 110810 54060
rect 110940 54050 111060 54060
rect 111190 54050 111310 54060
rect 111440 54050 111560 54060
rect 111690 54050 111810 54060
rect 111940 54050 112060 54060
rect 112190 54050 112310 54060
rect 112440 54050 112560 54060
rect 112690 54050 112810 54060
rect 112940 54050 113060 54060
rect 113190 54050 113310 54060
rect 113440 54050 113560 54060
rect 113690 54050 113810 54060
rect 113940 54050 114060 54060
rect 114190 54050 114310 54060
rect 114440 54050 114560 54060
rect 114690 54050 114810 54060
rect 114940 54050 115060 54060
rect 115190 54050 115310 54060
rect 115440 54050 115560 54060
rect 115690 54050 115810 54060
rect 115940 54050 116000 54060
rect 89000 53950 116000 54050
rect 89000 53940 89060 53950
rect 89190 53940 89310 53950
rect 89440 53940 89560 53950
rect 89690 53940 89810 53950
rect 89940 53940 90060 53950
rect 90190 53940 90310 53950
rect 90440 53940 90560 53950
rect 90690 53940 90810 53950
rect 90940 53940 91060 53950
rect 91190 53940 91310 53950
rect 91440 53940 91560 53950
rect 91690 53940 91810 53950
rect 91940 53940 92060 53950
rect 92190 53940 92310 53950
rect 92440 53940 92560 53950
rect 92690 53940 92810 53950
rect 92940 53940 93060 53950
rect 93190 53940 93310 53950
rect 93440 53940 93560 53950
rect 93690 53940 93810 53950
rect 93940 53940 94060 53950
rect 94190 53940 94310 53950
rect 94440 53940 94560 53950
rect 94690 53940 94810 53950
rect 94940 53940 95060 53950
rect 95190 53940 95310 53950
rect 95440 53940 95560 53950
rect 95690 53940 95810 53950
rect 95940 53940 96060 53950
rect 96190 53940 96310 53950
rect 96440 53940 96560 53950
rect 96690 53940 96810 53950
rect 96940 53940 97060 53950
rect 97190 53940 97310 53950
rect 97440 53940 97560 53950
rect 97690 53940 97810 53950
rect 97940 53940 98060 53950
rect 98190 53940 98310 53950
rect 98440 53940 98560 53950
rect 98690 53940 98810 53950
rect 98940 53940 99060 53950
rect 99190 53940 99310 53950
rect 99440 53940 99560 53950
rect 99690 53940 99810 53950
rect 99940 53940 100060 53950
rect 100190 53940 100310 53950
rect 100440 53940 100560 53950
rect 100690 53940 100810 53950
rect 100940 53940 101060 53950
rect 101190 53940 101310 53950
rect 101440 53940 101560 53950
rect 101690 53940 101810 53950
rect 101940 53940 102060 53950
rect 102190 53940 102310 53950
rect 102440 53940 102560 53950
rect 102690 53940 102810 53950
rect 102940 53940 103060 53950
rect 103190 53940 103310 53950
rect 103440 53940 103560 53950
rect 103690 53940 103810 53950
rect 103940 53940 104060 53950
rect 104190 53940 104310 53950
rect 104440 53940 104560 53950
rect 104690 53940 104810 53950
rect 104940 53940 105060 53950
rect 105190 53940 105310 53950
rect 105440 53940 105560 53950
rect 105690 53940 105810 53950
rect 105940 53940 106060 53950
rect 106190 53940 106310 53950
rect 106440 53940 106560 53950
rect 106690 53940 106810 53950
rect 106940 53940 107060 53950
rect 107190 53940 107310 53950
rect 107440 53940 107560 53950
rect 107690 53940 107810 53950
rect 107940 53940 108060 53950
rect 108190 53940 108310 53950
rect 108440 53940 108560 53950
rect 108690 53940 108810 53950
rect 108940 53940 109060 53950
rect 109190 53940 109310 53950
rect 109440 53940 109560 53950
rect 109690 53940 109810 53950
rect 109940 53940 110060 53950
rect 110190 53940 110310 53950
rect 110440 53940 110560 53950
rect 110690 53940 110810 53950
rect 110940 53940 111060 53950
rect 111190 53940 111310 53950
rect 111440 53940 111560 53950
rect 111690 53940 111810 53950
rect 111940 53940 112060 53950
rect 112190 53940 112310 53950
rect 112440 53940 112560 53950
rect 112690 53940 112810 53950
rect 112940 53940 113060 53950
rect 113190 53940 113310 53950
rect 113440 53940 113560 53950
rect 113690 53940 113810 53950
rect 113940 53940 114060 53950
rect 114190 53940 114310 53950
rect 114440 53940 114560 53950
rect 114690 53940 114810 53950
rect 114940 53940 115060 53950
rect 115190 53940 115310 53950
rect 115440 53940 115560 53950
rect 115690 53940 115810 53950
rect 115940 53940 116000 53950
rect 89000 53810 89050 53940
rect 89200 53810 89300 53940
rect 89450 53810 89550 53940
rect 89700 53810 89800 53940
rect 89950 53810 90050 53940
rect 90200 53810 90300 53940
rect 90450 53810 90550 53940
rect 90700 53810 90800 53940
rect 90950 53810 91050 53940
rect 91200 53810 91300 53940
rect 91450 53810 91550 53940
rect 91700 53810 91800 53940
rect 91950 53810 92050 53940
rect 92200 53810 92300 53940
rect 92450 53810 92550 53940
rect 92700 53810 92800 53940
rect 92950 53810 93050 53940
rect 93200 53810 93300 53940
rect 93450 53810 93550 53940
rect 93700 53810 93800 53940
rect 93950 53810 94050 53940
rect 94200 53810 94300 53940
rect 94450 53810 94550 53940
rect 94700 53810 94800 53940
rect 94950 53810 95050 53940
rect 95200 53810 95300 53940
rect 95450 53810 95550 53940
rect 95700 53810 95800 53940
rect 95950 53810 96050 53940
rect 96200 53810 96300 53940
rect 96450 53810 96550 53940
rect 96700 53810 96800 53940
rect 96950 53810 97050 53940
rect 97200 53810 97300 53940
rect 97450 53810 97550 53940
rect 97700 53810 97800 53940
rect 97950 53810 98050 53940
rect 98200 53810 98300 53940
rect 98450 53810 98550 53940
rect 98700 53810 98800 53940
rect 98950 53810 99050 53940
rect 99200 53810 99300 53940
rect 99450 53810 99550 53940
rect 99700 53810 99800 53940
rect 99950 53810 100050 53940
rect 100200 53810 100300 53940
rect 100450 53810 100550 53940
rect 100700 53810 100800 53940
rect 100950 53810 101050 53940
rect 101200 53810 101300 53940
rect 101450 53810 101550 53940
rect 101700 53810 101800 53940
rect 101950 53810 102050 53940
rect 102200 53810 102300 53940
rect 102450 53810 102550 53940
rect 102700 53810 102800 53940
rect 102950 53810 103050 53940
rect 103200 53810 103300 53940
rect 103450 53810 103550 53940
rect 103700 53810 103800 53940
rect 103950 53810 104050 53940
rect 104200 53810 104300 53940
rect 104450 53810 104550 53940
rect 104700 53810 104800 53940
rect 104950 53810 105050 53940
rect 105200 53810 105300 53940
rect 105450 53810 105550 53940
rect 105700 53810 105800 53940
rect 105950 53810 106050 53940
rect 106200 53810 106300 53940
rect 106450 53810 106550 53940
rect 106700 53810 106800 53940
rect 106950 53810 107050 53940
rect 107200 53810 107300 53940
rect 107450 53810 107550 53940
rect 107700 53810 107800 53940
rect 107950 53810 108050 53940
rect 108200 53810 108300 53940
rect 108450 53810 108550 53940
rect 108700 53810 108800 53940
rect 108950 53810 109050 53940
rect 109200 53810 109300 53940
rect 109450 53810 109550 53940
rect 109700 53810 109800 53940
rect 109950 53810 110050 53940
rect 110200 53810 110300 53940
rect 110450 53810 110550 53940
rect 110700 53810 110800 53940
rect 110950 53810 111050 53940
rect 111200 53810 111300 53940
rect 111450 53810 111550 53940
rect 111700 53810 111800 53940
rect 111950 53810 112050 53940
rect 112200 53810 112300 53940
rect 112450 53810 112550 53940
rect 112700 53810 112800 53940
rect 112950 53810 113050 53940
rect 113200 53810 113300 53940
rect 113450 53810 113550 53940
rect 113700 53810 113800 53940
rect 113950 53810 114050 53940
rect 114200 53810 114300 53940
rect 114450 53810 114550 53940
rect 114700 53810 114800 53940
rect 114950 53810 115050 53940
rect 115200 53810 115300 53940
rect 115450 53810 115550 53940
rect 115700 53810 115800 53940
rect 115950 53810 116000 53940
rect 89000 53800 89060 53810
rect 89190 53800 89310 53810
rect 89440 53800 89560 53810
rect 89690 53800 89810 53810
rect 89940 53800 90060 53810
rect 90190 53800 90310 53810
rect 90440 53800 90560 53810
rect 90690 53800 90810 53810
rect 90940 53800 91060 53810
rect 91190 53800 91310 53810
rect 91440 53800 91560 53810
rect 91690 53800 91810 53810
rect 91940 53800 92060 53810
rect 92190 53800 92310 53810
rect 92440 53800 92560 53810
rect 92690 53800 92810 53810
rect 92940 53800 93060 53810
rect 93190 53800 93310 53810
rect 93440 53800 93560 53810
rect 93690 53800 93810 53810
rect 93940 53800 94060 53810
rect 94190 53800 94310 53810
rect 94440 53800 94560 53810
rect 94690 53800 94810 53810
rect 94940 53800 95060 53810
rect 95190 53800 95310 53810
rect 95440 53800 95560 53810
rect 95690 53800 95810 53810
rect 95940 53800 96060 53810
rect 96190 53800 96310 53810
rect 96440 53800 96560 53810
rect 96690 53800 96810 53810
rect 96940 53800 97060 53810
rect 97190 53800 97310 53810
rect 97440 53800 97560 53810
rect 97690 53800 97810 53810
rect 97940 53800 98060 53810
rect 98190 53800 98310 53810
rect 98440 53800 98560 53810
rect 98690 53800 98810 53810
rect 98940 53800 99060 53810
rect 99190 53800 99310 53810
rect 99440 53800 99560 53810
rect 99690 53800 99810 53810
rect 99940 53800 100060 53810
rect 100190 53800 100310 53810
rect 100440 53800 100560 53810
rect 100690 53800 100810 53810
rect 100940 53800 101060 53810
rect 101190 53800 101310 53810
rect 101440 53800 101560 53810
rect 101690 53800 101810 53810
rect 101940 53800 102060 53810
rect 102190 53800 102310 53810
rect 102440 53800 102560 53810
rect 102690 53800 102810 53810
rect 102940 53800 103060 53810
rect 103190 53800 103310 53810
rect 103440 53800 103560 53810
rect 103690 53800 103810 53810
rect 103940 53800 104060 53810
rect 104190 53800 104310 53810
rect 104440 53800 104560 53810
rect 104690 53800 104810 53810
rect 104940 53800 105060 53810
rect 105190 53800 105310 53810
rect 105440 53800 105560 53810
rect 105690 53800 105810 53810
rect 105940 53800 106060 53810
rect 106190 53800 106310 53810
rect 106440 53800 106560 53810
rect 106690 53800 106810 53810
rect 106940 53800 107060 53810
rect 107190 53800 107310 53810
rect 107440 53800 107560 53810
rect 107690 53800 107810 53810
rect 107940 53800 108060 53810
rect 108190 53800 108310 53810
rect 108440 53800 108560 53810
rect 108690 53800 108810 53810
rect 108940 53800 109060 53810
rect 109190 53800 109310 53810
rect 109440 53800 109560 53810
rect 109690 53800 109810 53810
rect 109940 53800 110060 53810
rect 110190 53800 110310 53810
rect 110440 53800 110560 53810
rect 110690 53800 110810 53810
rect 110940 53800 111060 53810
rect 111190 53800 111310 53810
rect 111440 53800 111560 53810
rect 111690 53800 111810 53810
rect 111940 53800 112060 53810
rect 112190 53800 112310 53810
rect 112440 53800 112560 53810
rect 112690 53800 112810 53810
rect 112940 53800 113060 53810
rect 113190 53800 113310 53810
rect 113440 53800 113560 53810
rect 113690 53800 113810 53810
rect 113940 53800 114060 53810
rect 114190 53800 114310 53810
rect 114440 53800 114560 53810
rect 114690 53800 114810 53810
rect 114940 53800 115060 53810
rect 115190 53800 115310 53810
rect 115440 53800 115560 53810
rect 115690 53800 115810 53810
rect 115940 53800 116000 53810
rect 89000 53700 116000 53800
rect 89000 53690 89060 53700
rect 89190 53690 89310 53700
rect 89440 53690 89560 53700
rect 89690 53690 89810 53700
rect 89940 53690 90060 53700
rect 90190 53690 90310 53700
rect 90440 53690 90560 53700
rect 90690 53690 90810 53700
rect 90940 53690 91060 53700
rect 91190 53690 91310 53700
rect 91440 53690 91560 53700
rect 91690 53690 91810 53700
rect 91940 53690 92060 53700
rect 92190 53690 92310 53700
rect 92440 53690 92560 53700
rect 92690 53690 92810 53700
rect 92940 53690 93060 53700
rect 93190 53690 93310 53700
rect 93440 53690 93560 53700
rect 93690 53690 93810 53700
rect 93940 53690 94060 53700
rect 94190 53690 94310 53700
rect 94440 53690 94560 53700
rect 94690 53690 94810 53700
rect 94940 53690 95060 53700
rect 95190 53690 95310 53700
rect 95440 53690 95560 53700
rect 95690 53690 95810 53700
rect 95940 53690 96060 53700
rect 96190 53690 96310 53700
rect 96440 53690 96560 53700
rect 96690 53690 96810 53700
rect 96940 53690 97060 53700
rect 97190 53690 97310 53700
rect 97440 53690 97560 53700
rect 97690 53690 97810 53700
rect 97940 53690 98060 53700
rect 98190 53690 98310 53700
rect 98440 53690 98560 53700
rect 98690 53690 98810 53700
rect 98940 53690 99060 53700
rect 99190 53690 99310 53700
rect 99440 53690 99560 53700
rect 99690 53690 99810 53700
rect 99940 53690 100060 53700
rect 100190 53690 100310 53700
rect 100440 53690 100560 53700
rect 100690 53690 100810 53700
rect 100940 53690 101060 53700
rect 101190 53690 101310 53700
rect 101440 53690 101560 53700
rect 101690 53690 101810 53700
rect 101940 53690 102060 53700
rect 102190 53690 102310 53700
rect 102440 53690 102560 53700
rect 102690 53690 102810 53700
rect 102940 53690 103060 53700
rect 103190 53690 103310 53700
rect 103440 53690 103560 53700
rect 103690 53690 103810 53700
rect 103940 53690 104060 53700
rect 104190 53690 104310 53700
rect 104440 53690 104560 53700
rect 104690 53690 104810 53700
rect 104940 53690 105060 53700
rect 105190 53690 105310 53700
rect 105440 53690 105560 53700
rect 105690 53690 105810 53700
rect 105940 53690 106060 53700
rect 106190 53690 106310 53700
rect 106440 53690 106560 53700
rect 106690 53690 106810 53700
rect 106940 53690 107060 53700
rect 107190 53690 107310 53700
rect 107440 53690 107560 53700
rect 107690 53690 107810 53700
rect 107940 53690 108060 53700
rect 108190 53690 108310 53700
rect 108440 53690 108560 53700
rect 108690 53690 108810 53700
rect 108940 53690 109060 53700
rect 109190 53690 109310 53700
rect 109440 53690 109560 53700
rect 109690 53690 109810 53700
rect 109940 53690 110060 53700
rect 110190 53690 110310 53700
rect 110440 53690 110560 53700
rect 110690 53690 110810 53700
rect 110940 53690 111060 53700
rect 111190 53690 111310 53700
rect 111440 53690 111560 53700
rect 111690 53690 111810 53700
rect 111940 53690 112060 53700
rect 112190 53690 112310 53700
rect 112440 53690 112560 53700
rect 112690 53690 112810 53700
rect 112940 53690 113060 53700
rect 113190 53690 113310 53700
rect 113440 53690 113560 53700
rect 113690 53690 113810 53700
rect 113940 53690 114060 53700
rect 114190 53690 114310 53700
rect 114440 53690 114560 53700
rect 114690 53690 114810 53700
rect 114940 53690 115060 53700
rect 115190 53690 115310 53700
rect 115440 53690 115560 53700
rect 115690 53690 115810 53700
rect 115940 53690 116000 53700
rect 89000 53560 89050 53690
rect 89200 53560 89300 53690
rect 89450 53560 89550 53690
rect 89700 53560 89800 53690
rect 89950 53560 90050 53690
rect 90200 53560 90300 53690
rect 90450 53560 90550 53690
rect 90700 53560 90800 53690
rect 90950 53560 91050 53690
rect 91200 53560 91300 53690
rect 91450 53560 91550 53690
rect 91700 53560 91800 53690
rect 91950 53560 92050 53690
rect 92200 53560 92300 53690
rect 92450 53560 92550 53690
rect 92700 53560 92800 53690
rect 92950 53560 93050 53690
rect 93200 53560 93300 53690
rect 93450 53560 93550 53690
rect 93700 53560 93800 53690
rect 93950 53560 94050 53690
rect 94200 53560 94300 53690
rect 94450 53560 94550 53690
rect 94700 53560 94800 53690
rect 94950 53560 95050 53690
rect 95200 53560 95300 53690
rect 95450 53560 95550 53690
rect 95700 53560 95800 53690
rect 95950 53560 96050 53690
rect 96200 53560 96300 53690
rect 96450 53560 96550 53690
rect 96700 53560 96800 53690
rect 96950 53560 97050 53690
rect 97200 53560 97300 53690
rect 97450 53560 97550 53690
rect 97700 53560 97800 53690
rect 97950 53560 98050 53690
rect 98200 53560 98300 53690
rect 98450 53560 98550 53690
rect 98700 53560 98800 53690
rect 98950 53560 99050 53690
rect 99200 53560 99300 53690
rect 99450 53560 99550 53690
rect 99700 53560 99800 53690
rect 99950 53560 100050 53690
rect 100200 53560 100300 53690
rect 100450 53560 100550 53690
rect 100700 53560 100800 53690
rect 100950 53560 101050 53690
rect 101200 53560 101300 53690
rect 101450 53560 101550 53690
rect 101700 53560 101800 53690
rect 101950 53560 102050 53690
rect 102200 53560 102300 53690
rect 102450 53560 102550 53690
rect 102700 53560 102800 53690
rect 102950 53560 103050 53690
rect 103200 53560 103300 53690
rect 103450 53560 103550 53690
rect 103700 53560 103800 53690
rect 103950 53560 104050 53690
rect 104200 53560 104300 53690
rect 104450 53560 104550 53690
rect 104700 53560 104800 53690
rect 104950 53560 105050 53690
rect 105200 53560 105300 53690
rect 105450 53560 105550 53690
rect 105700 53560 105800 53690
rect 105950 53560 106050 53690
rect 106200 53560 106300 53690
rect 106450 53560 106550 53690
rect 106700 53560 106800 53690
rect 106950 53560 107050 53690
rect 107200 53560 107300 53690
rect 107450 53560 107550 53690
rect 107700 53560 107800 53690
rect 107950 53560 108050 53690
rect 108200 53560 108300 53690
rect 108450 53560 108550 53690
rect 108700 53560 108800 53690
rect 108950 53560 109050 53690
rect 109200 53560 109300 53690
rect 109450 53560 109550 53690
rect 109700 53560 109800 53690
rect 109950 53560 110050 53690
rect 110200 53560 110300 53690
rect 110450 53560 110550 53690
rect 110700 53560 110800 53690
rect 110950 53560 111050 53690
rect 111200 53560 111300 53690
rect 111450 53560 111550 53690
rect 111700 53560 111800 53690
rect 111950 53560 112050 53690
rect 112200 53560 112300 53690
rect 112450 53560 112550 53690
rect 112700 53560 112800 53690
rect 112950 53560 113050 53690
rect 113200 53560 113300 53690
rect 113450 53560 113550 53690
rect 113700 53560 113800 53690
rect 113950 53560 114050 53690
rect 114200 53560 114300 53690
rect 114450 53560 114550 53690
rect 114700 53560 114800 53690
rect 114950 53560 115050 53690
rect 115200 53560 115300 53690
rect 115450 53560 115550 53690
rect 115700 53560 115800 53690
rect 115950 53560 116000 53690
rect 89000 53550 89060 53560
rect 89190 53550 89310 53560
rect 89440 53550 89560 53560
rect 89690 53550 89810 53560
rect 89940 53550 90060 53560
rect 90190 53550 90310 53560
rect 90440 53550 90560 53560
rect 90690 53550 90810 53560
rect 90940 53550 91060 53560
rect 91190 53550 91310 53560
rect 91440 53550 91560 53560
rect 91690 53550 91810 53560
rect 91940 53550 92060 53560
rect 92190 53550 92310 53560
rect 92440 53550 92560 53560
rect 92690 53550 92810 53560
rect 92940 53550 93060 53560
rect 93190 53550 93310 53560
rect 93440 53550 93560 53560
rect 93690 53550 93810 53560
rect 93940 53550 94060 53560
rect 94190 53550 94310 53560
rect 94440 53550 94560 53560
rect 94690 53550 94810 53560
rect 94940 53550 95060 53560
rect 95190 53550 95310 53560
rect 95440 53550 95560 53560
rect 95690 53550 95810 53560
rect 95940 53550 96060 53560
rect 96190 53550 96310 53560
rect 96440 53550 96560 53560
rect 96690 53550 96810 53560
rect 96940 53550 97060 53560
rect 97190 53550 97310 53560
rect 97440 53550 97560 53560
rect 97690 53550 97810 53560
rect 97940 53550 98060 53560
rect 98190 53550 98310 53560
rect 98440 53550 98560 53560
rect 98690 53550 98810 53560
rect 98940 53550 99060 53560
rect 99190 53550 99310 53560
rect 99440 53550 99560 53560
rect 99690 53550 99810 53560
rect 99940 53550 100060 53560
rect 100190 53550 100310 53560
rect 100440 53550 100560 53560
rect 100690 53550 100810 53560
rect 100940 53550 101060 53560
rect 101190 53550 101310 53560
rect 101440 53550 101560 53560
rect 101690 53550 101810 53560
rect 101940 53550 102060 53560
rect 102190 53550 102310 53560
rect 102440 53550 102560 53560
rect 102690 53550 102810 53560
rect 102940 53550 103060 53560
rect 103190 53550 103310 53560
rect 103440 53550 103560 53560
rect 103690 53550 103810 53560
rect 103940 53550 104060 53560
rect 104190 53550 104310 53560
rect 104440 53550 104560 53560
rect 104690 53550 104810 53560
rect 104940 53550 105060 53560
rect 105190 53550 105310 53560
rect 105440 53550 105560 53560
rect 105690 53550 105810 53560
rect 105940 53550 106060 53560
rect 106190 53550 106310 53560
rect 106440 53550 106560 53560
rect 106690 53550 106810 53560
rect 106940 53550 107060 53560
rect 107190 53550 107310 53560
rect 107440 53550 107560 53560
rect 107690 53550 107810 53560
rect 107940 53550 108060 53560
rect 108190 53550 108310 53560
rect 108440 53550 108560 53560
rect 108690 53550 108810 53560
rect 108940 53550 109060 53560
rect 109190 53550 109310 53560
rect 109440 53550 109560 53560
rect 109690 53550 109810 53560
rect 109940 53550 110060 53560
rect 110190 53550 110310 53560
rect 110440 53550 110560 53560
rect 110690 53550 110810 53560
rect 110940 53550 111060 53560
rect 111190 53550 111310 53560
rect 111440 53550 111560 53560
rect 111690 53550 111810 53560
rect 111940 53550 112060 53560
rect 112190 53550 112310 53560
rect 112440 53550 112560 53560
rect 112690 53550 112810 53560
rect 112940 53550 113060 53560
rect 113190 53550 113310 53560
rect 113440 53550 113560 53560
rect 113690 53550 113810 53560
rect 113940 53550 114060 53560
rect 114190 53550 114310 53560
rect 114440 53550 114560 53560
rect 114690 53550 114810 53560
rect 114940 53550 115060 53560
rect 115190 53550 115310 53560
rect 115440 53550 115560 53560
rect 115690 53550 115810 53560
rect 115940 53550 116000 53560
rect 89000 53450 116000 53550
rect 89000 53440 89060 53450
rect 89190 53440 89310 53450
rect 89440 53440 89560 53450
rect 89690 53440 89810 53450
rect 89940 53440 90060 53450
rect 90190 53440 90310 53450
rect 90440 53440 90560 53450
rect 90690 53440 90810 53450
rect 90940 53440 91060 53450
rect 91190 53440 91310 53450
rect 91440 53440 91560 53450
rect 91690 53440 91810 53450
rect 91940 53440 92060 53450
rect 92190 53440 92310 53450
rect 92440 53440 92560 53450
rect 92690 53440 92810 53450
rect 92940 53440 93060 53450
rect 93190 53440 93310 53450
rect 93440 53440 93560 53450
rect 93690 53440 93810 53450
rect 93940 53440 94060 53450
rect 94190 53440 94310 53450
rect 94440 53440 94560 53450
rect 94690 53440 94810 53450
rect 94940 53440 95060 53450
rect 95190 53440 95310 53450
rect 95440 53440 95560 53450
rect 95690 53440 95810 53450
rect 95940 53440 96060 53450
rect 96190 53440 96310 53450
rect 96440 53440 96560 53450
rect 96690 53440 96810 53450
rect 96940 53440 97060 53450
rect 97190 53440 97310 53450
rect 97440 53440 97560 53450
rect 97690 53440 97810 53450
rect 97940 53440 98060 53450
rect 98190 53440 98310 53450
rect 98440 53440 98560 53450
rect 98690 53440 98810 53450
rect 98940 53440 99060 53450
rect 99190 53440 99310 53450
rect 99440 53440 99560 53450
rect 99690 53440 99810 53450
rect 99940 53440 100060 53450
rect 100190 53440 100310 53450
rect 100440 53440 100560 53450
rect 100690 53440 100810 53450
rect 100940 53440 101060 53450
rect 101190 53440 101310 53450
rect 101440 53440 101560 53450
rect 101690 53440 101810 53450
rect 101940 53440 102060 53450
rect 102190 53440 102310 53450
rect 102440 53440 102560 53450
rect 102690 53440 102810 53450
rect 102940 53440 103060 53450
rect 103190 53440 103310 53450
rect 103440 53440 103560 53450
rect 103690 53440 103810 53450
rect 103940 53440 104060 53450
rect 104190 53440 104310 53450
rect 104440 53440 104560 53450
rect 104690 53440 104810 53450
rect 104940 53440 105060 53450
rect 105190 53440 105310 53450
rect 105440 53440 105560 53450
rect 105690 53440 105810 53450
rect 105940 53440 106060 53450
rect 106190 53440 106310 53450
rect 106440 53440 106560 53450
rect 106690 53440 106810 53450
rect 106940 53440 107060 53450
rect 107190 53440 107310 53450
rect 107440 53440 107560 53450
rect 107690 53440 107810 53450
rect 107940 53440 108060 53450
rect 108190 53440 108310 53450
rect 108440 53440 108560 53450
rect 108690 53440 108810 53450
rect 108940 53440 109060 53450
rect 109190 53440 109310 53450
rect 109440 53440 109560 53450
rect 109690 53440 109810 53450
rect 109940 53440 110060 53450
rect 110190 53440 110310 53450
rect 110440 53440 110560 53450
rect 110690 53440 110810 53450
rect 110940 53440 111060 53450
rect 111190 53440 111310 53450
rect 111440 53440 111560 53450
rect 111690 53440 111810 53450
rect 111940 53440 112060 53450
rect 112190 53440 112310 53450
rect 112440 53440 112560 53450
rect 112690 53440 112810 53450
rect 112940 53440 113060 53450
rect 113190 53440 113310 53450
rect 113440 53440 113560 53450
rect 113690 53440 113810 53450
rect 113940 53440 114060 53450
rect 114190 53440 114310 53450
rect 114440 53440 114560 53450
rect 114690 53440 114810 53450
rect 114940 53440 115060 53450
rect 115190 53440 115310 53450
rect 115440 53440 115560 53450
rect 115690 53440 115810 53450
rect 115940 53440 116000 53450
rect 89000 53310 89050 53440
rect 89200 53310 89300 53440
rect 89450 53310 89550 53440
rect 89700 53310 89800 53440
rect 89950 53310 90050 53440
rect 90200 53310 90300 53440
rect 90450 53310 90550 53440
rect 90700 53310 90800 53440
rect 90950 53310 91050 53440
rect 91200 53310 91300 53440
rect 91450 53310 91550 53440
rect 91700 53310 91800 53440
rect 91950 53310 92050 53440
rect 92200 53310 92300 53440
rect 92450 53310 92550 53440
rect 92700 53310 92800 53440
rect 92950 53310 93050 53440
rect 93200 53310 93300 53440
rect 93450 53310 93550 53440
rect 93700 53310 93800 53440
rect 93950 53310 94050 53440
rect 94200 53310 94300 53440
rect 94450 53310 94550 53440
rect 94700 53310 94800 53440
rect 94950 53310 95050 53440
rect 95200 53310 95300 53440
rect 95450 53310 95550 53440
rect 95700 53310 95800 53440
rect 95950 53310 96050 53440
rect 96200 53310 96300 53440
rect 96450 53310 96550 53440
rect 96700 53310 96800 53440
rect 96950 53310 97050 53440
rect 97200 53310 97300 53440
rect 97450 53310 97550 53440
rect 97700 53310 97800 53440
rect 97950 53310 98050 53440
rect 98200 53310 98300 53440
rect 98450 53310 98550 53440
rect 98700 53310 98800 53440
rect 98950 53310 99050 53440
rect 99200 53310 99300 53440
rect 99450 53310 99550 53440
rect 99700 53310 99800 53440
rect 99950 53310 100050 53440
rect 100200 53310 100300 53440
rect 100450 53310 100550 53440
rect 100700 53310 100800 53440
rect 100950 53310 101050 53440
rect 101200 53310 101300 53440
rect 101450 53310 101550 53440
rect 101700 53310 101800 53440
rect 101950 53310 102050 53440
rect 102200 53310 102300 53440
rect 102450 53310 102550 53440
rect 102700 53310 102800 53440
rect 102950 53310 103050 53440
rect 103200 53310 103300 53440
rect 103450 53310 103550 53440
rect 103700 53310 103800 53440
rect 103950 53310 104050 53440
rect 104200 53310 104300 53440
rect 104450 53310 104550 53440
rect 104700 53310 104800 53440
rect 104950 53310 105050 53440
rect 105200 53310 105300 53440
rect 105450 53310 105550 53440
rect 105700 53310 105800 53440
rect 105950 53310 106050 53440
rect 106200 53310 106300 53440
rect 106450 53310 106550 53440
rect 106700 53310 106800 53440
rect 106950 53310 107050 53440
rect 107200 53310 107300 53440
rect 107450 53310 107550 53440
rect 107700 53310 107800 53440
rect 107950 53310 108050 53440
rect 108200 53310 108300 53440
rect 108450 53310 108550 53440
rect 108700 53310 108800 53440
rect 108950 53310 109050 53440
rect 109200 53310 109300 53440
rect 109450 53310 109550 53440
rect 109700 53310 109800 53440
rect 109950 53310 110050 53440
rect 110200 53310 110300 53440
rect 110450 53310 110550 53440
rect 110700 53310 110800 53440
rect 110950 53310 111050 53440
rect 111200 53310 111300 53440
rect 111450 53310 111550 53440
rect 111700 53310 111800 53440
rect 111950 53310 112050 53440
rect 112200 53310 112300 53440
rect 112450 53310 112550 53440
rect 112700 53310 112800 53440
rect 112950 53310 113050 53440
rect 113200 53310 113300 53440
rect 113450 53310 113550 53440
rect 113700 53310 113800 53440
rect 113950 53310 114050 53440
rect 114200 53310 114300 53440
rect 114450 53310 114550 53440
rect 114700 53310 114800 53440
rect 114950 53310 115050 53440
rect 115200 53310 115300 53440
rect 115450 53310 115550 53440
rect 115700 53310 115800 53440
rect 115950 53310 116000 53440
rect 89000 53300 89060 53310
rect 89190 53300 89310 53310
rect 89440 53300 89560 53310
rect 89690 53300 89810 53310
rect 89940 53300 90060 53310
rect 90190 53300 90310 53310
rect 90440 53300 90560 53310
rect 90690 53300 90810 53310
rect 90940 53300 91060 53310
rect 91190 53300 91310 53310
rect 91440 53300 91560 53310
rect 91690 53300 91810 53310
rect 91940 53300 92060 53310
rect 92190 53300 92310 53310
rect 92440 53300 92560 53310
rect 92690 53300 92810 53310
rect 92940 53300 93060 53310
rect 93190 53300 93310 53310
rect 93440 53300 93560 53310
rect 93690 53300 93810 53310
rect 93940 53300 94060 53310
rect 94190 53300 94310 53310
rect 94440 53300 94560 53310
rect 94690 53300 94810 53310
rect 94940 53300 95060 53310
rect 95190 53300 95310 53310
rect 95440 53300 95560 53310
rect 95690 53300 95810 53310
rect 95940 53300 96060 53310
rect 96190 53300 96310 53310
rect 96440 53300 96560 53310
rect 96690 53300 96810 53310
rect 96940 53300 97060 53310
rect 97190 53300 97310 53310
rect 97440 53300 97560 53310
rect 97690 53300 97810 53310
rect 97940 53300 98060 53310
rect 98190 53300 98310 53310
rect 98440 53300 98560 53310
rect 98690 53300 98810 53310
rect 98940 53300 99060 53310
rect 99190 53300 99310 53310
rect 99440 53300 99560 53310
rect 99690 53300 99810 53310
rect 99940 53300 100060 53310
rect 100190 53300 100310 53310
rect 100440 53300 100560 53310
rect 100690 53300 100810 53310
rect 100940 53300 101060 53310
rect 101190 53300 101310 53310
rect 101440 53300 101560 53310
rect 101690 53300 101810 53310
rect 101940 53300 102060 53310
rect 102190 53300 102310 53310
rect 102440 53300 102560 53310
rect 102690 53300 102810 53310
rect 102940 53300 103060 53310
rect 103190 53300 103310 53310
rect 103440 53300 103560 53310
rect 103690 53300 103810 53310
rect 103940 53300 104060 53310
rect 104190 53300 104310 53310
rect 104440 53300 104560 53310
rect 104690 53300 104810 53310
rect 104940 53300 105060 53310
rect 105190 53300 105310 53310
rect 105440 53300 105560 53310
rect 105690 53300 105810 53310
rect 105940 53300 106060 53310
rect 106190 53300 106310 53310
rect 106440 53300 106560 53310
rect 106690 53300 106810 53310
rect 106940 53300 107060 53310
rect 107190 53300 107310 53310
rect 107440 53300 107560 53310
rect 107690 53300 107810 53310
rect 107940 53300 108060 53310
rect 108190 53300 108310 53310
rect 108440 53300 108560 53310
rect 108690 53300 108810 53310
rect 108940 53300 109060 53310
rect 109190 53300 109310 53310
rect 109440 53300 109560 53310
rect 109690 53300 109810 53310
rect 109940 53300 110060 53310
rect 110190 53300 110310 53310
rect 110440 53300 110560 53310
rect 110690 53300 110810 53310
rect 110940 53300 111060 53310
rect 111190 53300 111310 53310
rect 111440 53300 111560 53310
rect 111690 53300 111810 53310
rect 111940 53300 112060 53310
rect 112190 53300 112310 53310
rect 112440 53300 112560 53310
rect 112690 53300 112810 53310
rect 112940 53300 113060 53310
rect 113190 53300 113310 53310
rect 113440 53300 113560 53310
rect 113690 53300 113810 53310
rect 113940 53300 114060 53310
rect 114190 53300 114310 53310
rect 114440 53300 114560 53310
rect 114690 53300 114810 53310
rect 114940 53300 115060 53310
rect 115190 53300 115310 53310
rect 115440 53300 115560 53310
rect 115690 53300 115810 53310
rect 115940 53300 116000 53310
rect 89000 53200 116000 53300
rect 89000 53190 89060 53200
rect 89190 53190 89310 53200
rect 89440 53190 89560 53200
rect 89690 53190 89810 53200
rect 89940 53190 90060 53200
rect 90190 53190 90310 53200
rect 90440 53190 90560 53200
rect 90690 53190 90810 53200
rect 90940 53190 91060 53200
rect 91190 53190 91310 53200
rect 91440 53190 91560 53200
rect 91690 53190 91810 53200
rect 91940 53190 92060 53200
rect 92190 53190 92310 53200
rect 92440 53190 92560 53200
rect 92690 53190 92810 53200
rect 92940 53190 93060 53200
rect 93190 53190 93310 53200
rect 93440 53190 93560 53200
rect 93690 53190 93810 53200
rect 93940 53190 94060 53200
rect 94190 53190 94310 53200
rect 94440 53190 94560 53200
rect 94690 53190 94810 53200
rect 94940 53190 95060 53200
rect 95190 53190 95310 53200
rect 95440 53190 95560 53200
rect 95690 53190 95810 53200
rect 95940 53190 96060 53200
rect 96190 53190 96310 53200
rect 96440 53190 96560 53200
rect 96690 53190 96810 53200
rect 96940 53190 97060 53200
rect 97190 53190 97310 53200
rect 97440 53190 97560 53200
rect 97690 53190 97810 53200
rect 97940 53190 98060 53200
rect 98190 53190 98310 53200
rect 98440 53190 98560 53200
rect 98690 53190 98810 53200
rect 98940 53190 99060 53200
rect 99190 53190 99310 53200
rect 99440 53190 99560 53200
rect 99690 53190 99810 53200
rect 99940 53190 100060 53200
rect 100190 53190 100310 53200
rect 100440 53190 100560 53200
rect 100690 53190 100810 53200
rect 100940 53190 101060 53200
rect 101190 53190 101310 53200
rect 101440 53190 101560 53200
rect 101690 53190 101810 53200
rect 101940 53190 102060 53200
rect 102190 53190 102310 53200
rect 102440 53190 102560 53200
rect 102690 53190 102810 53200
rect 102940 53190 103060 53200
rect 103190 53190 103310 53200
rect 103440 53190 103560 53200
rect 103690 53190 103810 53200
rect 103940 53190 104060 53200
rect 104190 53190 104310 53200
rect 104440 53190 104560 53200
rect 104690 53190 104810 53200
rect 104940 53190 105060 53200
rect 105190 53190 105310 53200
rect 105440 53190 105560 53200
rect 105690 53190 105810 53200
rect 105940 53190 106060 53200
rect 106190 53190 106310 53200
rect 106440 53190 106560 53200
rect 106690 53190 106810 53200
rect 106940 53190 107060 53200
rect 107190 53190 107310 53200
rect 107440 53190 107560 53200
rect 107690 53190 107810 53200
rect 107940 53190 108060 53200
rect 108190 53190 108310 53200
rect 108440 53190 108560 53200
rect 108690 53190 108810 53200
rect 108940 53190 109060 53200
rect 109190 53190 109310 53200
rect 109440 53190 109560 53200
rect 109690 53190 109810 53200
rect 109940 53190 110060 53200
rect 110190 53190 110310 53200
rect 110440 53190 110560 53200
rect 110690 53190 110810 53200
rect 110940 53190 111060 53200
rect 111190 53190 111310 53200
rect 111440 53190 111560 53200
rect 111690 53190 111810 53200
rect 111940 53190 112060 53200
rect 112190 53190 112310 53200
rect 112440 53190 112560 53200
rect 112690 53190 112810 53200
rect 112940 53190 113060 53200
rect 113190 53190 113310 53200
rect 113440 53190 113560 53200
rect 113690 53190 113810 53200
rect 113940 53190 114060 53200
rect 114190 53190 114310 53200
rect 114440 53190 114560 53200
rect 114690 53190 114810 53200
rect 114940 53190 115060 53200
rect 115190 53190 115310 53200
rect 115440 53190 115560 53200
rect 115690 53190 115810 53200
rect 115940 53190 116000 53200
rect 89000 53060 89050 53190
rect 89200 53060 89300 53190
rect 89450 53060 89550 53190
rect 89700 53060 89800 53190
rect 89950 53060 90050 53190
rect 90200 53060 90300 53190
rect 90450 53060 90550 53190
rect 90700 53060 90800 53190
rect 90950 53060 91050 53190
rect 91200 53060 91300 53190
rect 91450 53060 91550 53190
rect 91700 53060 91800 53190
rect 91950 53060 92050 53190
rect 92200 53060 92300 53190
rect 92450 53060 92550 53190
rect 92700 53060 92800 53190
rect 92950 53060 93050 53190
rect 93200 53060 93300 53190
rect 93450 53060 93550 53190
rect 93700 53060 93800 53190
rect 93950 53060 94050 53190
rect 94200 53060 94300 53190
rect 94450 53060 94550 53190
rect 94700 53060 94800 53190
rect 94950 53060 95050 53190
rect 95200 53060 95300 53190
rect 95450 53060 95550 53190
rect 95700 53060 95800 53190
rect 95950 53060 96050 53190
rect 96200 53060 96300 53190
rect 96450 53060 96550 53190
rect 96700 53060 96800 53190
rect 96950 53060 97050 53190
rect 97200 53060 97300 53190
rect 97450 53060 97550 53190
rect 97700 53060 97800 53190
rect 97950 53060 98050 53190
rect 98200 53060 98300 53190
rect 98450 53060 98550 53190
rect 98700 53060 98800 53190
rect 98950 53060 99050 53190
rect 99200 53060 99300 53190
rect 99450 53060 99550 53190
rect 99700 53060 99800 53190
rect 99950 53060 100050 53190
rect 100200 53060 100300 53190
rect 100450 53060 100550 53190
rect 100700 53060 100800 53190
rect 100950 53060 101050 53190
rect 101200 53060 101300 53190
rect 101450 53060 101550 53190
rect 101700 53060 101800 53190
rect 101950 53060 102050 53190
rect 102200 53060 102300 53190
rect 102450 53060 102550 53190
rect 102700 53060 102800 53190
rect 102950 53060 103050 53190
rect 103200 53060 103300 53190
rect 103450 53060 103550 53190
rect 103700 53060 103800 53190
rect 103950 53060 104050 53190
rect 104200 53060 104300 53190
rect 104450 53060 104550 53190
rect 104700 53060 104800 53190
rect 104950 53060 105050 53190
rect 105200 53060 105300 53190
rect 105450 53060 105550 53190
rect 105700 53060 105800 53190
rect 105950 53060 106050 53190
rect 106200 53060 106300 53190
rect 106450 53060 106550 53190
rect 106700 53060 106800 53190
rect 106950 53060 107050 53190
rect 107200 53060 107300 53190
rect 107450 53060 107550 53190
rect 107700 53060 107800 53190
rect 107950 53060 108050 53190
rect 108200 53060 108300 53190
rect 108450 53060 108550 53190
rect 108700 53060 108800 53190
rect 108950 53060 109050 53190
rect 109200 53060 109300 53190
rect 109450 53060 109550 53190
rect 109700 53060 109800 53190
rect 109950 53060 110050 53190
rect 110200 53060 110300 53190
rect 110450 53060 110550 53190
rect 110700 53060 110800 53190
rect 110950 53060 111050 53190
rect 111200 53060 111300 53190
rect 111450 53060 111550 53190
rect 111700 53060 111800 53190
rect 111950 53060 112050 53190
rect 112200 53060 112300 53190
rect 112450 53060 112550 53190
rect 112700 53060 112800 53190
rect 112950 53060 113050 53190
rect 113200 53060 113300 53190
rect 113450 53060 113550 53190
rect 113700 53060 113800 53190
rect 113950 53060 114050 53190
rect 114200 53060 114300 53190
rect 114450 53060 114550 53190
rect 114700 53060 114800 53190
rect 114950 53060 115050 53190
rect 115200 53060 115300 53190
rect 115450 53060 115550 53190
rect 115700 53060 115800 53190
rect 115950 53060 116000 53190
rect 89000 53050 89060 53060
rect 89190 53050 89310 53060
rect 89440 53050 89560 53060
rect 89690 53050 89810 53060
rect 89940 53050 90060 53060
rect 90190 53050 90310 53060
rect 90440 53050 90560 53060
rect 90690 53050 90810 53060
rect 90940 53050 91060 53060
rect 91190 53050 91310 53060
rect 91440 53050 91560 53060
rect 91690 53050 91810 53060
rect 91940 53050 92060 53060
rect 92190 53050 92310 53060
rect 92440 53050 92560 53060
rect 92690 53050 92810 53060
rect 92940 53050 93060 53060
rect 93190 53050 93310 53060
rect 93440 53050 93560 53060
rect 93690 53050 93810 53060
rect 93940 53050 94060 53060
rect 94190 53050 94310 53060
rect 94440 53050 94560 53060
rect 94690 53050 94810 53060
rect 94940 53050 95060 53060
rect 95190 53050 95310 53060
rect 95440 53050 95560 53060
rect 95690 53050 95810 53060
rect 95940 53050 96060 53060
rect 96190 53050 96310 53060
rect 96440 53050 96560 53060
rect 96690 53050 96810 53060
rect 96940 53050 97060 53060
rect 97190 53050 97310 53060
rect 97440 53050 97560 53060
rect 97690 53050 97810 53060
rect 97940 53050 98060 53060
rect 98190 53050 98310 53060
rect 98440 53050 98560 53060
rect 98690 53050 98810 53060
rect 98940 53050 99060 53060
rect 99190 53050 99310 53060
rect 99440 53050 99560 53060
rect 99690 53050 99810 53060
rect 99940 53050 100060 53060
rect 100190 53050 100310 53060
rect 100440 53050 100560 53060
rect 100690 53050 100810 53060
rect 100940 53050 101060 53060
rect 101190 53050 101310 53060
rect 101440 53050 101560 53060
rect 101690 53050 101810 53060
rect 101940 53050 102060 53060
rect 102190 53050 102310 53060
rect 102440 53050 102560 53060
rect 102690 53050 102810 53060
rect 102940 53050 103060 53060
rect 103190 53050 103310 53060
rect 103440 53050 103560 53060
rect 103690 53050 103810 53060
rect 103940 53050 104060 53060
rect 104190 53050 104310 53060
rect 104440 53050 104560 53060
rect 104690 53050 104810 53060
rect 104940 53050 105060 53060
rect 105190 53050 105310 53060
rect 105440 53050 105560 53060
rect 105690 53050 105810 53060
rect 105940 53050 106060 53060
rect 106190 53050 106310 53060
rect 106440 53050 106560 53060
rect 106690 53050 106810 53060
rect 106940 53050 107060 53060
rect 107190 53050 107310 53060
rect 107440 53050 107560 53060
rect 107690 53050 107810 53060
rect 107940 53050 108060 53060
rect 108190 53050 108310 53060
rect 108440 53050 108560 53060
rect 108690 53050 108810 53060
rect 108940 53050 109060 53060
rect 109190 53050 109310 53060
rect 109440 53050 109560 53060
rect 109690 53050 109810 53060
rect 109940 53050 110060 53060
rect 110190 53050 110310 53060
rect 110440 53050 110560 53060
rect 110690 53050 110810 53060
rect 110940 53050 111060 53060
rect 111190 53050 111310 53060
rect 111440 53050 111560 53060
rect 111690 53050 111810 53060
rect 111940 53050 112060 53060
rect 112190 53050 112310 53060
rect 112440 53050 112560 53060
rect 112690 53050 112810 53060
rect 112940 53050 113060 53060
rect 113190 53050 113310 53060
rect 113440 53050 113560 53060
rect 113690 53050 113810 53060
rect 113940 53050 114060 53060
rect 114190 53050 114310 53060
rect 114440 53050 114560 53060
rect 114690 53050 114810 53060
rect 114940 53050 115060 53060
rect 115190 53050 115310 53060
rect 115440 53050 115560 53060
rect 115690 53050 115810 53060
rect 115940 53050 116000 53060
rect 89000 52950 116000 53050
rect 89000 52940 89060 52950
rect 89190 52940 89310 52950
rect 89440 52940 89560 52950
rect 89690 52940 89810 52950
rect 89940 52940 90060 52950
rect 90190 52940 90310 52950
rect 90440 52940 90560 52950
rect 90690 52940 90810 52950
rect 90940 52940 91060 52950
rect 91190 52940 91310 52950
rect 91440 52940 91560 52950
rect 91690 52940 91810 52950
rect 91940 52940 92060 52950
rect 92190 52940 92310 52950
rect 92440 52940 92560 52950
rect 92690 52940 92810 52950
rect 92940 52940 93060 52950
rect 93190 52940 93310 52950
rect 93440 52940 93560 52950
rect 93690 52940 93810 52950
rect 93940 52940 94060 52950
rect 94190 52940 94310 52950
rect 94440 52940 94560 52950
rect 94690 52940 94810 52950
rect 94940 52940 95060 52950
rect 95190 52940 95310 52950
rect 95440 52940 95560 52950
rect 95690 52940 95810 52950
rect 95940 52940 96060 52950
rect 96190 52940 96310 52950
rect 96440 52940 96560 52950
rect 96690 52940 96810 52950
rect 96940 52940 97060 52950
rect 97190 52940 97310 52950
rect 97440 52940 97560 52950
rect 97690 52940 97810 52950
rect 97940 52940 98060 52950
rect 98190 52940 98310 52950
rect 98440 52940 98560 52950
rect 98690 52940 98810 52950
rect 98940 52940 99060 52950
rect 99190 52940 99310 52950
rect 99440 52940 99560 52950
rect 99690 52940 99810 52950
rect 99940 52940 100060 52950
rect 100190 52940 100310 52950
rect 100440 52940 100560 52950
rect 100690 52940 100810 52950
rect 100940 52940 101060 52950
rect 101190 52940 101310 52950
rect 101440 52940 101560 52950
rect 101690 52940 101810 52950
rect 101940 52940 102060 52950
rect 102190 52940 102310 52950
rect 102440 52940 102560 52950
rect 102690 52940 102810 52950
rect 102940 52940 103060 52950
rect 103190 52940 103310 52950
rect 103440 52940 103560 52950
rect 103690 52940 103810 52950
rect 103940 52940 104060 52950
rect 104190 52940 104310 52950
rect 104440 52940 104560 52950
rect 104690 52940 104810 52950
rect 104940 52940 105060 52950
rect 105190 52940 105310 52950
rect 105440 52940 105560 52950
rect 105690 52940 105810 52950
rect 105940 52940 106060 52950
rect 106190 52940 106310 52950
rect 106440 52940 106560 52950
rect 106690 52940 106810 52950
rect 106940 52940 107060 52950
rect 107190 52940 107310 52950
rect 107440 52940 107560 52950
rect 107690 52940 107810 52950
rect 107940 52940 108060 52950
rect 108190 52940 108310 52950
rect 108440 52940 108560 52950
rect 108690 52940 108810 52950
rect 108940 52940 109060 52950
rect 109190 52940 109310 52950
rect 109440 52940 109560 52950
rect 109690 52940 109810 52950
rect 109940 52940 110060 52950
rect 110190 52940 110310 52950
rect 110440 52940 110560 52950
rect 110690 52940 110810 52950
rect 110940 52940 111060 52950
rect 111190 52940 111310 52950
rect 111440 52940 111560 52950
rect 111690 52940 111810 52950
rect 111940 52940 112060 52950
rect 112190 52940 112310 52950
rect 112440 52940 112560 52950
rect 112690 52940 112810 52950
rect 112940 52940 113060 52950
rect 113190 52940 113310 52950
rect 113440 52940 113560 52950
rect 113690 52940 113810 52950
rect 113940 52940 114060 52950
rect 114190 52940 114310 52950
rect 114440 52940 114560 52950
rect 114690 52940 114810 52950
rect 114940 52940 115060 52950
rect 115190 52940 115310 52950
rect 115440 52940 115560 52950
rect 115690 52940 115810 52950
rect 115940 52940 116000 52950
rect 89000 52810 89050 52940
rect 89200 52810 89300 52940
rect 89450 52810 89550 52940
rect 89700 52810 89800 52940
rect 89950 52810 90050 52940
rect 90200 52810 90300 52940
rect 90450 52810 90550 52940
rect 90700 52810 90800 52940
rect 90950 52810 91050 52940
rect 91200 52810 91300 52940
rect 91450 52810 91550 52940
rect 91700 52810 91800 52940
rect 91950 52810 92050 52940
rect 92200 52810 92300 52940
rect 92450 52810 92550 52940
rect 92700 52810 92800 52940
rect 92950 52810 93050 52940
rect 93200 52810 93300 52940
rect 93450 52810 93550 52940
rect 93700 52810 93800 52940
rect 93950 52810 94050 52940
rect 94200 52810 94300 52940
rect 94450 52810 94550 52940
rect 94700 52810 94800 52940
rect 94950 52810 95050 52940
rect 95200 52810 95300 52940
rect 95450 52810 95550 52940
rect 95700 52810 95800 52940
rect 95950 52810 96050 52940
rect 96200 52810 96300 52940
rect 96450 52810 96550 52940
rect 96700 52810 96800 52940
rect 96950 52810 97050 52940
rect 97200 52810 97300 52940
rect 97450 52810 97550 52940
rect 97700 52810 97800 52940
rect 97950 52810 98050 52940
rect 98200 52810 98300 52940
rect 98450 52810 98550 52940
rect 98700 52810 98800 52940
rect 98950 52810 99050 52940
rect 99200 52810 99300 52940
rect 99450 52810 99550 52940
rect 99700 52810 99800 52940
rect 99950 52810 100050 52940
rect 100200 52810 100300 52940
rect 100450 52810 100550 52940
rect 100700 52810 100800 52940
rect 100950 52810 101050 52940
rect 101200 52810 101300 52940
rect 101450 52810 101550 52940
rect 101700 52810 101800 52940
rect 101950 52810 102050 52940
rect 102200 52810 102300 52940
rect 102450 52810 102550 52940
rect 102700 52810 102800 52940
rect 102950 52810 103050 52940
rect 103200 52810 103300 52940
rect 103450 52810 103550 52940
rect 103700 52810 103800 52940
rect 103950 52810 104050 52940
rect 104200 52810 104300 52940
rect 104450 52810 104550 52940
rect 104700 52810 104800 52940
rect 104950 52810 105050 52940
rect 105200 52810 105300 52940
rect 105450 52810 105550 52940
rect 105700 52810 105800 52940
rect 105950 52810 106050 52940
rect 106200 52810 106300 52940
rect 106450 52810 106550 52940
rect 106700 52810 106800 52940
rect 106950 52810 107050 52940
rect 107200 52810 107300 52940
rect 107450 52810 107550 52940
rect 107700 52810 107800 52940
rect 107950 52810 108050 52940
rect 108200 52810 108300 52940
rect 108450 52810 108550 52940
rect 108700 52810 108800 52940
rect 108950 52810 109050 52940
rect 109200 52810 109300 52940
rect 109450 52810 109550 52940
rect 109700 52810 109800 52940
rect 109950 52810 110050 52940
rect 110200 52810 110300 52940
rect 110450 52810 110550 52940
rect 110700 52810 110800 52940
rect 110950 52810 111050 52940
rect 111200 52810 111300 52940
rect 111450 52810 111550 52940
rect 111700 52810 111800 52940
rect 111950 52810 112050 52940
rect 112200 52810 112300 52940
rect 112450 52810 112550 52940
rect 112700 52810 112800 52940
rect 112950 52810 113050 52940
rect 113200 52810 113300 52940
rect 113450 52810 113550 52940
rect 113700 52810 113800 52940
rect 113950 52810 114050 52940
rect 114200 52810 114300 52940
rect 114450 52810 114550 52940
rect 114700 52810 114800 52940
rect 114950 52810 115050 52940
rect 115200 52810 115300 52940
rect 115450 52810 115550 52940
rect 115700 52810 115800 52940
rect 115950 52810 116000 52940
rect 89000 52800 89060 52810
rect 89190 52800 89310 52810
rect 89440 52800 89560 52810
rect 89690 52800 89810 52810
rect 89940 52800 90060 52810
rect 90190 52800 90310 52810
rect 90440 52800 90560 52810
rect 90690 52800 90810 52810
rect 90940 52800 91060 52810
rect 91190 52800 91310 52810
rect 91440 52800 91560 52810
rect 91690 52800 91810 52810
rect 91940 52800 92060 52810
rect 92190 52800 92310 52810
rect 92440 52800 92560 52810
rect 92690 52800 92810 52810
rect 92940 52800 93060 52810
rect 93190 52800 93310 52810
rect 93440 52800 93560 52810
rect 93690 52800 93810 52810
rect 93940 52800 94060 52810
rect 94190 52800 94310 52810
rect 94440 52800 94560 52810
rect 94690 52800 94810 52810
rect 94940 52800 95060 52810
rect 95190 52800 95310 52810
rect 95440 52800 95560 52810
rect 95690 52800 95810 52810
rect 95940 52800 96060 52810
rect 96190 52800 96310 52810
rect 96440 52800 96560 52810
rect 96690 52800 96810 52810
rect 96940 52800 97060 52810
rect 97190 52800 97310 52810
rect 97440 52800 97560 52810
rect 97690 52800 97810 52810
rect 97940 52800 98060 52810
rect 98190 52800 98310 52810
rect 98440 52800 98560 52810
rect 98690 52800 98810 52810
rect 98940 52800 99060 52810
rect 99190 52800 99310 52810
rect 99440 52800 99560 52810
rect 99690 52800 99810 52810
rect 99940 52800 100060 52810
rect 100190 52800 100310 52810
rect 100440 52800 100560 52810
rect 100690 52800 100810 52810
rect 100940 52800 101060 52810
rect 101190 52800 101310 52810
rect 101440 52800 101560 52810
rect 101690 52800 101810 52810
rect 101940 52800 102060 52810
rect 102190 52800 102310 52810
rect 102440 52800 102560 52810
rect 102690 52800 102810 52810
rect 102940 52800 103060 52810
rect 103190 52800 103310 52810
rect 103440 52800 103560 52810
rect 103690 52800 103810 52810
rect 103940 52800 104060 52810
rect 104190 52800 104310 52810
rect 104440 52800 104560 52810
rect 104690 52800 104810 52810
rect 104940 52800 105060 52810
rect 105190 52800 105310 52810
rect 105440 52800 105560 52810
rect 105690 52800 105810 52810
rect 105940 52800 106060 52810
rect 106190 52800 106310 52810
rect 106440 52800 106560 52810
rect 106690 52800 106810 52810
rect 106940 52800 107060 52810
rect 107190 52800 107310 52810
rect 107440 52800 107560 52810
rect 107690 52800 107810 52810
rect 107940 52800 108060 52810
rect 108190 52800 108310 52810
rect 108440 52800 108560 52810
rect 108690 52800 108810 52810
rect 108940 52800 109060 52810
rect 109190 52800 109310 52810
rect 109440 52800 109560 52810
rect 109690 52800 109810 52810
rect 109940 52800 110060 52810
rect 110190 52800 110310 52810
rect 110440 52800 110560 52810
rect 110690 52800 110810 52810
rect 110940 52800 111060 52810
rect 111190 52800 111310 52810
rect 111440 52800 111560 52810
rect 111690 52800 111810 52810
rect 111940 52800 112060 52810
rect 112190 52800 112310 52810
rect 112440 52800 112560 52810
rect 112690 52800 112810 52810
rect 112940 52800 113060 52810
rect 113190 52800 113310 52810
rect 113440 52800 113560 52810
rect 113690 52800 113810 52810
rect 113940 52800 114060 52810
rect 114190 52800 114310 52810
rect 114440 52800 114560 52810
rect 114690 52800 114810 52810
rect 114940 52800 115060 52810
rect 115190 52800 115310 52810
rect 115440 52800 115560 52810
rect 115690 52800 115810 52810
rect 115940 52800 116000 52810
rect 89000 52700 116000 52800
rect 89000 52690 89060 52700
rect 89190 52690 89310 52700
rect 89440 52690 89560 52700
rect 89690 52690 89810 52700
rect 89940 52690 90060 52700
rect 90190 52690 90310 52700
rect 90440 52690 90560 52700
rect 90690 52690 90810 52700
rect 90940 52690 91060 52700
rect 91190 52690 91310 52700
rect 91440 52690 91560 52700
rect 91690 52690 91810 52700
rect 91940 52690 92060 52700
rect 92190 52690 92310 52700
rect 92440 52690 92560 52700
rect 92690 52690 92810 52700
rect 92940 52690 93060 52700
rect 93190 52690 93310 52700
rect 93440 52690 93560 52700
rect 93690 52690 93810 52700
rect 93940 52690 94060 52700
rect 94190 52690 94310 52700
rect 94440 52690 94560 52700
rect 94690 52690 94810 52700
rect 94940 52690 95060 52700
rect 95190 52690 95310 52700
rect 95440 52690 95560 52700
rect 95690 52690 95810 52700
rect 95940 52690 96060 52700
rect 96190 52690 96310 52700
rect 96440 52690 96560 52700
rect 96690 52690 96810 52700
rect 96940 52690 97060 52700
rect 97190 52690 97310 52700
rect 97440 52690 97560 52700
rect 97690 52690 97810 52700
rect 97940 52690 98060 52700
rect 98190 52690 98310 52700
rect 98440 52690 98560 52700
rect 98690 52690 98810 52700
rect 98940 52690 99060 52700
rect 99190 52690 99310 52700
rect 99440 52690 99560 52700
rect 99690 52690 99810 52700
rect 99940 52690 100060 52700
rect 100190 52690 100310 52700
rect 100440 52690 100560 52700
rect 100690 52690 100810 52700
rect 100940 52690 101060 52700
rect 101190 52690 101310 52700
rect 101440 52690 101560 52700
rect 101690 52690 101810 52700
rect 101940 52690 102060 52700
rect 102190 52690 102310 52700
rect 102440 52690 102560 52700
rect 102690 52690 102810 52700
rect 102940 52690 103060 52700
rect 103190 52690 103310 52700
rect 103440 52690 103560 52700
rect 103690 52690 103810 52700
rect 103940 52690 104060 52700
rect 104190 52690 104310 52700
rect 104440 52690 104560 52700
rect 104690 52690 104810 52700
rect 104940 52690 105060 52700
rect 105190 52690 105310 52700
rect 105440 52690 105560 52700
rect 105690 52690 105810 52700
rect 105940 52690 106060 52700
rect 106190 52690 106310 52700
rect 106440 52690 106560 52700
rect 106690 52690 106810 52700
rect 106940 52690 107060 52700
rect 107190 52690 107310 52700
rect 107440 52690 107560 52700
rect 107690 52690 107810 52700
rect 107940 52690 108060 52700
rect 108190 52690 108310 52700
rect 108440 52690 108560 52700
rect 108690 52690 108810 52700
rect 108940 52690 109060 52700
rect 109190 52690 109310 52700
rect 109440 52690 109560 52700
rect 109690 52690 109810 52700
rect 109940 52690 110060 52700
rect 110190 52690 110310 52700
rect 110440 52690 110560 52700
rect 110690 52690 110810 52700
rect 110940 52690 111060 52700
rect 111190 52690 111310 52700
rect 111440 52690 111560 52700
rect 111690 52690 111810 52700
rect 111940 52690 112060 52700
rect 112190 52690 112310 52700
rect 112440 52690 112560 52700
rect 112690 52690 112810 52700
rect 112940 52690 113060 52700
rect 113190 52690 113310 52700
rect 113440 52690 113560 52700
rect 113690 52690 113810 52700
rect 113940 52690 114060 52700
rect 114190 52690 114310 52700
rect 114440 52690 114560 52700
rect 114690 52690 114810 52700
rect 114940 52690 115060 52700
rect 115190 52690 115310 52700
rect 115440 52690 115560 52700
rect 115690 52690 115810 52700
rect 115940 52690 116000 52700
rect 89000 52560 89050 52690
rect 89200 52560 89300 52690
rect 89450 52560 89550 52690
rect 89700 52560 89800 52690
rect 89950 52560 90050 52690
rect 90200 52560 90300 52690
rect 90450 52560 90550 52690
rect 90700 52560 90800 52690
rect 90950 52560 91050 52690
rect 91200 52560 91300 52690
rect 91450 52560 91550 52690
rect 91700 52560 91800 52690
rect 91950 52560 92050 52690
rect 92200 52560 92300 52690
rect 92450 52560 92550 52690
rect 92700 52560 92800 52690
rect 92950 52560 93050 52690
rect 93200 52560 93300 52690
rect 93450 52560 93550 52690
rect 93700 52560 93800 52690
rect 93950 52560 94050 52690
rect 94200 52560 94300 52690
rect 94450 52560 94550 52690
rect 94700 52560 94800 52690
rect 94950 52560 95050 52690
rect 95200 52560 95300 52690
rect 95450 52560 95550 52690
rect 95700 52560 95800 52690
rect 95950 52560 96050 52690
rect 96200 52560 96300 52690
rect 96450 52560 96550 52690
rect 96700 52560 96800 52690
rect 96950 52560 97050 52690
rect 97200 52560 97300 52690
rect 97450 52560 97550 52690
rect 97700 52560 97800 52690
rect 97950 52560 98050 52690
rect 98200 52560 98300 52690
rect 98450 52560 98550 52690
rect 98700 52560 98800 52690
rect 98950 52560 99050 52690
rect 99200 52560 99300 52690
rect 99450 52560 99550 52690
rect 99700 52560 99800 52690
rect 99950 52560 100050 52690
rect 100200 52560 100300 52690
rect 100450 52560 100550 52690
rect 100700 52560 100800 52690
rect 100950 52560 101050 52690
rect 101200 52560 101300 52690
rect 101450 52560 101550 52690
rect 101700 52560 101800 52690
rect 101950 52560 102050 52690
rect 102200 52560 102300 52690
rect 102450 52560 102550 52690
rect 102700 52560 102800 52690
rect 102950 52560 103050 52690
rect 103200 52560 103300 52690
rect 103450 52560 103550 52690
rect 103700 52560 103800 52690
rect 103950 52560 104050 52690
rect 104200 52560 104300 52690
rect 104450 52560 104550 52690
rect 104700 52560 104800 52690
rect 104950 52560 105050 52690
rect 105200 52560 105300 52690
rect 105450 52560 105550 52690
rect 105700 52560 105800 52690
rect 105950 52560 106050 52690
rect 106200 52560 106300 52690
rect 106450 52560 106550 52690
rect 106700 52560 106800 52690
rect 106950 52560 107050 52690
rect 107200 52560 107300 52690
rect 107450 52560 107550 52690
rect 107700 52560 107800 52690
rect 107950 52560 108050 52690
rect 108200 52560 108300 52690
rect 108450 52560 108550 52690
rect 108700 52560 108800 52690
rect 108950 52560 109050 52690
rect 109200 52560 109300 52690
rect 109450 52560 109550 52690
rect 109700 52560 109800 52690
rect 109950 52560 110050 52690
rect 110200 52560 110300 52690
rect 110450 52560 110550 52690
rect 110700 52560 110800 52690
rect 110950 52560 111050 52690
rect 111200 52560 111300 52690
rect 111450 52560 111550 52690
rect 111700 52560 111800 52690
rect 111950 52560 112050 52690
rect 112200 52560 112300 52690
rect 112450 52560 112550 52690
rect 112700 52560 112800 52690
rect 112950 52560 113050 52690
rect 113200 52560 113300 52690
rect 113450 52560 113550 52690
rect 113700 52560 113800 52690
rect 113950 52560 114050 52690
rect 114200 52560 114300 52690
rect 114450 52560 114550 52690
rect 114700 52560 114800 52690
rect 114950 52560 115050 52690
rect 115200 52560 115300 52690
rect 115450 52560 115550 52690
rect 115700 52560 115800 52690
rect 115950 52560 116000 52690
rect 89000 52550 89060 52560
rect 89190 52550 89310 52560
rect 89440 52550 89560 52560
rect 89690 52550 89810 52560
rect 89940 52550 90060 52560
rect 90190 52550 90310 52560
rect 90440 52550 90560 52560
rect 90690 52550 90810 52560
rect 90940 52550 91060 52560
rect 91190 52550 91310 52560
rect 91440 52550 91560 52560
rect 91690 52550 91810 52560
rect 91940 52550 92060 52560
rect 92190 52550 92310 52560
rect 92440 52550 92560 52560
rect 92690 52550 92810 52560
rect 92940 52550 93060 52560
rect 93190 52550 93310 52560
rect 93440 52550 93560 52560
rect 93690 52550 93810 52560
rect 93940 52550 94060 52560
rect 94190 52550 94310 52560
rect 94440 52550 94560 52560
rect 94690 52550 94810 52560
rect 94940 52550 95060 52560
rect 95190 52550 95310 52560
rect 95440 52550 95560 52560
rect 95690 52550 95810 52560
rect 95940 52550 96060 52560
rect 96190 52550 96310 52560
rect 96440 52550 96560 52560
rect 96690 52550 96810 52560
rect 96940 52550 97060 52560
rect 97190 52550 97310 52560
rect 97440 52550 97560 52560
rect 97690 52550 97810 52560
rect 97940 52550 98060 52560
rect 98190 52550 98310 52560
rect 98440 52550 98560 52560
rect 98690 52550 98810 52560
rect 98940 52550 99060 52560
rect 99190 52550 99310 52560
rect 99440 52550 99560 52560
rect 99690 52550 99810 52560
rect 99940 52550 100060 52560
rect 100190 52550 100310 52560
rect 100440 52550 100560 52560
rect 100690 52550 100810 52560
rect 100940 52550 101060 52560
rect 101190 52550 101310 52560
rect 101440 52550 101560 52560
rect 101690 52550 101810 52560
rect 101940 52550 102060 52560
rect 102190 52550 102310 52560
rect 102440 52550 102560 52560
rect 102690 52550 102810 52560
rect 102940 52550 103060 52560
rect 103190 52550 103310 52560
rect 103440 52550 103560 52560
rect 103690 52550 103810 52560
rect 103940 52550 104060 52560
rect 104190 52550 104310 52560
rect 104440 52550 104560 52560
rect 104690 52550 104810 52560
rect 104940 52550 105060 52560
rect 105190 52550 105310 52560
rect 105440 52550 105560 52560
rect 105690 52550 105810 52560
rect 105940 52550 106060 52560
rect 106190 52550 106310 52560
rect 106440 52550 106560 52560
rect 106690 52550 106810 52560
rect 106940 52550 107060 52560
rect 107190 52550 107310 52560
rect 107440 52550 107560 52560
rect 107690 52550 107810 52560
rect 107940 52550 108060 52560
rect 108190 52550 108310 52560
rect 108440 52550 108560 52560
rect 108690 52550 108810 52560
rect 108940 52550 109060 52560
rect 109190 52550 109310 52560
rect 109440 52550 109560 52560
rect 109690 52550 109810 52560
rect 109940 52550 110060 52560
rect 110190 52550 110310 52560
rect 110440 52550 110560 52560
rect 110690 52550 110810 52560
rect 110940 52550 111060 52560
rect 111190 52550 111310 52560
rect 111440 52550 111560 52560
rect 111690 52550 111810 52560
rect 111940 52550 112060 52560
rect 112190 52550 112310 52560
rect 112440 52550 112560 52560
rect 112690 52550 112810 52560
rect 112940 52550 113060 52560
rect 113190 52550 113310 52560
rect 113440 52550 113560 52560
rect 113690 52550 113810 52560
rect 113940 52550 114060 52560
rect 114190 52550 114310 52560
rect 114440 52550 114560 52560
rect 114690 52550 114810 52560
rect 114940 52550 115060 52560
rect 115190 52550 115310 52560
rect 115440 52550 115560 52560
rect 115690 52550 115810 52560
rect 115940 52550 116000 52560
rect 89000 52450 116000 52550
rect 89000 52440 89060 52450
rect 89190 52440 89310 52450
rect 89440 52440 89560 52450
rect 89690 52440 89810 52450
rect 89940 52440 90060 52450
rect 90190 52440 90310 52450
rect 90440 52440 90560 52450
rect 90690 52440 90810 52450
rect 90940 52440 91060 52450
rect 91190 52440 91310 52450
rect 91440 52440 91560 52450
rect 91690 52440 91810 52450
rect 91940 52440 92060 52450
rect 92190 52440 92310 52450
rect 92440 52440 92560 52450
rect 92690 52440 92810 52450
rect 92940 52440 93060 52450
rect 93190 52440 93310 52450
rect 93440 52440 93560 52450
rect 93690 52440 93810 52450
rect 93940 52440 94060 52450
rect 94190 52440 94310 52450
rect 94440 52440 94560 52450
rect 94690 52440 94810 52450
rect 94940 52440 95060 52450
rect 95190 52440 95310 52450
rect 95440 52440 95560 52450
rect 95690 52440 95810 52450
rect 95940 52440 96060 52450
rect 96190 52440 96310 52450
rect 96440 52440 96560 52450
rect 96690 52440 96810 52450
rect 96940 52440 97060 52450
rect 97190 52440 97310 52450
rect 97440 52440 97560 52450
rect 97690 52440 97810 52450
rect 97940 52440 98060 52450
rect 98190 52440 98310 52450
rect 98440 52440 98560 52450
rect 98690 52440 98810 52450
rect 98940 52440 99060 52450
rect 99190 52440 99310 52450
rect 99440 52440 99560 52450
rect 99690 52440 99810 52450
rect 99940 52440 100060 52450
rect 100190 52440 100310 52450
rect 100440 52440 100560 52450
rect 100690 52440 100810 52450
rect 100940 52440 101060 52450
rect 101190 52440 101310 52450
rect 101440 52440 101560 52450
rect 101690 52440 101810 52450
rect 101940 52440 102060 52450
rect 102190 52440 102310 52450
rect 102440 52440 102560 52450
rect 102690 52440 102810 52450
rect 102940 52440 103060 52450
rect 103190 52440 103310 52450
rect 103440 52440 103560 52450
rect 103690 52440 103810 52450
rect 103940 52440 104060 52450
rect 104190 52440 104310 52450
rect 104440 52440 104560 52450
rect 104690 52440 104810 52450
rect 104940 52440 105060 52450
rect 105190 52440 105310 52450
rect 105440 52440 105560 52450
rect 105690 52440 105810 52450
rect 105940 52440 106060 52450
rect 106190 52440 106310 52450
rect 106440 52440 106560 52450
rect 106690 52440 106810 52450
rect 106940 52440 107060 52450
rect 107190 52440 107310 52450
rect 107440 52440 107560 52450
rect 107690 52440 107810 52450
rect 107940 52440 108060 52450
rect 108190 52440 108310 52450
rect 108440 52440 108560 52450
rect 108690 52440 108810 52450
rect 108940 52440 109060 52450
rect 109190 52440 109310 52450
rect 109440 52440 109560 52450
rect 109690 52440 109810 52450
rect 109940 52440 110060 52450
rect 110190 52440 110310 52450
rect 110440 52440 110560 52450
rect 110690 52440 110810 52450
rect 110940 52440 111060 52450
rect 111190 52440 111310 52450
rect 111440 52440 111560 52450
rect 111690 52440 111810 52450
rect 111940 52440 112060 52450
rect 112190 52440 112310 52450
rect 112440 52440 112560 52450
rect 112690 52440 112810 52450
rect 112940 52440 113060 52450
rect 113190 52440 113310 52450
rect 113440 52440 113560 52450
rect 113690 52440 113810 52450
rect 113940 52440 114060 52450
rect 114190 52440 114310 52450
rect 114440 52440 114560 52450
rect 114690 52440 114810 52450
rect 114940 52440 115060 52450
rect 115190 52440 115310 52450
rect 115440 52440 115560 52450
rect 115690 52440 115810 52450
rect 115940 52440 116000 52450
rect 89000 52310 89050 52440
rect 89200 52310 89300 52440
rect 89450 52310 89550 52440
rect 89700 52310 89800 52440
rect 89950 52310 90050 52440
rect 90200 52310 90300 52440
rect 90450 52310 90550 52440
rect 90700 52310 90800 52440
rect 90950 52310 91050 52440
rect 91200 52310 91300 52440
rect 91450 52310 91550 52440
rect 91700 52310 91800 52440
rect 91950 52310 92050 52440
rect 92200 52310 92300 52440
rect 92450 52310 92550 52440
rect 92700 52310 92800 52440
rect 92950 52310 93050 52440
rect 93200 52310 93300 52440
rect 93450 52310 93550 52440
rect 93700 52310 93800 52440
rect 93950 52310 94050 52440
rect 94200 52310 94300 52440
rect 94450 52310 94550 52440
rect 94700 52310 94800 52440
rect 94950 52310 95050 52440
rect 95200 52310 95300 52440
rect 95450 52310 95550 52440
rect 95700 52310 95800 52440
rect 95950 52310 96050 52440
rect 96200 52310 96300 52440
rect 96450 52310 96550 52440
rect 96700 52310 96800 52440
rect 96950 52310 97050 52440
rect 97200 52310 97300 52440
rect 97450 52310 97550 52440
rect 97700 52310 97800 52440
rect 97950 52310 98050 52440
rect 98200 52310 98300 52440
rect 98450 52310 98550 52440
rect 98700 52310 98800 52440
rect 98950 52310 99050 52440
rect 99200 52310 99300 52440
rect 99450 52310 99550 52440
rect 99700 52310 99800 52440
rect 99950 52310 100050 52440
rect 100200 52310 100300 52440
rect 100450 52310 100550 52440
rect 100700 52310 100800 52440
rect 100950 52310 101050 52440
rect 101200 52310 101300 52440
rect 101450 52310 101550 52440
rect 101700 52310 101800 52440
rect 101950 52310 102050 52440
rect 102200 52310 102300 52440
rect 102450 52310 102550 52440
rect 102700 52310 102800 52440
rect 102950 52310 103050 52440
rect 103200 52310 103300 52440
rect 103450 52310 103550 52440
rect 103700 52310 103800 52440
rect 103950 52310 104050 52440
rect 104200 52310 104300 52440
rect 104450 52310 104550 52440
rect 104700 52310 104800 52440
rect 104950 52310 105050 52440
rect 105200 52310 105300 52440
rect 105450 52310 105550 52440
rect 105700 52310 105800 52440
rect 105950 52310 106050 52440
rect 106200 52310 106300 52440
rect 106450 52310 106550 52440
rect 106700 52310 106800 52440
rect 106950 52310 107050 52440
rect 107200 52310 107300 52440
rect 107450 52310 107550 52440
rect 107700 52310 107800 52440
rect 107950 52310 108050 52440
rect 108200 52310 108300 52440
rect 108450 52310 108550 52440
rect 108700 52310 108800 52440
rect 108950 52310 109050 52440
rect 109200 52310 109300 52440
rect 109450 52310 109550 52440
rect 109700 52310 109800 52440
rect 109950 52310 110050 52440
rect 110200 52310 110300 52440
rect 110450 52310 110550 52440
rect 110700 52310 110800 52440
rect 110950 52310 111050 52440
rect 111200 52310 111300 52440
rect 111450 52310 111550 52440
rect 111700 52310 111800 52440
rect 111950 52310 112050 52440
rect 112200 52310 112300 52440
rect 112450 52310 112550 52440
rect 112700 52310 112800 52440
rect 112950 52310 113050 52440
rect 113200 52310 113300 52440
rect 113450 52310 113550 52440
rect 113700 52310 113800 52440
rect 113950 52310 114050 52440
rect 114200 52310 114300 52440
rect 114450 52310 114550 52440
rect 114700 52310 114800 52440
rect 114950 52310 115050 52440
rect 115200 52310 115300 52440
rect 115450 52310 115550 52440
rect 115700 52310 115800 52440
rect 115950 52310 116000 52440
rect 89000 52300 89060 52310
rect 89190 52300 89310 52310
rect 89440 52300 89560 52310
rect 89690 52300 89810 52310
rect 89940 52300 90060 52310
rect 90190 52300 90310 52310
rect 90440 52300 90560 52310
rect 90690 52300 90810 52310
rect 90940 52300 91060 52310
rect 91190 52300 91310 52310
rect 91440 52300 91560 52310
rect 91690 52300 91810 52310
rect 91940 52300 92060 52310
rect 92190 52300 92310 52310
rect 92440 52300 92560 52310
rect 92690 52300 92810 52310
rect 92940 52300 93060 52310
rect 93190 52300 93310 52310
rect 93440 52300 93560 52310
rect 93690 52300 93810 52310
rect 93940 52300 94060 52310
rect 94190 52300 94310 52310
rect 94440 52300 94560 52310
rect 94690 52300 94810 52310
rect 94940 52300 95060 52310
rect 95190 52300 95310 52310
rect 95440 52300 95560 52310
rect 95690 52300 95810 52310
rect 95940 52300 96060 52310
rect 96190 52300 96310 52310
rect 96440 52300 96560 52310
rect 96690 52300 96810 52310
rect 96940 52300 97060 52310
rect 97190 52300 97310 52310
rect 97440 52300 97560 52310
rect 97690 52300 97810 52310
rect 97940 52300 98060 52310
rect 98190 52300 98310 52310
rect 98440 52300 98560 52310
rect 98690 52300 98810 52310
rect 98940 52300 99060 52310
rect 99190 52300 99310 52310
rect 99440 52300 99560 52310
rect 99690 52300 99810 52310
rect 99940 52300 100060 52310
rect 100190 52300 100310 52310
rect 100440 52300 100560 52310
rect 100690 52300 100810 52310
rect 100940 52300 101060 52310
rect 101190 52300 101310 52310
rect 101440 52300 101560 52310
rect 101690 52300 101810 52310
rect 101940 52300 102060 52310
rect 102190 52300 102310 52310
rect 102440 52300 102560 52310
rect 102690 52300 102810 52310
rect 102940 52300 103060 52310
rect 103190 52300 103310 52310
rect 103440 52300 103560 52310
rect 103690 52300 103810 52310
rect 103940 52300 104060 52310
rect 104190 52300 104310 52310
rect 104440 52300 104560 52310
rect 104690 52300 104810 52310
rect 104940 52300 105060 52310
rect 105190 52300 105310 52310
rect 105440 52300 105560 52310
rect 105690 52300 105810 52310
rect 105940 52300 106060 52310
rect 106190 52300 106310 52310
rect 106440 52300 106560 52310
rect 106690 52300 106810 52310
rect 106940 52300 107060 52310
rect 107190 52300 107310 52310
rect 107440 52300 107560 52310
rect 107690 52300 107810 52310
rect 107940 52300 108060 52310
rect 108190 52300 108310 52310
rect 108440 52300 108560 52310
rect 108690 52300 108810 52310
rect 108940 52300 109060 52310
rect 109190 52300 109310 52310
rect 109440 52300 109560 52310
rect 109690 52300 109810 52310
rect 109940 52300 110060 52310
rect 110190 52300 110310 52310
rect 110440 52300 110560 52310
rect 110690 52300 110810 52310
rect 110940 52300 111060 52310
rect 111190 52300 111310 52310
rect 111440 52300 111560 52310
rect 111690 52300 111810 52310
rect 111940 52300 112060 52310
rect 112190 52300 112310 52310
rect 112440 52300 112560 52310
rect 112690 52300 112810 52310
rect 112940 52300 113060 52310
rect 113190 52300 113310 52310
rect 113440 52300 113560 52310
rect 113690 52300 113810 52310
rect 113940 52300 114060 52310
rect 114190 52300 114310 52310
rect 114440 52300 114560 52310
rect 114690 52300 114810 52310
rect 114940 52300 115060 52310
rect 115190 52300 115310 52310
rect 115440 52300 115560 52310
rect 115690 52300 115810 52310
rect 115940 52300 116000 52310
rect 89000 52200 116000 52300
rect 89000 52190 89060 52200
rect 89190 52190 89310 52200
rect 89440 52190 89560 52200
rect 89690 52190 89810 52200
rect 89940 52190 90060 52200
rect 90190 52190 90310 52200
rect 90440 52190 90560 52200
rect 90690 52190 90810 52200
rect 90940 52190 91060 52200
rect 91190 52190 91310 52200
rect 91440 52190 91560 52200
rect 91690 52190 91810 52200
rect 91940 52190 92060 52200
rect 92190 52190 92310 52200
rect 92440 52190 92560 52200
rect 92690 52190 92810 52200
rect 92940 52190 93060 52200
rect 93190 52190 93310 52200
rect 93440 52190 93560 52200
rect 93690 52190 93810 52200
rect 93940 52190 94060 52200
rect 94190 52190 94310 52200
rect 94440 52190 94560 52200
rect 94690 52190 94810 52200
rect 94940 52190 95060 52200
rect 95190 52190 95310 52200
rect 95440 52190 95560 52200
rect 95690 52190 95810 52200
rect 95940 52190 96060 52200
rect 96190 52190 96310 52200
rect 96440 52190 96560 52200
rect 96690 52190 96810 52200
rect 96940 52190 97060 52200
rect 97190 52190 97310 52200
rect 97440 52190 97560 52200
rect 97690 52190 97810 52200
rect 97940 52190 98060 52200
rect 98190 52190 98310 52200
rect 98440 52190 98560 52200
rect 98690 52190 98810 52200
rect 98940 52190 99060 52200
rect 99190 52190 99310 52200
rect 99440 52190 99560 52200
rect 99690 52190 99810 52200
rect 99940 52190 100060 52200
rect 100190 52190 100310 52200
rect 100440 52190 100560 52200
rect 100690 52190 100810 52200
rect 100940 52190 101060 52200
rect 101190 52190 101310 52200
rect 101440 52190 101560 52200
rect 101690 52190 101810 52200
rect 101940 52190 102060 52200
rect 102190 52190 102310 52200
rect 102440 52190 102560 52200
rect 102690 52190 102810 52200
rect 102940 52190 103060 52200
rect 103190 52190 103310 52200
rect 103440 52190 103560 52200
rect 103690 52190 103810 52200
rect 103940 52190 104060 52200
rect 104190 52190 104310 52200
rect 104440 52190 104560 52200
rect 104690 52190 104810 52200
rect 104940 52190 105060 52200
rect 105190 52190 105310 52200
rect 105440 52190 105560 52200
rect 105690 52190 105810 52200
rect 105940 52190 106060 52200
rect 106190 52190 106310 52200
rect 106440 52190 106560 52200
rect 106690 52190 106810 52200
rect 106940 52190 107060 52200
rect 107190 52190 107310 52200
rect 107440 52190 107560 52200
rect 107690 52190 107810 52200
rect 107940 52190 108060 52200
rect 108190 52190 108310 52200
rect 108440 52190 108560 52200
rect 108690 52190 108810 52200
rect 108940 52190 109060 52200
rect 109190 52190 109310 52200
rect 109440 52190 109560 52200
rect 109690 52190 109810 52200
rect 109940 52190 110060 52200
rect 110190 52190 110310 52200
rect 110440 52190 110560 52200
rect 110690 52190 110810 52200
rect 110940 52190 111060 52200
rect 111190 52190 111310 52200
rect 111440 52190 111560 52200
rect 111690 52190 111810 52200
rect 111940 52190 112060 52200
rect 112190 52190 112310 52200
rect 112440 52190 112560 52200
rect 112690 52190 112810 52200
rect 112940 52190 113060 52200
rect 113190 52190 113310 52200
rect 113440 52190 113560 52200
rect 113690 52190 113810 52200
rect 113940 52190 114060 52200
rect 114190 52190 114310 52200
rect 114440 52190 114560 52200
rect 114690 52190 114810 52200
rect 114940 52190 115060 52200
rect 115190 52190 115310 52200
rect 115440 52190 115560 52200
rect 115690 52190 115810 52200
rect 115940 52190 116000 52200
rect 89000 52060 89050 52190
rect 89200 52060 89300 52190
rect 89450 52060 89550 52190
rect 89700 52060 89800 52190
rect 89950 52060 90050 52190
rect 90200 52060 90300 52190
rect 90450 52060 90550 52190
rect 90700 52060 90800 52190
rect 90950 52060 91050 52190
rect 91200 52060 91300 52190
rect 91450 52060 91550 52190
rect 91700 52060 91800 52190
rect 91950 52060 92050 52190
rect 92200 52060 92300 52190
rect 92450 52060 92550 52190
rect 92700 52060 92800 52190
rect 92950 52060 93050 52190
rect 93200 52060 93300 52190
rect 93450 52060 93550 52190
rect 93700 52060 93800 52190
rect 93950 52060 94050 52190
rect 94200 52060 94300 52190
rect 94450 52060 94550 52190
rect 94700 52060 94800 52190
rect 94950 52060 95050 52190
rect 95200 52060 95300 52190
rect 95450 52060 95550 52190
rect 95700 52060 95800 52190
rect 95950 52060 96050 52190
rect 96200 52060 96300 52190
rect 96450 52060 96550 52190
rect 96700 52060 96800 52190
rect 96950 52060 97050 52190
rect 97200 52060 97300 52190
rect 97450 52060 97550 52190
rect 97700 52060 97800 52190
rect 97950 52060 98050 52190
rect 98200 52060 98300 52190
rect 98450 52060 98550 52190
rect 98700 52060 98800 52190
rect 98950 52060 99050 52190
rect 99200 52060 99300 52190
rect 99450 52060 99550 52190
rect 99700 52060 99800 52190
rect 99950 52060 100050 52190
rect 100200 52060 100300 52190
rect 100450 52060 100550 52190
rect 100700 52060 100800 52190
rect 100950 52060 101050 52190
rect 101200 52060 101300 52190
rect 101450 52060 101550 52190
rect 101700 52060 101800 52190
rect 101950 52060 102050 52190
rect 102200 52060 102300 52190
rect 102450 52060 102550 52190
rect 102700 52060 102800 52190
rect 102950 52060 103050 52190
rect 103200 52060 103300 52190
rect 103450 52060 103550 52190
rect 103700 52060 103800 52190
rect 103950 52060 104050 52190
rect 104200 52060 104300 52190
rect 104450 52060 104550 52190
rect 104700 52060 104800 52190
rect 104950 52060 105050 52190
rect 105200 52060 105300 52190
rect 105450 52060 105550 52190
rect 105700 52060 105800 52190
rect 105950 52060 106050 52190
rect 106200 52060 106300 52190
rect 106450 52060 106550 52190
rect 106700 52060 106800 52190
rect 106950 52060 107050 52190
rect 107200 52060 107300 52190
rect 107450 52060 107550 52190
rect 107700 52060 107800 52190
rect 107950 52060 108050 52190
rect 108200 52060 108300 52190
rect 108450 52060 108550 52190
rect 108700 52060 108800 52190
rect 108950 52060 109050 52190
rect 109200 52060 109300 52190
rect 109450 52060 109550 52190
rect 109700 52060 109800 52190
rect 109950 52060 110050 52190
rect 110200 52060 110300 52190
rect 110450 52060 110550 52190
rect 110700 52060 110800 52190
rect 110950 52060 111050 52190
rect 111200 52060 111300 52190
rect 111450 52060 111550 52190
rect 111700 52060 111800 52190
rect 111950 52060 112050 52190
rect 112200 52060 112300 52190
rect 112450 52060 112550 52190
rect 112700 52060 112800 52190
rect 112950 52060 113050 52190
rect 113200 52060 113300 52190
rect 113450 52060 113550 52190
rect 113700 52060 113800 52190
rect 113950 52060 114050 52190
rect 114200 52060 114300 52190
rect 114450 52060 114550 52190
rect 114700 52060 114800 52190
rect 114950 52060 115050 52190
rect 115200 52060 115300 52190
rect 115450 52060 115550 52190
rect 115700 52060 115800 52190
rect 115950 52060 116000 52190
rect 89000 52050 89060 52060
rect 89190 52050 89310 52060
rect 89440 52050 89560 52060
rect 89690 52050 89810 52060
rect 89940 52050 90060 52060
rect 90190 52050 90310 52060
rect 90440 52050 90560 52060
rect 90690 52050 90810 52060
rect 90940 52050 91060 52060
rect 91190 52050 91310 52060
rect 91440 52050 91560 52060
rect 91690 52050 91810 52060
rect 91940 52050 92060 52060
rect 92190 52050 92310 52060
rect 92440 52050 92560 52060
rect 92690 52050 92810 52060
rect 92940 52050 93060 52060
rect 93190 52050 93310 52060
rect 93440 52050 93560 52060
rect 93690 52050 93810 52060
rect 93940 52050 94060 52060
rect 94190 52050 94310 52060
rect 94440 52050 94560 52060
rect 94690 52050 94810 52060
rect 94940 52050 95060 52060
rect 95190 52050 95310 52060
rect 95440 52050 95560 52060
rect 95690 52050 95810 52060
rect 95940 52050 96060 52060
rect 96190 52050 96310 52060
rect 96440 52050 96560 52060
rect 96690 52050 96810 52060
rect 96940 52050 97060 52060
rect 97190 52050 97310 52060
rect 97440 52050 97560 52060
rect 97690 52050 97810 52060
rect 97940 52050 98060 52060
rect 98190 52050 98310 52060
rect 98440 52050 98560 52060
rect 98690 52050 98810 52060
rect 98940 52050 99060 52060
rect 99190 52050 99310 52060
rect 99440 52050 99560 52060
rect 99690 52050 99810 52060
rect 99940 52050 100060 52060
rect 100190 52050 100310 52060
rect 100440 52050 100560 52060
rect 100690 52050 100810 52060
rect 100940 52050 101060 52060
rect 101190 52050 101310 52060
rect 101440 52050 101560 52060
rect 101690 52050 101810 52060
rect 101940 52050 102060 52060
rect 102190 52050 102310 52060
rect 102440 52050 102560 52060
rect 102690 52050 102810 52060
rect 102940 52050 103060 52060
rect 103190 52050 103310 52060
rect 103440 52050 103560 52060
rect 103690 52050 103810 52060
rect 103940 52050 104060 52060
rect 104190 52050 104310 52060
rect 104440 52050 104560 52060
rect 104690 52050 104810 52060
rect 104940 52050 105060 52060
rect 105190 52050 105310 52060
rect 105440 52050 105560 52060
rect 105690 52050 105810 52060
rect 105940 52050 106060 52060
rect 106190 52050 106310 52060
rect 106440 52050 106560 52060
rect 106690 52050 106810 52060
rect 106940 52050 107060 52060
rect 107190 52050 107310 52060
rect 107440 52050 107560 52060
rect 107690 52050 107810 52060
rect 107940 52050 108060 52060
rect 108190 52050 108310 52060
rect 108440 52050 108560 52060
rect 108690 52050 108810 52060
rect 108940 52050 109060 52060
rect 109190 52050 109310 52060
rect 109440 52050 109560 52060
rect 109690 52050 109810 52060
rect 109940 52050 110060 52060
rect 110190 52050 110310 52060
rect 110440 52050 110560 52060
rect 110690 52050 110810 52060
rect 110940 52050 111060 52060
rect 111190 52050 111310 52060
rect 111440 52050 111560 52060
rect 111690 52050 111810 52060
rect 111940 52050 112060 52060
rect 112190 52050 112310 52060
rect 112440 52050 112560 52060
rect 112690 52050 112810 52060
rect 112940 52050 113060 52060
rect 113190 52050 113310 52060
rect 113440 52050 113560 52060
rect 113690 52050 113810 52060
rect 113940 52050 114060 52060
rect 114190 52050 114310 52060
rect 114440 52050 114560 52060
rect 114690 52050 114810 52060
rect 114940 52050 115060 52060
rect 115190 52050 115310 52060
rect 115440 52050 115560 52060
rect 115690 52050 115810 52060
rect 115940 52050 116000 52060
rect 89000 51950 116000 52050
rect 89000 51940 89060 51950
rect 89190 51940 89310 51950
rect 89440 51940 89560 51950
rect 89690 51940 89810 51950
rect 89940 51940 90060 51950
rect 90190 51940 90310 51950
rect 90440 51940 90560 51950
rect 90690 51940 90810 51950
rect 90940 51940 91060 51950
rect 91190 51940 91310 51950
rect 91440 51940 91560 51950
rect 91690 51940 91810 51950
rect 91940 51940 92060 51950
rect 92190 51940 92310 51950
rect 92440 51940 92560 51950
rect 92690 51940 92810 51950
rect 92940 51940 93060 51950
rect 93190 51940 93310 51950
rect 93440 51940 93560 51950
rect 93690 51940 93810 51950
rect 93940 51940 94060 51950
rect 94190 51940 94310 51950
rect 94440 51940 94560 51950
rect 94690 51940 94810 51950
rect 94940 51940 95060 51950
rect 95190 51940 95310 51950
rect 95440 51940 95560 51950
rect 95690 51940 95810 51950
rect 95940 51940 96060 51950
rect 96190 51940 96310 51950
rect 96440 51940 96560 51950
rect 96690 51940 96810 51950
rect 96940 51940 97060 51950
rect 97190 51940 97310 51950
rect 97440 51940 97560 51950
rect 97690 51940 97810 51950
rect 97940 51940 98060 51950
rect 98190 51940 98310 51950
rect 98440 51940 98560 51950
rect 98690 51940 98810 51950
rect 98940 51940 99060 51950
rect 99190 51940 99310 51950
rect 99440 51940 99560 51950
rect 99690 51940 99810 51950
rect 99940 51940 100060 51950
rect 100190 51940 100310 51950
rect 100440 51940 100560 51950
rect 100690 51940 100810 51950
rect 100940 51940 101060 51950
rect 101190 51940 101310 51950
rect 101440 51940 101560 51950
rect 101690 51940 101810 51950
rect 101940 51940 102060 51950
rect 102190 51940 102310 51950
rect 102440 51940 102560 51950
rect 102690 51940 102810 51950
rect 102940 51940 103060 51950
rect 103190 51940 103310 51950
rect 103440 51940 103560 51950
rect 103690 51940 103810 51950
rect 103940 51940 104060 51950
rect 104190 51940 104310 51950
rect 104440 51940 104560 51950
rect 104690 51940 104810 51950
rect 104940 51940 105060 51950
rect 105190 51940 105310 51950
rect 105440 51940 105560 51950
rect 105690 51940 105810 51950
rect 105940 51940 106060 51950
rect 106190 51940 106310 51950
rect 106440 51940 106560 51950
rect 106690 51940 106810 51950
rect 106940 51940 107060 51950
rect 107190 51940 107310 51950
rect 107440 51940 107560 51950
rect 107690 51940 107810 51950
rect 107940 51940 108060 51950
rect 108190 51940 108310 51950
rect 108440 51940 108560 51950
rect 108690 51940 108810 51950
rect 108940 51940 109060 51950
rect 109190 51940 109310 51950
rect 109440 51940 109560 51950
rect 109690 51940 109810 51950
rect 109940 51940 110060 51950
rect 110190 51940 110310 51950
rect 110440 51940 110560 51950
rect 110690 51940 110810 51950
rect 110940 51940 111060 51950
rect 111190 51940 111310 51950
rect 111440 51940 111560 51950
rect 111690 51940 111810 51950
rect 111940 51940 112060 51950
rect 112190 51940 112310 51950
rect 112440 51940 112560 51950
rect 112690 51940 112810 51950
rect 112940 51940 113060 51950
rect 113190 51940 113310 51950
rect 113440 51940 113560 51950
rect 113690 51940 113810 51950
rect 113940 51940 114060 51950
rect 114190 51940 114310 51950
rect 114440 51940 114560 51950
rect 114690 51940 114810 51950
rect 114940 51940 115060 51950
rect 115190 51940 115310 51950
rect 115440 51940 115560 51950
rect 115690 51940 115810 51950
rect 115940 51940 116000 51950
rect 89000 51810 89050 51940
rect 89200 51810 89300 51940
rect 89450 51810 89550 51940
rect 89700 51810 89800 51940
rect 89950 51810 90050 51940
rect 90200 51810 90300 51940
rect 90450 51810 90550 51940
rect 90700 51810 90800 51940
rect 90950 51810 91050 51940
rect 91200 51810 91300 51940
rect 91450 51810 91550 51940
rect 91700 51810 91800 51940
rect 91950 51810 92050 51940
rect 92200 51810 92300 51940
rect 92450 51810 92550 51940
rect 92700 51810 92800 51940
rect 92950 51810 93050 51940
rect 93200 51810 93300 51940
rect 93450 51810 93550 51940
rect 93700 51810 93800 51940
rect 93950 51810 94050 51940
rect 94200 51810 94300 51940
rect 94450 51810 94550 51940
rect 94700 51810 94800 51940
rect 94950 51810 95050 51940
rect 95200 51810 95300 51940
rect 95450 51810 95550 51940
rect 95700 51810 95800 51940
rect 95950 51810 96050 51940
rect 96200 51810 96300 51940
rect 96450 51810 96550 51940
rect 96700 51810 96800 51940
rect 96950 51810 97050 51940
rect 97200 51810 97300 51940
rect 97450 51810 97550 51940
rect 97700 51810 97800 51940
rect 97950 51810 98050 51940
rect 98200 51810 98300 51940
rect 98450 51810 98550 51940
rect 98700 51810 98800 51940
rect 98950 51810 99050 51940
rect 99200 51810 99300 51940
rect 99450 51810 99550 51940
rect 99700 51810 99800 51940
rect 99950 51810 100050 51940
rect 100200 51810 100300 51940
rect 100450 51810 100550 51940
rect 100700 51810 100800 51940
rect 100950 51810 101050 51940
rect 101200 51810 101300 51940
rect 101450 51810 101550 51940
rect 101700 51810 101800 51940
rect 101950 51810 102050 51940
rect 102200 51810 102300 51940
rect 102450 51810 102550 51940
rect 102700 51810 102800 51940
rect 102950 51810 103050 51940
rect 103200 51810 103300 51940
rect 103450 51810 103550 51940
rect 103700 51810 103800 51940
rect 103950 51810 104050 51940
rect 104200 51810 104300 51940
rect 104450 51810 104550 51940
rect 104700 51810 104800 51940
rect 104950 51810 105050 51940
rect 105200 51810 105300 51940
rect 105450 51810 105550 51940
rect 105700 51810 105800 51940
rect 105950 51810 106050 51940
rect 106200 51810 106300 51940
rect 106450 51810 106550 51940
rect 106700 51810 106800 51940
rect 106950 51810 107050 51940
rect 107200 51810 107300 51940
rect 107450 51810 107550 51940
rect 107700 51810 107800 51940
rect 107950 51810 108050 51940
rect 108200 51810 108300 51940
rect 108450 51810 108550 51940
rect 108700 51810 108800 51940
rect 108950 51810 109050 51940
rect 109200 51810 109300 51940
rect 109450 51810 109550 51940
rect 109700 51810 109800 51940
rect 109950 51810 110050 51940
rect 110200 51810 110300 51940
rect 110450 51810 110550 51940
rect 110700 51810 110800 51940
rect 110950 51810 111050 51940
rect 111200 51810 111300 51940
rect 111450 51810 111550 51940
rect 111700 51810 111800 51940
rect 111950 51810 112050 51940
rect 112200 51810 112300 51940
rect 112450 51810 112550 51940
rect 112700 51810 112800 51940
rect 112950 51810 113050 51940
rect 113200 51810 113300 51940
rect 113450 51810 113550 51940
rect 113700 51810 113800 51940
rect 113950 51810 114050 51940
rect 114200 51810 114300 51940
rect 114450 51810 114550 51940
rect 114700 51810 114800 51940
rect 114950 51810 115050 51940
rect 115200 51810 115300 51940
rect 115450 51810 115550 51940
rect 115700 51810 115800 51940
rect 115950 51810 116000 51940
rect 89000 51800 89060 51810
rect 89190 51800 89310 51810
rect 89440 51800 89560 51810
rect 89690 51800 89810 51810
rect 89940 51800 90060 51810
rect 90190 51800 90310 51810
rect 90440 51800 90560 51810
rect 90690 51800 90810 51810
rect 90940 51800 91060 51810
rect 91190 51800 91310 51810
rect 91440 51800 91560 51810
rect 91690 51800 91810 51810
rect 91940 51800 92060 51810
rect 92190 51800 92310 51810
rect 92440 51800 92560 51810
rect 92690 51800 92810 51810
rect 92940 51800 93060 51810
rect 93190 51800 93310 51810
rect 93440 51800 93560 51810
rect 93690 51800 93810 51810
rect 93940 51800 94060 51810
rect 94190 51800 94310 51810
rect 94440 51800 94560 51810
rect 94690 51800 94810 51810
rect 94940 51800 95060 51810
rect 95190 51800 95310 51810
rect 95440 51800 95560 51810
rect 95690 51800 95810 51810
rect 95940 51800 96060 51810
rect 96190 51800 96310 51810
rect 96440 51800 96560 51810
rect 96690 51800 96810 51810
rect 96940 51800 97060 51810
rect 97190 51800 97310 51810
rect 97440 51800 97560 51810
rect 97690 51800 97810 51810
rect 97940 51800 98060 51810
rect 98190 51800 98310 51810
rect 98440 51800 98560 51810
rect 98690 51800 98810 51810
rect 98940 51800 99060 51810
rect 99190 51800 99310 51810
rect 99440 51800 99560 51810
rect 99690 51800 99810 51810
rect 99940 51800 100060 51810
rect 100190 51800 100310 51810
rect 100440 51800 100560 51810
rect 100690 51800 100810 51810
rect 100940 51800 101060 51810
rect 101190 51800 101310 51810
rect 101440 51800 101560 51810
rect 101690 51800 101810 51810
rect 101940 51800 102060 51810
rect 102190 51800 102310 51810
rect 102440 51800 102560 51810
rect 102690 51800 102810 51810
rect 102940 51800 103060 51810
rect 103190 51800 103310 51810
rect 103440 51800 103560 51810
rect 103690 51800 103810 51810
rect 103940 51800 104060 51810
rect 104190 51800 104310 51810
rect 104440 51800 104560 51810
rect 104690 51800 104810 51810
rect 104940 51800 105060 51810
rect 105190 51800 105310 51810
rect 105440 51800 105560 51810
rect 105690 51800 105810 51810
rect 105940 51800 106060 51810
rect 106190 51800 106310 51810
rect 106440 51800 106560 51810
rect 106690 51800 106810 51810
rect 106940 51800 107060 51810
rect 107190 51800 107310 51810
rect 107440 51800 107560 51810
rect 107690 51800 107810 51810
rect 107940 51800 108060 51810
rect 108190 51800 108310 51810
rect 108440 51800 108560 51810
rect 108690 51800 108810 51810
rect 108940 51800 109060 51810
rect 109190 51800 109310 51810
rect 109440 51800 109560 51810
rect 109690 51800 109810 51810
rect 109940 51800 110060 51810
rect 110190 51800 110310 51810
rect 110440 51800 110560 51810
rect 110690 51800 110810 51810
rect 110940 51800 111060 51810
rect 111190 51800 111310 51810
rect 111440 51800 111560 51810
rect 111690 51800 111810 51810
rect 111940 51800 112060 51810
rect 112190 51800 112310 51810
rect 112440 51800 112560 51810
rect 112690 51800 112810 51810
rect 112940 51800 113060 51810
rect 113190 51800 113310 51810
rect 113440 51800 113560 51810
rect 113690 51800 113810 51810
rect 113940 51800 114060 51810
rect 114190 51800 114310 51810
rect 114440 51800 114560 51810
rect 114690 51800 114810 51810
rect 114940 51800 115060 51810
rect 115190 51800 115310 51810
rect 115440 51800 115560 51810
rect 115690 51800 115810 51810
rect 115940 51800 116000 51810
rect 89000 51700 116000 51800
rect 89000 51690 89060 51700
rect 89190 51690 89310 51700
rect 89440 51690 89560 51700
rect 89690 51690 89810 51700
rect 89940 51690 90060 51700
rect 90190 51690 90310 51700
rect 90440 51690 90560 51700
rect 90690 51690 90810 51700
rect 90940 51690 91060 51700
rect 91190 51690 91310 51700
rect 91440 51690 91560 51700
rect 91690 51690 91810 51700
rect 91940 51690 92060 51700
rect 92190 51690 92310 51700
rect 92440 51690 92560 51700
rect 92690 51690 92810 51700
rect 92940 51690 93060 51700
rect 93190 51690 93310 51700
rect 93440 51690 93560 51700
rect 93690 51690 93810 51700
rect 93940 51690 94060 51700
rect 94190 51690 94310 51700
rect 94440 51690 94560 51700
rect 94690 51690 94810 51700
rect 94940 51690 95060 51700
rect 95190 51690 95310 51700
rect 95440 51690 95560 51700
rect 95690 51690 95810 51700
rect 95940 51690 96060 51700
rect 96190 51690 96310 51700
rect 96440 51690 96560 51700
rect 96690 51690 96810 51700
rect 96940 51690 97060 51700
rect 97190 51690 97310 51700
rect 97440 51690 97560 51700
rect 97690 51690 97810 51700
rect 97940 51690 98060 51700
rect 98190 51690 98310 51700
rect 98440 51690 98560 51700
rect 98690 51690 98810 51700
rect 98940 51690 99060 51700
rect 99190 51690 99310 51700
rect 99440 51690 99560 51700
rect 99690 51690 99810 51700
rect 99940 51690 100060 51700
rect 100190 51690 100310 51700
rect 100440 51690 100560 51700
rect 100690 51690 100810 51700
rect 100940 51690 101060 51700
rect 101190 51690 101310 51700
rect 101440 51690 101560 51700
rect 101690 51690 101810 51700
rect 101940 51690 102060 51700
rect 102190 51690 102310 51700
rect 102440 51690 102560 51700
rect 102690 51690 102810 51700
rect 102940 51690 103060 51700
rect 103190 51690 103310 51700
rect 103440 51690 103560 51700
rect 103690 51690 103810 51700
rect 103940 51690 104060 51700
rect 104190 51690 104310 51700
rect 104440 51690 104560 51700
rect 104690 51690 104810 51700
rect 104940 51690 105060 51700
rect 105190 51690 105310 51700
rect 105440 51690 105560 51700
rect 105690 51690 105810 51700
rect 105940 51690 106060 51700
rect 106190 51690 106310 51700
rect 106440 51690 106560 51700
rect 106690 51690 106810 51700
rect 106940 51690 107060 51700
rect 107190 51690 107310 51700
rect 107440 51690 107560 51700
rect 107690 51690 107810 51700
rect 107940 51690 108060 51700
rect 108190 51690 108310 51700
rect 108440 51690 108560 51700
rect 108690 51690 108810 51700
rect 108940 51690 109060 51700
rect 109190 51690 109310 51700
rect 109440 51690 109560 51700
rect 109690 51690 109810 51700
rect 109940 51690 110060 51700
rect 110190 51690 110310 51700
rect 110440 51690 110560 51700
rect 110690 51690 110810 51700
rect 110940 51690 111060 51700
rect 111190 51690 111310 51700
rect 111440 51690 111560 51700
rect 111690 51690 111810 51700
rect 111940 51690 112060 51700
rect 112190 51690 112310 51700
rect 112440 51690 112560 51700
rect 112690 51690 112810 51700
rect 112940 51690 113060 51700
rect 113190 51690 113310 51700
rect 113440 51690 113560 51700
rect 113690 51690 113810 51700
rect 113940 51690 114060 51700
rect 114190 51690 114310 51700
rect 114440 51690 114560 51700
rect 114690 51690 114810 51700
rect 114940 51690 115060 51700
rect 115190 51690 115310 51700
rect 115440 51690 115560 51700
rect 115690 51690 115810 51700
rect 115940 51690 116000 51700
rect 89000 51560 89050 51690
rect 89200 51560 89300 51690
rect 89450 51560 89550 51690
rect 89700 51560 89800 51690
rect 89950 51560 90050 51690
rect 90200 51560 90300 51690
rect 90450 51560 90550 51690
rect 90700 51560 90800 51690
rect 90950 51560 91050 51690
rect 91200 51560 91300 51690
rect 91450 51560 91550 51690
rect 91700 51560 91800 51690
rect 91950 51560 92050 51690
rect 92200 51560 92300 51690
rect 92450 51560 92550 51690
rect 92700 51560 92800 51690
rect 92950 51560 93050 51690
rect 93200 51560 93300 51690
rect 93450 51560 93550 51690
rect 93700 51560 93800 51690
rect 93950 51560 94050 51690
rect 94200 51560 94300 51690
rect 94450 51560 94550 51690
rect 94700 51560 94800 51690
rect 94950 51560 95050 51690
rect 95200 51560 95300 51690
rect 95450 51560 95550 51690
rect 95700 51560 95800 51690
rect 95950 51560 96050 51690
rect 96200 51560 96300 51690
rect 96450 51560 96550 51690
rect 96700 51560 96800 51690
rect 96950 51560 97050 51690
rect 97200 51560 97300 51690
rect 97450 51560 97550 51690
rect 97700 51560 97800 51690
rect 97950 51560 98050 51690
rect 98200 51560 98300 51690
rect 98450 51560 98550 51690
rect 98700 51560 98800 51690
rect 98950 51560 99050 51690
rect 99200 51560 99300 51690
rect 99450 51560 99550 51690
rect 99700 51560 99800 51690
rect 99950 51560 100050 51690
rect 100200 51560 100300 51690
rect 100450 51560 100550 51690
rect 100700 51560 100800 51690
rect 100950 51560 101050 51690
rect 101200 51560 101300 51690
rect 101450 51560 101550 51690
rect 101700 51560 101800 51690
rect 101950 51560 102050 51690
rect 102200 51560 102300 51690
rect 102450 51560 102550 51690
rect 102700 51560 102800 51690
rect 102950 51560 103050 51690
rect 103200 51560 103300 51690
rect 103450 51560 103550 51690
rect 103700 51560 103800 51690
rect 103950 51560 104050 51690
rect 104200 51560 104300 51690
rect 104450 51560 104550 51690
rect 104700 51560 104800 51690
rect 104950 51560 105050 51690
rect 105200 51560 105300 51690
rect 105450 51560 105550 51690
rect 105700 51560 105800 51690
rect 105950 51560 106050 51690
rect 106200 51560 106300 51690
rect 106450 51560 106550 51690
rect 106700 51560 106800 51690
rect 106950 51560 107050 51690
rect 107200 51560 107300 51690
rect 107450 51560 107550 51690
rect 107700 51560 107800 51690
rect 107950 51560 108050 51690
rect 108200 51560 108300 51690
rect 108450 51560 108550 51690
rect 108700 51560 108800 51690
rect 108950 51560 109050 51690
rect 109200 51560 109300 51690
rect 109450 51560 109550 51690
rect 109700 51560 109800 51690
rect 109950 51560 110050 51690
rect 110200 51560 110300 51690
rect 110450 51560 110550 51690
rect 110700 51560 110800 51690
rect 110950 51560 111050 51690
rect 111200 51560 111300 51690
rect 111450 51560 111550 51690
rect 111700 51560 111800 51690
rect 111950 51560 112050 51690
rect 112200 51560 112300 51690
rect 112450 51560 112550 51690
rect 112700 51560 112800 51690
rect 112950 51560 113050 51690
rect 113200 51560 113300 51690
rect 113450 51560 113550 51690
rect 113700 51560 113800 51690
rect 113950 51560 114050 51690
rect 114200 51560 114300 51690
rect 114450 51560 114550 51690
rect 114700 51560 114800 51690
rect 114950 51560 115050 51690
rect 115200 51560 115300 51690
rect 115450 51560 115550 51690
rect 115700 51560 115800 51690
rect 115950 51560 116000 51690
rect 89000 51550 89060 51560
rect 89190 51550 89310 51560
rect 89440 51550 89560 51560
rect 89690 51550 89810 51560
rect 89940 51550 90060 51560
rect 90190 51550 90310 51560
rect 90440 51550 90560 51560
rect 90690 51550 90810 51560
rect 90940 51550 91060 51560
rect 91190 51550 91310 51560
rect 91440 51550 91560 51560
rect 91690 51550 91810 51560
rect 91940 51550 92060 51560
rect 92190 51550 92310 51560
rect 92440 51550 92560 51560
rect 92690 51550 92810 51560
rect 92940 51550 93060 51560
rect 93190 51550 93310 51560
rect 93440 51550 93560 51560
rect 93690 51550 93810 51560
rect 93940 51550 94060 51560
rect 94190 51550 94310 51560
rect 94440 51550 94560 51560
rect 94690 51550 94810 51560
rect 94940 51550 95060 51560
rect 95190 51550 95310 51560
rect 95440 51550 95560 51560
rect 95690 51550 95810 51560
rect 95940 51550 96060 51560
rect 96190 51550 96310 51560
rect 96440 51550 96560 51560
rect 96690 51550 96810 51560
rect 96940 51550 97060 51560
rect 97190 51550 97310 51560
rect 97440 51550 97560 51560
rect 97690 51550 97810 51560
rect 97940 51550 98060 51560
rect 98190 51550 98310 51560
rect 98440 51550 98560 51560
rect 98690 51550 98810 51560
rect 98940 51550 99060 51560
rect 99190 51550 99310 51560
rect 99440 51550 99560 51560
rect 99690 51550 99810 51560
rect 99940 51550 100060 51560
rect 100190 51550 100310 51560
rect 100440 51550 100560 51560
rect 100690 51550 100810 51560
rect 100940 51550 101060 51560
rect 101190 51550 101310 51560
rect 101440 51550 101560 51560
rect 101690 51550 101810 51560
rect 101940 51550 102060 51560
rect 102190 51550 102310 51560
rect 102440 51550 102560 51560
rect 102690 51550 102810 51560
rect 102940 51550 103060 51560
rect 103190 51550 103310 51560
rect 103440 51550 103560 51560
rect 103690 51550 103810 51560
rect 103940 51550 104060 51560
rect 104190 51550 104310 51560
rect 104440 51550 104560 51560
rect 104690 51550 104810 51560
rect 104940 51550 105060 51560
rect 105190 51550 105310 51560
rect 105440 51550 105560 51560
rect 105690 51550 105810 51560
rect 105940 51550 106060 51560
rect 106190 51550 106310 51560
rect 106440 51550 106560 51560
rect 106690 51550 106810 51560
rect 106940 51550 107060 51560
rect 107190 51550 107310 51560
rect 107440 51550 107560 51560
rect 107690 51550 107810 51560
rect 107940 51550 108060 51560
rect 108190 51550 108310 51560
rect 108440 51550 108560 51560
rect 108690 51550 108810 51560
rect 108940 51550 109060 51560
rect 109190 51550 109310 51560
rect 109440 51550 109560 51560
rect 109690 51550 109810 51560
rect 109940 51550 110060 51560
rect 110190 51550 110310 51560
rect 110440 51550 110560 51560
rect 110690 51550 110810 51560
rect 110940 51550 111060 51560
rect 111190 51550 111310 51560
rect 111440 51550 111560 51560
rect 111690 51550 111810 51560
rect 111940 51550 112060 51560
rect 112190 51550 112310 51560
rect 112440 51550 112560 51560
rect 112690 51550 112810 51560
rect 112940 51550 113060 51560
rect 113190 51550 113310 51560
rect 113440 51550 113560 51560
rect 113690 51550 113810 51560
rect 113940 51550 114060 51560
rect 114190 51550 114310 51560
rect 114440 51550 114560 51560
rect 114690 51550 114810 51560
rect 114940 51550 115060 51560
rect 115190 51550 115310 51560
rect 115440 51550 115560 51560
rect 115690 51550 115810 51560
rect 115940 51550 116000 51560
rect 89000 51450 116000 51550
rect 89000 51440 89060 51450
rect 89190 51440 89310 51450
rect 89440 51440 89560 51450
rect 89690 51440 89810 51450
rect 89940 51440 90060 51450
rect 90190 51440 90310 51450
rect 90440 51440 90560 51450
rect 90690 51440 90810 51450
rect 90940 51440 91060 51450
rect 91190 51440 91310 51450
rect 91440 51440 91560 51450
rect 91690 51440 91810 51450
rect 91940 51440 92060 51450
rect 92190 51440 92310 51450
rect 92440 51440 92560 51450
rect 92690 51440 92810 51450
rect 92940 51440 93060 51450
rect 93190 51440 93310 51450
rect 93440 51440 93560 51450
rect 93690 51440 93810 51450
rect 93940 51440 94060 51450
rect 94190 51440 94310 51450
rect 94440 51440 94560 51450
rect 94690 51440 94810 51450
rect 94940 51440 95060 51450
rect 95190 51440 95310 51450
rect 95440 51440 95560 51450
rect 95690 51440 95810 51450
rect 95940 51440 96060 51450
rect 96190 51440 96310 51450
rect 96440 51440 96560 51450
rect 96690 51440 96810 51450
rect 96940 51440 97060 51450
rect 97190 51440 97310 51450
rect 97440 51440 97560 51450
rect 97690 51440 97810 51450
rect 97940 51440 98060 51450
rect 98190 51440 98310 51450
rect 98440 51440 98560 51450
rect 98690 51440 98810 51450
rect 98940 51440 99060 51450
rect 99190 51440 99310 51450
rect 99440 51440 99560 51450
rect 99690 51440 99810 51450
rect 99940 51440 100060 51450
rect 100190 51440 100310 51450
rect 100440 51440 100560 51450
rect 100690 51440 100810 51450
rect 100940 51440 101060 51450
rect 101190 51440 101310 51450
rect 101440 51440 101560 51450
rect 101690 51440 101810 51450
rect 101940 51440 102060 51450
rect 102190 51440 102310 51450
rect 102440 51440 102560 51450
rect 102690 51440 102810 51450
rect 102940 51440 103060 51450
rect 103190 51440 103310 51450
rect 103440 51440 103560 51450
rect 103690 51440 103810 51450
rect 103940 51440 104060 51450
rect 104190 51440 104310 51450
rect 104440 51440 104560 51450
rect 104690 51440 104810 51450
rect 104940 51440 105060 51450
rect 105190 51440 105310 51450
rect 105440 51440 105560 51450
rect 105690 51440 105810 51450
rect 105940 51440 106060 51450
rect 106190 51440 106310 51450
rect 106440 51440 106560 51450
rect 106690 51440 106810 51450
rect 106940 51440 107060 51450
rect 107190 51440 107310 51450
rect 107440 51440 107560 51450
rect 107690 51440 107810 51450
rect 107940 51440 108060 51450
rect 108190 51440 108310 51450
rect 108440 51440 108560 51450
rect 108690 51440 108810 51450
rect 108940 51440 109060 51450
rect 109190 51440 109310 51450
rect 109440 51440 109560 51450
rect 109690 51440 109810 51450
rect 109940 51440 110060 51450
rect 110190 51440 110310 51450
rect 110440 51440 110560 51450
rect 110690 51440 110810 51450
rect 110940 51440 111060 51450
rect 111190 51440 111310 51450
rect 111440 51440 111560 51450
rect 111690 51440 111810 51450
rect 111940 51440 112060 51450
rect 112190 51440 112310 51450
rect 112440 51440 112560 51450
rect 112690 51440 112810 51450
rect 112940 51440 113060 51450
rect 113190 51440 113310 51450
rect 113440 51440 113560 51450
rect 113690 51440 113810 51450
rect 113940 51440 114060 51450
rect 114190 51440 114310 51450
rect 114440 51440 114560 51450
rect 114690 51440 114810 51450
rect 114940 51440 115060 51450
rect 115190 51440 115310 51450
rect 115440 51440 115560 51450
rect 115690 51440 115810 51450
rect 115940 51440 116000 51450
rect 89000 51310 89050 51440
rect 89200 51310 89300 51440
rect 89450 51310 89550 51440
rect 89700 51310 89800 51440
rect 89950 51310 90050 51440
rect 90200 51310 90300 51440
rect 90450 51310 90550 51440
rect 90700 51310 90800 51440
rect 90950 51310 91050 51440
rect 91200 51310 91300 51440
rect 91450 51310 91550 51440
rect 91700 51310 91800 51440
rect 91950 51310 92050 51440
rect 92200 51310 92300 51440
rect 92450 51310 92550 51440
rect 92700 51310 92800 51440
rect 92950 51310 93050 51440
rect 93200 51310 93300 51440
rect 93450 51310 93550 51440
rect 93700 51310 93800 51440
rect 93950 51310 94050 51440
rect 94200 51310 94300 51440
rect 94450 51310 94550 51440
rect 94700 51310 94800 51440
rect 94950 51310 95050 51440
rect 95200 51310 95300 51440
rect 95450 51310 95550 51440
rect 95700 51310 95800 51440
rect 95950 51310 96050 51440
rect 96200 51310 96300 51440
rect 96450 51310 96550 51440
rect 96700 51310 96800 51440
rect 96950 51310 97050 51440
rect 97200 51310 97300 51440
rect 97450 51310 97550 51440
rect 97700 51310 97800 51440
rect 97950 51310 98050 51440
rect 98200 51310 98300 51440
rect 98450 51310 98550 51440
rect 98700 51310 98800 51440
rect 98950 51310 99050 51440
rect 99200 51310 99300 51440
rect 99450 51310 99550 51440
rect 99700 51310 99800 51440
rect 99950 51310 100050 51440
rect 100200 51310 100300 51440
rect 100450 51310 100550 51440
rect 100700 51310 100800 51440
rect 100950 51310 101050 51440
rect 101200 51310 101300 51440
rect 101450 51310 101550 51440
rect 101700 51310 101800 51440
rect 101950 51310 102050 51440
rect 102200 51310 102300 51440
rect 102450 51310 102550 51440
rect 102700 51310 102800 51440
rect 102950 51310 103050 51440
rect 103200 51310 103300 51440
rect 103450 51310 103550 51440
rect 103700 51310 103800 51440
rect 103950 51310 104050 51440
rect 104200 51310 104300 51440
rect 104450 51310 104550 51440
rect 104700 51310 104800 51440
rect 104950 51310 105050 51440
rect 105200 51310 105300 51440
rect 105450 51310 105550 51440
rect 105700 51310 105800 51440
rect 105950 51310 106050 51440
rect 106200 51310 106300 51440
rect 106450 51310 106550 51440
rect 106700 51310 106800 51440
rect 106950 51310 107050 51440
rect 107200 51310 107300 51440
rect 107450 51310 107550 51440
rect 107700 51310 107800 51440
rect 107950 51310 108050 51440
rect 108200 51310 108300 51440
rect 108450 51310 108550 51440
rect 108700 51310 108800 51440
rect 108950 51310 109050 51440
rect 109200 51310 109300 51440
rect 109450 51310 109550 51440
rect 109700 51310 109800 51440
rect 109950 51310 110050 51440
rect 110200 51310 110300 51440
rect 110450 51310 110550 51440
rect 110700 51310 110800 51440
rect 110950 51310 111050 51440
rect 111200 51310 111300 51440
rect 111450 51310 111550 51440
rect 111700 51310 111800 51440
rect 111950 51310 112050 51440
rect 112200 51310 112300 51440
rect 112450 51310 112550 51440
rect 112700 51310 112800 51440
rect 112950 51310 113050 51440
rect 113200 51310 113300 51440
rect 113450 51310 113550 51440
rect 113700 51310 113800 51440
rect 113950 51310 114050 51440
rect 114200 51310 114300 51440
rect 114450 51310 114550 51440
rect 114700 51310 114800 51440
rect 114950 51310 115050 51440
rect 115200 51310 115300 51440
rect 115450 51310 115550 51440
rect 115700 51310 115800 51440
rect 115950 51310 116000 51440
rect 89000 51300 89060 51310
rect 89190 51300 89310 51310
rect 89440 51300 89560 51310
rect 89690 51300 89810 51310
rect 89940 51300 90060 51310
rect 90190 51300 90310 51310
rect 90440 51300 90560 51310
rect 90690 51300 90810 51310
rect 90940 51300 91060 51310
rect 91190 51300 91310 51310
rect 91440 51300 91560 51310
rect 91690 51300 91810 51310
rect 91940 51300 92060 51310
rect 92190 51300 92310 51310
rect 92440 51300 92560 51310
rect 92690 51300 92810 51310
rect 92940 51300 93060 51310
rect 93190 51300 93310 51310
rect 93440 51300 93560 51310
rect 93690 51300 93810 51310
rect 93940 51300 94060 51310
rect 94190 51300 94310 51310
rect 94440 51300 94560 51310
rect 94690 51300 94810 51310
rect 94940 51300 95060 51310
rect 95190 51300 95310 51310
rect 95440 51300 95560 51310
rect 95690 51300 95810 51310
rect 95940 51300 96060 51310
rect 96190 51300 96310 51310
rect 96440 51300 96560 51310
rect 96690 51300 96810 51310
rect 96940 51300 97060 51310
rect 97190 51300 97310 51310
rect 97440 51300 97560 51310
rect 97690 51300 97810 51310
rect 97940 51300 98060 51310
rect 98190 51300 98310 51310
rect 98440 51300 98560 51310
rect 98690 51300 98810 51310
rect 98940 51300 99060 51310
rect 99190 51300 99310 51310
rect 99440 51300 99560 51310
rect 99690 51300 99810 51310
rect 99940 51300 100060 51310
rect 100190 51300 100310 51310
rect 100440 51300 100560 51310
rect 100690 51300 100810 51310
rect 100940 51300 101060 51310
rect 101190 51300 101310 51310
rect 101440 51300 101560 51310
rect 101690 51300 101810 51310
rect 101940 51300 102060 51310
rect 102190 51300 102310 51310
rect 102440 51300 102560 51310
rect 102690 51300 102810 51310
rect 102940 51300 103060 51310
rect 103190 51300 103310 51310
rect 103440 51300 103560 51310
rect 103690 51300 103810 51310
rect 103940 51300 104060 51310
rect 104190 51300 104310 51310
rect 104440 51300 104560 51310
rect 104690 51300 104810 51310
rect 104940 51300 105060 51310
rect 105190 51300 105310 51310
rect 105440 51300 105560 51310
rect 105690 51300 105810 51310
rect 105940 51300 106060 51310
rect 106190 51300 106310 51310
rect 106440 51300 106560 51310
rect 106690 51300 106810 51310
rect 106940 51300 107060 51310
rect 107190 51300 107310 51310
rect 107440 51300 107560 51310
rect 107690 51300 107810 51310
rect 107940 51300 108060 51310
rect 108190 51300 108310 51310
rect 108440 51300 108560 51310
rect 108690 51300 108810 51310
rect 108940 51300 109060 51310
rect 109190 51300 109310 51310
rect 109440 51300 109560 51310
rect 109690 51300 109810 51310
rect 109940 51300 110060 51310
rect 110190 51300 110310 51310
rect 110440 51300 110560 51310
rect 110690 51300 110810 51310
rect 110940 51300 111060 51310
rect 111190 51300 111310 51310
rect 111440 51300 111560 51310
rect 111690 51300 111810 51310
rect 111940 51300 112060 51310
rect 112190 51300 112310 51310
rect 112440 51300 112560 51310
rect 112690 51300 112810 51310
rect 112940 51300 113060 51310
rect 113190 51300 113310 51310
rect 113440 51300 113560 51310
rect 113690 51300 113810 51310
rect 113940 51300 114060 51310
rect 114190 51300 114310 51310
rect 114440 51300 114560 51310
rect 114690 51300 114810 51310
rect 114940 51300 115060 51310
rect 115190 51300 115310 51310
rect 115440 51300 115560 51310
rect 115690 51300 115810 51310
rect 115940 51300 116000 51310
rect 89000 51200 116000 51300
rect 89000 51190 89060 51200
rect 89190 51190 89310 51200
rect 89440 51190 89560 51200
rect 89690 51190 89810 51200
rect 89940 51190 90060 51200
rect 90190 51190 90310 51200
rect 90440 51190 90560 51200
rect 90690 51190 90810 51200
rect 90940 51190 91060 51200
rect 91190 51190 91310 51200
rect 91440 51190 91560 51200
rect 91690 51190 91810 51200
rect 91940 51190 92060 51200
rect 92190 51190 92310 51200
rect 92440 51190 92560 51200
rect 92690 51190 92810 51200
rect 92940 51190 93060 51200
rect 93190 51190 93310 51200
rect 93440 51190 93560 51200
rect 93690 51190 93810 51200
rect 93940 51190 94060 51200
rect 94190 51190 94310 51200
rect 94440 51190 94560 51200
rect 94690 51190 94810 51200
rect 94940 51190 95060 51200
rect 95190 51190 95310 51200
rect 95440 51190 95560 51200
rect 95690 51190 95810 51200
rect 95940 51190 96060 51200
rect 96190 51190 96310 51200
rect 96440 51190 96560 51200
rect 96690 51190 96810 51200
rect 96940 51190 97060 51200
rect 97190 51190 97310 51200
rect 97440 51190 97560 51200
rect 97690 51190 97810 51200
rect 97940 51190 98060 51200
rect 98190 51190 98310 51200
rect 98440 51190 98560 51200
rect 98690 51190 98810 51200
rect 98940 51190 99060 51200
rect 99190 51190 99310 51200
rect 99440 51190 99560 51200
rect 99690 51190 99810 51200
rect 99940 51190 100060 51200
rect 100190 51190 100310 51200
rect 100440 51190 100560 51200
rect 100690 51190 100810 51200
rect 100940 51190 101060 51200
rect 101190 51190 101310 51200
rect 101440 51190 101560 51200
rect 101690 51190 101810 51200
rect 101940 51190 102060 51200
rect 102190 51190 102310 51200
rect 102440 51190 102560 51200
rect 102690 51190 102810 51200
rect 102940 51190 103060 51200
rect 103190 51190 103310 51200
rect 103440 51190 103560 51200
rect 103690 51190 103810 51200
rect 103940 51190 104060 51200
rect 104190 51190 104310 51200
rect 104440 51190 104560 51200
rect 104690 51190 104810 51200
rect 104940 51190 105060 51200
rect 105190 51190 105310 51200
rect 105440 51190 105560 51200
rect 105690 51190 105810 51200
rect 105940 51190 106060 51200
rect 106190 51190 106310 51200
rect 106440 51190 106560 51200
rect 106690 51190 106810 51200
rect 106940 51190 107060 51200
rect 107190 51190 107310 51200
rect 107440 51190 107560 51200
rect 107690 51190 107810 51200
rect 107940 51190 108060 51200
rect 108190 51190 108310 51200
rect 108440 51190 108560 51200
rect 108690 51190 108810 51200
rect 108940 51190 109060 51200
rect 109190 51190 109310 51200
rect 109440 51190 109560 51200
rect 109690 51190 109810 51200
rect 109940 51190 110060 51200
rect 110190 51190 110310 51200
rect 110440 51190 110560 51200
rect 110690 51190 110810 51200
rect 110940 51190 111060 51200
rect 111190 51190 111310 51200
rect 111440 51190 111560 51200
rect 111690 51190 111810 51200
rect 111940 51190 112060 51200
rect 112190 51190 112310 51200
rect 112440 51190 112560 51200
rect 112690 51190 112810 51200
rect 112940 51190 113060 51200
rect 113190 51190 113310 51200
rect 113440 51190 113560 51200
rect 113690 51190 113810 51200
rect 113940 51190 114060 51200
rect 114190 51190 114310 51200
rect 114440 51190 114560 51200
rect 114690 51190 114810 51200
rect 114940 51190 115060 51200
rect 115190 51190 115310 51200
rect 115440 51190 115560 51200
rect 115690 51190 115810 51200
rect 115940 51190 116000 51200
rect 89000 51060 89050 51190
rect 89200 51060 89300 51190
rect 89450 51060 89550 51190
rect 89700 51060 89800 51190
rect 89950 51060 90050 51190
rect 90200 51060 90300 51190
rect 90450 51060 90550 51190
rect 90700 51060 90800 51190
rect 90950 51060 91050 51190
rect 91200 51060 91300 51190
rect 91450 51060 91550 51190
rect 91700 51060 91800 51190
rect 91950 51060 92050 51190
rect 92200 51060 92300 51190
rect 92450 51060 92550 51190
rect 92700 51060 92800 51190
rect 92950 51060 93050 51190
rect 93200 51060 93300 51190
rect 93450 51060 93550 51190
rect 93700 51060 93800 51190
rect 93950 51060 94050 51190
rect 94200 51060 94300 51190
rect 94450 51060 94550 51190
rect 94700 51060 94800 51190
rect 94950 51060 95050 51190
rect 95200 51060 95300 51190
rect 95450 51060 95550 51190
rect 95700 51060 95800 51190
rect 95950 51060 96050 51190
rect 96200 51060 96300 51190
rect 96450 51060 96550 51190
rect 96700 51060 96800 51190
rect 96950 51060 97050 51190
rect 97200 51060 97300 51190
rect 97450 51060 97550 51190
rect 97700 51060 97800 51190
rect 97950 51060 98050 51190
rect 98200 51060 98300 51190
rect 98450 51060 98550 51190
rect 98700 51060 98800 51190
rect 98950 51060 99050 51190
rect 99200 51060 99300 51190
rect 99450 51060 99550 51190
rect 99700 51060 99800 51190
rect 99950 51060 100050 51190
rect 100200 51060 100300 51190
rect 100450 51060 100550 51190
rect 100700 51060 100800 51190
rect 100950 51060 101050 51190
rect 101200 51060 101300 51190
rect 101450 51060 101550 51190
rect 101700 51060 101800 51190
rect 101950 51060 102050 51190
rect 102200 51060 102300 51190
rect 102450 51060 102550 51190
rect 102700 51060 102800 51190
rect 102950 51060 103050 51190
rect 103200 51060 103300 51190
rect 103450 51060 103550 51190
rect 103700 51060 103800 51190
rect 103950 51060 104050 51190
rect 104200 51060 104300 51190
rect 104450 51060 104550 51190
rect 104700 51060 104800 51190
rect 104950 51060 105050 51190
rect 105200 51060 105300 51190
rect 105450 51060 105550 51190
rect 105700 51060 105800 51190
rect 105950 51060 106050 51190
rect 106200 51060 106300 51190
rect 106450 51060 106550 51190
rect 106700 51060 106800 51190
rect 106950 51060 107050 51190
rect 107200 51060 107300 51190
rect 107450 51060 107550 51190
rect 107700 51060 107800 51190
rect 107950 51060 108050 51190
rect 108200 51060 108300 51190
rect 108450 51060 108550 51190
rect 108700 51060 108800 51190
rect 108950 51060 109050 51190
rect 109200 51060 109300 51190
rect 109450 51060 109550 51190
rect 109700 51060 109800 51190
rect 109950 51060 110050 51190
rect 110200 51060 110300 51190
rect 110450 51060 110550 51190
rect 110700 51060 110800 51190
rect 110950 51060 111050 51190
rect 111200 51060 111300 51190
rect 111450 51060 111550 51190
rect 111700 51060 111800 51190
rect 111950 51060 112050 51190
rect 112200 51060 112300 51190
rect 112450 51060 112550 51190
rect 112700 51060 112800 51190
rect 112950 51060 113050 51190
rect 113200 51060 113300 51190
rect 113450 51060 113550 51190
rect 113700 51060 113800 51190
rect 113950 51060 114050 51190
rect 114200 51060 114300 51190
rect 114450 51060 114550 51190
rect 114700 51060 114800 51190
rect 114950 51060 115050 51190
rect 115200 51060 115300 51190
rect 115450 51060 115550 51190
rect 115700 51060 115800 51190
rect 115950 51060 116000 51190
rect 89000 51050 89060 51060
rect 89190 51050 89310 51060
rect 89440 51050 89560 51060
rect 89690 51050 89810 51060
rect 89940 51050 90060 51060
rect 90190 51050 90310 51060
rect 90440 51050 90560 51060
rect 90690 51050 90810 51060
rect 90940 51050 91060 51060
rect 91190 51050 91310 51060
rect 91440 51050 91560 51060
rect 91690 51050 91810 51060
rect 91940 51050 92060 51060
rect 92190 51050 92310 51060
rect 92440 51050 92560 51060
rect 92690 51050 92810 51060
rect 92940 51050 93060 51060
rect 93190 51050 93310 51060
rect 93440 51050 93560 51060
rect 93690 51050 93810 51060
rect 93940 51050 94060 51060
rect 94190 51050 94310 51060
rect 94440 51050 94560 51060
rect 94690 51050 94810 51060
rect 94940 51050 95060 51060
rect 95190 51050 95310 51060
rect 95440 51050 95560 51060
rect 95690 51050 95810 51060
rect 95940 51050 96060 51060
rect 96190 51050 96310 51060
rect 96440 51050 96560 51060
rect 96690 51050 96810 51060
rect 96940 51050 97060 51060
rect 97190 51050 97310 51060
rect 97440 51050 97560 51060
rect 97690 51050 97810 51060
rect 97940 51050 98060 51060
rect 98190 51050 98310 51060
rect 98440 51050 98560 51060
rect 98690 51050 98810 51060
rect 98940 51050 99060 51060
rect 99190 51050 99310 51060
rect 99440 51050 99560 51060
rect 99690 51050 99810 51060
rect 99940 51050 100060 51060
rect 100190 51050 100310 51060
rect 100440 51050 100560 51060
rect 100690 51050 100810 51060
rect 100940 51050 101060 51060
rect 101190 51050 101310 51060
rect 101440 51050 101560 51060
rect 101690 51050 101810 51060
rect 101940 51050 102060 51060
rect 102190 51050 102310 51060
rect 102440 51050 102560 51060
rect 102690 51050 102810 51060
rect 102940 51050 103060 51060
rect 103190 51050 103310 51060
rect 103440 51050 103560 51060
rect 103690 51050 103810 51060
rect 103940 51050 104060 51060
rect 104190 51050 104310 51060
rect 104440 51050 104560 51060
rect 104690 51050 104810 51060
rect 104940 51050 105060 51060
rect 105190 51050 105310 51060
rect 105440 51050 105560 51060
rect 105690 51050 105810 51060
rect 105940 51050 106060 51060
rect 106190 51050 106310 51060
rect 106440 51050 106560 51060
rect 106690 51050 106810 51060
rect 106940 51050 107060 51060
rect 107190 51050 107310 51060
rect 107440 51050 107560 51060
rect 107690 51050 107810 51060
rect 107940 51050 108060 51060
rect 108190 51050 108310 51060
rect 108440 51050 108560 51060
rect 108690 51050 108810 51060
rect 108940 51050 109060 51060
rect 109190 51050 109310 51060
rect 109440 51050 109560 51060
rect 109690 51050 109810 51060
rect 109940 51050 110060 51060
rect 110190 51050 110310 51060
rect 110440 51050 110560 51060
rect 110690 51050 110810 51060
rect 110940 51050 111060 51060
rect 111190 51050 111310 51060
rect 111440 51050 111560 51060
rect 111690 51050 111810 51060
rect 111940 51050 112060 51060
rect 112190 51050 112310 51060
rect 112440 51050 112560 51060
rect 112690 51050 112810 51060
rect 112940 51050 113060 51060
rect 113190 51050 113310 51060
rect 113440 51050 113560 51060
rect 113690 51050 113810 51060
rect 113940 51050 114060 51060
rect 114190 51050 114310 51060
rect 114440 51050 114560 51060
rect 114690 51050 114810 51060
rect 114940 51050 115060 51060
rect 115190 51050 115310 51060
rect 115440 51050 115560 51060
rect 115690 51050 115810 51060
rect 115940 51050 116000 51060
rect 89000 51000 116000 51050
<< metal3 >>
rect 8000 60900 11000 62000
rect 34097 61900 36597 62000
rect 34097 61150 36600 61900
rect 34100 61000 36600 61150
rect 8000 58100 8100 60900
rect 10900 58100 11000 60900
rect 8000 58000 11000 58100
rect 60000 60900 63000 62000
rect 82797 61150 85297 62000
rect 85447 61150 86547 62000
rect 86697 61150 87797 62000
rect 87947 61150 90447 62000
rect 108647 61150 111147 62000
rect 111297 61150 112397 62000
rect 112547 61150 113647 62000
rect 113797 61150 116297 62000
rect 159497 61150 161997 62000
rect 162147 61150 163247 62000
rect 163397 61150 164497 62000
rect 164647 61150 167147 62000
rect 206697 61150 209197 62000
rect 232697 61800 235200 62000
rect 232697 61150 232800 61800
rect 60000 58100 60100 60900
rect 62900 58100 63000 60900
rect 60000 58000 63000 58100
rect 83000 60900 85000 61150
rect 83000 57600 83100 60900
rect 84900 57600 85000 60900
rect 83000 57500 85000 57600
rect 109000 60900 111000 61150
rect 109000 57600 109100 60900
rect 110900 57600 111000 60900
rect 232700 60700 232800 61150
rect 234900 60700 235200 61800
rect 255297 61600 257697 62000
rect 255297 61170 257700 61600
rect 260297 61170 262697 62000
rect 232700 60600 235200 60700
rect 255300 61100 257700 61170
rect 283297 61150 285797 62000
rect 255300 58100 255400 61100
rect 257600 58100 257700 61100
rect 255300 57900 257700 58100
rect 109000 57500 111000 57600
rect 0 50121 850 52621
rect 291150 48992 292000 51492
rect 0 31921 830 34321
rect 291170 29892 292000 32292
rect 0 26921 830 29321
rect 291170 24892 292000 27292
rect 291760 4736 292400 4792
rect 291760 4145 292400 4201
rect 291760 3554 292400 3610
rect 291760 2963 292400 3019
rect 291760 2372 292400 2428
rect 291760 1781 292400 1837
rect 10000 0 10056 200
rect 13100 0 13156 200
rect 16200 0 16256 200
rect 19300 0 19356 200
rect 22400 0 22456 200
rect 25500 0 25556 200
rect 28600 0 28656 200
rect 31700 0 31756 200
rect 34800 0 34856 200
rect 37900 0 37956 200
rect 41000 0 41056 200
rect 44100 0 44156 200
rect 47200 0 47256 200
rect 50300 0 50356 200
rect 53400 0 53456 200
rect 56500 0 56556 200
rect 59600 0 59656 200
rect 62700 0 62756 200
rect 65800 0 65856 200
rect 68900 0 68956 200
rect 72000 0 72056 200
rect 75100 0 75156 200
rect 78200 0 78256 200
rect 81300 0 81356 200
rect 84400 0 84456 200
rect 87500 0 87556 200
rect 90600 0 90656 200
rect 93700 0 93756 200
rect 96800 0 96856 200
rect 99900 0 99956 200
rect 103000 0 103056 200
rect 106100 0 106156 200
rect 109200 0 109256 200
rect 112300 0 112356 200
rect 115400 0 115456 200
rect 118500 0 118556 200
rect 121600 0 121656 200
rect 124700 0 124756 200
rect 127800 0 127856 200
rect 130900 0 130956 200
rect 134000 0 134056 200
rect 137100 0 137156 200
rect 140200 0 140256 200
rect 143300 0 143356 200
rect 146400 0 146456 200
rect 149500 0 149556 200
rect 152600 0 152656 200
rect 155700 0 155756 200
rect 158800 0 158856 200
rect 161900 0 161956 200
rect 165000 0 165056 200
rect 168100 0 168156 200
rect 171200 0 171256 200
rect 174300 0 174356 200
rect 177400 0 177456 200
rect 180500 0 180556 200
rect 183600 0 183656 200
rect 186700 0 186756 200
rect 189800 0 189856 200
rect 192900 0 192956 200
rect 0 -10279 830 -7879
rect 0 -15279 830 -12879
rect 291170 -14719 292000 -12319
rect 291170 -19719 292000 -17319
<< via3 >>
rect 8100 58100 10900 60900
rect 60100 58100 62900 60900
rect 83100 57600 84900 60900
rect 109100 57600 110900 60900
rect 232800 60700 234900 61800
rect 255400 58100 257600 61100
<< metal4 >>
rect 232700 61800 235000 61900
rect 8000 60900 11000 61000
rect 8000 58100 8100 60900
rect 10900 58100 11000 60900
rect 8000 58000 11000 58100
rect 60000 60900 63000 61000
rect 60000 58100 60100 60900
rect 62900 58100 63000 60900
rect 60000 58000 63000 58100
rect 83000 60900 85000 61000
rect 83000 57600 83100 60900
rect 84900 57600 85000 60900
rect 83000 55000 85000 57600
rect 109000 60900 111000 61000
rect 109000 57600 109100 60900
rect 110900 57600 111000 60900
rect 232700 60700 232800 61800
rect 234900 60700 235000 61800
rect 232700 60600 235000 60700
rect 255300 61100 257700 61200
rect 255300 58100 255400 61100
rect 257600 58100 257700 61100
rect 255300 57900 257700 58100
rect 109000 54000 111000 57600
rect 85000 52500 111000 54000
rect 3049 0 6899 400
rect 7229 0 11079 400
rect 282049 0 285899 400
rect 286229 0 290079 400
<< via4 >>
rect 8100 58100 10900 60900
rect 60100 58100 62900 60900
rect 232800 60700 234900 61800
<< metal5 >>
rect 232700 61800 235000 61900
rect 8000 60900 11000 61000
rect 8000 58100 8100 60900
rect 10900 60000 11000 60900
rect 60000 60900 63000 61000
rect 10900 58100 28000 60000
rect 8000 58000 28000 58100
rect 60000 58100 60100 60900
rect 62900 60000 63000 60900
rect 232700 60700 232800 61800
rect 234900 60700 235000 61800
rect 232700 60600 235000 60700
rect 62900 58100 69000 60000
rect 233000 59900 234700 60600
rect 60000 58000 69000 58100
rect 26000 55000 28000 58000
rect 67000 55000 69000 58000
use RX_top  RX_top_0
timestamp 1662171338
transform 1 0 19000 0 -1 50000
box -18500 -11900 84000 49800
use TX_top  TX_top_0
timestamp 1662096097
transform 1 0 219650 0 -1 41900
box -41750 -18100 48250 27950
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501637
transform 1 0 5000 0 -1 61000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_38
timestamp 1659501637
transform 1 0 5000 0 -1 59000
box 0 0 2000 2000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660792292
transform 1 0 33000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_1
timestamp 1660792292
transform 1 0 37000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_2
timestamp 1660792292
transform 1 0 41000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_3
timestamp 1660792292
transform 1 0 45000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_4
timestamp 1660792292
transform 1 0 49000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_5
timestamp 1660792292
transform 1 0 53000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_6
timestamp 1660792292
transform 1 0 55000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_7
timestamp 1660792292
transform 1 0 71000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_8
timestamp 1660792292
transform 1 0 75000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_9
timestamp 1660792292
transform 1 0 77000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_10
timestamp 1660792292
transform 1 0 97000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_11
timestamp 1660792292
transform 1 0 93000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_12
timestamp 1660792292
transform 1 0 91000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_13
timestamp 1660792292
transform 1 0 101000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_14
timestamp 1660792292
transform 1 0 103000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_70
timestamp 1660792292
transform 1 0 29000 0 -1 61000
box 0 0 4000 4000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1662168084
transform 1 0 103000 0 1 43000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_1
timestamp 1662168084
transform 1 0 111000 0 1 43000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_2
timestamp 1662168084
transform 1 0 111000 0 1 35000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_3
timestamp 1662168084
transform 1 0 103000 0 1 35000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_4
timestamp 1662168084
transform 1 0 111000 0 1 27000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_5
timestamp 1662168084
transform 1 0 103000 0 1 27000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_6
timestamp 1662168084
transform 1 0 111000 0 1 19000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_7
timestamp 1662168084
transform 1 0 103000 0 1 19000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_8
timestamp 1662168084
transform 1 0 111000 0 1 11000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_9
timestamp 1662168084
transform 1 0 103000 0 1 11000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_10
timestamp 1662168084
transform 1 0 103000 0 1 3000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_11
timestamp 1662168084
transform 1 0 111000 0 1 3000
box 0 0 8000 8000
<< labels >>
rlabel metal3 s 10000 0 10056 200 0 analog_la_out[0]
port 1 nsew
rlabel metal3 s 13100 0 13156 200 0 analog_la_out[1]
port 2 nsew
rlabel metal3 s 16200 0 16256 200 0 analog_la_out[2]
port 3 nsew
rlabel metal3 s 19300 0 19356 200 0 analog_la_out[3]
port 4 nsew
rlabel metal3 s 22400 0 22456 200 0 analog_la_out[4]
port 5 nsew
rlabel metal3 s 25500 0 25556 200 0 analog_la_out[5]
port 6 nsew
rlabel metal3 s 28600 0 28656 200 0 analog_la_out[6]
port 7 nsew
rlabel metal3 s 31700 0 31756 200 0 analog_la_out[7]
port 8 nsew
rlabel metal3 s 34800 0 34856 200 0 analog_la_out[8]
port 9 nsew
rlabel metal3 s 37900 0 37956 200 0 analog_la_out[9]
port 10 nsew
rlabel metal3 s 41000 0 41056 200 0 analog_la_out[10]
port 11 nsew
rlabel metal3 s 44100 0 44156 200 0 analog_la_out[11]
port 12 nsew
rlabel metal3 s 47200 0 47256 200 0 analog_la_out[12]
port 13 nsew
rlabel metal3 s 50300 0 50356 200 0 analog_la_out[13]
port 14 nsew
rlabel metal3 s 53400 0 53456 200 0 analog_la_out[14]
port 15 nsew
rlabel metal3 s 56500 0 56556 200 0 analog_la_out[15]
port 16 nsew
rlabel metal3 s 59600 0 59656 200 0 analog_la_out[16]
port 17 nsew
rlabel metal3 s 62700 0 62756 200 0 analog_la_out[17]
port 18 nsew
rlabel metal3 s 65800 0 65856 200 0 analog_la_out[18]
port 19 nsew
rlabel metal3 s 68900 0 68956 200 0 analog_la_out[19]
port 20 nsew
rlabel metal3 s 72000 0 72056 200 0 analog_la_out[20]
port 21 nsew
rlabel metal3 s 75100 0 75156 200 0 analog_la_out[21]
port 22 nsew
rlabel metal3 s 78200 0 78256 200 0 analog_la_out[22]
port 23 nsew
rlabel metal3 s 81300 0 81356 200 0 analog_la_out[23]
port 24 nsew
rlabel metal3 s 84400 0 84456 200 0 analog_la_out[24]
port 25 nsew
rlabel metal3 s 87500 0 87556 200 0 analog_la_out[25]
port 26 nsew
rlabel metal3 s 90600 0 90656 200 0 analog_la_out[26]
port 27 nsew
rlabel metal3 s 93700 0 93756 200 0 analog_la_out[27]
port 28 nsew
rlabel metal3 s 96800 0 96856 200 0 analog_la_out[28]
port 29 nsew
rlabel metal3 s 99900 0 99956 200 0 analog_la_out[29]
port 30 nsew
rlabel metal3 s 103000 0 103056 200 0 analog_la_in[0]
port 31 nsew
rlabel metal3 s 106100 0 106156 200 0 analog_la_in[1]
port 32 nsew
rlabel metal3 s 109200 0 109256 200 0 analog_la_in[2]
port 33 nsew
rlabel metal3 s 112300 0 112356 200 0 analog_la_in[3]
port 34 nsew
rlabel metal3 s 115400 0 115456 200 0 analog_la_in[4]
port 35 nsew
rlabel metal3 s 118500 0 118556 200 0 analog_la_in[5]
port 36 nsew
rlabel metal3 s 121600 0 121656 200 0 analog_la_in[6]
port 37 nsew
rlabel metal3 s 124700 0 124756 200 0 analog_la_in[7]
port 38 nsew
rlabel metal3 s 127800 0 127856 200 0 analog_la_in[8]
port 39 nsew
rlabel metal3 s 130900 0 130956 200 0 analog_la_in[9]
port 40 nsew
rlabel metal3 s 134000 0 134056 200 0 analog_la_in[10]
port 41 nsew
rlabel metal3 s 137100 0 137156 200 0 analog_la_in[11]
port 42 nsew
rlabel metal3 s 140200 0 140256 200 0 analog_la_in[12]
port 43 nsew
rlabel metal3 s 143300 0 143356 200 0 analog_la_in[13]
port 44 nsew
rlabel metal3 s 146400 0 146456 200 0 analog_la_in[14]
port 45 nsew
rlabel metal3 s 149500 0 149556 200 0 analog_la_in[15]
port 46 nsew
rlabel metal3 s 152600 0 152656 200 0 analog_la_in[16]
port 47 nsew
rlabel metal3 s 155700 0 155756 200 0 analog_la_in[17]
port 48 nsew
rlabel metal3 s 158800 0 158856 200 0 analog_la_in[18]
port 49 nsew
rlabel metal3 s 161900 0 161956 200 0 analog_la_in[19]
port 50 nsew
rlabel metal3 s 165000 0 165056 200 0 analog_la_in[20]
port 51 nsew
rlabel metal3 s 168100 0 168156 200 0 analog_la_in[21]
port 52 nsew
rlabel metal3 s 171200 0 171256 200 0 analog_la_in[22]
port 53 nsew
rlabel metal3 s 174300 0 174356 200 0 analog_la_in[23]
port 54 nsew
rlabel metal3 s 177400 0 177456 200 0 analog_la_in[24]
port 55 nsew
rlabel metal3 s 180500 0 180556 200 0 analog_la_in[25]
port 56 nsew
rlabel metal3 s 183600 0 183656 200 0 analog_la_in[26]
port 57 nsew
rlabel metal3 s 186700 0 186756 200 0 analog_la_in[27]
port 58 nsew
rlabel metal3 s 189800 0 189856 200 0 analog_la_in[28]
port 59 nsew
rlabel metal3 s 192900 0 192956 200 0 analog_la_in[29]
port 60 nsew
rlabel metal4 s 282049 0 285899 400 0 vdda1
port 86 nsew
rlabel metal4 s 286229 0 290079 400 0 vssa1
port 87 nsew
rlabel metal4 s 3049 0 6899 400 0 vdda2
port 89 nsew
rlabel metal4 s 7229 0 11079 400 0 vssd2
port 90 nsew
rlabel metal3 s 291760 1781 292400 1837 0 gpio_analog[6]
port 61 nsew
rlabel metal3 s 291760 2372 292400 2428 0 gpio_noesd[6]
port 62 nsew
rlabel metal3 s 291150 48992 292000 51492 0 io_analog[0]
port 63 nsew
rlabel metal3 s 0 50121 850 52621 0 io_analog[10]
port 64 nsew
rlabel metal3 s 283297 61150 285797 62000 0 io_analog[1]
port 65 nsew
rlabel metal3 s 232697 61150 235197 62000 0 io_analog[2]
port 66 nsew
rlabel metal3 s 206697 61150 209197 62000 0 io_analog[3]
port 67 nsew
rlabel metal3 s 159497 61150 161997 62000 0 io_analog[4]
port 68 nsew
rlabel metal3 s 108647 61150 111147 62000 0 io_analog[5]
port 69 nsew
rlabel metal3 s 82797 61150 85297 62000 0 io_analog[6]
port 70 nsew
rlabel metal3 s 60097 61150 62597 62000 0 io_analog[7]
port 71 nsew
rlabel metal3 s 34097 61150 36597 62000 0 io_analog[8]
port 72 nsew
rlabel metal3 s 8097 61150 10597 62000 0 io_analog[9]
port 73 nsew
rlabel metal3 s 163397 61150 164497 62000 0 io_clamp_high[0]
port 74 nsew
rlabel metal3 s 112547 61150 113647 62000 0 io_clamp_high[1]
port 75 nsew
rlabel metal3 s 86697 61150 87797 62000 0 io_clamp_high[2]
port 76 nsew
rlabel metal3 s 162147 61150 163247 62000 0 io_clamp_low[0]
port 77 nsew
rlabel metal3 s 111297 61150 112397 62000 0 io_clamp_low[1]
port 78 nsew
rlabel metal3 s 85447 61150 86547 62000 0 io_clamp_low[2]
port 79 nsew
rlabel metal3 s 291760 3554 292400 3610 0 io_in[13]
port 80 nsew
rlabel metal3 s 291760 2963 292400 3019 0 io_in_3v3[13]
port 81 nsew
rlabel metal3 s 291760 4736 292400 4792 0 io_oeb[13]
port 82 nsew
rlabel metal3 s 291760 4145 292400 4201 0 io_out[13]
port 83 nsew
rlabel metal3 s 291170 24892 292000 27292 0 vccd1
port 84 nsew
rlabel metal3 s 0 26921 830 29321 0 vccd2
port 85 nsew
rlabel metal3 s 291170 -14719 292000 -12319 0 vdda1
port 86 nsew
rlabel metal3 s 255297 61170 257697 62000 0 vssa1
port 87 nsew
rlabel metal3 s 0 -15279 830 -12879 0 vssa2
port 88 nsew
<< properties >>
string FIXED_BBOX 0 0 292000 82000
string path 1929.280 0.000 1929.280 2.000 
<< end >>
