magic
tech sky130B
magscale 1 2
timestamp 1661374315
<< pwell >>
rect 0 126 2474 1188
<< nmos >>
rect 194 152 224 1162
rect 280 152 310 1162
rect 588 152 618 1162
rect 674 152 704 1162
rect 982 152 1012 1162
rect 1068 152 1098 1162
rect 1376 152 1406 1162
rect 1462 152 1492 1162
rect 1770 152 1800 1162
rect 1856 152 1886 1162
rect 2164 152 2194 1162
rect 2250 152 2280 1162
<< ndiff >>
rect 138 1150 194 1162
rect 138 1116 149 1150
rect 183 1116 194 1150
rect 138 1082 194 1116
rect 138 1048 149 1082
rect 183 1048 194 1082
rect 138 1014 194 1048
rect 138 980 149 1014
rect 183 980 194 1014
rect 138 946 194 980
rect 138 912 149 946
rect 183 912 194 946
rect 138 878 194 912
rect 138 844 149 878
rect 183 844 194 878
rect 138 810 194 844
rect 138 776 149 810
rect 183 776 194 810
rect 138 742 194 776
rect 138 708 149 742
rect 183 708 194 742
rect 138 674 194 708
rect 138 640 149 674
rect 183 640 194 674
rect 138 606 194 640
rect 138 572 149 606
rect 183 572 194 606
rect 138 538 194 572
rect 138 504 149 538
rect 183 504 194 538
rect 138 470 194 504
rect 138 436 149 470
rect 183 436 194 470
rect 138 402 194 436
rect 138 368 149 402
rect 183 368 194 402
rect 138 334 194 368
rect 138 300 149 334
rect 183 300 194 334
rect 138 266 194 300
rect 138 232 149 266
rect 183 232 194 266
rect 138 198 194 232
rect 138 164 149 198
rect 183 164 194 198
rect 138 152 194 164
rect 224 1150 280 1162
rect 224 1116 235 1150
rect 269 1116 280 1150
rect 224 1082 280 1116
rect 224 1048 235 1082
rect 269 1048 280 1082
rect 224 1014 280 1048
rect 224 980 235 1014
rect 269 980 280 1014
rect 224 946 280 980
rect 224 912 235 946
rect 269 912 280 946
rect 224 878 280 912
rect 224 844 235 878
rect 269 844 280 878
rect 224 810 280 844
rect 224 776 235 810
rect 269 776 280 810
rect 224 742 280 776
rect 224 708 235 742
rect 269 708 280 742
rect 224 674 280 708
rect 224 640 235 674
rect 269 640 280 674
rect 224 606 280 640
rect 224 572 235 606
rect 269 572 280 606
rect 224 538 280 572
rect 224 504 235 538
rect 269 504 280 538
rect 224 470 280 504
rect 224 436 235 470
rect 269 436 280 470
rect 224 402 280 436
rect 224 368 235 402
rect 269 368 280 402
rect 224 334 280 368
rect 224 300 235 334
rect 269 300 280 334
rect 224 266 280 300
rect 224 232 235 266
rect 269 232 280 266
rect 224 198 280 232
rect 224 164 235 198
rect 269 164 280 198
rect 224 152 280 164
rect 310 1150 366 1162
rect 310 1116 321 1150
rect 355 1116 366 1150
rect 310 1082 366 1116
rect 310 1048 321 1082
rect 355 1048 366 1082
rect 310 1014 366 1048
rect 310 980 321 1014
rect 355 980 366 1014
rect 310 946 366 980
rect 310 912 321 946
rect 355 912 366 946
rect 310 878 366 912
rect 310 844 321 878
rect 355 844 366 878
rect 310 810 366 844
rect 310 776 321 810
rect 355 776 366 810
rect 310 742 366 776
rect 310 708 321 742
rect 355 708 366 742
rect 310 674 366 708
rect 310 640 321 674
rect 355 640 366 674
rect 310 606 366 640
rect 310 572 321 606
rect 355 572 366 606
rect 310 538 366 572
rect 310 504 321 538
rect 355 504 366 538
rect 310 470 366 504
rect 310 436 321 470
rect 355 436 366 470
rect 310 402 366 436
rect 310 368 321 402
rect 355 368 366 402
rect 310 334 366 368
rect 310 300 321 334
rect 355 300 366 334
rect 310 266 366 300
rect 310 232 321 266
rect 355 232 366 266
rect 310 198 366 232
rect 310 164 321 198
rect 355 164 366 198
rect 310 152 366 164
rect 532 1150 588 1162
rect 532 1116 543 1150
rect 577 1116 588 1150
rect 532 1082 588 1116
rect 532 1048 543 1082
rect 577 1048 588 1082
rect 532 1014 588 1048
rect 532 980 543 1014
rect 577 980 588 1014
rect 532 946 588 980
rect 532 912 543 946
rect 577 912 588 946
rect 532 878 588 912
rect 532 844 543 878
rect 577 844 588 878
rect 532 810 588 844
rect 532 776 543 810
rect 577 776 588 810
rect 532 742 588 776
rect 532 708 543 742
rect 577 708 588 742
rect 532 674 588 708
rect 532 640 543 674
rect 577 640 588 674
rect 532 606 588 640
rect 532 572 543 606
rect 577 572 588 606
rect 532 538 588 572
rect 532 504 543 538
rect 577 504 588 538
rect 532 470 588 504
rect 532 436 543 470
rect 577 436 588 470
rect 532 402 588 436
rect 532 368 543 402
rect 577 368 588 402
rect 532 334 588 368
rect 532 300 543 334
rect 577 300 588 334
rect 532 266 588 300
rect 532 232 543 266
rect 577 232 588 266
rect 532 198 588 232
rect 532 164 543 198
rect 577 164 588 198
rect 532 152 588 164
rect 618 1150 674 1162
rect 618 1116 629 1150
rect 663 1116 674 1150
rect 618 1082 674 1116
rect 618 1048 629 1082
rect 663 1048 674 1082
rect 618 1014 674 1048
rect 618 980 629 1014
rect 663 980 674 1014
rect 618 946 674 980
rect 618 912 629 946
rect 663 912 674 946
rect 618 878 674 912
rect 618 844 629 878
rect 663 844 674 878
rect 618 810 674 844
rect 618 776 629 810
rect 663 776 674 810
rect 618 742 674 776
rect 618 708 629 742
rect 663 708 674 742
rect 618 674 674 708
rect 618 640 629 674
rect 663 640 674 674
rect 618 606 674 640
rect 618 572 629 606
rect 663 572 674 606
rect 618 538 674 572
rect 618 504 629 538
rect 663 504 674 538
rect 618 470 674 504
rect 618 436 629 470
rect 663 436 674 470
rect 618 402 674 436
rect 618 368 629 402
rect 663 368 674 402
rect 618 334 674 368
rect 618 300 629 334
rect 663 300 674 334
rect 618 266 674 300
rect 618 232 629 266
rect 663 232 674 266
rect 618 198 674 232
rect 618 164 629 198
rect 663 164 674 198
rect 618 152 674 164
rect 704 1150 760 1162
rect 704 1116 715 1150
rect 749 1116 760 1150
rect 704 1082 760 1116
rect 704 1048 715 1082
rect 749 1048 760 1082
rect 704 1014 760 1048
rect 704 980 715 1014
rect 749 980 760 1014
rect 704 946 760 980
rect 704 912 715 946
rect 749 912 760 946
rect 704 878 760 912
rect 704 844 715 878
rect 749 844 760 878
rect 704 810 760 844
rect 704 776 715 810
rect 749 776 760 810
rect 704 742 760 776
rect 704 708 715 742
rect 749 708 760 742
rect 704 674 760 708
rect 704 640 715 674
rect 749 640 760 674
rect 704 606 760 640
rect 704 572 715 606
rect 749 572 760 606
rect 704 538 760 572
rect 704 504 715 538
rect 749 504 760 538
rect 704 470 760 504
rect 704 436 715 470
rect 749 436 760 470
rect 704 402 760 436
rect 704 368 715 402
rect 749 368 760 402
rect 704 334 760 368
rect 704 300 715 334
rect 749 300 760 334
rect 704 266 760 300
rect 704 232 715 266
rect 749 232 760 266
rect 704 198 760 232
rect 704 164 715 198
rect 749 164 760 198
rect 704 152 760 164
rect 926 1150 982 1162
rect 926 1116 937 1150
rect 971 1116 982 1150
rect 926 1082 982 1116
rect 926 1048 937 1082
rect 971 1048 982 1082
rect 926 1014 982 1048
rect 926 980 937 1014
rect 971 980 982 1014
rect 926 946 982 980
rect 926 912 937 946
rect 971 912 982 946
rect 926 878 982 912
rect 926 844 937 878
rect 971 844 982 878
rect 926 810 982 844
rect 926 776 937 810
rect 971 776 982 810
rect 926 742 982 776
rect 926 708 937 742
rect 971 708 982 742
rect 926 674 982 708
rect 926 640 937 674
rect 971 640 982 674
rect 926 606 982 640
rect 926 572 937 606
rect 971 572 982 606
rect 926 538 982 572
rect 926 504 937 538
rect 971 504 982 538
rect 926 470 982 504
rect 926 436 937 470
rect 971 436 982 470
rect 926 402 982 436
rect 926 368 937 402
rect 971 368 982 402
rect 926 334 982 368
rect 926 300 937 334
rect 971 300 982 334
rect 926 266 982 300
rect 926 232 937 266
rect 971 232 982 266
rect 926 198 982 232
rect 926 164 937 198
rect 971 164 982 198
rect 926 152 982 164
rect 1012 1150 1068 1162
rect 1012 1116 1023 1150
rect 1057 1116 1068 1150
rect 1012 1082 1068 1116
rect 1012 1048 1023 1082
rect 1057 1048 1068 1082
rect 1012 1014 1068 1048
rect 1012 980 1023 1014
rect 1057 980 1068 1014
rect 1012 946 1068 980
rect 1012 912 1023 946
rect 1057 912 1068 946
rect 1012 878 1068 912
rect 1012 844 1023 878
rect 1057 844 1068 878
rect 1012 810 1068 844
rect 1012 776 1023 810
rect 1057 776 1068 810
rect 1012 742 1068 776
rect 1012 708 1023 742
rect 1057 708 1068 742
rect 1012 674 1068 708
rect 1012 640 1023 674
rect 1057 640 1068 674
rect 1012 606 1068 640
rect 1012 572 1023 606
rect 1057 572 1068 606
rect 1012 538 1068 572
rect 1012 504 1023 538
rect 1057 504 1068 538
rect 1012 470 1068 504
rect 1012 436 1023 470
rect 1057 436 1068 470
rect 1012 402 1068 436
rect 1012 368 1023 402
rect 1057 368 1068 402
rect 1012 334 1068 368
rect 1012 300 1023 334
rect 1057 300 1068 334
rect 1012 266 1068 300
rect 1012 232 1023 266
rect 1057 232 1068 266
rect 1012 198 1068 232
rect 1012 164 1023 198
rect 1057 164 1068 198
rect 1012 152 1068 164
rect 1098 1150 1154 1162
rect 1098 1116 1109 1150
rect 1143 1116 1154 1150
rect 1098 1082 1154 1116
rect 1098 1048 1109 1082
rect 1143 1048 1154 1082
rect 1098 1014 1154 1048
rect 1098 980 1109 1014
rect 1143 980 1154 1014
rect 1098 946 1154 980
rect 1098 912 1109 946
rect 1143 912 1154 946
rect 1098 878 1154 912
rect 1098 844 1109 878
rect 1143 844 1154 878
rect 1098 810 1154 844
rect 1098 776 1109 810
rect 1143 776 1154 810
rect 1098 742 1154 776
rect 1098 708 1109 742
rect 1143 708 1154 742
rect 1098 674 1154 708
rect 1098 640 1109 674
rect 1143 640 1154 674
rect 1098 606 1154 640
rect 1098 572 1109 606
rect 1143 572 1154 606
rect 1098 538 1154 572
rect 1098 504 1109 538
rect 1143 504 1154 538
rect 1098 470 1154 504
rect 1098 436 1109 470
rect 1143 436 1154 470
rect 1098 402 1154 436
rect 1098 368 1109 402
rect 1143 368 1154 402
rect 1098 334 1154 368
rect 1098 300 1109 334
rect 1143 300 1154 334
rect 1098 266 1154 300
rect 1098 232 1109 266
rect 1143 232 1154 266
rect 1098 198 1154 232
rect 1098 164 1109 198
rect 1143 164 1154 198
rect 1098 152 1154 164
rect 1320 1150 1376 1162
rect 1320 1116 1331 1150
rect 1365 1116 1376 1150
rect 1320 1082 1376 1116
rect 1320 1048 1331 1082
rect 1365 1048 1376 1082
rect 1320 1014 1376 1048
rect 1320 980 1331 1014
rect 1365 980 1376 1014
rect 1320 946 1376 980
rect 1320 912 1331 946
rect 1365 912 1376 946
rect 1320 878 1376 912
rect 1320 844 1331 878
rect 1365 844 1376 878
rect 1320 810 1376 844
rect 1320 776 1331 810
rect 1365 776 1376 810
rect 1320 742 1376 776
rect 1320 708 1331 742
rect 1365 708 1376 742
rect 1320 674 1376 708
rect 1320 640 1331 674
rect 1365 640 1376 674
rect 1320 606 1376 640
rect 1320 572 1331 606
rect 1365 572 1376 606
rect 1320 538 1376 572
rect 1320 504 1331 538
rect 1365 504 1376 538
rect 1320 470 1376 504
rect 1320 436 1331 470
rect 1365 436 1376 470
rect 1320 402 1376 436
rect 1320 368 1331 402
rect 1365 368 1376 402
rect 1320 334 1376 368
rect 1320 300 1331 334
rect 1365 300 1376 334
rect 1320 266 1376 300
rect 1320 232 1331 266
rect 1365 232 1376 266
rect 1320 198 1376 232
rect 1320 164 1331 198
rect 1365 164 1376 198
rect 1320 152 1376 164
rect 1406 1150 1462 1162
rect 1406 1116 1417 1150
rect 1451 1116 1462 1150
rect 1406 1082 1462 1116
rect 1406 1048 1417 1082
rect 1451 1048 1462 1082
rect 1406 1014 1462 1048
rect 1406 980 1417 1014
rect 1451 980 1462 1014
rect 1406 946 1462 980
rect 1406 912 1417 946
rect 1451 912 1462 946
rect 1406 878 1462 912
rect 1406 844 1417 878
rect 1451 844 1462 878
rect 1406 810 1462 844
rect 1406 776 1417 810
rect 1451 776 1462 810
rect 1406 742 1462 776
rect 1406 708 1417 742
rect 1451 708 1462 742
rect 1406 674 1462 708
rect 1406 640 1417 674
rect 1451 640 1462 674
rect 1406 606 1462 640
rect 1406 572 1417 606
rect 1451 572 1462 606
rect 1406 538 1462 572
rect 1406 504 1417 538
rect 1451 504 1462 538
rect 1406 470 1462 504
rect 1406 436 1417 470
rect 1451 436 1462 470
rect 1406 402 1462 436
rect 1406 368 1417 402
rect 1451 368 1462 402
rect 1406 334 1462 368
rect 1406 300 1417 334
rect 1451 300 1462 334
rect 1406 266 1462 300
rect 1406 232 1417 266
rect 1451 232 1462 266
rect 1406 198 1462 232
rect 1406 164 1417 198
rect 1451 164 1462 198
rect 1406 152 1462 164
rect 1492 1150 1548 1162
rect 1492 1116 1503 1150
rect 1537 1116 1548 1150
rect 1492 1082 1548 1116
rect 1492 1048 1503 1082
rect 1537 1048 1548 1082
rect 1492 1014 1548 1048
rect 1492 980 1503 1014
rect 1537 980 1548 1014
rect 1492 946 1548 980
rect 1492 912 1503 946
rect 1537 912 1548 946
rect 1492 878 1548 912
rect 1492 844 1503 878
rect 1537 844 1548 878
rect 1492 810 1548 844
rect 1492 776 1503 810
rect 1537 776 1548 810
rect 1492 742 1548 776
rect 1492 708 1503 742
rect 1537 708 1548 742
rect 1492 674 1548 708
rect 1492 640 1503 674
rect 1537 640 1548 674
rect 1492 606 1548 640
rect 1492 572 1503 606
rect 1537 572 1548 606
rect 1492 538 1548 572
rect 1492 504 1503 538
rect 1537 504 1548 538
rect 1492 470 1548 504
rect 1492 436 1503 470
rect 1537 436 1548 470
rect 1492 402 1548 436
rect 1492 368 1503 402
rect 1537 368 1548 402
rect 1492 334 1548 368
rect 1492 300 1503 334
rect 1537 300 1548 334
rect 1492 266 1548 300
rect 1492 232 1503 266
rect 1537 232 1548 266
rect 1492 198 1548 232
rect 1492 164 1503 198
rect 1537 164 1548 198
rect 1492 152 1548 164
rect 1714 1150 1770 1162
rect 1714 1116 1725 1150
rect 1759 1116 1770 1150
rect 1714 1082 1770 1116
rect 1714 1048 1725 1082
rect 1759 1048 1770 1082
rect 1714 1014 1770 1048
rect 1714 980 1725 1014
rect 1759 980 1770 1014
rect 1714 946 1770 980
rect 1714 912 1725 946
rect 1759 912 1770 946
rect 1714 878 1770 912
rect 1714 844 1725 878
rect 1759 844 1770 878
rect 1714 810 1770 844
rect 1714 776 1725 810
rect 1759 776 1770 810
rect 1714 742 1770 776
rect 1714 708 1725 742
rect 1759 708 1770 742
rect 1714 674 1770 708
rect 1714 640 1725 674
rect 1759 640 1770 674
rect 1714 606 1770 640
rect 1714 572 1725 606
rect 1759 572 1770 606
rect 1714 538 1770 572
rect 1714 504 1725 538
rect 1759 504 1770 538
rect 1714 470 1770 504
rect 1714 436 1725 470
rect 1759 436 1770 470
rect 1714 402 1770 436
rect 1714 368 1725 402
rect 1759 368 1770 402
rect 1714 334 1770 368
rect 1714 300 1725 334
rect 1759 300 1770 334
rect 1714 266 1770 300
rect 1714 232 1725 266
rect 1759 232 1770 266
rect 1714 198 1770 232
rect 1714 164 1725 198
rect 1759 164 1770 198
rect 1714 152 1770 164
rect 1800 1150 1856 1162
rect 1800 1116 1811 1150
rect 1845 1116 1856 1150
rect 1800 1082 1856 1116
rect 1800 1048 1811 1082
rect 1845 1048 1856 1082
rect 1800 1014 1856 1048
rect 1800 980 1811 1014
rect 1845 980 1856 1014
rect 1800 946 1856 980
rect 1800 912 1811 946
rect 1845 912 1856 946
rect 1800 878 1856 912
rect 1800 844 1811 878
rect 1845 844 1856 878
rect 1800 810 1856 844
rect 1800 776 1811 810
rect 1845 776 1856 810
rect 1800 742 1856 776
rect 1800 708 1811 742
rect 1845 708 1856 742
rect 1800 674 1856 708
rect 1800 640 1811 674
rect 1845 640 1856 674
rect 1800 606 1856 640
rect 1800 572 1811 606
rect 1845 572 1856 606
rect 1800 538 1856 572
rect 1800 504 1811 538
rect 1845 504 1856 538
rect 1800 470 1856 504
rect 1800 436 1811 470
rect 1845 436 1856 470
rect 1800 402 1856 436
rect 1800 368 1811 402
rect 1845 368 1856 402
rect 1800 334 1856 368
rect 1800 300 1811 334
rect 1845 300 1856 334
rect 1800 266 1856 300
rect 1800 232 1811 266
rect 1845 232 1856 266
rect 1800 198 1856 232
rect 1800 164 1811 198
rect 1845 164 1856 198
rect 1800 152 1856 164
rect 1886 1150 1942 1162
rect 1886 1116 1897 1150
rect 1931 1116 1942 1150
rect 1886 1082 1942 1116
rect 1886 1048 1897 1082
rect 1931 1048 1942 1082
rect 1886 1014 1942 1048
rect 1886 980 1897 1014
rect 1931 980 1942 1014
rect 1886 946 1942 980
rect 1886 912 1897 946
rect 1931 912 1942 946
rect 1886 878 1942 912
rect 1886 844 1897 878
rect 1931 844 1942 878
rect 1886 810 1942 844
rect 1886 776 1897 810
rect 1931 776 1942 810
rect 1886 742 1942 776
rect 1886 708 1897 742
rect 1931 708 1942 742
rect 1886 674 1942 708
rect 1886 640 1897 674
rect 1931 640 1942 674
rect 1886 606 1942 640
rect 1886 572 1897 606
rect 1931 572 1942 606
rect 1886 538 1942 572
rect 1886 504 1897 538
rect 1931 504 1942 538
rect 1886 470 1942 504
rect 1886 436 1897 470
rect 1931 436 1942 470
rect 1886 402 1942 436
rect 1886 368 1897 402
rect 1931 368 1942 402
rect 1886 334 1942 368
rect 1886 300 1897 334
rect 1931 300 1942 334
rect 1886 266 1942 300
rect 1886 232 1897 266
rect 1931 232 1942 266
rect 1886 198 1942 232
rect 1886 164 1897 198
rect 1931 164 1942 198
rect 1886 152 1942 164
rect 2108 1150 2164 1162
rect 2108 1116 2119 1150
rect 2153 1116 2164 1150
rect 2108 1082 2164 1116
rect 2108 1048 2119 1082
rect 2153 1048 2164 1082
rect 2108 1014 2164 1048
rect 2108 980 2119 1014
rect 2153 980 2164 1014
rect 2108 946 2164 980
rect 2108 912 2119 946
rect 2153 912 2164 946
rect 2108 878 2164 912
rect 2108 844 2119 878
rect 2153 844 2164 878
rect 2108 810 2164 844
rect 2108 776 2119 810
rect 2153 776 2164 810
rect 2108 742 2164 776
rect 2108 708 2119 742
rect 2153 708 2164 742
rect 2108 674 2164 708
rect 2108 640 2119 674
rect 2153 640 2164 674
rect 2108 606 2164 640
rect 2108 572 2119 606
rect 2153 572 2164 606
rect 2108 538 2164 572
rect 2108 504 2119 538
rect 2153 504 2164 538
rect 2108 470 2164 504
rect 2108 436 2119 470
rect 2153 436 2164 470
rect 2108 402 2164 436
rect 2108 368 2119 402
rect 2153 368 2164 402
rect 2108 334 2164 368
rect 2108 300 2119 334
rect 2153 300 2164 334
rect 2108 266 2164 300
rect 2108 232 2119 266
rect 2153 232 2164 266
rect 2108 198 2164 232
rect 2108 164 2119 198
rect 2153 164 2164 198
rect 2108 152 2164 164
rect 2194 1150 2250 1162
rect 2194 1116 2205 1150
rect 2239 1116 2250 1150
rect 2194 1082 2250 1116
rect 2194 1048 2205 1082
rect 2239 1048 2250 1082
rect 2194 1014 2250 1048
rect 2194 980 2205 1014
rect 2239 980 2250 1014
rect 2194 946 2250 980
rect 2194 912 2205 946
rect 2239 912 2250 946
rect 2194 878 2250 912
rect 2194 844 2205 878
rect 2239 844 2250 878
rect 2194 810 2250 844
rect 2194 776 2205 810
rect 2239 776 2250 810
rect 2194 742 2250 776
rect 2194 708 2205 742
rect 2239 708 2250 742
rect 2194 674 2250 708
rect 2194 640 2205 674
rect 2239 640 2250 674
rect 2194 606 2250 640
rect 2194 572 2205 606
rect 2239 572 2250 606
rect 2194 538 2250 572
rect 2194 504 2205 538
rect 2239 504 2250 538
rect 2194 470 2250 504
rect 2194 436 2205 470
rect 2239 436 2250 470
rect 2194 402 2250 436
rect 2194 368 2205 402
rect 2239 368 2250 402
rect 2194 334 2250 368
rect 2194 300 2205 334
rect 2239 300 2250 334
rect 2194 266 2250 300
rect 2194 232 2205 266
rect 2239 232 2250 266
rect 2194 198 2250 232
rect 2194 164 2205 198
rect 2239 164 2250 198
rect 2194 152 2250 164
rect 2280 1150 2336 1162
rect 2280 1116 2291 1150
rect 2325 1116 2336 1150
rect 2280 1082 2336 1116
rect 2280 1048 2291 1082
rect 2325 1048 2336 1082
rect 2280 1014 2336 1048
rect 2280 980 2291 1014
rect 2325 980 2336 1014
rect 2280 946 2336 980
rect 2280 912 2291 946
rect 2325 912 2336 946
rect 2280 878 2336 912
rect 2280 844 2291 878
rect 2325 844 2336 878
rect 2280 810 2336 844
rect 2280 776 2291 810
rect 2325 776 2336 810
rect 2280 742 2336 776
rect 2280 708 2291 742
rect 2325 708 2336 742
rect 2280 674 2336 708
rect 2280 640 2291 674
rect 2325 640 2336 674
rect 2280 606 2336 640
rect 2280 572 2291 606
rect 2325 572 2336 606
rect 2280 538 2336 572
rect 2280 504 2291 538
rect 2325 504 2336 538
rect 2280 470 2336 504
rect 2280 436 2291 470
rect 2325 436 2336 470
rect 2280 402 2336 436
rect 2280 368 2291 402
rect 2325 368 2336 402
rect 2280 334 2336 368
rect 2280 300 2291 334
rect 2325 300 2336 334
rect 2280 266 2336 300
rect 2280 232 2291 266
rect 2325 232 2336 266
rect 2280 198 2336 232
rect 2280 164 2291 198
rect 2325 164 2336 198
rect 2280 152 2336 164
<< ndiffc >>
rect 149 1116 183 1150
rect 149 1048 183 1082
rect 149 980 183 1014
rect 149 912 183 946
rect 149 844 183 878
rect 149 776 183 810
rect 149 708 183 742
rect 149 640 183 674
rect 149 572 183 606
rect 149 504 183 538
rect 149 436 183 470
rect 149 368 183 402
rect 149 300 183 334
rect 149 232 183 266
rect 149 164 183 198
rect 235 1116 269 1150
rect 235 1048 269 1082
rect 235 980 269 1014
rect 235 912 269 946
rect 235 844 269 878
rect 235 776 269 810
rect 235 708 269 742
rect 235 640 269 674
rect 235 572 269 606
rect 235 504 269 538
rect 235 436 269 470
rect 235 368 269 402
rect 235 300 269 334
rect 235 232 269 266
rect 235 164 269 198
rect 321 1116 355 1150
rect 321 1048 355 1082
rect 321 980 355 1014
rect 321 912 355 946
rect 321 844 355 878
rect 321 776 355 810
rect 321 708 355 742
rect 321 640 355 674
rect 321 572 355 606
rect 321 504 355 538
rect 321 436 355 470
rect 321 368 355 402
rect 321 300 355 334
rect 321 232 355 266
rect 321 164 355 198
rect 543 1116 577 1150
rect 543 1048 577 1082
rect 543 980 577 1014
rect 543 912 577 946
rect 543 844 577 878
rect 543 776 577 810
rect 543 708 577 742
rect 543 640 577 674
rect 543 572 577 606
rect 543 504 577 538
rect 543 436 577 470
rect 543 368 577 402
rect 543 300 577 334
rect 543 232 577 266
rect 543 164 577 198
rect 629 1116 663 1150
rect 629 1048 663 1082
rect 629 980 663 1014
rect 629 912 663 946
rect 629 844 663 878
rect 629 776 663 810
rect 629 708 663 742
rect 629 640 663 674
rect 629 572 663 606
rect 629 504 663 538
rect 629 436 663 470
rect 629 368 663 402
rect 629 300 663 334
rect 629 232 663 266
rect 629 164 663 198
rect 715 1116 749 1150
rect 715 1048 749 1082
rect 715 980 749 1014
rect 715 912 749 946
rect 715 844 749 878
rect 715 776 749 810
rect 715 708 749 742
rect 715 640 749 674
rect 715 572 749 606
rect 715 504 749 538
rect 715 436 749 470
rect 715 368 749 402
rect 715 300 749 334
rect 715 232 749 266
rect 715 164 749 198
rect 937 1116 971 1150
rect 937 1048 971 1082
rect 937 980 971 1014
rect 937 912 971 946
rect 937 844 971 878
rect 937 776 971 810
rect 937 708 971 742
rect 937 640 971 674
rect 937 572 971 606
rect 937 504 971 538
rect 937 436 971 470
rect 937 368 971 402
rect 937 300 971 334
rect 937 232 971 266
rect 937 164 971 198
rect 1023 1116 1057 1150
rect 1023 1048 1057 1082
rect 1023 980 1057 1014
rect 1023 912 1057 946
rect 1023 844 1057 878
rect 1023 776 1057 810
rect 1023 708 1057 742
rect 1023 640 1057 674
rect 1023 572 1057 606
rect 1023 504 1057 538
rect 1023 436 1057 470
rect 1023 368 1057 402
rect 1023 300 1057 334
rect 1023 232 1057 266
rect 1023 164 1057 198
rect 1109 1116 1143 1150
rect 1109 1048 1143 1082
rect 1109 980 1143 1014
rect 1109 912 1143 946
rect 1109 844 1143 878
rect 1109 776 1143 810
rect 1109 708 1143 742
rect 1109 640 1143 674
rect 1109 572 1143 606
rect 1109 504 1143 538
rect 1109 436 1143 470
rect 1109 368 1143 402
rect 1109 300 1143 334
rect 1109 232 1143 266
rect 1109 164 1143 198
rect 1331 1116 1365 1150
rect 1331 1048 1365 1082
rect 1331 980 1365 1014
rect 1331 912 1365 946
rect 1331 844 1365 878
rect 1331 776 1365 810
rect 1331 708 1365 742
rect 1331 640 1365 674
rect 1331 572 1365 606
rect 1331 504 1365 538
rect 1331 436 1365 470
rect 1331 368 1365 402
rect 1331 300 1365 334
rect 1331 232 1365 266
rect 1331 164 1365 198
rect 1417 1116 1451 1150
rect 1417 1048 1451 1082
rect 1417 980 1451 1014
rect 1417 912 1451 946
rect 1417 844 1451 878
rect 1417 776 1451 810
rect 1417 708 1451 742
rect 1417 640 1451 674
rect 1417 572 1451 606
rect 1417 504 1451 538
rect 1417 436 1451 470
rect 1417 368 1451 402
rect 1417 300 1451 334
rect 1417 232 1451 266
rect 1417 164 1451 198
rect 1503 1116 1537 1150
rect 1503 1048 1537 1082
rect 1503 980 1537 1014
rect 1503 912 1537 946
rect 1503 844 1537 878
rect 1503 776 1537 810
rect 1503 708 1537 742
rect 1503 640 1537 674
rect 1503 572 1537 606
rect 1503 504 1537 538
rect 1503 436 1537 470
rect 1503 368 1537 402
rect 1503 300 1537 334
rect 1503 232 1537 266
rect 1503 164 1537 198
rect 1725 1116 1759 1150
rect 1725 1048 1759 1082
rect 1725 980 1759 1014
rect 1725 912 1759 946
rect 1725 844 1759 878
rect 1725 776 1759 810
rect 1725 708 1759 742
rect 1725 640 1759 674
rect 1725 572 1759 606
rect 1725 504 1759 538
rect 1725 436 1759 470
rect 1725 368 1759 402
rect 1725 300 1759 334
rect 1725 232 1759 266
rect 1725 164 1759 198
rect 1811 1116 1845 1150
rect 1811 1048 1845 1082
rect 1811 980 1845 1014
rect 1811 912 1845 946
rect 1811 844 1845 878
rect 1811 776 1845 810
rect 1811 708 1845 742
rect 1811 640 1845 674
rect 1811 572 1845 606
rect 1811 504 1845 538
rect 1811 436 1845 470
rect 1811 368 1845 402
rect 1811 300 1845 334
rect 1811 232 1845 266
rect 1811 164 1845 198
rect 1897 1116 1931 1150
rect 1897 1048 1931 1082
rect 1897 980 1931 1014
rect 1897 912 1931 946
rect 1897 844 1931 878
rect 1897 776 1931 810
rect 1897 708 1931 742
rect 1897 640 1931 674
rect 1897 572 1931 606
rect 1897 504 1931 538
rect 1897 436 1931 470
rect 1897 368 1931 402
rect 1897 300 1931 334
rect 1897 232 1931 266
rect 1897 164 1931 198
rect 2119 1116 2153 1150
rect 2119 1048 2153 1082
rect 2119 980 2153 1014
rect 2119 912 2153 946
rect 2119 844 2153 878
rect 2119 776 2153 810
rect 2119 708 2153 742
rect 2119 640 2153 674
rect 2119 572 2153 606
rect 2119 504 2153 538
rect 2119 436 2153 470
rect 2119 368 2153 402
rect 2119 300 2153 334
rect 2119 232 2153 266
rect 2119 164 2153 198
rect 2205 1116 2239 1150
rect 2205 1048 2239 1082
rect 2205 980 2239 1014
rect 2205 912 2239 946
rect 2205 844 2239 878
rect 2205 776 2239 810
rect 2205 708 2239 742
rect 2205 640 2239 674
rect 2205 572 2239 606
rect 2205 504 2239 538
rect 2205 436 2239 470
rect 2205 368 2239 402
rect 2205 300 2239 334
rect 2205 232 2239 266
rect 2205 164 2239 198
rect 2291 1116 2325 1150
rect 2291 1048 2325 1082
rect 2291 980 2325 1014
rect 2291 912 2325 946
rect 2291 844 2325 878
rect 2291 776 2325 810
rect 2291 708 2325 742
rect 2291 640 2325 674
rect 2291 572 2325 606
rect 2291 504 2325 538
rect 2291 436 2325 470
rect 2291 368 2325 402
rect 2291 300 2325 334
rect 2291 232 2325 266
rect 2291 164 2325 198
<< psubdiff >>
rect 26 1116 84 1162
rect 26 1082 38 1116
rect 72 1082 84 1116
rect 26 1048 84 1082
rect 26 1014 38 1048
rect 72 1014 84 1048
rect 26 980 84 1014
rect 26 946 38 980
rect 72 946 84 980
rect 26 912 84 946
rect 26 878 38 912
rect 72 878 84 912
rect 26 844 84 878
rect 26 810 38 844
rect 72 810 84 844
rect 26 776 84 810
rect 26 742 38 776
rect 72 742 84 776
rect 26 708 84 742
rect 26 674 38 708
rect 72 674 84 708
rect 26 640 84 674
rect 26 606 38 640
rect 72 606 84 640
rect 26 572 84 606
rect 26 538 38 572
rect 72 538 84 572
rect 26 504 84 538
rect 26 470 38 504
rect 72 470 84 504
rect 26 436 84 470
rect 26 402 38 436
rect 72 402 84 436
rect 26 368 84 402
rect 26 334 38 368
rect 72 334 84 368
rect 26 300 84 334
rect 26 266 38 300
rect 72 266 84 300
rect 26 232 84 266
rect 26 198 38 232
rect 72 198 84 232
rect 26 152 84 198
rect 420 1116 478 1162
rect 420 1082 432 1116
rect 466 1082 478 1116
rect 420 1048 478 1082
rect 420 1014 432 1048
rect 466 1014 478 1048
rect 420 980 478 1014
rect 420 946 432 980
rect 466 946 478 980
rect 420 912 478 946
rect 420 878 432 912
rect 466 878 478 912
rect 420 844 478 878
rect 420 810 432 844
rect 466 810 478 844
rect 420 776 478 810
rect 420 742 432 776
rect 466 742 478 776
rect 420 708 478 742
rect 420 674 432 708
rect 466 674 478 708
rect 420 640 478 674
rect 420 606 432 640
rect 466 606 478 640
rect 420 572 478 606
rect 420 538 432 572
rect 466 538 478 572
rect 420 504 478 538
rect 420 470 432 504
rect 466 470 478 504
rect 420 436 478 470
rect 420 402 432 436
rect 466 402 478 436
rect 420 368 478 402
rect 420 334 432 368
rect 466 334 478 368
rect 420 300 478 334
rect 420 266 432 300
rect 466 266 478 300
rect 420 232 478 266
rect 420 198 432 232
rect 466 198 478 232
rect 420 152 478 198
rect 814 1116 872 1162
rect 814 1082 826 1116
rect 860 1082 872 1116
rect 814 1048 872 1082
rect 814 1014 826 1048
rect 860 1014 872 1048
rect 814 980 872 1014
rect 814 946 826 980
rect 860 946 872 980
rect 814 912 872 946
rect 814 878 826 912
rect 860 878 872 912
rect 814 844 872 878
rect 814 810 826 844
rect 860 810 872 844
rect 814 776 872 810
rect 814 742 826 776
rect 860 742 872 776
rect 814 708 872 742
rect 814 674 826 708
rect 860 674 872 708
rect 814 640 872 674
rect 814 606 826 640
rect 860 606 872 640
rect 814 572 872 606
rect 814 538 826 572
rect 860 538 872 572
rect 814 504 872 538
rect 814 470 826 504
rect 860 470 872 504
rect 814 436 872 470
rect 814 402 826 436
rect 860 402 872 436
rect 814 368 872 402
rect 814 334 826 368
rect 860 334 872 368
rect 814 300 872 334
rect 814 266 826 300
rect 860 266 872 300
rect 814 232 872 266
rect 814 198 826 232
rect 860 198 872 232
rect 814 152 872 198
rect 1208 1116 1266 1162
rect 1208 1082 1220 1116
rect 1254 1082 1266 1116
rect 1208 1048 1266 1082
rect 1208 1014 1220 1048
rect 1254 1014 1266 1048
rect 1208 980 1266 1014
rect 1208 946 1220 980
rect 1254 946 1266 980
rect 1208 912 1266 946
rect 1208 878 1220 912
rect 1254 878 1266 912
rect 1208 844 1266 878
rect 1208 810 1220 844
rect 1254 810 1266 844
rect 1208 776 1266 810
rect 1208 742 1220 776
rect 1254 742 1266 776
rect 1208 708 1266 742
rect 1208 674 1220 708
rect 1254 674 1266 708
rect 1208 640 1266 674
rect 1208 606 1220 640
rect 1254 606 1266 640
rect 1208 572 1266 606
rect 1208 538 1220 572
rect 1254 538 1266 572
rect 1208 504 1266 538
rect 1208 470 1220 504
rect 1254 470 1266 504
rect 1208 436 1266 470
rect 1208 402 1220 436
rect 1254 402 1266 436
rect 1208 368 1266 402
rect 1208 334 1220 368
rect 1254 334 1266 368
rect 1208 300 1266 334
rect 1208 266 1220 300
rect 1254 266 1266 300
rect 1208 232 1266 266
rect 1208 198 1220 232
rect 1254 198 1266 232
rect 1208 152 1266 198
rect 1602 1116 1660 1162
rect 1602 1082 1614 1116
rect 1648 1082 1660 1116
rect 1602 1048 1660 1082
rect 1602 1014 1614 1048
rect 1648 1014 1660 1048
rect 1602 980 1660 1014
rect 1602 946 1614 980
rect 1648 946 1660 980
rect 1602 912 1660 946
rect 1602 878 1614 912
rect 1648 878 1660 912
rect 1602 844 1660 878
rect 1602 810 1614 844
rect 1648 810 1660 844
rect 1602 776 1660 810
rect 1602 742 1614 776
rect 1648 742 1660 776
rect 1602 708 1660 742
rect 1602 674 1614 708
rect 1648 674 1660 708
rect 1602 640 1660 674
rect 1602 606 1614 640
rect 1648 606 1660 640
rect 1602 572 1660 606
rect 1602 538 1614 572
rect 1648 538 1660 572
rect 1602 504 1660 538
rect 1602 470 1614 504
rect 1648 470 1660 504
rect 1602 436 1660 470
rect 1602 402 1614 436
rect 1648 402 1660 436
rect 1602 368 1660 402
rect 1602 334 1614 368
rect 1648 334 1660 368
rect 1602 300 1660 334
rect 1602 266 1614 300
rect 1648 266 1660 300
rect 1602 232 1660 266
rect 1602 198 1614 232
rect 1648 198 1660 232
rect 1602 152 1660 198
rect 1996 1116 2054 1162
rect 1996 1082 2008 1116
rect 2042 1082 2054 1116
rect 1996 1048 2054 1082
rect 1996 1014 2008 1048
rect 2042 1014 2054 1048
rect 1996 980 2054 1014
rect 1996 946 2008 980
rect 2042 946 2054 980
rect 1996 912 2054 946
rect 1996 878 2008 912
rect 2042 878 2054 912
rect 1996 844 2054 878
rect 1996 810 2008 844
rect 2042 810 2054 844
rect 1996 776 2054 810
rect 1996 742 2008 776
rect 2042 742 2054 776
rect 1996 708 2054 742
rect 1996 674 2008 708
rect 2042 674 2054 708
rect 1996 640 2054 674
rect 1996 606 2008 640
rect 2042 606 2054 640
rect 1996 572 2054 606
rect 1996 538 2008 572
rect 2042 538 2054 572
rect 1996 504 2054 538
rect 1996 470 2008 504
rect 2042 470 2054 504
rect 1996 436 2054 470
rect 1996 402 2008 436
rect 2042 402 2054 436
rect 1996 368 2054 402
rect 1996 334 2008 368
rect 2042 334 2054 368
rect 1996 300 2054 334
rect 1996 266 2008 300
rect 2042 266 2054 300
rect 1996 232 2054 266
rect 1996 198 2008 232
rect 2042 198 2054 232
rect 1996 152 2054 198
rect 2390 1116 2448 1162
rect 2390 1082 2402 1116
rect 2436 1082 2448 1116
rect 2390 1048 2448 1082
rect 2390 1014 2402 1048
rect 2436 1014 2448 1048
rect 2390 980 2448 1014
rect 2390 946 2402 980
rect 2436 946 2448 980
rect 2390 912 2448 946
rect 2390 878 2402 912
rect 2436 878 2448 912
rect 2390 844 2448 878
rect 2390 810 2402 844
rect 2436 810 2448 844
rect 2390 776 2448 810
rect 2390 742 2402 776
rect 2436 742 2448 776
rect 2390 708 2448 742
rect 2390 674 2402 708
rect 2436 674 2448 708
rect 2390 640 2448 674
rect 2390 606 2402 640
rect 2436 606 2448 640
rect 2390 572 2448 606
rect 2390 538 2402 572
rect 2436 538 2448 572
rect 2390 504 2448 538
rect 2390 470 2402 504
rect 2436 470 2448 504
rect 2390 436 2448 470
rect 2390 402 2402 436
rect 2436 402 2448 436
rect 2390 368 2448 402
rect 2390 334 2402 368
rect 2436 334 2448 368
rect 2390 300 2448 334
rect 2390 266 2402 300
rect 2436 266 2448 300
rect 2390 232 2448 266
rect 2390 198 2402 232
rect 2436 198 2448 232
rect 2390 152 2448 198
<< psubdiffcont >>
rect 38 1082 72 1116
rect 38 1014 72 1048
rect 38 946 72 980
rect 38 878 72 912
rect 38 810 72 844
rect 38 742 72 776
rect 38 674 72 708
rect 38 606 72 640
rect 38 538 72 572
rect 38 470 72 504
rect 38 402 72 436
rect 38 334 72 368
rect 38 266 72 300
rect 38 198 72 232
rect 432 1082 466 1116
rect 432 1014 466 1048
rect 432 946 466 980
rect 432 878 466 912
rect 432 810 466 844
rect 432 742 466 776
rect 432 674 466 708
rect 432 606 466 640
rect 432 538 466 572
rect 432 470 466 504
rect 432 402 466 436
rect 432 334 466 368
rect 432 266 466 300
rect 432 198 466 232
rect 826 1082 860 1116
rect 826 1014 860 1048
rect 826 946 860 980
rect 826 878 860 912
rect 826 810 860 844
rect 826 742 860 776
rect 826 674 860 708
rect 826 606 860 640
rect 826 538 860 572
rect 826 470 860 504
rect 826 402 860 436
rect 826 334 860 368
rect 826 266 860 300
rect 826 198 860 232
rect 1220 1082 1254 1116
rect 1220 1014 1254 1048
rect 1220 946 1254 980
rect 1220 878 1254 912
rect 1220 810 1254 844
rect 1220 742 1254 776
rect 1220 674 1254 708
rect 1220 606 1254 640
rect 1220 538 1254 572
rect 1220 470 1254 504
rect 1220 402 1254 436
rect 1220 334 1254 368
rect 1220 266 1254 300
rect 1220 198 1254 232
rect 1614 1082 1648 1116
rect 1614 1014 1648 1048
rect 1614 946 1648 980
rect 1614 878 1648 912
rect 1614 810 1648 844
rect 1614 742 1648 776
rect 1614 674 1648 708
rect 1614 606 1648 640
rect 1614 538 1648 572
rect 1614 470 1648 504
rect 1614 402 1648 436
rect 1614 334 1648 368
rect 1614 266 1648 300
rect 1614 198 1648 232
rect 2008 1082 2042 1116
rect 2008 1014 2042 1048
rect 2008 946 2042 980
rect 2008 878 2042 912
rect 2008 810 2042 844
rect 2008 742 2042 776
rect 2008 674 2042 708
rect 2008 606 2042 640
rect 2008 538 2042 572
rect 2008 470 2042 504
rect 2008 402 2042 436
rect 2008 334 2042 368
rect 2008 266 2042 300
rect 2008 198 2042 232
rect 2402 1082 2436 1116
rect 2402 1014 2436 1048
rect 2402 946 2436 980
rect 2402 878 2436 912
rect 2402 810 2436 844
rect 2402 742 2436 776
rect 2402 674 2436 708
rect 2402 606 2436 640
rect 2402 538 2436 572
rect 2402 470 2436 504
rect 2402 402 2436 436
rect 2402 334 2436 368
rect 2402 266 2436 300
rect 2402 198 2436 232
<< poly >>
rect 151 1234 353 1254
rect 151 1200 167 1234
rect 201 1200 235 1234
rect 269 1200 303 1234
rect 337 1200 353 1234
rect 151 1184 353 1200
rect 545 1234 747 1254
rect 545 1200 561 1234
rect 595 1200 629 1234
rect 663 1200 697 1234
rect 731 1200 747 1234
rect 545 1184 747 1200
rect 939 1234 1141 1254
rect 939 1200 955 1234
rect 989 1200 1023 1234
rect 1057 1200 1091 1234
rect 1125 1200 1141 1234
rect 939 1184 1141 1200
rect 1333 1234 1535 1254
rect 1333 1200 1349 1234
rect 1383 1200 1417 1234
rect 1451 1200 1485 1234
rect 1519 1200 1535 1234
rect 1333 1184 1535 1200
rect 1727 1234 1929 1254
rect 1727 1200 1743 1234
rect 1777 1200 1811 1234
rect 1845 1200 1879 1234
rect 1913 1200 1929 1234
rect 1727 1184 1929 1200
rect 2121 1234 2323 1254
rect 2121 1200 2137 1234
rect 2171 1200 2205 1234
rect 2239 1200 2273 1234
rect 2307 1200 2323 1234
rect 2121 1184 2323 1200
rect 194 1162 224 1184
rect 280 1162 310 1184
rect 588 1162 618 1184
rect 674 1162 704 1184
rect 982 1162 1012 1184
rect 1068 1162 1098 1184
rect 1376 1162 1406 1184
rect 1462 1162 1492 1184
rect 1770 1162 1800 1184
rect 1856 1162 1886 1184
rect 2164 1162 2194 1184
rect 2250 1162 2280 1184
rect 194 130 224 152
rect 280 130 310 152
rect 588 130 618 152
rect 674 130 704 152
rect 982 130 1012 152
rect 1068 130 1098 152
rect 1376 130 1406 152
rect 1462 130 1492 152
rect 1770 130 1800 152
rect 1856 130 1886 152
rect 2164 130 2194 152
rect 2250 130 2280 152
rect 151 114 353 130
rect 151 80 167 114
rect 201 80 235 114
rect 269 80 303 114
rect 337 80 353 114
rect 151 60 353 80
rect 545 114 747 130
rect 545 80 561 114
rect 595 80 629 114
rect 663 80 697 114
rect 731 80 747 114
rect 545 60 747 80
rect 939 114 1141 130
rect 939 80 955 114
rect 989 80 1023 114
rect 1057 80 1091 114
rect 1125 80 1141 114
rect 939 60 1141 80
rect 1333 114 1535 130
rect 1333 80 1349 114
rect 1383 80 1417 114
rect 1451 80 1485 114
rect 1519 80 1535 114
rect 1333 60 1535 80
rect 1727 114 1929 130
rect 1727 80 1743 114
rect 1777 80 1811 114
rect 1845 80 1879 114
rect 1913 80 1929 114
rect 1727 60 1929 80
rect 2121 114 2323 130
rect 2121 80 2137 114
rect 2171 80 2205 114
rect 2239 80 2273 114
rect 2307 80 2323 114
rect 2121 60 2323 80
<< polycont >>
rect 167 1200 201 1234
rect 235 1200 269 1234
rect 303 1200 337 1234
rect 561 1200 595 1234
rect 629 1200 663 1234
rect 697 1200 731 1234
rect 955 1200 989 1234
rect 1023 1200 1057 1234
rect 1091 1200 1125 1234
rect 1349 1200 1383 1234
rect 1417 1200 1451 1234
rect 1485 1200 1519 1234
rect 1743 1200 1777 1234
rect 1811 1200 1845 1234
rect 1879 1200 1913 1234
rect 2137 1200 2171 1234
rect 2205 1200 2239 1234
rect 2273 1200 2307 1234
rect 167 80 201 114
rect 235 80 269 114
rect 303 80 337 114
rect 561 80 595 114
rect 629 80 663 114
rect 697 80 731 114
rect 955 80 989 114
rect 1023 80 1057 114
rect 1091 80 1125 114
rect 1349 80 1383 114
rect 1417 80 1451 114
rect 1485 80 1519 114
rect 1743 80 1777 114
rect 1811 80 1845 114
rect 1879 80 1913 114
rect 2137 80 2171 114
rect 2205 80 2239 114
rect 2273 80 2307 114
<< locali >>
rect 151 1200 163 1234
rect 201 1200 235 1234
rect 269 1200 303 1234
rect 341 1200 353 1234
rect 545 1200 557 1234
rect 595 1200 629 1234
rect 663 1200 697 1234
rect 735 1200 747 1234
rect 939 1200 951 1234
rect 989 1200 1023 1234
rect 1057 1200 1091 1234
rect 1129 1200 1141 1234
rect 1333 1200 1345 1234
rect 1383 1200 1417 1234
rect 1451 1200 1485 1234
rect 1523 1200 1535 1234
rect 1727 1200 1739 1234
rect 1777 1200 1811 1234
rect 1845 1200 1879 1234
rect 1917 1200 1929 1234
rect 2121 1200 2133 1234
rect 2171 1200 2205 1234
rect 2239 1200 2273 1234
rect 2311 1200 2323 1234
rect 149 1150 183 1166
rect 38 1070 72 1082
rect 38 998 72 1014
rect 38 926 72 946
rect 38 854 72 878
rect 38 782 72 810
rect 38 710 72 742
rect 38 640 72 674
rect 38 572 72 604
rect 38 504 72 532
rect 38 436 72 460
rect 38 368 72 388
rect 38 300 72 316
rect 38 232 72 244
rect 149 1082 183 1108
rect 149 1014 183 1036
rect 149 946 183 964
rect 149 878 183 892
rect 149 810 183 820
rect 149 742 183 748
rect 149 674 183 676
rect 149 638 183 640
rect 149 566 183 572
rect 149 494 183 504
rect 149 422 183 436
rect 149 350 183 368
rect 149 278 183 300
rect 149 206 183 232
rect 149 148 183 164
rect 235 1150 269 1166
rect 235 1082 269 1108
rect 235 1014 269 1036
rect 235 946 269 964
rect 235 878 269 892
rect 235 810 269 820
rect 235 742 269 748
rect 235 674 269 676
rect 235 638 269 640
rect 235 566 269 572
rect 235 494 269 504
rect 235 422 269 436
rect 235 350 269 368
rect 235 278 269 300
rect 235 206 269 232
rect 235 148 269 164
rect 321 1150 355 1166
rect 543 1150 577 1166
rect 321 1082 355 1108
rect 321 1014 355 1036
rect 321 946 355 964
rect 321 878 355 892
rect 321 810 355 820
rect 321 742 355 748
rect 321 674 355 676
rect 321 638 355 640
rect 321 566 355 572
rect 321 494 355 504
rect 321 422 355 436
rect 321 350 355 368
rect 321 278 355 300
rect 321 206 355 232
rect 432 1070 466 1082
rect 432 998 466 1014
rect 432 926 466 946
rect 432 854 466 878
rect 432 782 466 810
rect 432 710 466 742
rect 432 640 466 674
rect 432 572 466 604
rect 432 504 466 532
rect 432 436 466 460
rect 432 368 466 388
rect 432 300 466 316
rect 432 232 466 244
rect 543 1082 577 1108
rect 543 1014 577 1036
rect 543 946 577 964
rect 543 878 577 892
rect 543 810 577 820
rect 543 742 577 748
rect 543 674 577 676
rect 543 638 577 640
rect 543 566 577 572
rect 543 494 577 504
rect 543 422 577 436
rect 543 350 577 368
rect 543 278 577 300
rect 543 206 577 232
rect 321 148 355 164
rect 543 148 577 164
rect 629 1150 663 1166
rect 629 1082 663 1108
rect 629 1014 663 1036
rect 629 946 663 964
rect 629 878 663 892
rect 629 810 663 820
rect 629 742 663 748
rect 629 674 663 676
rect 629 638 663 640
rect 629 566 663 572
rect 629 494 663 504
rect 629 422 663 436
rect 629 350 663 368
rect 629 278 663 300
rect 629 206 663 232
rect 629 148 663 164
rect 715 1150 749 1166
rect 937 1150 971 1166
rect 715 1082 749 1108
rect 715 1014 749 1036
rect 715 946 749 964
rect 715 878 749 892
rect 715 810 749 820
rect 715 742 749 748
rect 715 674 749 676
rect 715 638 749 640
rect 715 566 749 572
rect 715 494 749 504
rect 715 422 749 436
rect 715 350 749 368
rect 715 278 749 300
rect 715 206 749 232
rect 826 1070 860 1082
rect 826 998 860 1014
rect 826 926 860 946
rect 826 854 860 878
rect 826 782 860 810
rect 826 710 860 742
rect 826 640 860 674
rect 826 572 860 604
rect 826 504 860 532
rect 826 436 860 460
rect 826 368 860 388
rect 826 300 860 316
rect 826 232 860 244
rect 937 1082 971 1108
rect 937 1014 971 1036
rect 937 946 971 964
rect 937 878 971 892
rect 937 810 971 820
rect 937 742 971 748
rect 937 674 971 676
rect 937 638 971 640
rect 937 566 971 572
rect 937 494 971 504
rect 937 422 971 436
rect 937 350 971 368
rect 937 278 971 300
rect 937 206 971 232
rect 715 148 749 164
rect 937 148 971 164
rect 1023 1150 1057 1166
rect 1023 1082 1057 1108
rect 1023 1014 1057 1036
rect 1023 946 1057 964
rect 1023 878 1057 892
rect 1023 810 1057 820
rect 1023 742 1057 748
rect 1023 674 1057 676
rect 1023 638 1057 640
rect 1023 566 1057 572
rect 1023 494 1057 504
rect 1023 422 1057 436
rect 1023 350 1057 368
rect 1023 278 1057 300
rect 1023 206 1057 232
rect 1023 148 1057 164
rect 1109 1150 1143 1166
rect 1331 1150 1365 1166
rect 1109 1082 1143 1108
rect 1109 1014 1143 1036
rect 1109 946 1143 964
rect 1109 878 1143 892
rect 1109 810 1143 820
rect 1109 742 1143 748
rect 1109 674 1143 676
rect 1109 638 1143 640
rect 1109 566 1143 572
rect 1109 494 1143 504
rect 1109 422 1143 436
rect 1109 350 1143 368
rect 1109 278 1143 300
rect 1109 206 1143 232
rect 1220 1070 1254 1082
rect 1220 998 1254 1014
rect 1220 926 1254 946
rect 1220 854 1254 878
rect 1220 782 1254 810
rect 1220 710 1254 742
rect 1220 640 1254 674
rect 1220 572 1254 604
rect 1220 504 1254 532
rect 1220 436 1254 460
rect 1220 368 1254 388
rect 1220 300 1254 316
rect 1220 232 1254 244
rect 1331 1082 1365 1108
rect 1331 1014 1365 1036
rect 1331 946 1365 964
rect 1331 878 1365 892
rect 1331 810 1365 820
rect 1331 742 1365 748
rect 1331 674 1365 676
rect 1331 638 1365 640
rect 1331 566 1365 572
rect 1331 494 1365 504
rect 1331 422 1365 436
rect 1331 350 1365 368
rect 1331 278 1365 300
rect 1331 206 1365 232
rect 1109 148 1143 164
rect 1331 148 1365 164
rect 1417 1150 1451 1166
rect 1417 1082 1451 1108
rect 1417 1014 1451 1036
rect 1417 946 1451 964
rect 1417 878 1451 892
rect 1417 810 1451 820
rect 1417 742 1451 748
rect 1417 674 1451 676
rect 1417 638 1451 640
rect 1417 566 1451 572
rect 1417 494 1451 504
rect 1417 422 1451 436
rect 1417 350 1451 368
rect 1417 278 1451 300
rect 1417 206 1451 232
rect 1417 148 1451 164
rect 1503 1150 1537 1166
rect 1725 1150 1759 1166
rect 1503 1082 1537 1108
rect 1503 1014 1537 1036
rect 1503 946 1537 964
rect 1503 878 1537 892
rect 1503 810 1537 820
rect 1503 742 1537 748
rect 1503 674 1537 676
rect 1503 638 1537 640
rect 1503 566 1537 572
rect 1503 494 1537 504
rect 1503 422 1537 436
rect 1503 350 1537 368
rect 1503 278 1537 300
rect 1503 206 1537 232
rect 1614 1070 1648 1082
rect 1614 998 1648 1014
rect 1614 926 1648 946
rect 1614 854 1648 878
rect 1614 782 1648 810
rect 1614 710 1648 742
rect 1614 640 1648 674
rect 1614 572 1648 604
rect 1614 504 1648 532
rect 1614 436 1648 460
rect 1614 368 1648 388
rect 1614 300 1648 316
rect 1614 232 1648 244
rect 1725 1082 1759 1108
rect 1725 1014 1759 1036
rect 1725 946 1759 964
rect 1725 878 1759 892
rect 1725 810 1759 820
rect 1725 742 1759 748
rect 1725 674 1759 676
rect 1725 638 1759 640
rect 1725 566 1759 572
rect 1725 494 1759 504
rect 1725 422 1759 436
rect 1725 350 1759 368
rect 1725 278 1759 300
rect 1725 206 1759 232
rect 1503 148 1537 164
rect 1725 148 1759 164
rect 1811 1150 1845 1166
rect 1811 1082 1845 1108
rect 1811 1014 1845 1036
rect 1811 946 1845 964
rect 1811 878 1845 892
rect 1811 810 1845 820
rect 1811 742 1845 748
rect 1811 674 1845 676
rect 1811 638 1845 640
rect 1811 566 1845 572
rect 1811 494 1845 504
rect 1811 422 1845 436
rect 1811 350 1845 368
rect 1811 278 1845 300
rect 1811 206 1845 232
rect 1811 148 1845 164
rect 1897 1150 1931 1166
rect 2119 1150 2153 1166
rect 1897 1082 1931 1108
rect 1897 1014 1931 1036
rect 1897 946 1931 964
rect 1897 878 1931 892
rect 1897 810 1931 820
rect 1897 742 1931 748
rect 1897 674 1931 676
rect 1897 638 1931 640
rect 1897 566 1931 572
rect 1897 494 1931 504
rect 1897 422 1931 436
rect 1897 350 1931 368
rect 1897 278 1931 300
rect 1897 206 1931 232
rect 2008 1070 2042 1082
rect 2008 998 2042 1014
rect 2008 926 2042 946
rect 2008 854 2042 878
rect 2008 782 2042 810
rect 2008 710 2042 742
rect 2008 640 2042 674
rect 2008 572 2042 604
rect 2008 504 2042 532
rect 2008 436 2042 460
rect 2008 368 2042 388
rect 2008 300 2042 316
rect 2008 232 2042 244
rect 2119 1082 2153 1108
rect 2119 1014 2153 1036
rect 2119 946 2153 964
rect 2119 878 2153 892
rect 2119 810 2153 820
rect 2119 742 2153 748
rect 2119 674 2153 676
rect 2119 638 2153 640
rect 2119 566 2153 572
rect 2119 494 2153 504
rect 2119 422 2153 436
rect 2119 350 2153 368
rect 2119 278 2153 300
rect 2119 206 2153 232
rect 1897 148 1931 164
rect 2119 148 2153 164
rect 2205 1150 2239 1166
rect 2205 1082 2239 1108
rect 2205 1014 2239 1036
rect 2205 946 2239 964
rect 2205 878 2239 892
rect 2205 810 2239 820
rect 2205 742 2239 748
rect 2205 674 2239 676
rect 2205 638 2239 640
rect 2205 566 2239 572
rect 2205 494 2239 504
rect 2205 422 2239 436
rect 2205 350 2239 368
rect 2205 278 2239 300
rect 2205 206 2239 232
rect 2205 148 2239 164
rect 2291 1150 2325 1166
rect 2291 1082 2325 1108
rect 2291 1014 2325 1036
rect 2291 946 2325 964
rect 2291 878 2325 892
rect 2291 810 2325 820
rect 2291 742 2325 748
rect 2291 674 2325 676
rect 2291 638 2325 640
rect 2291 566 2325 572
rect 2291 494 2325 504
rect 2291 422 2325 436
rect 2291 350 2325 368
rect 2291 278 2325 300
rect 2291 206 2325 232
rect 2402 1070 2436 1082
rect 2402 998 2436 1014
rect 2402 926 2436 946
rect 2402 854 2436 878
rect 2402 782 2436 810
rect 2402 710 2436 742
rect 2402 640 2436 674
rect 2402 572 2436 604
rect 2402 504 2436 532
rect 2402 436 2436 460
rect 2402 368 2436 388
rect 2402 300 2436 316
rect 2402 232 2436 244
rect 2291 148 2325 164
rect 151 80 163 114
rect 201 80 235 114
rect 269 80 303 114
rect 341 80 353 114
rect 545 80 557 114
rect 595 80 629 114
rect 663 80 697 114
rect 735 80 747 114
rect 939 80 951 114
rect 989 80 1023 114
rect 1057 80 1091 114
rect 1129 80 1141 114
rect 1333 80 1345 114
rect 1383 80 1417 114
rect 1451 80 1485 114
rect 1523 80 1535 114
rect 1727 80 1739 114
rect 1777 80 1811 114
rect 1845 80 1879 114
rect 1917 80 1929 114
rect 2121 80 2133 114
rect 2171 80 2205 114
rect 2239 80 2273 114
rect 2311 80 2323 114
<< viali >>
rect 163 1200 167 1234
rect 167 1200 197 1234
rect 235 1200 269 1234
rect 307 1200 337 1234
rect 337 1200 341 1234
rect 557 1200 561 1234
rect 561 1200 591 1234
rect 629 1200 663 1234
rect 701 1200 731 1234
rect 731 1200 735 1234
rect 951 1200 955 1234
rect 955 1200 985 1234
rect 1023 1200 1057 1234
rect 1095 1200 1125 1234
rect 1125 1200 1129 1234
rect 1345 1200 1349 1234
rect 1349 1200 1379 1234
rect 1417 1200 1451 1234
rect 1489 1200 1519 1234
rect 1519 1200 1523 1234
rect 1739 1200 1743 1234
rect 1743 1200 1773 1234
rect 1811 1200 1845 1234
rect 1883 1200 1913 1234
rect 1913 1200 1917 1234
rect 2133 1200 2137 1234
rect 2137 1200 2167 1234
rect 2205 1200 2239 1234
rect 2277 1200 2307 1234
rect 2307 1200 2311 1234
rect 38 1116 72 1142
rect 38 1108 72 1116
rect 38 1048 72 1070
rect 38 1036 72 1048
rect 38 980 72 998
rect 38 964 72 980
rect 38 912 72 926
rect 38 892 72 912
rect 38 844 72 854
rect 38 820 72 844
rect 38 776 72 782
rect 38 748 72 776
rect 38 708 72 710
rect 38 676 72 708
rect 38 606 72 638
rect 38 604 72 606
rect 38 538 72 566
rect 38 532 72 538
rect 38 470 72 494
rect 38 460 72 470
rect 38 402 72 422
rect 38 388 72 402
rect 38 334 72 350
rect 38 316 72 334
rect 38 266 72 278
rect 38 244 72 266
rect 38 198 72 206
rect 38 172 72 198
rect 149 1116 183 1142
rect 149 1108 183 1116
rect 149 1048 183 1070
rect 149 1036 183 1048
rect 149 980 183 998
rect 149 964 183 980
rect 149 912 183 926
rect 149 892 183 912
rect 149 844 183 854
rect 149 820 183 844
rect 149 776 183 782
rect 149 748 183 776
rect 149 708 183 710
rect 149 676 183 708
rect 149 606 183 638
rect 149 604 183 606
rect 149 538 183 566
rect 149 532 183 538
rect 149 470 183 494
rect 149 460 183 470
rect 149 402 183 422
rect 149 388 183 402
rect 149 334 183 350
rect 149 316 183 334
rect 149 266 183 278
rect 149 244 183 266
rect 149 198 183 206
rect 149 172 183 198
rect 235 1116 269 1142
rect 235 1108 269 1116
rect 235 1048 269 1070
rect 235 1036 269 1048
rect 235 980 269 998
rect 235 964 269 980
rect 235 912 269 926
rect 235 892 269 912
rect 235 844 269 854
rect 235 820 269 844
rect 235 776 269 782
rect 235 748 269 776
rect 235 708 269 710
rect 235 676 269 708
rect 235 606 269 638
rect 235 604 269 606
rect 235 538 269 566
rect 235 532 269 538
rect 235 470 269 494
rect 235 460 269 470
rect 235 402 269 422
rect 235 388 269 402
rect 235 334 269 350
rect 235 316 269 334
rect 235 266 269 278
rect 235 244 269 266
rect 235 198 269 206
rect 235 172 269 198
rect 321 1116 355 1142
rect 321 1108 355 1116
rect 321 1048 355 1070
rect 321 1036 355 1048
rect 321 980 355 998
rect 321 964 355 980
rect 321 912 355 926
rect 321 892 355 912
rect 321 844 355 854
rect 321 820 355 844
rect 321 776 355 782
rect 321 748 355 776
rect 321 708 355 710
rect 321 676 355 708
rect 321 606 355 638
rect 321 604 355 606
rect 321 538 355 566
rect 321 532 355 538
rect 321 470 355 494
rect 321 460 355 470
rect 321 402 355 422
rect 321 388 355 402
rect 321 334 355 350
rect 321 316 355 334
rect 321 266 355 278
rect 321 244 355 266
rect 321 198 355 206
rect 321 172 355 198
rect 432 1116 466 1142
rect 432 1108 466 1116
rect 432 1048 466 1070
rect 432 1036 466 1048
rect 432 980 466 998
rect 432 964 466 980
rect 432 912 466 926
rect 432 892 466 912
rect 432 844 466 854
rect 432 820 466 844
rect 432 776 466 782
rect 432 748 466 776
rect 432 708 466 710
rect 432 676 466 708
rect 432 606 466 638
rect 432 604 466 606
rect 432 538 466 566
rect 432 532 466 538
rect 432 470 466 494
rect 432 460 466 470
rect 432 402 466 422
rect 432 388 466 402
rect 432 334 466 350
rect 432 316 466 334
rect 432 266 466 278
rect 432 244 466 266
rect 432 198 466 206
rect 432 172 466 198
rect 543 1116 577 1142
rect 543 1108 577 1116
rect 543 1048 577 1070
rect 543 1036 577 1048
rect 543 980 577 998
rect 543 964 577 980
rect 543 912 577 926
rect 543 892 577 912
rect 543 844 577 854
rect 543 820 577 844
rect 543 776 577 782
rect 543 748 577 776
rect 543 708 577 710
rect 543 676 577 708
rect 543 606 577 638
rect 543 604 577 606
rect 543 538 577 566
rect 543 532 577 538
rect 543 470 577 494
rect 543 460 577 470
rect 543 402 577 422
rect 543 388 577 402
rect 543 334 577 350
rect 543 316 577 334
rect 543 266 577 278
rect 543 244 577 266
rect 543 198 577 206
rect 543 172 577 198
rect 629 1116 663 1142
rect 629 1108 663 1116
rect 629 1048 663 1070
rect 629 1036 663 1048
rect 629 980 663 998
rect 629 964 663 980
rect 629 912 663 926
rect 629 892 663 912
rect 629 844 663 854
rect 629 820 663 844
rect 629 776 663 782
rect 629 748 663 776
rect 629 708 663 710
rect 629 676 663 708
rect 629 606 663 638
rect 629 604 663 606
rect 629 538 663 566
rect 629 532 663 538
rect 629 470 663 494
rect 629 460 663 470
rect 629 402 663 422
rect 629 388 663 402
rect 629 334 663 350
rect 629 316 663 334
rect 629 266 663 278
rect 629 244 663 266
rect 629 198 663 206
rect 629 172 663 198
rect 715 1116 749 1142
rect 715 1108 749 1116
rect 715 1048 749 1070
rect 715 1036 749 1048
rect 715 980 749 998
rect 715 964 749 980
rect 715 912 749 926
rect 715 892 749 912
rect 715 844 749 854
rect 715 820 749 844
rect 715 776 749 782
rect 715 748 749 776
rect 715 708 749 710
rect 715 676 749 708
rect 715 606 749 638
rect 715 604 749 606
rect 715 538 749 566
rect 715 532 749 538
rect 715 470 749 494
rect 715 460 749 470
rect 715 402 749 422
rect 715 388 749 402
rect 715 334 749 350
rect 715 316 749 334
rect 715 266 749 278
rect 715 244 749 266
rect 715 198 749 206
rect 715 172 749 198
rect 826 1116 860 1142
rect 826 1108 860 1116
rect 826 1048 860 1070
rect 826 1036 860 1048
rect 826 980 860 998
rect 826 964 860 980
rect 826 912 860 926
rect 826 892 860 912
rect 826 844 860 854
rect 826 820 860 844
rect 826 776 860 782
rect 826 748 860 776
rect 826 708 860 710
rect 826 676 860 708
rect 826 606 860 638
rect 826 604 860 606
rect 826 538 860 566
rect 826 532 860 538
rect 826 470 860 494
rect 826 460 860 470
rect 826 402 860 422
rect 826 388 860 402
rect 826 334 860 350
rect 826 316 860 334
rect 826 266 860 278
rect 826 244 860 266
rect 826 198 860 206
rect 826 172 860 198
rect 937 1116 971 1142
rect 937 1108 971 1116
rect 937 1048 971 1070
rect 937 1036 971 1048
rect 937 980 971 998
rect 937 964 971 980
rect 937 912 971 926
rect 937 892 971 912
rect 937 844 971 854
rect 937 820 971 844
rect 937 776 971 782
rect 937 748 971 776
rect 937 708 971 710
rect 937 676 971 708
rect 937 606 971 638
rect 937 604 971 606
rect 937 538 971 566
rect 937 532 971 538
rect 937 470 971 494
rect 937 460 971 470
rect 937 402 971 422
rect 937 388 971 402
rect 937 334 971 350
rect 937 316 971 334
rect 937 266 971 278
rect 937 244 971 266
rect 937 198 971 206
rect 937 172 971 198
rect 1023 1116 1057 1142
rect 1023 1108 1057 1116
rect 1023 1048 1057 1070
rect 1023 1036 1057 1048
rect 1023 980 1057 998
rect 1023 964 1057 980
rect 1023 912 1057 926
rect 1023 892 1057 912
rect 1023 844 1057 854
rect 1023 820 1057 844
rect 1023 776 1057 782
rect 1023 748 1057 776
rect 1023 708 1057 710
rect 1023 676 1057 708
rect 1023 606 1057 638
rect 1023 604 1057 606
rect 1023 538 1057 566
rect 1023 532 1057 538
rect 1023 470 1057 494
rect 1023 460 1057 470
rect 1023 402 1057 422
rect 1023 388 1057 402
rect 1023 334 1057 350
rect 1023 316 1057 334
rect 1023 266 1057 278
rect 1023 244 1057 266
rect 1023 198 1057 206
rect 1023 172 1057 198
rect 1109 1116 1143 1142
rect 1109 1108 1143 1116
rect 1109 1048 1143 1070
rect 1109 1036 1143 1048
rect 1109 980 1143 998
rect 1109 964 1143 980
rect 1109 912 1143 926
rect 1109 892 1143 912
rect 1109 844 1143 854
rect 1109 820 1143 844
rect 1109 776 1143 782
rect 1109 748 1143 776
rect 1109 708 1143 710
rect 1109 676 1143 708
rect 1109 606 1143 638
rect 1109 604 1143 606
rect 1109 538 1143 566
rect 1109 532 1143 538
rect 1109 470 1143 494
rect 1109 460 1143 470
rect 1109 402 1143 422
rect 1109 388 1143 402
rect 1109 334 1143 350
rect 1109 316 1143 334
rect 1109 266 1143 278
rect 1109 244 1143 266
rect 1109 198 1143 206
rect 1109 172 1143 198
rect 1220 1116 1254 1142
rect 1220 1108 1254 1116
rect 1220 1048 1254 1070
rect 1220 1036 1254 1048
rect 1220 980 1254 998
rect 1220 964 1254 980
rect 1220 912 1254 926
rect 1220 892 1254 912
rect 1220 844 1254 854
rect 1220 820 1254 844
rect 1220 776 1254 782
rect 1220 748 1254 776
rect 1220 708 1254 710
rect 1220 676 1254 708
rect 1220 606 1254 638
rect 1220 604 1254 606
rect 1220 538 1254 566
rect 1220 532 1254 538
rect 1220 470 1254 494
rect 1220 460 1254 470
rect 1220 402 1254 422
rect 1220 388 1254 402
rect 1220 334 1254 350
rect 1220 316 1254 334
rect 1220 266 1254 278
rect 1220 244 1254 266
rect 1220 198 1254 206
rect 1220 172 1254 198
rect 1331 1116 1365 1142
rect 1331 1108 1365 1116
rect 1331 1048 1365 1070
rect 1331 1036 1365 1048
rect 1331 980 1365 998
rect 1331 964 1365 980
rect 1331 912 1365 926
rect 1331 892 1365 912
rect 1331 844 1365 854
rect 1331 820 1365 844
rect 1331 776 1365 782
rect 1331 748 1365 776
rect 1331 708 1365 710
rect 1331 676 1365 708
rect 1331 606 1365 638
rect 1331 604 1365 606
rect 1331 538 1365 566
rect 1331 532 1365 538
rect 1331 470 1365 494
rect 1331 460 1365 470
rect 1331 402 1365 422
rect 1331 388 1365 402
rect 1331 334 1365 350
rect 1331 316 1365 334
rect 1331 266 1365 278
rect 1331 244 1365 266
rect 1331 198 1365 206
rect 1331 172 1365 198
rect 1417 1116 1451 1142
rect 1417 1108 1451 1116
rect 1417 1048 1451 1070
rect 1417 1036 1451 1048
rect 1417 980 1451 998
rect 1417 964 1451 980
rect 1417 912 1451 926
rect 1417 892 1451 912
rect 1417 844 1451 854
rect 1417 820 1451 844
rect 1417 776 1451 782
rect 1417 748 1451 776
rect 1417 708 1451 710
rect 1417 676 1451 708
rect 1417 606 1451 638
rect 1417 604 1451 606
rect 1417 538 1451 566
rect 1417 532 1451 538
rect 1417 470 1451 494
rect 1417 460 1451 470
rect 1417 402 1451 422
rect 1417 388 1451 402
rect 1417 334 1451 350
rect 1417 316 1451 334
rect 1417 266 1451 278
rect 1417 244 1451 266
rect 1417 198 1451 206
rect 1417 172 1451 198
rect 1503 1116 1537 1142
rect 1503 1108 1537 1116
rect 1503 1048 1537 1070
rect 1503 1036 1537 1048
rect 1503 980 1537 998
rect 1503 964 1537 980
rect 1503 912 1537 926
rect 1503 892 1537 912
rect 1503 844 1537 854
rect 1503 820 1537 844
rect 1503 776 1537 782
rect 1503 748 1537 776
rect 1503 708 1537 710
rect 1503 676 1537 708
rect 1503 606 1537 638
rect 1503 604 1537 606
rect 1503 538 1537 566
rect 1503 532 1537 538
rect 1503 470 1537 494
rect 1503 460 1537 470
rect 1503 402 1537 422
rect 1503 388 1537 402
rect 1503 334 1537 350
rect 1503 316 1537 334
rect 1503 266 1537 278
rect 1503 244 1537 266
rect 1503 198 1537 206
rect 1503 172 1537 198
rect 1614 1116 1648 1142
rect 1614 1108 1648 1116
rect 1614 1048 1648 1070
rect 1614 1036 1648 1048
rect 1614 980 1648 998
rect 1614 964 1648 980
rect 1614 912 1648 926
rect 1614 892 1648 912
rect 1614 844 1648 854
rect 1614 820 1648 844
rect 1614 776 1648 782
rect 1614 748 1648 776
rect 1614 708 1648 710
rect 1614 676 1648 708
rect 1614 606 1648 638
rect 1614 604 1648 606
rect 1614 538 1648 566
rect 1614 532 1648 538
rect 1614 470 1648 494
rect 1614 460 1648 470
rect 1614 402 1648 422
rect 1614 388 1648 402
rect 1614 334 1648 350
rect 1614 316 1648 334
rect 1614 266 1648 278
rect 1614 244 1648 266
rect 1614 198 1648 206
rect 1614 172 1648 198
rect 1725 1116 1759 1142
rect 1725 1108 1759 1116
rect 1725 1048 1759 1070
rect 1725 1036 1759 1048
rect 1725 980 1759 998
rect 1725 964 1759 980
rect 1725 912 1759 926
rect 1725 892 1759 912
rect 1725 844 1759 854
rect 1725 820 1759 844
rect 1725 776 1759 782
rect 1725 748 1759 776
rect 1725 708 1759 710
rect 1725 676 1759 708
rect 1725 606 1759 638
rect 1725 604 1759 606
rect 1725 538 1759 566
rect 1725 532 1759 538
rect 1725 470 1759 494
rect 1725 460 1759 470
rect 1725 402 1759 422
rect 1725 388 1759 402
rect 1725 334 1759 350
rect 1725 316 1759 334
rect 1725 266 1759 278
rect 1725 244 1759 266
rect 1725 198 1759 206
rect 1725 172 1759 198
rect 1811 1116 1845 1142
rect 1811 1108 1845 1116
rect 1811 1048 1845 1070
rect 1811 1036 1845 1048
rect 1811 980 1845 998
rect 1811 964 1845 980
rect 1811 912 1845 926
rect 1811 892 1845 912
rect 1811 844 1845 854
rect 1811 820 1845 844
rect 1811 776 1845 782
rect 1811 748 1845 776
rect 1811 708 1845 710
rect 1811 676 1845 708
rect 1811 606 1845 638
rect 1811 604 1845 606
rect 1811 538 1845 566
rect 1811 532 1845 538
rect 1811 470 1845 494
rect 1811 460 1845 470
rect 1811 402 1845 422
rect 1811 388 1845 402
rect 1811 334 1845 350
rect 1811 316 1845 334
rect 1811 266 1845 278
rect 1811 244 1845 266
rect 1811 198 1845 206
rect 1811 172 1845 198
rect 1897 1116 1931 1142
rect 1897 1108 1931 1116
rect 1897 1048 1931 1070
rect 1897 1036 1931 1048
rect 1897 980 1931 998
rect 1897 964 1931 980
rect 1897 912 1931 926
rect 1897 892 1931 912
rect 1897 844 1931 854
rect 1897 820 1931 844
rect 1897 776 1931 782
rect 1897 748 1931 776
rect 1897 708 1931 710
rect 1897 676 1931 708
rect 1897 606 1931 638
rect 1897 604 1931 606
rect 1897 538 1931 566
rect 1897 532 1931 538
rect 1897 470 1931 494
rect 1897 460 1931 470
rect 1897 402 1931 422
rect 1897 388 1931 402
rect 1897 334 1931 350
rect 1897 316 1931 334
rect 1897 266 1931 278
rect 1897 244 1931 266
rect 1897 198 1931 206
rect 1897 172 1931 198
rect 2008 1116 2042 1142
rect 2008 1108 2042 1116
rect 2008 1048 2042 1070
rect 2008 1036 2042 1048
rect 2008 980 2042 998
rect 2008 964 2042 980
rect 2008 912 2042 926
rect 2008 892 2042 912
rect 2008 844 2042 854
rect 2008 820 2042 844
rect 2008 776 2042 782
rect 2008 748 2042 776
rect 2008 708 2042 710
rect 2008 676 2042 708
rect 2008 606 2042 638
rect 2008 604 2042 606
rect 2008 538 2042 566
rect 2008 532 2042 538
rect 2008 470 2042 494
rect 2008 460 2042 470
rect 2008 402 2042 422
rect 2008 388 2042 402
rect 2008 334 2042 350
rect 2008 316 2042 334
rect 2008 266 2042 278
rect 2008 244 2042 266
rect 2008 198 2042 206
rect 2008 172 2042 198
rect 2119 1116 2153 1142
rect 2119 1108 2153 1116
rect 2119 1048 2153 1070
rect 2119 1036 2153 1048
rect 2119 980 2153 998
rect 2119 964 2153 980
rect 2119 912 2153 926
rect 2119 892 2153 912
rect 2119 844 2153 854
rect 2119 820 2153 844
rect 2119 776 2153 782
rect 2119 748 2153 776
rect 2119 708 2153 710
rect 2119 676 2153 708
rect 2119 606 2153 638
rect 2119 604 2153 606
rect 2119 538 2153 566
rect 2119 532 2153 538
rect 2119 470 2153 494
rect 2119 460 2153 470
rect 2119 402 2153 422
rect 2119 388 2153 402
rect 2119 334 2153 350
rect 2119 316 2153 334
rect 2119 266 2153 278
rect 2119 244 2153 266
rect 2119 198 2153 206
rect 2119 172 2153 198
rect 2205 1116 2239 1142
rect 2205 1108 2239 1116
rect 2205 1048 2239 1070
rect 2205 1036 2239 1048
rect 2205 980 2239 998
rect 2205 964 2239 980
rect 2205 912 2239 926
rect 2205 892 2239 912
rect 2205 844 2239 854
rect 2205 820 2239 844
rect 2205 776 2239 782
rect 2205 748 2239 776
rect 2205 708 2239 710
rect 2205 676 2239 708
rect 2205 606 2239 638
rect 2205 604 2239 606
rect 2205 538 2239 566
rect 2205 532 2239 538
rect 2205 470 2239 494
rect 2205 460 2239 470
rect 2205 402 2239 422
rect 2205 388 2239 402
rect 2205 334 2239 350
rect 2205 316 2239 334
rect 2205 266 2239 278
rect 2205 244 2239 266
rect 2205 198 2239 206
rect 2205 172 2239 198
rect 2291 1116 2325 1142
rect 2291 1108 2325 1116
rect 2291 1048 2325 1070
rect 2291 1036 2325 1048
rect 2291 980 2325 998
rect 2291 964 2325 980
rect 2291 912 2325 926
rect 2291 892 2325 912
rect 2291 844 2325 854
rect 2291 820 2325 844
rect 2291 776 2325 782
rect 2291 748 2325 776
rect 2291 708 2325 710
rect 2291 676 2325 708
rect 2291 606 2325 638
rect 2291 604 2325 606
rect 2291 538 2325 566
rect 2291 532 2325 538
rect 2291 470 2325 494
rect 2291 460 2325 470
rect 2291 402 2325 422
rect 2291 388 2325 402
rect 2291 334 2325 350
rect 2291 316 2325 334
rect 2291 266 2325 278
rect 2291 244 2325 266
rect 2291 198 2325 206
rect 2291 172 2325 198
rect 2402 1116 2436 1142
rect 2402 1108 2436 1116
rect 2402 1048 2436 1070
rect 2402 1036 2436 1048
rect 2402 980 2436 998
rect 2402 964 2436 980
rect 2402 912 2436 926
rect 2402 892 2436 912
rect 2402 844 2436 854
rect 2402 820 2436 844
rect 2402 776 2436 782
rect 2402 748 2436 776
rect 2402 708 2436 710
rect 2402 676 2436 708
rect 2402 606 2436 638
rect 2402 604 2436 606
rect 2402 538 2436 566
rect 2402 532 2436 538
rect 2402 470 2436 494
rect 2402 460 2436 470
rect 2402 402 2436 422
rect 2402 388 2436 402
rect 2402 334 2436 350
rect 2402 316 2436 334
rect 2402 266 2436 278
rect 2402 244 2436 266
rect 2402 198 2436 206
rect 2402 172 2436 198
rect 163 80 167 114
rect 167 80 197 114
rect 235 80 269 114
rect 307 80 337 114
rect 337 80 341 114
rect 557 80 561 114
rect 561 80 591 114
rect 629 80 663 114
rect 701 80 731 114
rect 731 80 735 114
rect 951 80 955 114
rect 955 80 985 114
rect 1023 80 1057 114
rect 1095 80 1125 114
rect 1125 80 1129 114
rect 1345 80 1349 114
rect 1349 80 1379 114
rect 1417 80 1451 114
rect 1489 80 1519 114
rect 1519 80 1523 114
rect 1739 80 1743 114
rect 1743 80 1773 114
rect 1811 80 1845 114
rect 1883 80 1913 114
rect 1913 80 1917 114
rect 2133 80 2137 114
rect 2137 80 2167 114
rect 2205 80 2239 114
rect 2277 80 2307 114
rect 2307 80 2311 114
<< metal1 >>
rect 26 1370 2448 1440
rect 26 1142 84 1370
rect 140 1300 360 1320
rect 140 1220 160 1300
rect 240 1234 260 1300
rect 340 1234 360 1300
rect 140 1200 163 1220
rect 197 1200 235 1220
rect 269 1200 307 1220
rect 341 1200 360 1234
rect 151 1188 353 1200
rect 26 1108 38 1142
rect 72 1108 84 1142
rect 26 1070 84 1108
rect 26 1036 38 1070
rect 72 1036 84 1070
rect 26 998 84 1036
rect 26 964 38 998
rect 72 964 84 998
rect 26 926 84 964
rect 26 892 38 926
rect 72 892 84 926
rect 26 854 84 892
rect 26 820 38 854
rect 72 820 84 854
rect 26 782 84 820
rect 26 748 38 782
rect 72 748 84 782
rect 26 710 84 748
rect 26 676 38 710
rect 72 676 84 710
rect 26 638 84 676
rect 26 604 38 638
rect 72 604 84 638
rect 26 566 84 604
rect 26 532 38 566
rect 72 532 84 566
rect 26 494 84 532
rect 26 460 38 494
rect 72 460 84 494
rect 26 422 84 460
rect 26 388 38 422
rect 72 388 84 422
rect 26 350 84 388
rect 26 316 38 350
rect 72 316 84 350
rect 26 278 84 316
rect 26 244 38 278
rect 72 244 84 278
rect 26 206 84 244
rect 26 172 38 206
rect 72 172 84 206
rect 26 160 84 172
rect 140 1142 192 1154
rect 140 1108 149 1142
rect 183 1108 192 1142
rect 140 1070 192 1108
rect 140 1036 149 1070
rect 183 1036 192 1070
rect 140 998 192 1036
rect 140 964 149 998
rect 183 964 192 998
rect 140 926 192 964
rect 140 892 149 926
rect 183 892 192 926
rect 140 854 192 892
rect 140 820 149 854
rect 183 820 192 854
rect 140 782 192 820
rect 140 748 149 782
rect 183 748 192 782
rect 140 710 192 748
rect 140 676 149 710
rect 183 676 192 710
rect 140 638 192 676
rect 140 604 149 638
rect 183 604 192 638
rect 140 602 192 604
rect 140 538 149 550
rect 183 538 192 550
rect 140 474 149 486
rect 183 474 192 486
rect 140 410 149 422
rect 183 410 192 422
rect 140 350 192 358
rect 140 346 149 350
rect 183 346 192 350
rect 140 282 192 294
rect 140 218 192 230
rect 140 160 192 166
rect 226 1148 278 1154
rect 226 1084 278 1096
rect 226 1020 278 1032
rect 226 964 235 968
rect 269 964 278 968
rect 226 956 278 964
rect 226 892 235 904
rect 269 892 278 904
rect 226 828 235 840
rect 269 828 278 840
rect 226 764 235 776
rect 269 764 278 776
rect 226 710 278 712
rect 226 676 235 710
rect 269 676 278 710
rect 226 638 278 676
rect 226 604 235 638
rect 269 604 278 638
rect 226 566 278 604
rect 226 532 235 566
rect 269 532 278 566
rect 226 494 278 532
rect 226 460 235 494
rect 269 460 278 494
rect 226 422 278 460
rect 226 388 235 422
rect 269 388 278 422
rect 226 350 278 388
rect 226 316 235 350
rect 269 316 278 350
rect 226 278 278 316
rect 226 244 235 278
rect 269 244 278 278
rect 226 206 278 244
rect 226 172 235 206
rect 269 172 278 206
rect 226 160 278 172
rect 312 1142 364 1154
rect 312 1108 321 1142
rect 355 1108 364 1142
rect 312 1070 364 1108
rect 312 1036 321 1070
rect 355 1036 364 1070
rect 312 998 364 1036
rect 312 964 321 998
rect 355 964 364 998
rect 312 926 364 964
rect 312 892 321 926
rect 355 892 364 926
rect 312 854 364 892
rect 312 820 321 854
rect 355 820 364 854
rect 312 782 364 820
rect 312 748 321 782
rect 355 748 364 782
rect 312 710 364 748
rect 312 676 321 710
rect 355 676 364 710
rect 312 638 364 676
rect 312 604 321 638
rect 355 604 364 638
rect 312 602 364 604
rect 312 538 321 550
rect 355 538 364 550
rect 312 474 321 486
rect 355 474 364 486
rect 312 410 321 422
rect 355 410 364 422
rect 312 350 364 358
rect 312 346 321 350
rect 355 346 364 350
rect 312 282 364 294
rect 312 218 364 230
rect 312 160 364 166
rect 420 1142 478 1370
rect 530 1300 750 1320
rect 530 1220 550 1300
rect 630 1234 650 1300
rect 730 1234 750 1300
rect 530 1200 557 1220
rect 591 1200 629 1220
rect 663 1200 701 1220
rect 735 1200 750 1234
rect 541 1188 747 1200
rect 420 1108 432 1142
rect 466 1108 478 1142
rect 420 1070 478 1108
rect 420 1036 432 1070
rect 466 1036 478 1070
rect 420 998 478 1036
rect 420 964 432 998
rect 466 964 478 998
rect 420 926 478 964
rect 420 892 432 926
rect 466 892 478 926
rect 420 854 478 892
rect 420 820 432 854
rect 466 820 478 854
rect 420 782 478 820
rect 420 748 432 782
rect 466 748 478 782
rect 420 710 478 748
rect 420 676 432 710
rect 466 676 478 710
rect 420 638 478 676
rect 420 604 432 638
rect 466 604 478 638
rect 420 566 478 604
rect 420 532 432 566
rect 466 532 478 566
rect 420 494 478 532
rect 420 460 432 494
rect 466 460 478 494
rect 420 422 478 460
rect 420 388 432 422
rect 466 388 478 422
rect 420 350 478 388
rect 420 316 432 350
rect 466 316 478 350
rect 420 278 478 316
rect 420 244 432 278
rect 466 244 478 278
rect 420 206 478 244
rect 420 172 432 206
rect 466 172 478 206
rect 420 160 478 172
rect 534 1142 586 1154
rect 534 1108 543 1142
rect 577 1108 586 1142
rect 534 1070 586 1108
rect 534 1036 543 1070
rect 577 1036 586 1070
rect 534 998 586 1036
rect 534 964 543 998
rect 577 964 586 998
rect 534 926 586 964
rect 534 892 543 926
rect 577 892 586 926
rect 534 854 586 892
rect 534 820 543 854
rect 577 820 586 854
rect 534 782 586 820
rect 534 748 543 782
rect 577 748 586 782
rect 534 710 586 748
rect 534 676 543 710
rect 577 676 586 710
rect 534 638 586 676
rect 534 604 543 638
rect 577 604 586 638
rect 534 602 586 604
rect 534 538 543 550
rect 577 538 586 550
rect 534 474 543 486
rect 577 474 586 486
rect 534 410 543 422
rect 577 410 586 422
rect 534 350 586 358
rect 534 346 543 350
rect 577 346 586 350
rect 534 282 586 294
rect 534 218 586 230
rect 534 160 586 166
rect 620 1148 672 1154
rect 620 1084 672 1096
rect 620 1020 672 1032
rect 620 964 629 968
rect 663 964 672 968
rect 620 956 672 964
rect 620 892 629 904
rect 663 892 672 904
rect 620 828 629 840
rect 663 828 672 840
rect 620 764 629 776
rect 663 764 672 776
rect 620 710 672 712
rect 620 676 629 710
rect 663 676 672 710
rect 620 638 672 676
rect 620 604 629 638
rect 663 604 672 638
rect 620 566 672 604
rect 620 532 629 566
rect 663 532 672 566
rect 620 494 672 532
rect 620 460 629 494
rect 663 460 672 494
rect 620 422 672 460
rect 620 388 629 422
rect 663 388 672 422
rect 620 350 672 388
rect 620 316 629 350
rect 663 316 672 350
rect 620 278 672 316
rect 620 244 629 278
rect 663 244 672 278
rect 620 206 672 244
rect 620 172 629 206
rect 663 172 672 206
rect 620 160 672 172
rect 706 1142 758 1154
rect 706 1108 715 1142
rect 749 1108 758 1142
rect 706 1070 758 1108
rect 706 1036 715 1070
rect 749 1036 758 1070
rect 706 998 758 1036
rect 706 964 715 998
rect 749 964 758 998
rect 706 926 758 964
rect 706 892 715 926
rect 749 892 758 926
rect 706 854 758 892
rect 706 820 715 854
rect 749 820 758 854
rect 706 782 758 820
rect 706 748 715 782
rect 749 748 758 782
rect 706 710 758 748
rect 706 676 715 710
rect 749 676 758 710
rect 706 638 758 676
rect 706 604 715 638
rect 749 604 758 638
rect 706 602 758 604
rect 706 538 715 550
rect 749 538 758 550
rect 706 474 715 486
rect 749 474 758 486
rect 706 410 715 422
rect 749 410 758 422
rect 706 350 758 358
rect 706 346 715 350
rect 749 346 758 350
rect 706 282 758 294
rect 706 218 758 230
rect 706 160 758 166
rect 814 1142 872 1370
rect 930 1300 1150 1320
rect 930 1220 950 1300
rect 1030 1234 1050 1300
rect 1130 1220 1150 1300
rect 930 1200 951 1220
rect 985 1200 1023 1220
rect 1057 1200 1095 1220
rect 1129 1200 1150 1220
rect 939 1188 1143 1200
rect 814 1108 826 1142
rect 860 1108 872 1142
rect 814 1070 872 1108
rect 814 1036 826 1070
rect 860 1036 872 1070
rect 814 998 872 1036
rect 814 964 826 998
rect 860 964 872 998
rect 814 926 872 964
rect 814 892 826 926
rect 860 892 872 926
rect 814 854 872 892
rect 814 820 826 854
rect 860 820 872 854
rect 814 782 872 820
rect 814 748 826 782
rect 860 748 872 782
rect 814 710 872 748
rect 814 676 826 710
rect 860 676 872 710
rect 814 638 872 676
rect 814 604 826 638
rect 860 604 872 638
rect 814 566 872 604
rect 814 532 826 566
rect 860 532 872 566
rect 814 494 872 532
rect 814 460 826 494
rect 860 460 872 494
rect 814 422 872 460
rect 814 388 826 422
rect 860 388 872 422
rect 814 350 872 388
rect 814 316 826 350
rect 860 316 872 350
rect 814 278 872 316
rect 814 244 826 278
rect 860 244 872 278
rect 814 206 872 244
rect 814 172 826 206
rect 860 172 872 206
rect 814 160 872 172
rect 928 1142 980 1154
rect 928 1108 937 1142
rect 971 1108 980 1142
rect 928 1070 980 1108
rect 928 1036 937 1070
rect 971 1036 980 1070
rect 928 998 980 1036
rect 928 964 937 998
rect 971 964 980 998
rect 928 926 980 964
rect 928 892 937 926
rect 971 892 980 926
rect 928 854 980 892
rect 928 820 937 854
rect 971 820 980 854
rect 928 782 980 820
rect 928 748 937 782
rect 971 748 980 782
rect 928 710 980 748
rect 928 676 937 710
rect 971 676 980 710
rect 928 638 980 676
rect 928 604 937 638
rect 971 604 980 638
rect 928 602 980 604
rect 928 538 937 550
rect 971 538 980 550
rect 928 474 937 486
rect 971 474 980 486
rect 928 410 937 422
rect 971 410 980 422
rect 928 350 980 358
rect 928 346 937 350
rect 971 346 980 350
rect 928 282 980 294
rect 928 218 980 230
rect 928 160 980 166
rect 1014 1148 1066 1154
rect 1014 1084 1066 1096
rect 1014 1020 1066 1032
rect 1014 964 1023 968
rect 1057 964 1066 968
rect 1014 956 1066 964
rect 1014 892 1023 904
rect 1057 892 1066 904
rect 1014 828 1023 840
rect 1057 828 1066 840
rect 1014 764 1023 776
rect 1057 764 1066 776
rect 1014 710 1066 712
rect 1014 676 1023 710
rect 1057 676 1066 710
rect 1014 638 1066 676
rect 1014 604 1023 638
rect 1057 604 1066 638
rect 1014 566 1066 604
rect 1014 532 1023 566
rect 1057 532 1066 566
rect 1014 494 1066 532
rect 1014 460 1023 494
rect 1057 460 1066 494
rect 1014 422 1066 460
rect 1014 388 1023 422
rect 1057 388 1066 422
rect 1014 350 1066 388
rect 1014 316 1023 350
rect 1057 316 1066 350
rect 1014 278 1066 316
rect 1014 244 1023 278
rect 1057 244 1066 278
rect 1014 206 1066 244
rect 1014 172 1023 206
rect 1057 172 1066 206
rect 1014 160 1066 172
rect 1100 1142 1152 1154
rect 1100 1108 1109 1142
rect 1143 1108 1152 1142
rect 1100 1070 1152 1108
rect 1100 1036 1109 1070
rect 1143 1036 1152 1070
rect 1100 998 1152 1036
rect 1100 964 1109 998
rect 1143 964 1152 998
rect 1100 926 1152 964
rect 1100 892 1109 926
rect 1143 892 1152 926
rect 1100 854 1152 892
rect 1100 820 1109 854
rect 1143 820 1152 854
rect 1100 782 1152 820
rect 1100 748 1109 782
rect 1143 748 1152 782
rect 1100 710 1152 748
rect 1100 676 1109 710
rect 1143 676 1152 710
rect 1100 638 1152 676
rect 1100 604 1109 638
rect 1143 604 1152 638
rect 1100 602 1152 604
rect 1100 538 1109 550
rect 1143 538 1152 550
rect 1100 474 1109 486
rect 1143 474 1152 486
rect 1100 410 1109 422
rect 1143 410 1152 422
rect 1100 350 1152 358
rect 1100 346 1109 350
rect 1143 346 1152 350
rect 1100 282 1152 294
rect 1100 218 1152 230
rect 1100 160 1152 166
rect 1208 1142 1266 1370
rect 1322 1300 1542 1320
rect 1322 1220 1342 1300
rect 1422 1234 1442 1300
rect 1522 1234 1542 1300
rect 1322 1200 1345 1220
rect 1379 1200 1417 1220
rect 1451 1200 1489 1220
rect 1523 1200 1542 1234
rect 1333 1188 1535 1200
rect 1208 1108 1220 1142
rect 1254 1108 1266 1142
rect 1208 1070 1266 1108
rect 1208 1036 1220 1070
rect 1254 1036 1266 1070
rect 1208 998 1266 1036
rect 1208 964 1220 998
rect 1254 964 1266 998
rect 1208 926 1266 964
rect 1208 892 1220 926
rect 1254 892 1266 926
rect 1208 854 1266 892
rect 1208 820 1220 854
rect 1254 820 1266 854
rect 1208 782 1266 820
rect 1208 748 1220 782
rect 1254 748 1266 782
rect 1208 710 1266 748
rect 1208 676 1220 710
rect 1254 676 1266 710
rect 1208 638 1266 676
rect 1208 604 1220 638
rect 1254 604 1266 638
rect 1208 566 1266 604
rect 1208 532 1220 566
rect 1254 532 1266 566
rect 1208 494 1266 532
rect 1208 460 1220 494
rect 1254 460 1266 494
rect 1208 422 1266 460
rect 1208 388 1220 422
rect 1254 388 1266 422
rect 1208 350 1266 388
rect 1208 316 1220 350
rect 1254 316 1266 350
rect 1208 278 1266 316
rect 1208 244 1220 278
rect 1254 244 1266 278
rect 1208 206 1266 244
rect 1208 172 1220 206
rect 1254 172 1266 206
rect 1208 160 1266 172
rect 1322 1142 1374 1154
rect 1322 1108 1331 1142
rect 1365 1108 1374 1142
rect 1322 1070 1374 1108
rect 1322 1036 1331 1070
rect 1365 1036 1374 1070
rect 1322 998 1374 1036
rect 1322 964 1331 998
rect 1365 964 1374 998
rect 1322 926 1374 964
rect 1322 892 1331 926
rect 1365 892 1374 926
rect 1322 854 1374 892
rect 1322 820 1331 854
rect 1365 820 1374 854
rect 1322 782 1374 820
rect 1322 748 1331 782
rect 1365 748 1374 782
rect 1322 710 1374 748
rect 1322 676 1331 710
rect 1365 676 1374 710
rect 1322 638 1374 676
rect 1322 604 1331 638
rect 1365 604 1374 638
rect 1322 602 1374 604
rect 1322 538 1331 550
rect 1365 538 1374 550
rect 1322 474 1331 486
rect 1365 474 1374 486
rect 1322 410 1331 422
rect 1365 410 1374 422
rect 1322 350 1374 358
rect 1322 346 1331 350
rect 1365 346 1374 350
rect 1322 282 1374 294
rect 1322 218 1374 230
rect 1322 160 1374 166
rect 1408 1148 1460 1154
rect 1408 1084 1460 1096
rect 1408 1020 1460 1032
rect 1408 964 1417 968
rect 1451 964 1460 968
rect 1408 956 1460 964
rect 1408 892 1417 904
rect 1451 892 1460 904
rect 1408 828 1417 840
rect 1451 828 1460 840
rect 1408 764 1417 776
rect 1451 764 1460 776
rect 1408 710 1460 712
rect 1408 676 1417 710
rect 1451 676 1460 710
rect 1408 638 1460 676
rect 1408 604 1417 638
rect 1451 604 1460 638
rect 1408 566 1460 604
rect 1408 532 1417 566
rect 1451 532 1460 566
rect 1408 494 1460 532
rect 1408 460 1417 494
rect 1451 460 1460 494
rect 1408 422 1460 460
rect 1408 388 1417 422
rect 1451 388 1460 422
rect 1408 350 1460 388
rect 1408 316 1417 350
rect 1451 316 1460 350
rect 1408 278 1460 316
rect 1408 244 1417 278
rect 1451 244 1460 278
rect 1408 206 1460 244
rect 1408 172 1417 206
rect 1451 172 1460 206
rect 1408 160 1460 172
rect 1494 1142 1546 1154
rect 1494 1108 1503 1142
rect 1537 1108 1546 1142
rect 1494 1070 1546 1108
rect 1494 1036 1503 1070
rect 1537 1036 1546 1070
rect 1494 998 1546 1036
rect 1494 964 1503 998
rect 1537 964 1546 998
rect 1494 926 1546 964
rect 1494 892 1503 926
rect 1537 892 1546 926
rect 1494 854 1546 892
rect 1494 820 1503 854
rect 1537 820 1546 854
rect 1494 782 1546 820
rect 1494 748 1503 782
rect 1537 748 1546 782
rect 1494 710 1546 748
rect 1494 676 1503 710
rect 1537 676 1546 710
rect 1494 638 1546 676
rect 1494 604 1503 638
rect 1537 604 1546 638
rect 1494 602 1546 604
rect 1494 538 1503 550
rect 1537 538 1546 550
rect 1494 474 1503 486
rect 1537 474 1546 486
rect 1494 410 1503 422
rect 1537 410 1546 422
rect 1494 350 1546 358
rect 1494 346 1503 350
rect 1537 346 1546 350
rect 1494 282 1546 294
rect 1494 218 1546 230
rect 1494 160 1546 166
rect 1602 1142 1660 1370
rect 1712 1300 1932 1320
rect 1712 1220 1732 1300
rect 1812 1234 1832 1300
rect 1912 1234 1932 1300
rect 1712 1200 1739 1220
rect 1773 1200 1811 1220
rect 1845 1200 1883 1220
rect 1917 1200 1932 1234
rect 1723 1188 1929 1200
rect 1602 1108 1614 1142
rect 1648 1108 1660 1142
rect 1602 1070 1660 1108
rect 1602 1036 1614 1070
rect 1648 1036 1660 1070
rect 1602 998 1660 1036
rect 1602 964 1614 998
rect 1648 964 1660 998
rect 1602 926 1660 964
rect 1602 892 1614 926
rect 1648 892 1660 926
rect 1602 854 1660 892
rect 1602 820 1614 854
rect 1648 820 1660 854
rect 1602 782 1660 820
rect 1602 748 1614 782
rect 1648 748 1660 782
rect 1602 710 1660 748
rect 1602 676 1614 710
rect 1648 676 1660 710
rect 1602 638 1660 676
rect 1602 604 1614 638
rect 1648 604 1660 638
rect 1602 566 1660 604
rect 1602 532 1614 566
rect 1648 532 1660 566
rect 1602 494 1660 532
rect 1602 460 1614 494
rect 1648 460 1660 494
rect 1602 422 1660 460
rect 1602 388 1614 422
rect 1648 388 1660 422
rect 1602 350 1660 388
rect 1602 316 1614 350
rect 1648 316 1660 350
rect 1602 278 1660 316
rect 1602 244 1614 278
rect 1648 244 1660 278
rect 1602 206 1660 244
rect 1602 172 1614 206
rect 1648 172 1660 206
rect 1602 160 1660 172
rect 1716 1142 1768 1154
rect 1716 1108 1725 1142
rect 1759 1108 1768 1142
rect 1716 1070 1768 1108
rect 1716 1036 1725 1070
rect 1759 1036 1768 1070
rect 1716 998 1768 1036
rect 1716 964 1725 998
rect 1759 964 1768 998
rect 1716 926 1768 964
rect 1716 892 1725 926
rect 1759 892 1768 926
rect 1716 854 1768 892
rect 1716 820 1725 854
rect 1759 820 1768 854
rect 1716 782 1768 820
rect 1716 748 1725 782
rect 1759 748 1768 782
rect 1716 710 1768 748
rect 1716 676 1725 710
rect 1759 676 1768 710
rect 1716 638 1768 676
rect 1716 604 1725 638
rect 1759 604 1768 638
rect 1716 602 1768 604
rect 1716 538 1725 550
rect 1759 538 1768 550
rect 1716 474 1725 486
rect 1759 474 1768 486
rect 1716 410 1725 422
rect 1759 410 1768 422
rect 1716 350 1768 358
rect 1716 346 1725 350
rect 1759 346 1768 350
rect 1716 282 1768 294
rect 1716 218 1768 230
rect 1716 160 1768 166
rect 1802 1148 1854 1154
rect 1802 1084 1854 1096
rect 1802 1020 1854 1032
rect 1802 964 1811 968
rect 1845 964 1854 968
rect 1802 956 1854 964
rect 1802 892 1811 904
rect 1845 892 1854 904
rect 1802 828 1811 840
rect 1845 828 1854 840
rect 1802 764 1811 776
rect 1845 764 1854 776
rect 1802 710 1854 712
rect 1802 676 1811 710
rect 1845 676 1854 710
rect 1802 638 1854 676
rect 1802 604 1811 638
rect 1845 604 1854 638
rect 1802 566 1854 604
rect 1802 532 1811 566
rect 1845 532 1854 566
rect 1802 494 1854 532
rect 1802 460 1811 494
rect 1845 460 1854 494
rect 1802 422 1854 460
rect 1802 388 1811 422
rect 1845 388 1854 422
rect 1802 350 1854 388
rect 1802 316 1811 350
rect 1845 316 1854 350
rect 1802 278 1854 316
rect 1802 244 1811 278
rect 1845 244 1854 278
rect 1802 206 1854 244
rect 1802 172 1811 206
rect 1845 172 1854 206
rect 1802 160 1854 172
rect 1888 1142 1940 1154
rect 1888 1108 1897 1142
rect 1931 1108 1940 1142
rect 1888 1070 1940 1108
rect 1888 1036 1897 1070
rect 1931 1036 1940 1070
rect 1888 998 1940 1036
rect 1888 964 1897 998
rect 1931 964 1940 998
rect 1888 926 1940 964
rect 1888 892 1897 926
rect 1931 892 1940 926
rect 1888 854 1940 892
rect 1888 820 1897 854
rect 1931 820 1940 854
rect 1888 782 1940 820
rect 1888 748 1897 782
rect 1931 748 1940 782
rect 1888 710 1940 748
rect 1888 676 1897 710
rect 1931 676 1940 710
rect 1888 638 1940 676
rect 1888 604 1897 638
rect 1931 604 1940 638
rect 1888 602 1940 604
rect 1888 538 1897 550
rect 1931 538 1940 550
rect 1888 474 1897 486
rect 1931 474 1940 486
rect 1888 410 1897 422
rect 1931 410 1940 422
rect 1888 350 1940 358
rect 1888 346 1897 350
rect 1931 346 1940 350
rect 1888 282 1940 294
rect 1888 218 1940 230
rect 1888 160 1940 166
rect 1996 1142 2054 1370
rect 2112 1300 2332 1320
rect 2112 1220 2132 1300
rect 2212 1234 2232 1300
rect 2312 1220 2332 1300
rect 2112 1200 2133 1220
rect 2167 1200 2205 1220
rect 2239 1200 2277 1220
rect 2311 1200 2332 1220
rect 2121 1188 2325 1200
rect 1996 1108 2008 1142
rect 2042 1108 2054 1142
rect 1996 1070 2054 1108
rect 1996 1036 2008 1070
rect 2042 1036 2054 1070
rect 1996 998 2054 1036
rect 1996 964 2008 998
rect 2042 964 2054 998
rect 1996 926 2054 964
rect 1996 892 2008 926
rect 2042 892 2054 926
rect 1996 854 2054 892
rect 1996 820 2008 854
rect 2042 820 2054 854
rect 1996 782 2054 820
rect 1996 748 2008 782
rect 2042 748 2054 782
rect 1996 710 2054 748
rect 1996 676 2008 710
rect 2042 676 2054 710
rect 1996 638 2054 676
rect 1996 604 2008 638
rect 2042 604 2054 638
rect 1996 566 2054 604
rect 1996 532 2008 566
rect 2042 532 2054 566
rect 1996 494 2054 532
rect 1996 460 2008 494
rect 2042 460 2054 494
rect 1996 422 2054 460
rect 1996 388 2008 422
rect 2042 388 2054 422
rect 1996 350 2054 388
rect 1996 316 2008 350
rect 2042 316 2054 350
rect 1996 278 2054 316
rect 1996 244 2008 278
rect 2042 244 2054 278
rect 1996 206 2054 244
rect 1996 172 2008 206
rect 2042 172 2054 206
rect 1996 160 2054 172
rect 2110 1142 2162 1154
rect 2110 1108 2119 1142
rect 2153 1108 2162 1142
rect 2110 1070 2162 1108
rect 2110 1036 2119 1070
rect 2153 1036 2162 1070
rect 2110 998 2162 1036
rect 2110 964 2119 998
rect 2153 964 2162 998
rect 2110 926 2162 964
rect 2110 892 2119 926
rect 2153 892 2162 926
rect 2110 854 2162 892
rect 2110 820 2119 854
rect 2153 820 2162 854
rect 2110 782 2162 820
rect 2110 748 2119 782
rect 2153 748 2162 782
rect 2110 710 2162 748
rect 2110 676 2119 710
rect 2153 676 2162 710
rect 2110 638 2162 676
rect 2110 604 2119 638
rect 2153 604 2162 638
rect 2110 602 2162 604
rect 2110 538 2119 550
rect 2153 538 2162 550
rect 2110 474 2119 486
rect 2153 474 2162 486
rect 2110 410 2119 422
rect 2153 410 2162 422
rect 2110 350 2162 358
rect 2110 346 2119 350
rect 2153 346 2162 350
rect 2110 282 2162 294
rect 2110 218 2162 230
rect 2110 160 2162 166
rect 2196 1148 2248 1154
rect 2196 1084 2248 1096
rect 2196 1020 2248 1032
rect 2196 964 2205 968
rect 2239 964 2248 968
rect 2196 956 2248 964
rect 2196 892 2205 904
rect 2239 892 2248 904
rect 2196 828 2205 840
rect 2239 828 2248 840
rect 2196 764 2205 776
rect 2239 764 2248 776
rect 2196 710 2248 712
rect 2196 676 2205 710
rect 2239 676 2248 710
rect 2196 638 2248 676
rect 2196 604 2205 638
rect 2239 604 2248 638
rect 2196 566 2248 604
rect 2196 532 2205 566
rect 2239 532 2248 566
rect 2196 494 2248 532
rect 2196 460 2205 494
rect 2239 460 2248 494
rect 2196 422 2248 460
rect 2196 388 2205 422
rect 2239 388 2248 422
rect 2196 350 2248 388
rect 2196 316 2205 350
rect 2239 316 2248 350
rect 2196 278 2248 316
rect 2196 244 2205 278
rect 2239 244 2248 278
rect 2196 206 2248 244
rect 2196 172 2205 206
rect 2239 172 2248 206
rect 2196 160 2248 172
rect 2282 1142 2334 1154
rect 2282 1108 2291 1142
rect 2325 1108 2334 1142
rect 2282 1070 2334 1108
rect 2282 1036 2291 1070
rect 2325 1036 2334 1070
rect 2282 998 2334 1036
rect 2282 964 2291 998
rect 2325 964 2334 998
rect 2282 926 2334 964
rect 2282 892 2291 926
rect 2325 892 2334 926
rect 2282 854 2334 892
rect 2282 820 2291 854
rect 2325 820 2334 854
rect 2282 782 2334 820
rect 2282 748 2291 782
rect 2325 748 2334 782
rect 2282 710 2334 748
rect 2282 676 2291 710
rect 2325 676 2334 710
rect 2282 638 2334 676
rect 2282 604 2291 638
rect 2325 604 2334 638
rect 2282 602 2334 604
rect 2282 538 2291 550
rect 2325 538 2334 550
rect 2282 474 2291 486
rect 2325 474 2334 486
rect 2282 410 2291 422
rect 2325 410 2334 422
rect 2282 350 2334 358
rect 2282 346 2291 350
rect 2325 346 2334 350
rect 2282 282 2334 294
rect 2282 218 2334 230
rect 2282 160 2334 166
rect 2390 1142 2448 1370
rect 2390 1108 2402 1142
rect 2436 1108 2448 1142
rect 2390 1070 2448 1108
rect 2390 1036 2402 1070
rect 2436 1036 2448 1070
rect 2390 998 2448 1036
rect 2390 964 2402 998
rect 2436 964 2448 998
rect 2390 926 2448 964
rect 2390 892 2402 926
rect 2436 892 2448 926
rect 2390 854 2448 892
rect 2390 820 2402 854
rect 2436 820 2448 854
rect 2390 782 2448 820
rect 2390 748 2402 782
rect 2436 748 2448 782
rect 2390 710 2448 748
rect 2390 676 2402 710
rect 2436 676 2448 710
rect 2390 638 2448 676
rect 2390 604 2402 638
rect 2436 604 2448 638
rect 2390 566 2448 604
rect 2390 532 2402 566
rect 2436 532 2448 566
rect 2390 494 2448 532
rect 2390 460 2402 494
rect 2436 460 2448 494
rect 2390 422 2448 460
rect 2390 388 2402 422
rect 2436 388 2448 422
rect 2390 350 2448 388
rect 2390 316 2402 350
rect 2436 316 2448 350
rect 2390 278 2448 316
rect 2390 244 2402 278
rect 2436 244 2448 278
rect 2390 206 2448 244
rect 2390 172 2402 206
rect 2436 172 2448 206
rect 2390 160 2448 172
rect 151 120 353 132
rect 541 126 743 132
rect 941 126 1143 132
rect 541 120 747 126
rect 939 120 1143 126
rect 1333 120 1535 132
rect 1723 126 1925 132
rect 2123 126 2325 132
rect 1723 120 1929 126
rect 2121 120 2325 126
rect 140 114 360 120
rect 140 100 163 114
rect 197 100 235 114
rect 269 100 307 114
rect 140 20 160 100
rect 341 80 360 114
rect 240 20 260 80
rect 340 20 360 80
rect 140 0 360 20
rect 530 114 750 120
rect 530 100 557 114
rect 591 100 629 114
rect 663 100 701 114
rect 530 20 550 100
rect 735 80 750 114
rect 630 20 650 80
rect 730 20 750 80
rect 530 0 750 20
rect 930 114 1150 120
rect 930 100 951 114
rect 985 100 1023 114
rect 1057 100 1095 114
rect 1129 100 1150 114
rect 930 20 950 100
rect 1030 20 1050 80
rect 1130 20 1150 100
rect 930 0 1150 20
rect 1322 114 1542 120
rect 1322 100 1345 114
rect 1379 100 1417 114
rect 1451 100 1489 114
rect 1322 20 1342 100
rect 1523 80 1542 114
rect 1422 20 1442 80
rect 1522 20 1542 80
rect 1322 0 1542 20
rect 1712 114 1932 120
rect 1712 100 1739 114
rect 1773 100 1811 114
rect 1845 100 1883 114
rect 1712 20 1732 100
rect 1917 80 1932 114
rect 1812 20 1832 80
rect 1912 20 1932 80
rect 1712 0 1932 20
rect 2112 114 2332 120
rect 2112 100 2133 114
rect 2167 100 2205 114
rect 2239 100 2277 114
rect 2311 100 2332 114
rect 2112 20 2132 100
rect 2212 20 2232 80
rect 2312 20 2332 100
rect 2112 0 2332 20
<< via1 >>
rect 160 1234 240 1300
rect 260 1234 340 1300
rect 160 1220 163 1234
rect 163 1220 197 1234
rect 197 1220 235 1234
rect 235 1220 240 1234
rect 260 1220 269 1234
rect 269 1220 307 1234
rect 307 1220 340 1234
rect 140 566 192 602
rect 140 550 149 566
rect 149 550 183 566
rect 183 550 192 566
rect 140 532 149 538
rect 149 532 183 538
rect 183 532 192 538
rect 140 494 192 532
rect 140 486 149 494
rect 149 486 183 494
rect 183 486 192 494
rect 140 460 149 474
rect 149 460 183 474
rect 183 460 192 474
rect 140 422 192 460
rect 140 388 149 410
rect 149 388 183 410
rect 183 388 192 410
rect 140 358 192 388
rect 140 316 149 346
rect 149 316 183 346
rect 183 316 192 346
rect 140 294 192 316
rect 140 278 192 282
rect 140 244 149 278
rect 149 244 183 278
rect 183 244 192 278
rect 140 230 192 244
rect 140 206 192 218
rect 140 172 149 206
rect 149 172 183 206
rect 183 172 192 206
rect 140 166 192 172
rect 226 1142 278 1148
rect 226 1108 235 1142
rect 235 1108 269 1142
rect 269 1108 278 1142
rect 226 1096 278 1108
rect 226 1070 278 1084
rect 226 1036 235 1070
rect 235 1036 269 1070
rect 269 1036 278 1070
rect 226 1032 278 1036
rect 226 998 278 1020
rect 226 968 235 998
rect 235 968 269 998
rect 269 968 278 998
rect 226 926 278 956
rect 226 904 235 926
rect 235 904 269 926
rect 269 904 278 926
rect 226 854 278 892
rect 226 840 235 854
rect 235 840 269 854
rect 269 840 278 854
rect 226 820 235 828
rect 235 820 269 828
rect 269 820 278 828
rect 226 782 278 820
rect 226 776 235 782
rect 235 776 269 782
rect 269 776 278 782
rect 226 748 235 764
rect 235 748 269 764
rect 269 748 278 764
rect 226 712 278 748
rect 312 566 364 602
rect 312 550 321 566
rect 321 550 355 566
rect 355 550 364 566
rect 312 532 321 538
rect 321 532 355 538
rect 355 532 364 538
rect 312 494 364 532
rect 312 486 321 494
rect 321 486 355 494
rect 355 486 364 494
rect 312 460 321 474
rect 321 460 355 474
rect 355 460 364 474
rect 312 422 364 460
rect 312 388 321 410
rect 321 388 355 410
rect 355 388 364 410
rect 312 358 364 388
rect 312 316 321 346
rect 321 316 355 346
rect 355 316 364 346
rect 312 294 364 316
rect 312 278 364 282
rect 312 244 321 278
rect 321 244 355 278
rect 355 244 364 278
rect 312 230 364 244
rect 312 206 364 218
rect 312 172 321 206
rect 321 172 355 206
rect 355 172 364 206
rect 312 166 364 172
rect 550 1234 630 1300
rect 650 1234 730 1300
rect 550 1220 557 1234
rect 557 1220 591 1234
rect 591 1220 629 1234
rect 629 1220 630 1234
rect 650 1220 663 1234
rect 663 1220 701 1234
rect 701 1220 730 1234
rect 534 566 586 602
rect 534 550 543 566
rect 543 550 577 566
rect 577 550 586 566
rect 534 532 543 538
rect 543 532 577 538
rect 577 532 586 538
rect 534 494 586 532
rect 534 486 543 494
rect 543 486 577 494
rect 577 486 586 494
rect 534 460 543 474
rect 543 460 577 474
rect 577 460 586 474
rect 534 422 586 460
rect 534 388 543 410
rect 543 388 577 410
rect 577 388 586 410
rect 534 358 586 388
rect 534 316 543 346
rect 543 316 577 346
rect 577 316 586 346
rect 534 294 586 316
rect 534 278 586 282
rect 534 244 543 278
rect 543 244 577 278
rect 577 244 586 278
rect 534 230 586 244
rect 534 206 586 218
rect 534 172 543 206
rect 543 172 577 206
rect 577 172 586 206
rect 534 166 586 172
rect 620 1142 672 1148
rect 620 1108 629 1142
rect 629 1108 663 1142
rect 663 1108 672 1142
rect 620 1096 672 1108
rect 620 1070 672 1084
rect 620 1036 629 1070
rect 629 1036 663 1070
rect 663 1036 672 1070
rect 620 1032 672 1036
rect 620 998 672 1020
rect 620 968 629 998
rect 629 968 663 998
rect 663 968 672 998
rect 620 926 672 956
rect 620 904 629 926
rect 629 904 663 926
rect 663 904 672 926
rect 620 854 672 892
rect 620 840 629 854
rect 629 840 663 854
rect 663 840 672 854
rect 620 820 629 828
rect 629 820 663 828
rect 663 820 672 828
rect 620 782 672 820
rect 620 776 629 782
rect 629 776 663 782
rect 663 776 672 782
rect 620 748 629 764
rect 629 748 663 764
rect 663 748 672 764
rect 620 712 672 748
rect 706 566 758 602
rect 706 550 715 566
rect 715 550 749 566
rect 749 550 758 566
rect 706 532 715 538
rect 715 532 749 538
rect 749 532 758 538
rect 706 494 758 532
rect 706 486 715 494
rect 715 486 749 494
rect 749 486 758 494
rect 706 460 715 474
rect 715 460 749 474
rect 749 460 758 474
rect 706 422 758 460
rect 706 388 715 410
rect 715 388 749 410
rect 749 388 758 410
rect 706 358 758 388
rect 706 316 715 346
rect 715 316 749 346
rect 749 316 758 346
rect 706 294 758 316
rect 706 278 758 282
rect 706 244 715 278
rect 715 244 749 278
rect 749 244 758 278
rect 706 230 758 244
rect 706 206 758 218
rect 706 172 715 206
rect 715 172 749 206
rect 749 172 758 206
rect 706 166 758 172
rect 950 1234 1030 1300
rect 1050 1234 1130 1300
rect 950 1220 951 1234
rect 951 1220 985 1234
rect 985 1220 1023 1234
rect 1023 1220 1030 1234
rect 1050 1220 1057 1234
rect 1057 1220 1095 1234
rect 1095 1220 1129 1234
rect 1129 1220 1130 1234
rect 928 566 980 602
rect 928 550 937 566
rect 937 550 971 566
rect 971 550 980 566
rect 928 532 937 538
rect 937 532 971 538
rect 971 532 980 538
rect 928 494 980 532
rect 928 486 937 494
rect 937 486 971 494
rect 971 486 980 494
rect 928 460 937 474
rect 937 460 971 474
rect 971 460 980 474
rect 928 422 980 460
rect 928 388 937 410
rect 937 388 971 410
rect 971 388 980 410
rect 928 358 980 388
rect 928 316 937 346
rect 937 316 971 346
rect 971 316 980 346
rect 928 294 980 316
rect 928 278 980 282
rect 928 244 937 278
rect 937 244 971 278
rect 971 244 980 278
rect 928 230 980 244
rect 928 206 980 218
rect 928 172 937 206
rect 937 172 971 206
rect 971 172 980 206
rect 928 166 980 172
rect 1014 1142 1066 1148
rect 1014 1108 1023 1142
rect 1023 1108 1057 1142
rect 1057 1108 1066 1142
rect 1014 1096 1066 1108
rect 1014 1070 1066 1084
rect 1014 1036 1023 1070
rect 1023 1036 1057 1070
rect 1057 1036 1066 1070
rect 1014 1032 1066 1036
rect 1014 998 1066 1020
rect 1014 968 1023 998
rect 1023 968 1057 998
rect 1057 968 1066 998
rect 1014 926 1066 956
rect 1014 904 1023 926
rect 1023 904 1057 926
rect 1057 904 1066 926
rect 1014 854 1066 892
rect 1014 840 1023 854
rect 1023 840 1057 854
rect 1057 840 1066 854
rect 1014 820 1023 828
rect 1023 820 1057 828
rect 1057 820 1066 828
rect 1014 782 1066 820
rect 1014 776 1023 782
rect 1023 776 1057 782
rect 1057 776 1066 782
rect 1014 748 1023 764
rect 1023 748 1057 764
rect 1057 748 1066 764
rect 1014 712 1066 748
rect 1100 566 1152 602
rect 1100 550 1109 566
rect 1109 550 1143 566
rect 1143 550 1152 566
rect 1100 532 1109 538
rect 1109 532 1143 538
rect 1143 532 1152 538
rect 1100 494 1152 532
rect 1100 486 1109 494
rect 1109 486 1143 494
rect 1143 486 1152 494
rect 1100 460 1109 474
rect 1109 460 1143 474
rect 1143 460 1152 474
rect 1100 422 1152 460
rect 1100 388 1109 410
rect 1109 388 1143 410
rect 1143 388 1152 410
rect 1100 358 1152 388
rect 1100 316 1109 346
rect 1109 316 1143 346
rect 1143 316 1152 346
rect 1100 294 1152 316
rect 1100 278 1152 282
rect 1100 244 1109 278
rect 1109 244 1143 278
rect 1143 244 1152 278
rect 1100 230 1152 244
rect 1100 206 1152 218
rect 1100 172 1109 206
rect 1109 172 1143 206
rect 1143 172 1152 206
rect 1100 166 1152 172
rect 1342 1234 1422 1300
rect 1442 1234 1522 1300
rect 1342 1220 1345 1234
rect 1345 1220 1379 1234
rect 1379 1220 1417 1234
rect 1417 1220 1422 1234
rect 1442 1220 1451 1234
rect 1451 1220 1489 1234
rect 1489 1220 1522 1234
rect 1322 566 1374 602
rect 1322 550 1331 566
rect 1331 550 1365 566
rect 1365 550 1374 566
rect 1322 532 1331 538
rect 1331 532 1365 538
rect 1365 532 1374 538
rect 1322 494 1374 532
rect 1322 486 1331 494
rect 1331 486 1365 494
rect 1365 486 1374 494
rect 1322 460 1331 474
rect 1331 460 1365 474
rect 1365 460 1374 474
rect 1322 422 1374 460
rect 1322 388 1331 410
rect 1331 388 1365 410
rect 1365 388 1374 410
rect 1322 358 1374 388
rect 1322 316 1331 346
rect 1331 316 1365 346
rect 1365 316 1374 346
rect 1322 294 1374 316
rect 1322 278 1374 282
rect 1322 244 1331 278
rect 1331 244 1365 278
rect 1365 244 1374 278
rect 1322 230 1374 244
rect 1322 206 1374 218
rect 1322 172 1331 206
rect 1331 172 1365 206
rect 1365 172 1374 206
rect 1322 166 1374 172
rect 1408 1142 1460 1148
rect 1408 1108 1417 1142
rect 1417 1108 1451 1142
rect 1451 1108 1460 1142
rect 1408 1096 1460 1108
rect 1408 1070 1460 1084
rect 1408 1036 1417 1070
rect 1417 1036 1451 1070
rect 1451 1036 1460 1070
rect 1408 1032 1460 1036
rect 1408 998 1460 1020
rect 1408 968 1417 998
rect 1417 968 1451 998
rect 1451 968 1460 998
rect 1408 926 1460 956
rect 1408 904 1417 926
rect 1417 904 1451 926
rect 1451 904 1460 926
rect 1408 854 1460 892
rect 1408 840 1417 854
rect 1417 840 1451 854
rect 1451 840 1460 854
rect 1408 820 1417 828
rect 1417 820 1451 828
rect 1451 820 1460 828
rect 1408 782 1460 820
rect 1408 776 1417 782
rect 1417 776 1451 782
rect 1451 776 1460 782
rect 1408 748 1417 764
rect 1417 748 1451 764
rect 1451 748 1460 764
rect 1408 712 1460 748
rect 1494 566 1546 602
rect 1494 550 1503 566
rect 1503 550 1537 566
rect 1537 550 1546 566
rect 1494 532 1503 538
rect 1503 532 1537 538
rect 1537 532 1546 538
rect 1494 494 1546 532
rect 1494 486 1503 494
rect 1503 486 1537 494
rect 1537 486 1546 494
rect 1494 460 1503 474
rect 1503 460 1537 474
rect 1537 460 1546 474
rect 1494 422 1546 460
rect 1494 388 1503 410
rect 1503 388 1537 410
rect 1537 388 1546 410
rect 1494 358 1546 388
rect 1494 316 1503 346
rect 1503 316 1537 346
rect 1537 316 1546 346
rect 1494 294 1546 316
rect 1494 278 1546 282
rect 1494 244 1503 278
rect 1503 244 1537 278
rect 1537 244 1546 278
rect 1494 230 1546 244
rect 1494 206 1546 218
rect 1494 172 1503 206
rect 1503 172 1537 206
rect 1537 172 1546 206
rect 1494 166 1546 172
rect 1732 1234 1812 1300
rect 1832 1234 1912 1300
rect 1732 1220 1739 1234
rect 1739 1220 1773 1234
rect 1773 1220 1811 1234
rect 1811 1220 1812 1234
rect 1832 1220 1845 1234
rect 1845 1220 1883 1234
rect 1883 1220 1912 1234
rect 1716 566 1768 602
rect 1716 550 1725 566
rect 1725 550 1759 566
rect 1759 550 1768 566
rect 1716 532 1725 538
rect 1725 532 1759 538
rect 1759 532 1768 538
rect 1716 494 1768 532
rect 1716 486 1725 494
rect 1725 486 1759 494
rect 1759 486 1768 494
rect 1716 460 1725 474
rect 1725 460 1759 474
rect 1759 460 1768 474
rect 1716 422 1768 460
rect 1716 388 1725 410
rect 1725 388 1759 410
rect 1759 388 1768 410
rect 1716 358 1768 388
rect 1716 316 1725 346
rect 1725 316 1759 346
rect 1759 316 1768 346
rect 1716 294 1768 316
rect 1716 278 1768 282
rect 1716 244 1725 278
rect 1725 244 1759 278
rect 1759 244 1768 278
rect 1716 230 1768 244
rect 1716 206 1768 218
rect 1716 172 1725 206
rect 1725 172 1759 206
rect 1759 172 1768 206
rect 1716 166 1768 172
rect 1802 1142 1854 1148
rect 1802 1108 1811 1142
rect 1811 1108 1845 1142
rect 1845 1108 1854 1142
rect 1802 1096 1854 1108
rect 1802 1070 1854 1084
rect 1802 1036 1811 1070
rect 1811 1036 1845 1070
rect 1845 1036 1854 1070
rect 1802 1032 1854 1036
rect 1802 998 1854 1020
rect 1802 968 1811 998
rect 1811 968 1845 998
rect 1845 968 1854 998
rect 1802 926 1854 956
rect 1802 904 1811 926
rect 1811 904 1845 926
rect 1845 904 1854 926
rect 1802 854 1854 892
rect 1802 840 1811 854
rect 1811 840 1845 854
rect 1845 840 1854 854
rect 1802 820 1811 828
rect 1811 820 1845 828
rect 1845 820 1854 828
rect 1802 782 1854 820
rect 1802 776 1811 782
rect 1811 776 1845 782
rect 1845 776 1854 782
rect 1802 748 1811 764
rect 1811 748 1845 764
rect 1845 748 1854 764
rect 1802 712 1854 748
rect 1888 566 1940 602
rect 1888 550 1897 566
rect 1897 550 1931 566
rect 1931 550 1940 566
rect 1888 532 1897 538
rect 1897 532 1931 538
rect 1931 532 1940 538
rect 1888 494 1940 532
rect 1888 486 1897 494
rect 1897 486 1931 494
rect 1931 486 1940 494
rect 1888 460 1897 474
rect 1897 460 1931 474
rect 1931 460 1940 474
rect 1888 422 1940 460
rect 1888 388 1897 410
rect 1897 388 1931 410
rect 1931 388 1940 410
rect 1888 358 1940 388
rect 1888 316 1897 346
rect 1897 316 1931 346
rect 1931 316 1940 346
rect 1888 294 1940 316
rect 1888 278 1940 282
rect 1888 244 1897 278
rect 1897 244 1931 278
rect 1931 244 1940 278
rect 1888 230 1940 244
rect 1888 206 1940 218
rect 1888 172 1897 206
rect 1897 172 1931 206
rect 1931 172 1940 206
rect 1888 166 1940 172
rect 2132 1234 2212 1300
rect 2232 1234 2312 1300
rect 2132 1220 2133 1234
rect 2133 1220 2167 1234
rect 2167 1220 2205 1234
rect 2205 1220 2212 1234
rect 2232 1220 2239 1234
rect 2239 1220 2277 1234
rect 2277 1220 2311 1234
rect 2311 1220 2312 1234
rect 2110 566 2162 602
rect 2110 550 2119 566
rect 2119 550 2153 566
rect 2153 550 2162 566
rect 2110 532 2119 538
rect 2119 532 2153 538
rect 2153 532 2162 538
rect 2110 494 2162 532
rect 2110 486 2119 494
rect 2119 486 2153 494
rect 2153 486 2162 494
rect 2110 460 2119 474
rect 2119 460 2153 474
rect 2153 460 2162 474
rect 2110 422 2162 460
rect 2110 388 2119 410
rect 2119 388 2153 410
rect 2153 388 2162 410
rect 2110 358 2162 388
rect 2110 316 2119 346
rect 2119 316 2153 346
rect 2153 316 2162 346
rect 2110 294 2162 316
rect 2110 278 2162 282
rect 2110 244 2119 278
rect 2119 244 2153 278
rect 2153 244 2162 278
rect 2110 230 2162 244
rect 2110 206 2162 218
rect 2110 172 2119 206
rect 2119 172 2153 206
rect 2153 172 2162 206
rect 2110 166 2162 172
rect 2196 1142 2248 1148
rect 2196 1108 2205 1142
rect 2205 1108 2239 1142
rect 2239 1108 2248 1142
rect 2196 1096 2248 1108
rect 2196 1070 2248 1084
rect 2196 1036 2205 1070
rect 2205 1036 2239 1070
rect 2239 1036 2248 1070
rect 2196 1032 2248 1036
rect 2196 998 2248 1020
rect 2196 968 2205 998
rect 2205 968 2239 998
rect 2239 968 2248 998
rect 2196 926 2248 956
rect 2196 904 2205 926
rect 2205 904 2239 926
rect 2239 904 2248 926
rect 2196 854 2248 892
rect 2196 840 2205 854
rect 2205 840 2239 854
rect 2239 840 2248 854
rect 2196 820 2205 828
rect 2205 820 2239 828
rect 2239 820 2248 828
rect 2196 782 2248 820
rect 2196 776 2205 782
rect 2205 776 2239 782
rect 2239 776 2248 782
rect 2196 748 2205 764
rect 2205 748 2239 764
rect 2239 748 2248 764
rect 2196 712 2248 748
rect 2282 566 2334 602
rect 2282 550 2291 566
rect 2291 550 2325 566
rect 2325 550 2334 566
rect 2282 532 2291 538
rect 2291 532 2325 538
rect 2325 532 2334 538
rect 2282 494 2334 532
rect 2282 486 2291 494
rect 2291 486 2325 494
rect 2325 486 2334 494
rect 2282 460 2291 474
rect 2291 460 2325 474
rect 2325 460 2334 474
rect 2282 422 2334 460
rect 2282 388 2291 410
rect 2291 388 2325 410
rect 2325 388 2334 410
rect 2282 358 2334 388
rect 2282 316 2291 346
rect 2291 316 2325 346
rect 2325 316 2334 346
rect 2282 294 2334 316
rect 2282 278 2334 282
rect 2282 244 2291 278
rect 2291 244 2325 278
rect 2325 244 2334 278
rect 2282 230 2334 244
rect 2282 206 2334 218
rect 2282 172 2291 206
rect 2291 172 2325 206
rect 2325 172 2334 206
rect 2282 166 2334 172
rect 160 80 163 100
rect 163 80 197 100
rect 197 80 235 100
rect 235 80 240 100
rect 260 80 269 100
rect 269 80 307 100
rect 307 80 340 100
rect 160 20 240 80
rect 260 20 340 80
rect 550 80 557 100
rect 557 80 591 100
rect 591 80 629 100
rect 629 80 630 100
rect 650 80 663 100
rect 663 80 701 100
rect 701 80 730 100
rect 550 20 630 80
rect 650 20 730 80
rect 950 80 951 100
rect 951 80 985 100
rect 985 80 1023 100
rect 1023 80 1030 100
rect 1050 80 1057 100
rect 1057 80 1095 100
rect 1095 80 1129 100
rect 1129 80 1130 100
rect 950 20 1030 80
rect 1050 20 1130 80
rect 1342 80 1345 100
rect 1345 80 1379 100
rect 1379 80 1417 100
rect 1417 80 1422 100
rect 1442 80 1451 100
rect 1451 80 1489 100
rect 1489 80 1522 100
rect 1342 20 1422 80
rect 1442 20 1522 80
rect 1732 80 1739 100
rect 1739 80 1773 100
rect 1773 80 1811 100
rect 1811 80 1812 100
rect 1832 80 1845 100
rect 1845 80 1883 100
rect 1883 80 1912 100
rect 1732 20 1812 80
rect 1832 20 1912 80
rect 2132 80 2133 100
rect 2133 80 2167 100
rect 2167 80 2205 100
rect 2205 80 2212 100
rect 2232 80 2239 100
rect 2239 80 2277 100
rect 2277 80 2311 100
rect 2311 80 2312 100
rect 2132 20 2212 80
rect 2232 20 2312 80
<< metal2 >>
rect 140 1300 360 1320
rect 140 1220 160 1300
rect 240 1220 260 1300
rect 340 1220 360 1300
rect 140 1200 360 1220
rect 530 1300 750 1320
rect 530 1220 550 1300
rect 630 1220 650 1300
rect 730 1220 750 1300
rect 530 1200 750 1220
rect 930 1300 1150 1320
rect 930 1220 950 1300
rect 1030 1220 1050 1300
rect 1130 1220 1150 1300
rect 930 1200 1150 1220
rect 1322 1300 1542 1320
rect 1322 1220 1342 1300
rect 1422 1220 1442 1300
rect 1522 1220 1542 1300
rect 1322 1200 1542 1220
rect 1712 1300 1932 1320
rect 1712 1220 1732 1300
rect 1812 1220 1832 1300
rect 1912 1220 1932 1300
rect 1712 1200 1932 1220
rect 2112 1300 2332 1320
rect 2112 1220 2132 1300
rect 2212 1220 2232 1300
rect 2312 1220 2332 1300
rect 2112 1200 2332 1220
rect 0 1148 2474 1154
rect 0 1096 226 1148
rect 278 1096 620 1148
rect 672 1096 1014 1148
rect 1066 1096 1408 1148
rect 1460 1096 1802 1148
rect 1854 1096 2196 1148
rect 2248 1096 2474 1148
rect 0 1084 2474 1096
rect 0 1032 226 1084
rect 278 1032 620 1084
rect 672 1032 1014 1084
rect 1066 1032 1408 1084
rect 1460 1032 1802 1084
rect 1854 1032 2196 1084
rect 2248 1032 2474 1084
rect 0 1020 2474 1032
rect 0 968 226 1020
rect 278 968 620 1020
rect 672 968 1014 1020
rect 1066 968 1408 1020
rect 1460 968 1802 1020
rect 1854 968 2196 1020
rect 2248 968 2474 1020
rect 0 956 2474 968
rect 0 904 226 956
rect 278 904 620 956
rect 672 904 1014 956
rect 1066 904 1408 956
rect 1460 904 1802 956
rect 1854 904 2196 956
rect 2248 904 2474 956
rect 0 892 2474 904
rect 0 840 226 892
rect 278 840 620 892
rect 672 840 1014 892
rect 1066 840 1408 892
rect 1460 840 1802 892
rect 1854 840 2196 892
rect 2248 840 2474 892
rect 0 828 2474 840
rect 0 776 226 828
rect 278 776 620 828
rect 672 776 1014 828
rect 1066 776 1408 828
rect 1460 776 1802 828
rect 1854 776 2196 828
rect 2248 776 2474 828
rect 0 764 2474 776
rect 0 712 226 764
rect 278 712 620 764
rect 672 712 1014 764
rect 1066 712 1408 764
rect 1460 712 1802 764
rect 1854 712 2196 764
rect 2248 712 2474 764
rect 0 682 2474 712
rect 0 602 2474 632
rect 0 550 140 602
rect 192 550 312 602
rect 364 550 534 602
rect 586 550 706 602
rect 758 550 928 602
rect 980 550 1100 602
rect 1152 550 1322 602
rect 1374 550 1494 602
rect 1546 550 1716 602
rect 1768 550 1888 602
rect 1940 550 2110 602
rect 2162 550 2282 602
rect 2334 550 2474 602
rect 0 538 2474 550
rect 0 486 140 538
rect 192 486 312 538
rect 364 486 534 538
rect 586 486 706 538
rect 758 486 928 538
rect 980 486 1100 538
rect 1152 486 1322 538
rect 1374 486 1494 538
rect 1546 486 1716 538
rect 1768 486 1888 538
rect 1940 486 2110 538
rect 2162 486 2282 538
rect 2334 486 2474 538
rect 0 474 2474 486
rect 0 422 140 474
rect 192 422 312 474
rect 364 422 534 474
rect 586 422 706 474
rect 758 422 928 474
rect 980 422 1100 474
rect 1152 422 1322 474
rect 1374 422 1494 474
rect 1546 422 1716 474
rect 1768 422 1888 474
rect 1940 422 2110 474
rect 2162 422 2282 474
rect 2334 422 2474 474
rect 0 410 2474 422
rect 0 358 140 410
rect 192 358 312 410
rect 364 358 534 410
rect 586 358 706 410
rect 758 358 928 410
rect 980 358 1100 410
rect 1152 358 1322 410
rect 1374 358 1494 410
rect 1546 358 1716 410
rect 1768 358 1888 410
rect 1940 358 2110 410
rect 2162 358 2282 410
rect 2334 358 2474 410
rect 0 346 2474 358
rect 0 294 140 346
rect 192 294 312 346
rect 364 294 534 346
rect 586 294 706 346
rect 758 294 928 346
rect 980 294 1100 346
rect 1152 294 1322 346
rect 1374 294 1494 346
rect 1546 294 1716 346
rect 1768 294 1888 346
rect 1940 294 2110 346
rect 2162 294 2282 346
rect 2334 294 2474 346
rect 0 282 2474 294
rect 0 230 140 282
rect 192 230 312 282
rect 364 230 534 282
rect 586 230 706 282
rect 758 230 928 282
rect 980 230 1100 282
rect 1152 230 1322 282
rect 1374 230 1494 282
rect 1546 230 1716 282
rect 1768 230 1888 282
rect 1940 230 2110 282
rect 2162 230 2282 282
rect 2334 230 2474 282
rect 0 218 2474 230
rect 0 166 140 218
rect 192 166 312 218
rect 364 166 534 218
rect 586 166 706 218
rect 758 166 928 218
rect 980 166 1100 218
rect 1152 166 1322 218
rect 1374 166 1494 218
rect 1546 166 1716 218
rect 1768 166 1888 218
rect 1940 166 2110 218
rect 2162 166 2282 218
rect 2334 166 2474 218
rect 0 160 2474 166
rect 140 100 360 120
rect 140 20 160 100
rect 240 20 260 100
rect 340 20 360 100
rect 140 0 360 20
rect 530 100 750 120
rect 530 20 550 100
rect 630 20 650 100
rect 730 20 750 100
rect 530 0 750 20
rect 930 100 1150 120
rect 930 20 950 100
rect 1030 20 1050 100
rect 1130 20 1150 100
rect 930 0 1150 20
rect 1322 100 1542 120
rect 1322 20 1342 100
rect 1422 20 1442 100
rect 1522 20 1542 100
rect 1322 0 1542 20
rect 1712 100 1932 120
rect 1712 20 1732 100
rect 1812 20 1832 100
rect 1912 20 1932 100
rect 1712 0 1932 20
rect 2112 100 2332 120
rect 2112 20 2132 100
rect 2212 20 2232 100
rect 2312 20 2332 100
rect 2112 0 2332 20
<< via2 >>
rect 160 1220 230 1300
rect 270 1220 340 1300
rect 550 1220 620 1300
rect 660 1220 730 1300
rect 950 1220 1020 1300
rect 1060 1220 1130 1300
rect 1342 1220 1412 1300
rect 1452 1220 1522 1300
rect 1732 1220 1802 1300
rect 1842 1220 1912 1300
rect 2132 1220 2202 1300
rect 2242 1220 2312 1300
rect 160 20 230 100
rect 270 20 340 100
rect 550 20 620 100
rect 660 20 730 100
rect 950 20 1020 100
rect 1060 20 1130 100
rect 1342 20 1412 100
rect 1452 20 1522 100
rect 1732 20 1802 100
rect 1842 20 1912 100
rect 2132 20 2202 100
rect 2242 20 2312 100
<< metal3 >>
rect 140 1300 1150 1320
rect 140 1220 160 1300
rect 230 1220 270 1300
rect 340 1220 550 1300
rect 620 1220 660 1300
rect 730 1220 950 1300
rect 1020 1220 1060 1300
rect 1130 1220 1150 1300
rect 140 1200 1150 1220
rect 1322 1300 2332 1320
rect 1322 1220 1342 1300
rect 1412 1220 1452 1300
rect 1522 1220 1732 1300
rect 1802 1220 1842 1300
rect 1912 1220 2132 1300
rect 2202 1220 2242 1300
rect 2312 1220 2332 1300
rect 1322 1200 2332 1220
rect 400 700 500 1200
rect 800 700 900 1200
rect 1582 700 1682 1200
rect 1982 700 2082 1200
rect 400 600 2082 700
rect 400 120 500 600
rect 800 120 900 600
rect 1582 120 1682 600
rect 1982 120 2082 600
rect 140 100 1150 120
rect 140 20 160 100
rect 230 20 270 100
rect 340 20 550 100
rect 620 20 660 100
rect 730 20 950 100
rect 1020 20 1060 100
rect 1130 20 1150 100
rect 140 0 1150 20
rect 1322 100 2332 120
rect 1322 20 1342 100
rect 1412 20 1452 100
rect 1522 20 1732 100
rect 1802 20 1842 100
rect 1912 20 2132 100
rect 2202 20 2242 100
rect 2312 20 2332 100
rect 1322 0 2332 20
<< labels >>
rlabel metal2 0 682 20 1154 1 D
rlabel metal2 0 160 20 632 1 S
rlabel metal1 26 1370 86 1440 1 B
rlabel metal3 400 600 2082 700 1 G
rlabel metal1 1208 1370 2448 1440 1 nfet_3x_2_1/sub
rlabel metal3 1322 1200 2322 1320 1 nfet_3x_2_1/G
rlabel metal2 1182 682 2474 1154 1 nfet_3x_2_1/D
rlabel metal2 1182 160 2474 632 1 nfet_3x_2_1/S
flabel metal2 1970 682 1990 1154 7 FreeSans 300 180 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/DRAIN
flabel metal2 1970 160 1990 632 7 FreeSans 300 180 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SOURCE
flabel metal1 2390 160 2448 176 3 FreeSans 300 90 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SUBSTRATE
flabel metal1 1996 160 2054 176 3 FreeSans 300 90 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SUBSTRATE
flabel metal1 2121 1188 2323 1254 0 FreeSans 300 0 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE
flabel metal1 2121 60 2323 126 0 FreeSans 300 0 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE
flabel metal2 2060 682 2080 1154 3 FreeSans 300 180 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/DRAIN
flabel metal2 2060 160 2080 632 3 FreeSans 300 180 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SOURCE
flabel metal1 1602 160 1660 176 7 FreeSans 300 90 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SUBSTRATE
flabel metal1 1996 160 2054 176 7 FreeSans 300 90 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SUBSTRATE
flabel metal1 1727 1188 1929 1254 0 FreeSans 300 0 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE
flabel metal1 1727 60 1929 126 0 FreeSans 300 0 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE
flabel metal2 1182 682 1202 1154 7 FreeSans 300 180 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN
flabel metal2 1182 160 1202 632 7 FreeSans 300 180 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/SOURCE
flabel metal1 1602 160 1660 176 3 FreeSans 300 90 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/SUBSTRATE
flabel metal1 1208 160 1266 176 3 FreeSans 300 90 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/SUBSTRATE
flabel metal1 1333 1188 1535 1254 0 FreeSans 300 0 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE
flabel metal1 1333 60 1535 126 0 FreeSans 300 0 0 0 nfet_3x_2_1/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE
rlabel metal1 26 1370 1266 1440 1 nfet_3x_2_0/sub
rlabel metal3 140 1200 1140 1320 1 nfet_3x_2_0/G
rlabel metal2 0 682 1292 1154 1 nfet_3x_2_0/D
rlabel metal2 0 160 1292 632 1 nfet_3x_2_0/S
flabel metal2 788 682 808 1154 7 FreeSans 300 180 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/DRAIN
flabel metal2 788 160 808 632 7 FreeSans 300 180 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SOURCE
flabel metal1 1208 160 1266 176 3 FreeSans 300 90 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SUBSTRATE
flabel metal1 814 160 872 176 3 FreeSans 300 90 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SUBSTRATE
flabel metal1 939 1188 1141 1254 0 FreeSans 300 0 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE
flabel metal1 939 60 1141 126 0 FreeSans 300 0 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE
flabel metal2 878 682 898 1154 3 FreeSans 300 180 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/DRAIN
flabel metal2 878 160 898 632 3 FreeSans 300 180 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SOURCE
flabel metal1 420 160 478 176 7 FreeSans 300 90 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SUBSTRATE
flabel metal1 814 160 872 176 7 FreeSans 300 90 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SUBSTRATE
flabel metal1 545 1188 747 1254 0 FreeSans 300 0 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE
flabel metal1 545 60 747 126 0 FreeSans 300 0 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE
flabel metal2 0 682 20 1154 7 FreeSans 300 180 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN
flabel metal2 0 160 20 632 7 FreeSans 300 180 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/SOURCE
flabel metal1 420 160 478 176 3 FreeSans 300 90 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/SUBSTRATE
flabel metal1 26 160 84 176 3 FreeSans 300 90 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/SUBSTRATE
flabel metal1 151 1188 353 1254 0 FreeSans 300 0 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE
flabel metal1 151 60 353 126 0 FreeSans 300 0 0 0 nfet_3x_2_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE
<< end >>
