magic
tech sky130B
timestamp 1659901159
<< nwell >>
rect 0 -370 15 1110
rect 1190 -370 1205 1110
<< metal1 >>
rect 15 1060 110 1110
rect 160 1075 165 1110
rect 200 1075 205 1110
rect 280 1075 285 1110
rect 320 1075 325 1110
rect 400 1075 405 1110
rect 440 1075 445 1110
rect 520 1075 525 1110
rect 560 1075 565 1110
rect 640 1075 645 1110
rect 680 1075 685 1110
rect 760 1075 765 1110
rect 800 1075 805 1110
rect 880 1075 885 1110
rect 920 1075 925 1110
rect 1000 1075 1005 1110
rect 1040 1075 1045 1110
rect 1095 1060 1190 1110
rect 15 1055 45 1060
rect 15 960 19 1055
rect 15 955 45 960
rect 15 875 110 925
rect 160 890 165 925
rect 200 890 205 925
rect 280 890 285 925
rect 320 890 325 925
rect 400 890 405 925
rect 440 890 445 925
rect 520 890 525 925
rect 560 890 565 925
rect 640 890 645 925
rect 680 890 685 925
rect 760 890 765 925
rect 800 890 805 925
rect 880 890 885 925
rect 920 890 925 925
rect 1000 890 1005 925
rect 1040 890 1045 925
rect 1095 875 1190 925
rect 15 870 45 875
rect 15 775 19 870
rect 15 770 45 775
rect 15 690 110 740
rect 160 705 165 740
rect 200 705 205 740
rect 280 705 285 740
rect 320 705 325 740
rect 400 705 405 740
rect 440 705 445 740
rect 520 705 525 740
rect 560 705 565 740
rect 640 705 645 740
rect 680 705 685 740
rect 760 705 765 740
rect 800 705 805 740
rect 880 705 885 740
rect 920 705 925 740
rect 1000 705 1005 740
rect 1040 705 1045 740
rect 1095 690 1190 740
rect 15 685 45 690
rect 15 590 19 685
rect 15 585 45 590
rect 15 505 110 555
rect 160 520 165 555
rect 200 520 205 555
rect 280 520 285 555
rect 320 520 325 555
rect 400 520 405 555
rect 440 520 445 555
rect 520 520 525 555
rect 560 520 565 555
rect 640 520 645 555
rect 680 520 685 555
rect 760 520 765 555
rect 800 520 805 555
rect 880 520 885 555
rect 920 520 925 555
rect 1000 520 1005 555
rect 1040 520 1045 555
rect 1095 505 1190 555
rect 15 500 45 505
rect 15 405 19 500
rect 15 400 45 405
rect 15 335 45 340
rect 15 240 19 335
rect 15 235 45 240
rect 15 185 110 235
rect 160 185 165 220
rect 200 185 205 220
rect 280 185 285 220
rect 320 185 325 220
rect 400 185 405 220
rect 440 185 445 220
rect 520 185 525 220
rect 560 185 565 220
rect 640 185 645 220
rect 680 185 685 220
rect 760 185 765 220
rect 800 185 805 220
rect 880 185 885 220
rect 920 185 925 220
rect 1000 185 1005 220
rect 1040 185 1045 220
rect 1095 185 1190 235
rect 15 150 45 155
rect 15 55 19 150
rect 15 50 45 55
rect 15 0 110 50
rect 160 0 165 35
rect 200 0 205 35
rect 280 0 285 35
rect 320 0 325 35
rect 400 0 405 35
rect 440 0 445 35
rect 520 0 525 35
rect 560 0 565 35
rect 640 0 645 35
rect 680 0 685 35
rect 760 0 765 35
rect 800 0 805 35
rect 880 0 885 35
rect 920 0 925 35
rect 1000 0 1005 35
rect 1040 0 1045 35
rect 1095 0 1190 50
rect 15 -35 45 -30
rect 15 -130 19 -35
rect 15 -135 45 -130
rect 15 -185 110 -135
rect 160 -185 165 -150
rect 200 -185 205 -150
rect 280 -185 285 -150
rect 320 -185 325 -150
rect 400 -185 405 -150
rect 440 -185 445 -150
rect 520 -185 525 -150
rect 560 -185 565 -150
rect 640 -185 645 -150
rect 680 -185 685 -150
rect 760 -185 765 -150
rect 800 -185 805 -150
rect 880 -185 885 -150
rect 920 -185 925 -150
rect 1000 -185 1005 -150
rect 1040 -185 1045 -150
rect 1095 -185 1190 -135
rect 15 -220 45 -215
rect 15 -315 19 -220
rect 15 -320 45 -315
rect 15 -370 110 -320
rect 160 -370 165 -335
rect 200 -370 205 -335
rect 280 -370 285 -335
rect 320 -370 325 -335
rect 400 -370 405 -335
rect 440 -370 445 -335
rect 520 -370 525 -335
rect 560 -370 565 -335
rect 640 -370 645 -335
rect 680 -370 685 -335
rect 760 -370 765 -335
rect 800 -370 805 -335
rect 880 -370 885 -335
rect 920 -370 925 -335
rect 1000 -370 1005 -335
rect 1040 -370 1045 -335
rect 1095 -370 1190 -320
<< via1 >>
rect 165 1075 200 1110
rect 285 1075 320 1110
rect 405 1075 440 1110
rect 525 1075 560 1110
rect 645 1075 680 1110
rect 765 1075 800 1110
rect 885 1075 920 1110
rect 1005 1075 1040 1110
rect 19 960 45 1055
rect 165 890 200 925
rect 285 890 320 925
rect 405 890 440 925
rect 525 890 560 925
rect 645 890 680 925
rect 765 890 800 925
rect 885 890 920 925
rect 1005 890 1040 925
rect 19 775 45 870
rect 165 705 200 740
rect 285 705 320 740
rect 405 705 440 740
rect 525 705 560 740
rect 645 705 680 740
rect 765 705 800 740
rect 885 705 920 740
rect 1005 705 1040 740
rect 19 590 45 685
rect 165 520 200 555
rect 285 520 320 555
rect 405 520 440 555
rect 525 520 560 555
rect 645 520 680 555
rect 765 520 800 555
rect 885 520 920 555
rect 1005 520 1040 555
rect 19 405 45 500
rect 19 240 45 335
rect 165 185 200 220
rect 285 185 320 220
rect 405 185 440 220
rect 525 185 560 220
rect 645 185 680 220
rect 765 185 800 220
rect 885 185 920 220
rect 1005 185 1040 220
rect 19 55 45 150
rect 165 0 200 35
rect 285 0 320 35
rect 405 0 440 35
rect 525 0 560 35
rect 645 0 680 35
rect 765 0 800 35
rect 885 0 920 35
rect 1005 0 1040 35
rect 19 -130 45 -35
rect 165 -185 200 -150
rect 285 -185 320 -150
rect 405 -185 440 -150
rect 525 -185 560 -150
rect 645 -185 680 -150
rect 765 -185 800 -150
rect 885 -185 920 -150
rect 1005 -185 1040 -150
rect 19 -315 45 -220
rect 165 -370 200 -335
rect 285 -370 320 -335
rect 405 -370 440 -335
rect 525 -370 560 -335
rect 645 -370 680 -335
rect 765 -370 800 -335
rect 885 -370 920 -335
rect 1005 -370 1040 -335
<< metal2 >>
rect 225 1135 980 1185
rect 160 1110 205 1115
rect 225 1110 260 1135
rect 280 1110 325 1115
rect 160 1075 165 1110
rect 200 1075 205 1110
rect 280 1075 285 1110
rect 320 1075 325 1110
rect 400 1110 445 1115
rect 465 1110 500 1135
rect 520 1110 565 1115
rect 400 1075 405 1110
rect 440 1075 445 1110
rect 520 1075 525 1110
rect 560 1075 565 1110
rect 640 1110 685 1115
rect 705 1110 740 1135
rect 760 1110 805 1115
rect 640 1075 645 1110
rect 680 1075 685 1110
rect 760 1075 765 1110
rect 800 1075 805 1110
rect 880 1110 925 1115
rect 945 1110 980 1135
rect 1000 1110 1045 1115
rect 880 1075 885 1110
rect 920 1075 925 1110
rect 1000 1075 1005 1110
rect 1040 1075 1045 1110
rect 15 1055 45 1060
rect 15 960 19 1055
rect 15 870 45 960
rect 160 925 205 930
rect 160 890 165 925
rect 200 890 205 925
rect 280 925 325 930
rect 280 890 285 925
rect 320 890 325 925
rect 400 925 445 930
rect 400 890 405 925
rect 440 890 445 925
rect 520 925 565 930
rect 520 890 525 925
rect 560 890 565 925
rect 640 925 685 930
rect 640 890 645 925
rect 680 890 685 925
rect 760 925 805 930
rect 880 925 925 930
rect 760 890 765 925
rect 800 890 805 925
rect 825 915 860 925
rect 880 890 885 925
rect 920 890 925 925
rect 1000 925 1045 930
rect 1000 890 1005 925
rect 1040 890 1045 925
rect 15 775 19 870
rect 15 685 45 775
rect 160 740 205 745
rect 160 705 165 740
rect 200 705 205 740
rect 280 740 325 745
rect 280 705 285 740
rect 320 705 325 740
rect 400 740 445 745
rect 400 705 405 740
rect 440 705 445 740
rect 520 740 565 745
rect 520 705 525 740
rect 560 705 565 740
rect 640 740 685 745
rect 640 705 645 740
rect 680 705 685 740
rect 760 740 805 745
rect 760 705 765 740
rect 800 705 805 740
rect 880 740 925 745
rect 880 705 885 740
rect 920 705 925 740
rect 1000 740 1045 745
rect 1000 705 1005 740
rect 1040 705 1045 740
rect 15 590 19 685
rect 15 500 45 590
rect 160 555 205 560
rect 160 520 165 555
rect 200 520 205 555
rect 280 555 325 560
rect 280 520 285 555
rect 320 520 325 555
rect 400 555 445 560
rect 400 520 405 555
rect 440 520 445 555
rect 520 555 565 560
rect 520 520 525 555
rect 560 520 565 555
rect 640 555 685 560
rect 640 520 645 555
rect 680 520 685 555
rect 760 555 805 560
rect 760 520 765 555
rect 800 520 805 555
rect 880 555 925 560
rect 880 520 885 555
rect 920 520 925 555
rect 1000 555 1045 560
rect 1000 520 1005 555
rect 1040 520 1045 555
rect 15 405 19 500
rect 15 335 45 405
rect 15 240 19 335
rect 15 150 45 240
rect 160 185 165 220
rect 200 185 205 220
rect 160 180 205 185
rect 280 185 285 220
rect 320 185 325 220
rect 280 180 325 185
rect 400 185 405 220
rect 440 185 445 220
rect 400 180 445 185
rect 520 185 525 220
rect 560 185 565 220
rect 520 180 565 185
rect 640 185 645 220
rect 680 185 685 220
rect 640 180 685 185
rect 760 185 765 220
rect 800 185 805 220
rect 760 180 805 185
rect 880 185 885 220
rect 920 185 925 220
rect 880 180 925 185
rect 1000 185 1005 220
rect 1040 185 1045 220
rect 1000 180 1045 185
rect 15 55 19 150
rect 15 -35 45 55
rect 160 0 165 35
rect 200 0 205 35
rect 160 -5 205 0
rect 280 0 285 35
rect 320 0 325 35
rect 280 -5 325 0
rect 400 0 405 35
rect 440 0 445 35
rect 400 -5 445 0
rect 520 0 525 35
rect 560 0 565 35
rect 520 -5 565 0
rect 640 0 645 35
rect 680 0 685 35
rect 640 -5 685 0
rect 760 0 765 35
rect 800 0 805 35
rect 760 -5 805 0
rect 880 0 885 35
rect 920 0 925 35
rect 880 -5 925 0
rect 1000 0 1005 35
rect 1040 0 1045 35
rect 1000 -5 1045 0
rect 15 -130 19 -35
rect 15 -220 45 -130
rect 160 -185 165 -150
rect 200 -185 205 -150
rect 160 -190 205 -185
rect 280 -185 285 -150
rect 320 -185 325 -150
rect 280 -190 325 -185
rect 400 -185 405 -150
rect 440 -185 445 -150
rect 400 -190 445 -185
rect 520 -185 525 -150
rect 560 -185 565 -150
rect 520 -190 565 -185
rect 640 -185 645 -150
rect 680 -185 685 -150
rect 640 -190 685 -185
rect 760 -185 765 -150
rect 800 -185 805 -150
rect 760 -190 805 -185
rect 880 -185 885 -150
rect 920 -185 925 -150
rect 880 -190 925 -185
rect 1000 -185 1005 -150
rect 1040 -185 1045 -150
rect 1000 -190 1045 -185
rect 15 -315 19 -220
rect 15 -390 45 -315
rect 105 -390 140 -320
rect 160 -370 165 -335
rect 200 -370 205 -335
rect 160 -375 205 -370
rect 280 -370 285 -335
rect 320 -370 325 -335
rect 400 -370 405 -335
rect 440 -370 445 -335
rect 280 -375 325 -370
rect 345 -390 380 -370
rect 400 -375 445 -370
rect 520 -370 525 -335
rect 560 -370 565 -335
rect 640 -370 645 -335
rect 680 -370 685 -335
rect 520 -375 565 -370
rect 585 -390 620 -370
rect 640 -375 685 -370
rect 760 -370 765 -335
rect 800 -370 805 -335
rect 880 -370 885 -335
rect 920 -370 925 -335
rect 760 -375 805 -370
rect 825 -390 860 -370
rect 880 -375 925 -370
rect 1000 -370 1005 -335
rect 1040 -370 1045 -335
rect 1000 -375 1045 -370
rect 1065 -390 1100 -370
rect 1160 -390 1190 1060
rect 15 -440 1190 -390
<< via2 >>
rect 165 1080 200 1110
rect 285 1080 320 1110
rect 405 1080 440 1110
rect 525 1080 560 1110
rect 645 1080 680 1110
rect 765 1080 800 1110
rect 885 1080 920 1110
rect 1005 1080 1040 1110
rect 165 895 200 925
rect 285 895 320 925
rect 405 895 440 925
rect 525 895 560 925
rect 645 895 680 925
rect 765 895 800 925
rect 885 895 920 925
rect 1005 895 1040 925
rect 165 710 200 740
rect 285 710 320 740
rect 405 710 440 740
rect 525 710 560 740
rect 645 710 680 740
rect 765 710 800 740
rect 885 710 920 740
rect 1005 710 1040 740
rect 165 525 200 555
rect 285 525 320 555
rect 405 525 440 555
rect 525 525 560 555
rect 645 525 680 555
rect 765 525 800 555
rect 885 525 920 555
rect 1005 525 1040 555
rect 165 185 200 215
rect 285 185 320 215
rect 405 185 440 215
rect 525 185 560 215
rect 645 185 680 215
rect 765 185 800 215
rect 885 185 920 215
rect 1005 185 1040 215
rect 165 0 200 30
rect 285 0 320 30
rect 405 0 440 30
rect 525 0 560 30
rect 645 0 680 30
rect 765 0 800 30
rect 885 0 920 30
rect 1005 0 1040 30
rect 165 -185 200 -155
rect 285 -185 320 -155
rect 405 -185 440 -155
rect 525 -185 560 -155
rect 645 -185 680 -155
rect 765 -185 800 -155
rect 885 -185 920 -155
rect 1005 -185 1040 -155
rect 165 -370 200 -340
rect 285 -370 320 -340
rect 405 -370 440 -340
rect 525 -370 560 -340
rect 645 -370 680 -340
rect 765 -370 800 -340
rect 885 -370 920 -340
rect 1005 -370 1040 -340
<< metal3 >>
rect 160 1110 1165 1115
rect 160 1080 165 1110
rect 200 1080 285 1110
rect 320 1080 405 1110
rect 440 1080 525 1110
rect 560 1080 645 1110
rect 680 1080 765 1110
rect 800 1080 885 1110
rect 920 1080 1005 1110
rect 1040 1080 1165 1110
rect 160 1075 1165 1080
rect 1120 930 1165 1075
rect 1200 940 1280 945
rect 1200 930 1210 940
rect 160 925 1210 930
rect 160 895 165 925
rect 200 895 285 925
rect 320 895 405 925
rect 440 895 525 925
rect 560 895 645 925
rect 680 895 765 925
rect 800 895 885 925
rect 920 895 1005 925
rect 1040 895 1210 925
rect 160 890 1210 895
rect 1200 880 1210 890
rect 1275 880 1280 940
rect 1200 875 1280 880
rect 1100 755 1175 760
rect 1100 745 1105 755
rect 160 740 1105 745
rect 160 710 165 740
rect 200 710 285 740
rect 320 710 405 740
rect 440 710 525 740
rect 560 710 645 740
rect 680 710 765 740
rect 800 710 885 740
rect 920 710 1005 740
rect 1040 710 1105 740
rect 160 705 1105 710
rect 1100 695 1105 705
rect 1170 745 1175 755
rect 1170 705 1295 745
rect 1170 695 1175 705
rect 1100 690 1175 695
rect 280 615 925 655
rect 280 560 325 615
rect 880 560 925 615
rect 995 625 1070 630
rect 995 565 1000 625
rect 1065 565 1070 625
rect 995 560 1070 565
rect 160 555 325 560
rect 160 525 165 555
rect 200 525 285 555
rect 320 525 325 555
rect 160 520 325 525
rect 400 555 805 560
rect 400 525 405 555
rect 440 525 525 555
rect 560 525 645 555
rect 680 525 765 555
rect 800 525 805 555
rect 400 520 805 525
rect 880 555 1295 560
rect 880 525 885 555
rect 920 525 1005 555
rect 1040 525 1295 555
rect 880 520 1295 525
rect 760 490 805 520
rect 760 455 1295 490
rect 520 390 1295 425
rect 520 220 565 390
rect 160 215 325 220
rect 160 185 165 215
rect 200 185 285 215
rect 320 185 325 215
rect 160 180 325 185
rect 400 215 565 220
rect 400 185 405 215
rect 440 185 525 215
rect 560 185 565 215
rect 400 180 565 185
rect 640 325 1295 360
rect 640 215 685 325
rect 640 185 645 215
rect 680 185 685 215
rect 640 180 685 185
rect 760 255 1295 290
rect 760 215 805 255
rect 760 185 765 215
rect 800 185 805 215
rect 760 180 805 185
rect 880 215 1070 220
rect 880 185 885 215
rect 920 185 1005 215
rect 1040 185 1070 215
rect 880 180 1070 185
rect 280 125 325 180
rect 880 125 925 180
rect 280 85 925 125
rect 995 175 1070 180
rect 995 115 1000 175
rect 1065 115 1070 175
rect 995 110 1070 115
rect 1100 45 1175 50
rect 1100 35 1105 45
rect 160 30 1105 35
rect 160 0 165 30
rect 200 0 285 30
rect 320 0 405 30
rect 440 0 525 30
rect 560 0 645 30
rect 680 0 765 30
rect 800 0 885 30
rect 920 0 1005 30
rect 1040 0 1105 30
rect 160 -5 1105 0
rect 1100 -15 1105 -5
rect 1170 -15 1175 45
rect 1100 -20 1175 -15
rect 1205 -140 1280 -135
rect 1205 -150 1210 -140
rect 160 -155 1210 -150
rect 160 -185 165 -155
rect 200 -185 285 -155
rect 320 -185 405 -155
rect 440 -185 525 -155
rect 560 -185 645 -155
rect 680 -185 765 -155
rect 800 -185 885 -155
rect 920 -185 1005 -155
rect 1040 -185 1210 -155
rect 160 -190 1210 -185
rect 1120 -335 1165 -190
rect 1205 -200 1210 -190
rect 1275 -200 1280 -140
rect 1205 -205 1280 -200
rect 160 -340 1165 -335
rect 160 -370 165 -340
rect 200 -370 285 -340
rect 320 -370 405 -340
rect 440 -370 525 -340
rect 560 -370 645 -340
rect 680 -370 765 -340
rect 800 -370 885 -340
rect 920 -370 1005 -340
rect 1040 -370 1165 -340
rect 160 -375 1165 -370
<< via3 >>
rect 1210 880 1275 940
rect 1105 695 1170 755
rect 1000 565 1065 625
rect 1000 115 1065 175
rect 1105 -15 1170 45
rect 1210 -200 1275 -140
<< metal4 >>
rect 1205 940 1280 945
rect 1205 880 1210 940
rect 1275 880 1280 940
rect 1100 755 1175 760
rect 1100 695 1105 755
rect 1170 695 1175 755
rect 995 625 1070 630
rect 995 565 1000 625
rect 1065 565 1070 625
rect 995 175 1070 565
rect 995 115 1000 175
rect 1065 115 1070 175
rect 995 110 1070 115
rect 1100 45 1175 695
rect 1100 -15 1105 45
rect 1170 -15 1175 45
rect 1100 -20 1175 -15
rect 1205 -140 1280 880
rect 1205 -200 1210 -140
rect 1275 -200 1280 -140
rect 1205 -205 1280 -200
use pmirror_pfet_8xSlice  pmirror_pfet_8xSlice_0
timestamp 1659898741
transform 1 0 0 0 1 370
box 0 -740 244 740
use pmirror_pfet_8xSlice  pmirror_pfet_8xSlice_1
timestamp 1659898741
transform 1 0 120 0 1 370
box 0 -740 244 740
use pmirror_pfet_8xSlice  pmirror_pfet_8xSlice_2
timestamp 1659898741
transform 1 0 240 0 1 370
box 0 -740 244 740
use pmirror_pfet_8xSlice  pmirror_pfet_8xSlice_3
timestamp 1659898741
transform 1 0 360 0 1 370
box 0 -740 244 740
use pmirror_pfet_8xSlice  pmirror_pfet_8xSlice_4
timestamp 1659898741
transform 1 0 480 0 1 370
box 0 -740 244 740
use pmirror_pfet_8xSlice  pmirror_pfet_8xSlice_5
timestamp 1659898741
transform 1 0 600 0 1 370
box 0 -740 244 740
use pmirror_pfet_8xSlice  pmirror_pfet_8xSlice_6
timestamp 1659898741
transform 1 0 720 0 1 370
box 0 -740 244 740
use pmirror_pfet_8xSlice  pmirror_pfet_8xSlice_7
timestamp 1659898741
transform 1 0 840 0 1 370
box 0 -740 244 740
use pmirror_pfet_8xSlice  pmirror_pfet_8xSlice_8
timestamp 1659898741
transform 1 0 960 0 1 370
box 0 -740 244 740
<< end >>
