magic
tech sky130B
timestamp 1662014484
<< metal1 >>
rect 7000 80950 29000 81000
rect 7000 80940 7060 80950
rect 7190 80940 7310 80950
rect 7440 80940 7560 80950
rect 7690 80940 7810 80950
rect 7940 80940 8060 80950
rect 8190 80940 8310 80950
rect 8440 80940 8560 80950
rect 8690 80940 8810 80950
rect 8940 80940 9060 80950
rect 9190 80940 9310 80950
rect 9440 80940 9560 80950
rect 9690 80940 9810 80950
rect 9940 80940 10060 80950
rect 10190 80940 10310 80950
rect 10440 80940 10560 80950
rect 10690 80940 10810 80950
rect 10940 80940 11060 80950
rect 11190 80940 11310 80950
rect 11440 80940 11560 80950
rect 11690 80940 11810 80950
rect 11940 80940 12060 80950
rect 12190 80940 12310 80950
rect 12440 80940 12560 80950
rect 12690 80940 12810 80950
rect 12940 80940 13060 80950
rect 13190 80940 13310 80950
rect 13440 80940 13560 80950
rect 13690 80940 13810 80950
rect 13940 80940 14060 80950
rect 14190 80940 14310 80950
rect 14440 80940 14560 80950
rect 14690 80940 14810 80950
rect 14940 80940 15060 80950
rect 15190 80940 15310 80950
rect 15440 80940 15560 80950
rect 15690 80940 15810 80950
rect 15940 80940 16060 80950
rect 16190 80940 16310 80950
rect 16440 80940 16560 80950
rect 16690 80940 16810 80950
rect 16940 80940 17060 80950
rect 17190 80940 17310 80950
rect 17440 80940 17560 80950
rect 17690 80940 17810 80950
rect 17940 80940 18060 80950
rect 18190 80940 18310 80950
rect 18440 80940 18560 80950
rect 18690 80940 18810 80950
rect 18940 80940 19060 80950
rect 19190 80940 19310 80950
rect 19440 80940 19560 80950
rect 19690 80940 19810 80950
rect 19940 80940 20060 80950
rect 20190 80940 20310 80950
rect 20440 80940 20560 80950
rect 20690 80940 20810 80950
rect 20940 80940 21060 80950
rect 21190 80940 21310 80950
rect 21440 80940 21560 80950
rect 21690 80940 21810 80950
rect 21940 80940 22060 80950
rect 22190 80940 22310 80950
rect 22440 80940 22560 80950
rect 22690 80940 22810 80950
rect 22940 80940 23060 80950
rect 23190 80940 23310 80950
rect 23440 80940 23560 80950
rect 23690 80940 23810 80950
rect 23940 80940 24060 80950
rect 24190 80940 24310 80950
rect 24440 80940 24560 80950
rect 24690 80940 24810 80950
rect 24940 80940 25060 80950
rect 25190 80940 25310 80950
rect 25440 80940 25560 80950
rect 25690 80940 25810 80950
rect 25940 80940 26060 80950
rect 26190 80940 26310 80950
rect 26440 80940 26560 80950
rect 26690 80940 26810 80950
rect 26940 80940 27060 80950
rect 27190 80940 27310 80950
rect 27440 80940 27560 80950
rect 27690 80940 27810 80950
rect 27940 80940 28060 80950
rect 28190 80940 28310 80950
rect 28440 80940 28560 80950
rect 28690 80940 28810 80950
rect 28940 80940 29000 80950
rect 7000 80810 7050 80940
rect 7200 80810 7300 80940
rect 7450 80810 7550 80940
rect 7700 80810 7800 80940
rect 7950 80810 8050 80940
rect 8200 80810 8300 80940
rect 8450 80810 8550 80940
rect 8700 80810 8800 80940
rect 8950 80810 9050 80940
rect 9200 80810 9300 80940
rect 9450 80810 9550 80940
rect 9700 80810 9800 80940
rect 9950 80810 10050 80940
rect 10200 80810 10300 80940
rect 10450 80810 10550 80940
rect 10700 80810 10800 80940
rect 10950 80810 11050 80940
rect 11200 80810 11300 80940
rect 11450 80810 11550 80940
rect 11700 80810 11800 80940
rect 11950 80810 12050 80940
rect 12200 80810 12300 80940
rect 12450 80810 12550 80940
rect 12700 80810 12800 80940
rect 12950 80810 13050 80940
rect 13200 80810 13300 80940
rect 13450 80810 13550 80940
rect 13700 80810 13800 80940
rect 13950 80810 14050 80940
rect 14200 80810 14300 80940
rect 14450 80810 14550 80940
rect 14700 80810 14800 80940
rect 14950 80810 15050 80940
rect 15200 80810 15300 80940
rect 15450 80810 15550 80940
rect 15700 80810 15800 80940
rect 15950 80810 16050 80940
rect 16200 80810 16300 80940
rect 16450 80810 16550 80940
rect 16700 80810 16800 80940
rect 16950 80810 17050 80940
rect 17200 80810 17300 80940
rect 17450 80810 17550 80940
rect 17700 80810 17800 80940
rect 17950 80810 18050 80940
rect 18200 80810 18300 80940
rect 18450 80810 18550 80940
rect 18700 80810 18800 80940
rect 18950 80810 19050 80940
rect 19200 80810 19300 80940
rect 19450 80810 19550 80940
rect 19700 80810 19800 80940
rect 19950 80810 20050 80940
rect 20200 80810 20300 80940
rect 20450 80810 20550 80940
rect 20700 80810 20800 80940
rect 20950 80810 21050 80940
rect 21200 80810 21300 80940
rect 21450 80810 21550 80940
rect 21700 80810 21800 80940
rect 21950 80810 22050 80940
rect 22200 80810 22300 80940
rect 22450 80810 22550 80940
rect 22700 80810 22800 80940
rect 22950 80810 23050 80940
rect 23200 80810 23300 80940
rect 23450 80810 23550 80940
rect 23700 80810 23800 80940
rect 23950 80810 24050 80940
rect 24200 80810 24300 80940
rect 24450 80810 24550 80940
rect 24700 80810 24800 80940
rect 24950 80810 25050 80940
rect 25200 80810 25300 80940
rect 25450 80810 25550 80940
rect 25700 80810 25800 80940
rect 25950 80810 26050 80940
rect 26200 80810 26300 80940
rect 26450 80810 26550 80940
rect 26700 80810 26800 80940
rect 26950 80810 27050 80940
rect 27200 80810 27300 80940
rect 27450 80810 27550 80940
rect 27700 80810 27800 80940
rect 27950 80810 28050 80940
rect 28200 80810 28300 80940
rect 28450 80810 28550 80940
rect 28700 80810 28800 80940
rect 28950 80810 29000 80940
rect 7000 80800 7060 80810
rect 7190 80800 7310 80810
rect 7440 80800 7560 80810
rect 7690 80800 7810 80810
rect 7940 80800 8060 80810
rect 8190 80800 8310 80810
rect 8440 80800 8560 80810
rect 8690 80800 8810 80810
rect 8940 80800 9060 80810
rect 9190 80800 9310 80810
rect 9440 80800 9560 80810
rect 9690 80800 9810 80810
rect 9940 80800 10060 80810
rect 10190 80800 10310 80810
rect 10440 80800 10560 80810
rect 10690 80800 10810 80810
rect 10940 80800 11060 80810
rect 11190 80800 11310 80810
rect 11440 80800 11560 80810
rect 11690 80800 11810 80810
rect 11940 80800 12060 80810
rect 12190 80800 12310 80810
rect 12440 80800 12560 80810
rect 12690 80800 12810 80810
rect 12940 80800 13060 80810
rect 13190 80800 13310 80810
rect 13440 80800 13560 80810
rect 13690 80800 13810 80810
rect 13940 80800 14060 80810
rect 14190 80800 14310 80810
rect 14440 80800 14560 80810
rect 14690 80800 14810 80810
rect 14940 80800 15060 80810
rect 15190 80800 15310 80810
rect 15440 80800 15560 80810
rect 15690 80800 15810 80810
rect 15940 80800 16060 80810
rect 16190 80800 16310 80810
rect 16440 80800 16560 80810
rect 16690 80800 16810 80810
rect 16940 80800 17060 80810
rect 17190 80800 17310 80810
rect 17440 80800 17560 80810
rect 17690 80800 17810 80810
rect 17940 80800 18060 80810
rect 18190 80800 18310 80810
rect 18440 80800 18560 80810
rect 18690 80800 18810 80810
rect 18940 80800 19060 80810
rect 19190 80800 19310 80810
rect 19440 80800 19560 80810
rect 19690 80800 19810 80810
rect 19940 80800 20060 80810
rect 20190 80800 20310 80810
rect 20440 80800 20560 80810
rect 20690 80800 20810 80810
rect 20940 80800 21060 80810
rect 21190 80800 21310 80810
rect 21440 80800 21560 80810
rect 21690 80800 21810 80810
rect 21940 80800 22060 80810
rect 22190 80800 22310 80810
rect 22440 80800 22560 80810
rect 22690 80800 22810 80810
rect 22940 80800 23060 80810
rect 23190 80800 23310 80810
rect 23440 80800 23560 80810
rect 23690 80800 23810 80810
rect 23940 80800 24060 80810
rect 24190 80800 24310 80810
rect 24440 80800 24560 80810
rect 24690 80800 24810 80810
rect 24940 80800 25060 80810
rect 25190 80800 25310 80810
rect 25440 80800 25560 80810
rect 25690 80800 25810 80810
rect 25940 80800 26060 80810
rect 26190 80800 26310 80810
rect 26440 80800 26560 80810
rect 26690 80800 26810 80810
rect 26940 80800 27060 80810
rect 27190 80800 27310 80810
rect 27440 80800 27560 80810
rect 27690 80800 27810 80810
rect 27940 80800 28060 80810
rect 28190 80800 28310 80810
rect 28440 80800 28560 80810
rect 28690 80800 28810 80810
rect 28940 80800 29000 80810
rect 7000 80700 29000 80800
rect 7000 80690 7060 80700
rect 7190 80690 7310 80700
rect 7440 80690 7560 80700
rect 7690 80690 7810 80700
rect 7940 80690 8060 80700
rect 8190 80690 8310 80700
rect 8440 80690 8560 80700
rect 8690 80690 8810 80700
rect 8940 80690 9060 80700
rect 9190 80690 9310 80700
rect 9440 80690 9560 80700
rect 9690 80690 9810 80700
rect 9940 80690 10060 80700
rect 10190 80690 10310 80700
rect 10440 80690 10560 80700
rect 10690 80690 10810 80700
rect 10940 80690 11060 80700
rect 11190 80690 11310 80700
rect 11440 80690 11560 80700
rect 11690 80690 11810 80700
rect 11940 80690 12060 80700
rect 12190 80690 12310 80700
rect 12440 80690 12560 80700
rect 12690 80690 12810 80700
rect 12940 80690 13060 80700
rect 13190 80690 13310 80700
rect 13440 80690 13560 80700
rect 13690 80690 13810 80700
rect 13940 80690 14060 80700
rect 14190 80690 14310 80700
rect 14440 80690 14560 80700
rect 14690 80690 14810 80700
rect 14940 80690 15060 80700
rect 15190 80690 15310 80700
rect 15440 80690 15560 80700
rect 15690 80690 15810 80700
rect 15940 80690 16060 80700
rect 16190 80690 16310 80700
rect 16440 80690 16560 80700
rect 16690 80690 16810 80700
rect 16940 80690 17060 80700
rect 17190 80690 17310 80700
rect 17440 80690 17560 80700
rect 17690 80690 17810 80700
rect 17940 80690 18060 80700
rect 18190 80690 18310 80700
rect 18440 80690 18560 80700
rect 18690 80690 18810 80700
rect 18940 80690 19060 80700
rect 19190 80690 19310 80700
rect 19440 80690 19560 80700
rect 19690 80690 19810 80700
rect 19940 80690 20060 80700
rect 20190 80690 20310 80700
rect 20440 80690 20560 80700
rect 20690 80690 20810 80700
rect 20940 80690 21060 80700
rect 21190 80690 21310 80700
rect 21440 80690 21560 80700
rect 21690 80690 21810 80700
rect 21940 80690 22060 80700
rect 22190 80690 22310 80700
rect 22440 80690 22560 80700
rect 22690 80690 22810 80700
rect 22940 80690 23060 80700
rect 23190 80690 23310 80700
rect 23440 80690 23560 80700
rect 23690 80690 23810 80700
rect 23940 80690 24060 80700
rect 24190 80690 24310 80700
rect 24440 80690 24560 80700
rect 24690 80690 24810 80700
rect 24940 80690 25060 80700
rect 25190 80690 25310 80700
rect 25440 80690 25560 80700
rect 25690 80690 25810 80700
rect 25940 80690 26060 80700
rect 26190 80690 26310 80700
rect 26440 80690 26560 80700
rect 26690 80690 26810 80700
rect 26940 80690 27060 80700
rect 27190 80690 27310 80700
rect 27440 80690 27560 80700
rect 27690 80690 27810 80700
rect 27940 80690 28060 80700
rect 28190 80690 28310 80700
rect 28440 80690 28560 80700
rect 28690 80690 28810 80700
rect 28940 80690 29000 80700
rect 7000 80560 7050 80690
rect 7200 80560 7300 80690
rect 7450 80560 7550 80690
rect 7700 80560 7800 80690
rect 7950 80560 8050 80690
rect 8200 80560 8300 80690
rect 8450 80560 8550 80690
rect 8700 80560 8800 80690
rect 8950 80560 9050 80690
rect 9200 80560 9300 80690
rect 9450 80560 9550 80690
rect 9700 80560 9800 80690
rect 9950 80560 10050 80690
rect 10200 80560 10300 80690
rect 10450 80560 10550 80690
rect 10700 80560 10800 80690
rect 10950 80560 11050 80690
rect 11200 80560 11300 80690
rect 11450 80560 11550 80690
rect 11700 80560 11800 80690
rect 11950 80560 12050 80690
rect 12200 80560 12300 80690
rect 12450 80560 12550 80690
rect 12700 80560 12800 80690
rect 12950 80560 13050 80690
rect 13200 80560 13300 80690
rect 13450 80560 13550 80690
rect 13700 80560 13800 80690
rect 13950 80560 14050 80690
rect 14200 80560 14300 80690
rect 14450 80560 14550 80690
rect 14700 80560 14800 80690
rect 14950 80560 15050 80690
rect 15200 80560 15300 80690
rect 15450 80560 15550 80690
rect 15700 80560 15800 80690
rect 15950 80560 16050 80690
rect 16200 80560 16300 80690
rect 16450 80560 16550 80690
rect 16700 80560 16800 80690
rect 16950 80560 17050 80690
rect 17200 80560 17300 80690
rect 17450 80560 17550 80690
rect 17700 80560 17800 80690
rect 17950 80560 18050 80690
rect 18200 80560 18300 80690
rect 18450 80560 18550 80690
rect 18700 80560 18800 80690
rect 18950 80560 19050 80690
rect 19200 80560 19300 80690
rect 19450 80560 19550 80690
rect 19700 80560 19800 80690
rect 19950 80560 20050 80690
rect 20200 80560 20300 80690
rect 20450 80560 20550 80690
rect 20700 80560 20800 80690
rect 20950 80560 21050 80690
rect 21200 80560 21300 80690
rect 21450 80560 21550 80690
rect 21700 80560 21800 80690
rect 21950 80560 22050 80690
rect 22200 80560 22300 80690
rect 22450 80560 22550 80690
rect 22700 80560 22800 80690
rect 22950 80560 23050 80690
rect 23200 80560 23300 80690
rect 23450 80560 23550 80690
rect 23700 80560 23800 80690
rect 23950 80560 24050 80690
rect 24200 80560 24300 80690
rect 24450 80560 24550 80690
rect 24700 80560 24800 80690
rect 24950 80560 25050 80690
rect 25200 80560 25300 80690
rect 25450 80560 25550 80690
rect 25700 80560 25800 80690
rect 25950 80560 26050 80690
rect 26200 80560 26300 80690
rect 26450 80560 26550 80690
rect 26700 80560 26800 80690
rect 26950 80560 27050 80690
rect 27200 80560 27300 80690
rect 27450 80560 27550 80690
rect 27700 80560 27800 80690
rect 27950 80560 28050 80690
rect 28200 80560 28300 80690
rect 28450 80560 28550 80690
rect 28700 80560 28800 80690
rect 28950 80560 29000 80690
rect 7000 80550 7060 80560
rect 7190 80550 7310 80560
rect 7440 80550 7560 80560
rect 7690 80550 7810 80560
rect 7940 80550 8060 80560
rect 8190 80550 8310 80560
rect 8440 80550 8560 80560
rect 8690 80550 8810 80560
rect 8940 80550 9060 80560
rect 9190 80550 9310 80560
rect 9440 80550 9560 80560
rect 9690 80550 9810 80560
rect 9940 80550 10060 80560
rect 10190 80550 10310 80560
rect 10440 80550 10560 80560
rect 10690 80550 10810 80560
rect 10940 80550 11060 80560
rect 11190 80550 11310 80560
rect 11440 80550 11560 80560
rect 11690 80550 11810 80560
rect 11940 80550 12060 80560
rect 12190 80550 12310 80560
rect 12440 80550 12560 80560
rect 12690 80550 12810 80560
rect 12940 80550 13060 80560
rect 13190 80550 13310 80560
rect 13440 80550 13560 80560
rect 13690 80550 13810 80560
rect 13940 80550 14060 80560
rect 14190 80550 14310 80560
rect 14440 80550 14560 80560
rect 14690 80550 14810 80560
rect 14940 80550 15060 80560
rect 15190 80550 15310 80560
rect 15440 80550 15560 80560
rect 15690 80550 15810 80560
rect 15940 80550 16060 80560
rect 16190 80550 16310 80560
rect 16440 80550 16560 80560
rect 16690 80550 16810 80560
rect 16940 80550 17060 80560
rect 17190 80550 17310 80560
rect 17440 80550 17560 80560
rect 17690 80550 17810 80560
rect 17940 80550 18060 80560
rect 18190 80550 18310 80560
rect 18440 80550 18560 80560
rect 18690 80550 18810 80560
rect 18940 80550 19060 80560
rect 19190 80550 19310 80560
rect 19440 80550 19560 80560
rect 19690 80550 19810 80560
rect 19940 80550 20060 80560
rect 20190 80550 20310 80560
rect 20440 80550 20560 80560
rect 20690 80550 20810 80560
rect 20940 80550 21060 80560
rect 21190 80550 21310 80560
rect 21440 80550 21560 80560
rect 21690 80550 21810 80560
rect 21940 80550 22060 80560
rect 22190 80550 22310 80560
rect 22440 80550 22560 80560
rect 22690 80550 22810 80560
rect 22940 80550 23060 80560
rect 23190 80550 23310 80560
rect 23440 80550 23560 80560
rect 23690 80550 23810 80560
rect 23940 80550 24060 80560
rect 24190 80550 24310 80560
rect 24440 80550 24560 80560
rect 24690 80550 24810 80560
rect 24940 80550 25060 80560
rect 25190 80550 25310 80560
rect 25440 80550 25560 80560
rect 25690 80550 25810 80560
rect 25940 80550 26060 80560
rect 26190 80550 26310 80560
rect 26440 80550 26560 80560
rect 26690 80550 26810 80560
rect 26940 80550 27060 80560
rect 27190 80550 27310 80560
rect 27440 80550 27560 80560
rect 27690 80550 27810 80560
rect 27940 80550 28060 80560
rect 28190 80550 28310 80560
rect 28440 80550 28560 80560
rect 28690 80550 28810 80560
rect 28940 80550 29000 80560
rect 7000 80450 29000 80550
rect 7000 80440 7060 80450
rect 7190 80440 7310 80450
rect 7440 80440 7560 80450
rect 7690 80440 7810 80450
rect 7940 80440 8060 80450
rect 8190 80440 8310 80450
rect 8440 80440 8560 80450
rect 8690 80440 8810 80450
rect 8940 80440 9060 80450
rect 9190 80440 9310 80450
rect 9440 80440 9560 80450
rect 9690 80440 9810 80450
rect 9940 80440 10060 80450
rect 10190 80440 10310 80450
rect 10440 80440 10560 80450
rect 10690 80440 10810 80450
rect 10940 80440 11060 80450
rect 11190 80440 11310 80450
rect 11440 80440 11560 80450
rect 11690 80440 11810 80450
rect 11940 80440 12060 80450
rect 12190 80440 12310 80450
rect 12440 80440 12560 80450
rect 12690 80440 12810 80450
rect 12940 80440 13060 80450
rect 13190 80440 13310 80450
rect 13440 80440 13560 80450
rect 13690 80440 13810 80450
rect 13940 80440 14060 80450
rect 14190 80440 14310 80450
rect 14440 80440 14560 80450
rect 14690 80440 14810 80450
rect 14940 80440 15060 80450
rect 15190 80440 15310 80450
rect 15440 80440 15560 80450
rect 15690 80440 15810 80450
rect 15940 80440 16060 80450
rect 16190 80440 16310 80450
rect 16440 80440 16560 80450
rect 16690 80440 16810 80450
rect 16940 80440 17060 80450
rect 17190 80440 17310 80450
rect 17440 80440 17560 80450
rect 17690 80440 17810 80450
rect 17940 80440 18060 80450
rect 18190 80440 18310 80450
rect 18440 80440 18560 80450
rect 18690 80440 18810 80450
rect 18940 80440 19060 80450
rect 19190 80440 19310 80450
rect 19440 80440 19560 80450
rect 19690 80440 19810 80450
rect 19940 80440 20060 80450
rect 20190 80440 20310 80450
rect 20440 80440 20560 80450
rect 20690 80440 20810 80450
rect 20940 80440 21060 80450
rect 21190 80440 21310 80450
rect 21440 80440 21560 80450
rect 21690 80440 21810 80450
rect 21940 80440 22060 80450
rect 22190 80440 22310 80450
rect 22440 80440 22560 80450
rect 22690 80440 22810 80450
rect 22940 80440 23060 80450
rect 23190 80440 23310 80450
rect 23440 80440 23560 80450
rect 23690 80440 23810 80450
rect 23940 80440 24060 80450
rect 24190 80440 24310 80450
rect 24440 80440 24560 80450
rect 24690 80440 24810 80450
rect 24940 80440 25060 80450
rect 25190 80440 25310 80450
rect 25440 80440 25560 80450
rect 25690 80440 25810 80450
rect 25940 80440 26060 80450
rect 26190 80440 26310 80450
rect 26440 80440 26560 80450
rect 26690 80440 26810 80450
rect 26940 80440 27060 80450
rect 27190 80440 27310 80450
rect 27440 80440 27560 80450
rect 27690 80440 27810 80450
rect 27940 80440 28060 80450
rect 28190 80440 28310 80450
rect 28440 80440 28560 80450
rect 28690 80440 28810 80450
rect 28940 80440 29000 80450
rect 7000 80310 7050 80440
rect 7200 80310 7300 80440
rect 7450 80310 7550 80440
rect 7700 80310 7800 80440
rect 7950 80310 8050 80440
rect 8200 80310 8300 80440
rect 8450 80310 8550 80440
rect 8700 80310 8800 80440
rect 8950 80310 9050 80440
rect 9200 80310 9300 80440
rect 9450 80310 9550 80440
rect 9700 80310 9800 80440
rect 9950 80310 10050 80440
rect 10200 80310 10300 80440
rect 10450 80310 10550 80440
rect 10700 80310 10800 80440
rect 10950 80310 11050 80440
rect 11200 80310 11300 80440
rect 11450 80310 11550 80440
rect 11700 80310 11800 80440
rect 11950 80310 12050 80440
rect 12200 80310 12300 80440
rect 12450 80310 12550 80440
rect 12700 80310 12800 80440
rect 12950 80310 13050 80440
rect 13200 80310 13300 80440
rect 13450 80310 13550 80440
rect 13700 80310 13800 80440
rect 13950 80310 14050 80440
rect 14200 80310 14300 80440
rect 14450 80310 14550 80440
rect 14700 80310 14800 80440
rect 14950 80310 15050 80440
rect 15200 80310 15300 80440
rect 15450 80310 15550 80440
rect 15700 80310 15800 80440
rect 15950 80310 16050 80440
rect 16200 80310 16300 80440
rect 16450 80310 16550 80440
rect 16700 80310 16800 80440
rect 16950 80310 17050 80440
rect 17200 80310 17300 80440
rect 17450 80310 17550 80440
rect 17700 80310 17800 80440
rect 17950 80310 18050 80440
rect 18200 80310 18300 80440
rect 18450 80310 18550 80440
rect 18700 80310 18800 80440
rect 18950 80310 19050 80440
rect 19200 80310 19300 80440
rect 19450 80310 19550 80440
rect 19700 80310 19800 80440
rect 19950 80310 20050 80440
rect 20200 80310 20300 80440
rect 20450 80310 20550 80440
rect 20700 80310 20800 80440
rect 20950 80310 21050 80440
rect 21200 80310 21300 80440
rect 21450 80310 21550 80440
rect 21700 80310 21800 80440
rect 21950 80310 22050 80440
rect 22200 80310 22300 80440
rect 22450 80310 22550 80440
rect 22700 80310 22800 80440
rect 22950 80310 23050 80440
rect 23200 80310 23300 80440
rect 23450 80310 23550 80440
rect 23700 80310 23800 80440
rect 23950 80310 24050 80440
rect 24200 80310 24300 80440
rect 24450 80310 24550 80440
rect 24700 80310 24800 80440
rect 24950 80310 25050 80440
rect 25200 80310 25300 80440
rect 25450 80310 25550 80440
rect 25700 80310 25800 80440
rect 25950 80310 26050 80440
rect 26200 80310 26300 80440
rect 26450 80310 26550 80440
rect 26700 80310 26800 80440
rect 26950 80310 27050 80440
rect 27200 80310 27300 80440
rect 27450 80310 27550 80440
rect 27700 80310 27800 80440
rect 27950 80310 28050 80440
rect 28200 80310 28300 80440
rect 28450 80310 28550 80440
rect 28700 80310 28800 80440
rect 28950 80310 29000 80440
rect 7000 80300 7060 80310
rect 7190 80300 7310 80310
rect 7440 80300 7560 80310
rect 7690 80300 7810 80310
rect 7940 80300 8060 80310
rect 8190 80300 8310 80310
rect 8440 80300 8560 80310
rect 8690 80300 8810 80310
rect 8940 80300 9060 80310
rect 9190 80300 9310 80310
rect 9440 80300 9560 80310
rect 9690 80300 9810 80310
rect 9940 80300 10060 80310
rect 10190 80300 10310 80310
rect 10440 80300 10560 80310
rect 10690 80300 10810 80310
rect 10940 80300 11060 80310
rect 11190 80300 11310 80310
rect 11440 80300 11560 80310
rect 11690 80300 11810 80310
rect 11940 80300 12060 80310
rect 12190 80300 12310 80310
rect 12440 80300 12560 80310
rect 12690 80300 12810 80310
rect 12940 80300 13060 80310
rect 13190 80300 13310 80310
rect 13440 80300 13560 80310
rect 13690 80300 13810 80310
rect 13940 80300 14060 80310
rect 14190 80300 14310 80310
rect 14440 80300 14560 80310
rect 14690 80300 14810 80310
rect 14940 80300 15060 80310
rect 15190 80300 15310 80310
rect 15440 80300 15560 80310
rect 15690 80300 15810 80310
rect 15940 80300 16060 80310
rect 16190 80300 16310 80310
rect 16440 80300 16560 80310
rect 16690 80300 16810 80310
rect 16940 80300 17060 80310
rect 17190 80300 17310 80310
rect 17440 80300 17560 80310
rect 17690 80300 17810 80310
rect 17940 80300 18060 80310
rect 18190 80300 18310 80310
rect 18440 80300 18560 80310
rect 18690 80300 18810 80310
rect 18940 80300 19060 80310
rect 19190 80300 19310 80310
rect 19440 80300 19560 80310
rect 19690 80300 19810 80310
rect 19940 80300 20060 80310
rect 20190 80300 20310 80310
rect 20440 80300 20560 80310
rect 20690 80300 20810 80310
rect 20940 80300 21060 80310
rect 21190 80300 21310 80310
rect 21440 80300 21560 80310
rect 21690 80300 21810 80310
rect 21940 80300 22060 80310
rect 22190 80300 22310 80310
rect 22440 80300 22560 80310
rect 22690 80300 22810 80310
rect 22940 80300 23060 80310
rect 23190 80300 23310 80310
rect 23440 80300 23560 80310
rect 23690 80300 23810 80310
rect 23940 80300 24060 80310
rect 24190 80300 24310 80310
rect 24440 80300 24560 80310
rect 24690 80300 24810 80310
rect 24940 80300 25060 80310
rect 25190 80300 25310 80310
rect 25440 80300 25560 80310
rect 25690 80300 25810 80310
rect 25940 80300 26060 80310
rect 26190 80300 26310 80310
rect 26440 80300 26560 80310
rect 26690 80300 26810 80310
rect 26940 80300 27060 80310
rect 27190 80300 27310 80310
rect 27440 80300 27560 80310
rect 27690 80300 27810 80310
rect 27940 80300 28060 80310
rect 28190 80300 28310 80310
rect 28440 80300 28560 80310
rect 28690 80300 28810 80310
rect 28940 80300 29000 80310
rect 7000 80200 29000 80300
rect 7000 80190 7060 80200
rect 7190 80190 7310 80200
rect 7440 80190 7560 80200
rect 7690 80190 7810 80200
rect 7940 80190 8060 80200
rect 8190 80190 8310 80200
rect 8440 80190 8560 80200
rect 8690 80190 8810 80200
rect 8940 80190 9060 80200
rect 9190 80190 9310 80200
rect 9440 80190 9560 80200
rect 9690 80190 9810 80200
rect 9940 80190 10060 80200
rect 10190 80190 10310 80200
rect 10440 80190 10560 80200
rect 10690 80190 10810 80200
rect 10940 80190 11060 80200
rect 11190 80190 11310 80200
rect 11440 80190 11560 80200
rect 11690 80190 11810 80200
rect 11940 80190 12060 80200
rect 12190 80190 12310 80200
rect 12440 80190 12560 80200
rect 12690 80190 12810 80200
rect 12940 80190 13060 80200
rect 13190 80190 13310 80200
rect 13440 80190 13560 80200
rect 13690 80190 13810 80200
rect 13940 80190 14060 80200
rect 14190 80190 14310 80200
rect 14440 80190 14560 80200
rect 14690 80190 14810 80200
rect 14940 80190 15060 80200
rect 15190 80190 15310 80200
rect 15440 80190 15560 80200
rect 15690 80190 15810 80200
rect 15940 80190 16060 80200
rect 16190 80190 16310 80200
rect 16440 80190 16560 80200
rect 16690 80190 16810 80200
rect 16940 80190 17060 80200
rect 17190 80190 17310 80200
rect 17440 80190 17560 80200
rect 17690 80190 17810 80200
rect 17940 80190 18060 80200
rect 18190 80190 18310 80200
rect 18440 80190 18560 80200
rect 18690 80190 18810 80200
rect 18940 80190 19060 80200
rect 19190 80190 19310 80200
rect 19440 80190 19560 80200
rect 19690 80190 19810 80200
rect 19940 80190 20060 80200
rect 20190 80190 20310 80200
rect 20440 80190 20560 80200
rect 20690 80190 20810 80200
rect 20940 80190 21060 80200
rect 21190 80190 21310 80200
rect 21440 80190 21560 80200
rect 21690 80190 21810 80200
rect 21940 80190 22060 80200
rect 22190 80190 22310 80200
rect 22440 80190 22560 80200
rect 22690 80190 22810 80200
rect 22940 80190 23060 80200
rect 23190 80190 23310 80200
rect 23440 80190 23560 80200
rect 23690 80190 23810 80200
rect 23940 80190 24060 80200
rect 24190 80190 24310 80200
rect 24440 80190 24560 80200
rect 24690 80190 24810 80200
rect 24940 80190 25060 80200
rect 25190 80190 25310 80200
rect 25440 80190 25560 80200
rect 25690 80190 25810 80200
rect 25940 80190 26060 80200
rect 26190 80190 26310 80200
rect 26440 80190 26560 80200
rect 26690 80190 26810 80200
rect 26940 80190 27060 80200
rect 27190 80190 27310 80200
rect 27440 80190 27560 80200
rect 27690 80190 27810 80200
rect 27940 80190 28060 80200
rect 28190 80190 28310 80200
rect 28440 80190 28560 80200
rect 28690 80190 28810 80200
rect 28940 80190 29000 80200
rect 7000 80060 7050 80190
rect 7200 80060 7300 80190
rect 7450 80060 7550 80190
rect 7700 80060 7800 80190
rect 7950 80060 8050 80190
rect 8200 80060 8300 80190
rect 8450 80060 8550 80190
rect 8700 80060 8800 80190
rect 8950 80060 9050 80190
rect 9200 80060 9300 80190
rect 9450 80060 9550 80190
rect 9700 80060 9800 80190
rect 9950 80060 10050 80190
rect 10200 80060 10300 80190
rect 10450 80060 10550 80190
rect 10700 80060 10800 80190
rect 10950 80060 11050 80190
rect 11200 80060 11300 80190
rect 11450 80060 11550 80190
rect 11700 80060 11800 80190
rect 11950 80060 12050 80190
rect 12200 80060 12300 80190
rect 12450 80060 12550 80190
rect 12700 80060 12800 80190
rect 12950 80060 13050 80190
rect 13200 80060 13300 80190
rect 13450 80060 13550 80190
rect 13700 80060 13800 80190
rect 13950 80060 14050 80190
rect 14200 80060 14300 80190
rect 14450 80060 14550 80190
rect 14700 80060 14800 80190
rect 14950 80060 15050 80190
rect 15200 80060 15300 80190
rect 15450 80060 15550 80190
rect 15700 80060 15800 80190
rect 15950 80060 16050 80190
rect 16200 80060 16300 80190
rect 16450 80060 16550 80190
rect 16700 80060 16800 80190
rect 16950 80060 17050 80190
rect 17200 80060 17300 80190
rect 17450 80060 17550 80190
rect 17700 80060 17800 80190
rect 17950 80060 18050 80190
rect 18200 80060 18300 80190
rect 18450 80060 18550 80190
rect 18700 80060 18800 80190
rect 18950 80060 19050 80190
rect 19200 80060 19300 80190
rect 19450 80060 19550 80190
rect 19700 80060 19800 80190
rect 19950 80060 20050 80190
rect 20200 80060 20300 80190
rect 20450 80060 20550 80190
rect 20700 80060 20800 80190
rect 20950 80060 21050 80190
rect 21200 80060 21300 80190
rect 21450 80060 21550 80190
rect 21700 80060 21800 80190
rect 21950 80060 22050 80190
rect 22200 80060 22300 80190
rect 22450 80060 22550 80190
rect 22700 80060 22800 80190
rect 22950 80060 23050 80190
rect 23200 80060 23300 80190
rect 23450 80060 23550 80190
rect 23700 80060 23800 80190
rect 23950 80060 24050 80190
rect 24200 80060 24300 80190
rect 24450 80060 24550 80190
rect 24700 80060 24800 80190
rect 24950 80060 25050 80190
rect 25200 80060 25300 80190
rect 25450 80060 25550 80190
rect 25700 80060 25800 80190
rect 25950 80060 26050 80190
rect 26200 80060 26300 80190
rect 26450 80060 26550 80190
rect 26700 80060 26800 80190
rect 26950 80060 27050 80190
rect 27200 80060 27300 80190
rect 27450 80060 27550 80190
rect 27700 80060 27800 80190
rect 27950 80060 28050 80190
rect 28200 80060 28300 80190
rect 28450 80060 28550 80190
rect 28700 80060 28800 80190
rect 28950 80060 29000 80190
rect 7000 80050 7060 80060
rect 7190 80050 7310 80060
rect 7440 80050 7560 80060
rect 7690 80050 7810 80060
rect 7940 80050 8060 80060
rect 8190 80050 8310 80060
rect 8440 80050 8560 80060
rect 8690 80050 8810 80060
rect 8940 80050 9060 80060
rect 9190 80050 9310 80060
rect 9440 80050 9560 80060
rect 9690 80050 9810 80060
rect 9940 80050 10060 80060
rect 10190 80050 10310 80060
rect 10440 80050 10560 80060
rect 10690 80050 10810 80060
rect 10940 80050 11060 80060
rect 11190 80050 11310 80060
rect 11440 80050 11560 80060
rect 11690 80050 11810 80060
rect 11940 80050 12060 80060
rect 12190 80050 12310 80060
rect 12440 80050 12560 80060
rect 12690 80050 12810 80060
rect 12940 80050 13060 80060
rect 13190 80050 13310 80060
rect 13440 80050 13560 80060
rect 13690 80050 13810 80060
rect 13940 80050 14060 80060
rect 14190 80050 14310 80060
rect 14440 80050 14560 80060
rect 14690 80050 14810 80060
rect 14940 80050 15060 80060
rect 15190 80050 15310 80060
rect 15440 80050 15560 80060
rect 15690 80050 15810 80060
rect 15940 80050 16060 80060
rect 16190 80050 16310 80060
rect 16440 80050 16560 80060
rect 16690 80050 16810 80060
rect 16940 80050 17060 80060
rect 17190 80050 17310 80060
rect 17440 80050 17560 80060
rect 17690 80050 17810 80060
rect 17940 80050 18060 80060
rect 18190 80050 18310 80060
rect 18440 80050 18560 80060
rect 18690 80050 18810 80060
rect 18940 80050 19060 80060
rect 19190 80050 19310 80060
rect 19440 80050 19560 80060
rect 19690 80050 19810 80060
rect 19940 80050 20060 80060
rect 20190 80050 20310 80060
rect 20440 80050 20560 80060
rect 20690 80050 20810 80060
rect 20940 80050 21060 80060
rect 21190 80050 21310 80060
rect 21440 80050 21560 80060
rect 21690 80050 21810 80060
rect 21940 80050 22060 80060
rect 22190 80050 22310 80060
rect 22440 80050 22560 80060
rect 22690 80050 22810 80060
rect 22940 80050 23060 80060
rect 23190 80050 23310 80060
rect 23440 80050 23560 80060
rect 23690 80050 23810 80060
rect 23940 80050 24060 80060
rect 24190 80050 24310 80060
rect 24440 80050 24560 80060
rect 24690 80050 24810 80060
rect 24940 80050 25060 80060
rect 25190 80050 25310 80060
rect 25440 80050 25560 80060
rect 25690 80050 25810 80060
rect 25940 80050 26060 80060
rect 26190 80050 26310 80060
rect 26440 80050 26560 80060
rect 26690 80050 26810 80060
rect 26940 80050 27060 80060
rect 27190 80050 27310 80060
rect 27440 80050 27560 80060
rect 27690 80050 27810 80060
rect 27940 80050 28060 80060
rect 28190 80050 28310 80060
rect 28440 80050 28560 80060
rect 28690 80050 28810 80060
rect 28940 80050 29000 80060
rect 7000 79950 29000 80050
rect 7000 79940 7060 79950
rect 7190 79940 7310 79950
rect 7440 79940 7560 79950
rect 7690 79940 7810 79950
rect 7940 79940 8060 79950
rect 8190 79940 8310 79950
rect 8440 79940 8560 79950
rect 8690 79940 8810 79950
rect 8940 79940 9060 79950
rect 9190 79940 9310 79950
rect 9440 79940 9560 79950
rect 9690 79940 9810 79950
rect 9940 79940 10060 79950
rect 10190 79940 10310 79950
rect 10440 79940 10560 79950
rect 10690 79940 10810 79950
rect 10940 79940 11060 79950
rect 11190 79940 11310 79950
rect 11440 79940 11560 79950
rect 11690 79940 11810 79950
rect 11940 79940 12060 79950
rect 12190 79940 12310 79950
rect 12440 79940 12560 79950
rect 12690 79940 12810 79950
rect 12940 79940 13060 79950
rect 13190 79940 13310 79950
rect 13440 79940 13560 79950
rect 13690 79940 13810 79950
rect 13940 79940 14060 79950
rect 14190 79940 14310 79950
rect 14440 79940 14560 79950
rect 14690 79940 14810 79950
rect 14940 79940 15060 79950
rect 15190 79940 15310 79950
rect 15440 79940 15560 79950
rect 15690 79940 15810 79950
rect 15940 79940 16060 79950
rect 16190 79940 16310 79950
rect 16440 79940 16560 79950
rect 16690 79940 16810 79950
rect 16940 79940 17060 79950
rect 17190 79940 17310 79950
rect 17440 79940 17560 79950
rect 17690 79940 17810 79950
rect 17940 79940 18060 79950
rect 18190 79940 18310 79950
rect 18440 79940 18560 79950
rect 18690 79940 18810 79950
rect 18940 79940 19060 79950
rect 19190 79940 19310 79950
rect 19440 79940 19560 79950
rect 19690 79940 19810 79950
rect 19940 79940 20060 79950
rect 20190 79940 20310 79950
rect 20440 79940 20560 79950
rect 20690 79940 20810 79950
rect 20940 79940 21060 79950
rect 21190 79940 21310 79950
rect 21440 79940 21560 79950
rect 21690 79940 21810 79950
rect 21940 79940 22060 79950
rect 22190 79940 22310 79950
rect 22440 79940 22560 79950
rect 22690 79940 22810 79950
rect 22940 79940 23060 79950
rect 23190 79940 23310 79950
rect 23440 79940 23560 79950
rect 23690 79940 23810 79950
rect 23940 79940 24060 79950
rect 24190 79940 24310 79950
rect 24440 79940 24560 79950
rect 24690 79940 24810 79950
rect 24940 79940 25060 79950
rect 25190 79940 25310 79950
rect 25440 79940 25560 79950
rect 25690 79940 25810 79950
rect 25940 79940 26060 79950
rect 26190 79940 26310 79950
rect 26440 79940 26560 79950
rect 26690 79940 26810 79950
rect 26940 79940 27060 79950
rect 27190 79940 27310 79950
rect 27440 79940 27560 79950
rect 27690 79940 27810 79950
rect 27940 79940 28060 79950
rect 28190 79940 28310 79950
rect 28440 79940 28560 79950
rect 28690 79940 28810 79950
rect 28940 79940 29000 79950
rect 7000 79810 7050 79940
rect 7200 79810 7300 79940
rect 7450 79810 7550 79940
rect 7700 79810 7800 79940
rect 7950 79810 8050 79940
rect 8200 79810 8300 79940
rect 8450 79810 8550 79940
rect 8700 79810 8800 79940
rect 8950 79810 9050 79940
rect 9200 79810 9300 79940
rect 9450 79810 9550 79940
rect 9700 79810 9800 79940
rect 9950 79810 10050 79940
rect 10200 79810 10300 79940
rect 10450 79810 10550 79940
rect 10700 79810 10800 79940
rect 10950 79810 11050 79940
rect 11200 79810 11300 79940
rect 11450 79810 11550 79940
rect 11700 79810 11800 79940
rect 11950 79810 12050 79940
rect 12200 79810 12300 79940
rect 12450 79810 12550 79940
rect 12700 79810 12800 79940
rect 12950 79810 13050 79940
rect 13200 79810 13300 79940
rect 13450 79810 13550 79940
rect 13700 79810 13800 79940
rect 13950 79810 14050 79940
rect 14200 79810 14300 79940
rect 14450 79810 14550 79940
rect 14700 79810 14800 79940
rect 14950 79810 15050 79940
rect 15200 79810 15300 79940
rect 15450 79810 15550 79940
rect 15700 79810 15800 79940
rect 15950 79810 16050 79940
rect 16200 79810 16300 79940
rect 16450 79810 16550 79940
rect 16700 79810 16800 79940
rect 16950 79810 17050 79940
rect 17200 79810 17300 79940
rect 17450 79810 17550 79940
rect 17700 79810 17800 79940
rect 17950 79810 18050 79940
rect 18200 79810 18300 79940
rect 18450 79810 18550 79940
rect 18700 79810 18800 79940
rect 18950 79810 19050 79940
rect 19200 79810 19300 79940
rect 19450 79810 19550 79940
rect 19700 79810 19800 79940
rect 19950 79810 20050 79940
rect 20200 79810 20300 79940
rect 20450 79810 20550 79940
rect 20700 79810 20800 79940
rect 20950 79810 21050 79940
rect 21200 79810 21300 79940
rect 21450 79810 21550 79940
rect 21700 79810 21800 79940
rect 21950 79810 22050 79940
rect 22200 79810 22300 79940
rect 22450 79810 22550 79940
rect 22700 79810 22800 79940
rect 22950 79810 23050 79940
rect 23200 79810 23300 79940
rect 23450 79810 23550 79940
rect 23700 79810 23800 79940
rect 23950 79810 24050 79940
rect 24200 79810 24300 79940
rect 24450 79810 24550 79940
rect 24700 79810 24800 79940
rect 24950 79810 25050 79940
rect 25200 79810 25300 79940
rect 25450 79810 25550 79940
rect 25700 79810 25800 79940
rect 25950 79810 26050 79940
rect 26200 79810 26300 79940
rect 26450 79810 26550 79940
rect 26700 79810 26800 79940
rect 26950 79810 27050 79940
rect 27200 79810 27300 79940
rect 27450 79810 27550 79940
rect 27700 79810 27800 79940
rect 27950 79810 28050 79940
rect 28200 79810 28300 79940
rect 28450 79810 28550 79940
rect 28700 79810 28800 79940
rect 28950 79810 29000 79940
rect 7000 79800 7060 79810
rect 7190 79800 7310 79810
rect 7440 79800 7560 79810
rect 7690 79800 7810 79810
rect 7940 79800 8060 79810
rect 8190 79800 8310 79810
rect 8440 79800 8560 79810
rect 8690 79800 8810 79810
rect 8940 79800 9060 79810
rect 9190 79800 9310 79810
rect 9440 79800 9560 79810
rect 9690 79800 9810 79810
rect 9940 79800 10060 79810
rect 10190 79800 10310 79810
rect 10440 79800 10560 79810
rect 10690 79800 10810 79810
rect 10940 79800 11060 79810
rect 11190 79800 11310 79810
rect 11440 79800 11560 79810
rect 11690 79800 11810 79810
rect 11940 79800 12060 79810
rect 12190 79800 12310 79810
rect 12440 79800 12560 79810
rect 12690 79800 12810 79810
rect 12940 79800 13060 79810
rect 13190 79800 13310 79810
rect 13440 79800 13560 79810
rect 13690 79800 13810 79810
rect 13940 79800 14060 79810
rect 14190 79800 14310 79810
rect 14440 79800 14560 79810
rect 14690 79800 14810 79810
rect 14940 79800 15060 79810
rect 15190 79800 15310 79810
rect 15440 79800 15560 79810
rect 15690 79800 15810 79810
rect 15940 79800 16060 79810
rect 16190 79800 16310 79810
rect 16440 79800 16560 79810
rect 16690 79800 16810 79810
rect 16940 79800 17060 79810
rect 17190 79800 17310 79810
rect 17440 79800 17560 79810
rect 17690 79800 17810 79810
rect 17940 79800 18060 79810
rect 18190 79800 18310 79810
rect 18440 79800 18560 79810
rect 18690 79800 18810 79810
rect 18940 79800 19060 79810
rect 19190 79800 19310 79810
rect 19440 79800 19560 79810
rect 19690 79800 19810 79810
rect 19940 79800 20060 79810
rect 20190 79800 20310 79810
rect 20440 79800 20560 79810
rect 20690 79800 20810 79810
rect 20940 79800 21060 79810
rect 21190 79800 21310 79810
rect 21440 79800 21560 79810
rect 21690 79800 21810 79810
rect 21940 79800 22060 79810
rect 22190 79800 22310 79810
rect 22440 79800 22560 79810
rect 22690 79800 22810 79810
rect 22940 79800 23060 79810
rect 23190 79800 23310 79810
rect 23440 79800 23560 79810
rect 23690 79800 23810 79810
rect 23940 79800 24060 79810
rect 24190 79800 24310 79810
rect 24440 79800 24560 79810
rect 24690 79800 24810 79810
rect 24940 79800 25060 79810
rect 25190 79800 25310 79810
rect 25440 79800 25560 79810
rect 25690 79800 25810 79810
rect 25940 79800 26060 79810
rect 26190 79800 26310 79810
rect 26440 79800 26560 79810
rect 26690 79800 26810 79810
rect 26940 79800 27060 79810
rect 27190 79800 27310 79810
rect 27440 79800 27560 79810
rect 27690 79800 27810 79810
rect 27940 79800 28060 79810
rect 28190 79800 28310 79810
rect 28440 79800 28560 79810
rect 28690 79800 28810 79810
rect 28940 79800 29000 79810
rect 7000 79700 29000 79800
rect 7000 79690 7060 79700
rect 7190 79690 7310 79700
rect 7440 79690 7560 79700
rect 7690 79690 7810 79700
rect 7940 79690 8060 79700
rect 8190 79690 8310 79700
rect 8440 79690 8560 79700
rect 8690 79690 8810 79700
rect 8940 79690 9060 79700
rect 9190 79690 9310 79700
rect 9440 79690 9560 79700
rect 9690 79690 9810 79700
rect 9940 79690 10060 79700
rect 10190 79690 10310 79700
rect 10440 79690 10560 79700
rect 10690 79690 10810 79700
rect 10940 79690 11060 79700
rect 11190 79690 11310 79700
rect 11440 79690 11560 79700
rect 11690 79690 11810 79700
rect 11940 79690 12060 79700
rect 12190 79690 12310 79700
rect 12440 79690 12560 79700
rect 12690 79690 12810 79700
rect 12940 79690 13060 79700
rect 13190 79690 13310 79700
rect 13440 79690 13560 79700
rect 13690 79690 13810 79700
rect 13940 79690 14060 79700
rect 14190 79690 14310 79700
rect 14440 79690 14560 79700
rect 14690 79690 14810 79700
rect 14940 79690 15060 79700
rect 15190 79690 15310 79700
rect 15440 79690 15560 79700
rect 15690 79690 15810 79700
rect 15940 79690 16060 79700
rect 16190 79690 16310 79700
rect 16440 79690 16560 79700
rect 16690 79690 16810 79700
rect 16940 79690 17060 79700
rect 17190 79690 17310 79700
rect 17440 79690 17560 79700
rect 17690 79690 17810 79700
rect 17940 79690 18060 79700
rect 18190 79690 18310 79700
rect 18440 79690 18560 79700
rect 18690 79690 18810 79700
rect 18940 79690 19060 79700
rect 19190 79690 19310 79700
rect 19440 79690 19560 79700
rect 19690 79690 19810 79700
rect 19940 79690 20060 79700
rect 20190 79690 20310 79700
rect 20440 79690 20560 79700
rect 20690 79690 20810 79700
rect 20940 79690 21060 79700
rect 21190 79690 21310 79700
rect 21440 79690 21560 79700
rect 21690 79690 21810 79700
rect 21940 79690 22060 79700
rect 22190 79690 22310 79700
rect 22440 79690 22560 79700
rect 22690 79690 22810 79700
rect 22940 79690 23060 79700
rect 23190 79690 23310 79700
rect 23440 79690 23560 79700
rect 23690 79690 23810 79700
rect 23940 79690 24060 79700
rect 24190 79690 24310 79700
rect 24440 79690 24560 79700
rect 24690 79690 24810 79700
rect 24940 79690 25060 79700
rect 25190 79690 25310 79700
rect 25440 79690 25560 79700
rect 25690 79690 25810 79700
rect 25940 79690 26060 79700
rect 26190 79690 26310 79700
rect 26440 79690 26560 79700
rect 26690 79690 26810 79700
rect 26940 79690 27060 79700
rect 27190 79690 27310 79700
rect 27440 79690 27560 79700
rect 27690 79690 27810 79700
rect 27940 79690 28060 79700
rect 28190 79690 28310 79700
rect 28440 79690 28560 79700
rect 28690 79690 28810 79700
rect 28940 79690 29000 79700
rect 7000 79560 7050 79690
rect 7200 79560 7300 79690
rect 7450 79560 7550 79690
rect 7700 79560 7800 79690
rect 7950 79560 8050 79690
rect 8200 79560 8300 79690
rect 8450 79560 8550 79690
rect 8700 79560 8800 79690
rect 8950 79560 9050 79690
rect 9200 79560 9300 79690
rect 9450 79560 9550 79690
rect 9700 79560 9800 79690
rect 9950 79560 10050 79690
rect 10200 79560 10300 79690
rect 10450 79560 10550 79690
rect 10700 79560 10800 79690
rect 10950 79560 11050 79690
rect 11200 79560 11300 79690
rect 11450 79560 11550 79690
rect 11700 79560 11800 79690
rect 11950 79560 12050 79690
rect 12200 79560 12300 79690
rect 12450 79560 12550 79690
rect 12700 79560 12800 79690
rect 12950 79560 13050 79690
rect 13200 79560 13300 79690
rect 13450 79560 13550 79690
rect 13700 79560 13800 79690
rect 13950 79560 14050 79690
rect 14200 79560 14300 79690
rect 14450 79560 14550 79690
rect 14700 79560 14800 79690
rect 14950 79560 15050 79690
rect 15200 79560 15300 79690
rect 15450 79560 15550 79690
rect 15700 79560 15800 79690
rect 15950 79560 16050 79690
rect 16200 79560 16300 79690
rect 16450 79560 16550 79690
rect 16700 79560 16800 79690
rect 16950 79560 17050 79690
rect 17200 79560 17300 79690
rect 17450 79560 17550 79690
rect 17700 79560 17800 79690
rect 17950 79560 18050 79690
rect 18200 79560 18300 79690
rect 18450 79560 18550 79690
rect 18700 79560 18800 79690
rect 18950 79560 19050 79690
rect 19200 79560 19300 79690
rect 19450 79560 19550 79690
rect 19700 79560 19800 79690
rect 19950 79560 20050 79690
rect 20200 79560 20300 79690
rect 20450 79560 20550 79690
rect 20700 79560 20800 79690
rect 20950 79560 21050 79690
rect 21200 79560 21300 79690
rect 21450 79560 21550 79690
rect 21700 79560 21800 79690
rect 21950 79560 22050 79690
rect 22200 79560 22300 79690
rect 22450 79560 22550 79690
rect 22700 79560 22800 79690
rect 22950 79560 23050 79690
rect 23200 79560 23300 79690
rect 23450 79560 23550 79690
rect 23700 79560 23800 79690
rect 23950 79560 24050 79690
rect 24200 79560 24300 79690
rect 24450 79560 24550 79690
rect 24700 79560 24800 79690
rect 24950 79560 25050 79690
rect 25200 79560 25300 79690
rect 25450 79560 25550 79690
rect 25700 79560 25800 79690
rect 25950 79560 26050 79690
rect 26200 79560 26300 79690
rect 26450 79560 26550 79690
rect 26700 79560 26800 79690
rect 26950 79560 27050 79690
rect 27200 79560 27300 79690
rect 27450 79560 27550 79690
rect 27700 79560 27800 79690
rect 27950 79560 28050 79690
rect 28200 79560 28300 79690
rect 28450 79560 28550 79690
rect 28700 79560 28800 79690
rect 28950 79560 29000 79690
rect 7000 79550 7060 79560
rect 7190 79550 7310 79560
rect 7440 79550 7560 79560
rect 7690 79550 7810 79560
rect 7940 79550 8060 79560
rect 8190 79550 8310 79560
rect 8440 79550 8560 79560
rect 8690 79550 8810 79560
rect 8940 79550 9060 79560
rect 9190 79550 9310 79560
rect 9440 79550 9560 79560
rect 9690 79550 9810 79560
rect 9940 79550 10060 79560
rect 10190 79550 10310 79560
rect 10440 79550 10560 79560
rect 10690 79550 10810 79560
rect 10940 79550 11060 79560
rect 11190 79550 11310 79560
rect 11440 79550 11560 79560
rect 11690 79550 11810 79560
rect 11940 79550 12060 79560
rect 12190 79550 12310 79560
rect 12440 79550 12560 79560
rect 12690 79550 12810 79560
rect 12940 79550 13060 79560
rect 13190 79550 13310 79560
rect 13440 79550 13560 79560
rect 13690 79550 13810 79560
rect 13940 79550 14060 79560
rect 14190 79550 14310 79560
rect 14440 79550 14560 79560
rect 14690 79550 14810 79560
rect 14940 79550 15060 79560
rect 15190 79550 15310 79560
rect 15440 79550 15560 79560
rect 15690 79550 15810 79560
rect 15940 79550 16060 79560
rect 16190 79550 16310 79560
rect 16440 79550 16560 79560
rect 16690 79550 16810 79560
rect 16940 79550 17060 79560
rect 17190 79550 17310 79560
rect 17440 79550 17560 79560
rect 17690 79550 17810 79560
rect 17940 79550 18060 79560
rect 18190 79550 18310 79560
rect 18440 79550 18560 79560
rect 18690 79550 18810 79560
rect 18940 79550 19060 79560
rect 19190 79550 19310 79560
rect 19440 79550 19560 79560
rect 19690 79550 19810 79560
rect 19940 79550 20060 79560
rect 20190 79550 20310 79560
rect 20440 79550 20560 79560
rect 20690 79550 20810 79560
rect 20940 79550 21060 79560
rect 21190 79550 21310 79560
rect 21440 79550 21560 79560
rect 21690 79550 21810 79560
rect 21940 79550 22060 79560
rect 22190 79550 22310 79560
rect 22440 79550 22560 79560
rect 22690 79550 22810 79560
rect 22940 79550 23060 79560
rect 23190 79550 23310 79560
rect 23440 79550 23560 79560
rect 23690 79550 23810 79560
rect 23940 79550 24060 79560
rect 24190 79550 24310 79560
rect 24440 79550 24560 79560
rect 24690 79550 24810 79560
rect 24940 79550 25060 79560
rect 25190 79550 25310 79560
rect 25440 79550 25560 79560
rect 25690 79550 25810 79560
rect 25940 79550 26060 79560
rect 26190 79550 26310 79560
rect 26440 79550 26560 79560
rect 26690 79550 26810 79560
rect 26940 79550 27060 79560
rect 27190 79550 27310 79560
rect 27440 79550 27560 79560
rect 27690 79550 27810 79560
rect 27940 79550 28060 79560
rect 28190 79550 28310 79560
rect 28440 79550 28560 79560
rect 28690 79550 28810 79560
rect 28940 79550 29000 79560
rect 7000 79450 29000 79550
rect 7000 79440 7060 79450
rect 7190 79440 7310 79450
rect 7440 79440 7560 79450
rect 7690 79440 7810 79450
rect 7940 79440 8060 79450
rect 8190 79440 8310 79450
rect 8440 79440 8560 79450
rect 8690 79440 8810 79450
rect 8940 79440 9060 79450
rect 9190 79440 9310 79450
rect 9440 79440 9560 79450
rect 9690 79440 9810 79450
rect 9940 79440 10060 79450
rect 10190 79440 10310 79450
rect 10440 79440 10560 79450
rect 10690 79440 10810 79450
rect 10940 79440 11060 79450
rect 11190 79440 11310 79450
rect 11440 79440 11560 79450
rect 11690 79440 11810 79450
rect 11940 79440 12060 79450
rect 12190 79440 12310 79450
rect 12440 79440 12560 79450
rect 12690 79440 12810 79450
rect 12940 79440 13060 79450
rect 13190 79440 13310 79450
rect 13440 79440 13560 79450
rect 13690 79440 13810 79450
rect 13940 79440 14060 79450
rect 14190 79440 14310 79450
rect 14440 79440 14560 79450
rect 14690 79440 14810 79450
rect 14940 79440 15060 79450
rect 15190 79440 15310 79450
rect 15440 79440 15560 79450
rect 15690 79440 15810 79450
rect 15940 79440 16060 79450
rect 16190 79440 16310 79450
rect 16440 79440 16560 79450
rect 16690 79440 16810 79450
rect 16940 79440 17060 79450
rect 17190 79440 17310 79450
rect 17440 79440 17560 79450
rect 17690 79440 17810 79450
rect 17940 79440 18060 79450
rect 18190 79440 18310 79450
rect 18440 79440 18560 79450
rect 18690 79440 18810 79450
rect 18940 79440 19060 79450
rect 19190 79440 19310 79450
rect 19440 79440 19560 79450
rect 19690 79440 19810 79450
rect 19940 79440 20060 79450
rect 20190 79440 20310 79450
rect 20440 79440 20560 79450
rect 20690 79440 20810 79450
rect 20940 79440 21060 79450
rect 21190 79440 21310 79450
rect 21440 79440 21560 79450
rect 21690 79440 21810 79450
rect 21940 79440 22060 79450
rect 22190 79440 22310 79450
rect 22440 79440 22560 79450
rect 22690 79440 22810 79450
rect 22940 79440 23060 79450
rect 23190 79440 23310 79450
rect 23440 79440 23560 79450
rect 23690 79440 23810 79450
rect 23940 79440 24060 79450
rect 24190 79440 24310 79450
rect 24440 79440 24560 79450
rect 24690 79440 24810 79450
rect 24940 79440 25060 79450
rect 25190 79440 25310 79450
rect 25440 79440 25560 79450
rect 25690 79440 25810 79450
rect 25940 79440 26060 79450
rect 26190 79440 26310 79450
rect 26440 79440 26560 79450
rect 26690 79440 26810 79450
rect 26940 79440 27060 79450
rect 27190 79440 27310 79450
rect 27440 79440 27560 79450
rect 27690 79440 27810 79450
rect 27940 79440 28060 79450
rect 28190 79440 28310 79450
rect 28440 79440 28560 79450
rect 28690 79440 28810 79450
rect 28940 79440 29000 79450
rect 7000 79310 7050 79440
rect 7200 79310 7300 79440
rect 7450 79310 7550 79440
rect 7700 79310 7800 79440
rect 7950 79310 8050 79440
rect 8200 79310 8300 79440
rect 8450 79310 8550 79440
rect 8700 79310 8800 79440
rect 8950 79310 9050 79440
rect 9200 79310 9300 79440
rect 9450 79310 9550 79440
rect 9700 79310 9800 79440
rect 9950 79310 10050 79440
rect 10200 79310 10300 79440
rect 10450 79310 10550 79440
rect 10700 79310 10800 79440
rect 10950 79310 11050 79440
rect 11200 79310 11300 79440
rect 11450 79310 11550 79440
rect 11700 79310 11800 79440
rect 11950 79310 12050 79440
rect 12200 79310 12300 79440
rect 12450 79310 12550 79440
rect 12700 79310 12800 79440
rect 12950 79310 13050 79440
rect 13200 79310 13300 79440
rect 13450 79310 13550 79440
rect 13700 79310 13800 79440
rect 13950 79310 14050 79440
rect 14200 79310 14300 79440
rect 14450 79310 14550 79440
rect 14700 79310 14800 79440
rect 14950 79310 15050 79440
rect 15200 79310 15300 79440
rect 15450 79310 15550 79440
rect 15700 79310 15800 79440
rect 15950 79310 16050 79440
rect 16200 79310 16300 79440
rect 16450 79310 16550 79440
rect 16700 79310 16800 79440
rect 16950 79310 17050 79440
rect 17200 79310 17300 79440
rect 17450 79310 17550 79440
rect 17700 79310 17800 79440
rect 17950 79310 18050 79440
rect 18200 79310 18300 79440
rect 18450 79310 18550 79440
rect 18700 79310 18800 79440
rect 18950 79310 19050 79440
rect 19200 79310 19300 79440
rect 19450 79310 19550 79440
rect 19700 79310 19800 79440
rect 19950 79310 20050 79440
rect 20200 79310 20300 79440
rect 20450 79310 20550 79440
rect 20700 79310 20800 79440
rect 20950 79310 21050 79440
rect 21200 79310 21300 79440
rect 21450 79310 21550 79440
rect 21700 79310 21800 79440
rect 21950 79310 22050 79440
rect 22200 79310 22300 79440
rect 22450 79310 22550 79440
rect 22700 79310 22800 79440
rect 22950 79310 23050 79440
rect 23200 79310 23300 79440
rect 23450 79310 23550 79440
rect 23700 79310 23800 79440
rect 23950 79310 24050 79440
rect 24200 79310 24300 79440
rect 24450 79310 24550 79440
rect 24700 79310 24800 79440
rect 24950 79310 25050 79440
rect 25200 79310 25300 79440
rect 25450 79310 25550 79440
rect 25700 79310 25800 79440
rect 25950 79310 26050 79440
rect 26200 79310 26300 79440
rect 26450 79310 26550 79440
rect 26700 79310 26800 79440
rect 26950 79310 27050 79440
rect 27200 79310 27300 79440
rect 27450 79310 27550 79440
rect 27700 79310 27800 79440
rect 27950 79310 28050 79440
rect 28200 79310 28300 79440
rect 28450 79310 28550 79440
rect 28700 79310 28800 79440
rect 28950 79310 29000 79440
rect 7000 79300 7060 79310
rect 7190 79300 7310 79310
rect 7440 79300 7560 79310
rect 7690 79300 7810 79310
rect 7940 79300 8060 79310
rect 8190 79300 8310 79310
rect 8440 79300 8560 79310
rect 8690 79300 8810 79310
rect 8940 79300 9060 79310
rect 9190 79300 9310 79310
rect 9440 79300 9560 79310
rect 9690 79300 9810 79310
rect 9940 79300 10060 79310
rect 10190 79300 10310 79310
rect 10440 79300 10560 79310
rect 10690 79300 10810 79310
rect 10940 79300 11060 79310
rect 11190 79300 11310 79310
rect 11440 79300 11560 79310
rect 11690 79300 11810 79310
rect 11940 79300 12060 79310
rect 12190 79300 12310 79310
rect 12440 79300 12560 79310
rect 12690 79300 12810 79310
rect 12940 79300 13060 79310
rect 13190 79300 13310 79310
rect 13440 79300 13560 79310
rect 13690 79300 13810 79310
rect 13940 79300 14060 79310
rect 14190 79300 14310 79310
rect 14440 79300 14560 79310
rect 14690 79300 14810 79310
rect 14940 79300 15060 79310
rect 15190 79300 15310 79310
rect 15440 79300 15560 79310
rect 15690 79300 15810 79310
rect 15940 79300 16060 79310
rect 16190 79300 16310 79310
rect 16440 79300 16560 79310
rect 16690 79300 16810 79310
rect 16940 79300 17060 79310
rect 17190 79300 17310 79310
rect 17440 79300 17560 79310
rect 17690 79300 17810 79310
rect 17940 79300 18060 79310
rect 18190 79300 18310 79310
rect 18440 79300 18560 79310
rect 18690 79300 18810 79310
rect 18940 79300 19060 79310
rect 19190 79300 19310 79310
rect 19440 79300 19560 79310
rect 19690 79300 19810 79310
rect 19940 79300 20060 79310
rect 20190 79300 20310 79310
rect 20440 79300 20560 79310
rect 20690 79300 20810 79310
rect 20940 79300 21060 79310
rect 21190 79300 21310 79310
rect 21440 79300 21560 79310
rect 21690 79300 21810 79310
rect 21940 79300 22060 79310
rect 22190 79300 22310 79310
rect 22440 79300 22560 79310
rect 22690 79300 22810 79310
rect 22940 79300 23060 79310
rect 23190 79300 23310 79310
rect 23440 79300 23560 79310
rect 23690 79300 23810 79310
rect 23940 79300 24060 79310
rect 24190 79300 24310 79310
rect 24440 79300 24560 79310
rect 24690 79300 24810 79310
rect 24940 79300 25060 79310
rect 25190 79300 25310 79310
rect 25440 79300 25560 79310
rect 25690 79300 25810 79310
rect 25940 79300 26060 79310
rect 26190 79300 26310 79310
rect 26440 79300 26560 79310
rect 26690 79300 26810 79310
rect 26940 79300 27060 79310
rect 27190 79300 27310 79310
rect 27440 79300 27560 79310
rect 27690 79300 27810 79310
rect 27940 79300 28060 79310
rect 28190 79300 28310 79310
rect 28440 79300 28560 79310
rect 28690 79300 28810 79310
rect 28940 79300 29000 79310
rect 7000 79200 29000 79300
rect 7000 79190 7060 79200
rect 7190 79190 7310 79200
rect 7440 79190 7560 79200
rect 7690 79190 7810 79200
rect 7940 79190 8060 79200
rect 8190 79190 8310 79200
rect 8440 79190 8560 79200
rect 8690 79190 8810 79200
rect 8940 79190 9060 79200
rect 9190 79190 9310 79200
rect 9440 79190 9560 79200
rect 9690 79190 9810 79200
rect 9940 79190 10060 79200
rect 10190 79190 10310 79200
rect 10440 79190 10560 79200
rect 10690 79190 10810 79200
rect 10940 79190 11060 79200
rect 11190 79190 11310 79200
rect 11440 79190 11560 79200
rect 11690 79190 11810 79200
rect 11940 79190 12060 79200
rect 12190 79190 12310 79200
rect 12440 79190 12560 79200
rect 12690 79190 12810 79200
rect 12940 79190 13060 79200
rect 13190 79190 13310 79200
rect 13440 79190 13560 79200
rect 13690 79190 13810 79200
rect 13940 79190 14060 79200
rect 14190 79190 14310 79200
rect 14440 79190 14560 79200
rect 14690 79190 14810 79200
rect 14940 79190 15060 79200
rect 15190 79190 15310 79200
rect 15440 79190 15560 79200
rect 15690 79190 15810 79200
rect 15940 79190 16060 79200
rect 16190 79190 16310 79200
rect 16440 79190 16560 79200
rect 16690 79190 16810 79200
rect 16940 79190 17060 79200
rect 17190 79190 17310 79200
rect 17440 79190 17560 79200
rect 17690 79190 17810 79200
rect 17940 79190 18060 79200
rect 18190 79190 18310 79200
rect 18440 79190 18560 79200
rect 18690 79190 18810 79200
rect 18940 79190 19060 79200
rect 19190 79190 19310 79200
rect 19440 79190 19560 79200
rect 19690 79190 19810 79200
rect 19940 79190 20060 79200
rect 20190 79190 20310 79200
rect 20440 79190 20560 79200
rect 20690 79190 20810 79200
rect 20940 79190 21060 79200
rect 21190 79190 21310 79200
rect 21440 79190 21560 79200
rect 21690 79190 21810 79200
rect 21940 79190 22060 79200
rect 22190 79190 22310 79200
rect 22440 79190 22560 79200
rect 22690 79190 22810 79200
rect 22940 79190 23060 79200
rect 23190 79190 23310 79200
rect 23440 79190 23560 79200
rect 23690 79190 23810 79200
rect 23940 79190 24060 79200
rect 24190 79190 24310 79200
rect 24440 79190 24560 79200
rect 24690 79190 24810 79200
rect 24940 79190 25060 79200
rect 25190 79190 25310 79200
rect 25440 79190 25560 79200
rect 25690 79190 25810 79200
rect 25940 79190 26060 79200
rect 26190 79190 26310 79200
rect 26440 79190 26560 79200
rect 26690 79190 26810 79200
rect 26940 79190 27060 79200
rect 27190 79190 27310 79200
rect 27440 79190 27560 79200
rect 27690 79190 27810 79200
rect 27940 79190 28060 79200
rect 28190 79190 28310 79200
rect 28440 79190 28560 79200
rect 28690 79190 28810 79200
rect 28940 79190 29000 79200
rect 7000 79060 7050 79190
rect 7200 79060 7300 79190
rect 7450 79060 7550 79190
rect 7700 79060 7800 79190
rect 7950 79060 8050 79190
rect 8200 79060 8300 79190
rect 8450 79060 8550 79190
rect 8700 79060 8800 79190
rect 8950 79060 9050 79190
rect 9200 79060 9300 79190
rect 9450 79060 9550 79190
rect 9700 79060 9800 79190
rect 9950 79060 10050 79190
rect 10200 79060 10300 79190
rect 10450 79060 10550 79190
rect 10700 79060 10800 79190
rect 10950 79060 11050 79190
rect 11200 79060 11300 79190
rect 11450 79060 11550 79190
rect 11700 79060 11800 79190
rect 11950 79060 12050 79190
rect 12200 79060 12300 79190
rect 12450 79060 12550 79190
rect 12700 79060 12800 79190
rect 12950 79060 13050 79190
rect 13200 79060 13300 79190
rect 13450 79060 13550 79190
rect 13700 79060 13800 79190
rect 13950 79060 14050 79190
rect 14200 79060 14300 79190
rect 14450 79060 14550 79190
rect 14700 79060 14800 79190
rect 14950 79060 15050 79190
rect 15200 79060 15300 79190
rect 15450 79060 15550 79190
rect 15700 79060 15800 79190
rect 15950 79060 16050 79190
rect 16200 79060 16300 79190
rect 16450 79060 16550 79190
rect 16700 79060 16800 79190
rect 16950 79060 17050 79190
rect 17200 79060 17300 79190
rect 17450 79060 17550 79190
rect 17700 79060 17800 79190
rect 17950 79060 18050 79190
rect 18200 79060 18300 79190
rect 18450 79060 18550 79190
rect 18700 79060 18800 79190
rect 18950 79060 19050 79190
rect 19200 79060 19300 79190
rect 19450 79060 19550 79190
rect 19700 79060 19800 79190
rect 19950 79060 20050 79190
rect 20200 79060 20300 79190
rect 20450 79060 20550 79190
rect 20700 79060 20800 79190
rect 20950 79060 21050 79190
rect 21200 79060 21300 79190
rect 21450 79060 21550 79190
rect 21700 79060 21800 79190
rect 21950 79060 22050 79190
rect 22200 79060 22300 79190
rect 22450 79060 22550 79190
rect 22700 79060 22800 79190
rect 22950 79060 23050 79190
rect 23200 79060 23300 79190
rect 23450 79060 23550 79190
rect 23700 79060 23800 79190
rect 23950 79060 24050 79190
rect 24200 79060 24300 79190
rect 24450 79060 24550 79190
rect 24700 79060 24800 79190
rect 24950 79060 25050 79190
rect 25200 79060 25300 79190
rect 25450 79060 25550 79190
rect 25700 79060 25800 79190
rect 25950 79060 26050 79190
rect 26200 79060 26300 79190
rect 26450 79060 26550 79190
rect 26700 79060 26800 79190
rect 26950 79060 27050 79190
rect 27200 79060 27300 79190
rect 27450 79060 27550 79190
rect 27700 79060 27800 79190
rect 27950 79060 28050 79190
rect 28200 79060 28300 79190
rect 28450 79060 28550 79190
rect 28700 79060 28800 79190
rect 28950 79060 29000 79190
rect 7000 79050 7060 79060
rect 7190 79050 7310 79060
rect 7440 79050 7560 79060
rect 7690 79050 7810 79060
rect 7940 79050 8060 79060
rect 8190 79050 8310 79060
rect 8440 79050 8560 79060
rect 8690 79050 8810 79060
rect 8940 79050 9060 79060
rect 9190 79050 9310 79060
rect 9440 79050 9560 79060
rect 9690 79050 9810 79060
rect 9940 79050 10060 79060
rect 10190 79050 10310 79060
rect 10440 79050 10560 79060
rect 10690 79050 10810 79060
rect 10940 79050 11060 79060
rect 11190 79050 11310 79060
rect 11440 79050 11560 79060
rect 11690 79050 11810 79060
rect 11940 79050 12060 79060
rect 12190 79050 12310 79060
rect 12440 79050 12560 79060
rect 12690 79050 12810 79060
rect 12940 79050 13060 79060
rect 13190 79050 13310 79060
rect 13440 79050 13560 79060
rect 13690 79050 13810 79060
rect 13940 79050 14060 79060
rect 14190 79050 14310 79060
rect 14440 79050 14560 79060
rect 14690 79050 14810 79060
rect 14940 79050 15060 79060
rect 15190 79050 15310 79060
rect 15440 79050 15560 79060
rect 15690 79050 15810 79060
rect 15940 79050 16060 79060
rect 16190 79050 16310 79060
rect 16440 79050 16560 79060
rect 16690 79050 16810 79060
rect 16940 79050 17060 79060
rect 17190 79050 17310 79060
rect 17440 79050 17560 79060
rect 17690 79050 17810 79060
rect 17940 79050 18060 79060
rect 18190 79050 18310 79060
rect 18440 79050 18560 79060
rect 18690 79050 18810 79060
rect 18940 79050 19060 79060
rect 19190 79050 19310 79060
rect 19440 79050 19560 79060
rect 19690 79050 19810 79060
rect 19940 79050 20060 79060
rect 20190 79050 20310 79060
rect 20440 79050 20560 79060
rect 20690 79050 20810 79060
rect 20940 79050 21060 79060
rect 21190 79050 21310 79060
rect 21440 79050 21560 79060
rect 21690 79050 21810 79060
rect 21940 79050 22060 79060
rect 22190 79050 22310 79060
rect 22440 79050 22560 79060
rect 22690 79050 22810 79060
rect 22940 79050 23060 79060
rect 23190 79050 23310 79060
rect 23440 79050 23560 79060
rect 23690 79050 23810 79060
rect 23940 79050 24060 79060
rect 24190 79050 24310 79060
rect 24440 79050 24560 79060
rect 24690 79050 24810 79060
rect 24940 79050 25060 79060
rect 25190 79050 25310 79060
rect 25440 79050 25560 79060
rect 25690 79050 25810 79060
rect 25940 79050 26060 79060
rect 26190 79050 26310 79060
rect 26440 79050 26560 79060
rect 26690 79050 26810 79060
rect 26940 79050 27060 79060
rect 27190 79050 27310 79060
rect 27440 79050 27560 79060
rect 27690 79050 27810 79060
rect 27940 79050 28060 79060
rect 28190 79050 28310 79060
rect 28440 79050 28560 79060
rect 28690 79050 28810 79060
rect 28940 79050 29000 79060
rect 7000 78950 29000 79050
rect 7000 78940 7060 78950
rect 7190 78940 7310 78950
rect 7440 78940 7560 78950
rect 7690 78940 7810 78950
rect 7940 78940 8060 78950
rect 8190 78940 8310 78950
rect 8440 78940 8560 78950
rect 8690 78940 8810 78950
rect 8940 78940 9060 78950
rect 9190 78940 9310 78950
rect 9440 78940 9560 78950
rect 9690 78940 9810 78950
rect 9940 78940 10060 78950
rect 10190 78940 10310 78950
rect 10440 78940 10560 78950
rect 10690 78940 10810 78950
rect 10940 78940 11060 78950
rect 11190 78940 11310 78950
rect 11440 78940 11560 78950
rect 11690 78940 11810 78950
rect 11940 78940 12060 78950
rect 12190 78940 12310 78950
rect 12440 78940 12560 78950
rect 12690 78940 12810 78950
rect 12940 78940 13060 78950
rect 13190 78940 13310 78950
rect 13440 78940 13560 78950
rect 13690 78940 13810 78950
rect 13940 78940 14060 78950
rect 14190 78940 14310 78950
rect 14440 78940 14560 78950
rect 14690 78940 14810 78950
rect 14940 78940 15060 78950
rect 15190 78940 15310 78950
rect 15440 78940 15560 78950
rect 15690 78940 15810 78950
rect 15940 78940 16060 78950
rect 16190 78940 16310 78950
rect 16440 78940 16560 78950
rect 16690 78940 16810 78950
rect 16940 78940 17060 78950
rect 17190 78940 17310 78950
rect 17440 78940 17560 78950
rect 17690 78940 17810 78950
rect 17940 78940 18060 78950
rect 18190 78940 18310 78950
rect 18440 78940 18560 78950
rect 18690 78940 18810 78950
rect 18940 78940 19060 78950
rect 19190 78940 19310 78950
rect 19440 78940 19560 78950
rect 19690 78940 19810 78950
rect 19940 78940 20060 78950
rect 20190 78940 20310 78950
rect 20440 78940 20560 78950
rect 20690 78940 20810 78950
rect 20940 78940 21060 78950
rect 21190 78940 21310 78950
rect 21440 78940 21560 78950
rect 21690 78940 21810 78950
rect 21940 78940 22060 78950
rect 22190 78940 22310 78950
rect 22440 78940 22560 78950
rect 22690 78940 22810 78950
rect 22940 78940 23060 78950
rect 23190 78940 23310 78950
rect 23440 78940 23560 78950
rect 23690 78940 23810 78950
rect 23940 78940 24060 78950
rect 24190 78940 24310 78950
rect 24440 78940 24560 78950
rect 24690 78940 24810 78950
rect 24940 78940 25060 78950
rect 25190 78940 25310 78950
rect 25440 78940 25560 78950
rect 25690 78940 25810 78950
rect 25940 78940 26060 78950
rect 26190 78940 26310 78950
rect 26440 78940 26560 78950
rect 26690 78940 26810 78950
rect 26940 78940 27060 78950
rect 27190 78940 27310 78950
rect 27440 78940 27560 78950
rect 27690 78940 27810 78950
rect 27940 78940 28060 78950
rect 28190 78940 28310 78950
rect 28440 78940 28560 78950
rect 28690 78940 28810 78950
rect 28940 78940 29000 78950
rect 7000 78810 7050 78940
rect 7200 78810 7300 78940
rect 7450 78810 7550 78940
rect 7700 78810 7800 78940
rect 7950 78810 8050 78940
rect 8200 78810 8300 78940
rect 8450 78810 8550 78940
rect 8700 78810 8800 78940
rect 8950 78810 9050 78940
rect 9200 78810 9300 78940
rect 9450 78810 9550 78940
rect 9700 78810 9800 78940
rect 9950 78810 10050 78940
rect 10200 78810 10300 78940
rect 10450 78810 10550 78940
rect 10700 78810 10800 78940
rect 10950 78810 11050 78940
rect 11200 78810 11300 78940
rect 11450 78810 11550 78940
rect 11700 78810 11800 78940
rect 11950 78810 12050 78940
rect 12200 78810 12300 78940
rect 12450 78810 12550 78940
rect 12700 78810 12800 78940
rect 12950 78810 13050 78940
rect 13200 78810 13300 78940
rect 13450 78810 13550 78940
rect 13700 78810 13800 78940
rect 13950 78810 14050 78940
rect 14200 78810 14300 78940
rect 14450 78810 14550 78940
rect 14700 78810 14800 78940
rect 14950 78810 15050 78940
rect 15200 78810 15300 78940
rect 15450 78810 15550 78940
rect 15700 78810 15800 78940
rect 15950 78810 16050 78940
rect 16200 78810 16300 78940
rect 16450 78810 16550 78940
rect 16700 78810 16800 78940
rect 16950 78810 17050 78940
rect 17200 78810 17300 78940
rect 17450 78810 17550 78940
rect 17700 78810 17800 78940
rect 17950 78810 18050 78940
rect 18200 78810 18300 78940
rect 18450 78810 18550 78940
rect 18700 78810 18800 78940
rect 18950 78810 19050 78940
rect 19200 78810 19300 78940
rect 19450 78810 19550 78940
rect 19700 78810 19800 78940
rect 19950 78810 20050 78940
rect 20200 78810 20300 78940
rect 20450 78810 20550 78940
rect 20700 78810 20800 78940
rect 20950 78810 21050 78940
rect 21200 78810 21300 78940
rect 21450 78810 21550 78940
rect 21700 78810 21800 78940
rect 21950 78810 22050 78940
rect 22200 78810 22300 78940
rect 22450 78810 22550 78940
rect 22700 78810 22800 78940
rect 22950 78810 23050 78940
rect 23200 78810 23300 78940
rect 23450 78810 23550 78940
rect 23700 78810 23800 78940
rect 23950 78810 24050 78940
rect 24200 78810 24300 78940
rect 24450 78810 24550 78940
rect 24700 78810 24800 78940
rect 24950 78810 25050 78940
rect 25200 78810 25300 78940
rect 25450 78810 25550 78940
rect 25700 78810 25800 78940
rect 25950 78810 26050 78940
rect 26200 78810 26300 78940
rect 26450 78810 26550 78940
rect 26700 78810 26800 78940
rect 26950 78810 27050 78940
rect 27200 78810 27300 78940
rect 27450 78810 27550 78940
rect 27700 78810 27800 78940
rect 27950 78810 28050 78940
rect 28200 78810 28300 78940
rect 28450 78810 28550 78940
rect 28700 78810 28800 78940
rect 28950 78810 29000 78940
rect 7000 78800 7060 78810
rect 7190 78800 7310 78810
rect 7440 78800 7560 78810
rect 7690 78800 7810 78810
rect 7940 78800 8060 78810
rect 8190 78800 8310 78810
rect 8440 78800 8560 78810
rect 8690 78800 8810 78810
rect 8940 78800 9060 78810
rect 9190 78800 9310 78810
rect 9440 78800 9560 78810
rect 9690 78800 9810 78810
rect 9940 78800 10060 78810
rect 10190 78800 10310 78810
rect 10440 78800 10560 78810
rect 10690 78800 10810 78810
rect 10940 78800 11060 78810
rect 11190 78800 11310 78810
rect 11440 78800 11560 78810
rect 11690 78800 11810 78810
rect 11940 78800 12060 78810
rect 12190 78800 12310 78810
rect 12440 78800 12560 78810
rect 12690 78800 12810 78810
rect 12940 78800 13060 78810
rect 13190 78800 13310 78810
rect 13440 78800 13560 78810
rect 13690 78800 13810 78810
rect 13940 78800 14060 78810
rect 14190 78800 14310 78810
rect 14440 78800 14560 78810
rect 14690 78800 14810 78810
rect 14940 78800 15060 78810
rect 15190 78800 15310 78810
rect 15440 78800 15560 78810
rect 15690 78800 15810 78810
rect 15940 78800 16060 78810
rect 16190 78800 16310 78810
rect 16440 78800 16560 78810
rect 16690 78800 16810 78810
rect 16940 78800 17060 78810
rect 17190 78800 17310 78810
rect 17440 78800 17560 78810
rect 17690 78800 17810 78810
rect 17940 78800 18060 78810
rect 18190 78800 18310 78810
rect 18440 78800 18560 78810
rect 18690 78800 18810 78810
rect 18940 78800 19060 78810
rect 19190 78800 19310 78810
rect 19440 78800 19560 78810
rect 19690 78800 19810 78810
rect 19940 78800 20060 78810
rect 20190 78800 20310 78810
rect 20440 78800 20560 78810
rect 20690 78800 20810 78810
rect 20940 78800 21060 78810
rect 21190 78800 21310 78810
rect 21440 78800 21560 78810
rect 21690 78800 21810 78810
rect 21940 78800 22060 78810
rect 22190 78800 22310 78810
rect 22440 78800 22560 78810
rect 22690 78800 22810 78810
rect 22940 78800 23060 78810
rect 23190 78800 23310 78810
rect 23440 78800 23560 78810
rect 23690 78800 23810 78810
rect 23940 78800 24060 78810
rect 24190 78800 24310 78810
rect 24440 78800 24560 78810
rect 24690 78800 24810 78810
rect 24940 78800 25060 78810
rect 25190 78800 25310 78810
rect 25440 78800 25560 78810
rect 25690 78800 25810 78810
rect 25940 78800 26060 78810
rect 26190 78800 26310 78810
rect 26440 78800 26560 78810
rect 26690 78800 26810 78810
rect 26940 78800 27060 78810
rect 27190 78800 27310 78810
rect 27440 78800 27560 78810
rect 27690 78800 27810 78810
rect 27940 78800 28060 78810
rect 28190 78800 28310 78810
rect 28440 78800 28560 78810
rect 28690 78800 28810 78810
rect 28940 78800 29000 78810
rect 7000 78700 29000 78800
rect 7000 78690 7060 78700
rect 7190 78690 7310 78700
rect 7440 78690 7560 78700
rect 7690 78690 7810 78700
rect 7940 78690 8060 78700
rect 8190 78690 8310 78700
rect 8440 78690 8560 78700
rect 8690 78690 8810 78700
rect 8940 78690 9060 78700
rect 9190 78690 9310 78700
rect 9440 78690 9560 78700
rect 9690 78690 9810 78700
rect 9940 78690 10060 78700
rect 10190 78690 10310 78700
rect 10440 78690 10560 78700
rect 10690 78690 10810 78700
rect 10940 78690 11060 78700
rect 11190 78690 11310 78700
rect 11440 78690 11560 78700
rect 11690 78690 11810 78700
rect 11940 78690 12060 78700
rect 12190 78690 12310 78700
rect 12440 78690 12560 78700
rect 12690 78690 12810 78700
rect 12940 78690 13060 78700
rect 13190 78690 13310 78700
rect 13440 78690 13560 78700
rect 13690 78690 13810 78700
rect 13940 78690 14060 78700
rect 14190 78690 14310 78700
rect 14440 78690 14560 78700
rect 14690 78690 14810 78700
rect 14940 78690 15060 78700
rect 15190 78690 15310 78700
rect 15440 78690 15560 78700
rect 15690 78690 15810 78700
rect 15940 78690 16060 78700
rect 16190 78690 16310 78700
rect 16440 78690 16560 78700
rect 16690 78690 16810 78700
rect 16940 78690 17060 78700
rect 17190 78690 17310 78700
rect 17440 78690 17560 78700
rect 17690 78690 17810 78700
rect 17940 78690 18060 78700
rect 18190 78690 18310 78700
rect 18440 78690 18560 78700
rect 18690 78690 18810 78700
rect 18940 78690 19060 78700
rect 19190 78690 19310 78700
rect 19440 78690 19560 78700
rect 19690 78690 19810 78700
rect 19940 78690 20060 78700
rect 20190 78690 20310 78700
rect 20440 78690 20560 78700
rect 20690 78690 20810 78700
rect 20940 78690 21060 78700
rect 21190 78690 21310 78700
rect 21440 78690 21560 78700
rect 21690 78690 21810 78700
rect 21940 78690 22060 78700
rect 22190 78690 22310 78700
rect 22440 78690 22560 78700
rect 22690 78690 22810 78700
rect 22940 78690 23060 78700
rect 23190 78690 23310 78700
rect 23440 78690 23560 78700
rect 23690 78690 23810 78700
rect 23940 78690 24060 78700
rect 24190 78690 24310 78700
rect 24440 78690 24560 78700
rect 24690 78690 24810 78700
rect 24940 78690 25060 78700
rect 25190 78690 25310 78700
rect 25440 78690 25560 78700
rect 25690 78690 25810 78700
rect 25940 78690 26060 78700
rect 26190 78690 26310 78700
rect 26440 78690 26560 78700
rect 26690 78690 26810 78700
rect 26940 78690 27060 78700
rect 27190 78690 27310 78700
rect 27440 78690 27560 78700
rect 27690 78690 27810 78700
rect 27940 78690 28060 78700
rect 28190 78690 28310 78700
rect 28440 78690 28560 78700
rect 28690 78690 28810 78700
rect 28940 78690 29000 78700
rect 7000 78560 7050 78690
rect 7200 78560 7300 78690
rect 7450 78560 7550 78690
rect 7700 78560 7800 78690
rect 7950 78560 8050 78690
rect 8200 78560 8300 78690
rect 8450 78560 8550 78690
rect 8700 78560 8800 78690
rect 8950 78560 9050 78690
rect 9200 78560 9300 78690
rect 9450 78560 9550 78690
rect 9700 78560 9800 78690
rect 9950 78560 10050 78690
rect 10200 78560 10300 78690
rect 10450 78560 10550 78690
rect 10700 78560 10800 78690
rect 10950 78560 11050 78690
rect 11200 78560 11300 78690
rect 11450 78560 11550 78690
rect 11700 78560 11800 78690
rect 11950 78560 12050 78690
rect 12200 78560 12300 78690
rect 12450 78560 12550 78690
rect 12700 78560 12800 78690
rect 12950 78560 13050 78690
rect 13200 78560 13300 78690
rect 13450 78560 13550 78690
rect 13700 78560 13800 78690
rect 13950 78560 14050 78690
rect 14200 78560 14300 78690
rect 14450 78560 14550 78690
rect 14700 78560 14800 78690
rect 14950 78560 15050 78690
rect 15200 78560 15300 78690
rect 15450 78560 15550 78690
rect 15700 78560 15800 78690
rect 15950 78560 16050 78690
rect 16200 78560 16300 78690
rect 16450 78560 16550 78690
rect 16700 78560 16800 78690
rect 16950 78560 17050 78690
rect 17200 78560 17300 78690
rect 17450 78560 17550 78690
rect 17700 78560 17800 78690
rect 17950 78560 18050 78690
rect 18200 78560 18300 78690
rect 18450 78560 18550 78690
rect 18700 78560 18800 78690
rect 18950 78560 19050 78690
rect 19200 78560 19300 78690
rect 19450 78560 19550 78690
rect 19700 78560 19800 78690
rect 19950 78560 20050 78690
rect 20200 78560 20300 78690
rect 20450 78560 20550 78690
rect 20700 78560 20800 78690
rect 20950 78560 21050 78690
rect 21200 78560 21300 78690
rect 21450 78560 21550 78690
rect 21700 78560 21800 78690
rect 21950 78560 22050 78690
rect 22200 78560 22300 78690
rect 22450 78560 22550 78690
rect 22700 78560 22800 78690
rect 22950 78560 23050 78690
rect 23200 78560 23300 78690
rect 23450 78560 23550 78690
rect 23700 78560 23800 78690
rect 23950 78560 24050 78690
rect 24200 78560 24300 78690
rect 24450 78560 24550 78690
rect 24700 78560 24800 78690
rect 24950 78560 25050 78690
rect 25200 78560 25300 78690
rect 25450 78560 25550 78690
rect 25700 78560 25800 78690
rect 25950 78560 26050 78690
rect 26200 78560 26300 78690
rect 26450 78560 26550 78690
rect 26700 78560 26800 78690
rect 26950 78560 27050 78690
rect 27200 78560 27300 78690
rect 27450 78560 27550 78690
rect 27700 78560 27800 78690
rect 27950 78560 28050 78690
rect 28200 78560 28300 78690
rect 28450 78560 28550 78690
rect 28700 78560 28800 78690
rect 28950 78560 29000 78690
rect 7000 78550 7060 78560
rect 7190 78550 7310 78560
rect 7440 78550 7560 78560
rect 7690 78550 7810 78560
rect 7940 78550 8060 78560
rect 8190 78550 8310 78560
rect 8440 78550 8560 78560
rect 8690 78550 8810 78560
rect 8940 78550 9060 78560
rect 9190 78550 9310 78560
rect 9440 78550 9560 78560
rect 9690 78550 9810 78560
rect 9940 78550 10060 78560
rect 10190 78550 10310 78560
rect 10440 78550 10560 78560
rect 10690 78550 10810 78560
rect 10940 78550 11060 78560
rect 11190 78550 11310 78560
rect 11440 78550 11560 78560
rect 11690 78550 11810 78560
rect 11940 78550 12060 78560
rect 12190 78550 12310 78560
rect 12440 78550 12560 78560
rect 12690 78550 12810 78560
rect 12940 78550 13060 78560
rect 13190 78550 13310 78560
rect 13440 78550 13560 78560
rect 13690 78550 13810 78560
rect 13940 78550 14060 78560
rect 14190 78550 14310 78560
rect 14440 78550 14560 78560
rect 14690 78550 14810 78560
rect 14940 78550 15060 78560
rect 15190 78550 15310 78560
rect 15440 78550 15560 78560
rect 15690 78550 15810 78560
rect 15940 78550 16060 78560
rect 16190 78550 16310 78560
rect 16440 78550 16560 78560
rect 16690 78550 16810 78560
rect 16940 78550 17060 78560
rect 17190 78550 17310 78560
rect 17440 78550 17560 78560
rect 17690 78550 17810 78560
rect 17940 78550 18060 78560
rect 18190 78550 18310 78560
rect 18440 78550 18560 78560
rect 18690 78550 18810 78560
rect 18940 78550 19060 78560
rect 19190 78550 19310 78560
rect 19440 78550 19560 78560
rect 19690 78550 19810 78560
rect 19940 78550 20060 78560
rect 20190 78550 20310 78560
rect 20440 78550 20560 78560
rect 20690 78550 20810 78560
rect 20940 78550 21060 78560
rect 21190 78550 21310 78560
rect 21440 78550 21560 78560
rect 21690 78550 21810 78560
rect 21940 78550 22060 78560
rect 22190 78550 22310 78560
rect 22440 78550 22560 78560
rect 22690 78550 22810 78560
rect 22940 78550 23060 78560
rect 23190 78550 23310 78560
rect 23440 78550 23560 78560
rect 23690 78550 23810 78560
rect 23940 78550 24060 78560
rect 24190 78550 24310 78560
rect 24440 78550 24560 78560
rect 24690 78550 24810 78560
rect 24940 78550 25060 78560
rect 25190 78550 25310 78560
rect 25440 78550 25560 78560
rect 25690 78550 25810 78560
rect 25940 78550 26060 78560
rect 26190 78550 26310 78560
rect 26440 78550 26560 78560
rect 26690 78550 26810 78560
rect 26940 78550 27060 78560
rect 27190 78550 27310 78560
rect 27440 78550 27560 78560
rect 27690 78550 27810 78560
rect 27940 78550 28060 78560
rect 28190 78550 28310 78560
rect 28440 78550 28560 78560
rect 28690 78550 28810 78560
rect 28940 78550 29000 78560
rect 7000 78450 29000 78550
rect 7000 78440 7060 78450
rect 7190 78440 7310 78450
rect 7440 78440 7560 78450
rect 7690 78440 7810 78450
rect 7940 78440 8060 78450
rect 8190 78440 8310 78450
rect 8440 78440 8560 78450
rect 8690 78440 8810 78450
rect 8940 78440 9060 78450
rect 9190 78440 9310 78450
rect 9440 78440 9560 78450
rect 9690 78440 9810 78450
rect 9940 78440 10060 78450
rect 10190 78440 10310 78450
rect 10440 78440 10560 78450
rect 10690 78440 10810 78450
rect 10940 78440 11060 78450
rect 11190 78440 11310 78450
rect 11440 78440 11560 78450
rect 11690 78440 11810 78450
rect 11940 78440 12060 78450
rect 12190 78440 12310 78450
rect 12440 78440 12560 78450
rect 12690 78440 12810 78450
rect 12940 78440 13060 78450
rect 13190 78440 13310 78450
rect 13440 78440 13560 78450
rect 13690 78440 13810 78450
rect 13940 78440 14060 78450
rect 14190 78440 14310 78450
rect 14440 78440 14560 78450
rect 14690 78440 14810 78450
rect 14940 78440 15060 78450
rect 15190 78440 15310 78450
rect 15440 78440 15560 78450
rect 15690 78440 15810 78450
rect 15940 78440 16060 78450
rect 16190 78440 16310 78450
rect 16440 78440 16560 78450
rect 16690 78440 16810 78450
rect 16940 78440 17060 78450
rect 17190 78440 17310 78450
rect 17440 78440 17560 78450
rect 17690 78440 17810 78450
rect 17940 78440 18060 78450
rect 18190 78440 18310 78450
rect 18440 78440 18560 78450
rect 18690 78440 18810 78450
rect 18940 78440 19060 78450
rect 19190 78440 19310 78450
rect 19440 78440 19560 78450
rect 19690 78440 19810 78450
rect 19940 78440 20060 78450
rect 20190 78440 20310 78450
rect 20440 78440 20560 78450
rect 20690 78440 20810 78450
rect 20940 78440 21060 78450
rect 21190 78440 21310 78450
rect 21440 78440 21560 78450
rect 21690 78440 21810 78450
rect 21940 78440 22060 78450
rect 22190 78440 22310 78450
rect 22440 78440 22560 78450
rect 22690 78440 22810 78450
rect 22940 78440 23060 78450
rect 23190 78440 23310 78450
rect 23440 78440 23560 78450
rect 23690 78440 23810 78450
rect 23940 78440 24060 78450
rect 24190 78440 24310 78450
rect 24440 78440 24560 78450
rect 24690 78440 24810 78450
rect 24940 78440 25060 78450
rect 25190 78440 25310 78450
rect 25440 78440 25560 78450
rect 25690 78440 25810 78450
rect 25940 78440 26060 78450
rect 26190 78440 26310 78450
rect 26440 78440 26560 78450
rect 26690 78440 26810 78450
rect 26940 78440 27060 78450
rect 27190 78440 27310 78450
rect 27440 78440 27560 78450
rect 27690 78440 27810 78450
rect 27940 78440 28060 78450
rect 28190 78440 28310 78450
rect 28440 78440 28560 78450
rect 28690 78440 28810 78450
rect 28940 78440 29000 78450
rect 7000 78310 7050 78440
rect 7200 78310 7300 78440
rect 7450 78310 7550 78440
rect 7700 78310 7800 78440
rect 7950 78310 8050 78440
rect 8200 78310 8300 78440
rect 8450 78310 8550 78440
rect 8700 78310 8800 78440
rect 8950 78310 9050 78440
rect 9200 78310 9300 78440
rect 9450 78310 9550 78440
rect 9700 78310 9800 78440
rect 9950 78310 10050 78440
rect 10200 78310 10300 78440
rect 10450 78310 10550 78440
rect 10700 78310 10800 78440
rect 10950 78310 11050 78440
rect 11200 78310 11300 78440
rect 11450 78310 11550 78440
rect 11700 78310 11800 78440
rect 11950 78310 12050 78440
rect 12200 78310 12300 78440
rect 12450 78310 12550 78440
rect 12700 78310 12800 78440
rect 12950 78310 13050 78440
rect 13200 78310 13300 78440
rect 13450 78310 13550 78440
rect 13700 78310 13800 78440
rect 13950 78310 14050 78440
rect 14200 78310 14300 78440
rect 14450 78310 14550 78440
rect 14700 78310 14800 78440
rect 14950 78310 15050 78440
rect 15200 78310 15300 78440
rect 15450 78310 15550 78440
rect 15700 78310 15800 78440
rect 15950 78310 16050 78440
rect 16200 78310 16300 78440
rect 16450 78310 16550 78440
rect 16700 78310 16800 78440
rect 16950 78310 17050 78440
rect 17200 78310 17300 78440
rect 17450 78310 17550 78440
rect 17700 78310 17800 78440
rect 17950 78310 18050 78440
rect 18200 78310 18300 78440
rect 18450 78310 18550 78440
rect 18700 78310 18800 78440
rect 18950 78310 19050 78440
rect 19200 78310 19300 78440
rect 19450 78310 19550 78440
rect 19700 78310 19800 78440
rect 19950 78310 20050 78440
rect 20200 78310 20300 78440
rect 20450 78310 20550 78440
rect 20700 78310 20800 78440
rect 20950 78310 21050 78440
rect 21200 78310 21300 78440
rect 21450 78310 21550 78440
rect 21700 78310 21800 78440
rect 21950 78310 22050 78440
rect 22200 78310 22300 78440
rect 22450 78310 22550 78440
rect 22700 78310 22800 78440
rect 22950 78310 23050 78440
rect 23200 78310 23300 78440
rect 23450 78310 23550 78440
rect 23700 78310 23800 78440
rect 23950 78310 24050 78440
rect 24200 78310 24300 78440
rect 24450 78310 24550 78440
rect 24700 78310 24800 78440
rect 24950 78310 25050 78440
rect 25200 78310 25300 78440
rect 25450 78310 25550 78440
rect 25700 78310 25800 78440
rect 25950 78310 26050 78440
rect 26200 78310 26300 78440
rect 26450 78310 26550 78440
rect 26700 78310 26800 78440
rect 26950 78310 27050 78440
rect 27200 78310 27300 78440
rect 27450 78310 27550 78440
rect 27700 78310 27800 78440
rect 27950 78310 28050 78440
rect 28200 78310 28300 78440
rect 28450 78310 28550 78440
rect 28700 78310 28800 78440
rect 28950 78310 29000 78440
rect 7000 78300 7060 78310
rect 7190 78300 7310 78310
rect 7440 78300 7560 78310
rect 7690 78300 7810 78310
rect 7940 78300 8060 78310
rect 8190 78300 8310 78310
rect 8440 78300 8560 78310
rect 8690 78300 8810 78310
rect 8940 78300 9060 78310
rect 9190 78300 9310 78310
rect 9440 78300 9560 78310
rect 9690 78300 9810 78310
rect 9940 78300 10060 78310
rect 10190 78300 10310 78310
rect 10440 78300 10560 78310
rect 10690 78300 10810 78310
rect 10940 78300 11060 78310
rect 11190 78300 11310 78310
rect 11440 78300 11560 78310
rect 11690 78300 11810 78310
rect 11940 78300 12060 78310
rect 12190 78300 12310 78310
rect 12440 78300 12560 78310
rect 12690 78300 12810 78310
rect 12940 78300 13060 78310
rect 13190 78300 13310 78310
rect 13440 78300 13560 78310
rect 13690 78300 13810 78310
rect 13940 78300 14060 78310
rect 14190 78300 14310 78310
rect 14440 78300 14560 78310
rect 14690 78300 14810 78310
rect 14940 78300 15060 78310
rect 15190 78300 15310 78310
rect 15440 78300 15560 78310
rect 15690 78300 15810 78310
rect 15940 78300 16060 78310
rect 16190 78300 16310 78310
rect 16440 78300 16560 78310
rect 16690 78300 16810 78310
rect 16940 78300 17060 78310
rect 17190 78300 17310 78310
rect 17440 78300 17560 78310
rect 17690 78300 17810 78310
rect 17940 78300 18060 78310
rect 18190 78300 18310 78310
rect 18440 78300 18560 78310
rect 18690 78300 18810 78310
rect 18940 78300 19060 78310
rect 19190 78300 19310 78310
rect 19440 78300 19560 78310
rect 19690 78300 19810 78310
rect 19940 78300 20060 78310
rect 20190 78300 20310 78310
rect 20440 78300 20560 78310
rect 20690 78300 20810 78310
rect 20940 78300 21060 78310
rect 21190 78300 21310 78310
rect 21440 78300 21560 78310
rect 21690 78300 21810 78310
rect 21940 78300 22060 78310
rect 22190 78300 22310 78310
rect 22440 78300 22560 78310
rect 22690 78300 22810 78310
rect 22940 78300 23060 78310
rect 23190 78300 23310 78310
rect 23440 78300 23560 78310
rect 23690 78300 23810 78310
rect 23940 78300 24060 78310
rect 24190 78300 24310 78310
rect 24440 78300 24560 78310
rect 24690 78300 24810 78310
rect 24940 78300 25060 78310
rect 25190 78300 25310 78310
rect 25440 78300 25560 78310
rect 25690 78300 25810 78310
rect 25940 78300 26060 78310
rect 26190 78300 26310 78310
rect 26440 78300 26560 78310
rect 26690 78300 26810 78310
rect 26940 78300 27060 78310
rect 27190 78300 27310 78310
rect 27440 78300 27560 78310
rect 27690 78300 27810 78310
rect 27940 78300 28060 78310
rect 28190 78300 28310 78310
rect 28440 78300 28560 78310
rect 28690 78300 28810 78310
rect 28940 78300 29000 78310
rect 7000 78200 29000 78300
rect 7000 78190 7060 78200
rect 7190 78190 7310 78200
rect 7440 78190 7560 78200
rect 7690 78190 7810 78200
rect 7940 78190 8060 78200
rect 8190 78190 8310 78200
rect 8440 78190 8560 78200
rect 8690 78190 8810 78200
rect 8940 78190 9060 78200
rect 9190 78190 9310 78200
rect 9440 78190 9560 78200
rect 9690 78190 9810 78200
rect 9940 78190 10060 78200
rect 10190 78190 10310 78200
rect 10440 78190 10560 78200
rect 10690 78190 10810 78200
rect 10940 78190 11060 78200
rect 11190 78190 11310 78200
rect 11440 78190 11560 78200
rect 11690 78190 11810 78200
rect 11940 78190 12060 78200
rect 12190 78190 12310 78200
rect 12440 78190 12560 78200
rect 12690 78190 12810 78200
rect 12940 78190 13060 78200
rect 13190 78190 13310 78200
rect 13440 78190 13560 78200
rect 13690 78190 13810 78200
rect 13940 78190 14060 78200
rect 14190 78190 14310 78200
rect 14440 78190 14560 78200
rect 14690 78190 14810 78200
rect 14940 78190 15060 78200
rect 15190 78190 15310 78200
rect 15440 78190 15560 78200
rect 15690 78190 15810 78200
rect 15940 78190 16060 78200
rect 16190 78190 16310 78200
rect 16440 78190 16560 78200
rect 16690 78190 16810 78200
rect 16940 78190 17060 78200
rect 17190 78190 17310 78200
rect 17440 78190 17560 78200
rect 17690 78190 17810 78200
rect 17940 78190 18060 78200
rect 18190 78190 18310 78200
rect 18440 78190 18560 78200
rect 18690 78190 18810 78200
rect 18940 78190 19060 78200
rect 19190 78190 19310 78200
rect 19440 78190 19560 78200
rect 19690 78190 19810 78200
rect 19940 78190 20060 78200
rect 20190 78190 20310 78200
rect 20440 78190 20560 78200
rect 20690 78190 20810 78200
rect 20940 78190 21060 78200
rect 21190 78190 21310 78200
rect 21440 78190 21560 78200
rect 21690 78190 21810 78200
rect 21940 78190 22060 78200
rect 22190 78190 22310 78200
rect 22440 78190 22560 78200
rect 22690 78190 22810 78200
rect 22940 78190 23060 78200
rect 23190 78190 23310 78200
rect 23440 78190 23560 78200
rect 23690 78190 23810 78200
rect 23940 78190 24060 78200
rect 24190 78190 24310 78200
rect 24440 78190 24560 78200
rect 24690 78190 24810 78200
rect 24940 78190 25060 78200
rect 25190 78190 25310 78200
rect 25440 78190 25560 78200
rect 25690 78190 25810 78200
rect 25940 78190 26060 78200
rect 26190 78190 26310 78200
rect 26440 78190 26560 78200
rect 26690 78190 26810 78200
rect 26940 78190 27060 78200
rect 27190 78190 27310 78200
rect 27440 78190 27560 78200
rect 27690 78190 27810 78200
rect 27940 78190 28060 78200
rect 28190 78190 28310 78200
rect 28440 78190 28560 78200
rect 28690 78190 28810 78200
rect 28940 78190 29000 78200
rect 7000 78060 7050 78190
rect 7200 78060 7300 78190
rect 7450 78060 7550 78190
rect 7700 78060 7800 78190
rect 7950 78060 8050 78190
rect 8200 78060 8300 78190
rect 8450 78060 8550 78190
rect 8700 78060 8800 78190
rect 8950 78060 9050 78190
rect 9200 78060 9300 78190
rect 9450 78060 9550 78190
rect 9700 78060 9800 78190
rect 9950 78060 10050 78190
rect 10200 78060 10300 78190
rect 10450 78060 10550 78190
rect 10700 78060 10800 78190
rect 10950 78060 11050 78190
rect 11200 78060 11300 78190
rect 11450 78060 11550 78190
rect 11700 78060 11800 78190
rect 11950 78060 12050 78190
rect 12200 78060 12300 78190
rect 12450 78060 12550 78190
rect 12700 78060 12800 78190
rect 12950 78060 13050 78190
rect 13200 78060 13300 78190
rect 13450 78060 13550 78190
rect 13700 78060 13800 78190
rect 13950 78060 14050 78190
rect 14200 78060 14300 78190
rect 14450 78060 14550 78190
rect 14700 78060 14800 78190
rect 14950 78060 15050 78190
rect 15200 78060 15300 78190
rect 15450 78060 15550 78190
rect 15700 78060 15800 78190
rect 15950 78060 16050 78190
rect 16200 78060 16300 78190
rect 16450 78060 16550 78190
rect 16700 78060 16800 78190
rect 16950 78060 17050 78190
rect 17200 78060 17300 78190
rect 17450 78060 17550 78190
rect 17700 78060 17800 78190
rect 17950 78060 18050 78190
rect 18200 78060 18300 78190
rect 18450 78060 18550 78190
rect 18700 78060 18800 78190
rect 18950 78060 19050 78190
rect 19200 78060 19300 78190
rect 19450 78060 19550 78190
rect 19700 78060 19800 78190
rect 19950 78060 20050 78190
rect 20200 78060 20300 78190
rect 20450 78060 20550 78190
rect 20700 78060 20800 78190
rect 20950 78060 21050 78190
rect 21200 78060 21300 78190
rect 21450 78060 21550 78190
rect 21700 78060 21800 78190
rect 21950 78060 22050 78190
rect 22200 78060 22300 78190
rect 22450 78060 22550 78190
rect 22700 78060 22800 78190
rect 22950 78060 23050 78190
rect 23200 78060 23300 78190
rect 23450 78060 23550 78190
rect 23700 78060 23800 78190
rect 23950 78060 24050 78190
rect 24200 78060 24300 78190
rect 24450 78060 24550 78190
rect 24700 78060 24800 78190
rect 24950 78060 25050 78190
rect 25200 78060 25300 78190
rect 25450 78060 25550 78190
rect 25700 78060 25800 78190
rect 25950 78060 26050 78190
rect 26200 78060 26300 78190
rect 26450 78060 26550 78190
rect 26700 78060 26800 78190
rect 26950 78060 27050 78190
rect 27200 78060 27300 78190
rect 27450 78060 27550 78190
rect 27700 78060 27800 78190
rect 27950 78060 28050 78190
rect 28200 78060 28300 78190
rect 28450 78060 28550 78190
rect 28700 78060 28800 78190
rect 28950 78060 29000 78190
rect 7000 78050 7060 78060
rect 7190 78050 7310 78060
rect 7440 78050 7560 78060
rect 7690 78050 7810 78060
rect 7940 78050 8060 78060
rect 8190 78050 8310 78060
rect 8440 78050 8560 78060
rect 8690 78050 8810 78060
rect 8940 78050 9060 78060
rect 9190 78050 9310 78060
rect 9440 78050 9560 78060
rect 9690 78050 9810 78060
rect 9940 78050 10060 78060
rect 10190 78050 10310 78060
rect 10440 78050 10560 78060
rect 10690 78050 10810 78060
rect 10940 78050 11060 78060
rect 11190 78050 11310 78060
rect 11440 78050 11560 78060
rect 11690 78050 11810 78060
rect 11940 78050 12060 78060
rect 12190 78050 12310 78060
rect 12440 78050 12560 78060
rect 12690 78050 12810 78060
rect 12940 78050 13060 78060
rect 13190 78050 13310 78060
rect 13440 78050 13560 78060
rect 13690 78050 13810 78060
rect 13940 78050 14060 78060
rect 14190 78050 14310 78060
rect 14440 78050 14560 78060
rect 14690 78050 14810 78060
rect 14940 78050 15060 78060
rect 15190 78050 15310 78060
rect 15440 78050 15560 78060
rect 15690 78050 15810 78060
rect 15940 78050 16060 78060
rect 16190 78050 16310 78060
rect 16440 78050 16560 78060
rect 16690 78050 16810 78060
rect 16940 78050 17060 78060
rect 17190 78050 17310 78060
rect 17440 78050 17560 78060
rect 17690 78050 17810 78060
rect 17940 78050 18060 78060
rect 18190 78050 18310 78060
rect 18440 78050 18560 78060
rect 18690 78050 18810 78060
rect 18940 78050 19060 78060
rect 19190 78050 19310 78060
rect 19440 78050 19560 78060
rect 19690 78050 19810 78060
rect 19940 78050 20060 78060
rect 20190 78050 20310 78060
rect 20440 78050 20560 78060
rect 20690 78050 20810 78060
rect 20940 78050 21060 78060
rect 21190 78050 21310 78060
rect 21440 78050 21560 78060
rect 21690 78050 21810 78060
rect 21940 78050 22060 78060
rect 22190 78050 22310 78060
rect 22440 78050 22560 78060
rect 22690 78050 22810 78060
rect 22940 78050 23060 78060
rect 23190 78050 23310 78060
rect 23440 78050 23560 78060
rect 23690 78050 23810 78060
rect 23940 78050 24060 78060
rect 24190 78050 24310 78060
rect 24440 78050 24560 78060
rect 24690 78050 24810 78060
rect 24940 78050 25060 78060
rect 25190 78050 25310 78060
rect 25440 78050 25560 78060
rect 25690 78050 25810 78060
rect 25940 78050 26060 78060
rect 26190 78050 26310 78060
rect 26440 78050 26560 78060
rect 26690 78050 26810 78060
rect 26940 78050 27060 78060
rect 27190 78050 27310 78060
rect 27440 78050 27560 78060
rect 27690 78050 27810 78060
rect 27940 78050 28060 78060
rect 28190 78050 28310 78060
rect 28440 78050 28560 78060
rect 28690 78050 28810 78060
rect 28940 78050 29000 78060
rect 7000 77950 29000 78050
rect 7000 77940 7060 77950
rect 7190 77940 7310 77950
rect 7440 77940 7560 77950
rect 7690 77940 7810 77950
rect 7940 77940 8060 77950
rect 8190 77940 8310 77950
rect 8440 77940 8560 77950
rect 8690 77940 8810 77950
rect 8940 77940 9060 77950
rect 9190 77940 9310 77950
rect 9440 77940 9560 77950
rect 9690 77940 9810 77950
rect 9940 77940 10060 77950
rect 10190 77940 10310 77950
rect 10440 77940 10560 77950
rect 10690 77940 10810 77950
rect 10940 77940 11060 77950
rect 11190 77940 11310 77950
rect 11440 77940 11560 77950
rect 11690 77940 11810 77950
rect 11940 77940 12060 77950
rect 12190 77940 12310 77950
rect 12440 77940 12560 77950
rect 12690 77940 12810 77950
rect 12940 77940 13060 77950
rect 13190 77940 13310 77950
rect 13440 77940 13560 77950
rect 13690 77940 13810 77950
rect 13940 77940 14060 77950
rect 14190 77940 14310 77950
rect 14440 77940 14560 77950
rect 14690 77940 14810 77950
rect 14940 77940 15060 77950
rect 15190 77940 15310 77950
rect 15440 77940 15560 77950
rect 15690 77940 15810 77950
rect 15940 77940 16060 77950
rect 16190 77940 16310 77950
rect 16440 77940 16560 77950
rect 16690 77940 16810 77950
rect 16940 77940 17060 77950
rect 17190 77940 17310 77950
rect 17440 77940 17560 77950
rect 17690 77940 17810 77950
rect 17940 77940 18060 77950
rect 18190 77940 18310 77950
rect 18440 77940 18560 77950
rect 18690 77940 18810 77950
rect 18940 77940 19060 77950
rect 19190 77940 19310 77950
rect 19440 77940 19560 77950
rect 19690 77940 19810 77950
rect 19940 77940 20060 77950
rect 20190 77940 20310 77950
rect 20440 77940 20560 77950
rect 20690 77940 20810 77950
rect 20940 77940 21060 77950
rect 21190 77940 21310 77950
rect 21440 77940 21560 77950
rect 21690 77940 21810 77950
rect 21940 77940 22060 77950
rect 22190 77940 22310 77950
rect 22440 77940 22560 77950
rect 22690 77940 22810 77950
rect 22940 77940 23060 77950
rect 23190 77940 23310 77950
rect 23440 77940 23560 77950
rect 23690 77940 23810 77950
rect 23940 77940 24060 77950
rect 24190 77940 24310 77950
rect 24440 77940 24560 77950
rect 24690 77940 24810 77950
rect 24940 77940 25060 77950
rect 25190 77940 25310 77950
rect 25440 77940 25560 77950
rect 25690 77940 25810 77950
rect 25940 77940 26060 77950
rect 26190 77940 26310 77950
rect 26440 77940 26560 77950
rect 26690 77940 26810 77950
rect 26940 77940 27060 77950
rect 27190 77940 27310 77950
rect 27440 77940 27560 77950
rect 27690 77940 27810 77950
rect 27940 77940 28060 77950
rect 28190 77940 28310 77950
rect 28440 77940 28560 77950
rect 28690 77940 28810 77950
rect 28940 77940 29000 77950
rect 7000 77810 7050 77940
rect 7200 77810 7300 77940
rect 7450 77810 7550 77940
rect 7700 77810 7800 77940
rect 7950 77810 8050 77940
rect 8200 77810 8300 77940
rect 8450 77810 8550 77940
rect 8700 77810 8800 77940
rect 8950 77810 9050 77940
rect 9200 77810 9300 77940
rect 9450 77810 9550 77940
rect 9700 77810 9800 77940
rect 9950 77810 10050 77940
rect 10200 77810 10300 77940
rect 10450 77810 10550 77940
rect 10700 77810 10800 77940
rect 10950 77810 11050 77940
rect 11200 77810 11300 77940
rect 11450 77810 11550 77940
rect 11700 77810 11800 77940
rect 11950 77810 12050 77940
rect 12200 77810 12300 77940
rect 12450 77810 12550 77940
rect 12700 77810 12800 77940
rect 12950 77810 13050 77940
rect 13200 77810 13300 77940
rect 13450 77810 13550 77940
rect 13700 77810 13800 77940
rect 13950 77810 14050 77940
rect 14200 77810 14300 77940
rect 14450 77810 14550 77940
rect 14700 77810 14800 77940
rect 14950 77810 15050 77940
rect 15200 77810 15300 77940
rect 15450 77810 15550 77940
rect 15700 77810 15800 77940
rect 15950 77810 16050 77940
rect 16200 77810 16300 77940
rect 16450 77810 16550 77940
rect 16700 77810 16800 77940
rect 16950 77810 17050 77940
rect 17200 77810 17300 77940
rect 17450 77810 17550 77940
rect 17700 77810 17800 77940
rect 17950 77810 18050 77940
rect 18200 77810 18300 77940
rect 18450 77810 18550 77940
rect 18700 77810 18800 77940
rect 18950 77810 19050 77940
rect 19200 77810 19300 77940
rect 19450 77810 19550 77940
rect 19700 77810 19800 77940
rect 19950 77810 20050 77940
rect 20200 77810 20300 77940
rect 20450 77810 20550 77940
rect 20700 77810 20800 77940
rect 20950 77810 21050 77940
rect 21200 77810 21300 77940
rect 21450 77810 21550 77940
rect 21700 77810 21800 77940
rect 21950 77810 22050 77940
rect 22200 77810 22300 77940
rect 22450 77810 22550 77940
rect 22700 77810 22800 77940
rect 22950 77810 23050 77940
rect 23200 77810 23300 77940
rect 23450 77810 23550 77940
rect 23700 77810 23800 77940
rect 23950 77810 24050 77940
rect 24200 77810 24300 77940
rect 24450 77810 24550 77940
rect 24700 77810 24800 77940
rect 24950 77810 25050 77940
rect 25200 77810 25300 77940
rect 25450 77810 25550 77940
rect 25700 77810 25800 77940
rect 25950 77810 26050 77940
rect 26200 77810 26300 77940
rect 26450 77810 26550 77940
rect 26700 77810 26800 77940
rect 26950 77810 27050 77940
rect 27200 77810 27300 77940
rect 27450 77810 27550 77940
rect 27700 77810 27800 77940
rect 27950 77810 28050 77940
rect 28200 77810 28300 77940
rect 28450 77810 28550 77940
rect 28700 77810 28800 77940
rect 28950 77810 29000 77940
rect 7000 77800 7060 77810
rect 7190 77800 7310 77810
rect 7440 77800 7560 77810
rect 7690 77800 7810 77810
rect 7940 77800 8060 77810
rect 8190 77800 8310 77810
rect 8440 77800 8560 77810
rect 8690 77800 8810 77810
rect 8940 77800 9060 77810
rect 9190 77800 9310 77810
rect 9440 77800 9560 77810
rect 9690 77800 9810 77810
rect 9940 77800 10060 77810
rect 10190 77800 10310 77810
rect 10440 77800 10560 77810
rect 10690 77800 10810 77810
rect 10940 77800 11060 77810
rect 11190 77800 11310 77810
rect 11440 77800 11560 77810
rect 11690 77800 11810 77810
rect 11940 77800 12060 77810
rect 12190 77800 12310 77810
rect 12440 77800 12560 77810
rect 12690 77800 12810 77810
rect 12940 77800 13060 77810
rect 13190 77800 13310 77810
rect 13440 77800 13560 77810
rect 13690 77800 13810 77810
rect 13940 77800 14060 77810
rect 14190 77800 14310 77810
rect 14440 77800 14560 77810
rect 14690 77800 14810 77810
rect 14940 77800 15060 77810
rect 15190 77800 15310 77810
rect 15440 77800 15560 77810
rect 15690 77800 15810 77810
rect 15940 77800 16060 77810
rect 16190 77800 16310 77810
rect 16440 77800 16560 77810
rect 16690 77800 16810 77810
rect 16940 77800 17060 77810
rect 17190 77800 17310 77810
rect 17440 77800 17560 77810
rect 17690 77800 17810 77810
rect 17940 77800 18060 77810
rect 18190 77800 18310 77810
rect 18440 77800 18560 77810
rect 18690 77800 18810 77810
rect 18940 77800 19060 77810
rect 19190 77800 19310 77810
rect 19440 77800 19560 77810
rect 19690 77800 19810 77810
rect 19940 77800 20060 77810
rect 20190 77800 20310 77810
rect 20440 77800 20560 77810
rect 20690 77800 20810 77810
rect 20940 77800 21060 77810
rect 21190 77800 21310 77810
rect 21440 77800 21560 77810
rect 21690 77800 21810 77810
rect 21940 77800 22060 77810
rect 22190 77800 22310 77810
rect 22440 77800 22560 77810
rect 22690 77800 22810 77810
rect 22940 77800 23060 77810
rect 23190 77800 23310 77810
rect 23440 77800 23560 77810
rect 23690 77800 23810 77810
rect 23940 77800 24060 77810
rect 24190 77800 24310 77810
rect 24440 77800 24560 77810
rect 24690 77800 24810 77810
rect 24940 77800 25060 77810
rect 25190 77800 25310 77810
rect 25440 77800 25560 77810
rect 25690 77800 25810 77810
rect 25940 77800 26060 77810
rect 26190 77800 26310 77810
rect 26440 77800 26560 77810
rect 26690 77800 26810 77810
rect 26940 77800 27060 77810
rect 27190 77800 27310 77810
rect 27440 77800 27560 77810
rect 27690 77800 27810 77810
rect 27940 77800 28060 77810
rect 28190 77800 28310 77810
rect 28440 77800 28560 77810
rect 28690 77800 28810 77810
rect 28940 77800 29000 77810
rect 7000 77700 29000 77800
rect 7000 77690 7060 77700
rect 7190 77690 7310 77700
rect 7440 77690 7560 77700
rect 7690 77690 7810 77700
rect 7940 77690 8060 77700
rect 8190 77690 8310 77700
rect 8440 77690 8560 77700
rect 8690 77690 8810 77700
rect 8940 77690 9060 77700
rect 9190 77690 9310 77700
rect 9440 77690 9560 77700
rect 9690 77690 9810 77700
rect 9940 77690 10060 77700
rect 10190 77690 10310 77700
rect 10440 77690 10560 77700
rect 10690 77690 10810 77700
rect 10940 77690 11060 77700
rect 11190 77690 11310 77700
rect 11440 77690 11560 77700
rect 11690 77690 11810 77700
rect 11940 77690 12060 77700
rect 12190 77690 12310 77700
rect 12440 77690 12560 77700
rect 12690 77690 12810 77700
rect 12940 77690 13060 77700
rect 13190 77690 13310 77700
rect 13440 77690 13560 77700
rect 13690 77690 13810 77700
rect 13940 77690 14060 77700
rect 14190 77690 14310 77700
rect 14440 77690 14560 77700
rect 14690 77690 14810 77700
rect 14940 77690 15060 77700
rect 15190 77690 15310 77700
rect 15440 77690 15560 77700
rect 15690 77690 15810 77700
rect 15940 77690 16060 77700
rect 16190 77690 16310 77700
rect 16440 77690 16560 77700
rect 16690 77690 16810 77700
rect 16940 77690 17060 77700
rect 17190 77690 17310 77700
rect 17440 77690 17560 77700
rect 17690 77690 17810 77700
rect 17940 77690 18060 77700
rect 18190 77690 18310 77700
rect 18440 77690 18560 77700
rect 18690 77690 18810 77700
rect 18940 77690 19060 77700
rect 19190 77690 19310 77700
rect 19440 77690 19560 77700
rect 19690 77690 19810 77700
rect 19940 77690 20060 77700
rect 20190 77690 20310 77700
rect 20440 77690 20560 77700
rect 20690 77690 20810 77700
rect 20940 77690 21060 77700
rect 21190 77690 21310 77700
rect 21440 77690 21560 77700
rect 21690 77690 21810 77700
rect 21940 77690 22060 77700
rect 22190 77690 22310 77700
rect 22440 77690 22560 77700
rect 22690 77690 22810 77700
rect 22940 77690 23060 77700
rect 23190 77690 23310 77700
rect 23440 77690 23560 77700
rect 23690 77690 23810 77700
rect 23940 77690 24060 77700
rect 24190 77690 24310 77700
rect 24440 77690 24560 77700
rect 24690 77690 24810 77700
rect 24940 77690 25060 77700
rect 25190 77690 25310 77700
rect 25440 77690 25560 77700
rect 25690 77690 25810 77700
rect 25940 77690 26060 77700
rect 26190 77690 26310 77700
rect 26440 77690 26560 77700
rect 26690 77690 26810 77700
rect 26940 77690 27060 77700
rect 27190 77690 27310 77700
rect 27440 77690 27560 77700
rect 27690 77690 27810 77700
rect 27940 77690 28060 77700
rect 28190 77690 28310 77700
rect 28440 77690 28560 77700
rect 28690 77690 28810 77700
rect 28940 77690 29000 77700
rect 7000 77560 7050 77690
rect 7200 77560 7300 77690
rect 7450 77560 7550 77690
rect 7700 77560 7800 77690
rect 7950 77560 8050 77690
rect 8200 77560 8300 77690
rect 8450 77560 8550 77690
rect 8700 77560 8800 77690
rect 8950 77560 9050 77690
rect 9200 77560 9300 77690
rect 9450 77560 9550 77690
rect 9700 77560 9800 77690
rect 9950 77560 10050 77690
rect 10200 77560 10300 77690
rect 10450 77560 10550 77690
rect 10700 77560 10800 77690
rect 10950 77560 11050 77690
rect 11200 77560 11300 77690
rect 11450 77560 11550 77690
rect 11700 77560 11800 77690
rect 11950 77560 12050 77690
rect 12200 77560 12300 77690
rect 12450 77560 12550 77690
rect 12700 77560 12800 77690
rect 12950 77560 13050 77690
rect 13200 77560 13300 77690
rect 13450 77560 13550 77690
rect 13700 77560 13800 77690
rect 13950 77560 14050 77690
rect 14200 77560 14300 77690
rect 14450 77560 14550 77690
rect 14700 77560 14800 77690
rect 14950 77560 15050 77690
rect 15200 77560 15300 77690
rect 15450 77560 15550 77690
rect 15700 77560 15800 77690
rect 15950 77560 16050 77690
rect 16200 77560 16300 77690
rect 16450 77560 16550 77690
rect 16700 77560 16800 77690
rect 16950 77560 17050 77690
rect 17200 77560 17300 77690
rect 17450 77560 17550 77690
rect 17700 77560 17800 77690
rect 17950 77560 18050 77690
rect 18200 77560 18300 77690
rect 18450 77560 18550 77690
rect 18700 77560 18800 77690
rect 18950 77560 19050 77690
rect 19200 77560 19300 77690
rect 19450 77560 19550 77690
rect 19700 77560 19800 77690
rect 19950 77560 20050 77690
rect 20200 77560 20300 77690
rect 20450 77560 20550 77690
rect 20700 77560 20800 77690
rect 20950 77560 21050 77690
rect 21200 77560 21300 77690
rect 21450 77560 21550 77690
rect 21700 77560 21800 77690
rect 21950 77560 22050 77690
rect 22200 77560 22300 77690
rect 22450 77560 22550 77690
rect 22700 77560 22800 77690
rect 22950 77560 23050 77690
rect 23200 77560 23300 77690
rect 23450 77560 23550 77690
rect 23700 77560 23800 77690
rect 23950 77560 24050 77690
rect 24200 77560 24300 77690
rect 24450 77560 24550 77690
rect 24700 77560 24800 77690
rect 24950 77560 25050 77690
rect 25200 77560 25300 77690
rect 25450 77560 25550 77690
rect 25700 77560 25800 77690
rect 25950 77560 26050 77690
rect 26200 77560 26300 77690
rect 26450 77560 26550 77690
rect 26700 77560 26800 77690
rect 26950 77560 27050 77690
rect 27200 77560 27300 77690
rect 27450 77560 27550 77690
rect 27700 77560 27800 77690
rect 27950 77560 28050 77690
rect 28200 77560 28300 77690
rect 28450 77560 28550 77690
rect 28700 77560 28800 77690
rect 28950 77560 29000 77690
rect 7000 77550 7060 77560
rect 7190 77550 7310 77560
rect 7440 77550 7560 77560
rect 7690 77550 7810 77560
rect 7940 77550 8060 77560
rect 8190 77550 8310 77560
rect 8440 77550 8560 77560
rect 8690 77550 8810 77560
rect 8940 77550 9060 77560
rect 9190 77550 9310 77560
rect 9440 77550 9560 77560
rect 9690 77550 9810 77560
rect 9940 77550 10060 77560
rect 10190 77550 10310 77560
rect 10440 77550 10560 77560
rect 10690 77550 10810 77560
rect 10940 77550 11060 77560
rect 11190 77550 11310 77560
rect 11440 77550 11560 77560
rect 11690 77550 11810 77560
rect 11940 77550 12060 77560
rect 12190 77550 12310 77560
rect 12440 77550 12560 77560
rect 12690 77550 12810 77560
rect 12940 77550 13060 77560
rect 13190 77550 13310 77560
rect 13440 77550 13560 77560
rect 13690 77550 13810 77560
rect 13940 77550 14060 77560
rect 14190 77550 14310 77560
rect 14440 77550 14560 77560
rect 14690 77550 14810 77560
rect 14940 77550 15060 77560
rect 15190 77550 15310 77560
rect 15440 77550 15560 77560
rect 15690 77550 15810 77560
rect 15940 77550 16060 77560
rect 16190 77550 16310 77560
rect 16440 77550 16560 77560
rect 16690 77550 16810 77560
rect 16940 77550 17060 77560
rect 17190 77550 17310 77560
rect 17440 77550 17560 77560
rect 17690 77550 17810 77560
rect 17940 77550 18060 77560
rect 18190 77550 18310 77560
rect 18440 77550 18560 77560
rect 18690 77550 18810 77560
rect 18940 77550 19060 77560
rect 19190 77550 19310 77560
rect 19440 77550 19560 77560
rect 19690 77550 19810 77560
rect 19940 77550 20060 77560
rect 20190 77550 20310 77560
rect 20440 77550 20560 77560
rect 20690 77550 20810 77560
rect 20940 77550 21060 77560
rect 21190 77550 21310 77560
rect 21440 77550 21560 77560
rect 21690 77550 21810 77560
rect 21940 77550 22060 77560
rect 22190 77550 22310 77560
rect 22440 77550 22560 77560
rect 22690 77550 22810 77560
rect 22940 77550 23060 77560
rect 23190 77550 23310 77560
rect 23440 77550 23560 77560
rect 23690 77550 23810 77560
rect 23940 77550 24060 77560
rect 24190 77550 24310 77560
rect 24440 77550 24560 77560
rect 24690 77550 24810 77560
rect 24940 77550 25060 77560
rect 25190 77550 25310 77560
rect 25440 77550 25560 77560
rect 25690 77550 25810 77560
rect 25940 77550 26060 77560
rect 26190 77550 26310 77560
rect 26440 77550 26560 77560
rect 26690 77550 26810 77560
rect 26940 77550 27060 77560
rect 27190 77550 27310 77560
rect 27440 77550 27560 77560
rect 27690 77550 27810 77560
rect 27940 77550 28060 77560
rect 28190 77550 28310 77560
rect 28440 77550 28560 77560
rect 28690 77550 28810 77560
rect 28940 77550 29000 77560
rect 7000 77450 29000 77550
rect 7000 77440 7060 77450
rect 7190 77440 7310 77450
rect 7440 77440 7560 77450
rect 7690 77440 7810 77450
rect 7940 77440 8060 77450
rect 8190 77440 8310 77450
rect 8440 77440 8560 77450
rect 8690 77440 8810 77450
rect 8940 77440 9060 77450
rect 9190 77440 9310 77450
rect 9440 77440 9560 77450
rect 9690 77440 9810 77450
rect 9940 77440 10060 77450
rect 10190 77440 10310 77450
rect 10440 77440 10560 77450
rect 10690 77440 10810 77450
rect 10940 77440 11060 77450
rect 11190 77440 11310 77450
rect 11440 77440 11560 77450
rect 11690 77440 11810 77450
rect 11940 77440 12060 77450
rect 12190 77440 12310 77450
rect 12440 77440 12560 77450
rect 12690 77440 12810 77450
rect 12940 77440 13060 77450
rect 13190 77440 13310 77450
rect 13440 77440 13560 77450
rect 13690 77440 13810 77450
rect 13940 77440 14060 77450
rect 14190 77440 14310 77450
rect 14440 77440 14560 77450
rect 14690 77440 14810 77450
rect 14940 77440 15060 77450
rect 15190 77440 15310 77450
rect 15440 77440 15560 77450
rect 15690 77440 15810 77450
rect 15940 77440 16060 77450
rect 16190 77440 16310 77450
rect 16440 77440 16560 77450
rect 16690 77440 16810 77450
rect 16940 77440 17060 77450
rect 17190 77440 17310 77450
rect 17440 77440 17560 77450
rect 17690 77440 17810 77450
rect 17940 77440 18060 77450
rect 18190 77440 18310 77450
rect 18440 77440 18560 77450
rect 18690 77440 18810 77450
rect 18940 77440 19060 77450
rect 19190 77440 19310 77450
rect 19440 77440 19560 77450
rect 19690 77440 19810 77450
rect 19940 77440 20060 77450
rect 20190 77440 20310 77450
rect 20440 77440 20560 77450
rect 20690 77440 20810 77450
rect 20940 77440 21060 77450
rect 21190 77440 21310 77450
rect 21440 77440 21560 77450
rect 21690 77440 21810 77450
rect 21940 77440 22060 77450
rect 22190 77440 22310 77450
rect 22440 77440 22560 77450
rect 22690 77440 22810 77450
rect 22940 77440 23060 77450
rect 23190 77440 23310 77450
rect 23440 77440 23560 77450
rect 23690 77440 23810 77450
rect 23940 77440 24060 77450
rect 24190 77440 24310 77450
rect 24440 77440 24560 77450
rect 24690 77440 24810 77450
rect 24940 77440 25060 77450
rect 25190 77440 25310 77450
rect 25440 77440 25560 77450
rect 25690 77440 25810 77450
rect 25940 77440 26060 77450
rect 26190 77440 26310 77450
rect 26440 77440 26560 77450
rect 26690 77440 26810 77450
rect 26940 77440 27060 77450
rect 27190 77440 27310 77450
rect 27440 77440 27560 77450
rect 27690 77440 27810 77450
rect 27940 77440 28060 77450
rect 28190 77440 28310 77450
rect 28440 77440 28560 77450
rect 28690 77440 28810 77450
rect 28940 77440 29000 77450
rect 7000 77310 7050 77440
rect 7200 77310 7300 77440
rect 7450 77310 7550 77440
rect 7700 77310 7800 77440
rect 7950 77310 8050 77440
rect 8200 77310 8300 77440
rect 8450 77310 8550 77440
rect 8700 77310 8800 77440
rect 8950 77310 9050 77440
rect 9200 77310 9300 77440
rect 9450 77310 9550 77440
rect 9700 77310 9800 77440
rect 9950 77310 10050 77440
rect 10200 77310 10300 77440
rect 10450 77310 10550 77440
rect 10700 77310 10800 77440
rect 10950 77310 11050 77440
rect 11200 77310 11300 77440
rect 11450 77310 11550 77440
rect 11700 77310 11800 77440
rect 11950 77310 12050 77440
rect 12200 77310 12300 77440
rect 12450 77310 12550 77440
rect 12700 77310 12800 77440
rect 12950 77310 13050 77440
rect 13200 77310 13300 77440
rect 13450 77310 13550 77440
rect 13700 77310 13800 77440
rect 13950 77310 14050 77440
rect 14200 77310 14300 77440
rect 14450 77310 14550 77440
rect 14700 77310 14800 77440
rect 14950 77310 15050 77440
rect 15200 77310 15300 77440
rect 15450 77310 15550 77440
rect 15700 77310 15800 77440
rect 15950 77310 16050 77440
rect 16200 77310 16300 77440
rect 16450 77310 16550 77440
rect 16700 77310 16800 77440
rect 16950 77310 17050 77440
rect 17200 77310 17300 77440
rect 17450 77310 17550 77440
rect 17700 77310 17800 77440
rect 17950 77310 18050 77440
rect 18200 77310 18300 77440
rect 18450 77310 18550 77440
rect 18700 77310 18800 77440
rect 18950 77310 19050 77440
rect 19200 77310 19300 77440
rect 19450 77310 19550 77440
rect 19700 77310 19800 77440
rect 19950 77310 20050 77440
rect 20200 77310 20300 77440
rect 20450 77310 20550 77440
rect 20700 77310 20800 77440
rect 20950 77310 21050 77440
rect 21200 77310 21300 77440
rect 21450 77310 21550 77440
rect 21700 77310 21800 77440
rect 21950 77310 22050 77440
rect 22200 77310 22300 77440
rect 22450 77310 22550 77440
rect 22700 77310 22800 77440
rect 22950 77310 23050 77440
rect 23200 77310 23300 77440
rect 23450 77310 23550 77440
rect 23700 77310 23800 77440
rect 23950 77310 24050 77440
rect 24200 77310 24300 77440
rect 24450 77310 24550 77440
rect 24700 77310 24800 77440
rect 24950 77310 25050 77440
rect 25200 77310 25300 77440
rect 25450 77310 25550 77440
rect 25700 77310 25800 77440
rect 25950 77310 26050 77440
rect 26200 77310 26300 77440
rect 26450 77310 26550 77440
rect 26700 77310 26800 77440
rect 26950 77310 27050 77440
rect 27200 77310 27300 77440
rect 27450 77310 27550 77440
rect 27700 77310 27800 77440
rect 27950 77310 28050 77440
rect 28200 77310 28300 77440
rect 28450 77310 28550 77440
rect 28700 77310 28800 77440
rect 28950 77310 29000 77440
rect 7000 77300 7060 77310
rect 7190 77300 7310 77310
rect 7440 77300 7560 77310
rect 7690 77300 7810 77310
rect 7940 77300 8060 77310
rect 8190 77300 8310 77310
rect 8440 77300 8560 77310
rect 8690 77300 8810 77310
rect 8940 77300 9060 77310
rect 9190 77300 9310 77310
rect 9440 77300 9560 77310
rect 9690 77300 9810 77310
rect 9940 77300 10060 77310
rect 10190 77300 10310 77310
rect 10440 77300 10560 77310
rect 10690 77300 10810 77310
rect 10940 77300 11060 77310
rect 11190 77300 11310 77310
rect 11440 77300 11560 77310
rect 11690 77300 11810 77310
rect 11940 77300 12060 77310
rect 12190 77300 12310 77310
rect 12440 77300 12560 77310
rect 12690 77300 12810 77310
rect 12940 77300 13060 77310
rect 13190 77300 13310 77310
rect 13440 77300 13560 77310
rect 13690 77300 13810 77310
rect 13940 77300 14060 77310
rect 14190 77300 14310 77310
rect 14440 77300 14560 77310
rect 14690 77300 14810 77310
rect 14940 77300 15060 77310
rect 15190 77300 15310 77310
rect 15440 77300 15560 77310
rect 15690 77300 15810 77310
rect 15940 77300 16060 77310
rect 16190 77300 16310 77310
rect 16440 77300 16560 77310
rect 16690 77300 16810 77310
rect 16940 77300 17060 77310
rect 17190 77300 17310 77310
rect 17440 77300 17560 77310
rect 17690 77300 17810 77310
rect 17940 77300 18060 77310
rect 18190 77300 18310 77310
rect 18440 77300 18560 77310
rect 18690 77300 18810 77310
rect 18940 77300 19060 77310
rect 19190 77300 19310 77310
rect 19440 77300 19560 77310
rect 19690 77300 19810 77310
rect 19940 77300 20060 77310
rect 20190 77300 20310 77310
rect 20440 77300 20560 77310
rect 20690 77300 20810 77310
rect 20940 77300 21060 77310
rect 21190 77300 21310 77310
rect 21440 77300 21560 77310
rect 21690 77300 21810 77310
rect 21940 77300 22060 77310
rect 22190 77300 22310 77310
rect 22440 77300 22560 77310
rect 22690 77300 22810 77310
rect 22940 77300 23060 77310
rect 23190 77300 23310 77310
rect 23440 77300 23560 77310
rect 23690 77300 23810 77310
rect 23940 77300 24060 77310
rect 24190 77300 24310 77310
rect 24440 77300 24560 77310
rect 24690 77300 24810 77310
rect 24940 77300 25060 77310
rect 25190 77300 25310 77310
rect 25440 77300 25560 77310
rect 25690 77300 25810 77310
rect 25940 77300 26060 77310
rect 26190 77300 26310 77310
rect 26440 77300 26560 77310
rect 26690 77300 26810 77310
rect 26940 77300 27060 77310
rect 27190 77300 27310 77310
rect 27440 77300 27560 77310
rect 27690 77300 27810 77310
rect 27940 77300 28060 77310
rect 28190 77300 28310 77310
rect 28440 77300 28560 77310
rect 28690 77300 28810 77310
rect 28940 77300 29000 77310
rect 7000 77200 29000 77300
rect 7000 77190 7060 77200
rect 7190 77190 7310 77200
rect 7440 77190 7560 77200
rect 7690 77190 7810 77200
rect 7940 77190 8060 77200
rect 8190 77190 8310 77200
rect 8440 77190 8560 77200
rect 8690 77190 8810 77200
rect 8940 77190 9060 77200
rect 9190 77190 9310 77200
rect 9440 77190 9560 77200
rect 9690 77190 9810 77200
rect 9940 77190 10060 77200
rect 10190 77190 10310 77200
rect 10440 77190 10560 77200
rect 10690 77190 10810 77200
rect 10940 77190 11060 77200
rect 11190 77190 11310 77200
rect 11440 77190 11560 77200
rect 11690 77190 11810 77200
rect 11940 77190 12060 77200
rect 12190 77190 12310 77200
rect 12440 77190 12560 77200
rect 12690 77190 12810 77200
rect 12940 77190 13060 77200
rect 13190 77190 13310 77200
rect 13440 77190 13560 77200
rect 13690 77190 13810 77200
rect 13940 77190 14060 77200
rect 14190 77190 14310 77200
rect 14440 77190 14560 77200
rect 14690 77190 14810 77200
rect 14940 77190 15060 77200
rect 15190 77190 15310 77200
rect 15440 77190 15560 77200
rect 15690 77190 15810 77200
rect 15940 77190 16060 77200
rect 16190 77190 16310 77200
rect 16440 77190 16560 77200
rect 16690 77190 16810 77200
rect 16940 77190 17060 77200
rect 17190 77190 17310 77200
rect 17440 77190 17560 77200
rect 17690 77190 17810 77200
rect 17940 77190 18060 77200
rect 18190 77190 18310 77200
rect 18440 77190 18560 77200
rect 18690 77190 18810 77200
rect 18940 77190 19060 77200
rect 19190 77190 19310 77200
rect 19440 77190 19560 77200
rect 19690 77190 19810 77200
rect 19940 77190 20060 77200
rect 20190 77190 20310 77200
rect 20440 77190 20560 77200
rect 20690 77190 20810 77200
rect 20940 77190 21060 77200
rect 21190 77190 21310 77200
rect 21440 77190 21560 77200
rect 21690 77190 21810 77200
rect 21940 77190 22060 77200
rect 22190 77190 22310 77200
rect 22440 77190 22560 77200
rect 22690 77190 22810 77200
rect 22940 77190 23060 77200
rect 23190 77190 23310 77200
rect 23440 77190 23560 77200
rect 23690 77190 23810 77200
rect 23940 77190 24060 77200
rect 24190 77190 24310 77200
rect 24440 77190 24560 77200
rect 24690 77190 24810 77200
rect 24940 77190 25060 77200
rect 25190 77190 25310 77200
rect 25440 77190 25560 77200
rect 25690 77190 25810 77200
rect 25940 77190 26060 77200
rect 26190 77190 26310 77200
rect 26440 77190 26560 77200
rect 26690 77190 26810 77200
rect 26940 77190 27060 77200
rect 27190 77190 27310 77200
rect 27440 77190 27560 77200
rect 27690 77190 27810 77200
rect 27940 77190 28060 77200
rect 28190 77190 28310 77200
rect 28440 77190 28560 77200
rect 28690 77190 28810 77200
rect 28940 77190 29000 77200
rect 7000 77060 7050 77190
rect 7200 77060 7300 77190
rect 7450 77060 7550 77190
rect 7700 77060 7800 77190
rect 7950 77060 8050 77190
rect 8200 77060 8300 77190
rect 8450 77060 8550 77190
rect 8700 77060 8800 77190
rect 8950 77060 9050 77190
rect 9200 77060 9300 77190
rect 9450 77060 9550 77190
rect 9700 77060 9800 77190
rect 9950 77060 10050 77190
rect 10200 77060 10300 77190
rect 10450 77060 10550 77190
rect 10700 77060 10800 77190
rect 10950 77060 11050 77190
rect 11200 77060 11300 77190
rect 11450 77060 11550 77190
rect 11700 77060 11800 77190
rect 11950 77060 12050 77190
rect 12200 77060 12300 77190
rect 12450 77060 12550 77190
rect 12700 77060 12800 77190
rect 12950 77060 13050 77190
rect 13200 77060 13300 77190
rect 13450 77060 13550 77190
rect 13700 77060 13800 77190
rect 13950 77060 14050 77190
rect 14200 77060 14300 77190
rect 14450 77060 14550 77190
rect 14700 77060 14800 77190
rect 14950 77060 15050 77190
rect 15200 77060 15300 77190
rect 15450 77060 15550 77190
rect 15700 77060 15800 77190
rect 15950 77060 16050 77190
rect 16200 77060 16300 77190
rect 16450 77060 16550 77190
rect 16700 77060 16800 77190
rect 16950 77060 17050 77190
rect 17200 77060 17300 77190
rect 17450 77060 17550 77190
rect 17700 77060 17800 77190
rect 17950 77060 18050 77190
rect 18200 77060 18300 77190
rect 18450 77060 18550 77190
rect 18700 77060 18800 77190
rect 18950 77060 19050 77190
rect 19200 77060 19300 77190
rect 19450 77060 19550 77190
rect 19700 77060 19800 77190
rect 19950 77060 20050 77190
rect 20200 77060 20300 77190
rect 20450 77060 20550 77190
rect 20700 77060 20800 77190
rect 20950 77060 21050 77190
rect 21200 77060 21300 77190
rect 21450 77060 21550 77190
rect 21700 77060 21800 77190
rect 21950 77060 22050 77190
rect 22200 77060 22300 77190
rect 22450 77060 22550 77190
rect 22700 77060 22800 77190
rect 22950 77060 23050 77190
rect 23200 77060 23300 77190
rect 23450 77060 23550 77190
rect 23700 77060 23800 77190
rect 23950 77060 24050 77190
rect 24200 77060 24300 77190
rect 24450 77060 24550 77190
rect 24700 77060 24800 77190
rect 24950 77060 25050 77190
rect 25200 77060 25300 77190
rect 25450 77060 25550 77190
rect 25700 77060 25800 77190
rect 25950 77060 26050 77190
rect 26200 77060 26300 77190
rect 26450 77060 26550 77190
rect 26700 77060 26800 77190
rect 26950 77060 27050 77190
rect 27200 77060 27300 77190
rect 27450 77060 27550 77190
rect 27700 77060 27800 77190
rect 27950 77060 28050 77190
rect 28200 77060 28300 77190
rect 28450 77060 28550 77190
rect 28700 77060 28800 77190
rect 28950 77060 29000 77190
rect 7000 77050 7060 77060
rect 7190 77050 7310 77060
rect 7440 77050 7560 77060
rect 7690 77050 7810 77060
rect 7940 77050 8060 77060
rect 8190 77050 8310 77060
rect 8440 77050 8560 77060
rect 8690 77050 8810 77060
rect 8940 77050 9060 77060
rect 9190 77050 9310 77060
rect 9440 77050 9560 77060
rect 9690 77050 9810 77060
rect 9940 77050 10060 77060
rect 10190 77050 10310 77060
rect 10440 77050 10560 77060
rect 10690 77050 10810 77060
rect 10940 77050 11060 77060
rect 11190 77050 11310 77060
rect 11440 77050 11560 77060
rect 11690 77050 11810 77060
rect 11940 77050 12060 77060
rect 12190 77050 12310 77060
rect 12440 77050 12560 77060
rect 12690 77050 12810 77060
rect 12940 77050 13060 77060
rect 13190 77050 13310 77060
rect 13440 77050 13560 77060
rect 13690 77050 13810 77060
rect 13940 77050 14060 77060
rect 14190 77050 14310 77060
rect 14440 77050 14560 77060
rect 14690 77050 14810 77060
rect 14940 77050 15060 77060
rect 15190 77050 15310 77060
rect 15440 77050 15560 77060
rect 15690 77050 15810 77060
rect 15940 77050 16060 77060
rect 16190 77050 16310 77060
rect 16440 77050 16560 77060
rect 16690 77050 16810 77060
rect 16940 77050 17060 77060
rect 17190 77050 17310 77060
rect 17440 77050 17560 77060
rect 17690 77050 17810 77060
rect 17940 77050 18060 77060
rect 18190 77050 18310 77060
rect 18440 77050 18560 77060
rect 18690 77050 18810 77060
rect 18940 77050 19060 77060
rect 19190 77050 19310 77060
rect 19440 77050 19560 77060
rect 19690 77050 19810 77060
rect 19940 77050 20060 77060
rect 20190 77050 20310 77060
rect 20440 77050 20560 77060
rect 20690 77050 20810 77060
rect 20940 77050 21060 77060
rect 21190 77050 21310 77060
rect 21440 77050 21560 77060
rect 21690 77050 21810 77060
rect 21940 77050 22060 77060
rect 22190 77050 22310 77060
rect 22440 77050 22560 77060
rect 22690 77050 22810 77060
rect 22940 77050 23060 77060
rect 23190 77050 23310 77060
rect 23440 77050 23560 77060
rect 23690 77050 23810 77060
rect 23940 77050 24060 77060
rect 24190 77050 24310 77060
rect 24440 77050 24560 77060
rect 24690 77050 24810 77060
rect 24940 77050 25060 77060
rect 25190 77050 25310 77060
rect 25440 77050 25560 77060
rect 25690 77050 25810 77060
rect 25940 77050 26060 77060
rect 26190 77050 26310 77060
rect 26440 77050 26560 77060
rect 26690 77050 26810 77060
rect 26940 77050 27060 77060
rect 27190 77050 27310 77060
rect 27440 77050 27560 77060
rect 27690 77050 27810 77060
rect 27940 77050 28060 77060
rect 28190 77050 28310 77060
rect 28440 77050 28560 77060
rect 28690 77050 28810 77060
rect 28940 77050 29000 77060
rect 7000 77000 29000 77050
rect 59000 80950 71000 81000
rect 59000 80940 59060 80950
rect 59190 80940 59310 80950
rect 59440 80940 59560 80950
rect 59690 80940 59810 80950
rect 59940 80940 60060 80950
rect 60190 80940 60310 80950
rect 60440 80940 60560 80950
rect 60690 80940 60810 80950
rect 60940 80940 61060 80950
rect 61190 80940 61310 80950
rect 61440 80940 61560 80950
rect 61690 80940 61810 80950
rect 61940 80940 62060 80950
rect 62190 80940 62310 80950
rect 62440 80940 62560 80950
rect 62690 80940 62810 80950
rect 62940 80940 63060 80950
rect 63190 80940 63310 80950
rect 63440 80940 63560 80950
rect 63690 80940 63810 80950
rect 63940 80940 64060 80950
rect 64190 80940 64310 80950
rect 64440 80940 64560 80950
rect 64690 80940 64810 80950
rect 64940 80940 65060 80950
rect 65190 80940 65310 80950
rect 65440 80940 65560 80950
rect 65690 80940 65810 80950
rect 65940 80940 66060 80950
rect 66190 80940 66310 80950
rect 66440 80940 66560 80950
rect 66690 80940 66810 80950
rect 66940 80940 67060 80950
rect 67190 80940 67310 80950
rect 67440 80940 67560 80950
rect 67690 80940 67810 80950
rect 67940 80940 68060 80950
rect 68190 80940 68310 80950
rect 68440 80940 68560 80950
rect 68690 80940 68810 80950
rect 68940 80940 69060 80950
rect 69190 80940 69310 80950
rect 69440 80940 69560 80950
rect 69690 80940 69810 80950
rect 69940 80940 70060 80950
rect 70190 80940 70310 80950
rect 70440 80940 70560 80950
rect 70690 80940 70810 80950
rect 70940 80940 71000 80950
rect 59000 80810 59050 80940
rect 59200 80810 59300 80940
rect 59450 80810 59550 80940
rect 59700 80810 59800 80940
rect 59950 80810 60050 80940
rect 60200 80810 60300 80940
rect 60450 80810 60550 80940
rect 60700 80810 60800 80940
rect 60950 80810 61050 80940
rect 61200 80810 61300 80940
rect 61450 80810 61550 80940
rect 61700 80810 61800 80940
rect 61950 80810 62050 80940
rect 62200 80810 62300 80940
rect 62450 80810 62550 80940
rect 62700 80810 62800 80940
rect 62950 80810 63050 80940
rect 63200 80810 63300 80940
rect 63450 80810 63550 80940
rect 63700 80810 63800 80940
rect 63950 80810 64050 80940
rect 64200 80810 64300 80940
rect 64450 80810 64550 80940
rect 64700 80810 64800 80940
rect 64950 80810 65050 80940
rect 65200 80810 65300 80940
rect 65450 80810 65550 80940
rect 65700 80810 65800 80940
rect 65950 80810 66050 80940
rect 66200 80810 66300 80940
rect 66450 80810 66550 80940
rect 66700 80810 66800 80940
rect 66950 80810 67050 80940
rect 67200 80810 67300 80940
rect 67450 80810 67550 80940
rect 67700 80810 67800 80940
rect 67950 80810 68050 80940
rect 68200 80810 68300 80940
rect 68450 80810 68550 80940
rect 68700 80810 68800 80940
rect 68950 80810 69050 80940
rect 69200 80810 69300 80940
rect 69450 80810 69550 80940
rect 69700 80810 69800 80940
rect 69950 80810 70050 80940
rect 70200 80810 70300 80940
rect 70450 80810 70550 80940
rect 70700 80810 70800 80940
rect 70950 80810 71000 80940
rect 59000 80800 59060 80810
rect 59190 80800 59310 80810
rect 59440 80800 59560 80810
rect 59690 80800 59810 80810
rect 59940 80800 60060 80810
rect 60190 80800 60310 80810
rect 60440 80800 60560 80810
rect 60690 80800 60810 80810
rect 60940 80800 61060 80810
rect 61190 80800 61310 80810
rect 61440 80800 61560 80810
rect 61690 80800 61810 80810
rect 61940 80800 62060 80810
rect 62190 80800 62310 80810
rect 62440 80800 62560 80810
rect 62690 80800 62810 80810
rect 62940 80800 63060 80810
rect 63190 80800 63310 80810
rect 63440 80800 63560 80810
rect 63690 80800 63810 80810
rect 63940 80800 64060 80810
rect 64190 80800 64310 80810
rect 64440 80800 64560 80810
rect 64690 80800 64810 80810
rect 64940 80800 65060 80810
rect 65190 80800 65310 80810
rect 65440 80800 65560 80810
rect 65690 80800 65810 80810
rect 65940 80800 66060 80810
rect 66190 80800 66310 80810
rect 66440 80800 66560 80810
rect 66690 80800 66810 80810
rect 66940 80800 67060 80810
rect 67190 80800 67310 80810
rect 67440 80800 67560 80810
rect 67690 80800 67810 80810
rect 67940 80800 68060 80810
rect 68190 80800 68310 80810
rect 68440 80800 68560 80810
rect 68690 80800 68810 80810
rect 68940 80800 69060 80810
rect 69190 80800 69310 80810
rect 69440 80800 69560 80810
rect 69690 80800 69810 80810
rect 69940 80800 70060 80810
rect 70190 80800 70310 80810
rect 70440 80800 70560 80810
rect 70690 80800 70810 80810
rect 70940 80800 71000 80810
rect 59000 80700 71000 80800
rect 59000 80690 59060 80700
rect 59190 80690 59310 80700
rect 59440 80690 59560 80700
rect 59690 80690 59810 80700
rect 59940 80690 60060 80700
rect 60190 80690 60310 80700
rect 60440 80690 60560 80700
rect 60690 80690 60810 80700
rect 60940 80690 61060 80700
rect 61190 80690 61310 80700
rect 61440 80690 61560 80700
rect 61690 80690 61810 80700
rect 61940 80690 62060 80700
rect 62190 80690 62310 80700
rect 62440 80690 62560 80700
rect 62690 80690 62810 80700
rect 62940 80690 63060 80700
rect 63190 80690 63310 80700
rect 63440 80690 63560 80700
rect 63690 80690 63810 80700
rect 63940 80690 64060 80700
rect 64190 80690 64310 80700
rect 64440 80690 64560 80700
rect 64690 80690 64810 80700
rect 64940 80690 65060 80700
rect 65190 80690 65310 80700
rect 65440 80690 65560 80700
rect 65690 80690 65810 80700
rect 65940 80690 66060 80700
rect 66190 80690 66310 80700
rect 66440 80690 66560 80700
rect 66690 80690 66810 80700
rect 66940 80690 67060 80700
rect 67190 80690 67310 80700
rect 67440 80690 67560 80700
rect 67690 80690 67810 80700
rect 67940 80690 68060 80700
rect 68190 80690 68310 80700
rect 68440 80690 68560 80700
rect 68690 80690 68810 80700
rect 68940 80690 69060 80700
rect 69190 80690 69310 80700
rect 69440 80690 69560 80700
rect 69690 80690 69810 80700
rect 69940 80690 70060 80700
rect 70190 80690 70310 80700
rect 70440 80690 70560 80700
rect 70690 80690 70810 80700
rect 70940 80690 71000 80700
rect 59000 80560 59050 80690
rect 59200 80560 59300 80690
rect 59450 80560 59550 80690
rect 59700 80560 59800 80690
rect 59950 80560 60050 80690
rect 60200 80560 60300 80690
rect 60450 80560 60550 80690
rect 60700 80560 60800 80690
rect 60950 80560 61050 80690
rect 61200 80560 61300 80690
rect 61450 80560 61550 80690
rect 61700 80560 61800 80690
rect 61950 80560 62050 80690
rect 62200 80560 62300 80690
rect 62450 80560 62550 80690
rect 62700 80560 62800 80690
rect 62950 80560 63050 80690
rect 63200 80560 63300 80690
rect 63450 80560 63550 80690
rect 63700 80560 63800 80690
rect 63950 80560 64050 80690
rect 64200 80560 64300 80690
rect 64450 80560 64550 80690
rect 64700 80560 64800 80690
rect 64950 80560 65050 80690
rect 65200 80560 65300 80690
rect 65450 80560 65550 80690
rect 65700 80560 65800 80690
rect 65950 80560 66050 80690
rect 66200 80560 66300 80690
rect 66450 80560 66550 80690
rect 66700 80560 66800 80690
rect 66950 80560 67050 80690
rect 67200 80560 67300 80690
rect 67450 80560 67550 80690
rect 67700 80560 67800 80690
rect 67950 80560 68050 80690
rect 68200 80560 68300 80690
rect 68450 80560 68550 80690
rect 68700 80560 68800 80690
rect 68950 80560 69050 80690
rect 69200 80560 69300 80690
rect 69450 80560 69550 80690
rect 69700 80560 69800 80690
rect 69950 80560 70050 80690
rect 70200 80560 70300 80690
rect 70450 80560 70550 80690
rect 70700 80560 70800 80690
rect 70950 80560 71000 80690
rect 59000 80550 59060 80560
rect 59190 80550 59310 80560
rect 59440 80550 59560 80560
rect 59690 80550 59810 80560
rect 59940 80550 60060 80560
rect 60190 80550 60310 80560
rect 60440 80550 60560 80560
rect 60690 80550 60810 80560
rect 60940 80550 61060 80560
rect 61190 80550 61310 80560
rect 61440 80550 61560 80560
rect 61690 80550 61810 80560
rect 61940 80550 62060 80560
rect 62190 80550 62310 80560
rect 62440 80550 62560 80560
rect 62690 80550 62810 80560
rect 62940 80550 63060 80560
rect 63190 80550 63310 80560
rect 63440 80550 63560 80560
rect 63690 80550 63810 80560
rect 63940 80550 64060 80560
rect 64190 80550 64310 80560
rect 64440 80550 64560 80560
rect 64690 80550 64810 80560
rect 64940 80550 65060 80560
rect 65190 80550 65310 80560
rect 65440 80550 65560 80560
rect 65690 80550 65810 80560
rect 65940 80550 66060 80560
rect 66190 80550 66310 80560
rect 66440 80550 66560 80560
rect 66690 80550 66810 80560
rect 66940 80550 67060 80560
rect 67190 80550 67310 80560
rect 67440 80550 67560 80560
rect 67690 80550 67810 80560
rect 67940 80550 68060 80560
rect 68190 80550 68310 80560
rect 68440 80550 68560 80560
rect 68690 80550 68810 80560
rect 68940 80550 69060 80560
rect 69190 80550 69310 80560
rect 69440 80550 69560 80560
rect 69690 80550 69810 80560
rect 69940 80550 70060 80560
rect 70190 80550 70310 80560
rect 70440 80550 70560 80560
rect 70690 80550 70810 80560
rect 70940 80550 71000 80560
rect 59000 80450 71000 80550
rect 59000 80440 59060 80450
rect 59190 80440 59310 80450
rect 59440 80440 59560 80450
rect 59690 80440 59810 80450
rect 59940 80440 60060 80450
rect 60190 80440 60310 80450
rect 60440 80440 60560 80450
rect 60690 80440 60810 80450
rect 60940 80440 61060 80450
rect 61190 80440 61310 80450
rect 61440 80440 61560 80450
rect 61690 80440 61810 80450
rect 61940 80440 62060 80450
rect 62190 80440 62310 80450
rect 62440 80440 62560 80450
rect 62690 80440 62810 80450
rect 62940 80440 63060 80450
rect 63190 80440 63310 80450
rect 63440 80440 63560 80450
rect 63690 80440 63810 80450
rect 63940 80440 64060 80450
rect 64190 80440 64310 80450
rect 64440 80440 64560 80450
rect 64690 80440 64810 80450
rect 64940 80440 65060 80450
rect 65190 80440 65310 80450
rect 65440 80440 65560 80450
rect 65690 80440 65810 80450
rect 65940 80440 66060 80450
rect 66190 80440 66310 80450
rect 66440 80440 66560 80450
rect 66690 80440 66810 80450
rect 66940 80440 67060 80450
rect 67190 80440 67310 80450
rect 67440 80440 67560 80450
rect 67690 80440 67810 80450
rect 67940 80440 68060 80450
rect 68190 80440 68310 80450
rect 68440 80440 68560 80450
rect 68690 80440 68810 80450
rect 68940 80440 69060 80450
rect 69190 80440 69310 80450
rect 69440 80440 69560 80450
rect 69690 80440 69810 80450
rect 69940 80440 70060 80450
rect 70190 80440 70310 80450
rect 70440 80440 70560 80450
rect 70690 80440 70810 80450
rect 70940 80440 71000 80450
rect 59000 80310 59050 80440
rect 59200 80310 59300 80440
rect 59450 80310 59550 80440
rect 59700 80310 59800 80440
rect 59950 80310 60050 80440
rect 60200 80310 60300 80440
rect 60450 80310 60550 80440
rect 60700 80310 60800 80440
rect 60950 80310 61050 80440
rect 61200 80310 61300 80440
rect 61450 80310 61550 80440
rect 61700 80310 61800 80440
rect 61950 80310 62050 80440
rect 62200 80310 62300 80440
rect 62450 80310 62550 80440
rect 62700 80310 62800 80440
rect 62950 80310 63050 80440
rect 63200 80310 63300 80440
rect 63450 80310 63550 80440
rect 63700 80310 63800 80440
rect 63950 80310 64050 80440
rect 64200 80310 64300 80440
rect 64450 80310 64550 80440
rect 64700 80310 64800 80440
rect 64950 80310 65050 80440
rect 65200 80310 65300 80440
rect 65450 80310 65550 80440
rect 65700 80310 65800 80440
rect 65950 80310 66050 80440
rect 66200 80310 66300 80440
rect 66450 80310 66550 80440
rect 66700 80310 66800 80440
rect 66950 80310 67050 80440
rect 67200 80310 67300 80440
rect 67450 80310 67550 80440
rect 67700 80310 67800 80440
rect 67950 80310 68050 80440
rect 68200 80310 68300 80440
rect 68450 80310 68550 80440
rect 68700 80310 68800 80440
rect 68950 80310 69050 80440
rect 69200 80310 69300 80440
rect 69450 80310 69550 80440
rect 69700 80310 69800 80440
rect 69950 80310 70050 80440
rect 70200 80310 70300 80440
rect 70450 80310 70550 80440
rect 70700 80310 70800 80440
rect 70950 80310 71000 80440
rect 59000 80300 59060 80310
rect 59190 80300 59310 80310
rect 59440 80300 59560 80310
rect 59690 80300 59810 80310
rect 59940 80300 60060 80310
rect 60190 80300 60310 80310
rect 60440 80300 60560 80310
rect 60690 80300 60810 80310
rect 60940 80300 61060 80310
rect 61190 80300 61310 80310
rect 61440 80300 61560 80310
rect 61690 80300 61810 80310
rect 61940 80300 62060 80310
rect 62190 80300 62310 80310
rect 62440 80300 62560 80310
rect 62690 80300 62810 80310
rect 62940 80300 63060 80310
rect 63190 80300 63310 80310
rect 63440 80300 63560 80310
rect 63690 80300 63810 80310
rect 63940 80300 64060 80310
rect 64190 80300 64310 80310
rect 64440 80300 64560 80310
rect 64690 80300 64810 80310
rect 64940 80300 65060 80310
rect 65190 80300 65310 80310
rect 65440 80300 65560 80310
rect 65690 80300 65810 80310
rect 65940 80300 66060 80310
rect 66190 80300 66310 80310
rect 66440 80300 66560 80310
rect 66690 80300 66810 80310
rect 66940 80300 67060 80310
rect 67190 80300 67310 80310
rect 67440 80300 67560 80310
rect 67690 80300 67810 80310
rect 67940 80300 68060 80310
rect 68190 80300 68310 80310
rect 68440 80300 68560 80310
rect 68690 80300 68810 80310
rect 68940 80300 69060 80310
rect 69190 80300 69310 80310
rect 69440 80300 69560 80310
rect 69690 80300 69810 80310
rect 69940 80300 70060 80310
rect 70190 80300 70310 80310
rect 70440 80300 70560 80310
rect 70690 80300 70810 80310
rect 70940 80300 71000 80310
rect 59000 80200 71000 80300
rect 59000 80190 59060 80200
rect 59190 80190 59310 80200
rect 59440 80190 59560 80200
rect 59690 80190 59810 80200
rect 59940 80190 60060 80200
rect 60190 80190 60310 80200
rect 60440 80190 60560 80200
rect 60690 80190 60810 80200
rect 60940 80190 61060 80200
rect 61190 80190 61310 80200
rect 61440 80190 61560 80200
rect 61690 80190 61810 80200
rect 61940 80190 62060 80200
rect 62190 80190 62310 80200
rect 62440 80190 62560 80200
rect 62690 80190 62810 80200
rect 62940 80190 63060 80200
rect 63190 80190 63310 80200
rect 63440 80190 63560 80200
rect 63690 80190 63810 80200
rect 63940 80190 64060 80200
rect 64190 80190 64310 80200
rect 64440 80190 64560 80200
rect 64690 80190 64810 80200
rect 64940 80190 65060 80200
rect 65190 80190 65310 80200
rect 65440 80190 65560 80200
rect 65690 80190 65810 80200
rect 65940 80190 66060 80200
rect 66190 80190 66310 80200
rect 66440 80190 66560 80200
rect 66690 80190 66810 80200
rect 66940 80190 67060 80200
rect 67190 80190 67310 80200
rect 67440 80190 67560 80200
rect 67690 80190 67810 80200
rect 67940 80190 68060 80200
rect 68190 80190 68310 80200
rect 68440 80190 68560 80200
rect 68690 80190 68810 80200
rect 68940 80190 69060 80200
rect 69190 80190 69310 80200
rect 69440 80190 69560 80200
rect 69690 80190 69810 80200
rect 69940 80190 70060 80200
rect 70190 80190 70310 80200
rect 70440 80190 70560 80200
rect 70690 80190 70810 80200
rect 70940 80190 71000 80200
rect 59000 80060 59050 80190
rect 59200 80060 59300 80190
rect 59450 80060 59550 80190
rect 59700 80060 59800 80190
rect 59950 80060 60050 80190
rect 60200 80060 60300 80190
rect 60450 80060 60550 80190
rect 60700 80060 60800 80190
rect 60950 80060 61050 80190
rect 61200 80060 61300 80190
rect 61450 80060 61550 80190
rect 61700 80060 61800 80190
rect 61950 80060 62050 80190
rect 62200 80060 62300 80190
rect 62450 80060 62550 80190
rect 62700 80060 62800 80190
rect 62950 80060 63050 80190
rect 63200 80060 63300 80190
rect 63450 80060 63550 80190
rect 63700 80060 63800 80190
rect 63950 80060 64050 80190
rect 64200 80060 64300 80190
rect 64450 80060 64550 80190
rect 64700 80060 64800 80190
rect 64950 80060 65050 80190
rect 65200 80060 65300 80190
rect 65450 80060 65550 80190
rect 65700 80060 65800 80190
rect 65950 80060 66050 80190
rect 66200 80060 66300 80190
rect 66450 80060 66550 80190
rect 66700 80060 66800 80190
rect 66950 80060 67050 80190
rect 67200 80060 67300 80190
rect 67450 80060 67550 80190
rect 67700 80060 67800 80190
rect 67950 80060 68050 80190
rect 68200 80060 68300 80190
rect 68450 80060 68550 80190
rect 68700 80060 68800 80190
rect 68950 80060 69050 80190
rect 69200 80060 69300 80190
rect 69450 80060 69550 80190
rect 69700 80060 69800 80190
rect 69950 80060 70050 80190
rect 70200 80060 70300 80190
rect 70450 80060 70550 80190
rect 70700 80060 70800 80190
rect 70950 80060 71000 80190
rect 59000 80050 59060 80060
rect 59190 80050 59310 80060
rect 59440 80050 59560 80060
rect 59690 80050 59810 80060
rect 59940 80050 60060 80060
rect 60190 80050 60310 80060
rect 60440 80050 60560 80060
rect 60690 80050 60810 80060
rect 60940 80050 61060 80060
rect 61190 80050 61310 80060
rect 61440 80050 61560 80060
rect 61690 80050 61810 80060
rect 61940 80050 62060 80060
rect 62190 80050 62310 80060
rect 62440 80050 62560 80060
rect 62690 80050 62810 80060
rect 62940 80050 63060 80060
rect 63190 80050 63310 80060
rect 63440 80050 63560 80060
rect 63690 80050 63810 80060
rect 63940 80050 64060 80060
rect 64190 80050 64310 80060
rect 64440 80050 64560 80060
rect 64690 80050 64810 80060
rect 64940 80050 65060 80060
rect 65190 80050 65310 80060
rect 65440 80050 65560 80060
rect 65690 80050 65810 80060
rect 65940 80050 66060 80060
rect 66190 80050 66310 80060
rect 66440 80050 66560 80060
rect 66690 80050 66810 80060
rect 66940 80050 67060 80060
rect 67190 80050 67310 80060
rect 67440 80050 67560 80060
rect 67690 80050 67810 80060
rect 67940 80050 68060 80060
rect 68190 80050 68310 80060
rect 68440 80050 68560 80060
rect 68690 80050 68810 80060
rect 68940 80050 69060 80060
rect 69190 80050 69310 80060
rect 69440 80050 69560 80060
rect 69690 80050 69810 80060
rect 69940 80050 70060 80060
rect 70190 80050 70310 80060
rect 70440 80050 70560 80060
rect 70690 80050 70810 80060
rect 70940 80050 71000 80060
rect 59000 79950 71000 80050
rect 59000 79940 59060 79950
rect 59190 79940 59310 79950
rect 59440 79940 59560 79950
rect 59690 79940 59810 79950
rect 59940 79940 60060 79950
rect 60190 79940 60310 79950
rect 60440 79940 60560 79950
rect 60690 79940 60810 79950
rect 60940 79940 61060 79950
rect 61190 79940 61310 79950
rect 61440 79940 61560 79950
rect 61690 79940 61810 79950
rect 61940 79940 62060 79950
rect 62190 79940 62310 79950
rect 62440 79940 62560 79950
rect 62690 79940 62810 79950
rect 62940 79940 63060 79950
rect 63190 79940 63310 79950
rect 63440 79940 63560 79950
rect 63690 79940 63810 79950
rect 63940 79940 64060 79950
rect 64190 79940 64310 79950
rect 64440 79940 64560 79950
rect 64690 79940 64810 79950
rect 64940 79940 65060 79950
rect 65190 79940 65310 79950
rect 65440 79940 65560 79950
rect 65690 79940 65810 79950
rect 65940 79940 66060 79950
rect 66190 79940 66310 79950
rect 66440 79940 66560 79950
rect 66690 79940 66810 79950
rect 66940 79940 67060 79950
rect 67190 79940 67310 79950
rect 67440 79940 67560 79950
rect 67690 79940 67810 79950
rect 67940 79940 68060 79950
rect 68190 79940 68310 79950
rect 68440 79940 68560 79950
rect 68690 79940 68810 79950
rect 68940 79940 69060 79950
rect 69190 79940 69310 79950
rect 69440 79940 69560 79950
rect 69690 79940 69810 79950
rect 69940 79940 70060 79950
rect 70190 79940 70310 79950
rect 70440 79940 70560 79950
rect 70690 79940 70810 79950
rect 70940 79940 71000 79950
rect 59000 79810 59050 79940
rect 59200 79810 59300 79940
rect 59450 79810 59550 79940
rect 59700 79810 59800 79940
rect 59950 79810 60050 79940
rect 60200 79810 60300 79940
rect 60450 79810 60550 79940
rect 60700 79810 60800 79940
rect 60950 79810 61050 79940
rect 61200 79810 61300 79940
rect 61450 79810 61550 79940
rect 61700 79810 61800 79940
rect 61950 79810 62050 79940
rect 62200 79810 62300 79940
rect 62450 79810 62550 79940
rect 62700 79810 62800 79940
rect 62950 79810 63050 79940
rect 63200 79810 63300 79940
rect 63450 79810 63550 79940
rect 63700 79810 63800 79940
rect 63950 79810 64050 79940
rect 64200 79810 64300 79940
rect 64450 79810 64550 79940
rect 64700 79810 64800 79940
rect 64950 79810 65050 79940
rect 65200 79810 65300 79940
rect 65450 79810 65550 79940
rect 65700 79810 65800 79940
rect 65950 79810 66050 79940
rect 66200 79810 66300 79940
rect 66450 79810 66550 79940
rect 66700 79810 66800 79940
rect 66950 79810 67050 79940
rect 67200 79810 67300 79940
rect 67450 79810 67550 79940
rect 67700 79810 67800 79940
rect 67950 79810 68050 79940
rect 68200 79810 68300 79940
rect 68450 79810 68550 79940
rect 68700 79810 68800 79940
rect 68950 79810 69050 79940
rect 69200 79810 69300 79940
rect 69450 79810 69550 79940
rect 69700 79810 69800 79940
rect 69950 79810 70050 79940
rect 70200 79810 70300 79940
rect 70450 79810 70550 79940
rect 70700 79810 70800 79940
rect 70950 79810 71000 79940
rect 59000 79800 59060 79810
rect 59190 79800 59310 79810
rect 59440 79800 59560 79810
rect 59690 79800 59810 79810
rect 59940 79800 60060 79810
rect 60190 79800 60310 79810
rect 60440 79800 60560 79810
rect 60690 79800 60810 79810
rect 60940 79800 61060 79810
rect 61190 79800 61310 79810
rect 61440 79800 61560 79810
rect 61690 79800 61810 79810
rect 61940 79800 62060 79810
rect 62190 79800 62310 79810
rect 62440 79800 62560 79810
rect 62690 79800 62810 79810
rect 62940 79800 63060 79810
rect 63190 79800 63310 79810
rect 63440 79800 63560 79810
rect 63690 79800 63810 79810
rect 63940 79800 64060 79810
rect 64190 79800 64310 79810
rect 64440 79800 64560 79810
rect 64690 79800 64810 79810
rect 64940 79800 65060 79810
rect 65190 79800 65310 79810
rect 65440 79800 65560 79810
rect 65690 79800 65810 79810
rect 65940 79800 66060 79810
rect 66190 79800 66310 79810
rect 66440 79800 66560 79810
rect 66690 79800 66810 79810
rect 66940 79800 67060 79810
rect 67190 79800 67310 79810
rect 67440 79800 67560 79810
rect 67690 79800 67810 79810
rect 67940 79800 68060 79810
rect 68190 79800 68310 79810
rect 68440 79800 68560 79810
rect 68690 79800 68810 79810
rect 68940 79800 69060 79810
rect 69190 79800 69310 79810
rect 69440 79800 69560 79810
rect 69690 79800 69810 79810
rect 69940 79800 70060 79810
rect 70190 79800 70310 79810
rect 70440 79800 70560 79810
rect 70690 79800 70810 79810
rect 70940 79800 71000 79810
rect 59000 79700 71000 79800
rect 59000 79690 59060 79700
rect 59190 79690 59310 79700
rect 59440 79690 59560 79700
rect 59690 79690 59810 79700
rect 59940 79690 60060 79700
rect 60190 79690 60310 79700
rect 60440 79690 60560 79700
rect 60690 79690 60810 79700
rect 60940 79690 61060 79700
rect 61190 79690 61310 79700
rect 61440 79690 61560 79700
rect 61690 79690 61810 79700
rect 61940 79690 62060 79700
rect 62190 79690 62310 79700
rect 62440 79690 62560 79700
rect 62690 79690 62810 79700
rect 62940 79690 63060 79700
rect 63190 79690 63310 79700
rect 63440 79690 63560 79700
rect 63690 79690 63810 79700
rect 63940 79690 64060 79700
rect 64190 79690 64310 79700
rect 64440 79690 64560 79700
rect 64690 79690 64810 79700
rect 64940 79690 65060 79700
rect 65190 79690 65310 79700
rect 65440 79690 65560 79700
rect 65690 79690 65810 79700
rect 65940 79690 66060 79700
rect 66190 79690 66310 79700
rect 66440 79690 66560 79700
rect 66690 79690 66810 79700
rect 66940 79690 67060 79700
rect 67190 79690 67310 79700
rect 67440 79690 67560 79700
rect 67690 79690 67810 79700
rect 67940 79690 68060 79700
rect 68190 79690 68310 79700
rect 68440 79690 68560 79700
rect 68690 79690 68810 79700
rect 68940 79690 69060 79700
rect 69190 79690 69310 79700
rect 69440 79690 69560 79700
rect 69690 79690 69810 79700
rect 69940 79690 70060 79700
rect 70190 79690 70310 79700
rect 70440 79690 70560 79700
rect 70690 79690 70810 79700
rect 70940 79690 71000 79700
rect 59000 79560 59050 79690
rect 59200 79560 59300 79690
rect 59450 79560 59550 79690
rect 59700 79560 59800 79690
rect 59950 79560 60050 79690
rect 60200 79560 60300 79690
rect 60450 79560 60550 79690
rect 60700 79560 60800 79690
rect 60950 79560 61050 79690
rect 61200 79560 61300 79690
rect 61450 79560 61550 79690
rect 61700 79560 61800 79690
rect 61950 79560 62050 79690
rect 62200 79560 62300 79690
rect 62450 79560 62550 79690
rect 62700 79560 62800 79690
rect 62950 79560 63050 79690
rect 63200 79560 63300 79690
rect 63450 79560 63550 79690
rect 63700 79560 63800 79690
rect 63950 79560 64050 79690
rect 64200 79560 64300 79690
rect 64450 79560 64550 79690
rect 64700 79560 64800 79690
rect 64950 79560 65050 79690
rect 65200 79560 65300 79690
rect 65450 79560 65550 79690
rect 65700 79560 65800 79690
rect 65950 79560 66050 79690
rect 66200 79560 66300 79690
rect 66450 79560 66550 79690
rect 66700 79560 66800 79690
rect 66950 79560 67050 79690
rect 67200 79560 67300 79690
rect 67450 79560 67550 79690
rect 67700 79560 67800 79690
rect 67950 79560 68050 79690
rect 68200 79560 68300 79690
rect 68450 79560 68550 79690
rect 68700 79560 68800 79690
rect 68950 79560 69050 79690
rect 69200 79560 69300 79690
rect 69450 79560 69550 79690
rect 69700 79560 69800 79690
rect 69950 79560 70050 79690
rect 70200 79560 70300 79690
rect 70450 79560 70550 79690
rect 70700 79560 70800 79690
rect 70950 79560 71000 79690
rect 59000 79550 59060 79560
rect 59190 79550 59310 79560
rect 59440 79550 59560 79560
rect 59690 79550 59810 79560
rect 59940 79550 60060 79560
rect 60190 79550 60310 79560
rect 60440 79550 60560 79560
rect 60690 79550 60810 79560
rect 60940 79550 61060 79560
rect 61190 79550 61310 79560
rect 61440 79550 61560 79560
rect 61690 79550 61810 79560
rect 61940 79550 62060 79560
rect 62190 79550 62310 79560
rect 62440 79550 62560 79560
rect 62690 79550 62810 79560
rect 62940 79550 63060 79560
rect 63190 79550 63310 79560
rect 63440 79550 63560 79560
rect 63690 79550 63810 79560
rect 63940 79550 64060 79560
rect 64190 79550 64310 79560
rect 64440 79550 64560 79560
rect 64690 79550 64810 79560
rect 64940 79550 65060 79560
rect 65190 79550 65310 79560
rect 65440 79550 65560 79560
rect 65690 79550 65810 79560
rect 65940 79550 66060 79560
rect 66190 79550 66310 79560
rect 66440 79550 66560 79560
rect 66690 79550 66810 79560
rect 66940 79550 67060 79560
rect 67190 79550 67310 79560
rect 67440 79550 67560 79560
rect 67690 79550 67810 79560
rect 67940 79550 68060 79560
rect 68190 79550 68310 79560
rect 68440 79550 68560 79560
rect 68690 79550 68810 79560
rect 68940 79550 69060 79560
rect 69190 79550 69310 79560
rect 69440 79550 69560 79560
rect 69690 79550 69810 79560
rect 69940 79550 70060 79560
rect 70190 79550 70310 79560
rect 70440 79550 70560 79560
rect 70690 79550 70810 79560
rect 70940 79550 71000 79560
rect 59000 79450 71000 79550
rect 59000 79440 59060 79450
rect 59190 79440 59310 79450
rect 59440 79440 59560 79450
rect 59690 79440 59810 79450
rect 59940 79440 60060 79450
rect 60190 79440 60310 79450
rect 60440 79440 60560 79450
rect 60690 79440 60810 79450
rect 60940 79440 61060 79450
rect 61190 79440 61310 79450
rect 61440 79440 61560 79450
rect 61690 79440 61810 79450
rect 61940 79440 62060 79450
rect 62190 79440 62310 79450
rect 62440 79440 62560 79450
rect 62690 79440 62810 79450
rect 62940 79440 63060 79450
rect 63190 79440 63310 79450
rect 63440 79440 63560 79450
rect 63690 79440 63810 79450
rect 63940 79440 64060 79450
rect 64190 79440 64310 79450
rect 64440 79440 64560 79450
rect 64690 79440 64810 79450
rect 64940 79440 65060 79450
rect 65190 79440 65310 79450
rect 65440 79440 65560 79450
rect 65690 79440 65810 79450
rect 65940 79440 66060 79450
rect 66190 79440 66310 79450
rect 66440 79440 66560 79450
rect 66690 79440 66810 79450
rect 66940 79440 67060 79450
rect 67190 79440 67310 79450
rect 67440 79440 67560 79450
rect 67690 79440 67810 79450
rect 67940 79440 68060 79450
rect 68190 79440 68310 79450
rect 68440 79440 68560 79450
rect 68690 79440 68810 79450
rect 68940 79440 69060 79450
rect 69190 79440 69310 79450
rect 69440 79440 69560 79450
rect 69690 79440 69810 79450
rect 69940 79440 70060 79450
rect 70190 79440 70310 79450
rect 70440 79440 70560 79450
rect 70690 79440 70810 79450
rect 70940 79440 71000 79450
rect 59000 79310 59050 79440
rect 59200 79310 59300 79440
rect 59450 79310 59550 79440
rect 59700 79310 59800 79440
rect 59950 79310 60050 79440
rect 60200 79310 60300 79440
rect 60450 79310 60550 79440
rect 60700 79310 60800 79440
rect 60950 79310 61050 79440
rect 61200 79310 61300 79440
rect 61450 79310 61550 79440
rect 61700 79310 61800 79440
rect 61950 79310 62050 79440
rect 62200 79310 62300 79440
rect 62450 79310 62550 79440
rect 62700 79310 62800 79440
rect 62950 79310 63050 79440
rect 63200 79310 63300 79440
rect 63450 79310 63550 79440
rect 63700 79310 63800 79440
rect 63950 79310 64050 79440
rect 64200 79310 64300 79440
rect 64450 79310 64550 79440
rect 64700 79310 64800 79440
rect 64950 79310 65050 79440
rect 65200 79310 65300 79440
rect 65450 79310 65550 79440
rect 65700 79310 65800 79440
rect 65950 79310 66050 79440
rect 66200 79310 66300 79440
rect 66450 79310 66550 79440
rect 66700 79310 66800 79440
rect 66950 79310 67050 79440
rect 67200 79310 67300 79440
rect 67450 79310 67550 79440
rect 67700 79310 67800 79440
rect 67950 79310 68050 79440
rect 68200 79310 68300 79440
rect 68450 79310 68550 79440
rect 68700 79310 68800 79440
rect 68950 79310 69050 79440
rect 69200 79310 69300 79440
rect 69450 79310 69550 79440
rect 69700 79310 69800 79440
rect 69950 79310 70050 79440
rect 70200 79310 70300 79440
rect 70450 79310 70550 79440
rect 70700 79310 70800 79440
rect 70950 79310 71000 79440
rect 59000 79300 59060 79310
rect 59190 79300 59310 79310
rect 59440 79300 59560 79310
rect 59690 79300 59810 79310
rect 59940 79300 60060 79310
rect 60190 79300 60310 79310
rect 60440 79300 60560 79310
rect 60690 79300 60810 79310
rect 60940 79300 61060 79310
rect 61190 79300 61310 79310
rect 61440 79300 61560 79310
rect 61690 79300 61810 79310
rect 61940 79300 62060 79310
rect 62190 79300 62310 79310
rect 62440 79300 62560 79310
rect 62690 79300 62810 79310
rect 62940 79300 63060 79310
rect 63190 79300 63310 79310
rect 63440 79300 63560 79310
rect 63690 79300 63810 79310
rect 63940 79300 64060 79310
rect 64190 79300 64310 79310
rect 64440 79300 64560 79310
rect 64690 79300 64810 79310
rect 64940 79300 65060 79310
rect 65190 79300 65310 79310
rect 65440 79300 65560 79310
rect 65690 79300 65810 79310
rect 65940 79300 66060 79310
rect 66190 79300 66310 79310
rect 66440 79300 66560 79310
rect 66690 79300 66810 79310
rect 66940 79300 67060 79310
rect 67190 79300 67310 79310
rect 67440 79300 67560 79310
rect 67690 79300 67810 79310
rect 67940 79300 68060 79310
rect 68190 79300 68310 79310
rect 68440 79300 68560 79310
rect 68690 79300 68810 79310
rect 68940 79300 69060 79310
rect 69190 79300 69310 79310
rect 69440 79300 69560 79310
rect 69690 79300 69810 79310
rect 69940 79300 70060 79310
rect 70190 79300 70310 79310
rect 70440 79300 70560 79310
rect 70690 79300 70810 79310
rect 70940 79300 71000 79310
rect 59000 79200 71000 79300
rect 59000 79190 59060 79200
rect 59190 79190 59310 79200
rect 59440 79190 59560 79200
rect 59690 79190 59810 79200
rect 59940 79190 60060 79200
rect 60190 79190 60310 79200
rect 60440 79190 60560 79200
rect 60690 79190 60810 79200
rect 60940 79190 61060 79200
rect 61190 79190 61310 79200
rect 61440 79190 61560 79200
rect 61690 79190 61810 79200
rect 61940 79190 62060 79200
rect 62190 79190 62310 79200
rect 62440 79190 62560 79200
rect 62690 79190 62810 79200
rect 62940 79190 63060 79200
rect 63190 79190 63310 79200
rect 63440 79190 63560 79200
rect 63690 79190 63810 79200
rect 63940 79190 64060 79200
rect 64190 79190 64310 79200
rect 64440 79190 64560 79200
rect 64690 79190 64810 79200
rect 64940 79190 65060 79200
rect 65190 79190 65310 79200
rect 65440 79190 65560 79200
rect 65690 79190 65810 79200
rect 65940 79190 66060 79200
rect 66190 79190 66310 79200
rect 66440 79190 66560 79200
rect 66690 79190 66810 79200
rect 66940 79190 67060 79200
rect 67190 79190 67310 79200
rect 67440 79190 67560 79200
rect 67690 79190 67810 79200
rect 67940 79190 68060 79200
rect 68190 79190 68310 79200
rect 68440 79190 68560 79200
rect 68690 79190 68810 79200
rect 68940 79190 69060 79200
rect 69190 79190 69310 79200
rect 69440 79190 69560 79200
rect 69690 79190 69810 79200
rect 69940 79190 70060 79200
rect 70190 79190 70310 79200
rect 70440 79190 70560 79200
rect 70690 79190 70810 79200
rect 70940 79190 71000 79200
rect 59000 79060 59050 79190
rect 59200 79060 59300 79190
rect 59450 79060 59550 79190
rect 59700 79060 59800 79190
rect 59950 79060 60050 79190
rect 60200 79060 60300 79190
rect 60450 79060 60550 79190
rect 60700 79060 60800 79190
rect 60950 79060 61050 79190
rect 61200 79060 61300 79190
rect 61450 79060 61550 79190
rect 61700 79060 61800 79190
rect 61950 79060 62050 79190
rect 62200 79060 62300 79190
rect 62450 79060 62550 79190
rect 62700 79060 62800 79190
rect 62950 79060 63050 79190
rect 63200 79060 63300 79190
rect 63450 79060 63550 79190
rect 63700 79060 63800 79190
rect 63950 79060 64050 79190
rect 64200 79060 64300 79190
rect 64450 79060 64550 79190
rect 64700 79060 64800 79190
rect 64950 79060 65050 79190
rect 65200 79060 65300 79190
rect 65450 79060 65550 79190
rect 65700 79060 65800 79190
rect 65950 79060 66050 79190
rect 66200 79060 66300 79190
rect 66450 79060 66550 79190
rect 66700 79060 66800 79190
rect 66950 79060 67050 79190
rect 67200 79060 67300 79190
rect 67450 79060 67550 79190
rect 67700 79060 67800 79190
rect 67950 79060 68050 79190
rect 68200 79060 68300 79190
rect 68450 79060 68550 79190
rect 68700 79060 68800 79190
rect 68950 79060 69050 79190
rect 69200 79060 69300 79190
rect 69450 79060 69550 79190
rect 69700 79060 69800 79190
rect 69950 79060 70050 79190
rect 70200 79060 70300 79190
rect 70450 79060 70550 79190
rect 70700 79060 70800 79190
rect 70950 79060 71000 79190
rect 59000 79050 59060 79060
rect 59190 79050 59310 79060
rect 59440 79050 59560 79060
rect 59690 79050 59810 79060
rect 59940 79050 60060 79060
rect 60190 79050 60310 79060
rect 60440 79050 60560 79060
rect 60690 79050 60810 79060
rect 60940 79050 61060 79060
rect 61190 79050 61310 79060
rect 61440 79050 61560 79060
rect 61690 79050 61810 79060
rect 61940 79050 62060 79060
rect 62190 79050 62310 79060
rect 62440 79050 62560 79060
rect 62690 79050 62810 79060
rect 62940 79050 63060 79060
rect 63190 79050 63310 79060
rect 63440 79050 63560 79060
rect 63690 79050 63810 79060
rect 63940 79050 64060 79060
rect 64190 79050 64310 79060
rect 64440 79050 64560 79060
rect 64690 79050 64810 79060
rect 64940 79050 65060 79060
rect 65190 79050 65310 79060
rect 65440 79050 65560 79060
rect 65690 79050 65810 79060
rect 65940 79050 66060 79060
rect 66190 79050 66310 79060
rect 66440 79050 66560 79060
rect 66690 79050 66810 79060
rect 66940 79050 67060 79060
rect 67190 79050 67310 79060
rect 67440 79050 67560 79060
rect 67690 79050 67810 79060
rect 67940 79050 68060 79060
rect 68190 79050 68310 79060
rect 68440 79050 68560 79060
rect 68690 79050 68810 79060
rect 68940 79050 69060 79060
rect 69190 79050 69310 79060
rect 69440 79050 69560 79060
rect 69690 79050 69810 79060
rect 69940 79050 70060 79060
rect 70190 79050 70310 79060
rect 70440 79050 70560 79060
rect 70690 79050 70810 79060
rect 70940 79050 71000 79060
rect 59000 78950 71000 79050
rect 59000 78940 59060 78950
rect 59190 78940 59310 78950
rect 59440 78940 59560 78950
rect 59690 78940 59810 78950
rect 59940 78940 60060 78950
rect 60190 78940 60310 78950
rect 60440 78940 60560 78950
rect 60690 78940 60810 78950
rect 60940 78940 61060 78950
rect 61190 78940 61310 78950
rect 61440 78940 61560 78950
rect 61690 78940 61810 78950
rect 61940 78940 62060 78950
rect 62190 78940 62310 78950
rect 62440 78940 62560 78950
rect 62690 78940 62810 78950
rect 62940 78940 63060 78950
rect 63190 78940 63310 78950
rect 63440 78940 63560 78950
rect 63690 78940 63810 78950
rect 63940 78940 64060 78950
rect 64190 78940 64310 78950
rect 64440 78940 64560 78950
rect 64690 78940 64810 78950
rect 64940 78940 65060 78950
rect 65190 78940 65310 78950
rect 65440 78940 65560 78950
rect 65690 78940 65810 78950
rect 65940 78940 66060 78950
rect 66190 78940 66310 78950
rect 66440 78940 66560 78950
rect 66690 78940 66810 78950
rect 66940 78940 67060 78950
rect 67190 78940 67310 78950
rect 67440 78940 67560 78950
rect 67690 78940 67810 78950
rect 67940 78940 68060 78950
rect 68190 78940 68310 78950
rect 68440 78940 68560 78950
rect 68690 78940 68810 78950
rect 68940 78940 69060 78950
rect 69190 78940 69310 78950
rect 69440 78940 69560 78950
rect 69690 78940 69810 78950
rect 69940 78940 70060 78950
rect 70190 78940 70310 78950
rect 70440 78940 70560 78950
rect 70690 78940 70810 78950
rect 70940 78940 71000 78950
rect 59000 78810 59050 78940
rect 59200 78810 59300 78940
rect 59450 78810 59550 78940
rect 59700 78810 59800 78940
rect 59950 78810 60050 78940
rect 60200 78810 60300 78940
rect 60450 78810 60550 78940
rect 60700 78810 60800 78940
rect 60950 78810 61050 78940
rect 61200 78810 61300 78940
rect 61450 78810 61550 78940
rect 61700 78810 61800 78940
rect 61950 78810 62050 78940
rect 62200 78810 62300 78940
rect 62450 78810 62550 78940
rect 62700 78810 62800 78940
rect 62950 78810 63050 78940
rect 63200 78810 63300 78940
rect 63450 78810 63550 78940
rect 63700 78810 63800 78940
rect 63950 78810 64050 78940
rect 64200 78810 64300 78940
rect 64450 78810 64550 78940
rect 64700 78810 64800 78940
rect 64950 78810 65050 78940
rect 65200 78810 65300 78940
rect 65450 78810 65550 78940
rect 65700 78810 65800 78940
rect 65950 78810 66050 78940
rect 66200 78810 66300 78940
rect 66450 78810 66550 78940
rect 66700 78810 66800 78940
rect 66950 78810 67050 78940
rect 67200 78810 67300 78940
rect 67450 78810 67550 78940
rect 67700 78810 67800 78940
rect 67950 78810 68050 78940
rect 68200 78810 68300 78940
rect 68450 78810 68550 78940
rect 68700 78810 68800 78940
rect 68950 78810 69050 78940
rect 69200 78810 69300 78940
rect 69450 78810 69550 78940
rect 69700 78810 69800 78940
rect 69950 78810 70050 78940
rect 70200 78810 70300 78940
rect 70450 78810 70550 78940
rect 70700 78810 70800 78940
rect 70950 78810 71000 78940
rect 59000 78800 59060 78810
rect 59190 78800 59310 78810
rect 59440 78800 59560 78810
rect 59690 78800 59810 78810
rect 59940 78800 60060 78810
rect 60190 78800 60310 78810
rect 60440 78800 60560 78810
rect 60690 78800 60810 78810
rect 60940 78800 61060 78810
rect 61190 78800 61310 78810
rect 61440 78800 61560 78810
rect 61690 78800 61810 78810
rect 61940 78800 62060 78810
rect 62190 78800 62310 78810
rect 62440 78800 62560 78810
rect 62690 78800 62810 78810
rect 62940 78800 63060 78810
rect 63190 78800 63310 78810
rect 63440 78800 63560 78810
rect 63690 78800 63810 78810
rect 63940 78800 64060 78810
rect 64190 78800 64310 78810
rect 64440 78800 64560 78810
rect 64690 78800 64810 78810
rect 64940 78800 65060 78810
rect 65190 78800 65310 78810
rect 65440 78800 65560 78810
rect 65690 78800 65810 78810
rect 65940 78800 66060 78810
rect 66190 78800 66310 78810
rect 66440 78800 66560 78810
rect 66690 78800 66810 78810
rect 66940 78800 67060 78810
rect 67190 78800 67310 78810
rect 67440 78800 67560 78810
rect 67690 78800 67810 78810
rect 67940 78800 68060 78810
rect 68190 78800 68310 78810
rect 68440 78800 68560 78810
rect 68690 78800 68810 78810
rect 68940 78800 69060 78810
rect 69190 78800 69310 78810
rect 69440 78800 69560 78810
rect 69690 78800 69810 78810
rect 69940 78800 70060 78810
rect 70190 78800 70310 78810
rect 70440 78800 70560 78810
rect 70690 78800 70810 78810
rect 70940 78800 71000 78810
rect 59000 78700 71000 78800
rect 59000 78690 59060 78700
rect 59190 78690 59310 78700
rect 59440 78690 59560 78700
rect 59690 78690 59810 78700
rect 59940 78690 60060 78700
rect 60190 78690 60310 78700
rect 60440 78690 60560 78700
rect 60690 78690 60810 78700
rect 60940 78690 61060 78700
rect 61190 78690 61310 78700
rect 61440 78690 61560 78700
rect 61690 78690 61810 78700
rect 61940 78690 62060 78700
rect 62190 78690 62310 78700
rect 62440 78690 62560 78700
rect 62690 78690 62810 78700
rect 62940 78690 63060 78700
rect 63190 78690 63310 78700
rect 63440 78690 63560 78700
rect 63690 78690 63810 78700
rect 63940 78690 64060 78700
rect 64190 78690 64310 78700
rect 64440 78690 64560 78700
rect 64690 78690 64810 78700
rect 64940 78690 65060 78700
rect 65190 78690 65310 78700
rect 65440 78690 65560 78700
rect 65690 78690 65810 78700
rect 65940 78690 66060 78700
rect 66190 78690 66310 78700
rect 66440 78690 66560 78700
rect 66690 78690 66810 78700
rect 66940 78690 67060 78700
rect 67190 78690 67310 78700
rect 67440 78690 67560 78700
rect 67690 78690 67810 78700
rect 67940 78690 68060 78700
rect 68190 78690 68310 78700
rect 68440 78690 68560 78700
rect 68690 78690 68810 78700
rect 68940 78690 69060 78700
rect 69190 78690 69310 78700
rect 69440 78690 69560 78700
rect 69690 78690 69810 78700
rect 69940 78690 70060 78700
rect 70190 78690 70310 78700
rect 70440 78690 70560 78700
rect 70690 78690 70810 78700
rect 70940 78690 71000 78700
rect 59000 78560 59050 78690
rect 59200 78560 59300 78690
rect 59450 78560 59550 78690
rect 59700 78560 59800 78690
rect 59950 78560 60050 78690
rect 60200 78560 60300 78690
rect 60450 78560 60550 78690
rect 60700 78560 60800 78690
rect 60950 78560 61050 78690
rect 61200 78560 61300 78690
rect 61450 78560 61550 78690
rect 61700 78560 61800 78690
rect 61950 78560 62050 78690
rect 62200 78560 62300 78690
rect 62450 78560 62550 78690
rect 62700 78560 62800 78690
rect 62950 78560 63050 78690
rect 63200 78560 63300 78690
rect 63450 78560 63550 78690
rect 63700 78560 63800 78690
rect 63950 78560 64050 78690
rect 64200 78560 64300 78690
rect 64450 78560 64550 78690
rect 64700 78560 64800 78690
rect 64950 78560 65050 78690
rect 65200 78560 65300 78690
rect 65450 78560 65550 78690
rect 65700 78560 65800 78690
rect 65950 78560 66050 78690
rect 66200 78560 66300 78690
rect 66450 78560 66550 78690
rect 66700 78560 66800 78690
rect 66950 78560 67050 78690
rect 67200 78560 67300 78690
rect 67450 78560 67550 78690
rect 67700 78560 67800 78690
rect 67950 78560 68050 78690
rect 68200 78560 68300 78690
rect 68450 78560 68550 78690
rect 68700 78560 68800 78690
rect 68950 78560 69050 78690
rect 69200 78560 69300 78690
rect 69450 78560 69550 78690
rect 69700 78560 69800 78690
rect 69950 78560 70050 78690
rect 70200 78560 70300 78690
rect 70450 78560 70550 78690
rect 70700 78560 70800 78690
rect 70950 78560 71000 78690
rect 59000 78550 59060 78560
rect 59190 78550 59310 78560
rect 59440 78550 59560 78560
rect 59690 78550 59810 78560
rect 59940 78550 60060 78560
rect 60190 78550 60310 78560
rect 60440 78550 60560 78560
rect 60690 78550 60810 78560
rect 60940 78550 61060 78560
rect 61190 78550 61310 78560
rect 61440 78550 61560 78560
rect 61690 78550 61810 78560
rect 61940 78550 62060 78560
rect 62190 78550 62310 78560
rect 62440 78550 62560 78560
rect 62690 78550 62810 78560
rect 62940 78550 63060 78560
rect 63190 78550 63310 78560
rect 63440 78550 63560 78560
rect 63690 78550 63810 78560
rect 63940 78550 64060 78560
rect 64190 78550 64310 78560
rect 64440 78550 64560 78560
rect 64690 78550 64810 78560
rect 64940 78550 65060 78560
rect 65190 78550 65310 78560
rect 65440 78550 65560 78560
rect 65690 78550 65810 78560
rect 65940 78550 66060 78560
rect 66190 78550 66310 78560
rect 66440 78550 66560 78560
rect 66690 78550 66810 78560
rect 66940 78550 67060 78560
rect 67190 78550 67310 78560
rect 67440 78550 67560 78560
rect 67690 78550 67810 78560
rect 67940 78550 68060 78560
rect 68190 78550 68310 78560
rect 68440 78550 68560 78560
rect 68690 78550 68810 78560
rect 68940 78550 69060 78560
rect 69190 78550 69310 78560
rect 69440 78550 69560 78560
rect 69690 78550 69810 78560
rect 69940 78550 70060 78560
rect 70190 78550 70310 78560
rect 70440 78550 70560 78560
rect 70690 78550 70810 78560
rect 70940 78550 71000 78560
rect 59000 78450 71000 78550
rect 59000 78440 59060 78450
rect 59190 78440 59310 78450
rect 59440 78440 59560 78450
rect 59690 78440 59810 78450
rect 59940 78440 60060 78450
rect 60190 78440 60310 78450
rect 60440 78440 60560 78450
rect 60690 78440 60810 78450
rect 60940 78440 61060 78450
rect 61190 78440 61310 78450
rect 61440 78440 61560 78450
rect 61690 78440 61810 78450
rect 61940 78440 62060 78450
rect 62190 78440 62310 78450
rect 62440 78440 62560 78450
rect 62690 78440 62810 78450
rect 62940 78440 63060 78450
rect 63190 78440 63310 78450
rect 63440 78440 63560 78450
rect 63690 78440 63810 78450
rect 63940 78440 64060 78450
rect 64190 78440 64310 78450
rect 64440 78440 64560 78450
rect 64690 78440 64810 78450
rect 64940 78440 65060 78450
rect 65190 78440 65310 78450
rect 65440 78440 65560 78450
rect 65690 78440 65810 78450
rect 65940 78440 66060 78450
rect 66190 78440 66310 78450
rect 66440 78440 66560 78450
rect 66690 78440 66810 78450
rect 66940 78440 67060 78450
rect 67190 78440 67310 78450
rect 67440 78440 67560 78450
rect 67690 78440 67810 78450
rect 67940 78440 68060 78450
rect 68190 78440 68310 78450
rect 68440 78440 68560 78450
rect 68690 78440 68810 78450
rect 68940 78440 69060 78450
rect 69190 78440 69310 78450
rect 69440 78440 69560 78450
rect 69690 78440 69810 78450
rect 69940 78440 70060 78450
rect 70190 78440 70310 78450
rect 70440 78440 70560 78450
rect 70690 78440 70810 78450
rect 70940 78440 71000 78450
rect 59000 78310 59050 78440
rect 59200 78310 59300 78440
rect 59450 78310 59550 78440
rect 59700 78310 59800 78440
rect 59950 78310 60050 78440
rect 60200 78310 60300 78440
rect 60450 78310 60550 78440
rect 60700 78310 60800 78440
rect 60950 78310 61050 78440
rect 61200 78310 61300 78440
rect 61450 78310 61550 78440
rect 61700 78310 61800 78440
rect 61950 78310 62050 78440
rect 62200 78310 62300 78440
rect 62450 78310 62550 78440
rect 62700 78310 62800 78440
rect 62950 78310 63050 78440
rect 63200 78310 63300 78440
rect 63450 78310 63550 78440
rect 63700 78310 63800 78440
rect 63950 78310 64050 78440
rect 64200 78310 64300 78440
rect 64450 78310 64550 78440
rect 64700 78310 64800 78440
rect 64950 78310 65050 78440
rect 65200 78310 65300 78440
rect 65450 78310 65550 78440
rect 65700 78310 65800 78440
rect 65950 78310 66050 78440
rect 66200 78310 66300 78440
rect 66450 78310 66550 78440
rect 66700 78310 66800 78440
rect 66950 78310 67050 78440
rect 67200 78310 67300 78440
rect 67450 78310 67550 78440
rect 67700 78310 67800 78440
rect 67950 78310 68050 78440
rect 68200 78310 68300 78440
rect 68450 78310 68550 78440
rect 68700 78310 68800 78440
rect 68950 78310 69050 78440
rect 69200 78310 69300 78440
rect 69450 78310 69550 78440
rect 69700 78310 69800 78440
rect 69950 78310 70050 78440
rect 70200 78310 70300 78440
rect 70450 78310 70550 78440
rect 70700 78310 70800 78440
rect 70950 78310 71000 78440
rect 59000 78300 59060 78310
rect 59190 78300 59310 78310
rect 59440 78300 59560 78310
rect 59690 78300 59810 78310
rect 59940 78300 60060 78310
rect 60190 78300 60310 78310
rect 60440 78300 60560 78310
rect 60690 78300 60810 78310
rect 60940 78300 61060 78310
rect 61190 78300 61310 78310
rect 61440 78300 61560 78310
rect 61690 78300 61810 78310
rect 61940 78300 62060 78310
rect 62190 78300 62310 78310
rect 62440 78300 62560 78310
rect 62690 78300 62810 78310
rect 62940 78300 63060 78310
rect 63190 78300 63310 78310
rect 63440 78300 63560 78310
rect 63690 78300 63810 78310
rect 63940 78300 64060 78310
rect 64190 78300 64310 78310
rect 64440 78300 64560 78310
rect 64690 78300 64810 78310
rect 64940 78300 65060 78310
rect 65190 78300 65310 78310
rect 65440 78300 65560 78310
rect 65690 78300 65810 78310
rect 65940 78300 66060 78310
rect 66190 78300 66310 78310
rect 66440 78300 66560 78310
rect 66690 78300 66810 78310
rect 66940 78300 67060 78310
rect 67190 78300 67310 78310
rect 67440 78300 67560 78310
rect 67690 78300 67810 78310
rect 67940 78300 68060 78310
rect 68190 78300 68310 78310
rect 68440 78300 68560 78310
rect 68690 78300 68810 78310
rect 68940 78300 69060 78310
rect 69190 78300 69310 78310
rect 69440 78300 69560 78310
rect 69690 78300 69810 78310
rect 69940 78300 70060 78310
rect 70190 78300 70310 78310
rect 70440 78300 70560 78310
rect 70690 78300 70810 78310
rect 70940 78300 71000 78310
rect 59000 78200 71000 78300
rect 59000 78190 59060 78200
rect 59190 78190 59310 78200
rect 59440 78190 59560 78200
rect 59690 78190 59810 78200
rect 59940 78190 60060 78200
rect 60190 78190 60310 78200
rect 60440 78190 60560 78200
rect 60690 78190 60810 78200
rect 60940 78190 61060 78200
rect 61190 78190 61310 78200
rect 61440 78190 61560 78200
rect 61690 78190 61810 78200
rect 61940 78190 62060 78200
rect 62190 78190 62310 78200
rect 62440 78190 62560 78200
rect 62690 78190 62810 78200
rect 62940 78190 63060 78200
rect 63190 78190 63310 78200
rect 63440 78190 63560 78200
rect 63690 78190 63810 78200
rect 63940 78190 64060 78200
rect 64190 78190 64310 78200
rect 64440 78190 64560 78200
rect 64690 78190 64810 78200
rect 64940 78190 65060 78200
rect 65190 78190 65310 78200
rect 65440 78190 65560 78200
rect 65690 78190 65810 78200
rect 65940 78190 66060 78200
rect 66190 78190 66310 78200
rect 66440 78190 66560 78200
rect 66690 78190 66810 78200
rect 66940 78190 67060 78200
rect 67190 78190 67310 78200
rect 67440 78190 67560 78200
rect 67690 78190 67810 78200
rect 67940 78190 68060 78200
rect 68190 78190 68310 78200
rect 68440 78190 68560 78200
rect 68690 78190 68810 78200
rect 68940 78190 69060 78200
rect 69190 78190 69310 78200
rect 69440 78190 69560 78200
rect 69690 78190 69810 78200
rect 69940 78190 70060 78200
rect 70190 78190 70310 78200
rect 70440 78190 70560 78200
rect 70690 78190 70810 78200
rect 70940 78190 71000 78200
rect 59000 78060 59050 78190
rect 59200 78060 59300 78190
rect 59450 78060 59550 78190
rect 59700 78060 59800 78190
rect 59950 78060 60050 78190
rect 60200 78060 60300 78190
rect 60450 78060 60550 78190
rect 60700 78060 60800 78190
rect 60950 78060 61050 78190
rect 61200 78060 61300 78190
rect 61450 78060 61550 78190
rect 61700 78060 61800 78190
rect 61950 78060 62050 78190
rect 62200 78060 62300 78190
rect 62450 78060 62550 78190
rect 62700 78060 62800 78190
rect 62950 78060 63050 78190
rect 63200 78060 63300 78190
rect 63450 78060 63550 78190
rect 63700 78060 63800 78190
rect 63950 78060 64050 78190
rect 64200 78060 64300 78190
rect 64450 78060 64550 78190
rect 64700 78060 64800 78190
rect 64950 78060 65050 78190
rect 65200 78060 65300 78190
rect 65450 78060 65550 78190
rect 65700 78060 65800 78190
rect 65950 78060 66050 78190
rect 66200 78060 66300 78190
rect 66450 78060 66550 78190
rect 66700 78060 66800 78190
rect 66950 78060 67050 78190
rect 67200 78060 67300 78190
rect 67450 78060 67550 78190
rect 67700 78060 67800 78190
rect 67950 78060 68050 78190
rect 68200 78060 68300 78190
rect 68450 78060 68550 78190
rect 68700 78060 68800 78190
rect 68950 78060 69050 78190
rect 69200 78060 69300 78190
rect 69450 78060 69550 78190
rect 69700 78060 69800 78190
rect 69950 78060 70050 78190
rect 70200 78060 70300 78190
rect 70450 78060 70550 78190
rect 70700 78060 70800 78190
rect 70950 78060 71000 78190
rect 59000 78050 59060 78060
rect 59190 78050 59310 78060
rect 59440 78050 59560 78060
rect 59690 78050 59810 78060
rect 59940 78050 60060 78060
rect 60190 78050 60310 78060
rect 60440 78050 60560 78060
rect 60690 78050 60810 78060
rect 60940 78050 61060 78060
rect 61190 78050 61310 78060
rect 61440 78050 61560 78060
rect 61690 78050 61810 78060
rect 61940 78050 62060 78060
rect 62190 78050 62310 78060
rect 62440 78050 62560 78060
rect 62690 78050 62810 78060
rect 62940 78050 63060 78060
rect 63190 78050 63310 78060
rect 63440 78050 63560 78060
rect 63690 78050 63810 78060
rect 63940 78050 64060 78060
rect 64190 78050 64310 78060
rect 64440 78050 64560 78060
rect 64690 78050 64810 78060
rect 64940 78050 65060 78060
rect 65190 78050 65310 78060
rect 65440 78050 65560 78060
rect 65690 78050 65810 78060
rect 65940 78050 66060 78060
rect 66190 78050 66310 78060
rect 66440 78050 66560 78060
rect 66690 78050 66810 78060
rect 66940 78050 67060 78060
rect 67190 78050 67310 78060
rect 67440 78050 67560 78060
rect 67690 78050 67810 78060
rect 67940 78050 68060 78060
rect 68190 78050 68310 78060
rect 68440 78050 68560 78060
rect 68690 78050 68810 78060
rect 68940 78050 69060 78060
rect 69190 78050 69310 78060
rect 69440 78050 69560 78060
rect 69690 78050 69810 78060
rect 69940 78050 70060 78060
rect 70190 78050 70310 78060
rect 70440 78050 70560 78060
rect 70690 78050 70810 78060
rect 70940 78050 71000 78060
rect 59000 77950 71000 78050
rect 59000 77940 59060 77950
rect 59190 77940 59310 77950
rect 59440 77940 59560 77950
rect 59690 77940 59810 77950
rect 59940 77940 60060 77950
rect 60190 77940 60310 77950
rect 60440 77940 60560 77950
rect 60690 77940 60810 77950
rect 60940 77940 61060 77950
rect 61190 77940 61310 77950
rect 61440 77940 61560 77950
rect 61690 77940 61810 77950
rect 61940 77940 62060 77950
rect 62190 77940 62310 77950
rect 62440 77940 62560 77950
rect 62690 77940 62810 77950
rect 62940 77940 63060 77950
rect 63190 77940 63310 77950
rect 63440 77940 63560 77950
rect 63690 77940 63810 77950
rect 63940 77940 64060 77950
rect 64190 77940 64310 77950
rect 64440 77940 64560 77950
rect 64690 77940 64810 77950
rect 64940 77940 65060 77950
rect 65190 77940 65310 77950
rect 65440 77940 65560 77950
rect 65690 77940 65810 77950
rect 65940 77940 66060 77950
rect 66190 77940 66310 77950
rect 66440 77940 66560 77950
rect 66690 77940 66810 77950
rect 66940 77940 67060 77950
rect 67190 77940 67310 77950
rect 67440 77940 67560 77950
rect 67690 77940 67810 77950
rect 67940 77940 68060 77950
rect 68190 77940 68310 77950
rect 68440 77940 68560 77950
rect 68690 77940 68810 77950
rect 68940 77940 69060 77950
rect 69190 77940 69310 77950
rect 69440 77940 69560 77950
rect 69690 77940 69810 77950
rect 69940 77940 70060 77950
rect 70190 77940 70310 77950
rect 70440 77940 70560 77950
rect 70690 77940 70810 77950
rect 70940 77940 71000 77950
rect 59000 77810 59050 77940
rect 59200 77810 59300 77940
rect 59450 77810 59550 77940
rect 59700 77810 59800 77940
rect 59950 77810 60050 77940
rect 60200 77810 60300 77940
rect 60450 77810 60550 77940
rect 60700 77810 60800 77940
rect 60950 77810 61050 77940
rect 61200 77810 61300 77940
rect 61450 77810 61550 77940
rect 61700 77810 61800 77940
rect 61950 77810 62050 77940
rect 62200 77810 62300 77940
rect 62450 77810 62550 77940
rect 62700 77810 62800 77940
rect 62950 77810 63050 77940
rect 63200 77810 63300 77940
rect 63450 77810 63550 77940
rect 63700 77810 63800 77940
rect 63950 77810 64050 77940
rect 64200 77810 64300 77940
rect 64450 77810 64550 77940
rect 64700 77810 64800 77940
rect 64950 77810 65050 77940
rect 65200 77810 65300 77940
rect 65450 77810 65550 77940
rect 65700 77810 65800 77940
rect 65950 77810 66050 77940
rect 66200 77810 66300 77940
rect 66450 77810 66550 77940
rect 66700 77810 66800 77940
rect 66950 77810 67050 77940
rect 67200 77810 67300 77940
rect 67450 77810 67550 77940
rect 67700 77810 67800 77940
rect 67950 77810 68050 77940
rect 68200 77810 68300 77940
rect 68450 77810 68550 77940
rect 68700 77810 68800 77940
rect 68950 77810 69050 77940
rect 69200 77810 69300 77940
rect 69450 77810 69550 77940
rect 69700 77810 69800 77940
rect 69950 77810 70050 77940
rect 70200 77810 70300 77940
rect 70450 77810 70550 77940
rect 70700 77810 70800 77940
rect 70950 77810 71000 77940
rect 59000 77800 59060 77810
rect 59190 77800 59310 77810
rect 59440 77800 59560 77810
rect 59690 77800 59810 77810
rect 59940 77800 60060 77810
rect 60190 77800 60310 77810
rect 60440 77800 60560 77810
rect 60690 77800 60810 77810
rect 60940 77800 61060 77810
rect 61190 77800 61310 77810
rect 61440 77800 61560 77810
rect 61690 77800 61810 77810
rect 61940 77800 62060 77810
rect 62190 77800 62310 77810
rect 62440 77800 62560 77810
rect 62690 77800 62810 77810
rect 62940 77800 63060 77810
rect 63190 77800 63310 77810
rect 63440 77800 63560 77810
rect 63690 77800 63810 77810
rect 63940 77800 64060 77810
rect 64190 77800 64310 77810
rect 64440 77800 64560 77810
rect 64690 77800 64810 77810
rect 64940 77800 65060 77810
rect 65190 77800 65310 77810
rect 65440 77800 65560 77810
rect 65690 77800 65810 77810
rect 65940 77800 66060 77810
rect 66190 77800 66310 77810
rect 66440 77800 66560 77810
rect 66690 77800 66810 77810
rect 66940 77800 67060 77810
rect 67190 77800 67310 77810
rect 67440 77800 67560 77810
rect 67690 77800 67810 77810
rect 67940 77800 68060 77810
rect 68190 77800 68310 77810
rect 68440 77800 68560 77810
rect 68690 77800 68810 77810
rect 68940 77800 69060 77810
rect 69190 77800 69310 77810
rect 69440 77800 69560 77810
rect 69690 77800 69810 77810
rect 69940 77800 70060 77810
rect 70190 77800 70310 77810
rect 70440 77800 70560 77810
rect 70690 77800 70810 77810
rect 70940 77800 71000 77810
rect 59000 77700 71000 77800
rect 59000 77690 59060 77700
rect 59190 77690 59310 77700
rect 59440 77690 59560 77700
rect 59690 77690 59810 77700
rect 59940 77690 60060 77700
rect 60190 77690 60310 77700
rect 60440 77690 60560 77700
rect 60690 77690 60810 77700
rect 60940 77690 61060 77700
rect 61190 77690 61310 77700
rect 61440 77690 61560 77700
rect 61690 77690 61810 77700
rect 61940 77690 62060 77700
rect 62190 77690 62310 77700
rect 62440 77690 62560 77700
rect 62690 77690 62810 77700
rect 62940 77690 63060 77700
rect 63190 77690 63310 77700
rect 63440 77690 63560 77700
rect 63690 77690 63810 77700
rect 63940 77690 64060 77700
rect 64190 77690 64310 77700
rect 64440 77690 64560 77700
rect 64690 77690 64810 77700
rect 64940 77690 65060 77700
rect 65190 77690 65310 77700
rect 65440 77690 65560 77700
rect 65690 77690 65810 77700
rect 65940 77690 66060 77700
rect 66190 77690 66310 77700
rect 66440 77690 66560 77700
rect 66690 77690 66810 77700
rect 66940 77690 67060 77700
rect 67190 77690 67310 77700
rect 67440 77690 67560 77700
rect 67690 77690 67810 77700
rect 67940 77690 68060 77700
rect 68190 77690 68310 77700
rect 68440 77690 68560 77700
rect 68690 77690 68810 77700
rect 68940 77690 69060 77700
rect 69190 77690 69310 77700
rect 69440 77690 69560 77700
rect 69690 77690 69810 77700
rect 69940 77690 70060 77700
rect 70190 77690 70310 77700
rect 70440 77690 70560 77700
rect 70690 77690 70810 77700
rect 70940 77690 71000 77700
rect 59000 77560 59050 77690
rect 59200 77560 59300 77690
rect 59450 77560 59550 77690
rect 59700 77560 59800 77690
rect 59950 77560 60050 77690
rect 60200 77560 60300 77690
rect 60450 77560 60550 77690
rect 60700 77560 60800 77690
rect 60950 77560 61050 77690
rect 61200 77560 61300 77690
rect 61450 77560 61550 77690
rect 61700 77560 61800 77690
rect 61950 77560 62050 77690
rect 62200 77560 62300 77690
rect 62450 77560 62550 77690
rect 62700 77560 62800 77690
rect 62950 77560 63050 77690
rect 63200 77560 63300 77690
rect 63450 77560 63550 77690
rect 63700 77560 63800 77690
rect 63950 77560 64050 77690
rect 64200 77560 64300 77690
rect 64450 77560 64550 77690
rect 64700 77560 64800 77690
rect 64950 77560 65050 77690
rect 65200 77560 65300 77690
rect 65450 77560 65550 77690
rect 65700 77560 65800 77690
rect 65950 77560 66050 77690
rect 66200 77560 66300 77690
rect 66450 77560 66550 77690
rect 66700 77560 66800 77690
rect 66950 77560 67050 77690
rect 67200 77560 67300 77690
rect 67450 77560 67550 77690
rect 67700 77560 67800 77690
rect 67950 77560 68050 77690
rect 68200 77560 68300 77690
rect 68450 77560 68550 77690
rect 68700 77560 68800 77690
rect 68950 77560 69050 77690
rect 69200 77560 69300 77690
rect 69450 77560 69550 77690
rect 69700 77560 69800 77690
rect 69950 77560 70050 77690
rect 70200 77560 70300 77690
rect 70450 77560 70550 77690
rect 70700 77560 70800 77690
rect 70950 77560 71000 77690
rect 59000 77550 59060 77560
rect 59190 77550 59310 77560
rect 59440 77550 59560 77560
rect 59690 77550 59810 77560
rect 59940 77550 60060 77560
rect 60190 77550 60310 77560
rect 60440 77550 60560 77560
rect 60690 77550 60810 77560
rect 60940 77550 61060 77560
rect 61190 77550 61310 77560
rect 61440 77550 61560 77560
rect 61690 77550 61810 77560
rect 61940 77550 62060 77560
rect 62190 77550 62310 77560
rect 62440 77550 62560 77560
rect 62690 77550 62810 77560
rect 62940 77550 63060 77560
rect 63190 77550 63310 77560
rect 63440 77550 63560 77560
rect 63690 77550 63810 77560
rect 63940 77550 64060 77560
rect 64190 77550 64310 77560
rect 64440 77550 64560 77560
rect 64690 77550 64810 77560
rect 64940 77550 65060 77560
rect 65190 77550 65310 77560
rect 65440 77550 65560 77560
rect 65690 77550 65810 77560
rect 65940 77550 66060 77560
rect 66190 77550 66310 77560
rect 66440 77550 66560 77560
rect 66690 77550 66810 77560
rect 66940 77550 67060 77560
rect 67190 77550 67310 77560
rect 67440 77550 67560 77560
rect 67690 77550 67810 77560
rect 67940 77550 68060 77560
rect 68190 77550 68310 77560
rect 68440 77550 68560 77560
rect 68690 77550 68810 77560
rect 68940 77550 69060 77560
rect 69190 77550 69310 77560
rect 69440 77550 69560 77560
rect 69690 77550 69810 77560
rect 69940 77550 70060 77560
rect 70190 77550 70310 77560
rect 70440 77550 70560 77560
rect 70690 77550 70810 77560
rect 70940 77550 71000 77560
rect 59000 77450 71000 77550
rect 59000 77440 59060 77450
rect 59190 77440 59310 77450
rect 59440 77440 59560 77450
rect 59690 77440 59810 77450
rect 59940 77440 60060 77450
rect 60190 77440 60310 77450
rect 60440 77440 60560 77450
rect 60690 77440 60810 77450
rect 60940 77440 61060 77450
rect 61190 77440 61310 77450
rect 61440 77440 61560 77450
rect 61690 77440 61810 77450
rect 61940 77440 62060 77450
rect 62190 77440 62310 77450
rect 62440 77440 62560 77450
rect 62690 77440 62810 77450
rect 62940 77440 63060 77450
rect 63190 77440 63310 77450
rect 63440 77440 63560 77450
rect 63690 77440 63810 77450
rect 63940 77440 64060 77450
rect 64190 77440 64310 77450
rect 64440 77440 64560 77450
rect 64690 77440 64810 77450
rect 64940 77440 65060 77450
rect 65190 77440 65310 77450
rect 65440 77440 65560 77450
rect 65690 77440 65810 77450
rect 65940 77440 66060 77450
rect 66190 77440 66310 77450
rect 66440 77440 66560 77450
rect 66690 77440 66810 77450
rect 66940 77440 67060 77450
rect 67190 77440 67310 77450
rect 67440 77440 67560 77450
rect 67690 77440 67810 77450
rect 67940 77440 68060 77450
rect 68190 77440 68310 77450
rect 68440 77440 68560 77450
rect 68690 77440 68810 77450
rect 68940 77440 69060 77450
rect 69190 77440 69310 77450
rect 69440 77440 69560 77450
rect 69690 77440 69810 77450
rect 69940 77440 70060 77450
rect 70190 77440 70310 77450
rect 70440 77440 70560 77450
rect 70690 77440 70810 77450
rect 70940 77440 71000 77450
rect 59000 77310 59050 77440
rect 59200 77310 59300 77440
rect 59450 77310 59550 77440
rect 59700 77310 59800 77440
rect 59950 77310 60050 77440
rect 60200 77310 60300 77440
rect 60450 77310 60550 77440
rect 60700 77310 60800 77440
rect 60950 77310 61050 77440
rect 61200 77310 61300 77440
rect 61450 77310 61550 77440
rect 61700 77310 61800 77440
rect 61950 77310 62050 77440
rect 62200 77310 62300 77440
rect 62450 77310 62550 77440
rect 62700 77310 62800 77440
rect 62950 77310 63050 77440
rect 63200 77310 63300 77440
rect 63450 77310 63550 77440
rect 63700 77310 63800 77440
rect 63950 77310 64050 77440
rect 64200 77310 64300 77440
rect 64450 77310 64550 77440
rect 64700 77310 64800 77440
rect 64950 77310 65050 77440
rect 65200 77310 65300 77440
rect 65450 77310 65550 77440
rect 65700 77310 65800 77440
rect 65950 77310 66050 77440
rect 66200 77310 66300 77440
rect 66450 77310 66550 77440
rect 66700 77310 66800 77440
rect 66950 77310 67050 77440
rect 67200 77310 67300 77440
rect 67450 77310 67550 77440
rect 67700 77310 67800 77440
rect 67950 77310 68050 77440
rect 68200 77310 68300 77440
rect 68450 77310 68550 77440
rect 68700 77310 68800 77440
rect 68950 77310 69050 77440
rect 69200 77310 69300 77440
rect 69450 77310 69550 77440
rect 69700 77310 69800 77440
rect 69950 77310 70050 77440
rect 70200 77310 70300 77440
rect 70450 77310 70550 77440
rect 70700 77310 70800 77440
rect 70950 77310 71000 77440
rect 59000 77300 59060 77310
rect 59190 77300 59310 77310
rect 59440 77300 59560 77310
rect 59690 77300 59810 77310
rect 59940 77300 60060 77310
rect 60190 77300 60310 77310
rect 60440 77300 60560 77310
rect 60690 77300 60810 77310
rect 60940 77300 61060 77310
rect 61190 77300 61310 77310
rect 61440 77300 61560 77310
rect 61690 77300 61810 77310
rect 61940 77300 62060 77310
rect 62190 77300 62310 77310
rect 62440 77300 62560 77310
rect 62690 77300 62810 77310
rect 62940 77300 63060 77310
rect 63190 77300 63310 77310
rect 63440 77300 63560 77310
rect 63690 77300 63810 77310
rect 63940 77300 64060 77310
rect 64190 77300 64310 77310
rect 64440 77300 64560 77310
rect 64690 77300 64810 77310
rect 64940 77300 65060 77310
rect 65190 77300 65310 77310
rect 65440 77300 65560 77310
rect 65690 77300 65810 77310
rect 65940 77300 66060 77310
rect 66190 77300 66310 77310
rect 66440 77300 66560 77310
rect 66690 77300 66810 77310
rect 66940 77300 67060 77310
rect 67190 77300 67310 77310
rect 67440 77300 67560 77310
rect 67690 77300 67810 77310
rect 67940 77300 68060 77310
rect 68190 77300 68310 77310
rect 68440 77300 68560 77310
rect 68690 77300 68810 77310
rect 68940 77300 69060 77310
rect 69190 77300 69310 77310
rect 69440 77300 69560 77310
rect 69690 77300 69810 77310
rect 69940 77300 70060 77310
rect 70190 77300 70310 77310
rect 70440 77300 70560 77310
rect 70690 77300 70810 77310
rect 70940 77300 71000 77310
rect 59000 77200 71000 77300
rect 59000 77190 59060 77200
rect 59190 77190 59310 77200
rect 59440 77190 59560 77200
rect 59690 77190 59810 77200
rect 59940 77190 60060 77200
rect 60190 77190 60310 77200
rect 60440 77190 60560 77200
rect 60690 77190 60810 77200
rect 60940 77190 61060 77200
rect 61190 77190 61310 77200
rect 61440 77190 61560 77200
rect 61690 77190 61810 77200
rect 61940 77190 62060 77200
rect 62190 77190 62310 77200
rect 62440 77190 62560 77200
rect 62690 77190 62810 77200
rect 62940 77190 63060 77200
rect 63190 77190 63310 77200
rect 63440 77190 63560 77200
rect 63690 77190 63810 77200
rect 63940 77190 64060 77200
rect 64190 77190 64310 77200
rect 64440 77190 64560 77200
rect 64690 77190 64810 77200
rect 64940 77190 65060 77200
rect 65190 77190 65310 77200
rect 65440 77190 65560 77200
rect 65690 77190 65810 77200
rect 65940 77190 66060 77200
rect 66190 77190 66310 77200
rect 66440 77190 66560 77200
rect 66690 77190 66810 77200
rect 66940 77190 67060 77200
rect 67190 77190 67310 77200
rect 67440 77190 67560 77200
rect 67690 77190 67810 77200
rect 67940 77190 68060 77200
rect 68190 77190 68310 77200
rect 68440 77190 68560 77200
rect 68690 77190 68810 77200
rect 68940 77190 69060 77200
rect 69190 77190 69310 77200
rect 69440 77190 69560 77200
rect 69690 77190 69810 77200
rect 69940 77190 70060 77200
rect 70190 77190 70310 77200
rect 70440 77190 70560 77200
rect 70690 77190 70810 77200
rect 70940 77190 71000 77200
rect 59000 77060 59050 77190
rect 59200 77060 59300 77190
rect 59450 77060 59550 77190
rect 59700 77060 59800 77190
rect 59950 77060 60050 77190
rect 60200 77060 60300 77190
rect 60450 77060 60550 77190
rect 60700 77060 60800 77190
rect 60950 77060 61050 77190
rect 61200 77060 61300 77190
rect 61450 77060 61550 77190
rect 61700 77060 61800 77190
rect 61950 77060 62050 77190
rect 62200 77060 62300 77190
rect 62450 77060 62550 77190
rect 62700 77060 62800 77190
rect 62950 77060 63050 77190
rect 63200 77060 63300 77190
rect 63450 77060 63550 77190
rect 63700 77060 63800 77190
rect 63950 77060 64050 77190
rect 64200 77060 64300 77190
rect 64450 77060 64550 77190
rect 64700 77060 64800 77190
rect 64950 77060 65050 77190
rect 65200 77060 65300 77190
rect 65450 77060 65550 77190
rect 65700 77060 65800 77190
rect 65950 77060 66050 77190
rect 66200 77060 66300 77190
rect 66450 77060 66550 77190
rect 66700 77060 66800 77190
rect 66950 77060 67050 77190
rect 67200 77060 67300 77190
rect 67450 77060 67550 77190
rect 67700 77060 67800 77190
rect 67950 77060 68050 77190
rect 68200 77060 68300 77190
rect 68450 77060 68550 77190
rect 68700 77060 68800 77190
rect 68950 77060 69050 77190
rect 69200 77060 69300 77190
rect 69450 77060 69550 77190
rect 69700 77060 69800 77190
rect 69950 77060 70050 77190
rect 70200 77060 70300 77190
rect 70450 77060 70550 77190
rect 70700 77060 70800 77190
rect 70950 77060 71000 77190
rect 59000 77050 59060 77060
rect 59190 77050 59310 77060
rect 59440 77050 59560 77060
rect 59690 77050 59810 77060
rect 59940 77050 60060 77060
rect 60190 77050 60310 77060
rect 60440 77050 60560 77060
rect 60690 77050 60810 77060
rect 60940 77050 61060 77060
rect 61190 77050 61310 77060
rect 61440 77050 61560 77060
rect 61690 77050 61810 77060
rect 61940 77050 62060 77060
rect 62190 77050 62310 77060
rect 62440 77050 62560 77060
rect 62690 77050 62810 77060
rect 62940 77050 63060 77060
rect 63190 77050 63310 77060
rect 63440 77050 63560 77060
rect 63690 77050 63810 77060
rect 63940 77050 64060 77060
rect 64190 77050 64310 77060
rect 64440 77050 64560 77060
rect 64690 77050 64810 77060
rect 64940 77050 65060 77060
rect 65190 77050 65310 77060
rect 65440 77050 65560 77060
rect 65690 77050 65810 77060
rect 65940 77050 66060 77060
rect 66190 77050 66310 77060
rect 66440 77050 66560 77060
rect 66690 77050 66810 77060
rect 66940 77050 67060 77060
rect 67190 77050 67310 77060
rect 67440 77050 67560 77060
rect 67690 77050 67810 77060
rect 67940 77050 68060 77060
rect 68190 77050 68310 77060
rect 68440 77050 68560 77060
rect 68690 77050 68810 77060
rect 68940 77050 69060 77060
rect 69190 77050 69310 77060
rect 69440 77050 69560 77060
rect 69690 77050 69810 77060
rect 69940 77050 70060 77060
rect 70190 77050 70310 77060
rect 70440 77050 70560 77060
rect 70690 77050 70810 77060
rect 70940 77050 71000 77060
rect 59000 77000 71000 77050
rect 81000 80950 92000 81000
rect 81000 80940 81060 80950
rect 81190 80940 81310 80950
rect 81440 80940 81560 80950
rect 81690 80940 81810 80950
rect 81940 80940 82060 80950
rect 82190 80940 82310 80950
rect 82440 80940 82560 80950
rect 82690 80940 82810 80950
rect 82940 80940 83060 80950
rect 83190 80940 83310 80950
rect 83440 80940 83560 80950
rect 83690 80940 83810 80950
rect 83940 80940 84060 80950
rect 84190 80940 84310 80950
rect 84440 80940 84560 80950
rect 84690 80940 84810 80950
rect 84940 80940 85060 80950
rect 85190 80940 85310 80950
rect 85440 80940 85560 80950
rect 85690 80940 85810 80950
rect 85940 80940 86060 80950
rect 86190 80940 86310 80950
rect 86440 80940 86560 80950
rect 86690 80940 86810 80950
rect 86940 80940 87060 80950
rect 87190 80940 87310 80950
rect 87440 80940 87560 80950
rect 87690 80940 87810 80950
rect 87940 80940 88060 80950
rect 88190 80940 88310 80950
rect 88440 80940 88560 80950
rect 88690 80940 88810 80950
rect 88940 80940 89060 80950
rect 89190 80940 89310 80950
rect 89440 80940 89560 80950
rect 89690 80940 89810 80950
rect 89940 80940 90060 80950
rect 90190 80940 90310 80950
rect 90440 80940 90560 80950
rect 90690 80940 90810 80950
rect 90940 80940 91060 80950
rect 91190 80940 91310 80950
rect 91440 80940 91560 80950
rect 91690 80940 91810 80950
rect 91940 80940 92000 80950
rect 81000 80810 81050 80940
rect 81200 80810 81300 80940
rect 81450 80810 81550 80940
rect 81700 80810 81800 80940
rect 81950 80810 82050 80940
rect 82200 80810 82300 80940
rect 82450 80810 82550 80940
rect 82700 80810 82800 80940
rect 82950 80810 83050 80940
rect 83200 80810 83300 80940
rect 83450 80810 83550 80940
rect 83700 80810 83800 80940
rect 83950 80810 84050 80940
rect 84200 80810 84300 80940
rect 84450 80810 84550 80940
rect 84700 80810 84800 80940
rect 84950 80810 85050 80940
rect 85200 80810 85300 80940
rect 85450 80810 85550 80940
rect 85700 80810 85800 80940
rect 85950 80810 86050 80940
rect 86200 80810 86300 80940
rect 86450 80810 86550 80940
rect 86700 80810 86800 80940
rect 86950 80810 87050 80940
rect 87200 80810 87300 80940
rect 87450 80810 87550 80940
rect 87700 80810 87800 80940
rect 87950 80810 88050 80940
rect 88200 80810 88300 80940
rect 88450 80810 88550 80940
rect 88700 80810 88800 80940
rect 88950 80810 89050 80940
rect 89200 80810 89300 80940
rect 89450 80810 89550 80940
rect 89700 80810 89800 80940
rect 89950 80810 90050 80940
rect 90200 80810 90300 80940
rect 90450 80810 90550 80940
rect 90700 80810 90800 80940
rect 90950 80810 91050 80940
rect 91200 80810 91300 80940
rect 91450 80810 91550 80940
rect 91700 80810 91800 80940
rect 91950 80810 92000 80940
rect 81000 80800 81060 80810
rect 81190 80800 81310 80810
rect 81440 80800 81560 80810
rect 81690 80800 81810 80810
rect 81940 80800 82060 80810
rect 82190 80800 82310 80810
rect 82440 80800 82560 80810
rect 82690 80800 82810 80810
rect 82940 80800 83060 80810
rect 83190 80800 83310 80810
rect 83440 80800 83560 80810
rect 83690 80800 83810 80810
rect 83940 80800 84060 80810
rect 84190 80800 84310 80810
rect 84440 80800 84560 80810
rect 84690 80800 84810 80810
rect 84940 80800 85060 80810
rect 85190 80800 85310 80810
rect 85440 80800 85560 80810
rect 85690 80800 85810 80810
rect 85940 80800 86060 80810
rect 86190 80800 86310 80810
rect 86440 80800 86560 80810
rect 86690 80800 86810 80810
rect 86940 80800 87060 80810
rect 87190 80800 87310 80810
rect 87440 80800 87560 80810
rect 87690 80800 87810 80810
rect 87940 80800 88060 80810
rect 88190 80800 88310 80810
rect 88440 80800 88560 80810
rect 88690 80800 88810 80810
rect 88940 80800 89060 80810
rect 89190 80800 89310 80810
rect 89440 80800 89560 80810
rect 89690 80800 89810 80810
rect 89940 80800 90060 80810
rect 90190 80800 90310 80810
rect 90440 80800 90560 80810
rect 90690 80800 90810 80810
rect 90940 80800 91060 80810
rect 91190 80800 91310 80810
rect 91440 80800 91560 80810
rect 91690 80800 91810 80810
rect 91940 80800 92000 80810
rect 81000 80700 92000 80800
rect 81000 80690 81060 80700
rect 81190 80690 81310 80700
rect 81440 80690 81560 80700
rect 81690 80690 81810 80700
rect 81940 80690 82060 80700
rect 82190 80690 82310 80700
rect 82440 80690 82560 80700
rect 82690 80690 82810 80700
rect 82940 80690 83060 80700
rect 83190 80690 83310 80700
rect 83440 80690 83560 80700
rect 83690 80690 83810 80700
rect 83940 80690 84060 80700
rect 84190 80690 84310 80700
rect 84440 80690 84560 80700
rect 84690 80690 84810 80700
rect 84940 80690 85060 80700
rect 85190 80690 85310 80700
rect 85440 80690 85560 80700
rect 85690 80690 85810 80700
rect 85940 80690 86060 80700
rect 86190 80690 86310 80700
rect 86440 80690 86560 80700
rect 86690 80690 86810 80700
rect 86940 80690 87060 80700
rect 87190 80690 87310 80700
rect 87440 80690 87560 80700
rect 87690 80690 87810 80700
rect 87940 80690 88060 80700
rect 88190 80690 88310 80700
rect 88440 80690 88560 80700
rect 88690 80690 88810 80700
rect 88940 80690 89060 80700
rect 89190 80690 89310 80700
rect 89440 80690 89560 80700
rect 89690 80690 89810 80700
rect 89940 80690 90060 80700
rect 90190 80690 90310 80700
rect 90440 80690 90560 80700
rect 90690 80690 90810 80700
rect 90940 80690 91060 80700
rect 91190 80690 91310 80700
rect 91440 80690 91560 80700
rect 91690 80690 91810 80700
rect 91940 80690 92000 80700
rect 81000 80560 81050 80690
rect 81200 80560 81300 80690
rect 81450 80560 81550 80690
rect 81700 80560 81800 80690
rect 81950 80560 82050 80690
rect 82200 80560 82300 80690
rect 82450 80560 82550 80690
rect 82700 80560 82800 80690
rect 82950 80560 83050 80690
rect 83200 80560 83300 80690
rect 83450 80560 83550 80690
rect 83700 80560 83800 80690
rect 83950 80560 84050 80690
rect 84200 80560 84300 80690
rect 84450 80560 84550 80690
rect 84700 80560 84800 80690
rect 84950 80560 85050 80690
rect 85200 80560 85300 80690
rect 85450 80560 85550 80690
rect 85700 80560 85800 80690
rect 85950 80560 86050 80690
rect 86200 80560 86300 80690
rect 86450 80560 86550 80690
rect 86700 80560 86800 80690
rect 86950 80560 87050 80690
rect 87200 80560 87300 80690
rect 87450 80560 87550 80690
rect 87700 80560 87800 80690
rect 87950 80560 88050 80690
rect 88200 80560 88300 80690
rect 88450 80560 88550 80690
rect 88700 80560 88800 80690
rect 88950 80560 89050 80690
rect 89200 80560 89300 80690
rect 89450 80560 89550 80690
rect 89700 80560 89800 80690
rect 89950 80560 90050 80690
rect 90200 80560 90300 80690
rect 90450 80560 90550 80690
rect 90700 80560 90800 80690
rect 90950 80560 91050 80690
rect 91200 80560 91300 80690
rect 91450 80560 91550 80690
rect 91700 80560 91800 80690
rect 91950 80560 92000 80690
rect 81000 80550 81060 80560
rect 81190 80550 81310 80560
rect 81440 80550 81560 80560
rect 81690 80550 81810 80560
rect 81940 80550 82060 80560
rect 82190 80550 82310 80560
rect 82440 80550 82560 80560
rect 82690 80550 82810 80560
rect 82940 80550 83060 80560
rect 83190 80550 83310 80560
rect 83440 80550 83560 80560
rect 83690 80550 83810 80560
rect 83940 80550 84060 80560
rect 84190 80550 84310 80560
rect 84440 80550 84560 80560
rect 84690 80550 84810 80560
rect 84940 80550 85060 80560
rect 85190 80550 85310 80560
rect 85440 80550 85560 80560
rect 85690 80550 85810 80560
rect 85940 80550 86060 80560
rect 86190 80550 86310 80560
rect 86440 80550 86560 80560
rect 86690 80550 86810 80560
rect 86940 80550 87060 80560
rect 87190 80550 87310 80560
rect 87440 80550 87560 80560
rect 87690 80550 87810 80560
rect 87940 80550 88060 80560
rect 88190 80550 88310 80560
rect 88440 80550 88560 80560
rect 88690 80550 88810 80560
rect 88940 80550 89060 80560
rect 89190 80550 89310 80560
rect 89440 80550 89560 80560
rect 89690 80550 89810 80560
rect 89940 80550 90060 80560
rect 90190 80550 90310 80560
rect 90440 80550 90560 80560
rect 90690 80550 90810 80560
rect 90940 80550 91060 80560
rect 91190 80550 91310 80560
rect 91440 80550 91560 80560
rect 91690 80550 91810 80560
rect 91940 80550 92000 80560
rect 81000 80450 92000 80550
rect 81000 80440 81060 80450
rect 81190 80440 81310 80450
rect 81440 80440 81560 80450
rect 81690 80440 81810 80450
rect 81940 80440 82060 80450
rect 82190 80440 82310 80450
rect 82440 80440 82560 80450
rect 82690 80440 82810 80450
rect 82940 80440 83060 80450
rect 83190 80440 83310 80450
rect 83440 80440 83560 80450
rect 83690 80440 83810 80450
rect 83940 80440 84060 80450
rect 84190 80440 84310 80450
rect 84440 80440 84560 80450
rect 84690 80440 84810 80450
rect 84940 80440 85060 80450
rect 85190 80440 85310 80450
rect 85440 80440 85560 80450
rect 85690 80440 85810 80450
rect 85940 80440 86060 80450
rect 86190 80440 86310 80450
rect 86440 80440 86560 80450
rect 86690 80440 86810 80450
rect 86940 80440 87060 80450
rect 87190 80440 87310 80450
rect 87440 80440 87560 80450
rect 87690 80440 87810 80450
rect 87940 80440 88060 80450
rect 88190 80440 88310 80450
rect 88440 80440 88560 80450
rect 88690 80440 88810 80450
rect 88940 80440 89060 80450
rect 89190 80440 89310 80450
rect 89440 80440 89560 80450
rect 89690 80440 89810 80450
rect 89940 80440 90060 80450
rect 90190 80440 90310 80450
rect 90440 80440 90560 80450
rect 90690 80440 90810 80450
rect 90940 80440 91060 80450
rect 91190 80440 91310 80450
rect 91440 80440 91560 80450
rect 91690 80440 91810 80450
rect 91940 80440 92000 80450
rect 81000 80310 81050 80440
rect 81200 80310 81300 80440
rect 81450 80310 81550 80440
rect 81700 80310 81800 80440
rect 81950 80310 82050 80440
rect 82200 80310 82300 80440
rect 82450 80310 82550 80440
rect 82700 80310 82800 80440
rect 82950 80310 83050 80440
rect 83200 80310 83300 80440
rect 83450 80310 83550 80440
rect 83700 80310 83800 80440
rect 83950 80310 84050 80440
rect 84200 80310 84300 80440
rect 84450 80310 84550 80440
rect 84700 80310 84800 80440
rect 84950 80310 85050 80440
rect 85200 80310 85300 80440
rect 85450 80310 85550 80440
rect 85700 80310 85800 80440
rect 85950 80310 86050 80440
rect 86200 80310 86300 80440
rect 86450 80310 86550 80440
rect 86700 80310 86800 80440
rect 86950 80310 87050 80440
rect 87200 80310 87300 80440
rect 87450 80310 87550 80440
rect 87700 80310 87800 80440
rect 87950 80310 88050 80440
rect 88200 80310 88300 80440
rect 88450 80310 88550 80440
rect 88700 80310 88800 80440
rect 88950 80310 89050 80440
rect 89200 80310 89300 80440
rect 89450 80310 89550 80440
rect 89700 80310 89800 80440
rect 89950 80310 90050 80440
rect 90200 80310 90300 80440
rect 90450 80310 90550 80440
rect 90700 80310 90800 80440
rect 90950 80310 91050 80440
rect 91200 80310 91300 80440
rect 91450 80310 91550 80440
rect 91700 80310 91800 80440
rect 91950 80310 92000 80440
rect 81000 80300 81060 80310
rect 81190 80300 81310 80310
rect 81440 80300 81560 80310
rect 81690 80300 81810 80310
rect 81940 80300 82060 80310
rect 82190 80300 82310 80310
rect 82440 80300 82560 80310
rect 82690 80300 82810 80310
rect 82940 80300 83060 80310
rect 83190 80300 83310 80310
rect 83440 80300 83560 80310
rect 83690 80300 83810 80310
rect 83940 80300 84060 80310
rect 84190 80300 84310 80310
rect 84440 80300 84560 80310
rect 84690 80300 84810 80310
rect 84940 80300 85060 80310
rect 85190 80300 85310 80310
rect 85440 80300 85560 80310
rect 85690 80300 85810 80310
rect 85940 80300 86060 80310
rect 86190 80300 86310 80310
rect 86440 80300 86560 80310
rect 86690 80300 86810 80310
rect 86940 80300 87060 80310
rect 87190 80300 87310 80310
rect 87440 80300 87560 80310
rect 87690 80300 87810 80310
rect 87940 80300 88060 80310
rect 88190 80300 88310 80310
rect 88440 80300 88560 80310
rect 88690 80300 88810 80310
rect 88940 80300 89060 80310
rect 89190 80300 89310 80310
rect 89440 80300 89560 80310
rect 89690 80300 89810 80310
rect 89940 80300 90060 80310
rect 90190 80300 90310 80310
rect 90440 80300 90560 80310
rect 90690 80300 90810 80310
rect 90940 80300 91060 80310
rect 91190 80300 91310 80310
rect 91440 80300 91560 80310
rect 91690 80300 91810 80310
rect 91940 80300 92000 80310
rect 81000 80200 92000 80300
rect 81000 80190 81060 80200
rect 81190 80190 81310 80200
rect 81440 80190 81560 80200
rect 81690 80190 81810 80200
rect 81940 80190 82060 80200
rect 82190 80190 82310 80200
rect 82440 80190 82560 80200
rect 82690 80190 82810 80200
rect 82940 80190 83060 80200
rect 83190 80190 83310 80200
rect 83440 80190 83560 80200
rect 83690 80190 83810 80200
rect 83940 80190 84060 80200
rect 84190 80190 84310 80200
rect 84440 80190 84560 80200
rect 84690 80190 84810 80200
rect 84940 80190 85060 80200
rect 85190 80190 85310 80200
rect 85440 80190 85560 80200
rect 85690 80190 85810 80200
rect 85940 80190 86060 80200
rect 86190 80190 86310 80200
rect 86440 80190 86560 80200
rect 86690 80190 86810 80200
rect 86940 80190 87060 80200
rect 87190 80190 87310 80200
rect 87440 80190 87560 80200
rect 87690 80190 87810 80200
rect 87940 80190 88060 80200
rect 88190 80190 88310 80200
rect 88440 80190 88560 80200
rect 88690 80190 88810 80200
rect 88940 80190 89060 80200
rect 89190 80190 89310 80200
rect 89440 80190 89560 80200
rect 89690 80190 89810 80200
rect 89940 80190 90060 80200
rect 90190 80190 90310 80200
rect 90440 80190 90560 80200
rect 90690 80190 90810 80200
rect 90940 80190 91060 80200
rect 91190 80190 91310 80200
rect 91440 80190 91560 80200
rect 91690 80190 91810 80200
rect 91940 80190 92000 80200
rect 81000 80060 81050 80190
rect 81200 80060 81300 80190
rect 81450 80060 81550 80190
rect 81700 80060 81800 80190
rect 81950 80060 82050 80190
rect 82200 80060 82300 80190
rect 82450 80060 82550 80190
rect 82700 80060 82800 80190
rect 82950 80060 83050 80190
rect 83200 80060 83300 80190
rect 83450 80060 83550 80190
rect 83700 80060 83800 80190
rect 83950 80060 84050 80190
rect 84200 80060 84300 80190
rect 84450 80060 84550 80190
rect 84700 80060 84800 80190
rect 84950 80060 85050 80190
rect 85200 80060 85300 80190
rect 85450 80060 85550 80190
rect 85700 80060 85800 80190
rect 85950 80060 86050 80190
rect 86200 80060 86300 80190
rect 86450 80060 86550 80190
rect 86700 80060 86800 80190
rect 86950 80060 87050 80190
rect 87200 80060 87300 80190
rect 87450 80060 87550 80190
rect 87700 80060 87800 80190
rect 87950 80060 88050 80190
rect 88200 80060 88300 80190
rect 88450 80060 88550 80190
rect 88700 80060 88800 80190
rect 88950 80060 89050 80190
rect 89200 80060 89300 80190
rect 89450 80060 89550 80190
rect 89700 80060 89800 80190
rect 89950 80060 90050 80190
rect 90200 80060 90300 80190
rect 90450 80060 90550 80190
rect 90700 80060 90800 80190
rect 90950 80060 91050 80190
rect 91200 80060 91300 80190
rect 91450 80060 91550 80190
rect 91700 80060 91800 80190
rect 91950 80060 92000 80190
rect 81000 80050 81060 80060
rect 81190 80050 81310 80060
rect 81440 80050 81560 80060
rect 81690 80050 81810 80060
rect 81940 80050 82060 80060
rect 82190 80050 82310 80060
rect 82440 80050 82560 80060
rect 82690 80050 82810 80060
rect 82940 80050 83060 80060
rect 83190 80050 83310 80060
rect 83440 80050 83560 80060
rect 83690 80050 83810 80060
rect 83940 80050 84060 80060
rect 84190 80050 84310 80060
rect 84440 80050 84560 80060
rect 84690 80050 84810 80060
rect 84940 80050 85060 80060
rect 85190 80050 85310 80060
rect 85440 80050 85560 80060
rect 85690 80050 85810 80060
rect 85940 80050 86060 80060
rect 86190 80050 86310 80060
rect 86440 80050 86560 80060
rect 86690 80050 86810 80060
rect 86940 80050 87060 80060
rect 87190 80050 87310 80060
rect 87440 80050 87560 80060
rect 87690 80050 87810 80060
rect 87940 80050 88060 80060
rect 88190 80050 88310 80060
rect 88440 80050 88560 80060
rect 88690 80050 88810 80060
rect 88940 80050 89060 80060
rect 89190 80050 89310 80060
rect 89440 80050 89560 80060
rect 89690 80050 89810 80060
rect 89940 80050 90060 80060
rect 90190 80050 90310 80060
rect 90440 80050 90560 80060
rect 90690 80050 90810 80060
rect 90940 80050 91060 80060
rect 91190 80050 91310 80060
rect 91440 80050 91560 80060
rect 91690 80050 91810 80060
rect 91940 80050 92000 80060
rect 81000 79950 92000 80050
rect 81000 79940 81060 79950
rect 81190 79940 81310 79950
rect 81440 79940 81560 79950
rect 81690 79940 81810 79950
rect 81940 79940 82060 79950
rect 82190 79940 82310 79950
rect 82440 79940 82560 79950
rect 82690 79940 82810 79950
rect 82940 79940 83060 79950
rect 83190 79940 83310 79950
rect 83440 79940 83560 79950
rect 83690 79940 83810 79950
rect 83940 79940 84060 79950
rect 84190 79940 84310 79950
rect 84440 79940 84560 79950
rect 84690 79940 84810 79950
rect 84940 79940 85060 79950
rect 85190 79940 85310 79950
rect 85440 79940 85560 79950
rect 85690 79940 85810 79950
rect 85940 79940 86060 79950
rect 86190 79940 86310 79950
rect 86440 79940 86560 79950
rect 86690 79940 86810 79950
rect 86940 79940 87060 79950
rect 87190 79940 87310 79950
rect 87440 79940 87560 79950
rect 87690 79940 87810 79950
rect 87940 79940 88060 79950
rect 88190 79940 88310 79950
rect 88440 79940 88560 79950
rect 88690 79940 88810 79950
rect 88940 79940 89060 79950
rect 89190 79940 89310 79950
rect 89440 79940 89560 79950
rect 89690 79940 89810 79950
rect 89940 79940 90060 79950
rect 90190 79940 90310 79950
rect 90440 79940 90560 79950
rect 90690 79940 90810 79950
rect 90940 79940 91060 79950
rect 91190 79940 91310 79950
rect 91440 79940 91560 79950
rect 91690 79940 91810 79950
rect 91940 79940 92000 79950
rect 81000 79810 81050 79940
rect 81200 79810 81300 79940
rect 81450 79810 81550 79940
rect 81700 79810 81800 79940
rect 81950 79810 82050 79940
rect 82200 79810 82300 79940
rect 82450 79810 82550 79940
rect 82700 79810 82800 79940
rect 82950 79810 83050 79940
rect 83200 79810 83300 79940
rect 83450 79810 83550 79940
rect 83700 79810 83800 79940
rect 83950 79810 84050 79940
rect 84200 79810 84300 79940
rect 84450 79810 84550 79940
rect 84700 79810 84800 79940
rect 84950 79810 85050 79940
rect 85200 79810 85300 79940
rect 85450 79810 85550 79940
rect 85700 79810 85800 79940
rect 85950 79810 86050 79940
rect 86200 79810 86300 79940
rect 86450 79810 86550 79940
rect 86700 79810 86800 79940
rect 86950 79810 87050 79940
rect 87200 79810 87300 79940
rect 87450 79810 87550 79940
rect 87700 79810 87800 79940
rect 87950 79810 88050 79940
rect 88200 79810 88300 79940
rect 88450 79810 88550 79940
rect 88700 79810 88800 79940
rect 88950 79810 89050 79940
rect 89200 79810 89300 79940
rect 89450 79810 89550 79940
rect 89700 79810 89800 79940
rect 89950 79810 90050 79940
rect 90200 79810 90300 79940
rect 90450 79810 90550 79940
rect 90700 79810 90800 79940
rect 90950 79810 91050 79940
rect 91200 79810 91300 79940
rect 91450 79810 91550 79940
rect 91700 79810 91800 79940
rect 91950 79810 92000 79940
rect 81000 79800 81060 79810
rect 81190 79800 81310 79810
rect 81440 79800 81560 79810
rect 81690 79800 81810 79810
rect 81940 79800 82060 79810
rect 82190 79800 82310 79810
rect 82440 79800 82560 79810
rect 82690 79800 82810 79810
rect 82940 79800 83060 79810
rect 83190 79800 83310 79810
rect 83440 79800 83560 79810
rect 83690 79800 83810 79810
rect 83940 79800 84060 79810
rect 84190 79800 84310 79810
rect 84440 79800 84560 79810
rect 84690 79800 84810 79810
rect 84940 79800 85060 79810
rect 85190 79800 85310 79810
rect 85440 79800 85560 79810
rect 85690 79800 85810 79810
rect 85940 79800 86060 79810
rect 86190 79800 86310 79810
rect 86440 79800 86560 79810
rect 86690 79800 86810 79810
rect 86940 79800 87060 79810
rect 87190 79800 87310 79810
rect 87440 79800 87560 79810
rect 87690 79800 87810 79810
rect 87940 79800 88060 79810
rect 88190 79800 88310 79810
rect 88440 79800 88560 79810
rect 88690 79800 88810 79810
rect 88940 79800 89060 79810
rect 89190 79800 89310 79810
rect 89440 79800 89560 79810
rect 89690 79800 89810 79810
rect 89940 79800 90060 79810
rect 90190 79800 90310 79810
rect 90440 79800 90560 79810
rect 90690 79800 90810 79810
rect 90940 79800 91060 79810
rect 91190 79800 91310 79810
rect 91440 79800 91560 79810
rect 91690 79800 91810 79810
rect 91940 79800 92000 79810
rect 81000 79700 92000 79800
rect 81000 79690 81060 79700
rect 81190 79690 81310 79700
rect 81440 79690 81560 79700
rect 81690 79690 81810 79700
rect 81940 79690 82060 79700
rect 82190 79690 82310 79700
rect 82440 79690 82560 79700
rect 82690 79690 82810 79700
rect 82940 79690 83060 79700
rect 83190 79690 83310 79700
rect 83440 79690 83560 79700
rect 83690 79690 83810 79700
rect 83940 79690 84060 79700
rect 84190 79690 84310 79700
rect 84440 79690 84560 79700
rect 84690 79690 84810 79700
rect 84940 79690 85060 79700
rect 85190 79690 85310 79700
rect 85440 79690 85560 79700
rect 85690 79690 85810 79700
rect 85940 79690 86060 79700
rect 86190 79690 86310 79700
rect 86440 79690 86560 79700
rect 86690 79690 86810 79700
rect 86940 79690 87060 79700
rect 87190 79690 87310 79700
rect 87440 79690 87560 79700
rect 87690 79690 87810 79700
rect 87940 79690 88060 79700
rect 88190 79690 88310 79700
rect 88440 79690 88560 79700
rect 88690 79690 88810 79700
rect 88940 79690 89060 79700
rect 89190 79690 89310 79700
rect 89440 79690 89560 79700
rect 89690 79690 89810 79700
rect 89940 79690 90060 79700
rect 90190 79690 90310 79700
rect 90440 79690 90560 79700
rect 90690 79690 90810 79700
rect 90940 79690 91060 79700
rect 91190 79690 91310 79700
rect 91440 79690 91560 79700
rect 91690 79690 91810 79700
rect 91940 79690 92000 79700
rect 81000 79560 81050 79690
rect 81200 79560 81300 79690
rect 81450 79560 81550 79690
rect 81700 79560 81800 79690
rect 81950 79560 82050 79690
rect 82200 79560 82300 79690
rect 82450 79560 82550 79690
rect 82700 79560 82800 79690
rect 82950 79560 83050 79690
rect 83200 79560 83300 79690
rect 83450 79560 83550 79690
rect 83700 79560 83800 79690
rect 83950 79560 84050 79690
rect 84200 79560 84300 79690
rect 84450 79560 84550 79690
rect 84700 79560 84800 79690
rect 84950 79560 85050 79690
rect 85200 79560 85300 79690
rect 85450 79560 85550 79690
rect 85700 79560 85800 79690
rect 85950 79560 86050 79690
rect 86200 79560 86300 79690
rect 86450 79560 86550 79690
rect 86700 79560 86800 79690
rect 86950 79560 87050 79690
rect 87200 79560 87300 79690
rect 87450 79560 87550 79690
rect 87700 79560 87800 79690
rect 87950 79560 88050 79690
rect 88200 79560 88300 79690
rect 88450 79560 88550 79690
rect 88700 79560 88800 79690
rect 88950 79560 89050 79690
rect 89200 79560 89300 79690
rect 89450 79560 89550 79690
rect 89700 79560 89800 79690
rect 89950 79560 90050 79690
rect 90200 79560 90300 79690
rect 90450 79560 90550 79690
rect 90700 79560 90800 79690
rect 90950 79560 91050 79690
rect 91200 79560 91300 79690
rect 91450 79560 91550 79690
rect 91700 79560 91800 79690
rect 91950 79560 92000 79690
rect 81000 79550 81060 79560
rect 81190 79550 81310 79560
rect 81440 79550 81560 79560
rect 81690 79550 81810 79560
rect 81940 79550 82060 79560
rect 82190 79550 82310 79560
rect 82440 79550 82560 79560
rect 82690 79550 82810 79560
rect 82940 79550 83060 79560
rect 83190 79550 83310 79560
rect 83440 79550 83560 79560
rect 83690 79550 83810 79560
rect 83940 79550 84060 79560
rect 84190 79550 84310 79560
rect 84440 79550 84560 79560
rect 84690 79550 84810 79560
rect 84940 79550 85060 79560
rect 85190 79550 85310 79560
rect 85440 79550 85560 79560
rect 85690 79550 85810 79560
rect 85940 79550 86060 79560
rect 86190 79550 86310 79560
rect 86440 79550 86560 79560
rect 86690 79550 86810 79560
rect 86940 79550 87060 79560
rect 87190 79550 87310 79560
rect 87440 79550 87560 79560
rect 87690 79550 87810 79560
rect 87940 79550 88060 79560
rect 88190 79550 88310 79560
rect 88440 79550 88560 79560
rect 88690 79550 88810 79560
rect 88940 79550 89060 79560
rect 89190 79550 89310 79560
rect 89440 79550 89560 79560
rect 89690 79550 89810 79560
rect 89940 79550 90060 79560
rect 90190 79550 90310 79560
rect 90440 79550 90560 79560
rect 90690 79550 90810 79560
rect 90940 79550 91060 79560
rect 91190 79550 91310 79560
rect 91440 79550 91560 79560
rect 91690 79550 91810 79560
rect 91940 79550 92000 79560
rect 81000 79450 92000 79550
rect 81000 79440 81060 79450
rect 81190 79440 81310 79450
rect 81440 79440 81560 79450
rect 81690 79440 81810 79450
rect 81940 79440 82060 79450
rect 82190 79440 82310 79450
rect 82440 79440 82560 79450
rect 82690 79440 82810 79450
rect 82940 79440 83060 79450
rect 83190 79440 83310 79450
rect 83440 79440 83560 79450
rect 83690 79440 83810 79450
rect 83940 79440 84060 79450
rect 84190 79440 84310 79450
rect 84440 79440 84560 79450
rect 84690 79440 84810 79450
rect 84940 79440 85060 79450
rect 85190 79440 85310 79450
rect 85440 79440 85560 79450
rect 85690 79440 85810 79450
rect 85940 79440 86060 79450
rect 86190 79440 86310 79450
rect 86440 79440 86560 79450
rect 86690 79440 86810 79450
rect 86940 79440 87060 79450
rect 87190 79440 87310 79450
rect 87440 79440 87560 79450
rect 87690 79440 87810 79450
rect 87940 79440 88060 79450
rect 88190 79440 88310 79450
rect 88440 79440 88560 79450
rect 88690 79440 88810 79450
rect 88940 79440 89060 79450
rect 89190 79440 89310 79450
rect 89440 79440 89560 79450
rect 89690 79440 89810 79450
rect 89940 79440 90060 79450
rect 90190 79440 90310 79450
rect 90440 79440 90560 79450
rect 90690 79440 90810 79450
rect 90940 79440 91060 79450
rect 91190 79440 91310 79450
rect 91440 79440 91560 79450
rect 91690 79440 91810 79450
rect 91940 79440 92000 79450
rect 81000 79310 81050 79440
rect 81200 79310 81300 79440
rect 81450 79310 81550 79440
rect 81700 79310 81800 79440
rect 81950 79310 82050 79440
rect 82200 79310 82300 79440
rect 82450 79310 82550 79440
rect 82700 79310 82800 79440
rect 82950 79310 83050 79440
rect 83200 79310 83300 79440
rect 83450 79310 83550 79440
rect 83700 79310 83800 79440
rect 83950 79310 84050 79440
rect 84200 79310 84300 79440
rect 84450 79310 84550 79440
rect 84700 79310 84800 79440
rect 84950 79310 85050 79440
rect 85200 79310 85300 79440
rect 85450 79310 85550 79440
rect 85700 79310 85800 79440
rect 85950 79310 86050 79440
rect 86200 79310 86300 79440
rect 86450 79310 86550 79440
rect 86700 79310 86800 79440
rect 86950 79310 87050 79440
rect 87200 79310 87300 79440
rect 87450 79310 87550 79440
rect 87700 79310 87800 79440
rect 87950 79310 88050 79440
rect 88200 79310 88300 79440
rect 88450 79310 88550 79440
rect 88700 79310 88800 79440
rect 88950 79310 89050 79440
rect 89200 79310 89300 79440
rect 89450 79310 89550 79440
rect 89700 79310 89800 79440
rect 89950 79310 90050 79440
rect 90200 79310 90300 79440
rect 90450 79310 90550 79440
rect 90700 79310 90800 79440
rect 90950 79310 91050 79440
rect 91200 79310 91300 79440
rect 91450 79310 91550 79440
rect 91700 79310 91800 79440
rect 91950 79310 92000 79440
rect 81000 79300 81060 79310
rect 81190 79300 81310 79310
rect 81440 79300 81560 79310
rect 81690 79300 81810 79310
rect 81940 79300 82060 79310
rect 82190 79300 82310 79310
rect 82440 79300 82560 79310
rect 82690 79300 82810 79310
rect 82940 79300 83060 79310
rect 83190 79300 83310 79310
rect 83440 79300 83560 79310
rect 83690 79300 83810 79310
rect 83940 79300 84060 79310
rect 84190 79300 84310 79310
rect 84440 79300 84560 79310
rect 84690 79300 84810 79310
rect 84940 79300 85060 79310
rect 85190 79300 85310 79310
rect 85440 79300 85560 79310
rect 85690 79300 85810 79310
rect 85940 79300 86060 79310
rect 86190 79300 86310 79310
rect 86440 79300 86560 79310
rect 86690 79300 86810 79310
rect 86940 79300 87060 79310
rect 87190 79300 87310 79310
rect 87440 79300 87560 79310
rect 87690 79300 87810 79310
rect 87940 79300 88060 79310
rect 88190 79300 88310 79310
rect 88440 79300 88560 79310
rect 88690 79300 88810 79310
rect 88940 79300 89060 79310
rect 89190 79300 89310 79310
rect 89440 79300 89560 79310
rect 89690 79300 89810 79310
rect 89940 79300 90060 79310
rect 90190 79300 90310 79310
rect 90440 79300 90560 79310
rect 90690 79300 90810 79310
rect 90940 79300 91060 79310
rect 91190 79300 91310 79310
rect 91440 79300 91560 79310
rect 91690 79300 91810 79310
rect 91940 79300 92000 79310
rect 81000 79200 92000 79300
rect 81000 79190 81060 79200
rect 81190 79190 81310 79200
rect 81440 79190 81560 79200
rect 81690 79190 81810 79200
rect 81940 79190 82060 79200
rect 82190 79190 82310 79200
rect 82440 79190 82560 79200
rect 82690 79190 82810 79200
rect 82940 79190 83060 79200
rect 83190 79190 83310 79200
rect 83440 79190 83560 79200
rect 83690 79190 83810 79200
rect 83940 79190 84060 79200
rect 84190 79190 84310 79200
rect 84440 79190 84560 79200
rect 84690 79190 84810 79200
rect 84940 79190 85060 79200
rect 85190 79190 85310 79200
rect 85440 79190 85560 79200
rect 85690 79190 85810 79200
rect 85940 79190 86060 79200
rect 86190 79190 86310 79200
rect 86440 79190 86560 79200
rect 86690 79190 86810 79200
rect 86940 79190 87060 79200
rect 87190 79190 87310 79200
rect 87440 79190 87560 79200
rect 87690 79190 87810 79200
rect 87940 79190 88060 79200
rect 88190 79190 88310 79200
rect 88440 79190 88560 79200
rect 88690 79190 88810 79200
rect 88940 79190 89060 79200
rect 89190 79190 89310 79200
rect 89440 79190 89560 79200
rect 89690 79190 89810 79200
rect 89940 79190 90060 79200
rect 90190 79190 90310 79200
rect 90440 79190 90560 79200
rect 90690 79190 90810 79200
rect 90940 79190 91060 79200
rect 91190 79190 91310 79200
rect 91440 79190 91560 79200
rect 91690 79190 91810 79200
rect 91940 79190 92000 79200
rect 81000 79060 81050 79190
rect 81200 79060 81300 79190
rect 81450 79060 81550 79190
rect 81700 79060 81800 79190
rect 81950 79060 82050 79190
rect 82200 79060 82300 79190
rect 82450 79060 82550 79190
rect 82700 79060 82800 79190
rect 82950 79060 83050 79190
rect 83200 79060 83300 79190
rect 83450 79060 83550 79190
rect 83700 79060 83800 79190
rect 83950 79060 84050 79190
rect 84200 79060 84300 79190
rect 84450 79060 84550 79190
rect 84700 79060 84800 79190
rect 84950 79060 85050 79190
rect 85200 79060 85300 79190
rect 85450 79060 85550 79190
rect 85700 79060 85800 79190
rect 85950 79060 86050 79190
rect 86200 79060 86300 79190
rect 86450 79060 86550 79190
rect 86700 79060 86800 79190
rect 86950 79060 87050 79190
rect 87200 79060 87300 79190
rect 87450 79060 87550 79190
rect 87700 79060 87800 79190
rect 87950 79060 88050 79190
rect 88200 79060 88300 79190
rect 88450 79060 88550 79190
rect 88700 79060 88800 79190
rect 88950 79060 89050 79190
rect 89200 79060 89300 79190
rect 89450 79060 89550 79190
rect 89700 79060 89800 79190
rect 89950 79060 90050 79190
rect 90200 79060 90300 79190
rect 90450 79060 90550 79190
rect 90700 79060 90800 79190
rect 90950 79060 91050 79190
rect 91200 79060 91300 79190
rect 91450 79060 91550 79190
rect 91700 79060 91800 79190
rect 91950 79060 92000 79190
rect 81000 79050 81060 79060
rect 81190 79050 81310 79060
rect 81440 79050 81560 79060
rect 81690 79050 81810 79060
rect 81940 79050 82060 79060
rect 82190 79050 82310 79060
rect 82440 79050 82560 79060
rect 82690 79050 82810 79060
rect 82940 79050 83060 79060
rect 83190 79050 83310 79060
rect 83440 79050 83560 79060
rect 83690 79050 83810 79060
rect 83940 79050 84060 79060
rect 84190 79050 84310 79060
rect 84440 79050 84560 79060
rect 84690 79050 84810 79060
rect 84940 79050 85060 79060
rect 85190 79050 85310 79060
rect 85440 79050 85560 79060
rect 85690 79050 85810 79060
rect 85940 79050 86060 79060
rect 86190 79050 86310 79060
rect 86440 79050 86560 79060
rect 86690 79050 86810 79060
rect 86940 79050 87060 79060
rect 87190 79050 87310 79060
rect 87440 79050 87560 79060
rect 87690 79050 87810 79060
rect 87940 79050 88060 79060
rect 88190 79050 88310 79060
rect 88440 79050 88560 79060
rect 88690 79050 88810 79060
rect 88940 79050 89060 79060
rect 89190 79050 89310 79060
rect 89440 79050 89560 79060
rect 89690 79050 89810 79060
rect 89940 79050 90060 79060
rect 90190 79050 90310 79060
rect 90440 79050 90560 79060
rect 90690 79050 90810 79060
rect 90940 79050 91060 79060
rect 91190 79050 91310 79060
rect 91440 79050 91560 79060
rect 91690 79050 91810 79060
rect 91940 79050 92000 79060
rect 81000 78950 92000 79050
rect 81000 78940 81060 78950
rect 81190 78940 81310 78950
rect 81440 78940 81560 78950
rect 81690 78940 81810 78950
rect 81940 78940 82060 78950
rect 82190 78940 82310 78950
rect 82440 78940 82560 78950
rect 82690 78940 82810 78950
rect 82940 78940 83060 78950
rect 83190 78940 83310 78950
rect 83440 78940 83560 78950
rect 83690 78940 83810 78950
rect 83940 78940 84060 78950
rect 84190 78940 84310 78950
rect 84440 78940 84560 78950
rect 84690 78940 84810 78950
rect 84940 78940 85060 78950
rect 85190 78940 85310 78950
rect 85440 78940 85560 78950
rect 85690 78940 85810 78950
rect 85940 78940 86060 78950
rect 86190 78940 86310 78950
rect 86440 78940 86560 78950
rect 86690 78940 86810 78950
rect 86940 78940 87060 78950
rect 87190 78940 87310 78950
rect 87440 78940 87560 78950
rect 87690 78940 87810 78950
rect 87940 78940 88060 78950
rect 88190 78940 88310 78950
rect 88440 78940 88560 78950
rect 88690 78940 88810 78950
rect 88940 78940 89060 78950
rect 89190 78940 89310 78950
rect 89440 78940 89560 78950
rect 89690 78940 89810 78950
rect 89940 78940 90060 78950
rect 90190 78940 90310 78950
rect 90440 78940 90560 78950
rect 90690 78940 90810 78950
rect 90940 78940 91060 78950
rect 91190 78940 91310 78950
rect 91440 78940 91560 78950
rect 91690 78940 91810 78950
rect 91940 78940 92000 78950
rect 81000 78810 81050 78940
rect 81200 78810 81300 78940
rect 81450 78810 81550 78940
rect 81700 78810 81800 78940
rect 81950 78810 82050 78940
rect 82200 78810 82300 78940
rect 82450 78810 82550 78940
rect 82700 78810 82800 78940
rect 82950 78810 83050 78940
rect 83200 78810 83300 78940
rect 83450 78810 83550 78940
rect 83700 78810 83800 78940
rect 83950 78810 84050 78940
rect 84200 78810 84300 78940
rect 84450 78810 84550 78940
rect 84700 78810 84800 78940
rect 84950 78810 85050 78940
rect 85200 78810 85300 78940
rect 85450 78810 85550 78940
rect 85700 78810 85800 78940
rect 85950 78810 86050 78940
rect 86200 78810 86300 78940
rect 86450 78810 86550 78940
rect 86700 78810 86800 78940
rect 86950 78810 87050 78940
rect 87200 78810 87300 78940
rect 87450 78810 87550 78940
rect 87700 78810 87800 78940
rect 87950 78810 88050 78940
rect 88200 78810 88300 78940
rect 88450 78810 88550 78940
rect 88700 78810 88800 78940
rect 88950 78810 89050 78940
rect 89200 78810 89300 78940
rect 89450 78810 89550 78940
rect 89700 78810 89800 78940
rect 89950 78810 90050 78940
rect 90200 78810 90300 78940
rect 90450 78810 90550 78940
rect 90700 78810 90800 78940
rect 90950 78810 91050 78940
rect 91200 78810 91300 78940
rect 91450 78810 91550 78940
rect 91700 78810 91800 78940
rect 91950 78810 92000 78940
rect 81000 78800 81060 78810
rect 81190 78800 81310 78810
rect 81440 78800 81560 78810
rect 81690 78800 81810 78810
rect 81940 78800 82060 78810
rect 82190 78800 82310 78810
rect 82440 78800 82560 78810
rect 82690 78800 82810 78810
rect 82940 78800 83060 78810
rect 83190 78800 83310 78810
rect 83440 78800 83560 78810
rect 83690 78800 83810 78810
rect 83940 78800 84060 78810
rect 84190 78800 84310 78810
rect 84440 78800 84560 78810
rect 84690 78800 84810 78810
rect 84940 78800 85060 78810
rect 85190 78800 85310 78810
rect 85440 78800 85560 78810
rect 85690 78800 85810 78810
rect 85940 78800 86060 78810
rect 86190 78800 86310 78810
rect 86440 78800 86560 78810
rect 86690 78800 86810 78810
rect 86940 78800 87060 78810
rect 87190 78800 87310 78810
rect 87440 78800 87560 78810
rect 87690 78800 87810 78810
rect 87940 78800 88060 78810
rect 88190 78800 88310 78810
rect 88440 78800 88560 78810
rect 88690 78800 88810 78810
rect 88940 78800 89060 78810
rect 89190 78800 89310 78810
rect 89440 78800 89560 78810
rect 89690 78800 89810 78810
rect 89940 78800 90060 78810
rect 90190 78800 90310 78810
rect 90440 78800 90560 78810
rect 90690 78800 90810 78810
rect 90940 78800 91060 78810
rect 91190 78800 91310 78810
rect 91440 78800 91560 78810
rect 91690 78800 91810 78810
rect 91940 78800 92000 78810
rect 81000 78700 92000 78800
rect 81000 78690 81060 78700
rect 81190 78690 81310 78700
rect 81440 78690 81560 78700
rect 81690 78690 81810 78700
rect 81940 78690 82060 78700
rect 82190 78690 82310 78700
rect 82440 78690 82560 78700
rect 82690 78690 82810 78700
rect 82940 78690 83060 78700
rect 83190 78690 83310 78700
rect 83440 78690 83560 78700
rect 83690 78690 83810 78700
rect 83940 78690 84060 78700
rect 84190 78690 84310 78700
rect 84440 78690 84560 78700
rect 84690 78690 84810 78700
rect 84940 78690 85060 78700
rect 85190 78690 85310 78700
rect 85440 78690 85560 78700
rect 85690 78690 85810 78700
rect 85940 78690 86060 78700
rect 86190 78690 86310 78700
rect 86440 78690 86560 78700
rect 86690 78690 86810 78700
rect 86940 78690 87060 78700
rect 87190 78690 87310 78700
rect 87440 78690 87560 78700
rect 87690 78690 87810 78700
rect 87940 78690 88060 78700
rect 88190 78690 88310 78700
rect 88440 78690 88560 78700
rect 88690 78690 88810 78700
rect 88940 78690 89060 78700
rect 89190 78690 89310 78700
rect 89440 78690 89560 78700
rect 89690 78690 89810 78700
rect 89940 78690 90060 78700
rect 90190 78690 90310 78700
rect 90440 78690 90560 78700
rect 90690 78690 90810 78700
rect 90940 78690 91060 78700
rect 91190 78690 91310 78700
rect 91440 78690 91560 78700
rect 91690 78690 91810 78700
rect 91940 78690 92000 78700
rect 81000 78560 81050 78690
rect 81200 78560 81300 78690
rect 81450 78560 81550 78690
rect 81700 78560 81800 78690
rect 81950 78560 82050 78690
rect 82200 78560 82300 78690
rect 82450 78560 82550 78690
rect 82700 78560 82800 78690
rect 82950 78560 83050 78690
rect 83200 78560 83300 78690
rect 83450 78560 83550 78690
rect 83700 78560 83800 78690
rect 83950 78560 84050 78690
rect 84200 78560 84300 78690
rect 84450 78560 84550 78690
rect 84700 78560 84800 78690
rect 84950 78560 85050 78690
rect 85200 78560 85300 78690
rect 85450 78560 85550 78690
rect 85700 78560 85800 78690
rect 85950 78560 86050 78690
rect 86200 78560 86300 78690
rect 86450 78560 86550 78690
rect 86700 78560 86800 78690
rect 86950 78560 87050 78690
rect 87200 78560 87300 78690
rect 87450 78560 87550 78690
rect 87700 78560 87800 78690
rect 87950 78560 88050 78690
rect 88200 78560 88300 78690
rect 88450 78560 88550 78690
rect 88700 78560 88800 78690
rect 88950 78560 89050 78690
rect 89200 78560 89300 78690
rect 89450 78560 89550 78690
rect 89700 78560 89800 78690
rect 89950 78560 90050 78690
rect 90200 78560 90300 78690
rect 90450 78560 90550 78690
rect 90700 78560 90800 78690
rect 90950 78560 91050 78690
rect 91200 78560 91300 78690
rect 91450 78560 91550 78690
rect 91700 78560 91800 78690
rect 91950 78560 92000 78690
rect 81000 78550 81060 78560
rect 81190 78550 81310 78560
rect 81440 78550 81560 78560
rect 81690 78550 81810 78560
rect 81940 78550 82060 78560
rect 82190 78550 82310 78560
rect 82440 78550 82560 78560
rect 82690 78550 82810 78560
rect 82940 78550 83060 78560
rect 83190 78550 83310 78560
rect 83440 78550 83560 78560
rect 83690 78550 83810 78560
rect 83940 78550 84060 78560
rect 84190 78550 84310 78560
rect 84440 78550 84560 78560
rect 84690 78550 84810 78560
rect 84940 78550 85060 78560
rect 85190 78550 85310 78560
rect 85440 78550 85560 78560
rect 85690 78550 85810 78560
rect 85940 78550 86060 78560
rect 86190 78550 86310 78560
rect 86440 78550 86560 78560
rect 86690 78550 86810 78560
rect 86940 78550 87060 78560
rect 87190 78550 87310 78560
rect 87440 78550 87560 78560
rect 87690 78550 87810 78560
rect 87940 78550 88060 78560
rect 88190 78550 88310 78560
rect 88440 78550 88560 78560
rect 88690 78550 88810 78560
rect 88940 78550 89060 78560
rect 89190 78550 89310 78560
rect 89440 78550 89560 78560
rect 89690 78550 89810 78560
rect 89940 78550 90060 78560
rect 90190 78550 90310 78560
rect 90440 78550 90560 78560
rect 90690 78550 90810 78560
rect 90940 78550 91060 78560
rect 91190 78550 91310 78560
rect 91440 78550 91560 78560
rect 91690 78550 91810 78560
rect 91940 78550 92000 78560
rect 81000 78450 92000 78550
rect 81000 78440 81060 78450
rect 81190 78440 81310 78450
rect 81440 78440 81560 78450
rect 81690 78440 81810 78450
rect 81940 78440 82060 78450
rect 82190 78440 82310 78450
rect 82440 78440 82560 78450
rect 82690 78440 82810 78450
rect 82940 78440 83060 78450
rect 83190 78440 83310 78450
rect 83440 78440 83560 78450
rect 83690 78440 83810 78450
rect 83940 78440 84060 78450
rect 84190 78440 84310 78450
rect 84440 78440 84560 78450
rect 84690 78440 84810 78450
rect 84940 78440 85060 78450
rect 85190 78440 85310 78450
rect 85440 78440 85560 78450
rect 85690 78440 85810 78450
rect 85940 78440 86060 78450
rect 86190 78440 86310 78450
rect 86440 78440 86560 78450
rect 86690 78440 86810 78450
rect 86940 78440 87060 78450
rect 87190 78440 87310 78450
rect 87440 78440 87560 78450
rect 87690 78440 87810 78450
rect 87940 78440 88060 78450
rect 88190 78440 88310 78450
rect 88440 78440 88560 78450
rect 88690 78440 88810 78450
rect 88940 78440 89060 78450
rect 89190 78440 89310 78450
rect 89440 78440 89560 78450
rect 89690 78440 89810 78450
rect 89940 78440 90060 78450
rect 90190 78440 90310 78450
rect 90440 78440 90560 78450
rect 90690 78440 90810 78450
rect 90940 78440 91060 78450
rect 91190 78440 91310 78450
rect 91440 78440 91560 78450
rect 91690 78440 91810 78450
rect 91940 78440 92000 78450
rect 81000 78310 81050 78440
rect 81200 78310 81300 78440
rect 81450 78310 81550 78440
rect 81700 78310 81800 78440
rect 81950 78310 82050 78440
rect 82200 78310 82300 78440
rect 82450 78310 82550 78440
rect 82700 78310 82800 78440
rect 82950 78310 83050 78440
rect 83200 78310 83300 78440
rect 83450 78310 83550 78440
rect 83700 78310 83800 78440
rect 83950 78310 84050 78440
rect 84200 78310 84300 78440
rect 84450 78310 84550 78440
rect 84700 78310 84800 78440
rect 84950 78310 85050 78440
rect 85200 78310 85300 78440
rect 85450 78310 85550 78440
rect 85700 78310 85800 78440
rect 85950 78310 86050 78440
rect 86200 78310 86300 78440
rect 86450 78310 86550 78440
rect 86700 78310 86800 78440
rect 86950 78310 87050 78440
rect 87200 78310 87300 78440
rect 87450 78310 87550 78440
rect 87700 78310 87800 78440
rect 87950 78310 88050 78440
rect 88200 78310 88300 78440
rect 88450 78310 88550 78440
rect 88700 78310 88800 78440
rect 88950 78310 89050 78440
rect 89200 78310 89300 78440
rect 89450 78310 89550 78440
rect 89700 78310 89800 78440
rect 89950 78310 90050 78440
rect 90200 78310 90300 78440
rect 90450 78310 90550 78440
rect 90700 78310 90800 78440
rect 90950 78310 91050 78440
rect 91200 78310 91300 78440
rect 91450 78310 91550 78440
rect 91700 78310 91800 78440
rect 91950 78310 92000 78440
rect 81000 78300 81060 78310
rect 81190 78300 81310 78310
rect 81440 78300 81560 78310
rect 81690 78300 81810 78310
rect 81940 78300 82060 78310
rect 82190 78300 82310 78310
rect 82440 78300 82560 78310
rect 82690 78300 82810 78310
rect 82940 78300 83060 78310
rect 83190 78300 83310 78310
rect 83440 78300 83560 78310
rect 83690 78300 83810 78310
rect 83940 78300 84060 78310
rect 84190 78300 84310 78310
rect 84440 78300 84560 78310
rect 84690 78300 84810 78310
rect 84940 78300 85060 78310
rect 85190 78300 85310 78310
rect 85440 78300 85560 78310
rect 85690 78300 85810 78310
rect 85940 78300 86060 78310
rect 86190 78300 86310 78310
rect 86440 78300 86560 78310
rect 86690 78300 86810 78310
rect 86940 78300 87060 78310
rect 87190 78300 87310 78310
rect 87440 78300 87560 78310
rect 87690 78300 87810 78310
rect 87940 78300 88060 78310
rect 88190 78300 88310 78310
rect 88440 78300 88560 78310
rect 88690 78300 88810 78310
rect 88940 78300 89060 78310
rect 89190 78300 89310 78310
rect 89440 78300 89560 78310
rect 89690 78300 89810 78310
rect 89940 78300 90060 78310
rect 90190 78300 90310 78310
rect 90440 78300 90560 78310
rect 90690 78300 90810 78310
rect 90940 78300 91060 78310
rect 91190 78300 91310 78310
rect 91440 78300 91560 78310
rect 91690 78300 91810 78310
rect 91940 78300 92000 78310
rect 81000 78200 92000 78300
rect 81000 78190 81060 78200
rect 81190 78190 81310 78200
rect 81440 78190 81560 78200
rect 81690 78190 81810 78200
rect 81940 78190 82060 78200
rect 82190 78190 82310 78200
rect 82440 78190 82560 78200
rect 82690 78190 82810 78200
rect 82940 78190 83060 78200
rect 83190 78190 83310 78200
rect 83440 78190 83560 78200
rect 83690 78190 83810 78200
rect 83940 78190 84060 78200
rect 84190 78190 84310 78200
rect 84440 78190 84560 78200
rect 84690 78190 84810 78200
rect 84940 78190 85060 78200
rect 85190 78190 85310 78200
rect 85440 78190 85560 78200
rect 85690 78190 85810 78200
rect 85940 78190 86060 78200
rect 86190 78190 86310 78200
rect 86440 78190 86560 78200
rect 86690 78190 86810 78200
rect 86940 78190 87060 78200
rect 87190 78190 87310 78200
rect 87440 78190 87560 78200
rect 87690 78190 87810 78200
rect 87940 78190 88060 78200
rect 88190 78190 88310 78200
rect 88440 78190 88560 78200
rect 88690 78190 88810 78200
rect 88940 78190 89060 78200
rect 89190 78190 89310 78200
rect 89440 78190 89560 78200
rect 89690 78190 89810 78200
rect 89940 78190 90060 78200
rect 90190 78190 90310 78200
rect 90440 78190 90560 78200
rect 90690 78190 90810 78200
rect 90940 78190 91060 78200
rect 91190 78190 91310 78200
rect 91440 78190 91560 78200
rect 91690 78190 91810 78200
rect 91940 78190 92000 78200
rect 81000 78060 81050 78190
rect 81200 78060 81300 78190
rect 81450 78060 81550 78190
rect 81700 78060 81800 78190
rect 81950 78060 82050 78190
rect 82200 78060 82300 78190
rect 82450 78060 82550 78190
rect 82700 78060 82800 78190
rect 82950 78060 83050 78190
rect 83200 78060 83300 78190
rect 83450 78060 83550 78190
rect 83700 78060 83800 78190
rect 83950 78060 84050 78190
rect 84200 78060 84300 78190
rect 84450 78060 84550 78190
rect 84700 78060 84800 78190
rect 84950 78060 85050 78190
rect 85200 78060 85300 78190
rect 85450 78060 85550 78190
rect 85700 78060 85800 78190
rect 85950 78060 86050 78190
rect 86200 78060 86300 78190
rect 86450 78060 86550 78190
rect 86700 78060 86800 78190
rect 86950 78060 87050 78190
rect 87200 78060 87300 78190
rect 87450 78060 87550 78190
rect 87700 78060 87800 78190
rect 87950 78060 88050 78190
rect 88200 78060 88300 78190
rect 88450 78060 88550 78190
rect 88700 78060 88800 78190
rect 88950 78060 89050 78190
rect 89200 78060 89300 78190
rect 89450 78060 89550 78190
rect 89700 78060 89800 78190
rect 89950 78060 90050 78190
rect 90200 78060 90300 78190
rect 90450 78060 90550 78190
rect 90700 78060 90800 78190
rect 90950 78060 91050 78190
rect 91200 78060 91300 78190
rect 91450 78060 91550 78190
rect 91700 78060 91800 78190
rect 91950 78060 92000 78190
rect 81000 78050 81060 78060
rect 81190 78050 81310 78060
rect 81440 78050 81560 78060
rect 81690 78050 81810 78060
rect 81940 78050 82060 78060
rect 82190 78050 82310 78060
rect 82440 78050 82560 78060
rect 82690 78050 82810 78060
rect 82940 78050 83060 78060
rect 83190 78050 83310 78060
rect 83440 78050 83560 78060
rect 83690 78050 83810 78060
rect 83940 78050 84060 78060
rect 84190 78050 84310 78060
rect 84440 78050 84560 78060
rect 84690 78050 84810 78060
rect 84940 78050 85060 78060
rect 85190 78050 85310 78060
rect 85440 78050 85560 78060
rect 85690 78050 85810 78060
rect 85940 78050 86060 78060
rect 86190 78050 86310 78060
rect 86440 78050 86560 78060
rect 86690 78050 86810 78060
rect 86940 78050 87060 78060
rect 87190 78050 87310 78060
rect 87440 78050 87560 78060
rect 87690 78050 87810 78060
rect 87940 78050 88060 78060
rect 88190 78050 88310 78060
rect 88440 78050 88560 78060
rect 88690 78050 88810 78060
rect 88940 78050 89060 78060
rect 89190 78050 89310 78060
rect 89440 78050 89560 78060
rect 89690 78050 89810 78060
rect 89940 78050 90060 78060
rect 90190 78050 90310 78060
rect 90440 78050 90560 78060
rect 90690 78050 90810 78060
rect 90940 78050 91060 78060
rect 91190 78050 91310 78060
rect 91440 78050 91560 78060
rect 91690 78050 91810 78060
rect 91940 78050 92000 78060
rect 81000 77950 92000 78050
rect 81000 77940 81060 77950
rect 81190 77940 81310 77950
rect 81440 77940 81560 77950
rect 81690 77940 81810 77950
rect 81940 77940 82060 77950
rect 82190 77940 82310 77950
rect 82440 77940 82560 77950
rect 82690 77940 82810 77950
rect 82940 77940 83060 77950
rect 83190 77940 83310 77950
rect 83440 77940 83560 77950
rect 83690 77940 83810 77950
rect 83940 77940 84060 77950
rect 84190 77940 84310 77950
rect 84440 77940 84560 77950
rect 84690 77940 84810 77950
rect 84940 77940 85060 77950
rect 85190 77940 85310 77950
rect 85440 77940 85560 77950
rect 85690 77940 85810 77950
rect 85940 77940 86060 77950
rect 86190 77940 86310 77950
rect 86440 77940 86560 77950
rect 86690 77940 86810 77950
rect 86940 77940 87060 77950
rect 87190 77940 87310 77950
rect 87440 77940 87560 77950
rect 87690 77940 87810 77950
rect 87940 77940 88060 77950
rect 88190 77940 88310 77950
rect 88440 77940 88560 77950
rect 88690 77940 88810 77950
rect 88940 77940 89060 77950
rect 89190 77940 89310 77950
rect 89440 77940 89560 77950
rect 89690 77940 89810 77950
rect 89940 77940 90060 77950
rect 90190 77940 90310 77950
rect 90440 77940 90560 77950
rect 90690 77940 90810 77950
rect 90940 77940 91060 77950
rect 91190 77940 91310 77950
rect 91440 77940 91560 77950
rect 91690 77940 91810 77950
rect 91940 77940 92000 77950
rect 81000 77810 81050 77940
rect 81200 77810 81300 77940
rect 81450 77810 81550 77940
rect 81700 77810 81800 77940
rect 81950 77810 82050 77940
rect 82200 77810 82300 77940
rect 82450 77810 82550 77940
rect 82700 77810 82800 77940
rect 82950 77810 83050 77940
rect 83200 77810 83300 77940
rect 83450 77810 83550 77940
rect 83700 77810 83800 77940
rect 83950 77810 84050 77940
rect 84200 77810 84300 77940
rect 84450 77810 84550 77940
rect 84700 77810 84800 77940
rect 84950 77810 85050 77940
rect 85200 77810 85300 77940
rect 85450 77810 85550 77940
rect 85700 77810 85800 77940
rect 85950 77810 86050 77940
rect 86200 77810 86300 77940
rect 86450 77810 86550 77940
rect 86700 77810 86800 77940
rect 86950 77810 87050 77940
rect 87200 77810 87300 77940
rect 87450 77810 87550 77940
rect 87700 77810 87800 77940
rect 87950 77810 88050 77940
rect 88200 77810 88300 77940
rect 88450 77810 88550 77940
rect 88700 77810 88800 77940
rect 88950 77810 89050 77940
rect 89200 77810 89300 77940
rect 89450 77810 89550 77940
rect 89700 77810 89800 77940
rect 89950 77810 90050 77940
rect 90200 77810 90300 77940
rect 90450 77810 90550 77940
rect 90700 77810 90800 77940
rect 90950 77810 91050 77940
rect 91200 77810 91300 77940
rect 91450 77810 91550 77940
rect 91700 77810 91800 77940
rect 91950 77810 92000 77940
rect 81000 77800 81060 77810
rect 81190 77800 81310 77810
rect 81440 77800 81560 77810
rect 81690 77800 81810 77810
rect 81940 77800 82060 77810
rect 82190 77800 82310 77810
rect 82440 77800 82560 77810
rect 82690 77800 82810 77810
rect 82940 77800 83060 77810
rect 83190 77800 83310 77810
rect 83440 77800 83560 77810
rect 83690 77800 83810 77810
rect 83940 77800 84060 77810
rect 84190 77800 84310 77810
rect 84440 77800 84560 77810
rect 84690 77800 84810 77810
rect 84940 77800 85060 77810
rect 85190 77800 85310 77810
rect 85440 77800 85560 77810
rect 85690 77800 85810 77810
rect 85940 77800 86060 77810
rect 86190 77800 86310 77810
rect 86440 77800 86560 77810
rect 86690 77800 86810 77810
rect 86940 77800 87060 77810
rect 87190 77800 87310 77810
rect 87440 77800 87560 77810
rect 87690 77800 87810 77810
rect 87940 77800 88060 77810
rect 88190 77800 88310 77810
rect 88440 77800 88560 77810
rect 88690 77800 88810 77810
rect 88940 77800 89060 77810
rect 89190 77800 89310 77810
rect 89440 77800 89560 77810
rect 89690 77800 89810 77810
rect 89940 77800 90060 77810
rect 90190 77800 90310 77810
rect 90440 77800 90560 77810
rect 90690 77800 90810 77810
rect 90940 77800 91060 77810
rect 91190 77800 91310 77810
rect 91440 77800 91560 77810
rect 91690 77800 91810 77810
rect 91940 77800 92000 77810
rect 81000 77700 92000 77800
rect 81000 77690 81060 77700
rect 81190 77690 81310 77700
rect 81440 77690 81560 77700
rect 81690 77690 81810 77700
rect 81940 77690 82060 77700
rect 82190 77690 82310 77700
rect 82440 77690 82560 77700
rect 82690 77690 82810 77700
rect 82940 77690 83060 77700
rect 83190 77690 83310 77700
rect 83440 77690 83560 77700
rect 83690 77690 83810 77700
rect 83940 77690 84060 77700
rect 84190 77690 84310 77700
rect 84440 77690 84560 77700
rect 84690 77690 84810 77700
rect 84940 77690 85060 77700
rect 85190 77690 85310 77700
rect 85440 77690 85560 77700
rect 85690 77690 85810 77700
rect 85940 77690 86060 77700
rect 86190 77690 86310 77700
rect 86440 77690 86560 77700
rect 86690 77690 86810 77700
rect 86940 77690 87060 77700
rect 87190 77690 87310 77700
rect 87440 77690 87560 77700
rect 87690 77690 87810 77700
rect 87940 77690 88060 77700
rect 88190 77690 88310 77700
rect 88440 77690 88560 77700
rect 88690 77690 88810 77700
rect 88940 77690 89060 77700
rect 89190 77690 89310 77700
rect 89440 77690 89560 77700
rect 89690 77690 89810 77700
rect 89940 77690 90060 77700
rect 90190 77690 90310 77700
rect 90440 77690 90560 77700
rect 90690 77690 90810 77700
rect 90940 77690 91060 77700
rect 91190 77690 91310 77700
rect 91440 77690 91560 77700
rect 91690 77690 91810 77700
rect 91940 77690 92000 77700
rect 81000 77560 81050 77690
rect 81200 77560 81300 77690
rect 81450 77560 81550 77690
rect 81700 77560 81800 77690
rect 81950 77560 82050 77690
rect 82200 77560 82300 77690
rect 82450 77560 82550 77690
rect 82700 77560 82800 77690
rect 82950 77560 83050 77690
rect 83200 77560 83300 77690
rect 83450 77560 83550 77690
rect 83700 77560 83800 77690
rect 83950 77560 84050 77690
rect 84200 77560 84300 77690
rect 84450 77560 84550 77690
rect 84700 77560 84800 77690
rect 84950 77560 85050 77690
rect 85200 77560 85300 77690
rect 85450 77560 85550 77690
rect 85700 77560 85800 77690
rect 85950 77560 86050 77690
rect 86200 77560 86300 77690
rect 86450 77560 86550 77690
rect 86700 77560 86800 77690
rect 86950 77560 87050 77690
rect 87200 77560 87300 77690
rect 87450 77560 87550 77690
rect 87700 77560 87800 77690
rect 87950 77560 88050 77690
rect 88200 77560 88300 77690
rect 88450 77560 88550 77690
rect 88700 77560 88800 77690
rect 88950 77560 89050 77690
rect 89200 77560 89300 77690
rect 89450 77560 89550 77690
rect 89700 77560 89800 77690
rect 89950 77560 90050 77690
rect 90200 77560 90300 77690
rect 90450 77560 90550 77690
rect 90700 77560 90800 77690
rect 90950 77560 91050 77690
rect 91200 77560 91300 77690
rect 91450 77560 91550 77690
rect 91700 77560 91800 77690
rect 91950 77560 92000 77690
rect 81000 77550 81060 77560
rect 81190 77550 81310 77560
rect 81440 77550 81560 77560
rect 81690 77550 81810 77560
rect 81940 77550 82060 77560
rect 82190 77550 82310 77560
rect 82440 77550 82560 77560
rect 82690 77550 82810 77560
rect 82940 77550 83060 77560
rect 83190 77550 83310 77560
rect 83440 77550 83560 77560
rect 83690 77550 83810 77560
rect 83940 77550 84060 77560
rect 84190 77550 84310 77560
rect 84440 77550 84560 77560
rect 84690 77550 84810 77560
rect 84940 77550 85060 77560
rect 85190 77550 85310 77560
rect 85440 77550 85560 77560
rect 85690 77550 85810 77560
rect 85940 77550 86060 77560
rect 86190 77550 86310 77560
rect 86440 77550 86560 77560
rect 86690 77550 86810 77560
rect 86940 77550 87060 77560
rect 87190 77550 87310 77560
rect 87440 77550 87560 77560
rect 87690 77550 87810 77560
rect 87940 77550 88060 77560
rect 88190 77550 88310 77560
rect 88440 77550 88560 77560
rect 88690 77550 88810 77560
rect 88940 77550 89060 77560
rect 89190 77550 89310 77560
rect 89440 77550 89560 77560
rect 89690 77550 89810 77560
rect 89940 77550 90060 77560
rect 90190 77550 90310 77560
rect 90440 77550 90560 77560
rect 90690 77550 90810 77560
rect 90940 77550 91060 77560
rect 91190 77550 91310 77560
rect 91440 77550 91560 77560
rect 91690 77550 91810 77560
rect 91940 77550 92000 77560
rect 81000 77450 92000 77550
rect 81000 77440 81060 77450
rect 81190 77440 81310 77450
rect 81440 77440 81560 77450
rect 81690 77440 81810 77450
rect 81940 77440 82060 77450
rect 82190 77440 82310 77450
rect 82440 77440 82560 77450
rect 82690 77440 82810 77450
rect 82940 77440 83060 77450
rect 83190 77440 83310 77450
rect 83440 77440 83560 77450
rect 83690 77440 83810 77450
rect 83940 77440 84060 77450
rect 84190 77440 84310 77450
rect 84440 77440 84560 77450
rect 84690 77440 84810 77450
rect 84940 77440 85060 77450
rect 85190 77440 85310 77450
rect 85440 77440 85560 77450
rect 85690 77440 85810 77450
rect 85940 77440 86060 77450
rect 86190 77440 86310 77450
rect 86440 77440 86560 77450
rect 86690 77440 86810 77450
rect 86940 77440 87060 77450
rect 87190 77440 87310 77450
rect 87440 77440 87560 77450
rect 87690 77440 87810 77450
rect 87940 77440 88060 77450
rect 88190 77440 88310 77450
rect 88440 77440 88560 77450
rect 88690 77440 88810 77450
rect 88940 77440 89060 77450
rect 89190 77440 89310 77450
rect 89440 77440 89560 77450
rect 89690 77440 89810 77450
rect 89940 77440 90060 77450
rect 90190 77440 90310 77450
rect 90440 77440 90560 77450
rect 90690 77440 90810 77450
rect 90940 77440 91060 77450
rect 91190 77440 91310 77450
rect 91440 77440 91560 77450
rect 91690 77440 91810 77450
rect 91940 77440 92000 77450
rect 81000 77310 81050 77440
rect 81200 77310 81300 77440
rect 81450 77310 81550 77440
rect 81700 77310 81800 77440
rect 81950 77310 82050 77440
rect 82200 77310 82300 77440
rect 82450 77310 82550 77440
rect 82700 77310 82800 77440
rect 82950 77310 83050 77440
rect 83200 77310 83300 77440
rect 83450 77310 83550 77440
rect 83700 77310 83800 77440
rect 83950 77310 84050 77440
rect 84200 77310 84300 77440
rect 84450 77310 84550 77440
rect 84700 77310 84800 77440
rect 84950 77310 85050 77440
rect 85200 77310 85300 77440
rect 85450 77310 85550 77440
rect 85700 77310 85800 77440
rect 85950 77310 86050 77440
rect 86200 77310 86300 77440
rect 86450 77310 86550 77440
rect 86700 77310 86800 77440
rect 86950 77310 87050 77440
rect 87200 77310 87300 77440
rect 87450 77310 87550 77440
rect 87700 77310 87800 77440
rect 87950 77310 88050 77440
rect 88200 77310 88300 77440
rect 88450 77310 88550 77440
rect 88700 77310 88800 77440
rect 88950 77310 89050 77440
rect 89200 77310 89300 77440
rect 89450 77310 89550 77440
rect 89700 77310 89800 77440
rect 89950 77310 90050 77440
rect 90200 77310 90300 77440
rect 90450 77310 90550 77440
rect 90700 77310 90800 77440
rect 90950 77310 91050 77440
rect 91200 77310 91300 77440
rect 91450 77310 91550 77440
rect 91700 77310 91800 77440
rect 91950 77310 92000 77440
rect 81000 77300 81060 77310
rect 81190 77300 81310 77310
rect 81440 77300 81560 77310
rect 81690 77300 81810 77310
rect 81940 77300 82060 77310
rect 82190 77300 82310 77310
rect 82440 77300 82560 77310
rect 82690 77300 82810 77310
rect 82940 77300 83060 77310
rect 83190 77300 83310 77310
rect 83440 77300 83560 77310
rect 83690 77300 83810 77310
rect 83940 77300 84060 77310
rect 84190 77300 84310 77310
rect 84440 77300 84560 77310
rect 84690 77300 84810 77310
rect 84940 77300 85060 77310
rect 85190 77300 85310 77310
rect 85440 77300 85560 77310
rect 85690 77300 85810 77310
rect 85940 77300 86060 77310
rect 86190 77300 86310 77310
rect 86440 77300 86560 77310
rect 86690 77300 86810 77310
rect 86940 77300 87060 77310
rect 87190 77300 87310 77310
rect 87440 77300 87560 77310
rect 87690 77300 87810 77310
rect 87940 77300 88060 77310
rect 88190 77300 88310 77310
rect 88440 77300 88560 77310
rect 88690 77300 88810 77310
rect 88940 77300 89060 77310
rect 89190 77300 89310 77310
rect 89440 77300 89560 77310
rect 89690 77300 89810 77310
rect 89940 77300 90060 77310
rect 90190 77300 90310 77310
rect 90440 77300 90560 77310
rect 90690 77300 90810 77310
rect 90940 77300 91060 77310
rect 91190 77300 91310 77310
rect 91440 77300 91560 77310
rect 91690 77300 91810 77310
rect 91940 77300 92000 77310
rect 81000 77200 92000 77300
rect 81000 77190 81060 77200
rect 81190 77190 81310 77200
rect 81440 77190 81560 77200
rect 81690 77190 81810 77200
rect 81940 77190 82060 77200
rect 82190 77190 82310 77200
rect 82440 77190 82560 77200
rect 82690 77190 82810 77200
rect 82940 77190 83060 77200
rect 83190 77190 83310 77200
rect 83440 77190 83560 77200
rect 83690 77190 83810 77200
rect 83940 77190 84060 77200
rect 84190 77190 84310 77200
rect 84440 77190 84560 77200
rect 84690 77190 84810 77200
rect 84940 77190 85060 77200
rect 85190 77190 85310 77200
rect 85440 77190 85560 77200
rect 85690 77190 85810 77200
rect 85940 77190 86060 77200
rect 86190 77190 86310 77200
rect 86440 77190 86560 77200
rect 86690 77190 86810 77200
rect 86940 77190 87060 77200
rect 87190 77190 87310 77200
rect 87440 77190 87560 77200
rect 87690 77190 87810 77200
rect 87940 77190 88060 77200
rect 88190 77190 88310 77200
rect 88440 77190 88560 77200
rect 88690 77190 88810 77200
rect 88940 77190 89060 77200
rect 89190 77190 89310 77200
rect 89440 77190 89560 77200
rect 89690 77190 89810 77200
rect 89940 77190 90060 77200
rect 90190 77190 90310 77200
rect 90440 77190 90560 77200
rect 90690 77190 90810 77200
rect 90940 77190 91060 77200
rect 91190 77190 91310 77200
rect 91440 77190 91560 77200
rect 91690 77190 91810 77200
rect 91940 77190 92000 77200
rect 81000 77060 81050 77190
rect 81200 77060 81300 77190
rect 81450 77060 81550 77190
rect 81700 77060 81800 77190
rect 81950 77060 82050 77190
rect 82200 77060 82300 77190
rect 82450 77060 82550 77190
rect 82700 77060 82800 77190
rect 82950 77060 83050 77190
rect 83200 77060 83300 77190
rect 83450 77060 83550 77190
rect 83700 77060 83800 77190
rect 83950 77060 84050 77190
rect 84200 77060 84300 77190
rect 84450 77060 84550 77190
rect 84700 77060 84800 77190
rect 84950 77060 85050 77190
rect 85200 77060 85300 77190
rect 85450 77060 85550 77190
rect 85700 77060 85800 77190
rect 85950 77060 86050 77190
rect 86200 77060 86300 77190
rect 86450 77060 86550 77190
rect 86700 77060 86800 77190
rect 86950 77060 87050 77190
rect 87200 77060 87300 77190
rect 87450 77060 87550 77190
rect 87700 77060 87800 77190
rect 87950 77060 88050 77190
rect 88200 77060 88300 77190
rect 88450 77060 88550 77190
rect 88700 77060 88800 77190
rect 88950 77060 89050 77190
rect 89200 77060 89300 77190
rect 89450 77060 89550 77190
rect 89700 77060 89800 77190
rect 89950 77060 90050 77190
rect 90200 77060 90300 77190
rect 90450 77060 90550 77190
rect 90700 77060 90800 77190
rect 90950 77060 91050 77190
rect 91200 77060 91300 77190
rect 91450 77060 91550 77190
rect 91700 77060 91800 77190
rect 91950 77060 92000 77190
rect 81000 77050 81060 77060
rect 81190 77050 81310 77060
rect 81440 77050 81560 77060
rect 81690 77050 81810 77060
rect 81940 77050 82060 77060
rect 82190 77050 82310 77060
rect 82440 77050 82560 77060
rect 82690 77050 82810 77060
rect 82940 77050 83060 77060
rect 83190 77050 83310 77060
rect 83440 77050 83560 77060
rect 83690 77050 83810 77060
rect 83940 77050 84060 77060
rect 84190 77050 84310 77060
rect 84440 77050 84560 77060
rect 84690 77050 84810 77060
rect 84940 77050 85060 77060
rect 85190 77050 85310 77060
rect 85440 77050 85560 77060
rect 85690 77050 85810 77060
rect 85940 77050 86060 77060
rect 86190 77050 86310 77060
rect 86440 77050 86560 77060
rect 86690 77050 86810 77060
rect 86940 77050 87060 77060
rect 87190 77050 87310 77060
rect 87440 77050 87560 77060
rect 87690 77050 87810 77060
rect 87940 77050 88060 77060
rect 88190 77050 88310 77060
rect 88440 77050 88560 77060
rect 88690 77050 88810 77060
rect 88940 77050 89060 77060
rect 89190 77050 89310 77060
rect 89440 77050 89560 77060
rect 89690 77050 89810 77060
rect 89940 77050 90060 77060
rect 90190 77050 90310 77060
rect 90440 77050 90560 77060
rect 90690 77050 90810 77060
rect 90940 77050 91060 77060
rect 91190 77050 91310 77060
rect 91440 77050 91560 77060
rect 91690 77050 91810 77060
rect 91940 77050 92000 77060
rect 81000 77000 92000 77050
rect 107000 80950 116000 81000
rect 107000 80940 107060 80950
rect 107190 80940 107310 80950
rect 107440 80940 107560 80950
rect 107690 80940 107810 80950
rect 107940 80940 108060 80950
rect 108190 80940 108310 80950
rect 108440 80940 108560 80950
rect 108690 80940 108810 80950
rect 108940 80940 109060 80950
rect 109190 80940 109310 80950
rect 109440 80940 109560 80950
rect 109690 80940 109810 80950
rect 109940 80940 110060 80950
rect 110190 80940 110310 80950
rect 110440 80940 110560 80950
rect 110690 80940 110810 80950
rect 110940 80940 111060 80950
rect 111190 80940 111310 80950
rect 111440 80940 111560 80950
rect 111690 80940 111810 80950
rect 111940 80940 112060 80950
rect 112190 80940 112310 80950
rect 112440 80940 112560 80950
rect 112690 80940 112810 80950
rect 112940 80940 113060 80950
rect 113190 80940 113310 80950
rect 113440 80940 113560 80950
rect 113690 80940 113810 80950
rect 113940 80940 114060 80950
rect 114190 80940 114310 80950
rect 114440 80940 114560 80950
rect 114690 80940 114810 80950
rect 114940 80940 115060 80950
rect 115190 80940 115310 80950
rect 115440 80940 115560 80950
rect 115690 80940 115810 80950
rect 115940 80940 116000 80950
rect 107000 80810 107050 80940
rect 107200 80810 107300 80940
rect 107450 80810 107550 80940
rect 107700 80810 107800 80940
rect 107950 80810 108050 80940
rect 108200 80810 108300 80940
rect 108450 80810 108550 80940
rect 108700 80810 108800 80940
rect 108950 80810 109050 80940
rect 109200 80810 109300 80940
rect 109450 80810 109550 80940
rect 109700 80810 109800 80940
rect 109950 80810 110050 80940
rect 110200 80810 110300 80940
rect 110450 80810 110550 80940
rect 110700 80810 110800 80940
rect 110950 80810 111050 80940
rect 111200 80810 111300 80940
rect 111450 80810 111550 80940
rect 111700 80810 111800 80940
rect 111950 80810 112050 80940
rect 112200 80810 112300 80940
rect 112450 80810 112550 80940
rect 112700 80810 112800 80940
rect 112950 80810 113050 80940
rect 113200 80810 113300 80940
rect 113450 80810 113550 80940
rect 113700 80810 113800 80940
rect 113950 80810 114050 80940
rect 114200 80810 114300 80940
rect 114450 80810 114550 80940
rect 114700 80810 114800 80940
rect 114950 80810 115050 80940
rect 115200 80810 115300 80940
rect 115450 80810 115550 80940
rect 115700 80810 115800 80940
rect 115950 80810 116000 80940
rect 107000 80800 107060 80810
rect 107190 80800 107310 80810
rect 107440 80800 107560 80810
rect 107690 80800 107810 80810
rect 107940 80800 108060 80810
rect 108190 80800 108310 80810
rect 108440 80800 108560 80810
rect 108690 80800 108810 80810
rect 108940 80800 109060 80810
rect 109190 80800 109310 80810
rect 109440 80800 109560 80810
rect 109690 80800 109810 80810
rect 109940 80800 110060 80810
rect 110190 80800 110310 80810
rect 110440 80800 110560 80810
rect 110690 80800 110810 80810
rect 110940 80800 111060 80810
rect 111190 80800 111310 80810
rect 111440 80800 111560 80810
rect 111690 80800 111810 80810
rect 111940 80800 112060 80810
rect 112190 80800 112310 80810
rect 112440 80800 112560 80810
rect 112690 80800 112810 80810
rect 112940 80800 113060 80810
rect 113190 80800 113310 80810
rect 113440 80800 113560 80810
rect 113690 80800 113810 80810
rect 113940 80800 114060 80810
rect 114190 80800 114310 80810
rect 114440 80800 114560 80810
rect 114690 80800 114810 80810
rect 114940 80800 115060 80810
rect 115190 80800 115310 80810
rect 115440 80800 115560 80810
rect 115690 80800 115810 80810
rect 115940 80800 116000 80810
rect 107000 80700 116000 80800
rect 107000 80690 107060 80700
rect 107190 80690 107310 80700
rect 107440 80690 107560 80700
rect 107690 80690 107810 80700
rect 107940 80690 108060 80700
rect 108190 80690 108310 80700
rect 108440 80690 108560 80700
rect 108690 80690 108810 80700
rect 108940 80690 109060 80700
rect 109190 80690 109310 80700
rect 109440 80690 109560 80700
rect 109690 80690 109810 80700
rect 109940 80690 110060 80700
rect 110190 80690 110310 80700
rect 110440 80690 110560 80700
rect 110690 80690 110810 80700
rect 110940 80690 111060 80700
rect 111190 80690 111310 80700
rect 111440 80690 111560 80700
rect 111690 80690 111810 80700
rect 111940 80690 112060 80700
rect 112190 80690 112310 80700
rect 112440 80690 112560 80700
rect 112690 80690 112810 80700
rect 112940 80690 113060 80700
rect 113190 80690 113310 80700
rect 113440 80690 113560 80700
rect 113690 80690 113810 80700
rect 113940 80690 114060 80700
rect 114190 80690 114310 80700
rect 114440 80690 114560 80700
rect 114690 80690 114810 80700
rect 114940 80690 115060 80700
rect 115190 80690 115310 80700
rect 115440 80690 115560 80700
rect 115690 80690 115810 80700
rect 115940 80690 116000 80700
rect 107000 80560 107050 80690
rect 107200 80560 107300 80690
rect 107450 80560 107550 80690
rect 107700 80560 107800 80690
rect 107950 80560 108050 80690
rect 108200 80560 108300 80690
rect 108450 80560 108550 80690
rect 108700 80560 108800 80690
rect 108950 80560 109050 80690
rect 109200 80560 109300 80690
rect 109450 80560 109550 80690
rect 109700 80560 109800 80690
rect 109950 80560 110050 80690
rect 110200 80560 110300 80690
rect 110450 80560 110550 80690
rect 110700 80560 110800 80690
rect 110950 80560 111050 80690
rect 111200 80560 111300 80690
rect 111450 80560 111550 80690
rect 111700 80560 111800 80690
rect 111950 80560 112050 80690
rect 112200 80560 112300 80690
rect 112450 80560 112550 80690
rect 112700 80560 112800 80690
rect 112950 80560 113050 80690
rect 113200 80560 113300 80690
rect 113450 80560 113550 80690
rect 113700 80560 113800 80690
rect 113950 80560 114050 80690
rect 114200 80560 114300 80690
rect 114450 80560 114550 80690
rect 114700 80560 114800 80690
rect 114950 80560 115050 80690
rect 115200 80560 115300 80690
rect 115450 80560 115550 80690
rect 115700 80560 115800 80690
rect 115950 80560 116000 80690
rect 107000 80550 107060 80560
rect 107190 80550 107310 80560
rect 107440 80550 107560 80560
rect 107690 80550 107810 80560
rect 107940 80550 108060 80560
rect 108190 80550 108310 80560
rect 108440 80550 108560 80560
rect 108690 80550 108810 80560
rect 108940 80550 109060 80560
rect 109190 80550 109310 80560
rect 109440 80550 109560 80560
rect 109690 80550 109810 80560
rect 109940 80550 110060 80560
rect 110190 80550 110310 80560
rect 110440 80550 110560 80560
rect 110690 80550 110810 80560
rect 110940 80550 111060 80560
rect 111190 80550 111310 80560
rect 111440 80550 111560 80560
rect 111690 80550 111810 80560
rect 111940 80550 112060 80560
rect 112190 80550 112310 80560
rect 112440 80550 112560 80560
rect 112690 80550 112810 80560
rect 112940 80550 113060 80560
rect 113190 80550 113310 80560
rect 113440 80550 113560 80560
rect 113690 80550 113810 80560
rect 113940 80550 114060 80560
rect 114190 80550 114310 80560
rect 114440 80550 114560 80560
rect 114690 80550 114810 80560
rect 114940 80550 115060 80560
rect 115190 80550 115310 80560
rect 115440 80550 115560 80560
rect 115690 80550 115810 80560
rect 115940 80550 116000 80560
rect 107000 80450 116000 80550
rect 107000 80440 107060 80450
rect 107190 80440 107310 80450
rect 107440 80440 107560 80450
rect 107690 80440 107810 80450
rect 107940 80440 108060 80450
rect 108190 80440 108310 80450
rect 108440 80440 108560 80450
rect 108690 80440 108810 80450
rect 108940 80440 109060 80450
rect 109190 80440 109310 80450
rect 109440 80440 109560 80450
rect 109690 80440 109810 80450
rect 109940 80440 110060 80450
rect 110190 80440 110310 80450
rect 110440 80440 110560 80450
rect 110690 80440 110810 80450
rect 110940 80440 111060 80450
rect 111190 80440 111310 80450
rect 111440 80440 111560 80450
rect 111690 80440 111810 80450
rect 111940 80440 112060 80450
rect 112190 80440 112310 80450
rect 112440 80440 112560 80450
rect 112690 80440 112810 80450
rect 112940 80440 113060 80450
rect 113190 80440 113310 80450
rect 113440 80440 113560 80450
rect 113690 80440 113810 80450
rect 113940 80440 114060 80450
rect 114190 80440 114310 80450
rect 114440 80440 114560 80450
rect 114690 80440 114810 80450
rect 114940 80440 115060 80450
rect 115190 80440 115310 80450
rect 115440 80440 115560 80450
rect 115690 80440 115810 80450
rect 115940 80440 116000 80450
rect 107000 80310 107050 80440
rect 107200 80310 107300 80440
rect 107450 80310 107550 80440
rect 107700 80310 107800 80440
rect 107950 80310 108050 80440
rect 108200 80310 108300 80440
rect 108450 80310 108550 80440
rect 108700 80310 108800 80440
rect 108950 80310 109050 80440
rect 109200 80310 109300 80440
rect 109450 80310 109550 80440
rect 109700 80310 109800 80440
rect 109950 80310 110050 80440
rect 110200 80310 110300 80440
rect 110450 80310 110550 80440
rect 110700 80310 110800 80440
rect 110950 80310 111050 80440
rect 111200 80310 111300 80440
rect 111450 80310 111550 80440
rect 111700 80310 111800 80440
rect 111950 80310 112050 80440
rect 112200 80310 112300 80440
rect 112450 80310 112550 80440
rect 112700 80310 112800 80440
rect 112950 80310 113050 80440
rect 113200 80310 113300 80440
rect 113450 80310 113550 80440
rect 113700 80310 113800 80440
rect 113950 80310 114050 80440
rect 114200 80310 114300 80440
rect 114450 80310 114550 80440
rect 114700 80310 114800 80440
rect 114950 80310 115050 80440
rect 115200 80310 115300 80440
rect 115450 80310 115550 80440
rect 115700 80310 115800 80440
rect 115950 80310 116000 80440
rect 107000 80300 107060 80310
rect 107190 80300 107310 80310
rect 107440 80300 107560 80310
rect 107690 80300 107810 80310
rect 107940 80300 108060 80310
rect 108190 80300 108310 80310
rect 108440 80300 108560 80310
rect 108690 80300 108810 80310
rect 108940 80300 109060 80310
rect 109190 80300 109310 80310
rect 109440 80300 109560 80310
rect 109690 80300 109810 80310
rect 109940 80300 110060 80310
rect 110190 80300 110310 80310
rect 110440 80300 110560 80310
rect 110690 80300 110810 80310
rect 110940 80300 111060 80310
rect 111190 80300 111310 80310
rect 111440 80300 111560 80310
rect 111690 80300 111810 80310
rect 111940 80300 112060 80310
rect 112190 80300 112310 80310
rect 112440 80300 112560 80310
rect 112690 80300 112810 80310
rect 112940 80300 113060 80310
rect 113190 80300 113310 80310
rect 113440 80300 113560 80310
rect 113690 80300 113810 80310
rect 113940 80300 114060 80310
rect 114190 80300 114310 80310
rect 114440 80300 114560 80310
rect 114690 80300 114810 80310
rect 114940 80300 115060 80310
rect 115190 80300 115310 80310
rect 115440 80300 115560 80310
rect 115690 80300 115810 80310
rect 115940 80300 116000 80310
rect 107000 80200 116000 80300
rect 107000 80190 107060 80200
rect 107190 80190 107310 80200
rect 107440 80190 107560 80200
rect 107690 80190 107810 80200
rect 107940 80190 108060 80200
rect 108190 80190 108310 80200
rect 108440 80190 108560 80200
rect 108690 80190 108810 80200
rect 108940 80190 109060 80200
rect 109190 80190 109310 80200
rect 109440 80190 109560 80200
rect 109690 80190 109810 80200
rect 109940 80190 110060 80200
rect 110190 80190 110310 80200
rect 110440 80190 110560 80200
rect 110690 80190 110810 80200
rect 110940 80190 111060 80200
rect 111190 80190 111310 80200
rect 111440 80190 111560 80200
rect 111690 80190 111810 80200
rect 111940 80190 112060 80200
rect 112190 80190 112310 80200
rect 112440 80190 112560 80200
rect 112690 80190 112810 80200
rect 112940 80190 113060 80200
rect 113190 80190 113310 80200
rect 113440 80190 113560 80200
rect 113690 80190 113810 80200
rect 113940 80190 114060 80200
rect 114190 80190 114310 80200
rect 114440 80190 114560 80200
rect 114690 80190 114810 80200
rect 114940 80190 115060 80200
rect 115190 80190 115310 80200
rect 115440 80190 115560 80200
rect 115690 80190 115810 80200
rect 115940 80190 116000 80200
rect 107000 80060 107050 80190
rect 107200 80060 107300 80190
rect 107450 80060 107550 80190
rect 107700 80060 107800 80190
rect 107950 80060 108050 80190
rect 108200 80060 108300 80190
rect 108450 80060 108550 80190
rect 108700 80060 108800 80190
rect 108950 80060 109050 80190
rect 109200 80060 109300 80190
rect 109450 80060 109550 80190
rect 109700 80060 109800 80190
rect 109950 80060 110050 80190
rect 110200 80060 110300 80190
rect 110450 80060 110550 80190
rect 110700 80060 110800 80190
rect 110950 80060 111050 80190
rect 111200 80060 111300 80190
rect 111450 80060 111550 80190
rect 111700 80060 111800 80190
rect 111950 80060 112050 80190
rect 112200 80060 112300 80190
rect 112450 80060 112550 80190
rect 112700 80060 112800 80190
rect 112950 80060 113050 80190
rect 113200 80060 113300 80190
rect 113450 80060 113550 80190
rect 113700 80060 113800 80190
rect 113950 80060 114050 80190
rect 114200 80060 114300 80190
rect 114450 80060 114550 80190
rect 114700 80060 114800 80190
rect 114950 80060 115050 80190
rect 115200 80060 115300 80190
rect 115450 80060 115550 80190
rect 115700 80060 115800 80190
rect 115950 80060 116000 80190
rect 107000 80050 107060 80060
rect 107190 80050 107310 80060
rect 107440 80050 107560 80060
rect 107690 80050 107810 80060
rect 107940 80050 108060 80060
rect 108190 80050 108310 80060
rect 108440 80050 108560 80060
rect 108690 80050 108810 80060
rect 108940 80050 109060 80060
rect 109190 80050 109310 80060
rect 109440 80050 109560 80060
rect 109690 80050 109810 80060
rect 109940 80050 110060 80060
rect 110190 80050 110310 80060
rect 110440 80050 110560 80060
rect 110690 80050 110810 80060
rect 110940 80050 111060 80060
rect 111190 80050 111310 80060
rect 111440 80050 111560 80060
rect 111690 80050 111810 80060
rect 111940 80050 112060 80060
rect 112190 80050 112310 80060
rect 112440 80050 112560 80060
rect 112690 80050 112810 80060
rect 112940 80050 113060 80060
rect 113190 80050 113310 80060
rect 113440 80050 113560 80060
rect 113690 80050 113810 80060
rect 113940 80050 114060 80060
rect 114190 80050 114310 80060
rect 114440 80050 114560 80060
rect 114690 80050 114810 80060
rect 114940 80050 115060 80060
rect 115190 80050 115310 80060
rect 115440 80050 115560 80060
rect 115690 80050 115810 80060
rect 115940 80050 116000 80060
rect 107000 79950 116000 80050
rect 107000 79940 107060 79950
rect 107190 79940 107310 79950
rect 107440 79940 107560 79950
rect 107690 79940 107810 79950
rect 107940 79940 108060 79950
rect 108190 79940 108310 79950
rect 108440 79940 108560 79950
rect 108690 79940 108810 79950
rect 108940 79940 109060 79950
rect 109190 79940 109310 79950
rect 109440 79940 109560 79950
rect 109690 79940 109810 79950
rect 109940 79940 110060 79950
rect 110190 79940 110310 79950
rect 110440 79940 110560 79950
rect 110690 79940 110810 79950
rect 110940 79940 111060 79950
rect 111190 79940 111310 79950
rect 111440 79940 111560 79950
rect 111690 79940 111810 79950
rect 111940 79940 112060 79950
rect 112190 79940 112310 79950
rect 112440 79940 112560 79950
rect 112690 79940 112810 79950
rect 112940 79940 113060 79950
rect 113190 79940 113310 79950
rect 113440 79940 113560 79950
rect 113690 79940 113810 79950
rect 113940 79940 114060 79950
rect 114190 79940 114310 79950
rect 114440 79940 114560 79950
rect 114690 79940 114810 79950
rect 114940 79940 115060 79950
rect 115190 79940 115310 79950
rect 115440 79940 115560 79950
rect 115690 79940 115810 79950
rect 115940 79940 116000 79950
rect 107000 79810 107050 79940
rect 107200 79810 107300 79940
rect 107450 79810 107550 79940
rect 107700 79810 107800 79940
rect 107950 79810 108050 79940
rect 108200 79810 108300 79940
rect 108450 79810 108550 79940
rect 108700 79810 108800 79940
rect 108950 79810 109050 79940
rect 109200 79810 109300 79940
rect 109450 79810 109550 79940
rect 109700 79810 109800 79940
rect 109950 79810 110050 79940
rect 110200 79810 110300 79940
rect 110450 79810 110550 79940
rect 110700 79810 110800 79940
rect 110950 79810 111050 79940
rect 111200 79810 111300 79940
rect 111450 79810 111550 79940
rect 111700 79810 111800 79940
rect 111950 79810 112050 79940
rect 112200 79810 112300 79940
rect 112450 79810 112550 79940
rect 112700 79810 112800 79940
rect 112950 79810 113050 79940
rect 113200 79810 113300 79940
rect 113450 79810 113550 79940
rect 113700 79810 113800 79940
rect 113950 79810 114050 79940
rect 114200 79810 114300 79940
rect 114450 79810 114550 79940
rect 114700 79810 114800 79940
rect 114950 79810 115050 79940
rect 115200 79810 115300 79940
rect 115450 79810 115550 79940
rect 115700 79810 115800 79940
rect 115950 79810 116000 79940
rect 107000 79800 107060 79810
rect 107190 79800 107310 79810
rect 107440 79800 107560 79810
rect 107690 79800 107810 79810
rect 107940 79800 108060 79810
rect 108190 79800 108310 79810
rect 108440 79800 108560 79810
rect 108690 79800 108810 79810
rect 108940 79800 109060 79810
rect 109190 79800 109310 79810
rect 109440 79800 109560 79810
rect 109690 79800 109810 79810
rect 109940 79800 110060 79810
rect 110190 79800 110310 79810
rect 110440 79800 110560 79810
rect 110690 79800 110810 79810
rect 110940 79800 111060 79810
rect 111190 79800 111310 79810
rect 111440 79800 111560 79810
rect 111690 79800 111810 79810
rect 111940 79800 112060 79810
rect 112190 79800 112310 79810
rect 112440 79800 112560 79810
rect 112690 79800 112810 79810
rect 112940 79800 113060 79810
rect 113190 79800 113310 79810
rect 113440 79800 113560 79810
rect 113690 79800 113810 79810
rect 113940 79800 114060 79810
rect 114190 79800 114310 79810
rect 114440 79800 114560 79810
rect 114690 79800 114810 79810
rect 114940 79800 115060 79810
rect 115190 79800 115310 79810
rect 115440 79800 115560 79810
rect 115690 79800 115810 79810
rect 115940 79800 116000 79810
rect 107000 79700 116000 79800
rect 107000 79690 107060 79700
rect 107190 79690 107310 79700
rect 107440 79690 107560 79700
rect 107690 79690 107810 79700
rect 107940 79690 108060 79700
rect 108190 79690 108310 79700
rect 108440 79690 108560 79700
rect 108690 79690 108810 79700
rect 108940 79690 109060 79700
rect 109190 79690 109310 79700
rect 109440 79690 109560 79700
rect 109690 79690 109810 79700
rect 109940 79690 110060 79700
rect 110190 79690 110310 79700
rect 110440 79690 110560 79700
rect 110690 79690 110810 79700
rect 110940 79690 111060 79700
rect 111190 79690 111310 79700
rect 111440 79690 111560 79700
rect 111690 79690 111810 79700
rect 111940 79690 112060 79700
rect 112190 79690 112310 79700
rect 112440 79690 112560 79700
rect 112690 79690 112810 79700
rect 112940 79690 113060 79700
rect 113190 79690 113310 79700
rect 113440 79690 113560 79700
rect 113690 79690 113810 79700
rect 113940 79690 114060 79700
rect 114190 79690 114310 79700
rect 114440 79690 114560 79700
rect 114690 79690 114810 79700
rect 114940 79690 115060 79700
rect 115190 79690 115310 79700
rect 115440 79690 115560 79700
rect 115690 79690 115810 79700
rect 115940 79690 116000 79700
rect 107000 79560 107050 79690
rect 107200 79560 107300 79690
rect 107450 79560 107550 79690
rect 107700 79560 107800 79690
rect 107950 79560 108050 79690
rect 108200 79560 108300 79690
rect 108450 79560 108550 79690
rect 108700 79560 108800 79690
rect 108950 79560 109050 79690
rect 109200 79560 109300 79690
rect 109450 79560 109550 79690
rect 109700 79560 109800 79690
rect 109950 79560 110050 79690
rect 110200 79560 110300 79690
rect 110450 79560 110550 79690
rect 110700 79560 110800 79690
rect 110950 79560 111050 79690
rect 111200 79560 111300 79690
rect 111450 79560 111550 79690
rect 111700 79560 111800 79690
rect 111950 79560 112050 79690
rect 112200 79560 112300 79690
rect 112450 79560 112550 79690
rect 112700 79560 112800 79690
rect 112950 79560 113050 79690
rect 113200 79560 113300 79690
rect 113450 79560 113550 79690
rect 113700 79560 113800 79690
rect 113950 79560 114050 79690
rect 114200 79560 114300 79690
rect 114450 79560 114550 79690
rect 114700 79560 114800 79690
rect 114950 79560 115050 79690
rect 115200 79560 115300 79690
rect 115450 79560 115550 79690
rect 115700 79560 115800 79690
rect 115950 79560 116000 79690
rect 107000 79550 107060 79560
rect 107190 79550 107310 79560
rect 107440 79550 107560 79560
rect 107690 79550 107810 79560
rect 107940 79550 108060 79560
rect 108190 79550 108310 79560
rect 108440 79550 108560 79560
rect 108690 79550 108810 79560
rect 108940 79550 109060 79560
rect 109190 79550 109310 79560
rect 109440 79550 109560 79560
rect 109690 79550 109810 79560
rect 109940 79550 110060 79560
rect 110190 79550 110310 79560
rect 110440 79550 110560 79560
rect 110690 79550 110810 79560
rect 110940 79550 111060 79560
rect 111190 79550 111310 79560
rect 111440 79550 111560 79560
rect 111690 79550 111810 79560
rect 111940 79550 112060 79560
rect 112190 79550 112310 79560
rect 112440 79550 112560 79560
rect 112690 79550 112810 79560
rect 112940 79550 113060 79560
rect 113190 79550 113310 79560
rect 113440 79550 113560 79560
rect 113690 79550 113810 79560
rect 113940 79550 114060 79560
rect 114190 79550 114310 79560
rect 114440 79550 114560 79560
rect 114690 79550 114810 79560
rect 114940 79550 115060 79560
rect 115190 79550 115310 79560
rect 115440 79550 115560 79560
rect 115690 79550 115810 79560
rect 115940 79550 116000 79560
rect 107000 79450 116000 79550
rect 107000 79440 107060 79450
rect 107190 79440 107310 79450
rect 107440 79440 107560 79450
rect 107690 79440 107810 79450
rect 107940 79440 108060 79450
rect 108190 79440 108310 79450
rect 108440 79440 108560 79450
rect 108690 79440 108810 79450
rect 108940 79440 109060 79450
rect 109190 79440 109310 79450
rect 109440 79440 109560 79450
rect 109690 79440 109810 79450
rect 109940 79440 110060 79450
rect 110190 79440 110310 79450
rect 110440 79440 110560 79450
rect 110690 79440 110810 79450
rect 110940 79440 111060 79450
rect 111190 79440 111310 79450
rect 111440 79440 111560 79450
rect 111690 79440 111810 79450
rect 111940 79440 112060 79450
rect 112190 79440 112310 79450
rect 112440 79440 112560 79450
rect 112690 79440 112810 79450
rect 112940 79440 113060 79450
rect 113190 79440 113310 79450
rect 113440 79440 113560 79450
rect 113690 79440 113810 79450
rect 113940 79440 114060 79450
rect 114190 79440 114310 79450
rect 114440 79440 114560 79450
rect 114690 79440 114810 79450
rect 114940 79440 115060 79450
rect 115190 79440 115310 79450
rect 115440 79440 115560 79450
rect 115690 79440 115810 79450
rect 115940 79440 116000 79450
rect 107000 79310 107050 79440
rect 107200 79310 107300 79440
rect 107450 79310 107550 79440
rect 107700 79310 107800 79440
rect 107950 79310 108050 79440
rect 108200 79310 108300 79440
rect 108450 79310 108550 79440
rect 108700 79310 108800 79440
rect 108950 79310 109050 79440
rect 109200 79310 109300 79440
rect 109450 79310 109550 79440
rect 109700 79310 109800 79440
rect 109950 79310 110050 79440
rect 110200 79310 110300 79440
rect 110450 79310 110550 79440
rect 110700 79310 110800 79440
rect 110950 79310 111050 79440
rect 111200 79310 111300 79440
rect 111450 79310 111550 79440
rect 111700 79310 111800 79440
rect 111950 79310 112050 79440
rect 112200 79310 112300 79440
rect 112450 79310 112550 79440
rect 112700 79310 112800 79440
rect 112950 79310 113050 79440
rect 113200 79310 113300 79440
rect 113450 79310 113550 79440
rect 113700 79310 113800 79440
rect 113950 79310 114050 79440
rect 114200 79310 114300 79440
rect 114450 79310 114550 79440
rect 114700 79310 114800 79440
rect 114950 79310 115050 79440
rect 115200 79310 115300 79440
rect 115450 79310 115550 79440
rect 115700 79310 115800 79440
rect 115950 79310 116000 79440
rect 107000 79300 107060 79310
rect 107190 79300 107310 79310
rect 107440 79300 107560 79310
rect 107690 79300 107810 79310
rect 107940 79300 108060 79310
rect 108190 79300 108310 79310
rect 108440 79300 108560 79310
rect 108690 79300 108810 79310
rect 108940 79300 109060 79310
rect 109190 79300 109310 79310
rect 109440 79300 109560 79310
rect 109690 79300 109810 79310
rect 109940 79300 110060 79310
rect 110190 79300 110310 79310
rect 110440 79300 110560 79310
rect 110690 79300 110810 79310
rect 110940 79300 111060 79310
rect 111190 79300 111310 79310
rect 111440 79300 111560 79310
rect 111690 79300 111810 79310
rect 111940 79300 112060 79310
rect 112190 79300 112310 79310
rect 112440 79300 112560 79310
rect 112690 79300 112810 79310
rect 112940 79300 113060 79310
rect 113190 79300 113310 79310
rect 113440 79300 113560 79310
rect 113690 79300 113810 79310
rect 113940 79300 114060 79310
rect 114190 79300 114310 79310
rect 114440 79300 114560 79310
rect 114690 79300 114810 79310
rect 114940 79300 115060 79310
rect 115190 79300 115310 79310
rect 115440 79300 115560 79310
rect 115690 79300 115810 79310
rect 115940 79300 116000 79310
rect 107000 79200 116000 79300
rect 107000 79190 107060 79200
rect 107190 79190 107310 79200
rect 107440 79190 107560 79200
rect 107690 79190 107810 79200
rect 107940 79190 108060 79200
rect 108190 79190 108310 79200
rect 108440 79190 108560 79200
rect 108690 79190 108810 79200
rect 108940 79190 109060 79200
rect 109190 79190 109310 79200
rect 109440 79190 109560 79200
rect 109690 79190 109810 79200
rect 109940 79190 110060 79200
rect 110190 79190 110310 79200
rect 110440 79190 110560 79200
rect 110690 79190 110810 79200
rect 110940 79190 111060 79200
rect 111190 79190 111310 79200
rect 111440 79190 111560 79200
rect 111690 79190 111810 79200
rect 111940 79190 112060 79200
rect 112190 79190 112310 79200
rect 112440 79190 112560 79200
rect 112690 79190 112810 79200
rect 112940 79190 113060 79200
rect 113190 79190 113310 79200
rect 113440 79190 113560 79200
rect 113690 79190 113810 79200
rect 113940 79190 114060 79200
rect 114190 79190 114310 79200
rect 114440 79190 114560 79200
rect 114690 79190 114810 79200
rect 114940 79190 115060 79200
rect 115190 79190 115310 79200
rect 115440 79190 115560 79200
rect 115690 79190 115810 79200
rect 115940 79190 116000 79200
rect 107000 79060 107050 79190
rect 107200 79060 107300 79190
rect 107450 79060 107550 79190
rect 107700 79060 107800 79190
rect 107950 79060 108050 79190
rect 108200 79060 108300 79190
rect 108450 79060 108550 79190
rect 108700 79060 108800 79190
rect 108950 79060 109050 79190
rect 109200 79060 109300 79190
rect 109450 79060 109550 79190
rect 109700 79060 109800 79190
rect 109950 79060 110050 79190
rect 110200 79060 110300 79190
rect 110450 79060 110550 79190
rect 110700 79060 110800 79190
rect 110950 79060 111050 79190
rect 111200 79060 111300 79190
rect 111450 79060 111550 79190
rect 111700 79060 111800 79190
rect 111950 79060 112050 79190
rect 112200 79060 112300 79190
rect 112450 79060 112550 79190
rect 112700 79060 112800 79190
rect 112950 79060 113050 79190
rect 113200 79060 113300 79190
rect 113450 79060 113550 79190
rect 113700 79060 113800 79190
rect 113950 79060 114050 79190
rect 114200 79060 114300 79190
rect 114450 79060 114550 79190
rect 114700 79060 114800 79190
rect 114950 79060 115050 79190
rect 115200 79060 115300 79190
rect 115450 79060 115550 79190
rect 115700 79060 115800 79190
rect 115950 79060 116000 79190
rect 107000 79050 107060 79060
rect 107190 79050 107310 79060
rect 107440 79050 107560 79060
rect 107690 79050 107810 79060
rect 107940 79050 108060 79060
rect 108190 79050 108310 79060
rect 108440 79050 108560 79060
rect 108690 79050 108810 79060
rect 108940 79050 109060 79060
rect 109190 79050 109310 79060
rect 109440 79050 109560 79060
rect 109690 79050 109810 79060
rect 109940 79050 110060 79060
rect 110190 79050 110310 79060
rect 110440 79050 110560 79060
rect 110690 79050 110810 79060
rect 110940 79050 111060 79060
rect 111190 79050 111310 79060
rect 111440 79050 111560 79060
rect 111690 79050 111810 79060
rect 111940 79050 112060 79060
rect 112190 79050 112310 79060
rect 112440 79050 112560 79060
rect 112690 79050 112810 79060
rect 112940 79050 113060 79060
rect 113190 79050 113310 79060
rect 113440 79050 113560 79060
rect 113690 79050 113810 79060
rect 113940 79050 114060 79060
rect 114190 79050 114310 79060
rect 114440 79050 114560 79060
rect 114690 79050 114810 79060
rect 114940 79050 115060 79060
rect 115190 79050 115310 79060
rect 115440 79050 115560 79060
rect 115690 79050 115810 79060
rect 115940 79050 116000 79060
rect 107000 78950 116000 79050
rect 107000 78940 107060 78950
rect 107190 78940 107310 78950
rect 107440 78940 107560 78950
rect 107690 78940 107810 78950
rect 107940 78940 108060 78950
rect 108190 78940 108310 78950
rect 108440 78940 108560 78950
rect 108690 78940 108810 78950
rect 108940 78940 109060 78950
rect 109190 78940 109310 78950
rect 109440 78940 109560 78950
rect 109690 78940 109810 78950
rect 109940 78940 110060 78950
rect 110190 78940 110310 78950
rect 110440 78940 110560 78950
rect 110690 78940 110810 78950
rect 110940 78940 111060 78950
rect 111190 78940 111310 78950
rect 111440 78940 111560 78950
rect 111690 78940 111810 78950
rect 111940 78940 112060 78950
rect 112190 78940 112310 78950
rect 112440 78940 112560 78950
rect 112690 78940 112810 78950
rect 112940 78940 113060 78950
rect 113190 78940 113310 78950
rect 113440 78940 113560 78950
rect 113690 78940 113810 78950
rect 113940 78940 114060 78950
rect 114190 78940 114310 78950
rect 114440 78940 114560 78950
rect 114690 78940 114810 78950
rect 114940 78940 115060 78950
rect 115190 78940 115310 78950
rect 115440 78940 115560 78950
rect 115690 78940 115810 78950
rect 115940 78940 116000 78950
rect 107000 78810 107050 78940
rect 107200 78810 107300 78940
rect 107450 78810 107550 78940
rect 107700 78810 107800 78940
rect 107950 78810 108050 78940
rect 108200 78810 108300 78940
rect 108450 78810 108550 78940
rect 108700 78810 108800 78940
rect 108950 78810 109050 78940
rect 109200 78810 109300 78940
rect 109450 78810 109550 78940
rect 109700 78810 109800 78940
rect 109950 78810 110050 78940
rect 110200 78810 110300 78940
rect 110450 78810 110550 78940
rect 110700 78810 110800 78940
rect 110950 78810 111050 78940
rect 111200 78810 111300 78940
rect 111450 78810 111550 78940
rect 111700 78810 111800 78940
rect 111950 78810 112050 78940
rect 112200 78810 112300 78940
rect 112450 78810 112550 78940
rect 112700 78810 112800 78940
rect 112950 78810 113050 78940
rect 113200 78810 113300 78940
rect 113450 78810 113550 78940
rect 113700 78810 113800 78940
rect 113950 78810 114050 78940
rect 114200 78810 114300 78940
rect 114450 78810 114550 78940
rect 114700 78810 114800 78940
rect 114950 78810 115050 78940
rect 115200 78810 115300 78940
rect 115450 78810 115550 78940
rect 115700 78810 115800 78940
rect 115950 78810 116000 78940
rect 107000 78800 107060 78810
rect 107190 78800 107310 78810
rect 107440 78800 107560 78810
rect 107690 78800 107810 78810
rect 107940 78800 108060 78810
rect 108190 78800 108310 78810
rect 108440 78800 108560 78810
rect 108690 78800 108810 78810
rect 108940 78800 109060 78810
rect 109190 78800 109310 78810
rect 109440 78800 109560 78810
rect 109690 78800 109810 78810
rect 109940 78800 110060 78810
rect 110190 78800 110310 78810
rect 110440 78800 110560 78810
rect 110690 78800 110810 78810
rect 110940 78800 111060 78810
rect 111190 78800 111310 78810
rect 111440 78800 111560 78810
rect 111690 78800 111810 78810
rect 111940 78800 112060 78810
rect 112190 78800 112310 78810
rect 112440 78800 112560 78810
rect 112690 78800 112810 78810
rect 112940 78800 113060 78810
rect 113190 78800 113310 78810
rect 113440 78800 113560 78810
rect 113690 78800 113810 78810
rect 113940 78800 114060 78810
rect 114190 78800 114310 78810
rect 114440 78800 114560 78810
rect 114690 78800 114810 78810
rect 114940 78800 115060 78810
rect 115190 78800 115310 78810
rect 115440 78800 115560 78810
rect 115690 78800 115810 78810
rect 115940 78800 116000 78810
rect 107000 78700 116000 78800
rect 107000 78690 107060 78700
rect 107190 78690 107310 78700
rect 107440 78690 107560 78700
rect 107690 78690 107810 78700
rect 107940 78690 108060 78700
rect 108190 78690 108310 78700
rect 108440 78690 108560 78700
rect 108690 78690 108810 78700
rect 108940 78690 109060 78700
rect 109190 78690 109310 78700
rect 109440 78690 109560 78700
rect 109690 78690 109810 78700
rect 109940 78690 110060 78700
rect 110190 78690 110310 78700
rect 110440 78690 110560 78700
rect 110690 78690 110810 78700
rect 110940 78690 111060 78700
rect 111190 78690 111310 78700
rect 111440 78690 111560 78700
rect 111690 78690 111810 78700
rect 111940 78690 112060 78700
rect 112190 78690 112310 78700
rect 112440 78690 112560 78700
rect 112690 78690 112810 78700
rect 112940 78690 113060 78700
rect 113190 78690 113310 78700
rect 113440 78690 113560 78700
rect 113690 78690 113810 78700
rect 113940 78690 114060 78700
rect 114190 78690 114310 78700
rect 114440 78690 114560 78700
rect 114690 78690 114810 78700
rect 114940 78690 115060 78700
rect 115190 78690 115310 78700
rect 115440 78690 115560 78700
rect 115690 78690 115810 78700
rect 115940 78690 116000 78700
rect 107000 78560 107050 78690
rect 107200 78560 107300 78690
rect 107450 78560 107550 78690
rect 107700 78560 107800 78690
rect 107950 78560 108050 78690
rect 108200 78560 108300 78690
rect 108450 78560 108550 78690
rect 108700 78560 108800 78690
rect 108950 78560 109050 78690
rect 109200 78560 109300 78690
rect 109450 78560 109550 78690
rect 109700 78560 109800 78690
rect 109950 78560 110050 78690
rect 110200 78560 110300 78690
rect 110450 78560 110550 78690
rect 110700 78560 110800 78690
rect 110950 78560 111050 78690
rect 111200 78560 111300 78690
rect 111450 78560 111550 78690
rect 111700 78560 111800 78690
rect 111950 78560 112050 78690
rect 112200 78560 112300 78690
rect 112450 78560 112550 78690
rect 112700 78560 112800 78690
rect 112950 78560 113050 78690
rect 113200 78560 113300 78690
rect 113450 78560 113550 78690
rect 113700 78560 113800 78690
rect 113950 78560 114050 78690
rect 114200 78560 114300 78690
rect 114450 78560 114550 78690
rect 114700 78560 114800 78690
rect 114950 78560 115050 78690
rect 115200 78560 115300 78690
rect 115450 78560 115550 78690
rect 115700 78560 115800 78690
rect 115950 78560 116000 78690
rect 107000 78550 107060 78560
rect 107190 78550 107310 78560
rect 107440 78550 107560 78560
rect 107690 78550 107810 78560
rect 107940 78550 108060 78560
rect 108190 78550 108310 78560
rect 108440 78550 108560 78560
rect 108690 78550 108810 78560
rect 108940 78550 109060 78560
rect 109190 78550 109310 78560
rect 109440 78550 109560 78560
rect 109690 78550 109810 78560
rect 109940 78550 110060 78560
rect 110190 78550 110310 78560
rect 110440 78550 110560 78560
rect 110690 78550 110810 78560
rect 110940 78550 111060 78560
rect 111190 78550 111310 78560
rect 111440 78550 111560 78560
rect 111690 78550 111810 78560
rect 111940 78550 112060 78560
rect 112190 78550 112310 78560
rect 112440 78550 112560 78560
rect 112690 78550 112810 78560
rect 112940 78550 113060 78560
rect 113190 78550 113310 78560
rect 113440 78550 113560 78560
rect 113690 78550 113810 78560
rect 113940 78550 114060 78560
rect 114190 78550 114310 78560
rect 114440 78550 114560 78560
rect 114690 78550 114810 78560
rect 114940 78550 115060 78560
rect 115190 78550 115310 78560
rect 115440 78550 115560 78560
rect 115690 78550 115810 78560
rect 115940 78550 116000 78560
rect 107000 78450 116000 78550
rect 107000 78440 107060 78450
rect 107190 78440 107310 78450
rect 107440 78440 107560 78450
rect 107690 78440 107810 78450
rect 107940 78440 108060 78450
rect 108190 78440 108310 78450
rect 108440 78440 108560 78450
rect 108690 78440 108810 78450
rect 108940 78440 109060 78450
rect 109190 78440 109310 78450
rect 109440 78440 109560 78450
rect 109690 78440 109810 78450
rect 109940 78440 110060 78450
rect 110190 78440 110310 78450
rect 110440 78440 110560 78450
rect 110690 78440 110810 78450
rect 110940 78440 111060 78450
rect 111190 78440 111310 78450
rect 111440 78440 111560 78450
rect 111690 78440 111810 78450
rect 111940 78440 112060 78450
rect 112190 78440 112310 78450
rect 112440 78440 112560 78450
rect 112690 78440 112810 78450
rect 112940 78440 113060 78450
rect 113190 78440 113310 78450
rect 113440 78440 113560 78450
rect 113690 78440 113810 78450
rect 113940 78440 114060 78450
rect 114190 78440 114310 78450
rect 114440 78440 114560 78450
rect 114690 78440 114810 78450
rect 114940 78440 115060 78450
rect 115190 78440 115310 78450
rect 115440 78440 115560 78450
rect 115690 78440 115810 78450
rect 115940 78440 116000 78450
rect 107000 78310 107050 78440
rect 107200 78310 107300 78440
rect 107450 78310 107550 78440
rect 107700 78310 107800 78440
rect 107950 78310 108050 78440
rect 108200 78310 108300 78440
rect 108450 78310 108550 78440
rect 108700 78310 108800 78440
rect 108950 78310 109050 78440
rect 109200 78310 109300 78440
rect 109450 78310 109550 78440
rect 109700 78310 109800 78440
rect 109950 78310 110050 78440
rect 110200 78310 110300 78440
rect 110450 78310 110550 78440
rect 110700 78310 110800 78440
rect 110950 78310 111050 78440
rect 111200 78310 111300 78440
rect 111450 78310 111550 78440
rect 111700 78310 111800 78440
rect 111950 78310 112050 78440
rect 112200 78310 112300 78440
rect 112450 78310 112550 78440
rect 112700 78310 112800 78440
rect 112950 78310 113050 78440
rect 113200 78310 113300 78440
rect 113450 78310 113550 78440
rect 113700 78310 113800 78440
rect 113950 78310 114050 78440
rect 114200 78310 114300 78440
rect 114450 78310 114550 78440
rect 114700 78310 114800 78440
rect 114950 78310 115050 78440
rect 115200 78310 115300 78440
rect 115450 78310 115550 78440
rect 115700 78310 115800 78440
rect 115950 78310 116000 78440
rect 107000 78300 107060 78310
rect 107190 78300 107310 78310
rect 107440 78300 107560 78310
rect 107690 78300 107810 78310
rect 107940 78300 108060 78310
rect 108190 78300 108310 78310
rect 108440 78300 108560 78310
rect 108690 78300 108810 78310
rect 108940 78300 109060 78310
rect 109190 78300 109310 78310
rect 109440 78300 109560 78310
rect 109690 78300 109810 78310
rect 109940 78300 110060 78310
rect 110190 78300 110310 78310
rect 110440 78300 110560 78310
rect 110690 78300 110810 78310
rect 110940 78300 111060 78310
rect 111190 78300 111310 78310
rect 111440 78300 111560 78310
rect 111690 78300 111810 78310
rect 111940 78300 112060 78310
rect 112190 78300 112310 78310
rect 112440 78300 112560 78310
rect 112690 78300 112810 78310
rect 112940 78300 113060 78310
rect 113190 78300 113310 78310
rect 113440 78300 113560 78310
rect 113690 78300 113810 78310
rect 113940 78300 114060 78310
rect 114190 78300 114310 78310
rect 114440 78300 114560 78310
rect 114690 78300 114810 78310
rect 114940 78300 115060 78310
rect 115190 78300 115310 78310
rect 115440 78300 115560 78310
rect 115690 78300 115810 78310
rect 115940 78300 116000 78310
rect 107000 78200 116000 78300
rect 107000 78190 107060 78200
rect 107190 78190 107310 78200
rect 107440 78190 107560 78200
rect 107690 78190 107810 78200
rect 107940 78190 108060 78200
rect 108190 78190 108310 78200
rect 108440 78190 108560 78200
rect 108690 78190 108810 78200
rect 108940 78190 109060 78200
rect 109190 78190 109310 78200
rect 109440 78190 109560 78200
rect 109690 78190 109810 78200
rect 109940 78190 110060 78200
rect 110190 78190 110310 78200
rect 110440 78190 110560 78200
rect 110690 78190 110810 78200
rect 110940 78190 111060 78200
rect 111190 78190 111310 78200
rect 111440 78190 111560 78200
rect 111690 78190 111810 78200
rect 111940 78190 112060 78200
rect 112190 78190 112310 78200
rect 112440 78190 112560 78200
rect 112690 78190 112810 78200
rect 112940 78190 113060 78200
rect 113190 78190 113310 78200
rect 113440 78190 113560 78200
rect 113690 78190 113810 78200
rect 113940 78190 114060 78200
rect 114190 78190 114310 78200
rect 114440 78190 114560 78200
rect 114690 78190 114810 78200
rect 114940 78190 115060 78200
rect 115190 78190 115310 78200
rect 115440 78190 115560 78200
rect 115690 78190 115810 78200
rect 115940 78190 116000 78200
rect 107000 78060 107050 78190
rect 107200 78060 107300 78190
rect 107450 78060 107550 78190
rect 107700 78060 107800 78190
rect 107950 78060 108050 78190
rect 108200 78060 108300 78190
rect 108450 78060 108550 78190
rect 108700 78060 108800 78190
rect 108950 78060 109050 78190
rect 109200 78060 109300 78190
rect 109450 78060 109550 78190
rect 109700 78060 109800 78190
rect 109950 78060 110050 78190
rect 110200 78060 110300 78190
rect 110450 78060 110550 78190
rect 110700 78060 110800 78190
rect 110950 78060 111050 78190
rect 111200 78060 111300 78190
rect 111450 78060 111550 78190
rect 111700 78060 111800 78190
rect 111950 78060 112050 78190
rect 112200 78060 112300 78190
rect 112450 78060 112550 78190
rect 112700 78060 112800 78190
rect 112950 78060 113050 78190
rect 113200 78060 113300 78190
rect 113450 78060 113550 78190
rect 113700 78060 113800 78190
rect 113950 78060 114050 78190
rect 114200 78060 114300 78190
rect 114450 78060 114550 78190
rect 114700 78060 114800 78190
rect 114950 78060 115050 78190
rect 115200 78060 115300 78190
rect 115450 78060 115550 78190
rect 115700 78060 115800 78190
rect 115950 78060 116000 78190
rect 107000 78050 107060 78060
rect 107190 78050 107310 78060
rect 107440 78050 107560 78060
rect 107690 78050 107810 78060
rect 107940 78050 108060 78060
rect 108190 78050 108310 78060
rect 108440 78050 108560 78060
rect 108690 78050 108810 78060
rect 108940 78050 109060 78060
rect 109190 78050 109310 78060
rect 109440 78050 109560 78060
rect 109690 78050 109810 78060
rect 109940 78050 110060 78060
rect 110190 78050 110310 78060
rect 110440 78050 110560 78060
rect 110690 78050 110810 78060
rect 110940 78050 111060 78060
rect 111190 78050 111310 78060
rect 111440 78050 111560 78060
rect 111690 78050 111810 78060
rect 111940 78050 112060 78060
rect 112190 78050 112310 78060
rect 112440 78050 112560 78060
rect 112690 78050 112810 78060
rect 112940 78050 113060 78060
rect 113190 78050 113310 78060
rect 113440 78050 113560 78060
rect 113690 78050 113810 78060
rect 113940 78050 114060 78060
rect 114190 78050 114310 78060
rect 114440 78050 114560 78060
rect 114690 78050 114810 78060
rect 114940 78050 115060 78060
rect 115190 78050 115310 78060
rect 115440 78050 115560 78060
rect 115690 78050 115810 78060
rect 115940 78050 116000 78060
rect 107000 77950 116000 78050
rect 107000 77940 107060 77950
rect 107190 77940 107310 77950
rect 107440 77940 107560 77950
rect 107690 77940 107810 77950
rect 107940 77940 108060 77950
rect 108190 77940 108310 77950
rect 108440 77940 108560 77950
rect 108690 77940 108810 77950
rect 108940 77940 109060 77950
rect 109190 77940 109310 77950
rect 109440 77940 109560 77950
rect 109690 77940 109810 77950
rect 109940 77940 110060 77950
rect 110190 77940 110310 77950
rect 110440 77940 110560 77950
rect 110690 77940 110810 77950
rect 110940 77940 111060 77950
rect 111190 77940 111310 77950
rect 111440 77940 111560 77950
rect 111690 77940 111810 77950
rect 111940 77940 112060 77950
rect 112190 77940 112310 77950
rect 112440 77940 112560 77950
rect 112690 77940 112810 77950
rect 112940 77940 113060 77950
rect 113190 77940 113310 77950
rect 113440 77940 113560 77950
rect 113690 77940 113810 77950
rect 113940 77940 114060 77950
rect 114190 77940 114310 77950
rect 114440 77940 114560 77950
rect 114690 77940 114810 77950
rect 114940 77940 115060 77950
rect 115190 77940 115310 77950
rect 115440 77940 115560 77950
rect 115690 77940 115810 77950
rect 115940 77940 116000 77950
rect 107000 77810 107050 77940
rect 107200 77810 107300 77940
rect 107450 77810 107550 77940
rect 107700 77810 107800 77940
rect 107950 77810 108050 77940
rect 108200 77810 108300 77940
rect 108450 77810 108550 77940
rect 108700 77810 108800 77940
rect 108950 77810 109050 77940
rect 109200 77810 109300 77940
rect 109450 77810 109550 77940
rect 109700 77810 109800 77940
rect 109950 77810 110050 77940
rect 110200 77810 110300 77940
rect 110450 77810 110550 77940
rect 110700 77810 110800 77940
rect 110950 77810 111050 77940
rect 111200 77810 111300 77940
rect 111450 77810 111550 77940
rect 111700 77810 111800 77940
rect 111950 77810 112050 77940
rect 112200 77810 112300 77940
rect 112450 77810 112550 77940
rect 112700 77810 112800 77940
rect 112950 77810 113050 77940
rect 113200 77810 113300 77940
rect 113450 77810 113550 77940
rect 113700 77810 113800 77940
rect 113950 77810 114050 77940
rect 114200 77810 114300 77940
rect 114450 77810 114550 77940
rect 114700 77810 114800 77940
rect 114950 77810 115050 77940
rect 115200 77810 115300 77940
rect 115450 77810 115550 77940
rect 115700 77810 115800 77940
rect 115950 77810 116000 77940
rect 107000 77800 107060 77810
rect 107190 77800 107310 77810
rect 107440 77800 107560 77810
rect 107690 77800 107810 77810
rect 107940 77800 108060 77810
rect 108190 77800 108310 77810
rect 108440 77800 108560 77810
rect 108690 77800 108810 77810
rect 108940 77800 109060 77810
rect 109190 77800 109310 77810
rect 109440 77800 109560 77810
rect 109690 77800 109810 77810
rect 109940 77800 110060 77810
rect 110190 77800 110310 77810
rect 110440 77800 110560 77810
rect 110690 77800 110810 77810
rect 110940 77800 111060 77810
rect 111190 77800 111310 77810
rect 111440 77800 111560 77810
rect 111690 77800 111810 77810
rect 111940 77800 112060 77810
rect 112190 77800 112310 77810
rect 112440 77800 112560 77810
rect 112690 77800 112810 77810
rect 112940 77800 113060 77810
rect 113190 77800 113310 77810
rect 113440 77800 113560 77810
rect 113690 77800 113810 77810
rect 113940 77800 114060 77810
rect 114190 77800 114310 77810
rect 114440 77800 114560 77810
rect 114690 77800 114810 77810
rect 114940 77800 115060 77810
rect 115190 77800 115310 77810
rect 115440 77800 115560 77810
rect 115690 77800 115810 77810
rect 115940 77800 116000 77810
rect 107000 77700 116000 77800
rect 107000 77690 107060 77700
rect 107190 77690 107310 77700
rect 107440 77690 107560 77700
rect 107690 77690 107810 77700
rect 107940 77690 108060 77700
rect 108190 77690 108310 77700
rect 108440 77690 108560 77700
rect 108690 77690 108810 77700
rect 108940 77690 109060 77700
rect 109190 77690 109310 77700
rect 109440 77690 109560 77700
rect 109690 77690 109810 77700
rect 109940 77690 110060 77700
rect 110190 77690 110310 77700
rect 110440 77690 110560 77700
rect 110690 77690 110810 77700
rect 110940 77690 111060 77700
rect 111190 77690 111310 77700
rect 111440 77690 111560 77700
rect 111690 77690 111810 77700
rect 111940 77690 112060 77700
rect 112190 77690 112310 77700
rect 112440 77690 112560 77700
rect 112690 77690 112810 77700
rect 112940 77690 113060 77700
rect 113190 77690 113310 77700
rect 113440 77690 113560 77700
rect 113690 77690 113810 77700
rect 113940 77690 114060 77700
rect 114190 77690 114310 77700
rect 114440 77690 114560 77700
rect 114690 77690 114810 77700
rect 114940 77690 115060 77700
rect 115190 77690 115310 77700
rect 115440 77690 115560 77700
rect 115690 77690 115810 77700
rect 115940 77690 116000 77700
rect 107000 77560 107050 77690
rect 107200 77560 107300 77690
rect 107450 77560 107550 77690
rect 107700 77560 107800 77690
rect 107950 77560 108050 77690
rect 108200 77560 108300 77690
rect 108450 77560 108550 77690
rect 108700 77560 108800 77690
rect 108950 77560 109050 77690
rect 109200 77560 109300 77690
rect 109450 77560 109550 77690
rect 109700 77560 109800 77690
rect 109950 77560 110050 77690
rect 110200 77560 110300 77690
rect 110450 77560 110550 77690
rect 110700 77560 110800 77690
rect 110950 77560 111050 77690
rect 111200 77560 111300 77690
rect 111450 77560 111550 77690
rect 111700 77560 111800 77690
rect 111950 77560 112050 77690
rect 112200 77560 112300 77690
rect 112450 77560 112550 77690
rect 112700 77560 112800 77690
rect 112950 77560 113050 77690
rect 113200 77560 113300 77690
rect 113450 77560 113550 77690
rect 113700 77560 113800 77690
rect 113950 77560 114050 77690
rect 114200 77560 114300 77690
rect 114450 77560 114550 77690
rect 114700 77560 114800 77690
rect 114950 77560 115050 77690
rect 115200 77560 115300 77690
rect 115450 77560 115550 77690
rect 115700 77560 115800 77690
rect 115950 77560 116000 77690
rect 107000 77550 107060 77560
rect 107190 77550 107310 77560
rect 107440 77550 107560 77560
rect 107690 77550 107810 77560
rect 107940 77550 108060 77560
rect 108190 77550 108310 77560
rect 108440 77550 108560 77560
rect 108690 77550 108810 77560
rect 108940 77550 109060 77560
rect 109190 77550 109310 77560
rect 109440 77550 109560 77560
rect 109690 77550 109810 77560
rect 109940 77550 110060 77560
rect 110190 77550 110310 77560
rect 110440 77550 110560 77560
rect 110690 77550 110810 77560
rect 110940 77550 111060 77560
rect 111190 77550 111310 77560
rect 111440 77550 111560 77560
rect 111690 77550 111810 77560
rect 111940 77550 112060 77560
rect 112190 77550 112310 77560
rect 112440 77550 112560 77560
rect 112690 77550 112810 77560
rect 112940 77550 113060 77560
rect 113190 77550 113310 77560
rect 113440 77550 113560 77560
rect 113690 77550 113810 77560
rect 113940 77550 114060 77560
rect 114190 77550 114310 77560
rect 114440 77550 114560 77560
rect 114690 77550 114810 77560
rect 114940 77550 115060 77560
rect 115190 77550 115310 77560
rect 115440 77550 115560 77560
rect 115690 77550 115810 77560
rect 115940 77550 116000 77560
rect 107000 77450 116000 77550
rect 107000 77440 107060 77450
rect 107190 77440 107310 77450
rect 107440 77440 107560 77450
rect 107690 77440 107810 77450
rect 107940 77440 108060 77450
rect 108190 77440 108310 77450
rect 108440 77440 108560 77450
rect 108690 77440 108810 77450
rect 108940 77440 109060 77450
rect 109190 77440 109310 77450
rect 109440 77440 109560 77450
rect 109690 77440 109810 77450
rect 109940 77440 110060 77450
rect 110190 77440 110310 77450
rect 110440 77440 110560 77450
rect 110690 77440 110810 77450
rect 110940 77440 111060 77450
rect 111190 77440 111310 77450
rect 111440 77440 111560 77450
rect 111690 77440 111810 77450
rect 111940 77440 112060 77450
rect 112190 77440 112310 77450
rect 112440 77440 112560 77450
rect 112690 77440 112810 77450
rect 112940 77440 113060 77450
rect 113190 77440 113310 77450
rect 113440 77440 113560 77450
rect 113690 77440 113810 77450
rect 113940 77440 114060 77450
rect 114190 77440 114310 77450
rect 114440 77440 114560 77450
rect 114690 77440 114810 77450
rect 114940 77440 115060 77450
rect 115190 77440 115310 77450
rect 115440 77440 115560 77450
rect 115690 77440 115810 77450
rect 115940 77440 116000 77450
rect 107000 77310 107050 77440
rect 107200 77310 107300 77440
rect 107450 77310 107550 77440
rect 107700 77310 107800 77440
rect 107950 77310 108050 77440
rect 108200 77310 108300 77440
rect 108450 77310 108550 77440
rect 108700 77310 108800 77440
rect 108950 77310 109050 77440
rect 109200 77310 109300 77440
rect 109450 77310 109550 77440
rect 109700 77310 109800 77440
rect 109950 77310 110050 77440
rect 110200 77310 110300 77440
rect 110450 77310 110550 77440
rect 110700 77310 110800 77440
rect 110950 77310 111050 77440
rect 111200 77310 111300 77440
rect 111450 77310 111550 77440
rect 111700 77310 111800 77440
rect 111950 77310 112050 77440
rect 112200 77310 112300 77440
rect 112450 77310 112550 77440
rect 112700 77310 112800 77440
rect 112950 77310 113050 77440
rect 113200 77310 113300 77440
rect 113450 77310 113550 77440
rect 113700 77310 113800 77440
rect 113950 77310 114050 77440
rect 114200 77310 114300 77440
rect 114450 77310 114550 77440
rect 114700 77310 114800 77440
rect 114950 77310 115050 77440
rect 115200 77310 115300 77440
rect 115450 77310 115550 77440
rect 115700 77310 115800 77440
rect 115950 77310 116000 77440
rect 107000 77300 107060 77310
rect 107190 77300 107310 77310
rect 107440 77300 107560 77310
rect 107690 77300 107810 77310
rect 107940 77300 108060 77310
rect 108190 77300 108310 77310
rect 108440 77300 108560 77310
rect 108690 77300 108810 77310
rect 108940 77300 109060 77310
rect 109190 77300 109310 77310
rect 109440 77300 109560 77310
rect 109690 77300 109810 77310
rect 109940 77300 110060 77310
rect 110190 77300 110310 77310
rect 110440 77300 110560 77310
rect 110690 77300 110810 77310
rect 110940 77300 111060 77310
rect 111190 77300 111310 77310
rect 111440 77300 111560 77310
rect 111690 77300 111810 77310
rect 111940 77300 112060 77310
rect 112190 77300 112310 77310
rect 112440 77300 112560 77310
rect 112690 77300 112810 77310
rect 112940 77300 113060 77310
rect 113190 77300 113310 77310
rect 113440 77300 113560 77310
rect 113690 77300 113810 77310
rect 113940 77300 114060 77310
rect 114190 77300 114310 77310
rect 114440 77300 114560 77310
rect 114690 77300 114810 77310
rect 114940 77300 115060 77310
rect 115190 77300 115310 77310
rect 115440 77300 115560 77310
rect 115690 77300 115810 77310
rect 115940 77300 116000 77310
rect 107000 77200 116000 77300
rect 107000 77190 107060 77200
rect 107190 77190 107310 77200
rect 107440 77190 107560 77200
rect 107690 77190 107810 77200
rect 107940 77190 108060 77200
rect 108190 77190 108310 77200
rect 108440 77190 108560 77200
rect 108690 77190 108810 77200
rect 108940 77190 109060 77200
rect 109190 77190 109310 77200
rect 109440 77190 109560 77200
rect 109690 77190 109810 77200
rect 109940 77190 110060 77200
rect 110190 77190 110310 77200
rect 110440 77190 110560 77200
rect 110690 77190 110810 77200
rect 110940 77190 111060 77200
rect 111190 77190 111310 77200
rect 111440 77190 111560 77200
rect 111690 77190 111810 77200
rect 111940 77190 112060 77200
rect 112190 77190 112310 77200
rect 112440 77190 112560 77200
rect 112690 77190 112810 77200
rect 112940 77190 113060 77200
rect 113190 77190 113310 77200
rect 113440 77190 113560 77200
rect 113690 77190 113810 77200
rect 113940 77190 114060 77200
rect 114190 77190 114310 77200
rect 114440 77190 114560 77200
rect 114690 77190 114810 77200
rect 114940 77190 115060 77200
rect 115190 77190 115310 77200
rect 115440 77190 115560 77200
rect 115690 77190 115810 77200
rect 115940 77190 116000 77200
rect 107000 77060 107050 77190
rect 107200 77060 107300 77190
rect 107450 77060 107550 77190
rect 107700 77060 107800 77190
rect 107950 77060 108050 77190
rect 108200 77060 108300 77190
rect 108450 77060 108550 77190
rect 108700 77060 108800 77190
rect 108950 77060 109050 77190
rect 109200 77060 109300 77190
rect 109450 77060 109550 77190
rect 109700 77060 109800 77190
rect 109950 77060 110050 77190
rect 110200 77060 110300 77190
rect 110450 77060 110550 77190
rect 110700 77060 110800 77190
rect 110950 77060 111050 77190
rect 111200 77060 111300 77190
rect 111450 77060 111550 77190
rect 111700 77060 111800 77190
rect 111950 77060 112050 77190
rect 112200 77060 112300 77190
rect 112450 77060 112550 77190
rect 112700 77060 112800 77190
rect 112950 77060 113050 77190
rect 113200 77060 113300 77190
rect 113450 77060 113550 77190
rect 113700 77060 113800 77190
rect 113950 77060 114050 77190
rect 114200 77060 114300 77190
rect 114450 77060 114550 77190
rect 114700 77060 114800 77190
rect 114950 77060 115050 77190
rect 115200 77060 115300 77190
rect 115450 77060 115550 77190
rect 115700 77060 115800 77190
rect 115950 77060 116000 77190
rect 107000 77050 107060 77060
rect 107190 77050 107310 77060
rect 107440 77050 107560 77060
rect 107690 77050 107810 77060
rect 107940 77050 108060 77060
rect 108190 77050 108310 77060
rect 108440 77050 108560 77060
rect 108690 77050 108810 77060
rect 108940 77050 109060 77060
rect 109190 77050 109310 77060
rect 109440 77050 109560 77060
rect 109690 77050 109810 77060
rect 109940 77050 110060 77060
rect 110190 77050 110310 77060
rect 110440 77050 110560 77060
rect 110690 77050 110810 77060
rect 110940 77050 111060 77060
rect 111190 77050 111310 77060
rect 111440 77050 111560 77060
rect 111690 77050 111810 77060
rect 111940 77050 112060 77060
rect 112190 77050 112310 77060
rect 112440 77050 112560 77060
rect 112690 77050 112810 77060
rect 112940 77050 113060 77060
rect 113190 77050 113310 77060
rect 113440 77050 113560 77060
rect 113690 77050 113810 77060
rect 113940 77050 114060 77060
rect 114190 77050 114310 77060
rect 114440 77050 114560 77060
rect 114690 77050 114810 77060
rect 114940 77050 115060 77060
rect 115190 77050 115310 77060
rect 115440 77050 115560 77060
rect 115690 77050 115810 77060
rect 115940 77050 116000 77060
rect 107000 77000 116000 77050
rect 89000 76950 116000 77000
rect 89000 76940 89060 76950
rect 89190 76940 89310 76950
rect 89440 76940 89560 76950
rect 89690 76940 89810 76950
rect 89940 76940 90060 76950
rect 90190 76940 90310 76950
rect 90440 76940 90560 76950
rect 90690 76940 90810 76950
rect 90940 76940 91060 76950
rect 91190 76940 91310 76950
rect 91440 76940 91560 76950
rect 91690 76940 91810 76950
rect 91940 76940 92060 76950
rect 92190 76940 92310 76950
rect 92440 76940 92560 76950
rect 92690 76940 92810 76950
rect 92940 76940 93060 76950
rect 93190 76940 93310 76950
rect 93440 76940 93560 76950
rect 93690 76940 93810 76950
rect 93940 76940 94060 76950
rect 94190 76940 94310 76950
rect 94440 76940 94560 76950
rect 94690 76940 94810 76950
rect 94940 76940 95060 76950
rect 95190 76940 95310 76950
rect 95440 76940 95560 76950
rect 95690 76940 95810 76950
rect 95940 76940 96060 76950
rect 96190 76940 96310 76950
rect 96440 76940 96560 76950
rect 96690 76940 96810 76950
rect 96940 76940 97060 76950
rect 97190 76940 97310 76950
rect 97440 76940 97560 76950
rect 97690 76940 97810 76950
rect 97940 76940 98060 76950
rect 98190 76940 98310 76950
rect 98440 76940 98560 76950
rect 98690 76940 98810 76950
rect 98940 76940 99060 76950
rect 99190 76940 99310 76950
rect 99440 76940 99560 76950
rect 99690 76940 99810 76950
rect 99940 76940 100060 76950
rect 100190 76940 100310 76950
rect 100440 76940 100560 76950
rect 100690 76940 100810 76950
rect 100940 76940 101060 76950
rect 101190 76940 101310 76950
rect 101440 76940 101560 76950
rect 101690 76940 101810 76950
rect 101940 76940 102060 76950
rect 102190 76940 102310 76950
rect 102440 76940 102560 76950
rect 102690 76940 102810 76950
rect 102940 76940 103060 76950
rect 103190 76940 103310 76950
rect 103440 76940 103560 76950
rect 103690 76940 103810 76950
rect 103940 76940 104060 76950
rect 104190 76940 104310 76950
rect 104440 76940 104560 76950
rect 104690 76940 104810 76950
rect 104940 76940 105060 76950
rect 105190 76940 105310 76950
rect 105440 76940 105560 76950
rect 105690 76940 105810 76950
rect 105940 76940 106060 76950
rect 106190 76940 106310 76950
rect 106440 76940 106560 76950
rect 106690 76940 106810 76950
rect 106940 76940 107060 76950
rect 107190 76940 107310 76950
rect 107440 76940 107560 76950
rect 107690 76940 107810 76950
rect 107940 76940 108060 76950
rect 108190 76940 108310 76950
rect 108440 76940 108560 76950
rect 108690 76940 108810 76950
rect 108940 76940 109060 76950
rect 109190 76940 109310 76950
rect 109440 76940 109560 76950
rect 109690 76940 109810 76950
rect 109940 76940 110060 76950
rect 110190 76940 110310 76950
rect 110440 76940 110560 76950
rect 110690 76940 110810 76950
rect 110940 76940 111060 76950
rect 111190 76940 111310 76950
rect 111440 76940 111560 76950
rect 111690 76940 111810 76950
rect 111940 76940 112060 76950
rect 112190 76940 112310 76950
rect 112440 76940 112560 76950
rect 112690 76940 112810 76950
rect 112940 76940 113060 76950
rect 113190 76940 113310 76950
rect 113440 76940 113560 76950
rect 113690 76940 113810 76950
rect 113940 76940 114060 76950
rect 114190 76940 114310 76950
rect 114440 76940 114560 76950
rect 114690 76940 114810 76950
rect 114940 76940 115060 76950
rect 115190 76940 115310 76950
rect 115440 76940 115560 76950
rect 115690 76940 115810 76950
rect 115940 76940 116000 76950
rect 89000 76810 89050 76940
rect 89200 76810 89300 76940
rect 89450 76810 89550 76940
rect 89700 76810 89800 76940
rect 89950 76810 90050 76940
rect 90200 76810 90300 76940
rect 90450 76810 90550 76940
rect 90700 76810 90800 76940
rect 90950 76810 91050 76940
rect 91200 76810 91300 76940
rect 91450 76810 91550 76940
rect 91700 76810 91800 76940
rect 91950 76810 92050 76940
rect 92200 76810 92300 76940
rect 92450 76810 92550 76940
rect 92700 76810 92800 76940
rect 92950 76810 93050 76940
rect 93200 76810 93300 76940
rect 93450 76810 93550 76940
rect 93700 76810 93800 76940
rect 93950 76810 94050 76940
rect 94200 76810 94300 76940
rect 94450 76810 94550 76940
rect 94700 76810 94800 76940
rect 94950 76810 95050 76940
rect 95200 76810 95300 76940
rect 95450 76810 95550 76940
rect 95700 76810 95800 76940
rect 95950 76810 96050 76940
rect 96200 76810 96300 76940
rect 96450 76810 96550 76940
rect 96700 76810 96800 76940
rect 96950 76810 97050 76940
rect 97200 76810 97300 76940
rect 97450 76810 97550 76940
rect 97700 76810 97800 76940
rect 97950 76810 98050 76940
rect 98200 76810 98300 76940
rect 98450 76810 98550 76940
rect 98700 76810 98800 76940
rect 98950 76810 99050 76940
rect 99200 76810 99300 76940
rect 99450 76810 99550 76940
rect 99700 76810 99800 76940
rect 99950 76810 100050 76940
rect 100200 76810 100300 76940
rect 100450 76810 100550 76940
rect 100700 76810 100800 76940
rect 100950 76810 101050 76940
rect 101200 76810 101300 76940
rect 101450 76810 101550 76940
rect 101700 76810 101800 76940
rect 101950 76810 102050 76940
rect 102200 76810 102300 76940
rect 102450 76810 102550 76940
rect 102700 76810 102800 76940
rect 102950 76810 103050 76940
rect 103200 76810 103300 76940
rect 103450 76810 103550 76940
rect 103700 76810 103800 76940
rect 103950 76810 104050 76940
rect 104200 76810 104300 76940
rect 104450 76810 104550 76940
rect 104700 76810 104800 76940
rect 104950 76810 105050 76940
rect 105200 76810 105300 76940
rect 105450 76810 105550 76940
rect 105700 76810 105800 76940
rect 105950 76810 106050 76940
rect 106200 76810 106300 76940
rect 106450 76810 106550 76940
rect 106700 76810 106800 76940
rect 106950 76810 107050 76940
rect 107200 76810 107300 76940
rect 107450 76810 107550 76940
rect 107700 76810 107800 76940
rect 107950 76810 108050 76940
rect 108200 76810 108300 76940
rect 108450 76810 108550 76940
rect 108700 76810 108800 76940
rect 108950 76810 109050 76940
rect 109200 76810 109300 76940
rect 109450 76810 109550 76940
rect 109700 76810 109800 76940
rect 109950 76810 110050 76940
rect 110200 76810 110300 76940
rect 110450 76810 110550 76940
rect 110700 76810 110800 76940
rect 110950 76810 111050 76940
rect 111200 76810 111300 76940
rect 111450 76810 111550 76940
rect 111700 76810 111800 76940
rect 111950 76810 112050 76940
rect 112200 76810 112300 76940
rect 112450 76810 112550 76940
rect 112700 76810 112800 76940
rect 112950 76810 113050 76940
rect 113200 76810 113300 76940
rect 113450 76810 113550 76940
rect 113700 76810 113800 76940
rect 113950 76810 114050 76940
rect 114200 76810 114300 76940
rect 114450 76810 114550 76940
rect 114700 76810 114800 76940
rect 114950 76810 115050 76940
rect 115200 76810 115300 76940
rect 115450 76810 115550 76940
rect 115700 76810 115800 76940
rect 115950 76810 116000 76940
rect 89000 76800 89060 76810
rect 89190 76800 89310 76810
rect 89440 76800 89560 76810
rect 89690 76800 89810 76810
rect 89940 76800 90060 76810
rect 90190 76800 90310 76810
rect 90440 76800 90560 76810
rect 90690 76800 90810 76810
rect 90940 76800 91060 76810
rect 91190 76800 91310 76810
rect 91440 76800 91560 76810
rect 91690 76800 91810 76810
rect 91940 76800 92060 76810
rect 92190 76800 92310 76810
rect 92440 76800 92560 76810
rect 92690 76800 92810 76810
rect 92940 76800 93060 76810
rect 93190 76800 93310 76810
rect 93440 76800 93560 76810
rect 93690 76800 93810 76810
rect 93940 76800 94060 76810
rect 94190 76800 94310 76810
rect 94440 76800 94560 76810
rect 94690 76800 94810 76810
rect 94940 76800 95060 76810
rect 95190 76800 95310 76810
rect 95440 76800 95560 76810
rect 95690 76800 95810 76810
rect 95940 76800 96060 76810
rect 96190 76800 96310 76810
rect 96440 76800 96560 76810
rect 96690 76800 96810 76810
rect 96940 76800 97060 76810
rect 97190 76800 97310 76810
rect 97440 76800 97560 76810
rect 97690 76800 97810 76810
rect 97940 76800 98060 76810
rect 98190 76800 98310 76810
rect 98440 76800 98560 76810
rect 98690 76800 98810 76810
rect 98940 76800 99060 76810
rect 99190 76800 99310 76810
rect 99440 76800 99560 76810
rect 99690 76800 99810 76810
rect 99940 76800 100060 76810
rect 100190 76800 100310 76810
rect 100440 76800 100560 76810
rect 100690 76800 100810 76810
rect 100940 76800 101060 76810
rect 101190 76800 101310 76810
rect 101440 76800 101560 76810
rect 101690 76800 101810 76810
rect 101940 76800 102060 76810
rect 102190 76800 102310 76810
rect 102440 76800 102560 76810
rect 102690 76800 102810 76810
rect 102940 76800 103060 76810
rect 103190 76800 103310 76810
rect 103440 76800 103560 76810
rect 103690 76800 103810 76810
rect 103940 76800 104060 76810
rect 104190 76800 104310 76810
rect 104440 76800 104560 76810
rect 104690 76800 104810 76810
rect 104940 76800 105060 76810
rect 105190 76800 105310 76810
rect 105440 76800 105560 76810
rect 105690 76800 105810 76810
rect 105940 76800 106060 76810
rect 106190 76800 106310 76810
rect 106440 76800 106560 76810
rect 106690 76800 106810 76810
rect 106940 76800 107060 76810
rect 107190 76800 107310 76810
rect 107440 76800 107560 76810
rect 107690 76800 107810 76810
rect 107940 76800 108060 76810
rect 108190 76800 108310 76810
rect 108440 76800 108560 76810
rect 108690 76800 108810 76810
rect 108940 76800 109060 76810
rect 109190 76800 109310 76810
rect 109440 76800 109560 76810
rect 109690 76800 109810 76810
rect 109940 76800 110060 76810
rect 110190 76800 110310 76810
rect 110440 76800 110560 76810
rect 110690 76800 110810 76810
rect 110940 76800 111060 76810
rect 111190 76800 111310 76810
rect 111440 76800 111560 76810
rect 111690 76800 111810 76810
rect 111940 76800 112060 76810
rect 112190 76800 112310 76810
rect 112440 76800 112560 76810
rect 112690 76800 112810 76810
rect 112940 76800 113060 76810
rect 113190 76800 113310 76810
rect 113440 76800 113560 76810
rect 113690 76800 113810 76810
rect 113940 76800 114060 76810
rect 114190 76800 114310 76810
rect 114440 76800 114560 76810
rect 114690 76800 114810 76810
rect 114940 76800 115060 76810
rect 115190 76800 115310 76810
rect 115440 76800 115560 76810
rect 115690 76800 115810 76810
rect 115940 76800 116000 76810
rect 89000 76700 116000 76800
rect 89000 76690 89060 76700
rect 89190 76690 89310 76700
rect 89440 76690 89560 76700
rect 89690 76690 89810 76700
rect 89940 76690 90060 76700
rect 90190 76690 90310 76700
rect 90440 76690 90560 76700
rect 90690 76690 90810 76700
rect 90940 76690 91060 76700
rect 91190 76690 91310 76700
rect 91440 76690 91560 76700
rect 91690 76690 91810 76700
rect 91940 76690 92060 76700
rect 92190 76690 92310 76700
rect 92440 76690 92560 76700
rect 92690 76690 92810 76700
rect 92940 76690 93060 76700
rect 93190 76690 93310 76700
rect 93440 76690 93560 76700
rect 93690 76690 93810 76700
rect 93940 76690 94060 76700
rect 94190 76690 94310 76700
rect 94440 76690 94560 76700
rect 94690 76690 94810 76700
rect 94940 76690 95060 76700
rect 95190 76690 95310 76700
rect 95440 76690 95560 76700
rect 95690 76690 95810 76700
rect 95940 76690 96060 76700
rect 96190 76690 96310 76700
rect 96440 76690 96560 76700
rect 96690 76690 96810 76700
rect 96940 76690 97060 76700
rect 97190 76690 97310 76700
rect 97440 76690 97560 76700
rect 97690 76690 97810 76700
rect 97940 76690 98060 76700
rect 98190 76690 98310 76700
rect 98440 76690 98560 76700
rect 98690 76690 98810 76700
rect 98940 76690 99060 76700
rect 99190 76690 99310 76700
rect 99440 76690 99560 76700
rect 99690 76690 99810 76700
rect 99940 76690 100060 76700
rect 100190 76690 100310 76700
rect 100440 76690 100560 76700
rect 100690 76690 100810 76700
rect 100940 76690 101060 76700
rect 101190 76690 101310 76700
rect 101440 76690 101560 76700
rect 101690 76690 101810 76700
rect 101940 76690 102060 76700
rect 102190 76690 102310 76700
rect 102440 76690 102560 76700
rect 102690 76690 102810 76700
rect 102940 76690 103060 76700
rect 103190 76690 103310 76700
rect 103440 76690 103560 76700
rect 103690 76690 103810 76700
rect 103940 76690 104060 76700
rect 104190 76690 104310 76700
rect 104440 76690 104560 76700
rect 104690 76690 104810 76700
rect 104940 76690 105060 76700
rect 105190 76690 105310 76700
rect 105440 76690 105560 76700
rect 105690 76690 105810 76700
rect 105940 76690 106060 76700
rect 106190 76690 106310 76700
rect 106440 76690 106560 76700
rect 106690 76690 106810 76700
rect 106940 76690 107060 76700
rect 107190 76690 107310 76700
rect 107440 76690 107560 76700
rect 107690 76690 107810 76700
rect 107940 76690 108060 76700
rect 108190 76690 108310 76700
rect 108440 76690 108560 76700
rect 108690 76690 108810 76700
rect 108940 76690 109060 76700
rect 109190 76690 109310 76700
rect 109440 76690 109560 76700
rect 109690 76690 109810 76700
rect 109940 76690 110060 76700
rect 110190 76690 110310 76700
rect 110440 76690 110560 76700
rect 110690 76690 110810 76700
rect 110940 76690 111060 76700
rect 111190 76690 111310 76700
rect 111440 76690 111560 76700
rect 111690 76690 111810 76700
rect 111940 76690 112060 76700
rect 112190 76690 112310 76700
rect 112440 76690 112560 76700
rect 112690 76690 112810 76700
rect 112940 76690 113060 76700
rect 113190 76690 113310 76700
rect 113440 76690 113560 76700
rect 113690 76690 113810 76700
rect 113940 76690 114060 76700
rect 114190 76690 114310 76700
rect 114440 76690 114560 76700
rect 114690 76690 114810 76700
rect 114940 76690 115060 76700
rect 115190 76690 115310 76700
rect 115440 76690 115560 76700
rect 115690 76690 115810 76700
rect 115940 76690 116000 76700
rect 89000 76560 89050 76690
rect 89200 76560 89300 76690
rect 89450 76560 89550 76690
rect 89700 76560 89800 76690
rect 89950 76560 90050 76690
rect 90200 76560 90300 76690
rect 90450 76560 90550 76690
rect 90700 76560 90800 76690
rect 90950 76560 91050 76690
rect 91200 76560 91300 76690
rect 91450 76560 91550 76690
rect 91700 76560 91800 76690
rect 91950 76560 92050 76690
rect 92200 76560 92300 76690
rect 92450 76560 92550 76690
rect 92700 76560 92800 76690
rect 92950 76560 93050 76690
rect 93200 76560 93300 76690
rect 93450 76560 93550 76690
rect 93700 76560 93800 76690
rect 93950 76560 94050 76690
rect 94200 76560 94300 76690
rect 94450 76560 94550 76690
rect 94700 76560 94800 76690
rect 94950 76560 95050 76690
rect 95200 76560 95300 76690
rect 95450 76560 95550 76690
rect 95700 76560 95800 76690
rect 95950 76560 96050 76690
rect 96200 76560 96300 76690
rect 96450 76560 96550 76690
rect 96700 76560 96800 76690
rect 96950 76560 97050 76690
rect 97200 76560 97300 76690
rect 97450 76560 97550 76690
rect 97700 76560 97800 76690
rect 97950 76560 98050 76690
rect 98200 76560 98300 76690
rect 98450 76560 98550 76690
rect 98700 76560 98800 76690
rect 98950 76560 99050 76690
rect 99200 76560 99300 76690
rect 99450 76560 99550 76690
rect 99700 76560 99800 76690
rect 99950 76560 100050 76690
rect 100200 76560 100300 76690
rect 100450 76560 100550 76690
rect 100700 76560 100800 76690
rect 100950 76560 101050 76690
rect 101200 76560 101300 76690
rect 101450 76560 101550 76690
rect 101700 76560 101800 76690
rect 101950 76560 102050 76690
rect 102200 76560 102300 76690
rect 102450 76560 102550 76690
rect 102700 76560 102800 76690
rect 102950 76560 103050 76690
rect 103200 76560 103300 76690
rect 103450 76560 103550 76690
rect 103700 76560 103800 76690
rect 103950 76560 104050 76690
rect 104200 76560 104300 76690
rect 104450 76560 104550 76690
rect 104700 76560 104800 76690
rect 104950 76560 105050 76690
rect 105200 76560 105300 76690
rect 105450 76560 105550 76690
rect 105700 76560 105800 76690
rect 105950 76560 106050 76690
rect 106200 76560 106300 76690
rect 106450 76560 106550 76690
rect 106700 76560 106800 76690
rect 106950 76560 107050 76690
rect 107200 76560 107300 76690
rect 107450 76560 107550 76690
rect 107700 76560 107800 76690
rect 107950 76560 108050 76690
rect 108200 76560 108300 76690
rect 108450 76560 108550 76690
rect 108700 76560 108800 76690
rect 108950 76560 109050 76690
rect 109200 76560 109300 76690
rect 109450 76560 109550 76690
rect 109700 76560 109800 76690
rect 109950 76560 110050 76690
rect 110200 76560 110300 76690
rect 110450 76560 110550 76690
rect 110700 76560 110800 76690
rect 110950 76560 111050 76690
rect 111200 76560 111300 76690
rect 111450 76560 111550 76690
rect 111700 76560 111800 76690
rect 111950 76560 112050 76690
rect 112200 76560 112300 76690
rect 112450 76560 112550 76690
rect 112700 76560 112800 76690
rect 112950 76560 113050 76690
rect 113200 76560 113300 76690
rect 113450 76560 113550 76690
rect 113700 76560 113800 76690
rect 113950 76560 114050 76690
rect 114200 76560 114300 76690
rect 114450 76560 114550 76690
rect 114700 76560 114800 76690
rect 114950 76560 115050 76690
rect 115200 76560 115300 76690
rect 115450 76560 115550 76690
rect 115700 76560 115800 76690
rect 115950 76560 116000 76690
rect 89000 76550 89060 76560
rect 89190 76550 89310 76560
rect 89440 76550 89560 76560
rect 89690 76550 89810 76560
rect 89940 76550 90060 76560
rect 90190 76550 90310 76560
rect 90440 76550 90560 76560
rect 90690 76550 90810 76560
rect 90940 76550 91060 76560
rect 91190 76550 91310 76560
rect 91440 76550 91560 76560
rect 91690 76550 91810 76560
rect 91940 76550 92060 76560
rect 92190 76550 92310 76560
rect 92440 76550 92560 76560
rect 92690 76550 92810 76560
rect 92940 76550 93060 76560
rect 93190 76550 93310 76560
rect 93440 76550 93560 76560
rect 93690 76550 93810 76560
rect 93940 76550 94060 76560
rect 94190 76550 94310 76560
rect 94440 76550 94560 76560
rect 94690 76550 94810 76560
rect 94940 76550 95060 76560
rect 95190 76550 95310 76560
rect 95440 76550 95560 76560
rect 95690 76550 95810 76560
rect 95940 76550 96060 76560
rect 96190 76550 96310 76560
rect 96440 76550 96560 76560
rect 96690 76550 96810 76560
rect 96940 76550 97060 76560
rect 97190 76550 97310 76560
rect 97440 76550 97560 76560
rect 97690 76550 97810 76560
rect 97940 76550 98060 76560
rect 98190 76550 98310 76560
rect 98440 76550 98560 76560
rect 98690 76550 98810 76560
rect 98940 76550 99060 76560
rect 99190 76550 99310 76560
rect 99440 76550 99560 76560
rect 99690 76550 99810 76560
rect 99940 76550 100060 76560
rect 100190 76550 100310 76560
rect 100440 76550 100560 76560
rect 100690 76550 100810 76560
rect 100940 76550 101060 76560
rect 101190 76550 101310 76560
rect 101440 76550 101560 76560
rect 101690 76550 101810 76560
rect 101940 76550 102060 76560
rect 102190 76550 102310 76560
rect 102440 76550 102560 76560
rect 102690 76550 102810 76560
rect 102940 76550 103060 76560
rect 103190 76550 103310 76560
rect 103440 76550 103560 76560
rect 103690 76550 103810 76560
rect 103940 76550 104060 76560
rect 104190 76550 104310 76560
rect 104440 76550 104560 76560
rect 104690 76550 104810 76560
rect 104940 76550 105060 76560
rect 105190 76550 105310 76560
rect 105440 76550 105560 76560
rect 105690 76550 105810 76560
rect 105940 76550 106060 76560
rect 106190 76550 106310 76560
rect 106440 76550 106560 76560
rect 106690 76550 106810 76560
rect 106940 76550 107060 76560
rect 107190 76550 107310 76560
rect 107440 76550 107560 76560
rect 107690 76550 107810 76560
rect 107940 76550 108060 76560
rect 108190 76550 108310 76560
rect 108440 76550 108560 76560
rect 108690 76550 108810 76560
rect 108940 76550 109060 76560
rect 109190 76550 109310 76560
rect 109440 76550 109560 76560
rect 109690 76550 109810 76560
rect 109940 76550 110060 76560
rect 110190 76550 110310 76560
rect 110440 76550 110560 76560
rect 110690 76550 110810 76560
rect 110940 76550 111060 76560
rect 111190 76550 111310 76560
rect 111440 76550 111560 76560
rect 111690 76550 111810 76560
rect 111940 76550 112060 76560
rect 112190 76550 112310 76560
rect 112440 76550 112560 76560
rect 112690 76550 112810 76560
rect 112940 76550 113060 76560
rect 113190 76550 113310 76560
rect 113440 76550 113560 76560
rect 113690 76550 113810 76560
rect 113940 76550 114060 76560
rect 114190 76550 114310 76560
rect 114440 76550 114560 76560
rect 114690 76550 114810 76560
rect 114940 76550 115060 76560
rect 115190 76550 115310 76560
rect 115440 76550 115560 76560
rect 115690 76550 115810 76560
rect 115940 76550 116000 76560
rect 89000 76450 116000 76550
rect 89000 76440 89060 76450
rect 89190 76440 89310 76450
rect 89440 76440 89560 76450
rect 89690 76440 89810 76450
rect 89940 76440 90060 76450
rect 90190 76440 90310 76450
rect 90440 76440 90560 76450
rect 90690 76440 90810 76450
rect 90940 76440 91060 76450
rect 91190 76440 91310 76450
rect 91440 76440 91560 76450
rect 91690 76440 91810 76450
rect 91940 76440 92060 76450
rect 92190 76440 92310 76450
rect 92440 76440 92560 76450
rect 92690 76440 92810 76450
rect 92940 76440 93060 76450
rect 93190 76440 93310 76450
rect 93440 76440 93560 76450
rect 93690 76440 93810 76450
rect 93940 76440 94060 76450
rect 94190 76440 94310 76450
rect 94440 76440 94560 76450
rect 94690 76440 94810 76450
rect 94940 76440 95060 76450
rect 95190 76440 95310 76450
rect 95440 76440 95560 76450
rect 95690 76440 95810 76450
rect 95940 76440 96060 76450
rect 96190 76440 96310 76450
rect 96440 76440 96560 76450
rect 96690 76440 96810 76450
rect 96940 76440 97060 76450
rect 97190 76440 97310 76450
rect 97440 76440 97560 76450
rect 97690 76440 97810 76450
rect 97940 76440 98060 76450
rect 98190 76440 98310 76450
rect 98440 76440 98560 76450
rect 98690 76440 98810 76450
rect 98940 76440 99060 76450
rect 99190 76440 99310 76450
rect 99440 76440 99560 76450
rect 99690 76440 99810 76450
rect 99940 76440 100060 76450
rect 100190 76440 100310 76450
rect 100440 76440 100560 76450
rect 100690 76440 100810 76450
rect 100940 76440 101060 76450
rect 101190 76440 101310 76450
rect 101440 76440 101560 76450
rect 101690 76440 101810 76450
rect 101940 76440 102060 76450
rect 102190 76440 102310 76450
rect 102440 76440 102560 76450
rect 102690 76440 102810 76450
rect 102940 76440 103060 76450
rect 103190 76440 103310 76450
rect 103440 76440 103560 76450
rect 103690 76440 103810 76450
rect 103940 76440 104060 76450
rect 104190 76440 104310 76450
rect 104440 76440 104560 76450
rect 104690 76440 104810 76450
rect 104940 76440 105060 76450
rect 105190 76440 105310 76450
rect 105440 76440 105560 76450
rect 105690 76440 105810 76450
rect 105940 76440 106060 76450
rect 106190 76440 106310 76450
rect 106440 76440 106560 76450
rect 106690 76440 106810 76450
rect 106940 76440 107060 76450
rect 107190 76440 107310 76450
rect 107440 76440 107560 76450
rect 107690 76440 107810 76450
rect 107940 76440 108060 76450
rect 108190 76440 108310 76450
rect 108440 76440 108560 76450
rect 108690 76440 108810 76450
rect 108940 76440 109060 76450
rect 109190 76440 109310 76450
rect 109440 76440 109560 76450
rect 109690 76440 109810 76450
rect 109940 76440 110060 76450
rect 110190 76440 110310 76450
rect 110440 76440 110560 76450
rect 110690 76440 110810 76450
rect 110940 76440 111060 76450
rect 111190 76440 111310 76450
rect 111440 76440 111560 76450
rect 111690 76440 111810 76450
rect 111940 76440 112060 76450
rect 112190 76440 112310 76450
rect 112440 76440 112560 76450
rect 112690 76440 112810 76450
rect 112940 76440 113060 76450
rect 113190 76440 113310 76450
rect 113440 76440 113560 76450
rect 113690 76440 113810 76450
rect 113940 76440 114060 76450
rect 114190 76440 114310 76450
rect 114440 76440 114560 76450
rect 114690 76440 114810 76450
rect 114940 76440 115060 76450
rect 115190 76440 115310 76450
rect 115440 76440 115560 76450
rect 115690 76440 115810 76450
rect 115940 76440 116000 76450
rect 89000 76310 89050 76440
rect 89200 76310 89300 76440
rect 89450 76310 89550 76440
rect 89700 76310 89800 76440
rect 89950 76310 90050 76440
rect 90200 76310 90300 76440
rect 90450 76310 90550 76440
rect 90700 76310 90800 76440
rect 90950 76310 91050 76440
rect 91200 76310 91300 76440
rect 91450 76310 91550 76440
rect 91700 76310 91800 76440
rect 91950 76310 92050 76440
rect 92200 76310 92300 76440
rect 92450 76310 92550 76440
rect 92700 76310 92800 76440
rect 92950 76310 93050 76440
rect 93200 76310 93300 76440
rect 93450 76310 93550 76440
rect 93700 76310 93800 76440
rect 93950 76310 94050 76440
rect 94200 76310 94300 76440
rect 94450 76310 94550 76440
rect 94700 76310 94800 76440
rect 94950 76310 95050 76440
rect 95200 76310 95300 76440
rect 95450 76310 95550 76440
rect 95700 76310 95800 76440
rect 95950 76310 96050 76440
rect 96200 76310 96300 76440
rect 96450 76310 96550 76440
rect 96700 76310 96800 76440
rect 96950 76310 97050 76440
rect 97200 76310 97300 76440
rect 97450 76310 97550 76440
rect 97700 76310 97800 76440
rect 97950 76310 98050 76440
rect 98200 76310 98300 76440
rect 98450 76310 98550 76440
rect 98700 76310 98800 76440
rect 98950 76310 99050 76440
rect 99200 76310 99300 76440
rect 99450 76310 99550 76440
rect 99700 76310 99800 76440
rect 99950 76310 100050 76440
rect 100200 76310 100300 76440
rect 100450 76310 100550 76440
rect 100700 76310 100800 76440
rect 100950 76310 101050 76440
rect 101200 76310 101300 76440
rect 101450 76310 101550 76440
rect 101700 76310 101800 76440
rect 101950 76310 102050 76440
rect 102200 76310 102300 76440
rect 102450 76310 102550 76440
rect 102700 76310 102800 76440
rect 102950 76310 103050 76440
rect 103200 76310 103300 76440
rect 103450 76310 103550 76440
rect 103700 76310 103800 76440
rect 103950 76310 104050 76440
rect 104200 76310 104300 76440
rect 104450 76310 104550 76440
rect 104700 76310 104800 76440
rect 104950 76310 105050 76440
rect 105200 76310 105300 76440
rect 105450 76310 105550 76440
rect 105700 76310 105800 76440
rect 105950 76310 106050 76440
rect 106200 76310 106300 76440
rect 106450 76310 106550 76440
rect 106700 76310 106800 76440
rect 106950 76310 107050 76440
rect 107200 76310 107300 76440
rect 107450 76310 107550 76440
rect 107700 76310 107800 76440
rect 107950 76310 108050 76440
rect 108200 76310 108300 76440
rect 108450 76310 108550 76440
rect 108700 76310 108800 76440
rect 108950 76310 109050 76440
rect 109200 76310 109300 76440
rect 109450 76310 109550 76440
rect 109700 76310 109800 76440
rect 109950 76310 110050 76440
rect 110200 76310 110300 76440
rect 110450 76310 110550 76440
rect 110700 76310 110800 76440
rect 110950 76310 111050 76440
rect 111200 76310 111300 76440
rect 111450 76310 111550 76440
rect 111700 76310 111800 76440
rect 111950 76310 112050 76440
rect 112200 76310 112300 76440
rect 112450 76310 112550 76440
rect 112700 76310 112800 76440
rect 112950 76310 113050 76440
rect 113200 76310 113300 76440
rect 113450 76310 113550 76440
rect 113700 76310 113800 76440
rect 113950 76310 114050 76440
rect 114200 76310 114300 76440
rect 114450 76310 114550 76440
rect 114700 76310 114800 76440
rect 114950 76310 115050 76440
rect 115200 76310 115300 76440
rect 115450 76310 115550 76440
rect 115700 76310 115800 76440
rect 115950 76310 116000 76440
rect 89000 76300 89060 76310
rect 89190 76300 89310 76310
rect 89440 76300 89560 76310
rect 89690 76300 89810 76310
rect 89940 76300 90060 76310
rect 90190 76300 90310 76310
rect 90440 76300 90560 76310
rect 90690 76300 90810 76310
rect 90940 76300 91060 76310
rect 91190 76300 91310 76310
rect 91440 76300 91560 76310
rect 91690 76300 91810 76310
rect 91940 76300 92060 76310
rect 92190 76300 92310 76310
rect 92440 76300 92560 76310
rect 92690 76300 92810 76310
rect 92940 76300 93060 76310
rect 93190 76300 93310 76310
rect 93440 76300 93560 76310
rect 93690 76300 93810 76310
rect 93940 76300 94060 76310
rect 94190 76300 94310 76310
rect 94440 76300 94560 76310
rect 94690 76300 94810 76310
rect 94940 76300 95060 76310
rect 95190 76300 95310 76310
rect 95440 76300 95560 76310
rect 95690 76300 95810 76310
rect 95940 76300 96060 76310
rect 96190 76300 96310 76310
rect 96440 76300 96560 76310
rect 96690 76300 96810 76310
rect 96940 76300 97060 76310
rect 97190 76300 97310 76310
rect 97440 76300 97560 76310
rect 97690 76300 97810 76310
rect 97940 76300 98060 76310
rect 98190 76300 98310 76310
rect 98440 76300 98560 76310
rect 98690 76300 98810 76310
rect 98940 76300 99060 76310
rect 99190 76300 99310 76310
rect 99440 76300 99560 76310
rect 99690 76300 99810 76310
rect 99940 76300 100060 76310
rect 100190 76300 100310 76310
rect 100440 76300 100560 76310
rect 100690 76300 100810 76310
rect 100940 76300 101060 76310
rect 101190 76300 101310 76310
rect 101440 76300 101560 76310
rect 101690 76300 101810 76310
rect 101940 76300 102060 76310
rect 102190 76300 102310 76310
rect 102440 76300 102560 76310
rect 102690 76300 102810 76310
rect 102940 76300 103060 76310
rect 103190 76300 103310 76310
rect 103440 76300 103560 76310
rect 103690 76300 103810 76310
rect 103940 76300 104060 76310
rect 104190 76300 104310 76310
rect 104440 76300 104560 76310
rect 104690 76300 104810 76310
rect 104940 76300 105060 76310
rect 105190 76300 105310 76310
rect 105440 76300 105560 76310
rect 105690 76300 105810 76310
rect 105940 76300 106060 76310
rect 106190 76300 106310 76310
rect 106440 76300 106560 76310
rect 106690 76300 106810 76310
rect 106940 76300 107060 76310
rect 107190 76300 107310 76310
rect 107440 76300 107560 76310
rect 107690 76300 107810 76310
rect 107940 76300 108060 76310
rect 108190 76300 108310 76310
rect 108440 76300 108560 76310
rect 108690 76300 108810 76310
rect 108940 76300 109060 76310
rect 109190 76300 109310 76310
rect 109440 76300 109560 76310
rect 109690 76300 109810 76310
rect 109940 76300 110060 76310
rect 110190 76300 110310 76310
rect 110440 76300 110560 76310
rect 110690 76300 110810 76310
rect 110940 76300 111060 76310
rect 111190 76300 111310 76310
rect 111440 76300 111560 76310
rect 111690 76300 111810 76310
rect 111940 76300 112060 76310
rect 112190 76300 112310 76310
rect 112440 76300 112560 76310
rect 112690 76300 112810 76310
rect 112940 76300 113060 76310
rect 113190 76300 113310 76310
rect 113440 76300 113560 76310
rect 113690 76300 113810 76310
rect 113940 76300 114060 76310
rect 114190 76300 114310 76310
rect 114440 76300 114560 76310
rect 114690 76300 114810 76310
rect 114940 76300 115060 76310
rect 115190 76300 115310 76310
rect 115440 76300 115560 76310
rect 115690 76300 115810 76310
rect 115940 76300 116000 76310
rect 89000 76200 116000 76300
rect 89000 76190 89060 76200
rect 89190 76190 89310 76200
rect 89440 76190 89560 76200
rect 89690 76190 89810 76200
rect 89940 76190 90060 76200
rect 90190 76190 90310 76200
rect 90440 76190 90560 76200
rect 90690 76190 90810 76200
rect 90940 76190 91060 76200
rect 91190 76190 91310 76200
rect 91440 76190 91560 76200
rect 91690 76190 91810 76200
rect 91940 76190 92060 76200
rect 92190 76190 92310 76200
rect 92440 76190 92560 76200
rect 92690 76190 92810 76200
rect 92940 76190 93060 76200
rect 93190 76190 93310 76200
rect 93440 76190 93560 76200
rect 93690 76190 93810 76200
rect 93940 76190 94060 76200
rect 94190 76190 94310 76200
rect 94440 76190 94560 76200
rect 94690 76190 94810 76200
rect 94940 76190 95060 76200
rect 95190 76190 95310 76200
rect 95440 76190 95560 76200
rect 95690 76190 95810 76200
rect 95940 76190 96060 76200
rect 96190 76190 96310 76200
rect 96440 76190 96560 76200
rect 96690 76190 96810 76200
rect 96940 76190 97060 76200
rect 97190 76190 97310 76200
rect 97440 76190 97560 76200
rect 97690 76190 97810 76200
rect 97940 76190 98060 76200
rect 98190 76190 98310 76200
rect 98440 76190 98560 76200
rect 98690 76190 98810 76200
rect 98940 76190 99060 76200
rect 99190 76190 99310 76200
rect 99440 76190 99560 76200
rect 99690 76190 99810 76200
rect 99940 76190 100060 76200
rect 100190 76190 100310 76200
rect 100440 76190 100560 76200
rect 100690 76190 100810 76200
rect 100940 76190 101060 76200
rect 101190 76190 101310 76200
rect 101440 76190 101560 76200
rect 101690 76190 101810 76200
rect 101940 76190 102060 76200
rect 102190 76190 102310 76200
rect 102440 76190 102560 76200
rect 102690 76190 102810 76200
rect 102940 76190 103060 76200
rect 103190 76190 103310 76200
rect 103440 76190 103560 76200
rect 103690 76190 103810 76200
rect 103940 76190 104060 76200
rect 104190 76190 104310 76200
rect 104440 76190 104560 76200
rect 104690 76190 104810 76200
rect 104940 76190 105060 76200
rect 105190 76190 105310 76200
rect 105440 76190 105560 76200
rect 105690 76190 105810 76200
rect 105940 76190 106060 76200
rect 106190 76190 106310 76200
rect 106440 76190 106560 76200
rect 106690 76190 106810 76200
rect 106940 76190 107060 76200
rect 107190 76190 107310 76200
rect 107440 76190 107560 76200
rect 107690 76190 107810 76200
rect 107940 76190 108060 76200
rect 108190 76190 108310 76200
rect 108440 76190 108560 76200
rect 108690 76190 108810 76200
rect 108940 76190 109060 76200
rect 109190 76190 109310 76200
rect 109440 76190 109560 76200
rect 109690 76190 109810 76200
rect 109940 76190 110060 76200
rect 110190 76190 110310 76200
rect 110440 76190 110560 76200
rect 110690 76190 110810 76200
rect 110940 76190 111060 76200
rect 111190 76190 111310 76200
rect 111440 76190 111560 76200
rect 111690 76190 111810 76200
rect 111940 76190 112060 76200
rect 112190 76190 112310 76200
rect 112440 76190 112560 76200
rect 112690 76190 112810 76200
rect 112940 76190 113060 76200
rect 113190 76190 113310 76200
rect 113440 76190 113560 76200
rect 113690 76190 113810 76200
rect 113940 76190 114060 76200
rect 114190 76190 114310 76200
rect 114440 76190 114560 76200
rect 114690 76190 114810 76200
rect 114940 76190 115060 76200
rect 115190 76190 115310 76200
rect 115440 76190 115560 76200
rect 115690 76190 115810 76200
rect 115940 76190 116000 76200
rect 89000 76060 89050 76190
rect 89200 76060 89300 76190
rect 89450 76060 89550 76190
rect 89700 76060 89800 76190
rect 89950 76060 90050 76190
rect 90200 76060 90300 76190
rect 90450 76060 90550 76190
rect 90700 76060 90800 76190
rect 90950 76060 91050 76190
rect 91200 76060 91300 76190
rect 91450 76060 91550 76190
rect 91700 76060 91800 76190
rect 91950 76060 92050 76190
rect 92200 76060 92300 76190
rect 92450 76060 92550 76190
rect 92700 76060 92800 76190
rect 92950 76060 93050 76190
rect 93200 76060 93300 76190
rect 93450 76060 93550 76190
rect 93700 76060 93800 76190
rect 93950 76060 94050 76190
rect 94200 76060 94300 76190
rect 94450 76060 94550 76190
rect 94700 76060 94800 76190
rect 94950 76060 95050 76190
rect 95200 76060 95300 76190
rect 95450 76060 95550 76190
rect 95700 76060 95800 76190
rect 95950 76060 96050 76190
rect 96200 76060 96300 76190
rect 96450 76060 96550 76190
rect 96700 76060 96800 76190
rect 96950 76060 97050 76190
rect 97200 76060 97300 76190
rect 97450 76060 97550 76190
rect 97700 76060 97800 76190
rect 97950 76060 98050 76190
rect 98200 76060 98300 76190
rect 98450 76060 98550 76190
rect 98700 76060 98800 76190
rect 98950 76060 99050 76190
rect 99200 76060 99300 76190
rect 99450 76060 99550 76190
rect 99700 76060 99800 76190
rect 99950 76060 100050 76190
rect 100200 76060 100300 76190
rect 100450 76060 100550 76190
rect 100700 76060 100800 76190
rect 100950 76060 101050 76190
rect 101200 76060 101300 76190
rect 101450 76060 101550 76190
rect 101700 76060 101800 76190
rect 101950 76060 102050 76190
rect 102200 76060 102300 76190
rect 102450 76060 102550 76190
rect 102700 76060 102800 76190
rect 102950 76060 103050 76190
rect 103200 76060 103300 76190
rect 103450 76060 103550 76190
rect 103700 76060 103800 76190
rect 103950 76060 104050 76190
rect 104200 76060 104300 76190
rect 104450 76060 104550 76190
rect 104700 76060 104800 76190
rect 104950 76060 105050 76190
rect 105200 76060 105300 76190
rect 105450 76060 105550 76190
rect 105700 76060 105800 76190
rect 105950 76060 106050 76190
rect 106200 76060 106300 76190
rect 106450 76060 106550 76190
rect 106700 76060 106800 76190
rect 106950 76060 107050 76190
rect 107200 76060 107300 76190
rect 107450 76060 107550 76190
rect 107700 76060 107800 76190
rect 107950 76060 108050 76190
rect 108200 76060 108300 76190
rect 108450 76060 108550 76190
rect 108700 76060 108800 76190
rect 108950 76060 109050 76190
rect 109200 76060 109300 76190
rect 109450 76060 109550 76190
rect 109700 76060 109800 76190
rect 109950 76060 110050 76190
rect 110200 76060 110300 76190
rect 110450 76060 110550 76190
rect 110700 76060 110800 76190
rect 110950 76060 111050 76190
rect 111200 76060 111300 76190
rect 111450 76060 111550 76190
rect 111700 76060 111800 76190
rect 111950 76060 112050 76190
rect 112200 76060 112300 76190
rect 112450 76060 112550 76190
rect 112700 76060 112800 76190
rect 112950 76060 113050 76190
rect 113200 76060 113300 76190
rect 113450 76060 113550 76190
rect 113700 76060 113800 76190
rect 113950 76060 114050 76190
rect 114200 76060 114300 76190
rect 114450 76060 114550 76190
rect 114700 76060 114800 76190
rect 114950 76060 115050 76190
rect 115200 76060 115300 76190
rect 115450 76060 115550 76190
rect 115700 76060 115800 76190
rect 115950 76060 116000 76190
rect 89000 76050 89060 76060
rect 89190 76050 89310 76060
rect 89440 76050 89560 76060
rect 89690 76050 89810 76060
rect 89940 76050 90060 76060
rect 90190 76050 90310 76060
rect 90440 76050 90560 76060
rect 90690 76050 90810 76060
rect 90940 76050 91060 76060
rect 91190 76050 91310 76060
rect 91440 76050 91560 76060
rect 91690 76050 91810 76060
rect 91940 76050 92060 76060
rect 92190 76050 92310 76060
rect 92440 76050 92560 76060
rect 92690 76050 92810 76060
rect 92940 76050 93060 76060
rect 93190 76050 93310 76060
rect 93440 76050 93560 76060
rect 93690 76050 93810 76060
rect 93940 76050 94060 76060
rect 94190 76050 94310 76060
rect 94440 76050 94560 76060
rect 94690 76050 94810 76060
rect 94940 76050 95060 76060
rect 95190 76050 95310 76060
rect 95440 76050 95560 76060
rect 95690 76050 95810 76060
rect 95940 76050 96060 76060
rect 96190 76050 96310 76060
rect 96440 76050 96560 76060
rect 96690 76050 96810 76060
rect 96940 76050 97060 76060
rect 97190 76050 97310 76060
rect 97440 76050 97560 76060
rect 97690 76050 97810 76060
rect 97940 76050 98060 76060
rect 98190 76050 98310 76060
rect 98440 76050 98560 76060
rect 98690 76050 98810 76060
rect 98940 76050 99060 76060
rect 99190 76050 99310 76060
rect 99440 76050 99560 76060
rect 99690 76050 99810 76060
rect 99940 76050 100060 76060
rect 100190 76050 100310 76060
rect 100440 76050 100560 76060
rect 100690 76050 100810 76060
rect 100940 76050 101060 76060
rect 101190 76050 101310 76060
rect 101440 76050 101560 76060
rect 101690 76050 101810 76060
rect 101940 76050 102060 76060
rect 102190 76050 102310 76060
rect 102440 76050 102560 76060
rect 102690 76050 102810 76060
rect 102940 76050 103060 76060
rect 103190 76050 103310 76060
rect 103440 76050 103560 76060
rect 103690 76050 103810 76060
rect 103940 76050 104060 76060
rect 104190 76050 104310 76060
rect 104440 76050 104560 76060
rect 104690 76050 104810 76060
rect 104940 76050 105060 76060
rect 105190 76050 105310 76060
rect 105440 76050 105560 76060
rect 105690 76050 105810 76060
rect 105940 76050 106060 76060
rect 106190 76050 106310 76060
rect 106440 76050 106560 76060
rect 106690 76050 106810 76060
rect 106940 76050 107060 76060
rect 107190 76050 107310 76060
rect 107440 76050 107560 76060
rect 107690 76050 107810 76060
rect 107940 76050 108060 76060
rect 108190 76050 108310 76060
rect 108440 76050 108560 76060
rect 108690 76050 108810 76060
rect 108940 76050 109060 76060
rect 109190 76050 109310 76060
rect 109440 76050 109560 76060
rect 109690 76050 109810 76060
rect 109940 76050 110060 76060
rect 110190 76050 110310 76060
rect 110440 76050 110560 76060
rect 110690 76050 110810 76060
rect 110940 76050 111060 76060
rect 111190 76050 111310 76060
rect 111440 76050 111560 76060
rect 111690 76050 111810 76060
rect 111940 76050 112060 76060
rect 112190 76050 112310 76060
rect 112440 76050 112560 76060
rect 112690 76050 112810 76060
rect 112940 76050 113060 76060
rect 113190 76050 113310 76060
rect 113440 76050 113560 76060
rect 113690 76050 113810 76060
rect 113940 76050 114060 76060
rect 114190 76050 114310 76060
rect 114440 76050 114560 76060
rect 114690 76050 114810 76060
rect 114940 76050 115060 76060
rect 115190 76050 115310 76060
rect 115440 76050 115560 76060
rect 115690 76050 115810 76060
rect 115940 76050 116000 76060
rect 89000 75950 116000 76050
rect 89000 75940 89060 75950
rect 89190 75940 89310 75950
rect 89440 75940 89560 75950
rect 89690 75940 89810 75950
rect 89940 75940 90060 75950
rect 90190 75940 90310 75950
rect 90440 75940 90560 75950
rect 90690 75940 90810 75950
rect 90940 75940 91060 75950
rect 91190 75940 91310 75950
rect 91440 75940 91560 75950
rect 91690 75940 91810 75950
rect 91940 75940 92060 75950
rect 92190 75940 92310 75950
rect 92440 75940 92560 75950
rect 92690 75940 92810 75950
rect 92940 75940 93060 75950
rect 93190 75940 93310 75950
rect 93440 75940 93560 75950
rect 93690 75940 93810 75950
rect 93940 75940 94060 75950
rect 94190 75940 94310 75950
rect 94440 75940 94560 75950
rect 94690 75940 94810 75950
rect 94940 75940 95060 75950
rect 95190 75940 95310 75950
rect 95440 75940 95560 75950
rect 95690 75940 95810 75950
rect 95940 75940 96060 75950
rect 96190 75940 96310 75950
rect 96440 75940 96560 75950
rect 96690 75940 96810 75950
rect 96940 75940 97060 75950
rect 97190 75940 97310 75950
rect 97440 75940 97560 75950
rect 97690 75940 97810 75950
rect 97940 75940 98060 75950
rect 98190 75940 98310 75950
rect 98440 75940 98560 75950
rect 98690 75940 98810 75950
rect 98940 75940 99060 75950
rect 99190 75940 99310 75950
rect 99440 75940 99560 75950
rect 99690 75940 99810 75950
rect 99940 75940 100060 75950
rect 100190 75940 100310 75950
rect 100440 75940 100560 75950
rect 100690 75940 100810 75950
rect 100940 75940 101060 75950
rect 101190 75940 101310 75950
rect 101440 75940 101560 75950
rect 101690 75940 101810 75950
rect 101940 75940 102060 75950
rect 102190 75940 102310 75950
rect 102440 75940 102560 75950
rect 102690 75940 102810 75950
rect 102940 75940 103060 75950
rect 103190 75940 103310 75950
rect 103440 75940 103560 75950
rect 103690 75940 103810 75950
rect 103940 75940 104060 75950
rect 104190 75940 104310 75950
rect 104440 75940 104560 75950
rect 104690 75940 104810 75950
rect 104940 75940 105060 75950
rect 105190 75940 105310 75950
rect 105440 75940 105560 75950
rect 105690 75940 105810 75950
rect 105940 75940 106060 75950
rect 106190 75940 106310 75950
rect 106440 75940 106560 75950
rect 106690 75940 106810 75950
rect 106940 75940 107060 75950
rect 107190 75940 107310 75950
rect 107440 75940 107560 75950
rect 107690 75940 107810 75950
rect 107940 75940 108060 75950
rect 108190 75940 108310 75950
rect 108440 75940 108560 75950
rect 108690 75940 108810 75950
rect 108940 75940 109060 75950
rect 109190 75940 109310 75950
rect 109440 75940 109560 75950
rect 109690 75940 109810 75950
rect 109940 75940 110060 75950
rect 110190 75940 110310 75950
rect 110440 75940 110560 75950
rect 110690 75940 110810 75950
rect 110940 75940 111060 75950
rect 111190 75940 111310 75950
rect 111440 75940 111560 75950
rect 111690 75940 111810 75950
rect 111940 75940 112060 75950
rect 112190 75940 112310 75950
rect 112440 75940 112560 75950
rect 112690 75940 112810 75950
rect 112940 75940 113060 75950
rect 113190 75940 113310 75950
rect 113440 75940 113560 75950
rect 113690 75940 113810 75950
rect 113940 75940 114060 75950
rect 114190 75940 114310 75950
rect 114440 75940 114560 75950
rect 114690 75940 114810 75950
rect 114940 75940 115060 75950
rect 115190 75940 115310 75950
rect 115440 75940 115560 75950
rect 115690 75940 115810 75950
rect 115940 75940 116000 75950
rect 89000 75810 89050 75940
rect 89200 75810 89300 75940
rect 89450 75810 89550 75940
rect 89700 75810 89800 75940
rect 89950 75810 90050 75940
rect 90200 75810 90300 75940
rect 90450 75810 90550 75940
rect 90700 75810 90800 75940
rect 90950 75810 91050 75940
rect 91200 75810 91300 75940
rect 91450 75810 91550 75940
rect 91700 75810 91800 75940
rect 91950 75810 92050 75940
rect 92200 75810 92300 75940
rect 92450 75810 92550 75940
rect 92700 75810 92800 75940
rect 92950 75810 93050 75940
rect 93200 75810 93300 75940
rect 93450 75810 93550 75940
rect 93700 75810 93800 75940
rect 93950 75810 94050 75940
rect 94200 75810 94300 75940
rect 94450 75810 94550 75940
rect 94700 75810 94800 75940
rect 94950 75810 95050 75940
rect 95200 75810 95300 75940
rect 95450 75810 95550 75940
rect 95700 75810 95800 75940
rect 95950 75810 96050 75940
rect 96200 75810 96300 75940
rect 96450 75810 96550 75940
rect 96700 75810 96800 75940
rect 96950 75810 97050 75940
rect 97200 75810 97300 75940
rect 97450 75810 97550 75940
rect 97700 75810 97800 75940
rect 97950 75810 98050 75940
rect 98200 75810 98300 75940
rect 98450 75810 98550 75940
rect 98700 75810 98800 75940
rect 98950 75810 99050 75940
rect 99200 75810 99300 75940
rect 99450 75810 99550 75940
rect 99700 75810 99800 75940
rect 99950 75810 100050 75940
rect 100200 75810 100300 75940
rect 100450 75810 100550 75940
rect 100700 75810 100800 75940
rect 100950 75810 101050 75940
rect 101200 75810 101300 75940
rect 101450 75810 101550 75940
rect 101700 75810 101800 75940
rect 101950 75810 102050 75940
rect 102200 75810 102300 75940
rect 102450 75810 102550 75940
rect 102700 75810 102800 75940
rect 102950 75810 103050 75940
rect 103200 75810 103300 75940
rect 103450 75810 103550 75940
rect 103700 75810 103800 75940
rect 103950 75810 104050 75940
rect 104200 75810 104300 75940
rect 104450 75810 104550 75940
rect 104700 75810 104800 75940
rect 104950 75810 105050 75940
rect 105200 75810 105300 75940
rect 105450 75810 105550 75940
rect 105700 75810 105800 75940
rect 105950 75810 106050 75940
rect 106200 75810 106300 75940
rect 106450 75810 106550 75940
rect 106700 75810 106800 75940
rect 106950 75810 107050 75940
rect 107200 75810 107300 75940
rect 107450 75810 107550 75940
rect 107700 75810 107800 75940
rect 107950 75810 108050 75940
rect 108200 75810 108300 75940
rect 108450 75810 108550 75940
rect 108700 75810 108800 75940
rect 108950 75810 109050 75940
rect 109200 75810 109300 75940
rect 109450 75810 109550 75940
rect 109700 75810 109800 75940
rect 109950 75810 110050 75940
rect 110200 75810 110300 75940
rect 110450 75810 110550 75940
rect 110700 75810 110800 75940
rect 110950 75810 111050 75940
rect 111200 75810 111300 75940
rect 111450 75810 111550 75940
rect 111700 75810 111800 75940
rect 111950 75810 112050 75940
rect 112200 75810 112300 75940
rect 112450 75810 112550 75940
rect 112700 75810 112800 75940
rect 112950 75810 113050 75940
rect 113200 75810 113300 75940
rect 113450 75810 113550 75940
rect 113700 75810 113800 75940
rect 113950 75810 114050 75940
rect 114200 75810 114300 75940
rect 114450 75810 114550 75940
rect 114700 75810 114800 75940
rect 114950 75810 115050 75940
rect 115200 75810 115300 75940
rect 115450 75810 115550 75940
rect 115700 75810 115800 75940
rect 115950 75810 116000 75940
rect 89000 75800 89060 75810
rect 89190 75800 89310 75810
rect 89440 75800 89560 75810
rect 89690 75800 89810 75810
rect 89940 75800 90060 75810
rect 90190 75800 90310 75810
rect 90440 75800 90560 75810
rect 90690 75800 90810 75810
rect 90940 75800 91060 75810
rect 91190 75800 91310 75810
rect 91440 75800 91560 75810
rect 91690 75800 91810 75810
rect 91940 75800 92060 75810
rect 92190 75800 92310 75810
rect 92440 75800 92560 75810
rect 92690 75800 92810 75810
rect 92940 75800 93060 75810
rect 93190 75800 93310 75810
rect 93440 75800 93560 75810
rect 93690 75800 93810 75810
rect 93940 75800 94060 75810
rect 94190 75800 94310 75810
rect 94440 75800 94560 75810
rect 94690 75800 94810 75810
rect 94940 75800 95060 75810
rect 95190 75800 95310 75810
rect 95440 75800 95560 75810
rect 95690 75800 95810 75810
rect 95940 75800 96060 75810
rect 96190 75800 96310 75810
rect 96440 75800 96560 75810
rect 96690 75800 96810 75810
rect 96940 75800 97060 75810
rect 97190 75800 97310 75810
rect 97440 75800 97560 75810
rect 97690 75800 97810 75810
rect 97940 75800 98060 75810
rect 98190 75800 98310 75810
rect 98440 75800 98560 75810
rect 98690 75800 98810 75810
rect 98940 75800 99060 75810
rect 99190 75800 99310 75810
rect 99440 75800 99560 75810
rect 99690 75800 99810 75810
rect 99940 75800 100060 75810
rect 100190 75800 100310 75810
rect 100440 75800 100560 75810
rect 100690 75800 100810 75810
rect 100940 75800 101060 75810
rect 101190 75800 101310 75810
rect 101440 75800 101560 75810
rect 101690 75800 101810 75810
rect 101940 75800 102060 75810
rect 102190 75800 102310 75810
rect 102440 75800 102560 75810
rect 102690 75800 102810 75810
rect 102940 75800 103060 75810
rect 103190 75800 103310 75810
rect 103440 75800 103560 75810
rect 103690 75800 103810 75810
rect 103940 75800 104060 75810
rect 104190 75800 104310 75810
rect 104440 75800 104560 75810
rect 104690 75800 104810 75810
rect 104940 75800 105060 75810
rect 105190 75800 105310 75810
rect 105440 75800 105560 75810
rect 105690 75800 105810 75810
rect 105940 75800 106060 75810
rect 106190 75800 106310 75810
rect 106440 75800 106560 75810
rect 106690 75800 106810 75810
rect 106940 75800 107060 75810
rect 107190 75800 107310 75810
rect 107440 75800 107560 75810
rect 107690 75800 107810 75810
rect 107940 75800 108060 75810
rect 108190 75800 108310 75810
rect 108440 75800 108560 75810
rect 108690 75800 108810 75810
rect 108940 75800 109060 75810
rect 109190 75800 109310 75810
rect 109440 75800 109560 75810
rect 109690 75800 109810 75810
rect 109940 75800 110060 75810
rect 110190 75800 110310 75810
rect 110440 75800 110560 75810
rect 110690 75800 110810 75810
rect 110940 75800 111060 75810
rect 111190 75800 111310 75810
rect 111440 75800 111560 75810
rect 111690 75800 111810 75810
rect 111940 75800 112060 75810
rect 112190 75800 112310 75810
rect 112440 75800 112560 75810
rect 112690 75800 112810 75810
rect 112940 75800 113060 75810
rect 113190 75800 113310 75810
rect 113440 75800 113560 75810
rect 113690 75800 113810 75810
rect 113940 75800 114060 75810
rect 114190 75800 114310 75810
rect 114440 75800 114560 75810
rect 114690 75800 114810 75810
rect 114940 75800 115060 75810
rect 115190 75800 115310 75810
rect 115440 75800 115560 75810
rect 115690 75800 115810 75810
rect 115940 75800 116000 75810
rect 89000 75700 116000 75800
rect 89000 75690 89060 75700
rect 89190 75690 89310 75700
rect 89440 75690 89560 75700
rect 89690 75690 89810 75700
rect 89940 75690 90060 75700
rect 90190 75690 90310 75700
rect 90440 75690 90560 75700
rect 90690 75690 90810 75700
rect 90940 75690 91060 75700
rect 91190 75690 91310 75700
rect 91440 75690 91560 75700
rect 91690 75690 91810 75700
rect 91940 75690 92060 75700
rect 92190 75690 92310 75700
rect 92440 75690 92560 75700
rect 92690 75690 92810 75700
rect 92940 75690 93060 75700
rect 93190 75690 93310 75700
rect 93440 75690 93560 75700
rect 93690 75690 93810 75700
rect 93940 75690 94060 75700
rect 94190 75690 94310 75700
rect 94440 75690 94560 75700
rect 94690 75690 94810 75700
rect 94940 75690 95060 75700
rect 95190 75690 95310 75700
rect 95440 75690 95560 75700
rect 95690 75690 95810 75700
rect 95940 75690 96060 75700
rect 96190 75690 96310 75700
rect 96440 75690 96560 75700
rect 96690 75690 96810 75700
rect 96940 75690 97060 75700
rect 97190 75690 97310 75700
rect 97440 75690 97560 75700
rect 97690 75690 97810 75700
rect 97940 75690 98060 75700
rect 98190 75690 98310 75700
rect 98440 75690 98560 75700
rect 98690 75690 98810 75700
rect 98940 75690 99060 75700
rect 99190 75690 99310 75700
rect 99440 75690 99560 75700
rect 99690 75690 99810 75700
rect 99940 75690 100060 75700
rect 100190 75690 100310 75700
rect 100440 75690 100560 75700
rect 100690 75690 100810 75700
rect 100940 75690 101060 75700
rect 101190 75690 101310 75700
rect 101440 75690 101560 75700
rect 101690 75690 101810 75700
rect 101940 75690 102060 75700
rect 102190 75690 102310 75700
rect 102440 75690 102560 75700
rect 102690 75690 102810 75700
rect 102940 75690 103060 75700
rect 103190 75690 103310 75700
rect 103440 75690 103560 75700
rect 103690 75690 103810 75700
rect 103940 75690 104060 75700
rect 104190 75690 104310 75700
rect 104440 75690 104560 75700
rect 104690 75690 104810 75700
rect 104940 75690 105060 75700
rect 105190 75690 105310 75700
rect 105440 75690 105560 75700
rect 105690 75690 105810 75700
rect 105940 75690 106060 75700
rect 106190 75690 106310 75700
rect 106440 75690 106560 75700
rect 106690 75690 106810 75700
rect 106940 75690 107060 75700
rect 107190 75690 107310 75700
rect 107440 75690 107560 75700
rect 107690 75690 107810 75700
rect 107940 75690 108060 75700
rect 108190 75690 108310 75700
rect 108440 75690 108560 75700
rect 108690 75690 108810 75700
rect 108940 75690 109060 75700
rect 109190 75690 109310 75700
rect 109440 75690 109560 75700
rect 109690 75690 109810 75700
rect 109940 75690 110060 75700
rect 110190 75690 110310 75700
rect 110440 75690 110560 75700
rect 110690 75690 110810 75700
rect 110940 75690 111060 75700
rect 111190 75690 111310 75700
rect 111440 75690 111560 75700
rect 111690 75690 111810 75700
rect 111940 75690 112060 75700
rect 112190 75690 112310 75700
rect 112440 75690 112560 75700
rect 112690 75690 112810 75700
rect 112940 75690 113060 75700
rect 113190 75690 113310 75700
rect 113440 75690 113560 75700
rect 113690 75690 113810 75700
rect 113940 75690 114060 75700
rect 114190 75690 114310 75700
rect 114440 75690 114560 75700
rect 114690 75690 114810 75700
rect 114940 75690 115060 75700
rect 115190 75690 115310 75700
rect 115440 75690 115560 75700
rect 115690 75690 115810 75700
rect 115940 75690 116000 75700
rect 89000 75560 89050 75690
rect 89200 75560 89300 75690
rect 89450 75560 89550 75690
rect 89700 75560 89800 75690
rect 89950 75560 90050 75690
rect 90200 75560 90300 75690
rect 90450 75560 90550 75690
rect 90700 75560 90800 75690
rect 90950 75560 91050 75690
rect 91200 75560 91300 75690
rect 91450 75560 91550 75690
rect 91700 75560 91800 75690
rect 91950 75560 92050 75690
rect 92200 75560 92300 75690
rect 92450 75560 92550 75690
rect 92700 75560 92800 75690
rect 92950 75560 93050 75690
rect 93200 75560 93300 75690
rect 93450 75560 93550 75690
rect 93700 75560 93800 75690
rect 93950 75560 94050 75690
rect 94200 75560 94300 75690
rect 94450 75560 94550 75690
rect 94700 75560 94800 75690
rect 94950 75560 95050 75690
rect 95200 75560 95300 75690
rect 95450 75560 95550 75690
rect 95700 75560 95800 75690
rect 95950 75560 96050 75690
rect 96200 75560 96300 75690
rect 96450 75560 96550 75690
rect 96700 75560 96800 75690
rect 96950 75560 97050 75690
rect 97200 75560 97300 75690
rect 97450 75560 97550 75690
rect 97700 75560 97800 75690
rect 97950 75560 98050 75690
rect 98200 75560 98300 75690
rect 98450 75560 98550 75690
rect 98700 75560 98800 75690
rect 98950 75560 99050 75690
rect 99200 75560 99300 75690
rect 99450 75560 99550 75690
rect 99700 75560 99800 75690
rect 99950 75560 100050 75690
rect 100200 75560 100300 75690
rect 100450 75560 100550 75690
rect 100700 75560 100800 75690
rect 100950 75560 101050 75690
rect 101200 75560 101300 75690
rect 101450 75560 101550 75690
rect 101700 75560 101800 75690
rect 101950 75560 102050 75690
rect 102200 75560 102300 75690
rect 102450 75560 102550 75690
rect 102700 75560 102800 75690
rect 102950 75560 103050 75690
rect 103200 75560 103300 75690
rect 103450 75560 103550 75690
rect 103700 75560 103800 75690
rect 103950 75560 104050 75690
rect 104200 75560 104300 75690
rect 104450 75560 104550 75690
rect 104700 75560 104800 75690
rect 104950 75560 105050 75690
rect 105200 75560 105300 75690
rect 105450 75560 105550 75690
rect 105700 75560 105800 75690
rect 105950 75560 106050 75690
rect 106200 75560 106300 75690
rect 106450 75560 106550 75690
rect 106700 75560 106800 75690
rect 106950 75560 107050 75690
rect 107200 75560 107300 75690
rect 107450 75560 107550 75690
rect 107700 75560 107800 75690
rect 107950 75560 108050 75690
rect 108200 75560 108300 75690
rect 108450 75560 108550 75690
rect 108700 75560 108800 75690
rect 108950 75560 109050 75690
rect 109200 75560 109300 75690
rect 109450 75560 109550 75690
rect 109700 75560 109800 75690
rect 109950 75560 110050 75690
rect 110200 75560 110300 75690
rect 110450 75560 110550 75690
rect 110700 75560 110800 75690
rect 110950 75560 111050 75690
rect 111200 75560 111300 75690
rect 111450 75560 111550 75690
rect 111700 75560 111800 75690
rect 111950 75560 112050 75690
rect 112200 75560 112300 75690
rect 112450 75560 112550 75690
rect 112700 75560 112800 75690
rect 112950 75560 113050 75690
rect 113200 75560 113300 75690
rect 113450 75560 113550 75690
rect 113700 75560 113800 75690
rect 113950 75560 114050 75690
rect 114200 75560 114300 75690
rect 114450 75560 114550 75690
rect 114700 75560 114800 75690
rect 114950 75560 115050 75690
rect 115200 75560 115300 75690
rect 115450 75560 115550 75690
rect 115700 75560 115800 75690
rect 115950 75560 116000 75690
rect 89000 75550 89060 75560
rect 89190 75550 89310 75560
rect 89440 75550 89560 75560
rect 89690 75550 89810 75560
rect 89940 75550 90060 75560
rect 90190 75550 90310 75560
rect 90440 75550 90560 75560
rect 90690 75550 90810 75560
rect 90940 75550 91060 75560
rect 91190 75550 91310 75560
rect 91440 75550 91560 75560
rect 91690 75550 91810 75560
rect 91940 75550 92060 75560
rect 92190 75550 92310 75560
rect 92440 75550 92560 75560
rect 92690 75550 92810 75560
rect 92940 75550 93060 75560
rect 93190 75550 93310 75560
rect 93440 75550 93560 75560
rect 93690 75550 93810 75560
rect 93940 75550 94060 75560
rect 94190 75550 94310 75560
rect 94440 75550 94560 75560
rect 94690 75550 94810 75560
rect 94940 75550 95060 75560
rect 95190 75550 95310 75560
rect 95440 75550 95560 75560
rect 95690 75550 95810 75560
rect 95940 75550 96060 75560
rect 96190 75550 96310 75560
rect 96440 75550 96560 75560
rect 96690 75550 96810 75560
rect 96940 75550 97060 75560
rect 97190 75550 97310 75560
rect 97440 75550 97560 75560
rect 97690 75550 97810 75560
rect 97940 75550 98060 75560
rect 98190 75550 98310 75560
rect 98440 75550 98560 75560
rect 98690 75550 98810 75560
rect 98940 75550 99060 75560
rect 99190 75550 99310 75560
rect 99440 75550 99560 75560
rect 99690 75550 99810 75560
rect 99940 75550 100060 75560
rect 100190 75550 100310 75560
rect 100440 75550 100560 75560
rect 100690 75550 100810 75560
rect 100940 75550 101060 75560
rect 101190 75550 101310 75560
rect 101440 75550 101560 75560
rect 101690 75550 101810 75560
rect 101940 75550 102060 75560
rect 102190 75550 102310 75560
rect 102440 75550 102560 75560
rect 102690 75550 102810 75560
rect 102940 75550 103060 75560
rect 103190 75550 103310 75560
rect 103440 75550 103560 75560
rect 103690 75550 103810 75560
rect 103940 75550 104060 75560
rect 104190 75550 104310 75560
rect 104440 75550 104560 75560
rect 104690 75550 104810 75560
rect 104940 75550 105060 75560
rect 105190 75550 105310 75560
rect 105440 75550 105560 75560
rect 105690 75550 105810 75560
rect 105940 75550 106060 75560
rect 106190 75550 106310 75560
rect 106440 75550 106560 75560
rect 106690 75550 106810 75560
rect 106940 75550 107060 75560
rect 107190 75550 107310 75560
rect 107440 75550 107560 75560
rect 107690 75550 107810 75560
rect 107940 75550 108060 75560
rect 108190 75550 108310 75560
rect 108440 75550 108560 75560
rect 108690 75550 108810 75560
rect 108940 75550 109060 75560
rect 109190 75550 109310 75560
rect 109440 75550 109560 75560
rect 109690 75550 109810 75560
rect 109940 75550 110060 75560
rect 110190 75550 110310 75560
rect 110440 75550 110560 75560
rect 110690 75550 110810 75560
rect 110940 75550 111060 75560
rect 111190 75550 111310 75560
rect 111440 75550 111560 75560
rect 111690 75550 111810 75560
rect 111940 75550 112060 75560
rect 112190 75550 112310 75560
rect 112440 75550 112560 75560
rect 112690 75550 112810 75560
rect 112940 75550 113060 75560
rect 113190 75550 113310 75560
rect 113440 75550 113560 75560
rect 113690 75550 113810 75560
rect 113940 75550 114060 75560
rect 114190 75550 114310 75560
rect 114440 75550 114560 75560
rect 114690 75550 114810 75560
rect 114940 75550 115060 75560
rect 115190 75550 115310 75560
rect 115440 75550 115560 75560
rect 115690 75550 115810 75560
rect 115940 75550 116000 75560
rect 89000 75450 116000 75550
rect 89000 75440 89060 75450
rect 89190 75440 89310 75450
rect 89440 75440 89560 75450
rect 89690 75440 89810 75450
rect 89940 75440 90060 75450
rect 90190 75440 90310 75450
rect 90440 75440 90560 75450
rect 90690 75440 90810 75450
rect 90940 75440 91060 75450
rect 91190 75440 91310 75450
rect 91440 75440 91560 75450
rect 91690 75440 91810 75450
rect 91940 75440 92060 75450
rect 92190 75440 92310 75450
rect 92440 75440 92560 75450
rect 92690 75440 92810 75450
rect 92940 75440 93060 75450
rect 93190 75440 93310 75450
rect 93440 75440 93560 75450
rect 93690 75440 93810 75450
rect 93940 75440 94060 75450
rect 94190 75440 94310 75450
rect 94440 75440 94560 75450
rect 94690 75440 94810 75450
rect 94940 75440 95060 75450
rect 95190 75440 95310 75450
rect 95440 75440 95560 75450
rect 95690 75440 95810 75450
rect 95940 75440 96060 75450
rect 96190 75440 96310 75450
rect 96440 75440 96560 75450
rect 96690 75440 96810 75450
rect 96940 75440 97060 75450
rect 97190 75440 97310 75450
rect 97440 75440 97560 75450
rect 97690 75440 97810 75450
rect 97940 75440 98060 75450
rect 98190 75440 98310 75450
rect 98440 75440 98560 75450
rect 98690 75440 98810 75450
rect 98940 75440 99060 75450
rect 99190 75440 99310 75450
rect 99440 75440 99560 75450
rect 99690 75440 99810 75450
rect 99940 75440 100060 75450
rect 100190 75440 100310 75450
rect 100440 75440 100560 75450
rect 100690 75440 100810 75450
rect 100940 75440 101060 75450
rect 101190 75440 101310 75450
rect 101440 75440 101560 75450
rect 101690 75440 101810 75450
rect 101940 75440 102060 75450
rect 102190 75440 102310 75450
rect 102440 75440 102560 75450
rect 102690 75440 102810 75450
rect 102940 75440 103060 75450
rect 103190 75440 103310 75450
rect 103440 75440 103560 75450
rect 103690 75440 103810 75450
rect 103940 75440 104060 75450
rect 104190 75440 104310 75450
rect 104440 75440 104560 75450
rect 104690 75440 104810 75450
rect 104940 75440 105060 75450
rect 105190 75440 105310 75450
rect 105440 75440 105560 75450
rect 105690 75440 105810 75450
rect 105940 75440 106060 75450
rect 106190 75440 106310 75450
rect 106440 75440 106560 75450
rect 106690 75440 106810 75450
rect 106940 75440 107060 75450
rect 107190 75440 107310 75450
rect 107440 75440 107560 75450
rect 107690 75440 107810 75450
rect 107940 75440 108060 75450
rect 108190 75440 108310 75450
rect 108440 75440 108560 75450
rect 108690 75440 108810 75450
rect 108940 75440 109060 75450
rect 109190 75440 109310 75450
rect 109440 75440 109560 75450
rect 109690 75440 109810 75450
rect 109940 75440 110060 75450
rect 110190 75440 110310 75450
rect 110440 75440 110560 75450
rect 110690 75440 110810 75450
rect 110940 75440 111060 75450
rect 111190 75440 111310 75450
rect 111440 75440 111560 75450
rect 111690 75440 111810 75450
rect 111940 75440 112060 75450
rect 112190 75440 112310 75450
rect 112440 75440 112560 75450
rect 112690 75440 112810 75450
rect 112940 75440 113060 75450
rect 113190 75440 113310 75450
rect 113440 75440 113560 75450
rect 113690 75440 113810 75450
rect 113940 75440 114060 75450
rect 114190 75440 114310 75450
rect 114440 75440 114560 75450
rect 114690 75440 114810 75450
rect 114940 75440 115060 75450
rect 115190 75440 115310 75450
rect 115440 75440 115560 75450
rect 115690 75440 115810 75450
rect 115940 75440 116000 75450
rect 89000 75310 89050 75440
rect 89200 75310 89300 75440
rect 89450 75310 89550 75440
rect 89700 75310 89800 75440
rect 89950 75310 90050 75440
rect 90200 75310 90300 75440
rect 90450 75310 90550 75440
rect 90700 75310 90800 75440
rect 90950 75310 91050 75440
rect 91200 75310 91300 75440
rect 91450 75310 91550 75440
rect 91700 75310 91800 75440
rect 91950 75310 92050 75440
rect 92200 75310 92300 75440
rect 92450 75310 92550 75440
rect 92700 75310 92800 75440
rect 92950 75310 93050 75440
rect 93200 75310 93300 75440
rect 93450 75310 93550 75440
rect 93700 75310 93800 75440
rect 93950 75310 94050 75440
rect 94200 75310 94300 75440
rect 94450 75310 94550 75440
rect 94700 75310 94800 75440
rect 94950 75310 95050 75440
rect 95200 75310 95300 75440
rect 95450 75310 95550 75440
rect 95700 75310 95800 75440
rect 95950 75310 96050 75440
rect 96200 75310 96300 75440
rect 96450 75310 96550 75440
rect 96700 75310 96800 75440
rect 96950 75310 97050 75440
rect 97200 75310 97300 75440
rect 97450 75310 97550 75440
rect 97700 75310 97800 75440
rect 97950 75310 98050 75440
rect 98200 75310 98300 75440
rect 98450 75310 98550 75440
rect 98700 75310 98800 75440
rect 98950 75310 99050 75440
rect 99200 75310 99300 75440
rect 99450 75310 99550 75440
rect 99700 75310 99800 75440
rect 99950 75310 100050 75440
rect 100200 75310 100300 75440
rect 100450 75310 100550 75440
rect 100700 75310 100800 75440
rect 100950 75310 101050 75440
rect 101200 75310 101300 75440
rect 101450 75310 101550 75440
rect 101700 75310 101800 75440
rect 101950 75310 102050 75440
rect 102200 75310 102300 75440
rect 102450 75310 102550 75440
rect 102700 75310 102800 75440
rect 102950 75310 103050 75440
rect 103200 75310 103300 75440
rect 103450 75310 103550 75440
rect 103700 75310 103800 75440
rect 103950 75310 104050 75440
rect 104200 75310 104300 75440
rect 104450 75310 104550 75440
rect 104700 75310 104800 75440
rect 104950 75310 105050 75440
rect 105200 75310 105300 75440
rect 105450 75310 105550 75440
rect 105700 75310 105800 75440
rect 105950 75310 106050 75440
rect 106200 75310 106300 75440
rect 106450 75310 106550 75440
rect 106700 75310 106800 75440
rect 106950 75310 107050 75440
rect 107200 75310 107300 75440
rect 107450 75310 107550 75440
rect 107700 75310 107800 75440
rect 107950 75310 108050 75440
rect 108200 75310 108300 75440
rect 108450 75310 108550 75440
rect 108700 75310 108800 75440
rect 108950 75310 109050 75440
rect 109200 75310 109300 75440
rect 109450 75310 109550 75440
rect 109700 75310 109800 75440
rect 109950 75310 110050 75440
rect 110200 75310 110300 75440
rect 110450 75310 110550 75440
rect 110700 75310 110800 75440
rect 110950 75310 111050 75440
rect 111200 75310 111300 75440
rect 111450 75310 111550 75440
rect 111700 75310 111800 75440
rect 111950 75310 112050 75440
rect 112200 75310 112300 75440
rect 112450 75310 112550 75440
rect 112700 75310 112800 75440
rect 112950 75310 113050 75440
rect 113200 75310 113300 75440
rect 113450 75310 113550 75440
rect 113700 75310 113800 75440
rect 113950 75310 114050 75440
rect 114200 75310 114300 75440
rect 114450 75310 114550 75440
rect 114700 75310 114800 75440
rect 114950 75310 115050 75440
rect 115200 75310 115300 75440
rect 115450 75310 115550 75440
rect 115700 75310 115800 75440
rect 115950 75310 116000 75440
rect 89000 75300 89060 75310
rect 89190 75300 89310 75310
rect 89440 75300 89560 75310
rect 89690 75300 89810 75310
rect 89940 75300 90060 75310
rect 90190 75300 90310 75310
rect 90440 75300 90560 75310
rect 90690 75300 90810 75310
rect 90940 75300 91060 75310
rect 91190 75300 91310 75310
rect 91440 75300 91560 75310
rect 91690 75300 91810 75310
rect 91940 75300 92060 75310
rect 92190 75300 92310 75310
rect 92440 75300 92560 75310
rect 92690 75300 92810 75310
rect 92940 75300 93060 75310
rect 93190 75300 93310 75310
rect 93440 75300 93560 75310
rect 93690 75300 93810 75310
rect 93940 75300 94060 75310
rect 94190 75300 94310 75310
rect 94440 75300 94560 75310
rect 94690 75300 94810 75310
rect 94940 75300 95060 75310
rect 95190 75300 95310 75310
rect 95440 75300 95560 75310
rect 95690 75300 95810 75310
rect 95940 75300 96060 75310
rect 96190 75300 96310 75310
rect 96440 75300 96560 75310
rect 96690 75300 96810 75310
rect 96940 75300 97060 75310
rect 97190 75300 97310 75310
rect 97440 75300 97560 75310
rect 97690 75300 97810 75310
rect 97940 75300 98060 75310
rect 98190 75300 98310 75310
rect 98440 75300 98560 75310
rect 98690 75300 98810 75310
rect 98940 75300 99060 75310
rect 99190 75300 99310 75310
rect 99440 75300 99560 75310
rect 99690 75300 99810 75310
rect 99940 75300 100060 75310
rect 100190 75300 100310 75310
rect 100440 75300 100560 75310
rect 100690 75300 100810 75310
rect 100940 75300 101060 75310
rect 101190 75300 101310 75310
rect 101440 75300 101560 75310
rect 101690 75300 101810 75310
rect 101940 75300 102060 75310
rect 102190 75300 102310 75310
rect 102440 75300 102560 75310
rect 102690 75300 102810 75310
rect 102940 75300 103060 75310
rect 103190 75300 103310 75310
rect 103440 75300 103560 75310
rect 103690 75300 103810 75310
rect 103940 75300 104060 75310
rect 104190 75300 104310 75310
rect 104440 75300 104560 75310
rect 104690 75300 104810 75310
rect 104940 75300 105060 75310
rect 105190 75300 105310 75310
rect 105440 75300 105560 75310
rect 105690 75300 105810 75310
rect 105940 75300 106060 75310
rect 106190 75300 106310 75310
rect 106440 75300 106560 75310
rect 106690 75300 106810 75310
rect 106940 75300 107060 75310
rect 107190 75300 107310 75310
rect 107440 75300 107560 75310
rect 107690 75300 107810 75310
rect 107940 75300 108060 75310
rect 108190 75300 108310 75310
rect 108440 75300 108560 75310
rect 108690 75300 108810 75310
rect 108940 75300 109060 75310
rect 109190 75300 109310 75310
rect 109440 75300 109560 75310
rect 109690 75300 109810 75310
rect 109940 75300 110060 75310
rect 110190 75300 110310 75310
rect 110440 75300 110560 75310
rect 110690 75300 110810 75310
rect 110940 75300 111060 75310
rect 111190 75300 111310 75310
rect 111440 75300 111560 75310
rect 111690 75300 111810 75310
rect 111940 75300 112060 75310
rect 112190 75300 112310 75310
rect 112440 75300 112560 75310
rect 112690 75300 112810 75310
rect 112940 75300 113060 75310
rect 113190 75300 113310 75310
rect 113440 75300 113560 75310
rect 113690 75300 113810 75310
rect 113940 75300 114060 75310
rect 114190 75300 114310 75310
rect 114440 75300 114560 75310
rect 114690 75300 114810 75310
rect 114940 75300 115060 75310
rect 115190 75300 115310 75310
rect 115440 75300 115560 75310
rect 115690 75300 115810 75310
rect 115940 75300 116000 75310
rect 89000 75200 116000 75300
rect 89000 75190 89060 75200
rect 89190 75190 89310 75200
rect 89440 75190 89560 75200
rect 89690 75190 89810 75200
rect 89940 75190 90060 75200
rect 90190 75190 90310 75200
rect 90440 75190 90560 75200
rect 90690 75190 90810 75200
rect 90940 75190 91060 75200
rect 91190 75190 91310 75200
rect 91440 75190 91560 75200
rect 91690 75190 91810 75200
rect 91940 75190 92060 75200
rect 92190 75190 92310 75200
rect 92440 75190 92560 75200
rect 92690 75190 92810 75200
rect 92940 75190 93060 75200
rect 93190 75190 93310 75200
rect 93440 75190 93560 75200
rect 93690 75190 93810 75200
rect 93940 75190 94060 75200
rect 94190 75190 94310 75200
rect 94440 75190 94560 75200
rect 94690 75190 94810 75200
rect 94940 75190 95060 75200
rect 95190 75190 95310 75200
rect 95440 75190 95560 75200
rect 95690 75190 95810 75200
rect 95940 75190 96060 75200
rect 96190 75190 96310 75200
rect 96440 75190 96560 75200
rect 96690 75190 96810 75200
rect 96940 75190 97060 75200
rect 97190 75190 97310 75200
rect 97440 75190 97560 75200
rect 97690 75190 97810 75200
rect 97940 75190 98060 75200
rect 98190 75190 98310 75200
rect 98440 75190 98560 75200
rect 98690 75190 98810 75200
rect 98940 75190 99060 75200
rect 99190 75190 99310 75200
rect 99440 75190 99560 75200
rect 99690 75190 99810 75200
rect 99940 75190 100060 75200
rect 100190 75190 100310 75200
rect 100440 75190 100560 75200
rect 100690 75190 100810 75200
rect 100940 75190 101060 75200
rect 101190 75190 101310 75200
rect 101440 75190 101560 75200
rect 101690 75190 101810 75200
rect 101940 75190 102060 75200
rect 102190 75190 102310 75200
rect 102440 75190 102560 75200
rect 102690 75190 102810 75200
rect 102940 75190 103060 75200
rect 103190 75190 103310 75200
rect 103440 75190 103560 75200
rect 103690 75190 103810 75200
rect 103940 75190 104060 75200
rect 104190 75190 104310 75200
rect 104440 75190 104560 75200
rect 104690 75190 104810 75200
rect 104940 75190 105060 75200
rect 105190 75190 105310 75200
rect 105440 75190 105560 75200
rect 105690 75190 105810 75200
rect 105940 75190 106060 75200
rect 106190 75190 106310 75200
rect 106440 75190 106560 75200
rect 106690 75190 106810 75200
rect 106940 75190 107060 75200
rect 107190 75190 107310 75200
rect 107440 75190 107560 75200
rect 107690 75190 107810 75200
rect 107940 75190 108060 75200
rect 108190 75190 108310 75200
rect 108440 75190 108560 75200
rect 108690 75190 108810 75200
rect 108940 75190 109060 75200
rect 109190 75190 109310 75200
rect 109440 75190 109560 75200
rect 109690 75190 109810 75200
rect 109940 75190 110060 75200
rect 110190 75190 110310 75200
rect 110440 75190 110560 75200
rect 110690 75190 110810 75200
rect 110940 75190 111060 75200
rect 111190 75190 111310 75200
rect 111440 75190 111560 75200
rect 111690 75190 111810 75200
rect 111940 75190 112060 75200
rect 112190 75190 112310 75200
rect 112440 75190 112560 75200
rect 112690 75190 112810 75200
rect 112940 75190 113060 75200
rect 113190 75190 113310 75200
rect 113440 75190 113560 75200
rect 113690 75190 113810 75200
rect 113940 75190 114060 75200
rect 114190 75190 114310 75200
rect 114440 75190 114560 75200
rect 114690 75190 114810 75200
rect 114940 75190 115060 75200
rect 115190 75190 115310 75200
rect 115440 75190 115560 75200
rect 115690 75190 115810 75200
rect 115940 75190 116000 75200
rect 89000 75060 89050 75190
rect 89200 75060 89300 75190
rect 89450 75060 89550 75190
rect 89700 75060 89800 75190
rect 89950 75060 90050 75190
rect 90200 75060 90300 75190
rect 90450 75060 90550 75190
rect 90700 75060 90800 75190
rect 90950 75060 91050 75190
rect 91200 75060 91300 75190
rect 91450 75060 91550 75190
rect 91700 75060 91800 75190
rect 91950 75060 92050 75190
rect 92200 75060 92300 75190
rect 92450 75060 92550 75190
rect 92700 75060 92800 75190
rect 92950 75060 93050 75190
rect 93200 75060 93300 75190
rect 93450 75060 93550 75190
rect 93700 75060 93800 75190
rect 93950 75060 94050 75190
rect 94200 75060 94300 75190
rect 94450 75060 94550 75190
rect 94700 75060 94800 75190
rect 94950 75060 95050 75190
rect 95200 75060 95300 75190
rect 95450 75060 95550 75190
rect 95700 75060 95800 75190
rect 95950 75060 96050 75190
rect 96200 75060 96300 75190
rect 96450 75060 96550 75190
rect 96700 75060 96800 75190
rect 96950 75060 97050 75190
rect 97200 75060 97300 75190
rect 97450 75060 97550 75190
rect 97700 75060 97800 75190
rect 97950 75060 98050 75190
rect 98200 75060 98300 75190
rect 98450 75060 98550 75190
rect 98700 75060 98800 75190
rect 98950 75060 99050 75190
rect 99200 75060 99300 75190
rect 99450 75060 99550 75190
rect 99700 75060 99800 75190
rect 99950 75060 100050 75190
rect 100200 75060 100300 75190
rect 100450 75060 100550 75190
rect 100700 75060 100800 75190
rect 100950 75060 101050 75190
rect 101200 75060 101300 75190
rect 101450 75060 101550 75190
rect 101700 75060 101800 75190
rect 101950 75060 102050 75190
rect 102200 75060 102300 75190
rect 102450 75060 102550 75190
rect 102700 75060 102800 75190
rect 102950 75060 103050 75190
rect 103200 75060 103300 75190
rect 103450 75060 103550 75190
rect 103700 75060 103800 75190
rect 103950 75060 104050 75190
rect 104200 75060 104300 75190
rect 104450 75060 104550 75190
rect 104700 75060 104800 75190
rect 104950 75060 105050 75190
rect 105200 75060 105300 75190
rect 105450 75060 105550 75190
rect 105700 75060 105800 75190
rect 105950 75060 106050 75190
rect 106200 75060 106300 75190
rect 106450 75060 106550 75190
rect 106700 75060 106800 75190
rect 106950 75060 107050 75190
rect 107200 75060 107300 75190
rect 107450 75060 107550 75190
rect 107700 75060 107800 75190
rect 107950 75060 108050 75190
rect 108200 75060 108300 75190
rect 108450 75060 108550 75190
rect 108700 75060 108800 75190
rect 108950 75060 109050 75190
rect 109200 75060 109300 75190
rect 109450 75060 109550 75190
rect 109700 75060 109800 75190
rect 109950 75060 110050 75190
rect 110200 75060 110300 75190
rect 110450 75060 110550 75190
rect 110700 75060 110800 75190
rect 110950 75060 111050 75190
rect 111200 75060 111300 75190
rect 111450 75060 111550 75190
rect 111700 75060 111800 75190
rect 111950 75060 112050 75190
rect 112200 75060 112300 75190
rect 112450 75060 112550 75190
rect 112700 75060 112800 75190
rect 112950 75060 113050 75190
rect 113200 75060 113300 75190
rect 113450 75060 113550 75190
rect 113700 75060 113800 75190
rect 113950 75060 114050 75190
rect 114200 75060 114300 75190
rect 114450 75060 114550 75190
rect 114700 75060 114800 75190
rect 114950 75060 115050 75190
rect 115200 75060 115300 75190
rect 115450 75060 115550 75190
rect 115700 75060 115800 75190
rect 115950 75060 116000 75190
rect 89000 75050 89060 75060
rect 89190 75050 89310 75060
rect 89440 75050 89560 75060
rect 89690 75050 89810 75060
rect 89940 75050 90060 75060
rect 90190 75050 90310 75060
rect 90440 75050 90560 75060
rect 90690 75050 90810 75060
rect 90940 75050 91060 75060
rect 91190 75050 91310 75060
rect 91440 75050 91560 75060
rect 91690 75050 91810 75060
rect 91940 75050 92060 75060
rect 92190 75050 92310 75060
rect 92440 75050 92560 75060
rect 92690 75050 92810 75060
rect 92940 75050 93060 75060
rect 93190 75050 93310 75060
rect 93440 75050 93560 75060
rect 93690 75050 93810 75060
rect 93940 75050 94060 75060
rect 94190 75050 94310 75060
rect 94440 75050 94560 75060
rect 94690 75050 94810 75060
rect 94940 75050 95060 75060
rect 95190 75050 95310 75060
rect 95440 75050 95560 75060
rect 95690 75050 95810 75060
rect 95940 75050 96060 75060
rect 96190 75050 96310 75060
rect 96440 75050 96560 75060
rect 96690 75050 96810 75060
rect 96940 75050 97060 75060
rect 97190 75050 97310 75060
rect 97440 75050 97560 75060
rect 97690 75050 97810 75060
rect 97940 75050 98060 75060
rect 98190 75050 98310 75060
rect 98440 75050 98560 75060
rect 98690 75050 98810 75060
rect 98940 75050 99060 75060
rect 99190 75050 99310 75060
rect 99440 75050 99560 75060
rect 99690 75050 99810 75060
rect 99940 75050 100060 75060
rect 100190 75050 100310 75060
rect 100440 75050 100560 75060
rect 100690 75050 100810 75060
rect 100940 75050 101060 75060
rect 101190 75050 101310 75060
rect 101440 75050 101560 75060
rect 101690 75050 101810 75060
rect 101940 75050 102060 75060
rect 102190 75050 102310 75060
rect 102440 75050 102560 75060
rect 102690 75050 102810 75060
rect 102940 75050 103060 75060
rect 103190 75050 103310 75060
rect 103440 75050 103560 75060
rect 103690 75050 103810 75060
rect 103940 75050 104060 75060
rect 104190 75050 104310 75060
rect 104440 75050 104560 75060
rect 104690 75050 104810 75060
rect 104940 75050 105060 75060
rect 105190 75050 105310 75060
rect 105440 75050 105560 75060
rect 105690 75050 105810 75060
rect 105940 75050 106060 75060
rect 106190 75050 106310 75060
rect 106440 75050 106560 75060
rect 106690 75050 106810 75060
rect 106940 75050 107060 75060
rect 107190 75050 107310 75060
rect 107440 75050 107560 75060
rect 107690 75050 107810 75060
rect 107940 75050 108060 75060
rect 108190 75050 108310 75060
rect 108440 75050 108560 75060
rect 108690 75050 108810 75060
rect 108940 75050 109060 75060
rect 109190 75050 109310 75060
rect 109440 75050 109560 75060
rect 109690 75050 109810 75060
rect 109940 75050 110060 75060
rect 110190 75050 110310 75060
rect 110440 75050 110560 75060
rect 110690 75050 110810 75060
rect 110940 75050 111060 75060
rect 111190 75050 111310 75060
rect 111440 75050 111560 75060
rect 111690 75050 111810 75060
rect 111940 75050 112060 75060
rect 112190 75050 112310 75060
rect 112440 75050 112560 75060
rect 112690 75050 112810 75060
rect 112940 75050 113060 75060
rect 113190 75050 113310 75060
rect 113440 75050 113560 75060
rect 113690 75050 113810 75060
rect 113940 75050 114060 75060
rect 114190 75050 114310 75060
rect 114440 75050 114560 75060
rect 114690 75050 114810 75060
rect 114940 75050 115060 75060
rect 115190 75050 115310 75060
rect 115440 75050 115560 75060
rect 115690 75050 115810 75060
rect 115940 75050 116000 75060
rect 89000 74950 116000 75050
rect 89000 74940 89060 74950
rect 89190 74940 89310 74950
rect 89440 74940 89560 74950
rect 89690 74940 89810 74950
rect 89940 74940 90060 74950
rect 90190 74940 90310 74950
rect 90440 74940 90560 74950
rect 90690 74940 90810 74950
rect 90940 74940 91060 74950
rect 91190 74940 91310 74950
rect 91440 74940 91560 74950
rect 91690 74940 91810 74950
rect 91940 74940 92060 74950
rect 92190 74940 92310 74950
rect 92440 74940 92560 74950
rect 92690 74940 92810 74950
rect 92940 74940 93060 74950
rect 93190 74940 93310 74950
rect 93440 74940 93560 74950
rect 93690 74940 93810 74950
rect 93940 74940 94060 74950
rect 94190 74940 94310 74950
rect 94440 74940 94560 74950
rect 94690 74940 94810 74950
rect 94940 74940 95060 74950
rect 95190 74940 95310 74950
rect 95440 74940 95560 74950
rect 95690 74940 95810 74950
rect 95940 74940 96060 74950
rect 96190 74940 96310 74950
rect 96440 74940 96560 74950
rect 96690 74940 96810 74950
rect 96940 74940 97060 74950
rect 97190 74940 97310 74950
rect 97440 74940 97560 74950
rect 97690 74940 97810 74950
rect 97940 74940 98060 74950
rect 98190 74940 98310 74950
rect 98440 74940 98560 74950
rect 98690 74940 98810 74950
rect 98940 74940 99060 74950
rect 99190 74940 99310 74950
rect 99440 74940 99560 74950
rect 99690 74940 99810 74950
rect 99940 74940 100060 74950
rect 100190 74940 100310 74950
rect 100440 74940 100560 74950
rect 100690 74940 100810 74950
rect 100940 74940 101060 74950
rect 101190 74940 101310 74950
rect 101440 74940 101560 74950
rect 101690 74940 101810 74950
rect 101940 74940 102060 74950
rect 102190 74940 102310 74950
rect 102440 74940 102560 74950
rect 102690 74940 102810 74950
rect 102940 74940 103060 74950
rect 103190 74940 103310 74950
rect 103440 74940 103560 74950
rect 103690 74940 103810 74950
rect 103940 74940 104060 74950
rect 104190 74940 104310 74950
rect 104440 74940 104560 74950
rect 104690 74940 104810 74950
rect 104940 74940 105060 74950
rect 105190 74940 105310 74950
rect 105440 74940 105560 74950
rect 105690 74940 105810 74950
rect 105940 74940 106060 74950
rect 106190 74940 106310 74950
rect 106440 74940 106560 74950
rect 106690 74940 106810 74950
rect 106940 74940 107060 74950
rect 107190 74940 107310 74950
rect 107440 74940 107560 74950
rect 107690 74940 107810 74950
rect 107940 74940 108060 74950
rect 108190 74940 108310 74950
rect 108440 74940 108560 74950
rect 108690 74940 108810 74950
rect 108940 74940 109060 74950
rect 109190 74940 109310 74950
rect 109440 74940 109560 74950
rect 109690 74940 109810 74950
rect 109940 74940 110060 74950
rect 110190 74940 110310 74950
rect 110440 74940 110560 74950
rect 110690 74940 110810 74950
rect 110940 74940 111060 74950
rect 111190 74940 111310 74950
rect 111440 74940 111560 74950
rect 111690 74940 111810 74950
rect 111940 74940 112060 74950
rect 112190 74940 112310 74950
rect 112440 74940 112560 74950
rect 112690 74940 112810 74950
rect 112940 74940 113060 74950
rect 113190 74940 113310 74950
rect 113440 74940 113560 74950
rect 113690 74940 113810 74950
rect 113940 74940 114060 74950
rect 114190 74940 114310 74950
rect 114440 74940 114560 74950
rect 114690 74940 114810 74950
rect 114940 74940 115060 74950
rect 115190 74940 115310 74950
rect 115440 74940 115560 74950
rect 115690 74940 115810 74950
rect 115940 74940 116000 74950
rect 89000 74810 89050 74940
rect 89200 74810 89300 74940
rect 89450 74810 89550 74940
rect 89700 74810 89800 74940
rect 89950 74810 90050 74940
rect 90200 74810 90300 74940
rect 90450 74810 90550 74940
rect 90700 74810 90800 74940
rect 90950 74810 91050 74940
rect 91200 74810 91300 74940
rect 91450 74810 91550 74940
rect 91700 74810 91800 74940
rect 91950 74810 92050 74940
rect 92200 74810 92300 74940
rect 92450 74810 92550 74940
rect 92700 74810 92800 74940
rect 92950 74810 93050 74940
rect 93200 74810 93300 74940
rect 93450 74810 93550 74940
rect 93700 74810 93800 74940
rect 93950 74810 94050 74940
rect 94200 74810 94300 74940
rect 94450 74810 94550 74940
rect 94700 74810 94800 74940
rect 94950 74810 95050 74940
rect 95200 74810 95300 74940
rect 95450 74810 95550 74940
rect 95700 74810 95800 74940
rect 95950 74810 96050 74940
rect 96200 74810 96300 74940
rect 96450 74810 96550 74940
rect 96700 74810 96800 74940
rect 96950 74810 97050 74940
rect 97200 74810 97300 74940
rect 97450 74810 97550 74940
rect 97700 74810 97800 74940
rect 97950 74810 98050 74940
rect 98200 74810 98300 74940
rect 98450 74810 98550 74940
rect 98700 74810 98800 74940
rect 98950 74810 99050 74940
rect 99200 74810 99300 74940
rect 99450 74810 99550 74940
rect 99700 74810 99800 74940
rect 99950 74810 100050 74940
rect 100200 74810 100300 74940
rect 100450 74810 100550 74940
rect 100700 74810 100800 74940
rect 100950 74810 101050 74940
rect 101200 74810 101300 74940
rect 101450 74810 101550 74940
rect 101700 74810 101800 74940
rect 101950 74810 102050 74940
rect 102200 74810 102300 74940
rect 102450 74810 102550 74940
rect 102700 74810 102800 74940
rect 102950 74810 103050 74940
rect 103200 74810 103300 74940
rect 103450 74810 103550 74940
rect 103700 74810 103800 74940
rect 103950 74810 104050 74940
rect 104200 74810 104300 74940
rect 104450 74810 104550 74940
rect 104700 74810 104800 74940
rect 104950 74810 105050 74940
rect 105200 74810 105300 74940
rect 105450 74810 105550 74940
rect 105700 74810 105800 74940
rect 105950 74810 106050 74940
rect 106200 74810 106300 74940
rect 106450 74810 106550 74940
rect 106700 74810 106800 74940
rect 106950 74810 107050 74940
rect 107200 74810 107300 74940
rect 107450 74810 107550 74940
rect 107700 74810 107800 74940
rect 107950 74810 108050 74940
rect 108200 74810 108300 74940
rect 108450 74810 108550 74940
rect 108700 74810 108800 74940
rect 108950 74810 109050 74940
rect 109200 74810 109300 74940
rect 109450 74810 109550 74940
rect 109700 74810 109800 74940
rect 109950 74810 110050 74940
rect 110200 74810 110300 74940
rect 110450 74810 110550 74940
rect 110700 74810 110800 74940
rect 110950 74810 111050 74940
rect 111200 74810 111300 74940
rect 111450 74810 111550 74940
rect 111700 74810 111800 74940
rect 111950 74810 112050 74940
rect 112200 74810 112300 74940
rect 112450 74810 112550 74940
rect 112700 74810 112800 74940
rect 112950 74810 113050 74940
rect 113200 74810 113300 74940
rect 113450 74810 113550 74940
rect 113700 74810 113800 74940
rect 113950 74810 114050 74940
rect 114200 74810 114300 74940
rect 114450 74810 114550 74940
rect 114700 74810 114800 74940
rect 114950 74810 115050 74940
rect 115200 74810 115300 74940
rect 115450 74810 115550 74940
rect 115700 74810 115800 74940
rect 115950 74810 116000 74940
rect 89000 74800 89060 74810
rect 89190 74800 89310 74810
rect 89440 74800 89560 74810
rect 89690 74800 89810 74810
rect 89940 74800 90060 74810
rect 90190 74800 90310 74810
rect 90440 74800 90560 74810
rect 90690 74800 90810 74810
rect 90940 74800 91060 74810
rect 91190 74800 91310 74810
rect 91440 74800 91560 74810
rect 91690 74800 91810 74810
rect 91940 74800 92060 74810
rect 92190 74800 92310 74810
rect 92440 74800 92560 74810
rect 92690 74800 92810 74810
rect 92940 74800 93060 74810
rect 93190 74800 93310 74810
rect 93440 74800 93560 74810
rect 93690 74800 93810 74810
rect 93940 74800 94060 74810
rect 94190 74800 94310 74810
rect 94440 74800 94560 74810
rect 94690 74800 94810 74810
rect 94940 74800 95060 74810
rect 95190 74800 95310 74810
rect 95440 74800 95560 74810
rect 95690 74800 95810 74810
rect 95940 74800 96060 74810
rect 96190 74800 96310 74810
rect 96440 74800 96560 74810
rect 96690 74800 96810 74810
rect 96940 74800 97060 74810
rect 97190 74800 97310 74810
rect 97440 74800 97560 74810
rect 97690 74800 97810 74810
rect 97940 74800 98060 74810
rect 98190 74800 98310 74810
rect 98440 74800 98560 74810
rect 98690 74800 98810 74810
rect 98940 74800 99060 74810
rect 99190 74800 99310 74810
rect 99440 74800 99560 74810
rect 99690 74800 99810 74810
rect 99940 74800 100060 74810
rect 100190 74800 100310 74810
rect 100440 74800 100560 74810
rect 100690 74800 100810 74810
rect 100940 74800 101060 74810
rect 101190 74800 101310 74810
rect 101440 74800 101560 74810
rect 101690 74800 101810 74810
rect 101940 74800 102060 74810
rect 102190 74800 102310 74810
rect 102440 74800 102560 74810
rect 102690 74800 102810 74810
rect 102940 74800 103060 74810
rect 103190 74800 103310 74810
rect 103440 74800 103560 74810
rect 103690 74800 103810 74810
rect 103940 74800 104060 74810
rect 104190 74800 104310 74810
rect 104440 74800 104560 74810
rect 104690 74800 104810 74810
rect 104940 74800 105060 74810
rect 105190 74800 105310 74810
rect 105440 74800 105560 74810
rect 105690 74800 105810 74810
rect 105940 74800 106060 74810
rect 106190 74800 106310 74810
rect 106440 74800 106560 74810
rect 106690 74800 106810 74810
rect 106940 74800 107060 74810
rect 107190 74800 107310 74810
rect 107440 74800 107560 74810
rect 107690 74800 107810 74810
rect 107940 74800 108060 74810
rect 108190 74800 108310 74810
rect 108440 74800 108560 74810
rect 108690 74800 108810 74810
rect 108940 74800 109060 74810
rect 109190 74800 109310 74810
rect 109440 74800 109560 74810
rect 109690 74800 109810 74810
rect 109940 74800 110060 74810
rect 110190 74800 110310 74810
rect 110440 74800 110560 74810
rect 110690 74800 110810 74810
rect 110940 74800 111060 74810
rect 111190 74800 111310 74810
rect 111440 74800 111560 74810
rect 111690 74800 111810 74810
rect 111940 74800 112060 74810
rect 112190 74800 112310 74810
rect 112440 74800 112560 74810
rect 112690 74800 112810 74810
rect 112940 74800 113060 74810
rect 113190 74800 113310 74810
rect 113440 74800 113560 74810
rect 113690 74800 113810 74810
rect 113940 74800 114060 74810
rect 114190 74800 114310 74810
rect 114440 74800 114560 74810
rect 114690 74800 114810 74810
rect 114940 74800 115060 74810
rect 115190 74800 115310 74810
rect 115440 74800 115560 74810
rect 115690 74800 115810 74810
rect 115940 74800 116000 74810
rect 89000 74700 116000 74800
rect 89000 74690 89060 74700
rect 89190 74690 89310 74700
rect 89440 74690 89560 74700
rect 89690 74690 89810 74700
rect 89940 74690 90060 74700
rect 90190 74690 90310 74700
rect 90440 74690 90560 74700
rect 90690 74690 90810 74700
rect 90940 74690 91060 74700
rect 91190 74690 91310 74700
rect 91440 74690 91560 74700
rect 91690 74690 91810 74700
rect 91940 74690 92060 74700
rect 92190 74690 92310 74700
rect 92440 74690 92560 74700
rect 92690 74690 92810 74700
rect 92940 74690 93060 74700
rect 93190 74690 93310 74700
rect 93440 74690 93560 74700
rect 93690 74690 93810 74700
rect 93940 74690 94060 74700
rect 94190 74690 94310 74700
rect 94440 74690 94560 74700
rect 94690 74690 94810 74700
rect 94940 74690 95060 74700
rect 95190 74690 95310 74700
rect 95440 74690 95560 74700
rect 95690 74690 95810 74700
rect 95940 74690 96060 74700
rect 96190 74690 96310 74700
rect 96440 74690 96560 74700
rect 96690 74690 96810 74700
rect 96940 74690 97060 74700
rect 97190 74690 97310 74700
rect 97440 74690 97560 74700
rect 97690 74690 97810 74700
rect 97940 74690 98060 74700
rect 98190 74690 98310 74700
rect 98440 74690 98560 74700
rect 98690 74690 98810 74700
rect 98940 74690 99060 74700
rect 99190 74690 99310 74700
rect 99440 74690 99560 74700
rect 99690 74690 99810 74700
rect 99940 74690 100060 74700
rect 100190 74690 100310 74700
rect 100440 74690 100560 74700
rect 100690 74690 100810 74700
rect 100940 74690 101060 74700
rect 101190 74690 101310 74700
rect 101440 74690 101560 74700
rect 101690 74690 101810 74700
rect 101940 74690 102060 74700
rect 102190 74690 102310 74700
rect 102440 74690 102560 74700
rect 102690 74690 102810 74700
rect 102940 74690 103060 74700
rect 103190 74690 103310 74700
rect 103440 74690 103560 74700
rect 103690 74690 103810 74700
rect 103940 74690 104060 74700
rect 104190 74690 104310 74700
rect 104440 74690 104560 74700
rect 104690 74690 104810 74700
rect 104940 74690 105060 74700
rect 105190 74690 105310 74700
rect 105440 74690 105560 74700
rect 105690 74690 105810 74700
rect 105940 74690 106060 74700
rect 106190 74690 106310 74700
rect 106440 74690 106560 74700
rect 106690 74690 106810 74700
rect 106940 74690 107060 74700
rect 107190 74690 107310 74700
rect 107440 74690 107560 74700
rect 107690 74690 107810 74700
rect 107940 74690 108060 74700
rect 108190 74690 108310 74700
rect 108440 74690 108560 74700
rect 108690 74690 108810 74700
rect 108940 74690 109060 74700
rect 109190 74690 109310 74700
rect 109440 74690 109560 74700
rect 109690 74690 109810 74700
rect 109940 74690 110060 74700
rect 110190 74690 110310 74700
rect 110440 74690 110560 74700
rect 110690 74690 110810 74700
rect 110940 74690 111060 74700
rect 111190 74690 111310 74700
rect 111440 74690 111560 74700
rect 111690 74690 111810 74700
rect 111940 74690 112060 74700
rect 112190 74690 112310 74700
rect 112440 74690 112560 74700
rect 112690 74690 112810 74700
rect 112940 74690 113060 74700
rect 113190 74690 113310 74700
rect 113440 74690 113560 74700
rect 113690 74690 113810 74700
rect 113940 74690 114060 74700
rect 114190 74690 114310 74700
rect 114440 74690 114560 74700
rect 114690 74690 114810 74700
rect 114940 74690 115060 74700
rect 115190 74690 115310 74700
rect 115440 74690 115560 74700
rect 115690 74690 115810 74700
rect 115940 74690 116000 74700
rect 89000 74560 89050 74690
rect 89200 74560 89300 74690
rect 89450 74560 89550 74690
rect 89700 74560 89800 74690
rect 89950 74560 90050 74690
rect 90200 74560 90300 74690
rect 90450 74560 90550 74690
rect 90700 74560 90800 74690
rect 90950 74560 91050 74690
rect 91200 74560 91300 74690
rect 91450 74560 91550 74690
rect 91700 74560 91800 74690
rect 91950 74560 92050 74690
rect 92200 74560 92300 74690
rect 92450 74560 92550 74690
rect 92700 74560 92800 74690
rect 92950 74560 93050 74690
rect 93200 74560 93300 74690
rect 93450 74560 93550 74690
rect 93700 74560 93800 74690
rect 93950 74560 94050 74690
rect 94200 74560 94300 74690
rect 94450 74560 94550 74690
rect 94700 74560 94800 74690
rect 94950 74560 95050 74690
rect 95200 74560 95300 74690
rect 95450 74560 95550 74690
rect 95700 74560 95800 74690
rect 95950 74560 96050 74690
rect 96200 74560 96300 74690
rect 96450 74560 96550 74690
rect 96700 74560 96800 74690
rect 96950 74560 97050 74690
rect 97200 74560 97300 74690
rect 97450 74560 97550 74690
rect 97700 74560 97800 74690
rect 97950 74560 98050 74690
rect 98200 74560 98300 74690
rect 98450 74560 98550 74690
rect 98700 74560 98800 74690
rect 98950 74560 99050 74690
rect 99200 74560 99300 74690
rect 99450 74560 99550 74690
rect 99700 74560 99800 74690
rect 99950 74560 100050 74690
rect 100200 74560 100300 74690
rect 100450 74560 100550 74690
rect 100700 74560 100800 74690
rect 100950 74560 101050 74690
rect 101200 74560 101300 74690
rect 101450 74560 101550 74690
rect 101700 74560 101800 74690
rect 101950 74560 102050 74690
rect 102200 74560 102300 74690
rect 102450 74560 102550 74690
rect 102700 74560 102800 74690
rect 102950 74560 103050 74690
rect 103200 74560 103300 74690
rect 103450 74560 103550 74690
rect 103700 74560 103800 74690
rect 103950 74560 104050 74690
rect 104200 74560 104300 74690
rect 104450 74560 104550 74690
rect 104700 74560 104800 74690
rect 104950 74560 105050 74690
rect 105200 74560 105300 74690
rect 105450 74560 105550 74690
rect 105700 74560 105800 74690
rect 105950 74560 106050 74690
rect 106200 74560 106300 74690
rect 106450 74560 106550 74690
rect 106700 74560 106800 74690
rect 106950 74560 107050 74690
rect 107200 74560 107300 74690
rect 107450 74560 107550 74690
rect 107700 74560 107800 74690
rect 107950 74560 108050 74690
rect 108200 74560 108300 74690
rect 108450 74560 108550 74690
rect 108700 74560 108800 74690
rect 108950 74560 109050 74690
rect 109200 74560 109300 74690
rect 109450 74560 109550 74690
rect 109700 74560 109800 74690
rect 109950 74560 110050 74690
rect 110200 74560 110300 74690
rect 110450 74560 110550 74690
rect 110700 74560 110800 74690
rect 110950 74560 111050 74690
rect 111200 74560 111300 74690
rect 111450 74560 111550 74690
rect 111700 74560 111800 74690
rect 111950 74560 112050 74690
rect 112200 74560 112300 74690
rect 112450 74560 112550 74690
rect 112700 74560 112800 74690
rect 112950 74560 113050 74690
rect 113200 74560 113300 74690
rect 113450 74560 113550 74690
rect 113700 74560 113800 74690
rect 113950 74560 114050 74690
rect 114200 74560 114300 74690
rect 114450 74560 114550 74690
rect 114700 74560 114800 74690
rect 114950 74560 115050 74690
rect 115200 74560 115300 74690
rect 115450 74560 115550 74690
rect 115700 74560 115800 74690
rect 115950 74560 116000 74690
rect 89000 74550 89060 74560
rect 89190 74550 89310 74560
rect 89440 74550 89560 74560
rect 89690 74550 89810 74560
rect 89940 74550 90060 74560
rect 90190 74550 90310 74560
rect 90440 74550 90560 74560
rect 90690 74550 90810 74560
rect 90940 74550 91060 74560
rect 91190 74550 91310 74560
rect 91440 74550 91560 74560
rect 91690 74550 91810 74560
rect 91940 74550 92060 74560
rect 92190 74550 92310 74560
rect 92440 74550 92560 74560
rect 92690 74550 92810 74560
rect 92940 74550 93060 74560
rect 93190 74550 93310 74560
rect 93440 74550 93560 74560
rect 93690 74550 93810 74560
rect 93940 74550 94060 74560
rect 94190 74550 94310 74560
rect 94440 74550 94560 74560
rect 94690 74550 94810 74560
rect 94940 74550 95060 74560
rect 95190 74550 95310 74560
rect 95440 74550 95560 74560
rect 95690 74550 95810 74560
rect 95940 74550 96060 74560
rect 96190 74550 96310 74560
rect 96440 74550 96560 74560
rect 96690 74550 96810 74560
rect 96940 74550 97060 74560
rect 97190 74550 97310 74560
rect 97440 74550 97560 74560
rect 97690 74550 97810 74560
rect 97940 74550 98060 74560
rect 98190 74550 98310 74560
rect 98440 74550 98560 74560
rect 98690 74550 98810 74560
rect 98940 74550 99060 74560
rect 99190 74550 99310 74560
rect 99440 74550 99560 74560
rect 99690 74550 99810 74560
rect 99940 74550 100060 74560
rect 100190 74550 100310 74560
rect 100440 74550 100560 74560
rect 100690 74550 100810 74560
rect 100940 74550 101060 74560
rect 101190 74550 101310 74560
rect 101440 74550 101560 74560
rect 101690 74550 101810 74560
rect 101940 74550 102060 74560
rect 102190 74550 102310 74560
rect 102440 74550 102560 74560
rect 102690 74550 102810 74560
rect 102940 74550 103060 74560
rect 103190 74550 103310 74560
rect 103440 74550 103560 74560
rect 103690 74550 103810 74560
rect 103940 74550 104060 74560
rect 104190 74550 104310 74560
rect 104440 74550 104560 74560
rect 104690 74550 104810 74560
rect 104940 74550 105060 74560
rect 105190 74550 105310 74560
rect 105440 74550 105560 74560
rect 105690 74550 105810 74560
rect 105940 74550 106060 74560
rect 106190 74550 106310 74560
rect 106440 74550 106560 74560
rect 106690 74550 106810 74560
rect 106940 74550 107060 74560
rect 107190 74550 107310 74560
rect 107440 74550 107560 74560
rect 107690 74550 107810 74560
rect 107940 74550 108060 74560
rect 108190 74550 108310 74560
rect 108440 74550 108560 74560
rect 108690 74550 108810 74560
rect 108940 74550 109060 74560
rect 109190 74550 109310 74560
rect 109440 74550 109560 74560
rect 109690 74550 109810 74560
rect 109940 74550 110060 74560
rect 110190 74550 110310 74560
rect 110440 74550 110560 74560
rect 110690 74550 110810 74560
rect 110940 74550 111060 74560
rect 111190 74550 111310 74560
rect 111440 74550 111560 74560
rect 111690 74550 111810 74560
rect 111940 74550 112060 74560
rect 112190 74550 112310 74560
rect 112440 74550 112560 74560
rect 112690 74550 112810 74560
rect 112940 74550 113060 74560
rect 113190 74550 113310 74560
rect 113440 74550 113560 74560
rect 113690 74550 113810 74560
rect 113940 74550 114060 74560
rect 114190 74550 114310 74560
rect 114440 74550 114560 74560
rect 114690 74550 114810 74560
rect 114940 74550 115060 74560
rect 115190 74550 115310 74560
rect 115440 74550 115560 74560
rect 115690 74550 115810 74560
rect 115940 74550 116000 74560
rect 89000 74450 116000 74550
rect 89000 74440 89060 74450
rect 89190 74440 89310 74450
rect 89440 74440 89560 74450
rect 89690 74440 89810 74450
rect 89940 74440 90060 74450
rect 90190 74440 90310 74450
rect 90440 74440 90560 74450
rect 90690 74440 90810 74450
rect 90940 74440 91060 74450
rect 91190 74440 91310 74450
rect 91440 74440 91560 74450
rect 91690 74440 91810 74450
rect 91940 74440 92060 74450
rect 92190 74440 92310 74450
rect 92440 74440 92560 74450
rect 92690 74440 92810 74450
rect 92940 74440 93060 74450
rect 93190 74440 93310 74450
rect 93440 74440 93560 74450
rect 93690 74440 93810 74450
rect 93940 74440 94060 74450
rect 94190 74440 94310 74450
rect 94440 74440 94560 74450
rect 94690 74440 94810 74450
rect 94940 74440 95060 74450
rect 95190 74440 95310 74450
rect 95440 74440 95560 74450
rect 95690 74440 95810 74450
rect 95940 74440 96060 74450
rect 96190 74440 96310 74450
rect 96440 74440 96560 74450
rect 96690 74440 96810 74450
rect 96940 74440 97060 74450
rect 97190 74440 97310 74450
rect 97440 74440 97560 74450
rect 97690 74440 97810 74450
rect 97940 74440 98060 74450
rect 98190 74440 98310 74450
rect 98440 74440 98560 74450
rect 98690 74440 98810 74450
rect 98940 74440 99060 74450
rect 99190 74440 99310 74450
rect 99440 74440 99560 74450
rect 99690 74440 99810 74450
rect 99940 74440 100060 74450
rect 100190 74440 100310 74450
rect 100440 74440 100560 74450
rect 100690 74440 100810 74450
rect 100940 74440 101060 74450
rect 101190 74440 101310 74450
rect 101440 74440 101560 74450
rect 101690 74440 101810 74450
rect 101940 74440 102060 74450
rect 102190 74440 102310 74450
rect 102440 74440 102560 74450
rect 102690 74440 102810 74450
rect 102940 74440 103060 74450
rect 103190 74440 103310 74450
rect 103440 74440 103560 74450
rect 103690 74440 103810 74450
rect 103940 74440 104060 74450
rect 104190 74440 104310 74450
rect 104440 74440 104560 74450
rect 104690 74440 104810 74450
rect 104940 74440 105060 74450
rect 105190 74440 105310 74450
rect 105440 74440 105560 74450
rect 105690 74440 105810 74450
rect 105940 74440 106060 74450
rect 106190 74440 106310 74450
rect 106440 74440 106560 74450
rect 106690 74440 106810 74450
rect 106940 74440 107060 74450
rect 107190 74440 107310 74450
rect 107440 74440 107560 74450
rect 107690 74440 107810 74450
rect 107940 74440 108060 74450
rect 108190 74440 108310 74450
rect 108440 74440 108560 74450
rect 108690 74440 108810 74450
rect 108940 74440 109060 74450
rect 109190 74440 109310 74450
rect 109440 74440 109560 74450
rect 109690 74440 109810 74450
rect 109940 74440 110060 74450
rect 110190 74440 110310 74450
rect 110440 74440 110560 74450
rect 110690 74440 110810 74450
rect 110940 74440 111060 74450
rect 111190 74440 111310 74450
rect 111440 74440 111560 74450
rect 111690 74440 111810 74450
rect 111940 74440 112060 74450
rect 112190 74440 112310 74450
rect 112440 74440 112560 74450
rect 112690 74440 112810 74450
rect 112940 74440 113060 74450
rect 113190 74440 113310 74450
rect 113440 74440 113560 74450
rect 113690 74440 113810 74450
rect 113940 74440 114060 74450
rect 114190 74440 114310 74450
rect 114440 74440 114560 74450
rect 114690 74440 114810 74450
rect 114940 74440 115060 74450
rect 115190 74440 115310 74450
rect 115440 74440 115560 74450
rect 115690 74440 115810 74450
rect 115940 74440 116000 74450
rect 89000 74310 89050 74440
rect 89200 74310 89300 74440
rect 89450 74310 89550 74440
rect 89700 74310 89800 74440
rect 89950 74310 90050 74440
rect 90200 74310 90300 74440
rect 90450 74310 90550 74440
rect 90700 74310 90800 74440
rect 90950 74310 91050 74440
rect 91200 74310 91300 74440
rect 91450 74310 91550 74440
rect 91700 74310 91800 74440
rect 91950 74310 92050 74440
rect 92200 74310 92300 74440
rect 92450 74310 92550 74440
rect 92700 74310 92800 74440
rect 92950 74310 93050 74440
rect 93200 74310 93300 74440
rect 93450 74310 93550 74440
rect 93700 74310 93800 74440
rect 93950 74310 94050 74440
rect 94200 74310 94300 74440
rect 94450 74310 94550 74440
rect 94700 74310 94800 74440
rect 94950 74310 95050 74440
rect 95200 74310 95300 74440
rect 95450 74310 95550 74440
rect 95700 74310 95800 74440
rect 95950 74310 96050 74440
rect 96200 74310 96300 74440
rect 96450 74310 96550 74440
rect 96700 74310 96800 74440
rect 96950 74310 97050 74440
rect 97200 74310 97300 74440
rect 97450 74310 97550 74440
rect 97700 74310 97800 74440
rect 97950 74310 98050 74440
rect 98200 74310 98300 74440
rect 98450 74310 98550 74440
rect 98700 74310 98800 74440
rect 98950 74310 99050 74440
rect 99200 74310 99300 74440
rect 99450 74310 99550 74440
rect 99700 74310 99800 74440
rect 99950 74310 100050 74440
rect 100200 74310 100300 74440
rect 100450 74310 100550 74440
rect 100700 74310 100800 74440
rect 100950 74310 101050 74440
rect 101200 74310 101300 74440
rect 101450 74310 101550 74440
rect 101700 74310 101800 74440
rect 101950 74310 102050 74440
rect 102200 74310 102300 74440
rect 102450 74310 102550 74440
rect 102700 74310 102800 74440
rect 102950 74310 103050 74440
rect 103200 74310 103300 74440
rect 103450 74310 103550 74440
rect 103700 74310 103800 74440
rect 103950 74310 104050 74440
rect 104200 74310 104300 74440
rect 104450 74310 104550 74440
rect 104700 74310 104800 74440
rect 104950 74310 105050 74440
rect 105200 74310 105300 74440
rect 105450 74310 105550 74440
rect 105700 74310 105800 74440
rect 105950 74310 106050 74440
rect 106200 74310 106300 74440
rect 106450 74310 106550 74440
rect 106700 74310 106800 74440
rect 106950 74310 107050 74440
rect 107200 74310 107300 74440
rect 107450 74310 107550 74440
rect 107700 74310 107800 74440
rect 107950 74310 108050 74440
rect 108200 74310 108300 74440
rect 108450 74310 108550 74440
rect 108700 74310 108800 74440
rect 108950 74310 109050 74440
rect 109200 74310 109300 74440
rect 109450 74310 109550 74440
rect 109700 74310 109800 74440
rect 109950 74310 110050 74440
rect 110200 74310 110300 74440
rect 110450 74310 110550 74440
rect 110700 74310 110800 74440
rect 110950 74310 111050 74440
rect 111200 74310 111300 74440
rect 111450 74310 111550 74440
rect 111700 74310 111800 74440
rect 111950 74310 112050 74440
rect 112200 74310 112300 74440
rect 112450 74310 112550 74440
rect 112700 74310 112800 74440
rect 112950 74310 113050 74440
rect 113200 74310 113300 74440
rect 113450 74310 113550 74440
rect 113700 74310 113800 74440
rect 113950 74310 114050 74440
rect 114200 74310 114300 74440
rect 114450 74310 114550 74440
rect 114700 74310 114800 74440
rect 114950 74310 115050 74440
rect 115200 74310 115300 74440
rect 115450 74310 115550 74440
rect 115700 74310 115800 74440
rect 115950 74310 116000 74440
rect 89000 74300 89060 74310
rect 89190 74300 89310 74310
rect 89440 74300 89560 74310
rect 89690 74300 89810 74310
rect 89940 74300 90060 74310
rect 90190 74300 90310 74310
rect 90440 74300 90560 74310
rect 90690 74300 90810 74310
rect 90940 74300 91060 74310
rect 91190 74300 91310 74310
rect 91440 74300 91560 74310
rect 91690 74300 91810 74310
rect 91940 74300 92060 74310
rect 92190 74300 92310 74310
rect 92440 74300 92560 74310
rect 92690 74300 92810 74310
rect 92940 74300 93060 74310
rect 93190 74300 93310 74310
rect 93440 74300 93560 74310
rect 93690 74300 93810 74310
rect 93940 74300 94060 74310
rect 94190 74300 94310 74310
rect 94440 74300 94560 74310
rect 94690 74300 94810 74310
rect 94940 74300 95060 74310
rect 95190 74300 95310 74310
rect 95440 74300 95560 74310
rect 95690 74300 95810 74310
rect 95940 74300 96060 74310
rect 96190 74300 96310 74310
rect 96440 74300 96560 74310
rect 96690 74300 96810 74310
rect 96940 74300 97060 74310
rect 97190 74300 97310 74310
rect 97440 74300 97560 74310
rect 97690 74300 97810 74310
rect 97940 74300 98060 74310
rect 98190 74300 98310 74310
rect 98440 74300 98560 74310
rect 98690 74300 98810 74310
rect 98940 74300 99060 74310
rect 99190 74300 99310 74310
rect 99440 74300 99560 74310
rect 99690 74300 99810 74310
rect 99940 74300 100060 74310
rect 100190 74300 100310 74310
rect 100440 74300 100560 74310
rect 100690 74300 100810 74310
rect 100940 74300 101060 74310
rect 101190 74300 101310 74310
rect 101440 74300 101560 74310
rect 101690 74300 101810 74310
rect 101940 74300 102060 74310
rect 102190 74300 102310 74310
rect 102440 74300 102560 74310
rect 102690 74300 102810 74310
rect 102940 74300 103060 74310
rect 103190 74300 103310 74310
rect 103440 74300 103560 74310
rect 103690 74300 103810 74310
rect 103940 74300 104060 74310
rect 104190 74300 104310 74310
rect 104440 74300 104560 74310
rect 104690 74300 104810 74310
rect 104940 74300 105060 74310
rect 105190 74300 105310 74310
rect 105440 74300 105560 74310
rect 105690 74300 105810 74310
rect 105940 74300 106060 74310
rect 106190 74300 106310 74310
rect 106440 74300 106560 74310
rect 106690 74300 106810 74310
rect 106940 74300 107060 74310
rect 107190 74300 107310 74310
rect 107440 74300 107560 74310
rect 107690 74300 107810 74310
rect 107940 74300 108060 74310
rect 108190 74300 108310 74310
rect 108440 74300 108560 74310
rect 108690 74300 108810 74310
rect 108940 74300 109060 74310
rect 109190 74300 109310 74310
rect 109440 74300 109560 74310
rect 109690 74300 109810 74310
rect 109940 74300 110060 74310
rect 110190 74300 110310 74310
rect 110440 74300 110560 74310
rect 110690 74300 110810 74310
rect 110940 74300 111060 74310
rect 111190 74300 111310 74310
rect 111440 74300 111560 74310
rect 111690 74300 111810 74310
rect 111940 74300 112060 74310
rect 112190 74300 112310 74310
rect 112440 74300 112560 74310
rect 112690 74300 112810 74310
rect 112940 74300 113060 74310
rect 113190 74300 113310 74310
rect 113440 74300 113560 74310
rect 113690 74300 113810 74310
rect 113940 74300 114060 74310
rect 114190 74300 114310 74310
rect 114440 74300 114560 74310
rect 114690 74300 114810 74310
rect 114940 74300 115060 74310
rect 115190 74300 115310 74310
rect 115440 74300 115560 74310
rect 115690 74300 115810 74310
rect 115940 74300 116000 74310
rect 89000 74200 116000 74300
rect 89000 74190 89060 74200
rect 89190 74190 89310 74200
rect 89440 74190 89560 74200
rect 89690 74190 89810 74200
rect 89940 74190 90060 74200
rect 90190 74190 90310 74200
rect 90440 74190 90560 74200
rect 90690 74190 90810 74200
rect 90940 74190 91060 74200
rect 91190 74190 91310 74200
rect 91440 74190 91560 74200
rect 91690 74190 91810 74200
rect 91940 74190 92060 74200
rect 92190 74190 92310 74200
rect 92440 74190 92560 74200
rect 92690 74190 92810 74200
rect 92940 74190 93060 74200
rect 93190 74190 93310 74200
rect 93440 74190 93560 74200
rect 93690 74190 93810 74200
rect 93940 74190 94060 74200
rect 94190 74190 94310 74200
rect 94440 74190 94560 74200
rect 94690 74190 94810 74200
rect 94940 74190 95060 74200
rect 95190 74190 95310 74200
rect 95440 74190 95560 74200
rect 95690 74190 95810 74200
rect 95940 74190 96060 74200
rect 96190 74190 96310 74200
rect 96440 74190 96560 74200
rect 96690 74190 96810 74200
rect 96940 74190 97060 74200
rect 97190 74190 97310 74200
rect 97440 74190 97560 74200
rect 97690 74190 97810 74200
rect 97940 74190 98060 74200
rect 98190 74190 98310 74200
rect 98440 74190 98560 74200
rect 98690 74190 98810 74200
rect 98940 74190 99060 74200
rect 99190 74190 99310 74200
rect 99440 74190 99560 74200
rect 99690 74190 99810 74200
rect 99940 74190 100060 74200
rect 100190 74190 100310 74200
rect 100440 74190 100560 74200
rect 100690 74190 100810 74200
rect 100940 74190 101060 74200
rect 101190 74190 101310 74200
rect 101440 74190 101560 74200
rect 101690 74190 101810 74200
rect 101940 74190 102060 74200
rect 102190 74190 102310 74200
rect 102440 74190 102560 74200
rect 102690 74190 102810 74200
rect 102940 74190 103060 74200
rect 103190 74190 103310 74200
rect 103440 74190 103560 74200
rect 103690 74190 103810 74200
rect 103940 74190 104060 74200
rect 104190 74190 104310 74200
rect 104440 74190 104560 74200
rect 104690 74190 104810 74200
rect 104940 74190 105060 74200
rect 105190 74190 105310 74200
rect 105440 74190 105560 74200
rect 105690 74190 105810 74200
rect 105940 74190 106060 74200
rect 106190 74190 106310 74200
rect 106440 74190 106560 74200
rect 106690 74190 106810 74200
rect 106940 74190 107060 74200
rect 107190 74190 107310 74200
rect 107440 74190 107560 74200
rect 107690 74190 107810 74200
rect 107940 74190 108060 74200
rect 108190 74190 108310 74200
rect 108440 74190 108560 74200
rect 108690 74190 108810 74200
rect 108940 74190 109060 74200
rect 109190 74190 109310 74200
rect 109440 74190 109560 74200
rect 109690 74190 109810 74200
rect 109940 74190 110060 74200
rect 110190 74190 110310 74200
rect 110440 74190 110560 74200
rect 110690 74190 110810 74200
rect 110940 74190 111060 74200
rect 111190 74190 111310 74200
rect 111440 74190 111560 74200
rect 111690 74190 111810 74200
rect 111940 74190 112060 74200
rect 112190 74190 112310 74200
rect 112440 74190 112560 74200
rect 112690 74190 112810 74200
rect 112940 74190 113060 74200
rect 113190 74190 113310 74200
rect 113440 74190 113560 74200
rect 113690 74190 113810 74200
rect 113940 74190 114060 74200
rect 114190 74190 114310 74200
rect 114440 74190 114560 74200
rect 114690 74190 114810 74200
rect 114940 74190 115060 74200
rect 115190 74190 115310 74200
rect 115440 74190 115560 74200
rect 115690 74190 115810 74200
rect 115940 74190 116000 74200
rect 89000 74060 89050 74190
rect 89200 74060 89300 74190
rect 89450 74060 89550 74190
rect 89700 74060 89800 74190
rect 89950 74060 90050 74190
rect 90200 74060 90300 74190
rect 90450 74060 90550 74190
rect 90700 74060 90800 74190
rect 90950 74060 91050 74190
rect 91200 74060 91300 74190
rect 91450 74060 91550 74190
rect 91700 74060 91800 74190
rect 91950 74060 92050 74190
rect 92200 74060 92300 74190
rect 92450 74060 92550 74190
rect 92700 74060 92800 74190
rect 92950 74060 93050 74190
rect 93200 74060 93300 74190
rect 93450 74060 93550 74190
rect 93700 74060 93800 74190
rect 93950 74060 94050 74190
rect 94200 74060 94300 74190
rect 94450 74060 94550 74190
rect 94700 74060 94800 74190
rect 94950 74060 95050 74190
rect 95200 74060 95300 74190
rect 95450 74060 95550 74190
rect 95700 74060 95800 74190
rect 95950 74060 96050 74190
rect 96200 74060 96300 74190
rect 96450 74060 96550 74190
rect 96700 74060 96800 74190
rect 96950 74060 97050 74190
rect 97200 74060 97300 74190
rect 97450 74060 97550 74190
rect 97700 74060 97800 74190
rect 97950 74060 98050 74190
rect 98200 74060 98300 74190
rect 98450 74060 98550 74190
rect 98700 74060 98800 74190
rect 98950 74060 99050 74190
rect 99200 74060 99300 74190
rect 99450 74060 99550 74190
rect 99700 74060 99800 74190
rect 99950 74060 100050 74190
rect 100200 74060 100300 74190
rect 100450 74060 100550 74190
rect 100700 74060 100800 74190
rect 100950 74060 101050 74190
rect 101200 74060 101300 74190
rect 101450 74060 101550 74190
rect 101700 74060 101800 74190
rect 101950 74060 102050 74190
rect 102200 74060 102300 74190
rect 102450 74060 102550 74190
rect 102700 74060 102800 74190
rect 102950 74060 103050 74190
rect 103200 74060 103300 74190
rect 103450 74060 103550 74190
rect 103700 74060 103800 74190
rect 103950 74060 104050 74190
rect 104200 74060 104300 74190
rect 104450 74060 104550 74190
rect 104700 74060 104800 74190
rect 104950 74060 105050 74190
rect 105200 74060 105300 74190
rect 105450 74060 105550 74190
rect 105700 74060 105800 74190
rect 105950 74060 106050 74190
rect 106200 74060 106300 74190
rect 106450 74060 106550 74190
rect 106700 74060 106800 74190
rect 106950 74060 107050 74190
rect 107200 74060 107300 74190
rect 107450 74060 107550 74190
rect 107700 74060 107800 74190
rect 107950 74060 108050 74190
rect 108200 74060 108300 74190
rect 108450 74060 108550 74190
rect 108700 74060 108800 74190
rect 108950 74060 109050 74190
rect 109200 74060 109300 74190
rect 109450 74060 109550 74190
rect 109700 74060 109800 74190
rect 109950 74060 110050 74190
rect 110200 74060 110300 74190
rect 110450 74060 110550 74190
rect 110700 74060 110800 74190
rect 110950 74060 111050 74190
rect 111200 74060 111300 74190
rect 111450 74060 111550 74190
rect 111700 74060 111800 74190
rect 111950 74060 112050 74190
rect 112200 74060 112300 74190
rect 112450 74060 112550 74190
rect 112700 74060 112800 74190
rect 112950 74060 113050 74190
rect 113200 74060 113300 74190
rect 113450 74060 113550 74190
rect 113700 74060 113800 74190
rect 113950 74060 114050 74190
rect 114200 74060 114300 74190
rect 114450 74060 114550 74190
rect 114700 74060 114800 74190
rect 114950 74060 115050 74190
rect 115200 74060 115300 74190
rect 115450 74060 115550 74190
rect 115700 74060 115800 74190
rect 115950 74060 116000 74190
rect 89000 74050 89060 74060
rect 89190 74050 89310 74060
rect 89440 74050 89560 74060
rect 89690 74050 89810 74060
rect 89940 74050 90060 74060
rect 90190 74050 90310 74060
rect 90440 74050 90560 74060
rect 90690 74050 90810 74060
rect 90940 74050 91060 74060
rect 91190 74050 91310 74060
rect 91440 74050 91560 74060
rect 91690 74050 91810 74060
rect 91940 74050 92060 74060
rect 92190 74050 92310 74060
rect 92440 74050 92560 74060
rect 92690 74050 92810 74060
rect 92940 74050 93060 74060
rect 93190 74050 93310 74060
rect 93440 74050 93560 74060
rect 93690 74050 93810 74060
rect 93940 74050 94060 74060
rect 94190 74050 94310 74060
rect 94440 74050 94560 74060
rect 94690 74050 94810 74060
rect 94940 74050 95060 74060
rect 95190 74050 95310 74060
rect 95440 74050 95560 74060
rect 95690 74050 95810 74060
rect 95940 74050 96060 74060
rect 96190 74050 96310 74060
rect 96440 74050 96560 74060
rect 96690 74050 96810 74060
rect 96940 74050 97060 74060
rect 97190 74050 97310 74060
rect 97440 74050 97560 74060
rect 97690 74050 97810 74060
rect 97940 74050 98060 74060
rect 98190 74050 98310 74060
rect 98440 74050 98560 74060
rect 98690 74050 98810 74060
rect 98940 74050 99060 74060
rect 99190 74050 99310 74060
rect 99440 74050 99560 74060
rect 99690 74050 99810 74060
rect 99940 74050 100060 74060
rect 100190 74050 100310 74060
rect 100440 74050 100560 74060
rect 100690 74050 100810 74060
rect 100940 74050 101060 74060
rect 101190 74050 101310 74060
rect 101440 74050 101560 74060
rect 101690 74050 101810 74060
rect 101940 74050 102060 74060
rect 102190 74050 102310 74060
rect 102440 74050 102560 74060
rect 102690 74050 102810 74060
rect 102940 74050 103060 74060
rect 103190 74050 103310 74060
rect 103440 74050 103560 74060
rect 103690 74050 103810 74060
rect 103940 74050 104060 74060
rect 104190 74050 104310 74060
rect 104440 74050 104560 74060
rect 104690 74050 104810 74060
rect 104940 74050 105060 74060
rect 105190 74050 105310 74060
rect 105440 74050 105560 74060
rect 105690 74050 105810 74060
rect 105940 74050 106060 74060
rect 106190 74050 106310 74060
rect 106440 74050 106560 74060
rect 106690 74050 106810 74060
rect 106940 74050 107060 74060
rect 107190 74050 107310 74060
rect 107440 74050 107560 74060
rect 107690 74050 107810 74060
rect 107940 74050 108060 74060
rect 108190 74050 108310 74060
rect 108440 74050 108560 74060
rect 108690 74050 108810 74060
rect 108940 74050 109060 74060
rect 109190 74050 109310 74060
rect 109440 74050 109560 74060
rect 109690 74050 109810 74060
rect 109940 74050 110060 74060
rect 110190 74050 110310 74060
rect 110440 74050 110560 74060
rect 110690 74050 110810 74060
rect 110940 74050 111060 74060
rect 111190 74050 111310 74060
rect 111440 74050 111560 74060
rect 111690 74050 111810 74060
rect 111940 74050 112060 74060
rect 112190 74050 112310 74060
rect 112440 74050 112560 74060
rect 112690 74050 112810 74060
rect 112940 74050 113060 74060
rect 113190 74050 113310 74060
rect 113440 74050 113560 74060
rect 113690 74050 113810 74060
rect 113940 74050 114060 74060
rect 114190 74050 114310 74060
rect 114440 74050 114560 74060
rect 114690 74050 114810 74060
rect 114940 74050 115060 74060
rect 115190 74050 115310 74060
rect 115440 74050 115560 74060
rect 115690 74050 115810 74060
rect 115940 74050 116000 74060
rect 89000 73950 116000 74050
rect 89000 73940 89060 73950
rect 89190 73940 89310 73950
rect 89440 73940 89560 73950
rect 89690 73940 89810 73950
rect 89940 73940 90060 73950
rect 90190 73940 90310 73950
rect 90440 73940 90560 73950
rect 90690 73940 90810 73950
rect 90940 73940 91060 73950
rect 91190 73940 91310 73950
rect 91440 73940 91560 73950
rect 91690 73940 91810 73950
rect 91940 73940 92060 73950
rect 92190 73940 92310 73950
rect 92440 73940 92560 73950
rect 92690 73940 92810 73950
rect 92940 73940 93060 73950
rect 93190 73940 93310 73950
rect 93440 73940 93560 73950
rect 93690 73940 93810 73950
rect 93940 73940 94060 73950
rect 94190 73940 94310 73950
rect 94440 73940 94560 73950
rect 94690 73940 94810 73950
rect 94940 73940 95060 73950
rect 95190 73940 95310 73950
rect 95440 73940 95560 73950
rect 95690 73940 95810 73950
rect 95940 73940 96060 73950
rect 96190 73940 96310 73950
rect 96440 73940 96560 73950
rect 96690 73940 96810 73950
rect 96940 73940 97060 73950
rect 97190 73940 97310 73950
rect 97440 73940 97560 73950
rect 97690 73940 97810 73950
rect 97940 73940 98060 73950
rect 98190 73940 98310 73950
rect 98440 73940 98560 73950
rect 98690 73940 98810 73950
rect 98940 73940 99060 73950
rect 99190 73940 99310 73950
rect 99440 73940 99560 73950
rect 99690 73940 99810 73950
rect 99940 73940 100060 73950
rect 100190 73940 100310 73950
rect 100440 73940 100560 73950
rect 100690 73940 100810 73950
rect 100940 73940 101060 73950
rect 101190 73940 101310 73950
rect 101440 73940 101560 73950
rect 101690 73940 101810 73950
rect 101940 73940 102060 73950
rect 102190 73940 102310 73950
rect 102440 73940 102560 73950
rect 102690 73940 102810 73950
rect 102940 73940 103060 73950
rect 103190 73940 103310 73950
rect 103440 73940 103560 73950
rect 103690 73940 103810 73950
rect 103940 73940 104060 73950
rect 104190 73940 104310 73950
rect 104440 73940 104560 73950
rect 104690 73940 104810 73950
rect 104940 73940 105060 73950
rect 105190 73940 105310 73950
rect 105440 73940 105560 73950
rect 105690 73940 105810 73950
rect 105940 73940 106060 73950
rect 106190 73940 106310 73950
rect 106440 73940 106560 73950
rect 106690 73940 106810 73950
rect 106940 73940 107060 73950
rect 107190 73940 107310 73950
rect 107440 73940 107560 73950
rect 107690 73940 107810 73950
rect 107940 73940 108060 73950
rect 108190 73940 108310 73950
rect 108440 73940 108560 73950
rect 108690 73940 108810 73950
rect 108940 73940 109060 73950
rect 109190 73940 109310 73950
rect 109440 73940 109560 73950
rect 109690 73940 109810 73950
rect 109940 73940 110060 73950
rect 110190 73940 110310 73950
rect 110440 73940 110560 73950
rect 110690 73940 110810 73950
rect 110940 73940 111060 73950
rect 111190 73940 111310 73950
rect 111440 73940 111560 73950
rect 111690 73940 111810 73950
rect 111940 73940 112060 73950
rect 112190 73940 112310 73950
rect 112440 73940 112560 73950
rect 112690 73940 112810 73950
rect 112940 73940 113060 73950
rect 113190 73940 113310 73950
rect 113440 73940 113560 73950
rect 113690 73940 113810 73950
rect 113940 73940 114060 73950
rect 114190 73940 114310 73950
rect 114440 73940 114560 73950
rect 114690 73940 114810 73950
rect 114940 73940 115060 73950
rect 115190 73940 115310 73950
rect 115440 73940 115560 73950
rect 115690 73940 115810 73950
rect 115940 73940 116000 73950
rect 89000 73810 89050 73940
rect 89200 73810 89300 73940
rect 89450 73810 89550 73940
rect 89700 73810 89800 73940
rect 89950 73810 90050 73940
rect 90200 73810 90300 73940
rect 90450 73810 90550 73940
rect 90700 73810 90800 73940
rect 90950 73810 91050 73940
rect 91200 73810 91300 73940
rect 91450 73810 91550 73940
rect 91700 73810 91800 73940
rect 91950 73810 92050 73940
rect 92200 73810 92300 73940
rect 92450 73810 92550 73940
rect 92700 73810 92800 73940
rect 92950 73810 93050 73940
rect 93200 73810 93300 73940
rect 93450 73810 93550 73940
rect 93700 73810 93800 73940
rect 93950 73810 94050 73940
rect 94200 73810 94300 73940
rect 94450 73810 94550 73940
rect 94700 73810 94800 73940
rect 94950 73810 95050 73940
rect 95200 73810 95300 73940
rect 95450 73810 95550 73940
rect 95700 73810 95800 73940
rect 95950 73810 96050 73940
rect 96200 73810 96300 73940
rect 96450 73810 96550 73940
rect 96700 73810 96800 73940
rect 96950 73810 97050 73940
rect 97200 73810 97300 73940
rect 97450 73810 97550 73940
rect 97700 73810 97800 73940
rect 97950 73810 98050 73940
rect 98200 73810 98300 73940
rect 98450 73810 98550 73940
rect 98700 73810 98800 73940
rect 98950 73810 99050 73940
rect 99200 73810 99300 73940
rect 99450 73810 99550 73940
rect 99700 73810 99800 73940
rect 99950 73810 100050 73940
rect 100200 73810 100300 73940
rect 100450 73810 100550 73940
rect 100700 73810 100800 73940
rect 100950 73810 101050 73940
rect 101200 73810 101300 73940
rect 101450 73810 101550 73940
rect 101700 73810 101800 73940
rect 101950 73810 102050 73940
rect 102200 73810 102300 73940
rect 102450 73810 102550 73940
rect 102700 73810 102800 73940
rect 102950 73810 103050 73940
rect 103200 73810 103300 73940
rect 103450 73810 103550 73940
rect 103700 73810 103800 73940
rect 103950 73810 104050 73940
rect 104200 73810 104300 73940
rect 104450 73810 104550 73940
rect 104700 73810 104800 73940
rect 104950 73810 105050 73940
rect 105200 73810 105300 73940
rect 105450 73810 105550 73940
rect 105700 73810 105800 73940
rect 105950 73810 106050 73940
rect 106200 73810 106300 73940
rect 106450 73810 106550 73940
rect 106700 73810 106800 73940
rect 106950 73810 107050 73940
rect 107200 73810 107300 73940
rect 107450 73810 107550 73940
rect 107700 73810 107800 73940
rect 107950 73810 108050 73940
rect 108200 73810 108300 73940
rect 108450 73810 108550 73940
rect 108700 73810 108800 73940
rect 108950 73810 109050 73940
rect 109200 73810 109300 73940
rect 109450 73810 109550 73940
rect 109700 73810 109800 73940
rect 109950 73810 110050 73940
rect 110200 73810 110300 73940
rect 110450 73810 110550 73940
rect 110700 73810 110800 73940
rect 110950 73810 111050 73940
rect 111200 73810 111300 73940
rect 111450 73810 111550 73940
rect 111700 73810 111800 73940
rect 111950 73810 112050 73940
rect 112200 73810 112300 73940
rect 112450 73810 112550 73940
rect 112700 73810 112800 73940
rect 112950 73810 113050 73940
rect 113200 73810 113300 73940
rect 113450 73810 113550 73940
rect 113700 73810 113800 73940
rect 113950 73810 114050 73940
rect 114200 73810 114300 73940
rect 114450 73810 114550 73940
rect 114700 73810 114800 73940
rect 114950 73810 115050 73940
rect 115200 73810 115300 73940
rect 115450 73810 115550 73940
rect 115700 73810 115800 73940
rect 115950 73810 116000 73940
rect 89000 73800 89060 73810
rect 89190 73800 89310 73810
rect 89440 73800 89560 73810
rect 89690 73800 89810 73810
rect 89940 73800 90060 73810
rect 90190 73800 90310 73810
rect 90440 73800 90560 73810
rect 90690 73800 90810 73810
rect 90940 73800 91060 73810
rect 91190 73800 91310 73810
rect 91440 73800 91560 73810
rect 91690 73800 91810 73810
rect 91940 73800 92060 73810
rect 92190 73800 92310 73810
rect 92440 73800 92560 73810
rect 92690 73800 92810 73810
rect 92940 73800 93060 73810
rect 93190 73800 93310 73810
rect 93440 73800 93560 73810
rect 93690 73800 93810 73810
rect 93940 73800 94060 73810
rect 94190 73800 94310 73810
rect 94440 73800 94560 73810
rect 94690 73800 94810 73810
rect 94940 73800 95060 73810
rect 95190 73800 95310 73810
rect 95440 73800 95560 73810
rect 95690 73800 95810 73810
rect 95940 73800 96060 73810
rect 96190 73800 96310 73810
rect 96440 73800 96560 73810
rect 96690 73800 96810 73810
rect 96940 73800 97060 73810
rect 97190 73800 97310 73810
rect 97440 73800 97560 73810
rect 97690 73800 97810 73810
rect 97940 73800 98060 73810
rect 98190 73800 98310 73810
rect 98440 73800 98560 73810
rect 98690 73800 98810 73810
rect 98940 73800 99060 73810
rect 99190 73800 99310 73810
rect 99440 73800 99560 73810
rect 99690 73800 99810 73810
rect 99940 73800 100060 73810
rect 100190 73800 100310 73810
rect 100440 73800 100560 73810
rect 100690 73800 100810 73810
rect 100940 73800 101060 73810
rect 101190 73800 101310 73810
rect 101440 73800 101560 73810
rect 101690 73800 101810 73810
rect 101940 73800 102060 73810
rect 102190 73800 102310 73810
rect 102440 73800 102560 73810
rect 102690 73800 102810 73810
rect 102940 73800 103060 73810
rect 103190 73800 103310 73810
rect 103440 73800 103560 73810
rect 103690 73800 103810 73810
rect 103940 73800 104060 73810
rect 104190 73800 104310 73810
rect 104440 73800 104560 73810
rect 104690 73800 104810 73810
rect 104940 73800 105060 73810
rect 105190 73800 105310 73810
rect 105440 73800 105560 73810
rect 105690 73800 105810 73810
rect 105940 73800 106060 73810
rect 106190 73800 106310 73810
rect 106440 73800 106560 73810
rect 106690 73800 106810 73810
rect 106940 73800 107060 73810
rect 107190 73800 107310 73810
rect 107440 73800 107560 73810
rect 107690 73800 107810 73810
rect 107940 73800 108060 73810
rect 108190 73800 108310 73810
rect 108440 73800 108560 73810
rect 108690 73800 108810 73810
rect 108940 73800 109060 73810
rect 109190 73800 109310 73810
rect 109440 73800 109560 73810
rect 109690 73800 109810 73810
rect 109940 73800 110060 73810
rect 110190 73800 110310 73810
rect 110440 73800 110560 73810
rect 110690 73800 110810 73810
rect 110940 73800 111060 73810
rect 111190 73800 111310 73810
rect 111440 73800 111560 73810
rect 111690 73800 111810 73810
rect 111940 73800 112060 73810
rect 112190 73800 112310 73810
rect 112440 73800 112560 73810
rect 112690 73800 112810 73810
rect 112940 73800 113060 73810
rect 113190 73800 113310 73810
rect 113440 73800 113560 73810
rect 113690 73800 113810 73810
rect 113940 73800 114060 73810
rect 114190 73800 114310 73810
rect 114440 73800 114560 73810
rect 114690 73800 114810 73810
rect 114940 73800 115060 73810
rect 115190 73800 115310 73810
rect 115440 73800 115560 73810
rect 115690 73800 115810 73810
rect 115940 73800 116000 73810
rect 89000 73700 116000 73800
rect 89000 73690 89060 73700
rect 89190 73690 89310 73700
rect 89440 73690 89560 73700
rect 89690 73690 89810 73700
rect 89940 73690 90060 73700
rect 90190 73690 90310 73700
rect 90440 73690 90560 73700
rect 90690 73690 90810 73700
rect 90940 73690 91060 73700
rect 91190 73690 91310 73700
rect 91440 73690 91560 73700
rect 91690 73690 91810 73700
rect 91940 73690 92060 73700
rect 92190 73690 92310 73700
rect 92440 73690 92560 73700
rect 92690 73690 92810 73700
rect 92940 73690 93060 73700
rect 93190 73690 93310 73700
rect 93440 73690 93560 73700
rect 93690 73690 93810 73700
rect 93940 73690 94060 73700
rect 94190 73690 94310 73700
rect 94440 73690 94560 73700
rect 94690 73690 94810 73700
rect 94940 73690 95060 73700
rect 95190 73690 95310 73700
rect 95440 73690 95560 73700
rect 95690 73690 95810 73700
rect 95940 73690 96060 73700
rect 96190 73690 96310 73700
rect 96440 73690 96560 73700
rect 96690 73690 96810 73700
rect 96940 73690 97060 73700
rect 97190 73690 97310 73700
rect 97440 73690 97560 73700
rect 97690 73690 97810 73700
rect 97940 73690 98060 73700
rect 98190 73690 98310 73700
rect 98440 73690 98560 73700
rect 98690 73690 98810 73700
rect 98940 73690 99060 73700
rect 99190 73690 99310 73700
rect 99440 73690 99560 73700
rect 99690 73690 99810 73700
rect 99940 73690 100060 73700
rect 100190 73690 100310 73700
rect 100440 73690 100560 73700
rect 100690 73690 100810 73700
rect 100940 73690 101060 73700
rect 101190 73690 101310 73700
rect 101440 73690 101560 73700
rect 101690 73690 101810 73700
rect 101940 73690 102060 73700
rect 102190 73690 102310 73700
rect 102440 73690 102560 73700
rect 102690 73690 102810 73700
rect 102940 73690 103060 73700
rect 103190 73690 103310 73700
rect 103440 73690 103560 73700
rect 103690 73690 103810 73700
rect 103940 73690 104060 73700
rect 104190 73690 104310 73700
rect 104440 73690 104560 73700
rect 104690 73690 104810 73700
rect 104940 73690 105060 73700
rect 105190 73690 105310 73700
rect 105440 73690 105560 73700
rect 105690 73690 105810 73700
rect 105940 73690 106060 73700
rect 106190 73690 106310 73700
rect 106440 73690 106560 73700
rect 106690 73690 106810 73700
rect 106940 73690 107060 73700
rect 107190 73690 107310 73700
rect 107440 73690 107560 73700
rect 107690 73690 107810 73700
rect 107940 73690 108060 73700
rect 108190 73690 108310 73700
rect 108440 73690 108560 73700
rect 108690 73690 108810 73700
rect 108940 73690 109060 73700
rect 109190 73690 109310 73700
rect 109440 73690 109560 73700
rect 109690 73690 109810 73700
rect 109940 73690 110060 73700
rect 110190 73690 110310 73700
rect 110440 73690 110560 73700
rect 110690 73690 110810 73700
rect 110940 73690 111060 73700
rect 111190 73690 111310 73700
rect 111440 73690 111560 73700
rect 111690 73690 111810 73700
rect 111940 73690 112060 73700
rect 112190 73690 112310 73700
rect 112440 73690 112560 73700
rect 112690 73690 112810 73700
rect 112940 73690 113060 73700
rect 113190 73690 113310 73700
rect 113440 73690 113560 73700
rect 113690 73690 113810 73700
rect 113940 73690 114060 73700
rect 114190 73690 114310 73700
rect 114440 73690 114560 73700
rect 114690 73690 114810 73700
rect 114940 73690 115060 73700
rect 115190 73690 115310 73700
rect 115440 73690 115560 73700
rect 115690 73690 115810 73700
rect 115940 73690 116000 73700
rect 89000 73560 89050 73690
rect 89200 73560 89300 73690
rect 89450 73560 89550 73690
rect 89700 73560 89800 73690
rect 89950 73560 90050 73690
rect 90200 73560 90300 73690
rect 90450 73560 90550 73690
rect 90700 73560 90800 73690
rect 90950 73560 91050 73690
rect 91200 73560 91300 73690
rect 91450 73560 91550 73690
rect 91700 73560 91800 73690
rect 91950 73560 92050 73690
rect 92200 73560 92300 73690
rect 92450 73560 92550 73690
rect 92700 73560 92800 73690
rect 92950 73560 93050 73690
rect 93200 73560 93300 73690
rect 93450 73560 93550 73690
rect 93700 73560 93800 73690
rect 93950 73560 94050 73690
rect 94200 73560 94300 73690
rect 94450 73560 94550 73690
rect 94700 73560 94800 73690
rect 94950 73560 95050 73690
rect 95200 73560 95300 73690
rect 95450 73560 95550 73690
rect 95700 73560 95800 73690
rect 95950 73560 96050 73690
rect 96200 73560 96300 73690
rect 96450 73560 96550 73690
rect 96700 73560 96800 73690
rect 96950 73560 97050 73690
rect 97200 73560 97300 73690
rect 97450 73560 97550 73690
rect 97700 73560 97800 73690
rect 97950 73560 98050 73690
rect 98200 73560 98300 73690
rect 98450 73560 98550 73690
rect 98700 73560 98800 73690
rect 98950 73560 99050 73690
rect 99200 73560 99300 73690
rect 99450 73560 99550 73690
rect 99700 73560 99800 73690
rect 99950 73560 100050 73690
rect 100200 73560 100300 73690
rect 100450 73560 100550 73690
rect 100700 73560 100800 73690
rect 100950 73560 101050 73690
rect 101200 73560 101300 73690
rect 101450 73560 101550 73690
rect 101700 73560 101800 73690
rect 101950 73560 102050 73690
rect 102200 73560 102300 73690
rect 102450 73560 102550 73690
rect 102700 73560 102800 73690
rect 102950 73560 103050 73690
rect 103200 73560 103300 73690
rect 103450 73560 103550 73690
rect 103700 73560 103800 73690
rect 103950 73560 104050 73690
rect 104200 73560 104300 73690
rect 104450 73560 104550 73690
rect 104700 73560 104800 73690
rect 104950 73560 105050 73690
rect 105200 73560 105300 73690
rect 105450 73560 105550 73690
rect 105700 73560 105800 73690
rect 105950 73560 106050 73690
rect 106200 73560 106300 73690
rect 106450 73560 106550 73690
rect 106700 73560 106800 73690
rect 106950 73560 107050 73690
rect 107200 73560 107300 73690
rect 107450 73560 107550 73690
rect 107700 73560 107800 73690
rect 107950 73560 108050 73690
rect 108200 73560 108300 73690
rect 108450 73560 108550 73690
rect 108700 73560 108800 73690
rect 108950 73560 109050 73690
rect 109200 73560 109300 73690
rect 109450 73560 109550 73690
rect 109700 73560 109800 73690
rect 109950 73560 110050 73690
rect 110200 73560 110300 73690
rect 110450 73560 110550 73690
rect 110700 73560 110800 73690
rect 110950 73560 111050 73690
rect 111200 73560 111300 73690
rect 111450 73560 111550 73690
rect 111700 73560 111800 73690
rect 111950 73560 112050 73690
rect 112200 73560 112300 73690
rect 112450 73560 112550 73690
rect 112700 73560 112800 73690
rect 112950 73560 113050 73690
rect 113200 73560 113300 73690
rect 113450 73560 113550 73690
rect 113700 73560 113800 73690
rect 113950 73560 114050 73690
rect 114200 73560 114300 73690
rect 114450 73560 114550 73690
rect 114700 73560 114800 73690
rect 114950 73560 115050 73690
rect 115200 73560 115300 73690
rect 115450 73560 115550 73690
rect 115700 73560 115800 73690
rect 115950 73560 116000 73690
rect 89000 73550 89060 73560
rect 89190 73550 89310 73560
rect 89440 73550 89560 73560
rect 89690 73550 89810 73560
rect 89940 73550 90060 73560
rect 90190 73550 90310 73560
rect 90440 73550 90560 73560
rect 90690 73550 90810 73560
rect 90940 73550 91060 73560
rect 91190 73550 91310 73560
rect 91440 73550 91560 73560
rect 91690 73550 91810 73560
rect 91940 73550 92060 73560
rect 92190 73550 92310 73560
rect 92440 73550 92560 73560
rect 92690 73550 92810 73560
rect 92940 73550 93060 73560
rect 93190 73550 93310 73560
rect 93440 73550 93560 73560
rect 93690 73550 93810 73560
rect 93940 73550 94060 73560
rect 94190 73550 94310 73560
rect 94440 73550 94560 73560
rect 94690 73550 94810 73560
rect 94940 73550 95060 73560
rect 95190 73550 95310 73560
rect 95440 73550 95560 73560
rect 95690 73550 95810 73560
rect 95940 73550 96060 73560
rect 96190 73550 96310 73560
rect 96440 73550 96560 73560
rect 96690 73550 96810 73560
rect 96940 73550 97060 73560
rect 97190 73550 97310 73560
rect 97440 73550 97560 73560
rect 97690 73550 97810 73560
rect 97940 73550 98060 73560
rect 98190 73550 98310 73560
rect 98440 73550 98560 73560
rect 98690 73550 98810 73560
rect 98940 73550 99060 73560
rect 99190 73550 99310 73560
rect 99440 73550 99560 73560
rect 99690 73550 99810 73560
rect 99940 73550 100060 73560
rect 100190 73550 100310 73560
rect 100440 73550 100560 73560
rect 100690 73550 100810 73560
rect 100940 73550 101060 73560
rect 101190 73550 101310 73560
rect 101440 73550 101560 73560
rect 101690 73550 101810 73560
rect 101940 73550 102060 73560
rect 102190 73550 102310 73560
rect 102440 73550 102560 73560
rect 102690 73550 102810 73560
rect 102940 73550 103060 73560
rect 103190 73550 103310 73560
rect 103440 73550 103560 73560
rect 103690 73550 103810 73560
rect 103940 73550 104060 73560
rect 104190 73550 104310 73560
rect 104440 73550 104560 73560
rect 104690 73550 104810 73560
rect 104940 73550 105060 73560
rect 105190 73550 105310 73560
rect 105440 73550 105560 73560
rect 105690 73550 105810 73560
rect 105940 73550 106060 73560
rect 106190 73550 106310 73560
rect 106440 73550 106560 73560
rect 106690 73550 106810 73560
rect 106940 73550 107060 73560
rect 107190 73550 107310 73560
rect 107440 73550 107560 73560
rect 107690 73550 107810 73560
rect 107940 73550 108060 73560
rect 108190 73550 108310 73560
rect 108440 73550 108560 73560
rect 108690 73550 108810 73560
rect 108940 73550 109060 73560
rect 109190 73550 109310 73560
rect 109440 73550 109560 73560
rect 109690 73550 109810 73560
rect 109940 73550 110060 73560
rect 110190 73550 110310 73560
rect 110440 73550 110560 73560
rect 110690 73550 110810 73560
rect 110940 73550 111060 73560
rect 111190 73550 111310 73560
rect 111440 73550 111560 73560
rect 111690 73550 111810 73560
rect 111940 73550 112060 73560
rect 112190 73550 112310 73560
rect 112440 73550 112560 73560
rect 112690 73550 112810 73560
rect 112940 73550 113060 73560
rect 113190 73550 113310 73560
rect 113440 73550 113560 73560
rect 113690 73550 113810 73560
rect 113940 73550 114060 73560
rect 114190 73550 114310 73560
rect 114440 73550 114560 73560
rect 114690 73550 114810 73560
rect 114940 73550 115060 73560
rect 115190 73550 115310 73560
rect 115440 73550 115560 73560
rect 115690 73550 115810 73560
rect 115940 73550 116000 73560
rect 89000 73450 116000 73550
rect 89000 73440 89060 73450
rect 89190 73440 89310 73450
rect 89440 73440 89560 73450
rect 89690 73440 89810 73450
rect 89940 73440 90060 73450
rect 90190 73440 90310 73450
rect 90440 73440 90560 73450
rect 90690 73440 90810 73450
rect 90940 73440 91060 73450
rect 91190 73440 91310 73450
rect 91440 73440 91560 73450
rect 91690 73440 91810 73450
rect 91940 73440 92060 73450
rect 92190 73440 92310 73450
rect 92440 73440 92560 73450
rect 92690 73440 92810 73450
rect 92940 73440 93060 73450
rect 93190 73440 93310 73450
rect 93440 73440 93560 73450
rect 93690 73440 93810 73450
rect 93940 73440 94060 73450
rect 94190 73440 94310 73450
rect 94440 73440 94560 73450
rect 94690 73440 94810 73450
rect 94940 73440 95060 73450
rect 95190 73440 95310 73450
rect 95440 73440 95560 73450
rect 95690 73440 95810 73450
rect 95940 73440 96060 73450
rect 96190 73440 96310 73450
rect 96440 73440 96560 73450
rect 96690 73440 96810 73450
rect 96940 73440 97060 73450
rect 97190 73440 97310 73450
rect 97440 73440 97560 73450
rect 97690 73440 97810 73450
rect 97940 73440 98060 73450
rect 98190 73440 98310 73450
rect 98440 73440 98560 73450
rect 98690 73440 98810 73450
rect 98940 73440 99060 73450
rect 99190 73440 99310 73450
rect 99440 73440 99560 73450
rect 99690 73440 99810 73450
rect 99940 73440 100060 73450
rect 100190 73440 100310 73450
rect 100440 73440 100560 73450
rect 100690 73440 100810 73450
rect 100940 73440 101060 73450
rect 101190 73440 101310 73450
rect 101440 73440 101560 73450
rect 101690 73440 101810 73450
rect 101940 73440 102060 73450
rect 102190 73440 102310 73450
rect 102440 73440 102560 73450
rect 102690 73440 102810 73450
rect 102940 73440 103060 73450
rect 103190 73440 103310 73450
rect 103440 73440 103560 73450
rect 103690 73440 103810 73450
rect 103940 73440 104060 73450
rect 104190 73440 104310 73450
rect 104440 73440 104560 73450
rect 104690 73440 104810 73450
rect 104940 73440 105060 73450
rect 105190 73440 105310 73450
rect 105440 73440 105560 73450
rect 105690 73440 105810 73450
rect 105940 73440 106060 73450
rect 106190 73440 106310 73450
rect 106440 73440 106560 73450
rect 106690 73440 106810 73450
rect 106940 73440 107060 73450
rect 107190 73440 107310 73450
rect 107440 73440 107560 73450
rect 107690 73440 107810 73450
rect 107940 73440 108060 73450
rect 108190 73440 108310 73450
rect 108440 73440 108560 73450
rect 108690 73440 108810 73450
rect 108940 73440 109060 73450
rect 109190 73440 109310 73450
rect 109440 73440 109560 73450
rect 109690 73440 109810 73450
rect 109940 73440 110060 73450
rect 110190 73440 110310 73450
rect 110440 73440 110560 73450
rect 110690 73440 110810 73450
rect 110940 73440 111060 73450
rect 111190 73440 111310 73450
rect 111440 73440 111560 73450
rect 111690 73440 111810 73450
rect 111940 73440 112060 73450
rect 112190 73440 112310 73450
rect 112440 73440 112560 73450
rect 112690 73440 112810 73450
rect 112940 73440 113060 73450
rect 113190 73440 113310 73450
rect 113440 73440 113560 73450
rect 113690 73440 113810 73450
rect 113940 73440 114060 73450
rect 114190 73440 114310 73450
rect 114440 73440 114560 73450
rect 114690 73440 114810 73450
rect 114940 73440 115060 73450
rect 115190 73440 115310 73450
rect 115440 73440 115560 73450
rect 115690 73440 115810 73450
rect 115940 73440 116000 73450
rect 89000 73310 89050 73440
rect 89200 73310 89300 73440
rect 89450 73310 89550 73440
rect 89700 73310 89800 73440
rect 89950 73310 90050 73440
rect 90200 73310 90300 73440
rect 90450 73310 90550 73440
rect 90700 73310 90800 73440
rect 90950 73310 91050 73440
rect 91200 73310 91300 73440
rect 91450 73310 91550 73440
rect 91700 73310 91800 73440
rect 91950 73310 92050 73440
rect 92200 73310 92300 73440
rect 92450 73310 92550 73440
rect 92700 73310 92800 73440
rect 92950 73310 93050 73440
rect 93200 73310 93300 73440
rect 93450 73310 93550 73440
rect 93700 73310 93800 73440
rect 93950 73310 94050 73440
rect 94200 73310 94300 73440
rect 94450 73310 94550 73440
rect 94700 73310 94800 73440
rect 94950 73310 95050 73440
rect 95200 73310 95300 73440
rect 95450 73310 95550 73440
rect 95700 73310 95800 73440
rect 95950 73310 96050 73440
rect 96200 73310 96300 73440
rect 96450 73310 96550 73440
rect 96700 73310 96800 73440
rect 96950 73310 97050 73440
rect 97200 73310 97300 73440
rect 97450 73310 97550 73440
rect 97700 73310 97800 73440
rect 97950 73310 98050 73440
rect 98200 73310 98300 73440
rect 98450 73310 98550 73440
rect 98700 73310 98800 73440
rect 98950 73310 99050 73440
rect 99200 73310 99300 73440
rect 99450 73310 99550 73440
rect 99700 73310 99800 73440
rect 99950 73310 100050 73440
rect 100200 73310 100300 73440
rect 100450 73310 100550 73440
rect 100700 73310 100800 73440
rect 100950 73310 101050 73440
rect 101200 73310 101300 73440
rect 101450 73310 101550 73440
rect 101700 73310 101800 73440
rect 101950 73310 102050 73440
rect 102200 73310 102300 73440
rect 102450 73310 102550 73440
rect 102700 73310 102800 73440
rect 102950 73310 103050 73440
rect 103200 73310 103300 73440
rect 103450 73310 103550 73440
rect 103700 73310 103800 73440
rect 103950 73310 104050 73440
rect 104200 73310 104300 73440
rect 104450 73310 104550 73440
rect 104700 73310 104800 73440
rect 104950 73310 105050 73440
rect 105200 73310 105300 73440
rect 105450 73310 105550 73440
rect 105700 73310 105800 73440
rect 105950 73310 106050 73440
rect 106200 73310 106300 73440
rect 106450 73310 106550 73440
rect 106700 73310 106800 73440
rect 106950 73310 107050 73440
rect 107200 73310 107300 73440
rect 107450 73310 107550 73440
rect 107700 73310 107800 73440
rect 107950 73310 108050 73440
rect 108200 73310 108300 73440
rect 108450 73310 108550 73440
rect 108700 73310 108800 73440
rect 108950 73310 109050 73440
rect 109200 73310 109300 73440
rect 109450 73310 109550 73440
rect 109700 73310 109800 73440
rect 109950 73310 110050 73440
rect 110200 73310 110300 73440
rect 110450 73310 110550 73440
rect 110700 73310 110800 73440
rect 110950 73310 111050 73440
rect 111200 73310 111300 73440
rect 111450 73310 111550 73440
rect 111700 73310 111800 73440
rect 111950 73310 112050 73440
rect 112200 73310 112300 73440
rect 112450 73310 112550 73440
rect 112700 73310 112800 73440
rect 112950 73310 113050 73440
rect 113200 73310 113300 73440
rect 113450 73310 113550 73440
rect 113700 73310 113800 73440
rect 113950 73310 114050 73440
rect 114200 73310 114300 73440
rect 114450 73310 114550 73440
rect 114700 73310 114800 73440
rect 114950 73310 115050 73440
rect 115200 73310 115300 73440
rect 115450 73310 115550 73440
rect 115700 73310 115800 73440
rect 115950 73310 116000 73440
rect 89000 73300 89060 73310
rect 89190 73300 89310 73310
rect 89440 73300 89560 73310
rect 89690 73300 89810 73310
rect 89940 73300 90060 73310
rect 90190 73300 90310 73310
rect 90440 73300 90560 73310
rect 90690 73300 90810 73310
rect 90940 73300 91060 73310
rect 91190 73300 91310 73310
rect 91440 73300 91560 73310
rect 91690 73300 91810 73310
rect 91940 73300 92060 73310
rect 92190 73300 92310 73310
rect 92440 73300 92560 73310
rect 92690 73300 92810 73310
rect 92940 73300 93060 73310
rect 93190 73300 93310 73310
rect 93440 73300 93560 73310
rect 93690 73300 93810 73310
rect 93940 73300 94060 73310
rect 94190 73300 94310 73310
rect 94440 73300 94560 73310
rect 94690 73300 94810 73310
rect 94940 73300 95060 73310
rect 95190 73300 95310 73310
rect 95440 73300 95560 73310
rect 95690 73300 95810 73310
rect 95940 73300 96060 73310
rect 96190 73300 96310 73310
rect 96440 73300 96560 73310
rect 96690 73300 96810 73310
rect 96940 73300 97060 73310
rect 97190 73300 97310 73310
rect 97440 73300 97560 73310
rect 97690 73300 97810 73310
rect 97940 73300 98060 73310
rect 98190 73300 98310 73310
rect 98440 73300 98560 73310
rect 98690 73300 98810 73310
rect 98940 73300 99060 73310
rect 99190 73300 99310 73310
rect 99440 73300 99560 73310
rect 99690 73300 99810 73310
rect 99940 73300 100060 73310
rect 100190 73300 100310 73310
rect 100440 73300 100560 73310
rect 100690 73300 100810 73310
rect 100940 73300 101060 73310
rect 101190 73300 101310 73310
rect 101440 73300 101560 73310
rect 101690 73300 101810 73310
rect 101940 73300 102060 73310
rect 102190 73300 102310 73310
rect 102440 73300 102560 73310
rect 102690 73300 102810 73310
rect 102940 73300 103060 73310
rect 103190 73300 103310 73310
rect 103440 73300 103560 73310
rect 103690 73300 103810 73310
rect 103940 73300 104060 73310
rect 104190 73300 104310 73310
rect 104440 73300 104560 73310
rect 104690 73300 104810 73310
rect 104940 73300 105060 73310
rect 105190 73300 105310 73310
rect 105440 73300 105560 73310
rect 105690 73300 105810 73310
rect 105940 73300 106060 73310
rect 106190 73300 106310 73310
rect 106440 73300 106560 73310
rect 106690 73300 106810 73310
rect 106940 73300 107060 73310
rect 107190 73300 107310 73310
rect 107440 73300 107560 73310
rect 107690 73300 107810 73310
rect 107940 73300 108060 73310
rect 108190 73300 108310 73310
rect 108440 73300 108560 73310
rect 108690 73300 108810 73310
rect 108940 73300 109060 73310
rect 109190 73300 109310 73310
rect 109440 73300 109560 73310
rect 109690 73300 109810 73310
rect 109940 73300 110060 73310
rect 110190 73300 110310 73310
rect 110440 73300 110560 73310
rect 110690 73300 110810 73310
rect 110940 73300 111060 73310
rect 111190 73300 111310 73310
rect 111440 73300 111560 73310
rect 111690 73300 111810 73310
rect 111940 73300 112060 73310
rect 112190 73300 112310 73310
rect 112440 73300 112560 73310
rect 112690 73300 112810 73310
rect 112940 73300 113060 73310
rect 113190 73300 113310 73310
rect 113440 73300 113560 73310
rect 113690 73300 113810 73310
rect 113940 73300 114060 73310
rect 114190 73300 114310 73310
rect 114440 73300 114560 73310
rect 114690 73300 114810 73310
rect 114940 73300 115060 73310
rect 115190 73300 115310 73310
rect 115440 73300 115560 73310
rect 115690 73300 115810 73310
rect 115940 73300 116000 73310
rect 89000 73200 116000 73300
rect 89000 73190 89060 73200
rect 89190 73190 89310 73200
rect 89440 73190 89560 73200
rect 89690 73190 89810 73200
rect 89940 73190 90060 73200
rect 90190 73190 90310 73200
rect 90440 73190 90560 73200
rect 90690 73190 90810 73200
rect 90940 73190 91060 73200
rect 91190 73190 91310 73200
rect 91440 73190 91560 73200
rect 91690 73190 91810 73200
rect 91940 73190 92060 73200
rect 92190 73190 92310 73200
rect 92440 73190 92560 73200
rect 92690 73190 92810 73200
rect 92940 73190 93060 73200
rect 93190 73190 93310 73200
rect 93440 73190 93560 73200
rect 93690 73190 93810 73200
rect 93940 73190 94060 73200
rect 94190 73190 94310 73200
rect 94440 73190 94560 73200
rect 94690 73190 94810 73200
rect 94940 73190 95060 73200
rect 95190 73190 95310 73200
rect 95440 73190 95560 73200
rect 95690 73190 95810 73200
rect 95940 73190 96060 73200
rect 96190 73190 96310 73200
rect 96440 73190 96560 73200
rect 96690 73190 96810 73200
rect 96940 73190 97060 73200
rect 97190 73190 97310 73200
rect 97440 73190 97560 73200
rect 97690 73190 97810 73200
rect 97940 73190 98060 73200
rect 98190 73190 98310 73200
rect 98440 73190 98560 73200
rect 98690 73190 98810 73200
rect 98940 73190 99060 73200
rect 99190 73190 99310 73200
rect 99440 73190 99560 73200
rect 99690 73190 99810 73200
rect 99940 73190 100060 73200
rect 100190 73190 100310 73200
rect 100440 73190 100560 73200
rect 100690 73190 100810 73200
rect 100940 73190 101060 73200
rect 101190 73190 101310 73200
rect 101440 73190 101560 73200
rect 101690 73190 101810 73200
rect 101940 73190 102060 73200
rect 102190 73190 102310 73200
rect 102440 73190 102560 73200
rect 102690 73190 102810 73200
rect 102940 73190 103060 73200
rect 103190 73190 103310 73200
rect 103440 73190 103560 73200
rect 103690 73190 103810 73200
rect 103940 73190 104060 73200
rect 104190 73190 104310 73200
rect 104440 73190 104560 73200
rect 104690 73190 104810 73200
rect 104940 73190 105060 73200
rect 105190 73190 105310 73200
rect 105440 73190 105560 73200
rect 105690 73190 105810 73200
rect 105940 73190 106060 73200
rect 106190 73190 106310 73200
rect 106440 73190 106560 73200
rect 106690 73190 106810 73200
rect 106940 73190 107060 73200
rect 107190 73190 107310 73200
rect 107440 73190 107560 73200
rect 107690 73190 107810 73200
rect 107940 73190 108060 73200
rect 108190 73190 108310 73200
rect 108440 73190 108560 73200
rect 108690 73190 108810 73200
rect 108940 73190 109060 73200
rect 109190 73190 109310 73200
rect 109440 73190 109560 73200
rect 109690 73190 109810 73200
rect 109940 73190 110060 73200
rect 110190 73190 110310 73200
rect 110440 73190 110560 73200
rect 110690 73190 110810 73200
rect 110940 73190 111060 73200
rect 111190 73190 111310 73200
rect 111440 73190 111560 73200
rect 111690 73190 111810 73200
rect 111940 73190 112060 73200
rect 112190 73190 112310 73200
rect 112440 73190 112560 73200
rect 112690 73190 112810 73200
rect 112940 73190 113060 73200
rect 113190 73190 113310 73200
rect 113440 73190 113560 73200
rect 113690 73190 113810 73200
rect 113940 73190 114060 73200
rect 114190 73190 114310 73200
rect 114440 73190 114560 73200
rect 114690 73190 114810 73200
rect 114940 73190 115060 73200
rect 115190 73190 115310 73200
rect 115440 73190 115560 73200
rect 115690 73190 115810 73200
rect 115940 73190 116000 73200
rect 89000 73060 89050 73190
rect 89200 73060 89300 73190
rect 89450 73060 89550 73190
rect 89700 73060 89800 73190
rect 89950 73060 90050 73190
rect 90200 73060 90300 73190
rect 90450 73060 90550 73190
rect 90700 73060 90800 73190
rect 90950 73060 91050 73190
rect 91200 73060 91300 73190
rect 91450 73060 91550 73190
rect 91700 73060 91800 73190
rect 91950 73060 92050 73190
rect 92200 73060 92300 73190
rect 92450 73060 92550 73190
rect 92700 73060 92800 73190
rect 92950 73060 93050 73190
rect 93200 73060 93300 73190
rect 93450 73060 93550 73190
rect 93700 73060 93800 73190
rect 93950 73060 94050 73190
rect 94200 73060 94300 73190
rect 94450 73060 94550 73190
rect 94700 73060 94800 73190
rect 94950 73060 95050 73190
rect 95200 73060 95300 73190
rect 95450 73060 95550 73190
rect 95700 73060 95800 73190
rect 95950 73060 96050 73190
rect 96200 73060 96300 73190
rect 96450 73060 96550 73190
rect 96700 73060 96800 73190
rect 96950 73060 97050 73190
rect 97200 73060 97300 73190
rect 97450 73060 97550 73190
rect 97700 73060 97800 73190
rect 97950 73060 98050 73190
rect 98200 73060 98300 73190
rect 98450 73060 98550 73190
rect 98700 73060 98800 73190
rect 98950 73060 99050 73190
rect 99200 73060 99300 73190
rect 99450 73060 99550 73190
rect 99700 73060 99800 73190
rect 99950 73060 100050 73190
rect 100200 73060 100300 73190
rect 100450 73060 100550 73190
rect 100700 73060 100800 73190
rect 100950 73060 101050 73190
rect 101200 73060 101300 73190
rect 101450 73060 101550 73190
rect 101700 73060 101800 73190
rect 101950 73060 102050 73190
rect 102200 73060 102300 73190
rect 102450 73060 102550 73190
rect 102700 73060 102800 73190
rect 102950 73060 103050 73190
rect 103200 73060 103300 73190
rect 103450 73060 103550 73190
rect 103700 73060 103800 73190
rect 103950 73060 104050 73190
rect 104200 73060 104300 73190
rect 104450 73060 104550 73190
rect 104700 73060 104800 73190
rect 104950 73060 105050 73190
rect 105200 73060 105300 73190
rect 105450 73060 105550 73190
rect 105700 73060 105800 73190
rect 105950 73060 106050 73190
rect 106200 73060 106300 73190
rect 106450 73060 106550 73190
rect 106700 73060 106800 73190
rect 106950 73060 107050 73190
rect 107200 73060 107300 73190
rect 107450 73060 107550 73190
rect 107700 73060 107800 73190
rect 107950 73060 108050 73190
rect 108200 73060 108300 73190
rect 108450 73060 108550 73190
rect 108700 73060 108800 73190
rect 108950 73060 109050 73190
rect 109200 73060 109300 73190
rect 109450 73060 109550 73190
rect 109700 73060 109800 73190
rect 109950 73060 110050 73190
rect 110200 73060 110300 73190
rect 110450 73060 110550 73190
rect 110700 73060 110800 73190
rect 110950 73060 111050 73190
rect 111200 73060 111300 73190
rect 111450 73060 111550 73190
rect 111700 73060 111800 73190
rect 111950 73060 112050 73190
rect 112200 73060 112300 73190
rect 112450 73060 112550 73190
rect 112700 73060 112800 73190
rect 112950 73060 113050 73190
rect 113200 73060 113300 73190
rect 113450 73060 113550 73190
rect 113700 73060 113800 73190
rect 113950 73060 114050 73190
rect 114200 73060 114300 73190
rect 114450 73060 114550 73190
rect 114700 73060 114800 73190
rect 114950 73060 115050 73190
rect 115200 73060 115300 73190
rect 115450 73060 115550 73190
rect 115700 73060 115800 73190
rect 115950 73060 116000 73190
rect 89000 73050 89060 73060
rect 89190 73050 89310 73060
rect 89440 73050 89560 73060
rect 89690 73050 89810 73060
rect 89940 73050 90060 73060
rect 90190 73050 90310 73060
rect 90440 73050 90560 73060
rect 90690 73050 90810 73060
rect 90940 73050 91060 73060
rect 91190 73050 91310 73060
rect 91440 73050 91560 73060
rect 91690 73050 91810 73060
rect 91940 73050 92060 73060
rect 92190 73050 92310 73060
rect 92440 73050 92560 73060
rect 92690 73050 92810 73060
rect 92940 73050 93060 73060
rect 93190 73050 93310 73060
rect 93440 73050 93560 73060
rect 93690 73050 93810 73060
rect 93940 73050 94060 73060
rect 94190 73050 94310 73060
rect 94440 73050 94560 73060
rect 94690 73050 94810 73060
rect 94940 73050 95060 73060
rect 95190 73050 95310 73060
rect 95440 73050 95560 73060
rect 95690 73050 95810 73060
rect 95940 73050 96060 73060
rect 96190 73050 96310 73060
rect 96440 73050 96560 73060
rect 96690 73050 96810 73060
rect 96940 73050 97060 73060
rect 97190 73050 97310 73060
rect 97440 73050 97560 73060
rect 97690 73050 97810 73060
rect 97940 73050 98060 73060
rect 98190 73050 98310 73060
rect 98440 73050 98560 73060
rect 98690 73050 98810 73060
rect 98940 73050 99060 73060
rect 99190 73050 99310 73060
rect 99440 73050 99560 73060
rect 99690 73050 99810 73060
rect 99940 73050 100060 73060
rect 100190 73050 100310 73060
rect 100440 73050 100560 73060
rect 100690 73050 100810 73060
rect 100940 73050 101060 73060
rect 101190 73050 101310 73060
rect 101440 73050 101560 73060
rect 101690 73050 101810 73060
rect 101940 73050 102060 73060
rect 102190 73050 102310 73060
rect 102440 73050 102560 73060
rect 102690 73050 102810 73060
rect 102940 73050 103060 73060
rect 103190 73050 103310 73060
rect 103440 73050 103560 73060
rect 103690 73050 103810 73060
rect 103940 73050 104060 73060
rect 104190 73050 104310 73060
rect 104440 73050 104560 73060
rect 104690 73050 104810 73060
rect 104940 73050 105060 73060
rect 105190 73050 105310 73060
rect 105440 73050 105560 73060
rect 105690 73050 105810 73060
rect 105940 73050 106060 73060
rect 106190 73050 106310 73060
rect 106440 73050 106560 73060
rect 106690 73050 106810 73060
rect 106940 73050 107060 73060
rect 107190 73050 107310 73060
rect 107440 73050 107560 73060
rect 107690 73050 107810 73060
rect 107940 73050 108060 73060
rect 108190 73050 108310 73060
rect 108440 73050 108560 73060
rect 108690 73050 108810 73060
rect 108940 73050 109060 73060
rect 109190 73050 109310 73060
rect 109440 73050 109560 73060
rect 109690 73050 109810 73060
rect 109940 73050 110060 73060
rect 110190 73050 110310 73060
rect 110440 73050 110560 73060
rect 110690 73050 110810 73060
rect 110940 73050 111060 73060
rect 111190 73050 111310 73060
rect 111440 73050 111560 73060
rect 111690 73050 111810 73060
rect 111940 73050 112060 73060
rect 112190 73050 112310 73060
rect 112440 73050 112560 73060
rect 112690 73050 112810 73060
rect 112940 73050 113060 73060
rect 113190 73050 113310 73060
rect 113440 73050 113560 73060
rect 113690 73050 113810 73060
rect 113940 73050 114060 73060
rect 114190 73050 114310 73060
rect 114440 73050 114560 73060
rect 114690 73050 114810 73060
rect 114940 73050 115060 73060
rect 115190 73050 115310 73060
rect 115440 73050 115560 73060
rect 115690 73050 115810 73060
rect 115940 73050 116000 73060
rect 89000 72950 116000 73050
rect 89000 72940 89060 72950
rect 89190 72940 89310 72950
rect 89440 72940 89560 72950
rect 89690 72940 89810 72950
rect 89940 72940 90060 72950
rect 90190 72940 90310 72950
rect 90440 72940 90560 72950
rect 90690 72940 90810 72950
rect 90940 72940 91060 72950
rect 91190 72940 91310 72950
rect 91440 72940 91560 72950
rect 91690 72940 91810 72950
rect 91940 72940 92060 72950
rect 92190 72940 92310 72950
rect 92440 72940 92560 72950
rect 92690 72940 92810 72950
rect 92940 72940 93060 72950
rect 93190 72940 93310 72950
rect 93440 72940 93560 72950
rect 93690 72940 93810 72950
rect 93940 72940 94060 72950
rect 94190 72940 94310 72950
rect 94440 72940 94560 72950
rect 94690 72940 94810 72950
rect 94940 72940 95060 72950
rect 95190 72940 95310 72950
rect 95440 72940 95560 72950
rect 95690 72940 95810 72950
rect 95940 72940 96060 72950
rect 96190 72940 96310 72950
rect 96440 72940 96560 72950
rect 96690 72940 96810 72950
rect 96940 72940 97060 72950
rect 97190 72940 97310 72950
rect 97440 72940 97560 72950
rect 97690 72940 97810 72950
rect 97940 72940 98060 72950
rect 98190 72940 98310 72950
rect 98440 72940 98560 72950
rect 98690 72940 98810 72950
rect 98940 72940 99060 72950
rect 99190 72940 99310 72950
rect 99440 72940 99560 72950
rect 99690 72940 99810 72950
rect 99940 72940 100060 72950
rect 100190 72940 100310 72950
rect 100440 72940 100560 72950
rect 100690 72940 100810 72950
rect 100940 72940 101060 72950
rect 101190 72940 101310 72950
rect 101440 72940 101560 72950
rect 101690 72940 101810 72950
rect 101940 72940 102060 72950
rect 102190 72940 102310 72950
rect 102440 72940 102560 72950
rect 102690 72940 102810 72950
rect 102940 72940 103060 72950
rect 103190 72940 103310 72950
rect 103440 72940 103560 72950
rect 103690 72940 103810 72950
rect 103940 72940 104060 72950
rect 104190 72940 104310 72950
rect 104440 72940 104560 72950
rect 104690 72940 104810 72950
rect 104940 72940 105060 72950
rect 105190 72940 105310 72950
rect 105440 72940 105560 72950
rect 105690 72940 105810 72950
rect 105940 72940 106060 72950
rect 106190 72940 106310 72950
rect 106440 72940 106560 72950
rect 106690 72940 106810 72950
rect 106940 72940 107060 72950
rect 107190 72940 107310 72950
rect 107440 72940 107560 72950
rect 107690 72940 107810 72950
rect 107940 72940 108060 72950
rect 108190 72940 108310 72950
rect 108440 72940 108560 72950
rect 108690 72940 108810 72950
rect 108940 72940 109060 72950
rect 109190 72940 109310 72950
rect 109440 72940 109560 72950
rect 109690 72940 109810 72950
rect 109940 72940 110060 72950
rect 110190 72940 110310 72950
rect 110440 72940 110560 72950
rect 110690 72940 110810 72950
rect 110940 72940 111060 72950
rect 111190 72940 111310 72950
rect 111440 72940 111560 72950
rect 111690 72940 111810 72950
rect 111940 72940 112060 72950
rect 112190 72940 112310 72950
rect 112440 72940 112560 72950
rect 112690 72940 112810 72950
rect 112940 72940 113060 72950
rect 113190 72940 113310 72950
rect 113440 72940 113560 72950
rect 113690 72940 113810 72950
rect 113940 72940 114060 72950
rect 114190 72940 114310 72950
rect 114440 72940 114560 72950
rect 114690 72940 114810 72950
rect 114940 72940 115060 72950
rect 115190 72940 115310 72950
rect 115440 72940 115560 72950
rect 115690 72940 115810 72950
rect 115940 72940 116000 72950
rect 89000 72810 89050 72940
rect 89200 72810 89300 72940
rect 89450 72810 89550 72940
rect 89700 72810 89800 72940
rect 89950 72810 90050 72940
rect 90200 72810 90300 72940
rect 90450 72810 90550 72940
rect 90700 72810 90800 72940
rect 90950 72810 91050 72940
rect 91200 72810 91300 72940
rect 91450 72810 91550 72940
rect 91700 72810 91800 72940
rect 91950 72810 92050 72940
rect 92200 72810 92300 72940
rect 92450 72810 92550 72940
rect 92700 72810 92800 72940
rect 92950 72810 93050 72940
rect 93200 72810 93300 72940
rect 93450 72810 93550 72940
rect 93700 72810 93800 72940
rect 93950 72810 94050 72940
rect 94200 72810 94300 72940
rect 94450 72810 94550 72940
rect 94700 72810 94800 72940
rect 94950 72810 95050 72940
rect 95200 72810 95300 72940
rect 95450 72810 95550 72940
rect 95700 72810 95800 72940
rect 95950 72810 96050 72940
rect 96200 72810 96300 72940
rect 96450 72810 96550 72940
rect 96700 72810 96800 72940
rect 96950 72810 97050 72940
rect 97200 72810 97300 72940
rect 97450 72810 97550 72940
rect 97700 72810 97800 72940
rect 97950 72810 98050 72940
rect 98200 72810 98300 72940
rect 98450 72810 98550 72940
rect 98700 72810 98800 72940
rect 98950 72810 99050 72940
rect 99200 72810 99300 72940
rect 99450 72810 99550 72940
rect 99700 72810 99800 72940
rect 99950 72810 100050 72940
rect 100200 72810 100300 72940
rect 100450 72810 100550 72940
rect 100700 72810 100800 72940
rect 100950 72810 101050 72940
rect 101200 72810 101300 72940
rect 101450 72810 101550 72940
rect 101700 72810 101800 72940
rect 101950 72810 102050 72940
rect 102200 72810 102300 72940
rect 102450 72810 102550 72940
rect 102700 72810 102800 72940
rect 102950 72810 103050 72940
rect 103200 72810 103300 72940
rect 103450 72810 103550 72940
rect 103700 72810 103800 72940
rect 103950 72810 104050 72940
rect 104200 72810 104300 72940
rect 104450 72810 104550 72940
rect 104700 72810 104800 72940
rect 104950 72810 105050 72940
rect 105200 72810 105300 72940
rect 105450 72810 105550 72940
rect 105700 72810 105800 72940
rect 105950 72810 106050 72940
rect 106200 72810 106300 72940
rect 106450 72810 106550 72940
rect 106700 72810 106800 72940
rect 106950 72810 107050 72940
rect 107200 72810 107300 72940
rect 107450 72810 107550 72940
rect 107700 72810 107800 72940
rect 107950 72810 108050 72940
rect 108200 72810 108300 72940
rect 108450 72810 108550 72940
rect 108700 72810 108800 72940
rect 108950 72810 109050 72940
rect 109200 72810 109300 72940
rect 109450 72810 109550 72940
rect 109700 72810 109800 72940
rect 109950 72810 110050 72940
rect 110200 72810 110300 72940
rect 110450 72810 110550 72940
rect 110700 72810 110800 72940
rect 110950 72810 111050 72940
rect 111200 72810 111300 72940
rect 111450 72810 111550 72940
rect 111700 72810 111800 72940
rect 111950 72810 112050 72940
rect 112200 72810 112300 72940
rect 112450 72810 112550 72940
rect 112700 72810 112800 72940
rect 112950 72810 113050 72940
rect 113200 72810 113300 72940
rect 113450 72810 113550 72940
rect 113700 72810 113800 72940
rect 113950 72810 114050 72940
rect 114200 72810 114300 72940
rect 114450 72810 114550 72940
rect 114700 72810 114800 72940
rect 114950 72810 115050 72940
rect 115200 72810 115300 72940
rect 115450 72810 115550 72940
rect 115700 72810 115800 72940
rect 115950 72810 116000 72940
rect 89000 72800 89060 72810
rect 89190 72800 89310 72810
rect 89440 72800 89560 72810
rect 89690 72800 89810 72810
rect 89940 72800 90060 72810
rect 90190 72800 90310 72810
rect 90440 72800 90560 72810
rect 90690 72800 90810 72810
rect 90940 72800 91060 72810
rect 91190 72800 91310 72810
rect 91440 72800 91560 72810
rect 91690 72800 91810 72810
rect 91940 72800 92060 72810
rect 92190 72800 92310 72810
rect 92440 72800 92560 72810
rect 92690 72800 92810 72810
rect 92940 72800 93060 72810
rect 93190 72800 93310 72810
rect 93440 72800 93560 72810
rect 93690 72800 93810 72810
rect 93940 72800 94060 72810
rect 94190 72800 94310 72810
rect 94440 72800 94560 72810
rect 94690 72800 94810 72810
rect 94940 72800 95060 72810
rect 95190 72800 95310 72810
rect 95440 72800 95560 72810
rect 95690 72800 95810 72810
rect 95940 72800 96060 72810
rect 96190 72800 96310 72810
rect 96440 72800 96560 72810
rect 96690 72800 96810 72810
rect 96940 72800 97060 72810
rect 97190 72800 97310 72810
rect 97440 72800 97560 72810
rect 97690 72800 97810 72810
rect 97940 72800 98060 72810
rect 98190 72800 98310 72810
rect 98440 72800 98560 72810
rect 98690 72800 98810 72810
rect 98940 72800 99060 72810
rect 99190 72800 99310 72810
rect 99440 72800 99560 72810
rect 99690 72800 99810 72810
rect 99940 72800 100060 72810
rect 100190 72800 100310 72810
rect 100440 72800 100560 72810
rect 100690 72800 100810 72810
rect 100940 72800 101060 72810
rect 101190 72800 101310 72810
rect 101440 72800 101560 72810
rect 101690 72800 101810 72810
rect 101940 72800 102060 72810
rect 102190 72800 102310 72810
rect 102440 72800 102560 72810
rect 102690 72800 102810 72810
rect 102940 72800 103060 72810
rect 103190 72800 103310 72810
rect 103440 72800 103560 72810
rect 103690 72800 103810 72810
rect 103940 72800 104060 72810
rect 104190 72800 104310 72810
rect 104440 72800 104560 72810
rect 104690 72800 104810 72810
rect 104940 72800 105060 72810
rect 105190 72800 105310 72810
rect 105440 72800 105560 72810
rect 105690 72800 105810 72810
rect 105940 72800 106060 72810
rect 106190 72800 106310 72810
rect 106440 72800 106560 72810
rect 106690 72800 106810 72810
rect 106940 72800 107060 72810
rect 107190 72800 107310 72810
rect 107440 72800 107560 72810
rect 107690 72800 107810 72810
rect 107940 72800 108060 72810
rect 108190 72800 108310 72810
rect 108440 72800 108560 72810
rect 108690 72800 108810 72810
rect 108940 72800 109060 72810
rect 109190 72800 109310 72810
rect 109440 72800 109560 72810
rect 109690 72800 109810 72810
rect 109940 72800 110060 72810
rect 110190 72800 110310 72810
rect 110440 72800 110560 72810
rect 110690 72800 110810 72810
rect 110940 72800 111060 72810
rect 111190 72800 111310 72810
rect 111440 72800 111560 72810
rect 111690 72800 111810 72810
rect 111940 72800 112060 72810
rect 112190 72800 112310 72810
rect 112440 72800 112560 72810
rect 112690 72800 112810 72810
rect 112940 72800 113060 72810
rect 113190 72800 113310 72810
rect 113440 72800 113560 72810
rect 113690 72800 113810 72810
rect 113940 72800 114060 72810
rect 114190 72800 114310 72810
rect 114440 72800 114560 72810
rect 114690 72800 114810 72810
rect 114940 72800 115060 72810
rect 115190 72800 115310 72810
rect 115440 72800 115560 72810
rect 115690 72800 115810 72810
rect 115940 72800 116000 72810
rect 89000 72700 116000 72800
rect 89000 72690 89060 72700
rect 89190 72690 89310 72700
rect 89440 72690 89560 72700
rect 89690 72690 89810 72700
rect 89940 72690 90060 72700
rect 90190 72690 90310 72700
rect 90440 72690 90560 72700
rect 90690 72690 90810 72700
rect 90940 72690 91060 72700
rect 91190 72690 91310 72700
rect 91440 72690 91560 72700
rect 91690 72690 91810 72700
rect 91940 72690 92060 72700
rect 92190 72690 92310 72700
rect 92440 72690 92560 72700
rect 92690 72690 92810 72700
rect 92940 72690 93060 72700
rect 93190 72690 93310 72700
rect 93440 72690 93560 72700
rect 93690 72690 93810 72700
rect 93940 72690 94060 72700
rect 94190 72690 94310 72700
rect 94440 72690 94560 72700
rect 94690 72690 94810 72700
rect 94940 72690 95060 72700
rect 95190 72690 95310 72700
rect 95440 72690 95560 72700
rect 95690 72690 95810 72700
rect 95940 72690 96060 72700
rect 96190 72690 96310 72700
rect 96440 72690 96560 72700
rect 96690 72690 96810 72700
rect 96940 72690 97060 72700
rect 97190 72690 97310 72700
rect 97440 72690 97560 72700
rect 97690 72690 97810 72700
rect 97940 72690 98060 72700
rect 98190 72690 98310 72700
rect 98440 72690 98560 72700
rect 98690 72690 98810 72700
rect 98940 72690 99060 72700
rect 99190 72690 99310 72700
rect 99440 72690 99560 72700
rect 99690 72690 99810 72700
rect 99940 72690 100060 72700
rect 100190 72690 100310 72700
rect 100440 72690 100560 72700
rect 100690 72690 100810 72700
rect 100940 72690 101060 72700
rect 101190 72690 101310 72700
rect 101440 72690 101560 72700
rect 101690 72690 101810 72700
rect 101940 72690 102060 72700
rect 102190 72690 102310 72700
rect 102440 72690 102560 72700
rect 102690 72690 102810 72700
rect 102940 72690 103060 72700
rect 103190 72690 103310 72700
rect 103440 72690 103560 72700
rect 103690 72690 103810 72700
rect 103940 72690 104060 72700
rect 104190 72690 104310 72700
rect 104440 72690 104560 72700
rect 104690 72690 104810 72700
rect 104940 72690 105060 72700
rect 105190 72690 105310 72700
rect 105440 72690 105560 72700
rect 105690 72690 105810 72700
rect 105940 72690 106060 72700
rect 106190 72690 106310 72700
rect 106440 72690 106560 72700
rect 106690 72690 106810 72700
rect 106940 72690 107060 72700
rect 107190 72690 107310 72700
rect 107440 72690 107560 72700
rect 107690 72690 107810 72700
rect 107940 72690 108060 72700
rect 108190 72690 108310 72700
rect 108440 72690 108560 72700
rect 108690 72690 108810 72700
rect 108940 72690 109060 72700
rect 109190 72690 109310 72700
rect 109440 72690 109560 72700
rect 109690 72690 109810 72700
rect 109940 72690 110060 72700
rect 110190 72690 110310 72700
rect 110440 72690 110560 72700
rect 110690 72690 110810 72700
rect 110940 72690 111060 72700
rect 111190 72690 111310 72700
rect 111440 72690 111560 72700
rect 111690 72690 111810 72700
rect 111940 72690 112060 72700
rect 112190 72690 112310 72700
rect 112440 72690 112560 72700
rect 112690 72690 112810 72700
rect 112940 72690 113060 72700
rect 113190 72690 113310 72700
rect 113440 72690 113560 72700
rect 113690 72690 113810 72700
rect 113940 72690 114060 72700
rect 114190 72690 114310 72700
rect 114440 72690 114560 72700
rect 114690 72690 114810 72700
rect 114940 72690 115060 72700
rect 115190 72690 115310 72700
rect 115440 72690 115560 72700
rect 115690 72690 115810 72700
rect 115940 72690 116000 72700
rect 89000 72560 89050 72690
rect 89200 72560 89300 72690
rect 89450 72560 89550 72690
rect 89700 72560 89800 72690
rect 89950 72560 90050 72690
rect 90200 72560 90300 72690
rect 90450 72560 90550 72690
rect 90700 72560 90800 72690
rect 90950 72560 91050 72690
rect 91200 72560 91300 72690
rect 91450 72560 91550 72690
rect 91700 72560 91800 72690
rect 91950 72560 92050 72690
rect 92200 72560 92300 72690
rect 92450 72560 92550 72690
rect 92700 72560 92800 72690
rect 92950 72560 93050 72690
rect 93200 72560 93300 72690
rect 93450 72560 93550 72690
rect 93700 72560 93800 72690
rect 93950 72560 94050 72690
rect 94200 72560 94300 72690
rect 94450 72560 94550 72690
rect 94700 72560 94800 72690
rect 94950 72560 95050 72690
rect 95200 72560 95300 72690
rect 95450 72560 95550 72690
rect 95700 72560 95800 72690
rect 95950 72560 96050 72690
rect 96200 72560 96300 72690
rect 96450 72560 96550 72690
rect 96700 72560 96800 72690
rect 96950 72560 97050 72690
rect 97200 72560 97300 72690
rect 97450 72560 97550 72690
rect 97700 72560 97800 72690
rect 97950 72560 98050 72690
rect 98200 72560 98300 72690
rect 98450 72560 98550 72690
rect 98700 72560 98800 72690
rect 98950 72560 99050 72690
rect 99200 72560 99300 72690
rect 99450 72560 99550 72690
rect 99700 72560 99800 72690
rect 99950 72560 100050 72690
rect 100200 72560 100300 72690
rect 100450 72560 100550 72690
rect 100700 72560 100800 72690
rect 100950 72560 101050 72690
rect 101200 72560 101300 72690
rect 101450 72560 101550 72690
rect 101700 72560 101800 72690
rect 101950 72560 102050 72690
rect 102200 72560 102300 72690
rect 102450 72560 102550 72690
rect 102700 72560 102800 72690
rect 102950 72560 103050 72690
rect 103200 72560 103300 72690
rect 103450 72560 103550 72690
rect 103700 72560 103800 72690
rect 103950 72560 104050 72690
rect 104200 72560 104300 72690
rect 104450 72560 104550 72690
rect 104700 72560 104800 72690
rect 104950 72560 105050 72690
rect 105200 72560 105300 72690
rect 105450 72560 105550 72690
rect 105700 72560 105800 72690
rect 105950 72560 106050 72690
rect 106200 72560 106300 72690
rect 106450 72560 106550 72690
rect 106700 72560 106800 72690
rect 106950 72560 107050 72690
rect 107200 72560 107300 72690
rect 107450 72560 107550 72690
rect 107700 72560 107800 72690
rect 107950 72560 108050 72690
rect 108200 72560 108300 72690
rect 108450 72560 108550 72690
rect 108700 72560 108800 72690
rect 108950 72560 109050 72690
rect 109200 72560 109300 72690
rect 109450 72560 109550 72690
rect 109700 72560 109800 72690
rect 109950 72560 110050 72690
rect 110200 72560 110300 72690
rect 110450 72560 110550 72690
rect 110700 72560 110800 72690
rect 110950 72560 111050 72690
rect 111200 72560 111300 72690
rect 111450 72560 111550 72690
rect 111700 72560 111800 72690
rect 111950 72560 112050 72690
rect 112200 72560 112300 72690
rect 112450 72560 112550 72690
rect 112700 72560 112800 72690
rect 112950 72560 113050 72690
rect 113200 72560 113300 72690
rect 113450 72560 113550 72690
rect 113700 72560 113800 72690
rect 113950 72560 114050 72690
rect 114200 72560 114300 72690
rect 114450 72560 114550 72690
rect 114700 72560 114800 72690
rect 114950 72560 115050 72690
rect 115200 72560 115300 72690
rect 115450 72560 115550 72690
rect 115700 72560 115800 72690
rect 115950 72560 116000 72690
rect 89000 72550 89060 72560
rect 89190 72550 89310 72560
rect 89440 72550 89560 72560
rect 89690 72550 89810 72560
rect 89940 72550 90060 72560
rect 90190 72550 90310 72560
rect 90440 72550 90560 72560
rect 90690 72550 90810 72560
rect 90940 72550 91060 72560
rect 91190 72550 91310 72560
rect 91440 72550 91560 72560
rect 91690 72550 91810 72560
rect 91940 72550 92060 72560
rect 92190 72550 92310 72560
rect 92440 72550 92560 72560
rect 92690 72550 92810 72560
rect 92940 72550 93060 72560
rect 93190 72550 93310 72560
rect 93440 72550 93560 72560
rect 93690 72550 93810 72560
rect 93940 72550 94060 72560
rect 94190 72550 94310 72560
rect 94440 72550 94560 72560
rect 94690 72550 94810 72560
rect 94940 72550 95060 72560
rect 95190 72550 95310 72560
rect 95440 72550 95560 72560
rect 95690 72550 95810 72560
rect 95940 72550 96060 72560
rect 96190 72550 96310 72560
rect 96440 72550 96560 72560
rect 96690 72550 96810 72560
rect 96940 72550 97060 72560
rect 97190 72550 97310 72560
rect 97440 72550 97560 72560
rect 97690 72550 97810 72560
rect 97940 72550 98060 72560
rect 98190 72550 98310 72560
rect 98440 72550 98560 72560
rect 98690 72550 98810 72560
rect 98940 72550 99060 72560
rect 99190 72550 99310 72560
rect 99440 72550 99560 72560
rect 99690 72550 99810 72560
rect 99940 72550 100060 72560
rect 100190 72550 100310 72560
rect 100440 72550 100560 72560
rect 100690 72550 100810 72560
rect 100940 72550 101060 72560
rect 101190 72550 101310 72560
rect 101440 72550 101560 72560
rect 101690 72550 101810 72560
rect 101940 72550 102060 72560
rect 102190 72550 102310 72560
rect 102440 72550 102560 72560
rect 102690 72550 102810 72560
rect 102940 72550 103060 72560
rect 103190 72550 103310 72560
rect 103440 72550 103560 72560
rect 103690 72550 103810 72560
rect 103940 72550 104060 72560
rect 104190 72550 104310 72560
rect 104440 72550 104560 72560
rect 104690 72550 104810 72560
rect 104940 72550 105060 72560
rect 105190 72550 105310 72560
rect 105440 72550 105560 72560
rect 105690 72550 105810 72560
rect 105940 72550 106060 72560
rect 106190 72550 106310 72560
rect 106440 72550 106560 72560
rect 106690 72550 106810 72560
rect 106940 72550 107060 72560
rect 107190 72550 107310 72560
rect 107440 72550 107560 72560
rect 107690 72550 107810 72560
rect 107940 72550 108060 72560
rect 108190 72550 108310 72560
rect 108440 72550 108560 72560
rect 108690 72550 108810 72560
rect 108940 72550 109060 72560
rect 109190 72550 109310 72560
rect 109440 72550 109560 72560
rect 109690 72550 109810 72560
rect 109940 72550 110060 72560
rect 110190 72550 110310 72560
rect 110440 72550 110560 72560
rect 110690 72550 110810 72560
rect 110940 72550 111060 72560
rect 111190 72550 111310 72560
rect 111440 72550 111560 72560
rect 111690 72550 111810 72560
rect 111940 72550 112060 72560
rect 112190 72550 112310 72560
rect 112440 72550 112560 72560
rect 112690 72550 112810 72560
rect 112940 72550 113060 72560
rect 113190 72550 113310 72560
rect 113440 72550 113560 72560
rect 113690 72550 113810 72560
rect 113940 72550 114060 72560
rect 114190 72550 114310 72560
rect 114440 72550 114560 72560
rect 114690 72550 114810 72560
rect 114940 72550 115060 72560
rect 115190 72550 115310 72560
rect 115440 72550 115560 72560
rect 115690 72550 115810 72560
rect 115940 72550 116000 72560
rect 89000 72450 116000 72550
rect 89000 72440 89060 72450
rect 89190 72440 89310 72450
rect 89440 72440 89560 72450
rect 89690 72440 89810 72450
rect 89940 72440 90060 72450
rect 90190 72440 90310 72450
rect 90440 72440 90560 72450
rect 90690 72440 90810 72450
rect 90940 72440 91060 72450
rect 91190 72440 91310 72450
rect 91440 72440 91560 72450
rect 91690 72440 91810 72450
rect 91940 72440 92060 72450
rect 92190 72440 92310 72450
rect 92440 72440 92560 72450
rect 92690 72440 92810 72450
rect 92940 72440 93060 72450
rect 93190 72440 93310 72450
rect 93440 72440 93560 72450
rect 93690 72440 93810 72450
rect 93940 72440 94060 72450
rect 94190 72440 94310 72450
rect 94440 72440 94560 72450
rect 94690 72440 94810 72450
rect 94940 72440 95060 72450
rect 95190 72440 95310 72450
rect 95440 72440 95560 72450
rect 95690 72440 95810 72450
rect 95940 72440 96060 72450
rect 96190 72440 96310 72450
rect 96440 72440 96560 72450
rect 96690 72440 96810 72450
rect 96940 72440 97060 72450
rect 97190 72440 97310 72450
rect 97440 72440 97560 72450
rect 97690 72440 97810 72450
rect 97940 72440 98060 72450
rect 98190 72440 98310 72450
rect 98440 72440 98560 72450
rect 98690 72440 98810 72450
rect 98940 72440 99060 72450
rect 99190 72440 99310 72450
rect 99440 72440 99560 72450
rect 99690 72440 99810 72450
rect 99940 72440 100060 72450
rect 100190 72440 100310 72450
rect 100440 72440 100560 72450
rect 100690 72440 100810 72450
rect 100940 72440 101060 72450
rect 101190 72440 101310 72450
rect 101440 72440 101560 72450
rect 101690 72440 101810 72450
rect 101940 72440 102060 72450
rect 102190 72440 102310 72450
rect 102440 72440 102560 72450
rect 102690 72440 102810 72450
rect 102940 72440 103060 72450
rect 103190 72440 103310 72450
rect 103440 72440 103560 72450
rect 103690 72440 103810 72450
rect 103940 72440 104060 72450
rect 104190 72440 104310 72450
rect 104440 72440 104560 72450
rect 104690 72440 104810 72450
rect 104940 72440 105060 72450
rect 105190 72440 105310 72450
rect 105440 72440 105560 72450
rect 105690 72440 105810 72450
rect 105940 72440 106060 72450
rect 106190 72440 106310 72450
rect 106440 72440 106560 72450
rect 106690 72440 106810 72450
rect 106940 72440 107060 72450
rect 107190 72440 107310 72450
rect 107440 72440 107560 72450
rect 107690 72440 107810 72450
rect 107940 72440 108060 72450
rect 108190 72440 108310 72450
rect 108440 72440 108560 72450
rect 108690 72440 108810 72450
rect 108940 72440 109060 72450
rect 109190 72440 109310 72450
rect 109440 72440 109560 72450
rect 109690 72440 109810 72450
rect 109940 72440 110060 72450
rect 110190 72440 110310 72450
rect 110440 72440 110560 72450
rect 110690 72440 110810 72450
rect 110940 72440 111060 72450
rect 111190 72440 111310 72450
rect 111440 72440 111560 72450
rect 111690 72440 111810 72450
rect 111940 72440 112060 72450
rect 112190 72440 112310 72450
rect 112440 72440 112560 72450
rect 112690 72440 112810 72450
rect 112940 72440 113060 72450
rect 113190 72440 113310 72450
rect 113440 72440 113560 72450
rect 113690 72440 113810 72450
rect 113940 72440 114060 72450
rect 114190 72440 114310 72450
rect 114440 72440 114560 72450
rect 114690 72440 114810 72450
rect 114940 72440 115060 72450
rect 115190 72440 115310 72450
rect 115440 72440 115560 72450
rect 115690 72440 115810 72450
rect 115940 72440 116000 72450
rect 89000 72310 89050 72440
rect 89200 72310 89300 72440
rect 89450 72310 89550 72440
rect 89700 72310 89800 72440
rect 89950 72310 90050 72440
rect 90200 72310 90300 72440
rect 90450 72310 90550 72440
rect 90700 72310 90800 72440
rect 90950 72310 91050 72440
rect 91200 72310 91300 72440
rect 91450 72310 91550 72440
rect 91700 72310 91800 72440
rect 91950 72310 92050 72440
rect 92200 72310 92300 72440
rect 92450 72310 92550 72440
rect 92700 72310 92800 72440
rect 92950 72310 93050 72440
rect 93200 72310 93300 72440
rect 93450 72310 93550 72440
rect 93700 72310 93800 72440
rect 93950 72310 94050 72440
rect 94200 72310 94300 72440
rect 94450 72310 94550 72440
rect 94700 72310 94800 72440
rect 94950 72310 95050 72440
rect 95200 72310 95300 72440
rect 95450 72310 95550 72440
rect 95700 72310 95800 72440
rect 95950 72310 96050 72440
rect 96200 72310 96300 72440
rect 96450 72310 96550 72440
rect 96700 72310 96800 72440
rect 96950 72310 97050 72440
rect 97200 72310 97300 72440
rect 97450 72310 97550 72440
rect 97700 72310 97800 72440
rect 97950 72310 98050 72440
rect 98200 72310 98300 72440
rect 98450 72310 98550 72440
rect 98700 72310 98800 72440
rect 98950 72310 99050 72440
rect 99200 72310 99300 72440
rect 99450 72310 99550 72440
rect 99700 72310 99800 72440
rect 99950 72310 100050 72440
rect 100200 72310 100300 72440
rect 100450 72310 100550 72440
rect 100700 72310 100800 72440
rect 100950 72310 101050 72440
rect 101200 72310 101300 72440
rect 101450 72310 101550 72440
rect 101700 72310 101800 72440
rect 101950 72310 102050 72440
rect 102200 72310 102300 72440
rect 102450 72310 102550 72440
rect 102700 72310 102800 72440
rect 102950 72310 103050 72440
rect 103200 72310 103300 72440
rect 103450 72310 103550 72440
rect 103700 72310 103800 72440
rect 103950 72310 104050 72440
rect 104200 72310 104300 72440
rect 104450 72310 104550 72440
rect 104700 72310 104800 72440
rect 104950 72310 105050 72440
rect 105200 72310 105300 72440
rect 105450 72310 105550 72440
rect 105700 72310 105800 72440
rect 105950 72310 106050 72440
rect 106200 72310 106300 72440
rect 106450 72310 106550 72440
rect 106700 72310 106800 72440
rect 106950 72310 107050 72440
rect 107200 72310 107300 72440
rect 107450 72310 107550 72440
rect 107700 72310 107800 72440
rect 107950 72310 108050 72440
rect 108200 72310 108300 72440
rect 108450 72310 108550 72440
rect 108700 72310 108800 72440
rect 108950 72310 109050 72440
rect 109200 72310 109300 72440
rect 109450 72310 109550 72440
rect 109700 72310 109800 72440
rect 109950 72310 110050 72440
rect 110200 72310 110300 72440
rect 110450 72310 110550 72440
rect 110700 72310 110800 72440
rect 110950 72310 111050 72440
rect 111200 72310 111300 72440
rect 111450 72310 111550 72440
rect 111700 72310 111800 72440
rect 111950 72310 112050 72440
rect 112200 72310 112300 72440
rect 112450 72310 112550 72440
rect 112700 72310 112800 72440
rect 112950 72310 113050 72440
rect 113200 72310 113300 72440
rect 113450 72310 113550 72440
rect 113700 72310 113800 72440
rect 113950 72310 114050 72440
rect 114200 72310 114300 72440
rect 114450 72310 114550 72440
rect 114700 72310 114800 72440
rect 114950 72310 115050 72440
rect 115200 72310 115300 72440
rect 115450 72310 115550 72440
rect 115700 72310 115800 72440
rect 115950 72310 116000 72440
rect 89000 72300 89060 72310
rect 89190 72300 89310 72310
rect 89440 72300 89560 72310
rect 89690 72300 89810 72310
rect 89940 72300 90060 72310
rect 90190 72300 90310 72310
rect 90440 72300 90560 72310
rect 90690 72300 90810 72310
rect 90940 72300 91060 72310
rect 91190 72300 91310 72310
rect 91440 72300 91560 72310
rect 91690 72300 91810 72310
rect 91940 72300 92060 72310
rect 92190 72300 92310 72310
rect 92440 72300 92560 72310
rect 92690 72300 92810 72310
rect 92940 72300 93060 72310
rect 93190 72300 93310 72310
rect 93440 72300 93560 72310
rect 93690 72300 93810 72310
rect 93940 72300 94060 72310
rect 94190 72300 94310 72310
rect 94440 72300 94560 72310
rect 94690 72300 94810 72310
rect 94940 72300 95060 72310
rect 95190 72300 95310 72310
rect 95440 72300 95560 72310
rect 95690 72300 95810 72310
rect 95940 72300 96060 72310
rect 96190 72300 96310 72310
rect 96440 72300 96560 72310
rect 96690 72300 96810 72310
rect 96940 72300 97060 72310
rect 97190 72300 97310 72310
rect 97440 72300 97560 72310
rect 97690 72300 97810 72310
rect 97940 72300 98060 72310
rect 98190 72300 98310 72310
rect 98440 72300 98560 72310
rect 98690 72300 98810 72310
rect 98940 72300 99060 72310
rect 99190 72300 99310 72310
rect 99440 72300 99560 72310
rect 99690 72300 99810 72310
rect 99940 72300 100060 72310
rect 100190 72300 100310 72310
rect 100440 72300 100560 72310
rect 100690 72300 100810 72310
rect 100940 72300 101060 72310
rect 101190 72300 101310 72310
rect 101440 72300 101560 72310
rect 101690 72300 101810 72310
rect 101940 72300 102060 72310
rect 102190 72300 102310 72310
rect 102440 72300 102560 72310
rect 102690 72300 102810 72310
rect 102940 72300 103060 72310
rect 103190 72300 103310 72310
rect 103440 72300 103560 72310
rect 103690 72300 103810 72310
rect 103940 72300 104060 72310
rect 104190 72300 104310 72310
rect 104440 72300 104560 72310
rect 104690 72300 104810 72310
rect 104940 72300 105060 72310
rect 105190 72300 105310 72310
rect 105440 72300 105560 72310
rect 105690 72300 105810 72310
rect 105940 72300 106060 72310
rect 106190 72300 106310 72310
rect 106440 72300 106560 72310
rect 106690 72300 106810 72310
rect 106940 72300 107060 72310
rect 107190 72300 107310 72310
rect 107440 72300 107560 72310
rect 107690 72300 107810 72310
rect 107940 72300 108060 72310
rect 108190 72300 108310 72310
rect 108440 72300 108560 72310
rect 108690 72300 108810 72310
rect 108940 72300 109060 72310
rect 109190 72300 109310 72310
rect 109440 72300 109560 72310
rect 109690 72300 109810 72310
rect 109940 72300 110060 72310
rect 110190 72300 110310 72310
rect 110440 72300 110560 72310
rect 110690 72300 110810 72310
rect 110940 72300 111060 72310
rect 111190 72300 111310 72310
rect 111440 72300 111560 72310
rect 111690 72300 111810 72310
rect 111940 72300 112060 72310
rect 112190 72300 112310 72310
rect 112440 72300 112560 72310
rect 112690 72300 112810 72310
rect 112940 72300 113060 72310
rect 113190 72300 113310 72310
rect 113440 72300 113560 72310
rect 113690 72300 113810 72310
rect 113940 72300 114060 72310
rect 114190 72300 114310 72310
rect 114440 72300 114560 72310
rect 114690 72300 114810 72310
rect 114940 72300 115060 72310
rect 115190 72300 115310 72310
rect 115440 72300 115560 72310
rect 115690 72300 115810 72310
rect 115940 72300 116000 72310
rect 89000 72200 116000 72300
rect 89000 72190 89060 72200
rect 89190 72190 89310 72200
rect 89440 72190 89560 72200
rect 89690 72190 89810 72200
rect 89940 72190 90060 72200
rect 90190 72190 90310 72200
rect 90440 72190 90560 72200
rect 90690 72190 90810 72200
rect 90940 72190 91060 72200
rect 91190 72190 91310 72200
rect 91440 72190 91560 72200
rect 91690 72190 91810 72200
rect 91940 72190 92060 72200
rect 92190 72190 92310 72200
rect 92440 72190 92560 72200
rect 92690 72190 92810 72200
rect 92940 72190 93060 72200
rect 93190 72190 93310 72200
rect 93440 72190 93560 72200
rect 93690 72190 93810 72200
rect 93940 72190 94060 72200
rect 94190 72190 94310 72200
rect 94440 72190 94560 72200
rect 94690 72190 94810 72200
rect 94940 72190 95060 72200
rect 95190 72190 95310 72200
rect 95440 72190 95560 72200
rect 95690 72190 95810 72200
rect 95940 72190 96060 72200
rect 96190 72190 96310 72200
rect 96440 72190 96560 72200
rect 96690 72190 96810 72200
rect 96940 72190 97060 72200
rect 97190 72190 97310 72200
rect 97440 72190 97560 72200
rect 97690 72190 97810 72200
rect 97940 72190 98060 72200
rect 98190 72190 98310 72200
rect 98440 72190 98560 72200
rect 98690 72190 98810 72200
rect 98940 72190 99060 72200
rect 99190 72190 99310 72200
rect 99440 72190 99560 72200
rect 99690 72190 99810 72200
rect 99940 72190 100060 72200
rect 100190 72190 100310 72200
rect 100440 72190 100560 72200
rect 100690 72190 100810 72200
rect 100940 72190 101060 72200
rect 101190 72190 101310 72200
rect 101440 72190 101560 72200
rect 101690 72190 101810 72200
rect 101940 72190 102060 72200
rect 102190 72190 102310 72200
rect 102440 72190 102560 72200
rect 102690 72190 102810 72200
rect 102940 72190 103060 72200
rect 103190 72190 103310 72200
rect 103440 72190 103560 72200
rect 103690 72190 103810 72200
rect 103940 72190 104060 72200
rect 104190 72190 104310 72200
rect 104440 72190 104560 72200
rect 104690 72190 104810 72200
rect 104940 72190 105060 72200
rect 105190 72190 105310 72200
rect 105440 72190 105560 72200
rect 105690 72190 105810 72200
rect 105940 72190 106060 72200
rect 106190 72190 106310 72200
rect 106440 72190 106560 72200
rect 106690 72190 106810 72200
rect 106940 72190 107060 72200
rect 107190 72190 107310 72200
rect 107440 72190 107560 72200
rect 107690 72190 107810 72200
rect 107940 72190 108060 72200
rect 108190 72190 108310 72200
rect 108440 72190 108560 72200
rect 108690 72190 108810 72200
rect 108940 72190 109060 72200
rect 109190 72190 109310 72200
rect 109440 72190 109560 72200
rect 109690 72190 109810 72200
rect 109940 72190 110060 72200
rect 110190 72190 110310 72200
rect 110440 72190 110560 72200
rect 110690 72190 110810 72200
rect 110940 72190 111060 72200
rect 111190 72190 111310 72200
rect 111440 72190 111560 72200
rect 111690 72190 111810 72200
rect 111940 72190 112060 72200
rect 112190 72190 112310 72200
rect 112440 72190 112560 72200
rect 112690 72190 112810 72200
rect 112940 72190 113060 72200
rect 113190 72190 113310 72200
rect 113440 72190 113560 72200
rect 113690 72190 113810 72200
rect 113940 72190 114060 72200
rect 114190 72190 114310 72200
rect 114440 72190 114560 72200
rect 114690 72190 114810 72200
rect 114940 72190 115060 72200
rect 115190 72190 115310 72200
rect 115440 72190 115560 72200
rect 115690 72190 115810 72200
rect 115940 72190 116000 72200
rect 89000 72060 89050 72190
rect 89200 72060 89300 72190
rect 89450 72060 89550 72190
rect 89700 72060 89800 72190
rect 89950 72060 90050 72190
rect 90200 72060 90300 72190
rect 90450 72060 90550 72190
rect 90700 72060 90800 72190
rect 90950 72060 91050 72190
rect 91200 72060 91300 72190
rect 91450 72060 91550 72190
rect 91700 72060 91800 72190
rect 91950 72060 92050 72190
rect 92200 72060 92300 72190
rect 92450 72060 92550 72190
rect 92700 72060 92800 72190
rect 92950 72060 93050 72190
rect 93200 72060 93300 72190
rect 93450 72060 93550 72190
rect 93700 72060 93800 72190
rect 93950 72060 94050 72190
rect 94200 72060 94300 72190
rect 94450 72060 94550 72190
rect 94700 72060 94800 72190
rect 94950 72060 95050 72190
rect 95200 72060 95300 72190
rect 95450 72060 95550 72190
rect 95700 72060 95800 72190
rect 95950 72060 96050 72190
rect 96200 72060 96300 72190
rect 96450 72060 96550 72190
rect 96700 72060 96800 72190
rect 96950 72060 97050 72190
rect 97200 72060 97300 72190
rect 97450 72060 97550 72190
rect 97700 72060 97800 72190
rect 97950 72060 98050 72190
rect 98200 72060 98300 72190
rect 98450 72060 98550 72190
rect 98700 72060 98800 72190
rect 98950 72060 99050 72190
rect 99200 72060 99300 72190
rect 99450 72060 99550 72190
rect 99700 72060 99800 72190
rect 99950 72060 100050 72190
rect 100200 72060 100300 72190
rect 100450 72060 100550 72190
rect 100700 72060 100800 72190
rect 100950 72060 101050 72190
rect 101200 72060 101300 72190
rect 101450 72060 101550 72190
rect 101700 72060 101800 72190
rect 101950 72060 102050 72190
rect 102200 72060 102300 72190
rect 102450 72060 102550 72190
rect 102700 72060 102800 72190
rect 102950 72060 103050 72190
rect 103200 72060 103300 72190
rect 103450 72060 103550 72190
rect 103700 72060 103800 72190
rect 103950 72060 104050 72190
rect 104200 72060 104300 72190
rect 104450 72060 104550 72190
rect 104700 72060 104800 72190
rect 104950 72060 105050 72190
rect 105200 72060 105300 72190
rect 105450 72060 105550 72190
rect 105700 72060 105800 72190
rect 105950 72060 106050 72190
rect 106200 72060 106300 72190
rect 106450 72060 106550 72190
rect 106700 72060 106800 72190
rect 106950 72060 107050 72190
rect 107200 72060 107300 72190
rect 107450 72060 107550 72190
rect 107700 72060 107800 72190
rect 107950 72060 108050 72190
rect 108200 72060 108300 72190
rect 108450 72060 108550 72190
rect 108700 72060 108800 72190
rect 108950 72060 109050 72190
rect 109200 72060 109300 72190
rect 109450 72060 109550 72190
rect 109700 72060 109800 72190
rect 109950 72060 110050 72190
rect 110200 72060 110300 72190
rect 110450 72060 110550 72190
rect 110700 72060 110800 72190
rect 110950 72060 111050 72190
rect 111200 72060 111300 72190
rect 111450 72060 111550 72190
rect 111700 72060 111800 72190
rect 111950 72060 112050 72190
rect 112200 72060 112300 72190
rect 112450 72060 112550 72190
rect 112700 72060 112800 72190
rect 112950 72060 113050 72190
rect 113200 72060 113300 72190
rect 113450 72060 113550 72190
rect 113700 72060 113800 72190
rect 113950 72060 114050 72190
rect 114200 72060 114300 72190
rect 114450 72060 114550 72190
rect 114700 72060 114800 72190
rect 114950 72060 115050 72190
rect 115200 72060 115300 72190
rect 115450 72060 115550 72190
rect 115700 72060 115800 72190
rect 115950 72060 116000 72190
rect 89000 72050 89060 72060
rect 89190 72050 89310 72060
rect 89440 72050 89560 72060
rect 89690 72050 89810 72060
rect 89940 72050 90060 72060
rect 90190 72050 90310 72060
rect 90440 72050 90560 72060
rect 90690 72050 90810 72060
rect 90940 72050 91060 72060
rect 91190 72050 91310 72060
rect 91440 72050 91560 72060
rect 91690 72050 91810 72060
rect 91940 72050 92060 72060
rect 92190 72050 92310 72060
rect 92440 72050 92560 72060
rect 92690 72050 92810 72060
rect 92940 72050 93060 72060
rect 93190 72050 93310 72060
rect 93440 72050 93560 72060
rect 93690 72050 93810 72060
rect 93940 72050 94060 72060
rect 94190 72050 94310 72060
rect 94440 72050 94560 72060
rect 94690 72050 94810 72060
rect 94940 72050 95060 72060
rect 95190 72050 95310 72060
rect 95440 72050 95560 72060
rect 95690 72050 95810 72060
rect 95940 72050 96060 72060
rect 96190 72050 96310 72060
rect 96440 72050 96560 72060
rect 96690 72050 96810 72060
rect 96940 72050 97060 72060
rect 97190 72050 97310 72060
rect 97440 72050 97560 72060
rect 97690 72050 97810 72060
rect 97940 72050 98060 72060
rect 98190 72050 98310 72060
rect 98440 72050 98560 72060
rect 98690 72050 98810 72060
rect 98940 72050 99060 72060
rect 99190 72050 99310 72060
rect 99440 72050 99560 72060
rect 99690 72050 99810 72060
rect 99940 72050 100060 72060
rect 100190 72050 100310 72060
rect 100440 72050 100560 72060
rect 100690 72050 100810 72060
rect 100940 72050 101060 72060
rect 101190 72050 101310 72060
rect 101440 72050 101560 72060
rect 101690 72050 101810 72060
rect 101940 72050 102060 72060
rect 102190 72050 102310 72060
rect 102440 72050 102560 72060
rect 102690 72050 102810 72060
rect 102940 72050 103060 72060
rect 103190 72050 103310 72060
rect 103440 72050 103560 72060
rect 103690 72050 103810 72060
rect 103940 72050 104060 72060
rect 104190 72050 104310 72060
rect 104440 72050 104560 72060
rect 104690 72050 104810 72060
rect 104940 72050 105060 72060
rect 105190 72050 105310 72060
rect 105440 72050 105560 72060
rect 105690 72050 105810 72060
rect 105940 72050 106060 72060
rect 106190 72050 106310 72060
rect 106440 72050 106560 72060
rect 106690 72050 106810 72060
rect 106940 72050 107060 72060
rect 107190 72050 107310 72060
rect 107440 72050 107560 72060
rect 107690 72050 107810 72060
rect 107940 72050 108060 72060
rect 108190 72050 108310 72060
rect 108440 72050 108560 72060
rect 108690 72050 108810 72060
rect 108940 72050 109060 72060
rect 109190 72050 109310 72060
rect 109440 72050 109560 72060
rect 109690 72050 109810 72060
rect 109940 72050 110060 72060
rect 110190 72050 110310 72060
rect 110440 72050 110560 72060
rect 110690 72050 110810 72060
rect 110940 72050 111060 72060
rect 111190 72050 111310 72060
rect 111440 72050 111560 72060
rect 111690 72050 111810 72060
rect 111940 72050 112060 72060
rect 112190 72050 112310 72060
rect 112440 72050 112560 72060
rect 112690 72050 112810 72060
rect 112940 72050 113060 72060
rect 113190 72050 113310 72060
rect 113440 72050 113560 72060
rect 113690 72050 113810 72060
rect 113940 72050 114060 72060
rect 114190 72050 114310 72060
rect 114440 72050 114560 72060
rect 114690 72050 114810 72060
rect 114940 72050 115060 72060
rect 115190 72050 115310 72060
rect 115440 72050 115560 72060
rect 115690 72050 115810 72060
rect 115940 72050 116000 72060
rect 89000 71950 116000 72050
rect 89000 71940 89060 71950
rect 89190 71940 89310 71950
rect 89440 71940 89560 71950
rect 89690 71940 89810 71950
rect 89940 71940 90060 71950
rect 90190 71940 90310 71950
rect 90440 71940 90560 71950
rect 90690 71940 90810 71950
rect 90940 71940 91060 71950
rect 91190 71940 91310 71950
rect 91440 71940 91560 71950
rect 91690 71940 91810 71950
rect 91940 71940 92060 71950
rect 92190 71940 92310 71950
rect 92440 71940 92560 71950
rect 92690 71940 92810 71950
rect 92940 71940 93060 71950
rect 93190 71940 93310 71950
rect 93440 71940 93560 71950
rect 93690 71940 93810 71950
rect 93940 71940 94060 71950
rect 94190 71940 94310 71950
rect 94440 71940 94560 71950
rect 94690 71940 94810 71950
rect 94940 71940 95060 71950
rect 95190 71940 95310 71950
rect 95440 71940 95560 71950
rect 95690 71940 95810 71950
rect 95940 71940 96060 71950
rect 96190 71940 96310 71950
rect 96440 71940 96560 71950
rect 96690 71940 96810 71950
rect 96940 71940 97060 71950
rect 97190 71940 97310 71950
rect 97440 71940 97560 71950
rect 97690 71940 97810 71950
rect 97940 71940 98060 71950
rect 98190 71940 98310 71950
rect 98440 71940 98560 71950
rect 98690 71940 98810 71950
rect 98940 71940 99060 71950
rect 99190 71940 99310 71950
rect 99440 71940 99560 71950
rect 99690 71940 99810 71950
rect 99940 71940 100060 71950
rect 100190 71940 100310 71950
rect 100440 71940 100560 71950
rect 100690 71940 100810 71950
rect 100940 71940 101060 71950
rect 101190 71940 101310 71950
rect 101440 71940 101560 71950
rect 101690 71940 101810 71950
rect 101940 71940 102060 71950
rect 102190 71940 102310 71950
rect 102440 71940 102560 71950
rect 102690 71940 102810 71950
rect 102940 71940 103060 71950
rect 103190 71940 103310 71950
rect 103440 71940 103560 71950
rect 103690 71940 103810 71950
rect 103940 71940 104060 71950
rect 104190 71940 104310 71950
rect 104440 71940 104560 71950
rect 104690 71940 104810 71950
rect 104940 71940 105060 71950
rect 105190 71940 105310 71950
rect 105440 71940 105560 71950
rect 105690 71940 105810 71950
rect 105940 71940 106060 71950
rect 106190 71940 106310 71950
rect 106440 71940 106560 71950
rect 106690 71940 106810 71950
rect 106940 71940 107060 71950
rect 107190 71940 107310 71950
rect 107440 71940 107560 71950
rect 107690 71940 107810 71950
rect 107940 71940 108060 71950
rect 108190 71940 108310 71950
rect 108440 71940 108560 71950
rect 108690 71940 108810 71950
rect 108940 71940 109060 71950
rect 109190 71940 109310 71950
rect 109440 71940 109560 71950
rect 109690 71940 109810 71950
rect 109940 71940 110060 71950
rect 110190 71940 110310 71950
rect 110440 71940 110560 71950
rect 110690 71940 110810 71950
rect 110940 71940 111060 71950
rect 111190 71940 111310 71950
rect 111440 71940 111560 71950
rect 111690 71940 111810 71950
rect 111940 71940 112060 71950
rect 112190 71940 112310 71950
rect 112440 71940 112560 71950
rect 112690 71940 112810 71950
rect 112940 71940 113060 71950
rect 113190 71940 113310 71950
rect 113440 71940 113560 71950
rect 113690 71940 113810 71950
rect 113940 71940 114060 71950
rect 114190 71940 114310 71950
rect 114440 71940 114560 71950
rect 114690 71940 114810 71950
rect 114940 71940 115060 71950
rect 115190 71940 115310 71950
rect 115440 71940 115560 71950
rect 115690 71940 115810 71950
rect 115940 71940 116000 71950
rect 89000 71810 89050 71940
rect 89200 71810 89300 71940
rect 89450 71810 89550 71940
rect 89700 71810 89800 71940
rect 89950 71810 90050 71940
rect 90200 71810 90300 71940
rect 90450 71810 90550 71940
rect 90700 71810 90800 71940
rect 90950 71810 91050 71940
rect 91200 71810 91300 71940
rect 91450 71810 91550 71940
rect 91700 71810 91800 71940
rect 91950 71810 92050 71940
rect 92200 71810 92300 71940
rect 92450 71810 92550 71940
rect 92700 71810 92800 71940
rect 92950 71810 93050 71940
rect 93200 71810 93300 71940
rect 93450 71810 93550 71940
rect 93700 71810 93800 71940
rect 93950 71810 94050 71940
rect 94200 71810 94300 71940
rect 94450 71810 94550 71940
rect 94700 71810 94800 71940
rect 94950 71810 95050 71940
rect 95200 71810 95300 71940
rect 95450 71810 95550 71940
rect 95700 71810 95800 71940
rect 95950 71810 96050 71940
rect 96200 71810 96300 71940
rect 96450 71810 96550 71940
rect 96700 71810 96800 71940
rect 96950 71810 97050 71940
rect 97200 71810 97300 71940
rect 97450 71810 97550 71940
rect 97700 71810 97800 71940
rect 97950 71810 98050 71940
rect 98200 71810 98300 71940
rect 98450 71810 98550 71940
rect 98700 71810 98800 71940
rect 98950 71810 99050 71940
rect 99200 71810 99300 71940
rect 99450 71810 99550 71940
rect 99700 71810 99800 71940
rect 99950 71810 100050 71940
rect 100200 71810 100300 71940
rect 100450 71810 100550 71940
rect 100700 71810 100800 71940
rect 100950 71810 101050 71940
rect 101200 71810 101300 71940
rect 101450 71810 101550 71940
rect 101700 71810 101800 71940
rect 101950 71810 102050 71940
rect 102200 71810 102300 71940
rect 102450 71810 102550 71940
rect 102700 71810 102800 71940
rect 102950 71810 103050 71940
rect 103200 71810 103300 71940
rect 103450 71810 103550 71940
rect 103700 71810 103800 71940
rect 103950 71810 104050 71940
rect 104200 71810 104300 71940
rect 104450 71810 104550 71940
rect 104700 71810 104800 71940
rect 104950 71810 105050 71940
rect 105200 71810 105300 71940
rect 105450 71810 105550 71940
rect 105700 71810 105800 71940
rect 105950 71810 106050 71940
rect 106200 71810 106300 71940
rect 106450 71810 106550 71940
rect 106700 71810 106800 71940
rect 106950 71810 107050 71940
rect 107200 71810 107300 71940
rect 107450 71810 107550 71940
rect 107700 71810 107800 71940
rect 107950 71810 108050 71940
rect 108200 71810 108300 71940
rect 108450 71810 108550 71940
rect 108700 71810 108800 71940
rect 108950 71810 109050 71940
rect 109200 71810 109300 71940
rect 109450 71810 109550 71940
rect 109700 71810 109800 71940
rect 109950 71810 110050 71940
rect 110200 71810 110300 71940
rect 110450 71810 110550 71940
rect 110700 71810 110800 71940
rect 110950 71810 111050 71940
rect 111200 71810 111300 71940
rect 111450 71810 111550 71940
rect 111700 71810 111800 71940
rect 111950 71810 112050 71940
rect 112200 71810 112300 71940
rect 112450 71810 112550 71940
rect 112700 71810 112800 71940
rect 112950 71810 113050 71940
rect 113200 71810 113300 71940
rect 113450 71810 113550 71940
rect 113700 71810 113800 71940
rect 113950 71810 114050 71940
rect 114200 71810 114300 71940
rect 114450 71810 114550 71940
rect 114700 71810 114800 71940
rect 114950 71810 115050 71940
rect 115200 71810 115300 71940
rect 115450 71810 115550 71940
rect 115700 71810 115800 71940
rect 115950 71810 116000 71940
rect 89000 71800 89060 71810
rect 89190 71800 89310 71810
rect 89440 71800 89560 71810
rect 89690 71800 89810 71810
rect 89940 71800 90060 71810
rect 90190 71800 90310 71810
rect 90440 71800 90560 71810
rect 90690 71800 90810 71810
rect 90940 71800 91060 71810
rect 91190 71800 91310 71810
rect 91440 71800 91560 71810
rect 91690 71800 91810 71810
rect 91940 71800 92060 71810
rect 92190 71800 92310 71810
rect 92440 71800 92560 71810
rect 92690 71800 92810 71810
rect 92940 71800 93060 71810
rect 93190 71800 93310 71810
rect 93440 71800 93560 71810
rect 93690 71800 93810 71810
rect 93940 71800 94060 71810
rect 94190 71800 94310 71810
rect 94440 71800 94560 71810
rect 94690 71800 94810 71810
rect 94940 71800 95060 71810
rect 95190 71800 95310 71810
rect 95440 71800 95560 71810
rect 95690 71800 95810 71810
rect 95940 71800 96060 71810
rect 96190 71800 96310 71810
rect 96440 71800 96560 71810
rect 96690 71800 96810 71810
rect 96940 71800 97060 71810
rect 97190 71800 97310 71810
rect 97440 71800 97560 71810
rect 97690 71800 97810 71810
rect 97940 71800 98060 71810
rect 98190 71800 98310 71810
rect 98440 71800 98560 71810
rect 98690 71800 98810 71810
rect 98940 71800 99060 71810
rect 99190 71800 99310 71810
rect 99440 71800 99560 71810
rect 99690 71800 99810 71810
rect 99940 71800 100060 71810
rect 100190 71800 100310 71810
rect 100440 71800 100560 71810
rect 100690 71800 100810 71810
rect 100940 71800 101060 71810
rect 101190 71800 101310 71810
rect 101440 71800 101560 71810
rect 101690 71800 101810 71810
rect 101940 71800 102060 71810
rect 102190 71800 102310 71810
rect 102440 71800 102560 71810
rect 102690 71800 102810 71810
rect 102940 71800 103060 71810
rect 103190 71800 103310 71810
rect 103440 71800 103560 71810
rect 103690 71800 103810 71810
rect 103940 71800 104060 71810
rect 104190 71800 104310 71810
rect 104440 71800 104560 71810
rect 104690 71800 104810 71810
rect 104940 71800 105060 71810
rect 105190 71800 105310 71810
rect 105440 71800 105560 71810
rect 105690 71800 105810 71810
rect 105940 71800 106060 71810
rect 106190 71800 106310 71810
rect 106440 71800 106560 71810
rect 106690 71800 106810 71810
rect 106940 71800 107060 71810
rect 107190 71800 107310 71810
rect 107440 71800 107560 71810
rect 107690 71800 107810 71810
rect 107940 71800 108060 71810
rect 108190 71800 108310 71810
rect 108440 71800 108560 71810
rect 108690 71800 108810 71810
rect 108940 71800 109060 71810
rect 109190 71800 109310 71810
rect 109440 71800 109560 71810
rect 109690 71800 109810 71810
rect 109940 71800 110060 71810
rect 110190 71800 110310 71810
rect 110440 71800 110560 71810
rect 110690 71800 110810 71810
rect 110940 71800 111060 71810
rect 111190 71800 111310 71810
rect 111440 71800 111560 71810
rect 111690 71800 111810 71810
rect 111940 71800 112060 71810
rect 112190 71800 112310 71810
rect 112440 71800 112560 71810
rect 112690 71800 112810 71810
rect 112940 71800 113060 71810
rect 113190 71800 113310 71810
rect 113440 71800 113560 71810
rect 113690 71800 113810 71810
rect 113940 71800 114060 71810
rect 114190 71800 114310 71810
rect 114440 71800 114560 71810
rect 114690 71800 114810 71810
rect 114940 71800 115060 71810
rect 115190 71800 115310 71810
rect 115440 71800 115560 71810
rect 115690 71800 115810 71810
rect 115940 71800 116000 71810
rect 89000 71700 116000 71800
rect 89000 71690 89060 71700
rect 89190 71690 89310 71700
rect 89440 71690 89560 71700
rect 89690 71690 89810 71700
rect 89940 71690 90060 71700
rect 90190 71690 90310 71700
rect 90440 71690 90560 71700
rect 90690 71690 90810 71700
rect 90940 71690 91060 71700
rect 91190 71690 91310 71700
rect 91440 71690 91560 71700
rect 91690 71690 91810 71700
rect 91940 71690 92060 71700
rect 92190 71690 92310 71700
rect 92440 71690 92560 71700
rect 92690 71690 92810 71700
rect 92940 71690 93060 71700
rect 93190 71690 93310 71700
rect 93440 71690 93560 71700
rect 93690 71690 93810 71700
rect 93940 71690 94060 71700
rect 94190 71690 94310 71700
rect 94440 71690 94560 71700
rect 94690 71690 94810 71700
rect 94940 71690 95060 71700
rect 95190 71690 95310 71700
rect 95440 71690 95560 71700
rect 95690 71690 95810 71700
rect 95940 71690 96060 71700
rect 96190 71690 96310 71700
rect 96440 71690 96560 71700
rect 96690 71690 96810 71700
rect 96940 71690 97060 71700
rect 97190 71690 97310 71700
rect 97440 71690 97560 71700
rect 97690 71690 97810 71700
rect 97940 71690 98060 71700
rect 98190 71690 98310 71700
rect 98440 71690 98560 71700
rect 98690 71690 98810 71700
rect 98940 71690 99060 71700
rect 99190 71690 99310 71700
rect 99440 71690 99560 71700
rect 99690 71690 99810 71700
rect 99940 71690 100060 71700
rect 100190 71690 100310 71700
rect 100440 71690 100560 71700
rect 100690 71690 100810 71700
rect 100940 71690 101060 71700
rect 101190 71690 101310 71700
rect 101440 71690 101560 71700
rect 101690 71690 101810 71700
rect 101940 71690 102060 71700
rect 102190 71690 102310 71700
rect 102440 71690 102560 71700
rect 102690 71690 102810 71700
rect 102940 71690 103060 71700
rect 103190 71690 103310 71700
rect 103440 71690 103560 71700
rect 103690 71690 103810 71700
rect 103940 71690 104060 71700
rect 104190 71690 104310 71700
rect 104440 71690 104560 71700
rect 104690 71690 104810 71700
rect 104940 71690 105060 71700
rect 105190 71690 105310 71700
rect 105440 71690 105560 71700
rect 105690 71690 105810 71700
rect 105940 71690 106060 71700
rect 106190 71690 106310 71700
rect 106440 71690 106560 71700
rect 106690 71690 106810 71700
rect 106940 71690 107060 71700
rect 107190 71690 107310 71700
rect 107440 71690 107560 71700
rect 107690 71690 107810 71700
rect 107940 71690 108060 71700
rect 108190 71690 108310 71700
rect 108440 71690 108560 71700
rect 108690 71690 108810 71700
rect 108940 71690 109060 71700
rect 109190 71690 109310 71700
rect 109440 71690 109560 71700
rect 109690 71690 109810 71700
rect 109940 71690 110060 71700
rect 110190 71690 110310 71700
rect 110440 71690 110560 71700
rect 110690 71690 110810 71700
rect 110940 71690 111060 71700
rect 111190 71690 111310 71700
rect 111440 71690 111560 71700
rect 111690 71690 111810 71700
rect 111940 71690 112060 71700
rect 112190 71690 112310 71700
rect 112440 71690 112560 71700
rect 112690 71690 112810 71700
rect 112940 71690 113060 71700
rect 113190 71690 113310 71700
rect 113440 71690 113560 71700
rect 113690 71690 113810 71700
rect 113940 71690 114060 71700
rect 114190 71690 114310 71700
rect 114440 71690 114560 71700
rect 114690 71690 114810 71700
rect 114940 71690 115060 71700
rect 115190 71690 115310 71700
rect 115440 71690 115560 71700
rect 115690 71690 115810 71700
rect 115940 71690 116000 71700
rect 89000 71560 89050 71690
rect 89200 71560 89300 71690
rect 89450 71560 89550 71690
rect 89700 71560 89800 71690
rect 89950 71560 90050 71690
rect 90200 71560 90300 71690
rect 90450 71560 90550 71690
rect 90700 71560 90800 71690
rect 90950 71560 91050 71690
rect 91200 71560 91300 71690
rect 91450 71560 91550 71690
rect 91700 71560 91800 71690
rect 91950 71560 92050 71690
rect 92200 71560 92300 71690
rect 92450 71560 92550 71690
rect 92700 71560 92800 71690
rect 92950 71560 93050 71690
rect 93200 71560 93300 71690
rect 93450 71560 93550 71690
rect 93700 71560 93800 71690
rect 93950 71560 94050 71690
rect 94200 71560 94300 71690
rect 94450 71560 94550 71690
rect 94700 71560 94800 71690
rect 94950 71560 95050 71690
rect 95200 71560 95300 71690
rect 95450 71560 95550 71690
rect 95700 71560 95800 71690
rect 95950 71560 96050 71690
rect 96200 71560 96300 71690
rect 96450 71560 96550 71690
rect 96700 71560 96800 71690
rect 96950 71560 97050 71690
rect 97200 71560 97300 71690
rect 97450 71560 97550 71690
rect 97700 71560 97800 71690
rect 97950 71560 98050 71690
rect 98200 71560 98300 71690
rect 98450 71560 98550 71690
rect 98700 71560 98800 71690
rect 98950 71560 99050 71690
rect 99200 71560 99300 71690
rect 99450 71560 99550 71690
rect 99700 71560 99800 71690
rect 99950 71560 100050 71690
rect 100200 71560 100300 71690
rect 100450 71560 100550 71690
rect 100700 71560 100800 71690
rect 100950 71560 101050 71690
rect 101200 71560 101300 71690
rect 101450 71560 101550 71690
rect 101700 71560 101800 71690
rect 101950 71560 102050 71690
rect 102200 71560 102300 71690
rect 102450 71560 102550 71690
rect 102700 71560 102800 71690
rect 102950 71560 103050 71690
rect 103200 71560 103300 71690
rect 103450 71560 103550 71690
rect 103700 71560 103800 71690
rect 103950 71560 104050 71690
rect 104200 71560 104300 71690
rect 104450 71560 104550 71690
rect 104700 71560 104800 71690
rect 104950 71560 105050 71690
rect 105200 71560 105300 71690
rect 105450 71560 105550 71690
rect 105700 71560 105800 71690
rect 105950 71560 106050 71690
rect 106200 71560 106300 71690
rect 106450 71560 106550 71690
rect 106700 71560 106800 71690
rect 106950 71560 107050 71690
rect 107200 71560 107300 71690
rect 107450 71560 107550 71690
rect 107700 71560 107800 71690
rect 107950 71560 108050 71690
rect 108200 71560 108300 71690
rect 108450 71560 108550 71690
rect 108700 71560 108800 71690
rect 108950 71560 109050 71690
rect 109200 71560 109300 71690
rect 109450 71560 109550 71690
rect 109700 71560 109800 71690
rect 109950 71560 110050 71690
rect 110200 71560 110300 71690
rect 110450 71560 110550 71690
rect 110700 71560 110800 71690
rect 110950 71560 111050 71690
rect 111200 71560 111300 71690
rect 111450 71560 111550 71690
rect 111700 71560 111800 71690
rect 111950 71560 112050 71690
rect 112200 71560 112300 71690
rect 112450 71560 112550 71690
rect 112700 71560 112800 71690
rect 112950 71560 113050 71690
rect 113200 71560 113300 71690
rect 113450 71560 113550 71690
rect 113700 71560 113800 71690
rect 113950 71560 114050 71690
rect 114200 71560 114300 71690
rect 114450 71560 114550 71690
rect 114700 71560 114800 71690
rect 114950 71560 115050 71690
rect 115200 71560 115300 71690
rect 115450 71560 115550 71690
rect 115700 71560 115800 71690
rect 115950 71560 116000 71690
rect 89000 71550 89060 71560
rect 89190 71550 89310 71560
rect 89440 71550 89560 71560
rect 89690 71550 89810 71560
rect 89940 71550 90060 71560
rect 90190 71550 90310 71560
rect 90440 71550 90560 71560
rect 90690 71550 90810 71560
rect 90940 71550 91060 71560
rect 91190 71550 91310 71560
rect 91440 71550 91560 71560
rect 91690 71550 91810 71560
rect 91940 71550 92060 71560
rect 92190 71550 92310 71560
rect 92440 71550 92560 71560
rect 92690 71550 92810 71560
rect 92940 71550 93060 71560
rect 93190 71550 93310 71560
rect 93440 71550 93560 71560
rect 93690 71550 93810 71560
rect 93940 71550 94060 71560
rect 94190 71550 94310 71560
rect 94440 71550 94560 71560
rect 94690 71550 94810 71560
rect 94940 71550 95060 71560
rect 95190 71550 95310 71560
rect 95440 71550 95560 71560
rect 95690 71550 95810 71560
rect 95940 71550 96060 71560
rect 96190 71550 96310 71560
rect 96440 71550 96560 71560
rect 96690 71550 96810 71560
rect 96940 71550 97060 71560
rect 97190 71550 97310 71560
rect 97440 71550 97560 71560
rect 97690 71550 97810 71560
rect 97940 71550 98060 71560
rect 98190 71550 98310 71560
rect 98440 71550 98560 71560
rect 98690 71550 98810 71560
rect 98940 71550 99060 71560
rect 99190 71550 99310 71560
rect 99440 71550 99560 71560
rect 99690 71550 99810 71560
rect 99940 71550 100060 71560
rect 100190 71550 100310 71560
rect 100440 71550 100560 71560
rect 100690 71550 100810 71560
rect 100940 71550 101060 71560
rect 101190 71550 101310 71560
rect 101440 71550 101560 71560
rect 101690 71550 101810 71560
rect 101940 71550 102060 71560
rect 102190 71550 102310 71560
rect 102440 71550 102560 71560
rect 102690 71550 102810 71560
rect 102940 71550 103060 71560
rect 103190 71550 103310 71560
rect 103440 71550 103560 71560
rect 103690 71550 103810 71560
rect 103940 71550 104060 71560
rect 104190 71550 104310 71560
rect 104440 71550 104560 71560
rect 104690 71550 104810 71560
rect 104940 71550 105060 71560
rect 105190 71550 105310 71560
rect 105440 71550 105560 71560
rect 105690 71550 105810 71560
rect 105940 71550 106060 71560
rect 106190 71550 106310 71560
rect 106440 71550 106560 71560
rect 106690 71550 106810 71560
rect 106940 71550 107060 71560
rect 107190 71550 107310 71560
rect 107440 71550 107560 71560
rect 107690 71550 107810 71560
rect 107940 71550 108060 71560
rect 108190 71550 108310 71560
rect 108440 71550 108560 71560
rect 108690 71550 108810 71560
rect 108940 71550 109060 71560
rect 109190 71550 109310 71560
rect 109440 71550 109560 71560
rect 109690 71550 109810 71560
rect 109940 71550 110060 71560
rect 110190 71550 110310 71560
rect 110440 71550 110560 71560
rect 110690 71550 110810 71560
rect 110940 71550 111060 71560
rect 111190 71550 111310 71560
rect 111440 71550 111560 71560
rect 111690 71550 111810 71560
rect 111940 71550 112060 71560
rect 112190 71550 112310 71560
rect 112440 71550 112560 71560
rect 112690 71550 112810 71560
rect 112940 71550 113060 71560
rect 113190 71550 113310 71560
rect 113440 71550 113560 71560
rect 113690 71550 113810 71560
rect 113940 71550 114060 71560
rect 114190 71550 114310 71560
rect 114440 71550 114560 71560
rect 114690 71550 114810 71560
rect 114940 71550 115060 71560
rect 115190 71550 115310 71560
rect 115440 71550 115560 71560
rect 115690 71550 115810 71560
rect 115940 71550 116000 71560
rect 89000 71450 116000 71550
rect 89000 71440 89060 71450
rect 89190 71440 89310 71450
rect 89440 71440 89560 71450
rect 89690 71440 89810 71450
rect 89940 71440 90060 71450
rect 90190 71440 90310 71450
rect 90440 71440 90560 71450
rect 90690 71440 90810 71450
rect 90940 71440 91060 71450
rect 91190 71440 91310 71450
rect 91440 71440 91560 71450
rect 91690 71440 91810 71450
rect 91940 71440 92060 71450
rect 92190 71440 92310 71450
rect 92440 71440 92560 71450
rect 92690 71440 92810 71450
rect 92940 71440 93060 71450
rect 93190 71440 93310 71450
rect 93440 71440 93560 71450
rect 93690 71440 93810 71450
rect 93940 71440 94060 71450
rect 94190 71440 94310 71450
rect 94440 71440 94560 71450
rect 94690 71440 94810 71450
rect 94940 71440 95060 71450
rect 95190 71440 95310 71450
rect 95440 71440 95560 71450
rect 95690 71440 95810 71450
rect 95940 71440 96060 71450
rect 96190 71440 96310 71450
rect 96440 71440 96560 71450
rect 96690 71440 96810 71450
rect 96940 71440 97060 71450
rect 97190 71440 97310 71450
rect 97440 71440 97560 71450
rect 97690 71440 97810 71450
rect 97940 71440 98060 71450
rect 98190 71440 98310 71450
rect 98440 71440 98560 71450
rect 98690 71440 98810 71450
rect 98940 71440 99060 71450
rect 99190 71440 99310 71450
rect 99440 71440 99560 71450
rect 99690 71440 99810 71450
rect 99940 71440 100060 71450
rect 100190 71440 100310 71450
rect 100440 71440 100560 71450
rect 100690 71440 100810 71450
rect 100940 71440 101060 71450
rect 101190 71440 101310 71450
rect 101440 71440 101560 71450
rect 101690 71440 101810 71450
rect 101940 71440 102060 71450
rect 102190 71440 102310 71450
rect 102440 71440 102560 71450
rect 102690 71440 102810 71450
rect 102940 71440 103060 71450
rect 103190 71440 103310 71450
rect 103440 71440 103560 71450
rect 103690 71440 103810 71450
rect 103940 71440 104060 71450
rect 104190 71440 104310 71450
rect 104440 71440 104560 71450
rect 104690 71440 104810 71450
rect 104940 71440 105060 71450
rect 105190 71440 105310 71450
rect 105440 71440 105560 71450
rect 105690 71440 105810 71450
rect 105940 71440 106060 71450
rect 106190 71440 106310 71450
rect 106440 71440 106560 71450
rect 106690 71440 106810 71450
rect 106940 71440 107060 71450
rect 107190 71440 107310 71450
rect 107440 71440 107560 71450
rect 107690 71440 107810 71450
rect 107940 71440 108060 71450
rect 108190 71440 108310 71450
rect 108440 71440 108560 71450
rect 108690 71440 108810 71450
rect 108940 71440 109060 71450
rect 109190 71440 109310 71450
rect 109440 71440 109560 71450
rect 109690 71440 109810 71450
rect 109940 71440 110060 71450
rect 110190 71440 110310 71450
rect 110440 71440 110560 71450
rect 110690 71440 110810 71450
rect 110940 71440 111060 71450
rect 111190 71440 111310 71450
rect 111440 71440 111560 71450
rect 111690 71440 111810 71450
rect 111940 71440 112060 71450
rect 112190 71440 112310 71450
rect 112440 71440 112560 71450
rect 112690 71440 112810 71450
rect 112940 71440 113060 71450
rect 113190 71440 113310 71450
rect 113440 71440 113560 71450
rect 113690 71440 113810 71450
rect 113940 71440 114060 71450
rect 114190 71440 114310 71450
rect 114440 71440 114560 71450
rect 114690 71440 114810 71450
rect 114940 71440 115060 71450
rect 115190 71440 115310 71450
rect 115440 71440 115560 71450
rect 115690 71440 115810 71450
rect 115940 71440 116000 71450
rect 89000 71310 89050 71440
rect 89200 71310 89300 71440
rect 89450 71310 89550 71440
rect 89700 71310 89800 71440
rect 89950 71310 90050 71440
rect 90200 71310 90300 71440
rect 90450 71310 90550 71440
rect 90700 71310 90800 71440
rect 90950 71310 91050 71440
rect 91200 71310 91300 71440
rect 91450 71310 91550 71440
rect 91700 71310 91800 71440
rect 91950 71310 92050 71440
rect 92200 71310 92300 71440
rect 92450 71310 92550 71440
rect 92700 71310 92800 71440
rect 92950 71310 93050 71440
rect 93200 71310 93300 71440
rect 93450 71310 93550 71440
rect 93700 71310 93800 71440
rect 93950 71310 94050 71440
rect 94200 71310 94300 71440
rect 94450 71310 94550 71440
rect 94700 71310 94800 71440
rect 94950 71310 95050 71440
rect 95200 71310 95300 71440
rect 95450 71310 95550 71440
rect 95700 71310 95800 71440
rect 95950 71310 96050 71440
rect 96200 71310 96300 71440
rect 96450 71310 96550 71440
rect 96700 71310 96800 71440
rect 96950 71310 97050 71440
rect 97200 71310 97300 71440
rect 97450 71310 97550 71440
rect 97700 71310 97800 71440
rect 97950 71310 98050 71440
rect 98200 71310 98300 71440
rect 98450 71310 98550 71440
rect 98700 71310 98800 71440
rect 98950 71310 99050 71440
rect 99200 71310 99300 71440
rect 99450 71310 99550 71440
rect 99700 71310 99800 71440
rect 99950 71310 100050 71440
rect 100200 71310 100300 71440
rect 100450 71310 100550 71440
rect 100700 71310 100800 71440
rect 100950 71310 101050 71440
rect 101200 71310 101300 71440
rect 101450 71310 101550 71440
rect 101700 71310 101800 71440
rect 101950 71310 102050 71440
rect 102200 71310 102300 71440
rect 102450 71310 102550 71440
rect 102700 71310 102800 71440
rect 102950 71310 103050 71440
rect 103200 71310 103300 71440
rect 103450 71310 103550 71440
rect 103700 71310 103800 71440
rect 103950 71310 104050 71440
rect 104200 71310 104300 71440
rect 104450 71310 104550 71440
rect 104700 71310 104800 71440
rect 104950 71310 105050 71440
rect 105200 71310 105300 71440
rect 105450 71310 105550 71440
rect 105700 71310 105800 71440
rect 105950 71310 106050 71440
rect 106200 71310 106300 71440
rect 106450 71310 106550 71440
rect 106700 71310 106800 71440
rect 106950 71310 107050 71440
rect 107200 71310 107300 71440
rect 107450 71310 107550 71440
rect 107700 71310 107800 71440
rect 107950 71310 108050 71440
rect 108200 71310 108300 71440
rect 108450 71310 108550 71440
rect 108700 71310 108800 71440
rect 108950 71310 109050 71440
rect 109200 71310 109300 71440
rect 109450 71310 109550 71440
rect 109700 71310 109800 71440
rect 109950 71310 110050 71440
rect 110200 71310 110300 71440
rect 110450 71310 110550 71440
rect 110700 71310 110800 71440
rect 110950 71310 111050 71440
rect 111200 71310 111300 71440
rect 111450 71310 111550 71440
rect 111700 71310 111800 71440
rect 111950 71310 112050 71440
rect 112200 71310 112300 71440
rect 112450 71310 112550 71440
rect 112700 71310 112800 71440
rect 112950 71310 113050 71440
rect 113200 71310 113300 71440
rect 113450 71310 113550 71440
rect 113700 71310 113800 71440
rect 113950 71310 114050 71440
rect 114200 71310 114300 71440
rect 114450 71310 114550 71440
rect 114700 71310 114800 71440
rect 114950 71310 115050 71440
rect 115200 71310 115300 71440
rect 115450 71310 115550 71440
rect 115700 71310 115800 71440
rect 115950 71310 116000 71440
rect 89000 71300 89060 71310
rect 89190 71300 89310 71310
rect 89440 71300 89560 71310
rect 89690 71300 89810 71310
rect 89940 71300 90060 71310
rect 90190 71300 90310 71310
rect 90440 71300 90560 71310
rect 90690 71300 90810 71310
rect 90940 71300 91060 71310
rect 91190 71300 91310 71310
rect 91440 71300 91560 71310
rect 91690 71300 91810 71310
rect 91940 71300 92060 71310
rect 92190 71300 92310 71310
rect 92440 71300 92560 71310
rect 92690 71300 92810 71310
rect 92940 71300 93060 71310
rect 93190 71300 93310 71310
rect 93440 71300 93560 71310
rect 93690 71300 93810 71310
rect 93940 71300 94060 71310
rect 94190 71300 94310 71310
rect 94440 71300 94560 71310
rect 94690 71300 94810 71310
rect 94940 71300 95060 71310
rect 95190 71300 95310 71310
rect 95440 71300 95560 71310
rect 95690 71300 95810 71310
rect 95940 71300 96060 71310
rect 96190 71300 96310 71310
rect 96440 71300 96560 71310
rect 96690 71300 96810 71310
rect 96940 71300 97060 71310
rect 97190 71300 97310 71310
rect 97440 71300 97560 71310
rect 97690 71300 97810 71310
rect 97940 71300 98060 71310
rect 98190 71300 98310 71310
rect 98440 71300 98560 71310
rect 98690 71300 98810 71310
rect 98940 71300 99060 71310
rect 99190 71300 99310 71310
rect 99440 71300 99560 71310
rect 99690 71300 99810 71310
rect 99940 71300 100060 71310
rect 100190 71300 100310 71310
rect 100440 71300 100560 71310
rect 100690 71300 100810 71310
rect 100940 71300 101060 71310
rect 101190 71300 101310 71310
rect 101440 71300 101560 71310
rect 101690 71300 101810 71310
rect 101940 71300 102060 71310
rect 102190 71300 102310 71310
rect 102440 71300 102560 71310
rect 102690 71300 102810 71310
rect 102940 71300 103060 71310
rect 103190 71300 103310 71310
rect 103440 71300 103560 71310
rect 103690 71300 103810 71310
rect 103940 71300 104060 71310
rect 104190 71300 104310 71310
rect 104440 71300 104560 71310
rect 104690 71300 104810 71310
rect 104940 71300 105060 71310
rect 105190 71300 105310 71310
rect 105440 71300 105560 71310
rect 105690 71300 105810 71310
rect 105940 71300 106060 71310
rect 106190 71300 106310 71310
rect 106440 71300 106560 71310
rect 106690 71300 106810 71310
rect 106940 71300 107060 71310
rect 107190 71300 107310 71310
rect 107440 71300 107560 71310
rect 107690 71300 107810 71310
rect 107940 71300 108060 71310
rect 108190 71300 108310 71310
rect 108440 71300 108560 71310
rect 108690 71300 108810 71310
rect 108940 71300 109060 71310
rect 109190 71300 109310 71310
rect 109440 71300 109560 71310
rect 109690 71300 109810 71310
rect 109940 71300 110060 71310
rect 110190 71300 110310 71310
rect 110440 71300 110560 71310
rect 110690 71300 110810 71310
rect 110940 71300 111060 71310
rect 111190 71300 111310 71310
rect 111440 71300 111560 71310
rect 111690 71300 111810 71310
rect 111940 71300 112060 71310
rect 112190 71300 112310 71310
rect 112440 71300 112560 71310
rect 112690 71300 112810 71310
rect 112940 71300 113060 71310
rect 113190 71300 113310 71310
rect 113440 71300 113560 71310
rect 113690 71300 113810 71310
rect 113940 71300 114060 71310
rect 114190 71300 114310 71310
rect 114440 71300 114560 71310
rect 114690 71300 114810 71310
rect 114940 71300 115060 71310
rect 115190 71300 115310 71310
rect 115440 71300 115560 71310
rect 115690 71300 115810 71310
rect 115940 71300 116000 71310
rect 89000 71200 116000 71300
rect 89000 71190 89060 71200
rect 89190 71190 89310 71200
rect 89440 71190 89560 71200
rect 89690 71190 89810 71200
rect 89940 71190 90060 71200
rect 90190 71190 90310 71200
rect 90440 71190 90560 71200
rect 90690 71190 90810 71200
rect 90940 71190 91060 71200
rect 91190 71190 91310 71200
rect 91440 71190 91560 71200
rect 91690 71190 91810 71200
rect 91940 71190 92060 71200
rect 92190 71190 92310 71200
rect 92440 71190 92560 71200
rect 92690 71190 92810 71200
rect 92940 71190 93060 71200
rect 93190 71190 93310 71200
rect 93440 71190 93560 71200
rect 93690 71190 93810 71200
rect 93940 71190 94060 71200
rect 94190 71190 94310 71200
rect 94440 71190 94560 71200
rect 94690 71190 94810 71200
rect 94940 71190 95060 71200
rect 95190 71190 95310 71200
rect 95440 71190 95560 71200
rect 95690 71190 95810 71200
rect 95940 71190 96060 71200
rect 96190 71190 96310 71200
rect 96440 71190 96560 71200
rect 96690 71190 96810 71200
rect 96940 71190 97060 71200
rect 97190 71190 97310 71200
rect 97440 71190 97560 71200
rect 97690 71190 97810 71200
rect 97940 71190 98060 71200
rect 98190 71190 98310 71200
rect 98440 71190 98560 71200
rect 98690 71190 98810 71200
rect 98940 71190 99060 71200
rect 99190 71190 99310 71200
rect 99440 71190 99560 71200
rect 99690 71190 99810 71200
rect 99940 71190 100060 71200
rect 100190 71190 100310 71200
rect 100440 71190 100560 71200
rect 100690 71190 100810 71200
rect 100940 71190 101060 71200
rect 101190 71190 101310 71200
rect 101440 71190 101560 71200
rect 101690 71190 101810 71200
rect 101940 71190 102060 71200
rect 102190 71190 102310 71200
rect 102440 71190 102560 71200
rect 102690 71190 102810 71200
rect 102940 71190 103060 71200
rect 103190 71190 103310 71200
rect 103440 71190 103560 71200
rect 103690 71190 103810 71200
rect 103940 71190 104060 71200
rect 104190 71190 104310 71200
rect 104440 71190 104560 71200
rect 104690 71190 104810 71200
rect 104940 71190 105060 71200
rect 105190 71190 105310 71200
rect 105440 71190 105560 71200
rect 105690 71190 105810 71200
rect 105940 71190 106060 71200
rect 106190 71190 106310 71200
rect 106440 71190 106560 71200
rect 106690 71190 106810 71200
rect 106940 71190 107060 71200
rect 107190 71190 107310 71200
rect 107440 71190 107560 71200
rect 107690 71190 107810 71200
rect 107940 71190 108060 71200
rect 108190 71190 108310 71200
rect 108440 71190 108560 71200
rect 108690 71190 108810 71200
rect 108940 71190 109060 71200
rect 109190 71190 109310 71200
rect 109440 71190 109560 71200
rect 109690 71190 109810 71200
rect 109940 71190 110060 71200
rect 110190 71190 110310 71200
rect 110440 71190 110560 71200
rect 110690 71190 110810 71200
rect 110940 71190 111060 71200
rect 111190 71190 111310 71200
rect 111440 71190 111560 71200
rect 111690 71190 111810 71200
rect 111940 71190 112060 71200
rect 112190 71190 112310 71200
rect 112440 71190 112560 71200
rect 112690 71190 112810 71200
rect 112940 71190 113060 71200
rect 113190 71190 113310 71200
rect 113440 71190 113560 71200
rect 113690 71190 113810 71200
rect 113940 71190 114060 71200
rect 114190 71190 114310 71200
rect 114440 71190 114560 71200
rect 114690 71190 114810 71200
rect 114940 71190 115060 71200
rect 115190 71190 115310 71200
rect 115440 71190 115560 71200
rect 115690 71190 115810 71200
rect 115940 71190 116000 71200
rect 89000 71060 89050 71190
rect 89200 71060 89300 71190
rect 89450 71060 89550 71190
rect 89700 71060 89800 71190
rect 89950 71060 90050 71190
rect 90200 71060 90300 71190
rect 90450 71060 90550 71190
rect 90700 71060 90800 71190
rect 90950 71060 91050 71190
rect 91200 71060 91300 71190
rect 91450 71060 91550 71190
rect 91700 71060 91800 71190
rect 91950 71060 92050 71190
rect 92200 71060 92300 71190
rect 92450 71060 92550 71190
rect 92700 71060 92800 71190
rect 92950 71060 93050 71190
rect 93200 71060 93300 71190
rect 93450 71060 93550 71190
rect 93700 71060 93800 71190
rect 93950 71060 94050 71190
rect 94200 71060 94300 71190
rect 94450 71060 94550 71190
rect 94700 71060 94800 71190
rect 94950 71060 95050 71190
rect 95200 71060 95300 71190
rect 95450 71060 95550 71190
rect 95700 71060 95800 71190
rect 95950 71060 96050 71190
rect 96200 71060 96300 71190
rect 96450 71060 96550 71190
rect 96700 71060 96800 71190
rect 96950 71060 97050 71190
rect 97200 71060 97300 71190
rect 97450 71060 97550 71190
rect 97700 71060 97800 71190
rect 97950 71060 98050 71190
rect 98200 71060 98300 71190
rect 98450 71060 98550 71190
rect 98700 71060 98800 71190
rect 98950 71060 99050 71190
rect 99200 71060 99300 71190
rect 99450 71060 99550 71190
rect 99700 71060 99800 71190
rect 99950 71060 100050 71190
rect 100200 71060 100300 71190
rect 100450 71060 100550 71190
rect 100700 71060 100800 71190
rect 100950 71060 101050 71190
rect 101200 71060 101300 71190
rect 101450 71060 101550 71190
rect 101700 71060 101800 71190
rect 101950 71060 102050 71190
rect 102200 71060 102300 71190
rect 102450 71060 102550 71190
rect 102700 71060 102800 71190
rect 102950 71060 103050 71190
rect 103200 71060 103300 71190
rect 103450 71060 103550 71190
rect 103700 71060 103800 71190
rect 103950 71060 104050 71190
rect 104200 71060 104300 71190
rect 104450 71060 104550 71190
rect 104700 71060 104800 71190
rect 104950 71060 105050 71190
rect 105200 71060 105300 71190
rect 105450 71060 105550 71190
rect 105700 71060 105800 71190
rect 105950 71060 106050 71190
rect 106200 71060 106300 71190
rect 106450 71060 106550 71190
rect 106700 71060 106800 71190
rect 106950 71060 107050 71190
rect 107200 71060 107300 71190
rect 107450 71060 107550 71190
rect 107700 71060 107800 71190
rect 107950 71060 108050 71190
rect 108200 71060 108300 71190
rect 108450 71060 108550 71190
rect 108700 71060 108800 71190
rect 108950 71060 109050 71190
rect 109200 71060 109300 71190
rect 109450 71060 109550 71190
rect 109700 71060 109800 71190
rect 109950 71060 110050 71190
rect 110200 71060 110300 71190
rect 110450 71060 110550 71190
rect 110700 71060 110800 71190
rect 110950 71060 111050 71190
rect 111200 71060 111300 71190
rect 111450 71060 111550 71190
rect 111700 71060 111800 71190
rect 111950 71060 112050 71190
rect 112200 71060 112300 71190
rect 112450 71060 112550 71190
rect 112700 71060 112800 71190
rect 112950 71060 113050 71190
rect 113200 71060 113300 71190
rect 113450 71060 113550 71190
rect 113700 71060 113800 71190
rect 113950 71060 114050 71190
rect 114200 71060 114300 71190
rect 114450 71060 114550 71190
rect 114700 71060 114800 71190
rect 114950 71060 115050 71190
rect 115200 71060 115300 71190
rect 115450 71060 115550 71190
rect 115700 71060 115800 71190
rect 115950 71060 116000 71190
rect 89000 71050 89060 71060
rect 89190 71050 89310 71060
rect 89440 71050 89560 71060
rect 89690 71050 89810 71060
rect 89940 71050 90060 71060
rect 90190 71050 90310 71060
rect 90440 71050 90560 71060
rect 90690 71050 90810 71060
rect 90940 71050 91060 71060
rect 91190 71050 91310 71060
rect 91440 71050 91560 71060
rect 91690 71050 91810 71060
rect 91940 71050 92060 71060
rect 92190 71050 92310 71060
rect 92440 71050 92560 71060
rect 92690 71050 92810 71060
rect 92940 71050 93060 71060
rect 93190 71050 93310 71060
rect 93440 71050 93560 71060
rect 93690 71050 93810 71060
rect 93940 71050 94060 71060
rect 94190 71050 94310 71060
rect 94440 71050 94560 71060
rect 94690 71050 94810 71060
rect 94940 71050 95060 71060
rect 95190 71050 95310 71060
rect 95440 71050 95560 71060
rect 95690 71050 95810 71060
rect 95940 71050 96060 71060
rect 96190 71050 96310 71060
rect 96440 71050 96560 71060
rect 96690 71050 96810 71060
rect 96940 71050 97060 71060
rect 97190 71050 97310 71060
rect 97440 71050 97560 71060
rect 97690 71050 97810 71060
rect 97940 71050 98060 71060
rect 98190 71050 98310 71060
rect 98440 71050 98560 71060
rect 98690 71050 98810 71060
rect 98940 71050 99060 71060
rect 99190 71050 99310 71060
rect 99440 71050 99560 71060
rect 99690 71050 99810 71060
rect 99940 71050 100060 71060
rect 100190 71050 100310 71060
rect 100440 71050 100560 71060
rect 100690 71050 100810 71060
rect 100940 71050 101060 71060
rect 101190 71050 101310 71060
rect 101440 71050 101560 71060
rect 101690 71050 101810 71060
rect 101940 71050 102060 71060
rect 102190 71050 102310 71060
rect 102440 71050 102560 71060
rect 102690 71050 102810 71060
rect 102940 71050 103060 71060
rect 103190 71050 103310 71060
rect 103440 71050 103560 71060
rect 103690 71050 103810 71060
rect 103940 71050 104060 71060
rect 104190 71050 104310 71060
rect 104440 71050 104560 71060
rect 104690 71050 104810 71060
rect 104940 71050 105060 71060
rect 105190 71050 105310 71060
rect 105440 71050 105560 71060
rect 105690 71050 105810 71060
rect 105940 71050 106060 71060
rect 106190 71050 106310 71060
rect 106440 71050 106560 71060
rect 106690 71050 106810 71060
rect 106940 71050 107060 71060
rect 107190 71050 107310 71060
rect 107440 71050 107560 71060
rect 107690 71050 107810 71060
rect 107940 71050 108060 71060
rect 108190 71050 108310 71060
rect 108440 71050 108560 71060
rect 108690 71050 108810 71060
rect 108940 71050 109060 71060
rect 109190 71050 109310 71060
rect 109440 71050 109560 71060
rect 109690 71050 109810 71060
rect 109940 71050 110060 71060
rect 110190 71050 110310 71060
rect 110440 71050 110560 71060
rect 110690 71050 110810 71060
rect 110940 71050 111060 71060
rect 111190 71050 111310 71060
rect 111440 71050 111560 71060
rect 111690 71050 111810 71060
rect 111940 71050 112060 71060
rect 112190 71050 112310 71060
rect 112440 71050 112560 71060
rect 112690 71050 112810 71060
rect 112940 71050 113060 71060
rect 113190 71050 113310 71060
rect 113440 71050 113560 71060
rect 113690 71050 113810 71060
rect 113940 71050 114060 71060
rect 114190 71050 114310 71060
rect 114440 71050 114560 71060
rect 114690 71050 114810 71060
rect 114940 71050 115060 71060
rect 115190 71050 115310 71060
rect 115440 71050 115560 71060
rect 115690 71050 115810 71060
rect 115940 71050 116000 71060
rect 89000 71000 116000 71050
<< metal3 >>
rect 8000 80900 11000 82000
rect 34097 81900 36597 82000
rect 34097 81150 36600 81900
rect 34100 81000 36600 81150
rect 8000 78100 8100 80900
rect 10900 78100 11000 80900
rect 8000 78000 11000 78100
rect 60000 80900 63000 82000
rect 82797 81150 85297 82000
rect 85447 81150 86547 82000
rect 86697 81150 87797 82000
rect 87947 81150 90447 82000
rect 108647 81150 111147 82000
rect 111297 81150 112397 82000
rect 112547 81150 113647 82000
rect 113797 81150 116297 82000
rect 159497 81150 161997 82000
rect 162147 81150 163247 82000
rect 163397 81150 164497 82000
rect 164647 81150 167147 82000
rect 206697 81150 209197 82000
rect 232697 81150 235197 82000
rect 255297 81170 257697 82000
rect 260297 81170 262697 82000
rect 283297 81150 285797 82000
rect 60000 78100 60100 80900
rect 62900 78100 63000 80900
rect 60000 78000 63000 78100
rect 83000 80900 85000 81150
rect 83000 77600 83100 80900
rect 84900 77600 85000 80900
rect 83000 77500 85000 77600
rect 109000 80900 111000 81150
rect 109000 77600 109100 80900
rect 110900 77600 111000 80900
rect 109000 77500 111000 77600
rect 0 70121 850 72621
rect 291150 68992 292000 71492
rect 0 51921 830 54321
rect 291170 49892 292000 52292
rect 0 46921 830 49321
rect 291170 44892 292000 47292
rect 291760 24736 292400 24792
rect 291760 24145 292400 24201
rect 291760 23554 292400 23610
rect 291760 22963 292400 23019
rect 291760 22372 292400 22428
rect 291760 21781 292400 21837
rect 0 9721 830 12121
rect 0 4721 830 7121
rect 291170 5281 292000 7681
rect 291170 281 292000 2681
rect 10000 0 10056 200
rect 13100 0 13156 200
rect 16200 0 16256 200
rect 19300 0 19356 200
rect 22400 0 22456 200
rect 25500 0 25556 200
rect 28600 0 28656 200
rect 31700 0 31756 200
rect 34800 0 34856 200
rect 37900 0 37956 200
rect 41000 0 41056 200
rect 44100 0 44156 200
rect 47200 0 47256 200
rect 50300 0 50356 200
rect 53400 0 53456 200
rect 56500 0 56556 200
rect 59600 0 59656 200
rect 62700 0 62756 200
rect 65800 0 65856 200
rect 68900 0 68956 200
rect 72000 0 72056 200
rect 75100 0 75156 200
rect 78200 0 78256 200
rect 81300 0 81356 200
rect 84400 0 84456 200
rect 87500 0 87556 200
rect 90600 0 90656 200
rect 93700 0 93756 200
rect 96800 0 96856 200
rect 99900 0 99956 200
rect 103000 0 103056 200
rect 106100 0 106156 200
rect 109200 0 109256 200
rect 112300 0 112356 200
rect 115400 0 115456 200
rect 118500 0 118556 200
rect 121600 0 121656 200
rect 124700 0 124756 200
rect 127800 0 127856 200
rect 130900 0 130956 200
rect 134000 0 134056 200
rect 137100 0 137156 200
rect 140200 0 140256 200
rect 143300 0 143356 200
rect 146400 0 146456 200
rect 149500 0 149556 200
rect 152600 0 152656 200
rect 155700 0 155756 200
rect 158800 0 158856 200
rect 161900 0 161956 200
rect 165000 0 165056 200
rect 168100 0 168156 200
rect 171200 0 171256 200
rect 174300 0 174356 200
rect 177400 0 177456 200
rect 180500 0 180556 200
rect 183600 0 183656 200
rect 186700 0 186756 200
rect 189800 0 189856 200
rect 192900 0 192956 200
<< via3 >>
rect 8100 78100 10900 80900
rect 60100 78100 62900 80900
rect 83100 77600 84900 80900
rect 109100 77600 110900 80900
<< metal4 >>
rect 8000 80900 11000 81000
rect 8000 78100 8100 80900
rect 10900 78100 11000 80900
rect 8000 78000 11000 78100
rect 60000 80900 63000 81000
rect 60000 78100 60100 80900
rect 62900 78100 63000 80900
rect 60000 78000 63000 78100
rect 83000 80900 85000 81000
rect 83000 77600 83100 80900
rect 84900 77600 85000 80900
rect 83000 75000 85000 77600
rect 109000 80900 111000 81000
rect 109000 77600 109100 80900
rect 110900 77600 111000 80900
rect 109000 74000 111000 77600
rect 85000 72500 111000 74000
rect 3049 0 6899 400
rect 7229 0 11079 400
rect 282049 0 285899 400
rect 286229 0 290079 400
<< via4 >>
rect 8100 78100 10900 80900
rect 60100 78100 62900 80900
<< metal5 >>
rect 8000 80900 11000 81000
rect 8000 78100 8100 80900
rect 10900 80000 11000 80900
rect 60000 80900 63000 81000
rect 10900 78100 28000 80000
rect 8000 78000 28000 78100
rect 60000 78100 60100 80900
rect 62900 80000 63000 80900
rect 62900 78100 69000 80000
rect 60000 78000 69000 78100
rect 26000 75000 28000 78000
rect 67000 75000 69000 78000
use RX_top  RX_top_0
timestamp 1662014484
transform 1 0 19000 0 -1 70000
box -18500 -11900 84000 70000
use TX_top  TX_top_0
timestamp 1661836362
transform 1 0 193750 0 -1 61900
box -41750 -18100 48250 27950
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501637
transform 1 0 5000 0 -1 81000
box 0 0 2000 2000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_38
timestamp 1659501637
transform 1 0 5000 0 -1 79000
box 0 0 2000 2000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660792292
transform 1 0 33000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_1
timestamp 1660792292
transform 1 0 37000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_2
timestamp 1660792292
transform 1 0 41000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_3
timestamp 1660792292
transform 1 0 45000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_4
timestamp 1660792292
transform 1 0 49000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_5
timestamp 1660792292
transform 1 0 53000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_6
timestamp 1660792292
transform 1 0 55000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_7
timestamp 1660792292
transform 1 0 71000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_8
timestamp 1660792292
transform 1 0 75000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_9
timestamp 1660792292
transform 1 0 77000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_10
timestamp 1660792292
transform 1 0 97000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_11
timestamp 1660792292
transform 1 0 93000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_12
timestamp 1660792292
transform 1 0 91000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_13
timestamp 1660792292
transform 1 0 101000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_14
timestamp 1660792292
transform 1 0 103000 0 -1 81000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_70
timestamp 1660792292
transform 1 0 29000 0 -1 81000
box 0 0 4000 4000
<< labels >>
rlabel metal3 s 10000 0 10056 200 0 analog_la_out[0]
port 1 nsew
rlabel metal3 s 13100 0 13156 200 0 analog_la_out[1]
port 2 nsew
rlabel metal3 s 16200 0 16256 200 0 analog_la_out[2]
port 3 nsew
rlabel metal3 s 19300 0 19356 200 0 analog_la_out[3]
port 4 nsew
rlabel metal3 s 22400 0 22456 200 0 analog_la_out[4]
port 5 nsew
rlabel metal3 s 25500 0 25556 200 0 analog_la_out[5]
port 6 nsew
rlabel metal3 s 28600 0 28656 200 0 analog_la_out[6]
port 7 nsew
rlabel metal3 s 31700 0 31756 200 0 analog_la_out[7]
port 8 nsew
rlabel metal3 s 34800 0 34856 200 0 analog_la_out[8]
port 9 nsew
rlabel metal3 s 37900 0 37956 200 0 analog_la_out[9]
port 10 nsew
rlabel metal3 s 41000 0 41056 200 0 analog_la_out[10]
port 11 nsew
rlabel metal3 s 44100 0 44156 200 0 analog_la_out[11]
port 12 nsew
rlabel metal3 s 47200 0 47256 200 0 analog_la_out[12]
port 13 nsew
rlabel metal3 s 50300 0 50356 200 0 analog_la_out[13]
port 14 nsew
rlabel metal3 s 53400 0 53456 200 0 analog_la_out[14]
port 15 nsew
rlabel metal3 s 56500 0 56556 200 0 analog_la_out[15]
port 16 nsew
rlabel metal3 s 59600 0 59656 200 0 analog_la_out[16]
port 17 nsew
rlabel metal3 s 62700 0 62756 200 0 analog_la_out[17]
port 18 nsew
rlabel metal3 s 65800 0 65856 200 0 analog_la_out[18]
port 19 nsew
rlabel metal3 s 68900 0 68956 200 0 analog_la_out[19]
port 20 nsew
rlabel metal3 s 72000 0 72056 200 0 analog_la_out[20]
port 21 nsew
rlabel metal3 s 75100 0 75156 200 0 analog_la_out[21]
port 22 nsew
rlabel metal3 s 78200 0 78256 200 0 analog_la_out[22]
port 23 nsew
rlabel metal3 s 81300 0 81356 200 0 analog_la_out[23]
port 24 nsew
rlabel metal3 s 84400 0 84456 200 0 analog_la_out[24]
port 25 nsew
rlabel metal3 s 87500 0 87556 200 0 analog_la_out[25]
port 26 nsew
rlabel metal3 s 90600 0 90656 200 0 analog_la_out[26]
port 27 nsew
rlabel metal3 s 93700 0 93756 200 0 analog_la_out[27]
port 28 nsew
rlabel metal3 s 96800 0 96856 200 0 analog_la_out[28]
port 29 nsew
rlabel metal3 s 99900 0 99956 200 0 analog_la_out[29]
port 30 nsew
rlabel metal3 s 103000 0 103056 200 0 analog_la_in[0]
port 31 nsew
rlabel metal3 s 106100 0 106156 200 0 analog_la_in[1]
port 32 nsew
rlabel metal3 s 109200 0 109256 200 0 analog_la_in[2]
port 33 nsew
rlabel metal3 s 112300 0 112356 200 0 analog_la_in[3]
port 34 nsew
rlabel metal3 s 115400 0 115456 200 0 analog_la_in[4]
port 35 nsew
rlabel metal3 s 118500 0 118556 200 0 analog_la_in[5]
port 36 nsew
rlabel metal3 s 121600 0 121656 200 0 analog_la_in[6]
port 37 nsew
rlabel metal3 s 124700 0 124756 200 0 analog_la_in[7]
port 38 nsew
rlabel metal3 s 127800 0 127856 200 0 analog_la_in[8]
port 39 nsew
rlabel metal3 s 130900 0 130956 200 0 analog_la_in[9]
port 40 nsew
rlabel metal3 s 134000 0 134056 200 0 analog_la_in[10]
port 41 nsew
rlabel metal3 s 137100 0 137156 200 0 analog_la_in[11]
port 42 nsew
rlabel metal3 s 140200 0 140256 200 0 analog_la_in[12]
port 43 nsew
rlabel metal3 s 143300 0 143356 200 0 analog_la_in[13]
port 44 nsew
rlabel metal3 s 146400 0 146456 200 0 analog_la_in[14]
port 45 nsew
rlabel metal3 s 149500 0 149556 200 0 analog_la_in[15]
port 46 nsew
rlabel metal3 s 152600 0 152656 200 0 analog_la_in[16]
port 47 nsew
rlabel metal3 s 155700 0 155756 200 0 analog_la_in[17]
port 48 nsew
rlabel metal3 s 158800 0 158856 200 0 analog_la_in[18]
port 49 nsew
rlabel metal3 s 161900 0 161956 200 0 analog_la_in[19]
port 50 nsew
rlabel metal3 s 165000 0 165056 200 0 analog_la_in[20]
port 51 nsew
rlabel metal3 s 168100 0 168156 200 0 analog_la_in[21]
port 52 nsew
rlabel metal3 s 171200 0 171256 200 0 analog_la_in[22]
port 53 nsew
rlabel metal3 s 174300 0 174356 200 0 analog_la_in[23]
port 54 nsew
rlabel metal3 s 177400 0 177456 200 0 analog_la_in[24]
port 55 nsew
rlabel metal3 s 180500 0 180556 200 0 analog_la_in[25]
port 56 nsew
rlabel metal3 s 183600 0 183656 200 0 analog_la_in[26]
port 57 nsew
rlabel metal3 s 186700 0 186756 200 0 analog_la_in[27]
port 58 nsew
rlabel metal3 s 189800 0 189856 200 0 analog_la_in[28]
port 59 nsew
rlabel metal3 s 192900 0 192956 200 0 analog_la_in[29]
port 60 nsew
rlabel metal3 s 291760 21781 292400 21837 0 gpio_analog[6]
port 61 nsew
rlabel metal3 s 291760 22372 292400 22428 0 gpio_noesd[6]
port 62 nsew
rlabel metal3 s 291150 68992 292000 71492 0 io_analog[0]
port 63 nsew
rlabel metal3 s 0 70121 850 72621 0 io_analog[10]
port 64 nsew
rlabel metal3 s 283297 81150 285797 82000 0 io_analog[1]
port 65 nsew
rlabel metal3 s 232697 81150 235197 82000 0 io_analog[2]
port 66 nsew
rlabel metal3 s 206697 81150 209197 82000 0 io_analog[3]
port 67 nsew
rlabel metal3 s 159497 81150 161997 82000 0 io_analog[4]
port 68 nsew
rlabel metal3 s 108647 81150 111147 82000 0 io_analog[5]
port 69 nsew
rlabel metal3 s 82797 81150 85297 82000 0 io_analog[6]
port 70 nsew
rlabel metal3 s 60097 81150 62597 82000 0 io_analog[7]
port 71 nsew
rlabel metal3 s 34097 81150 36597 82000 0 io_analog[8]
port 72 nsew
rlabel metal3 s 8097 81150 10597 82000 0 io_analog[9]
port 73 nsew
rlabel metal3 s 163397 81150 164497 82000 0 io_clamp_high[0]
port 74 nsew
rlabel metal3 s 112547 81150 113647 82000 0 io_clamp_high[1]
port 75 nsew
rlabel metal3 s 86697 81150 87797 82000 0 io_clamp_high[2]
port 76 nsew
rlabel metal3 s 162147 81150 163247 82000 0 io_clamp_low[0]
port 77 nsew
rlabel metal3 s 111297 81150 112397 82000 0 io_clamp_low[1]
port 78 nsew
rlabel metal3 s 85447 81150 86547 82000 0 io_clamp_low[2]
port 79 nsew
rlabel metal3 s 291760 23554 292400 23610 0 io_in[13]
port 80 nsew
rlabel metal3 s 291760 22963 292400 23019 0 io_in_3v3[13]
port 81 nsew
rlabel metal3 s 291760 24736 292400 24792 0 io_oeb[13]
port 82 nsew
rlabel metal3 s 291760 24145 292400 24201 0 io_out[13]
port 83 nsew
rlabel metal3 s 291170 44892 292000 47292 0 vccd1
port 84 nsew
rlabel metal3 s 0 46921 830 49321 0 vccd2
port 85 nsew
rlabel metal3 s 291170 5281 292000 7681 0 vdda1
port 86 nsew
rlabel metal3 s 255297 81170 257697 82000 0 vssa1
port 87 nsew
rlabel metal3 s 0 4721 830 7121 0 vssa2
port 88 nsew
rlabel metal4 s 282049 0 285899 400 0 vdda1
port 86 nsew
rlabel metal4 s 286229 0 290079 400 0 vssa1
port 87 nsew
rlabel metal4 s 3049 0 6899 400 0 vdda2
port 89 nsew
rlabel metal4 s 7229 0 11079 400 0 vssd2
port 90 nsew
<< properties >>
string FIXED_BBOX 0 0 292000 82000
string path 1929.280 0.000 1929.280 2.000 
<< end >>
