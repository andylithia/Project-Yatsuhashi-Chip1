magic
tech sky130A
timestamp 1658634298
<< metal1 >>
rect -162 -135 246 -35
<< end >>
