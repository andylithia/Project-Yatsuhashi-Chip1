magic
tech sky130B
magscale 1 2
timestamp 1660524083
<< metal4 >>
rect -17900 -2112 -7500 -2000
rect -17900 -3888 -17788 -2112
rect -16012 -3888 -9388 -2112
rect -7612 -3888 -7500 -2112
rect -17900 -4000 -7500 -3888
<< via4 >>
rect -17788 -3888 -16012 -2112
rect -9388 -3888 -7612 -2112
<< metal5 >>
tri -10100 12237 -8337 14000 se
rect -8337 12237 5737 14000
tri 5737 12237 7500 14000 sw
tri -10337 12000 -10100 12237 se
rect -10100 12000 7500 12237
tri 7500 12000 7737 12237 sw
tri -11012 11325 -10337 12000 se
rect -10337 11400 -8109 12000
tri -8109 11400 -7509 12000 nw
tri 4909 11400 5509 12000 ne
rect 5509 11400 7737 12000
rect -10337 11325 -8184 11400
tri -8184 11325 -8109 11400 nw
tri -7336 11325 -7261 11400 se
rect -7261 11325 4661 11400
tri -12700 9637 -11012 11325 se
rect -11012 10477 -9032 11325
tri -9032 10477 -8184 11325 nw
tri -8184 10477 -7336 11325 se
rect -7336 10552 4661 11325
tri 4661 10552 5509 11400 sw
tri 5509 10552 6357 11400 ne
rect 6357 10552 7737 11400
rect -7336 10477 5509 10552
tri 5509 10477 5584 10552 sw
tri 6357 10477 6432 10552 ne
rect 6432 10477 7737 10552
rect -11012 9637 -9880 10477
tri -12928 9409 -12700 9637 se
rect -12700 9629 -9880 9637
tri -9880 9629 -9032 10477 nw
tri -9032 9629 -8184 10477 se
rect -8184 10248 5584 10477
tri 5584 10248 5813 10477 sw
tri 6432 10248 6661 10477 ne
rect 6661 10248 7737 10477
rect -8184 9629 5813 10248
rect -12700 9409 -10100 9629
tri -10100 9409 -9880 9629 nw
tri -9252 9409 -9032 9629 se
rect -9032 9409 5813 9629
tri -15300 7037 -12928 9409 se
rect -12928 9400 -10109 9409
tri -10109 9400 -10100 9409 nw
tri -9261 9400 -9252 9409 se
rect -9252 9400 5813 9409
tri 5813 9400 6661 10248 sw
tri 6661 9400 7509 10248 ne
rect 7509 9400 7737 10248
tri 7737 9400 10337 12000 sw
rect -12928 8561 -10948 9400
tri -10948 8561 -10109 9400 nw
tri -10100 8561 -9261 9400 se
rect -9261 8800 -7032 9400
tri -7032 8800 -6432 9400 nw
tri 3832 8800 4432 9400 ne
rect 4432 8800 6661 9400
rect -9261 8561 -7880 8800
rect -12928 7713 -11796 8561
tri -11796 7713 -10948 8561 nw
tri -10948 7713 -10100 8561 se
rect -10100 7952 -7880 8561
tri -7880 7952 -7032 8800 nw
tri -7032 7952 -6184 8800 se
rect -6184 7952 3584 8800
tri 3584 7952 4432 8800 sw
tri 4432 7952 5280 8800 ne
rect 5280 8552 6661 8800
tri 6661 8552 7509 9400 sw
tri 7509 8552 8357 9400 ne
rect 8357 8552 10337 9400
rect 5280 8496 7509 8552
tri 7509 8496 7565 8552 sw
tri 8357 8496 8413 8552 ne
rect 8413 8496 10337 8552
rect 5280 7952 7565 8496
rect -10100 7713 -8184 7952
rect -12928 7648 -11861 7713
tri -11861 7648 -11796 7713 nw
tri -11013 7648 -10948 7713 se
rect -10948 7648 -8184 7713
tri -8184 7648 -7880 7952 nw
tri -7336 7648 -7032 7952 se
rect -7032 7648 4432 7952
tri 4432 7648 4736 7952 sw
tri 5280 7648 5584 7952 ne
rect 5584 7648 7565 7952
tri 7565 7648 8413 8496 sw
tri 8413 7648 9261 8496 ne
rect 9261 7648 10337 8496
rect -12928 7037 -12700 7648
tri -15528 6809 -15300 7037 se
rect -15300 6809 -12700 7037
tri -12700 6809 -11861 7648 nw
tri -11852 6809 -11013 7648 se
rect -11013 6809 -9032 7648
tri -17300 5037 -15528 6809 se
rect -15528 5961 -13548 6809
tri -13548 5961 -12700 6809 nw
tri -12700 5961 -11852 6809 se
rect -11852 6800 -9032 6809
tri -9032 6800 -8184 7648 nw
tri -8184 6800 -7336 7648 se
rect -7336 6800 4736 7648
tri 4736 6800 5584 7648 sw
tri 5584 6800 6432 7648 ne
rect 6432 6800 8413 7648
tri 8413 6800 9261 7648 sw
tri 9261 6800 10109 7648 ne
rect 10109 6800 10337 7648
tri 10337 6800 12937 9400 sw
rect -11852 5961 -9880 6800
rect -15528 5732 -13777 5961
tri -13777 5732 -13548 5961 nw
tri -12929 5732 -12700 5961 se
rect -12700 5952 -9880 5961
tri -9880 5952 -9032 6800 nw
tri -9032 5952 -8184 6800 se
rect -8184 5952 -7271 6800
rect -12700 5732 -10100 5952
tri -10100 5732 -9880 5952 nw
tri -9252 5732 -9032 5952 se
rect -9032 5732 -7271 5952
rect -15528 5037 -14625 5732
rect -17300 4884 -14625 5037
tri -14625 4884 -13777 5732 nw
tri -13777 4884 -12929 5732 se
rect -12929 4884 -10948 5732
tri -10948 4884 -10100 5732 nw
tri -10100 4884 -9252 5732 se
rect -9252 4884 -7271 5732
tri -7271 4884 -5355 6800 nw
tri 2755 4884 4671 6800 ne
rect 4671 5952 5584 6800
tri 5584 5952 6432 6800 sw
tri 6432 5952 7280 6800 ne
rect 7280 5952 9261 6800
tri 9261 5952 10109 6800 sw
tri 10109 5952 10957 6800 ne
rect 10957 5952 12937 6800
rect 4671 5732 6432 5952
tri 6432 5732 6652 5952 sw
tri 7280 5732 7500 5952 ne
rect 7500 5732 10109 5952
tri 10109 5732 10329 5952 sw
tri 10957 5732 11177 5952 ne
rect 11177 5732 12937 5952
rect 4671 4884 6652 5732
tri 6652 4884 7500 5732 sw
tri 7500 4884 8348 5732 ne
rect 8348 4884 10329 5732
tri 10329 4884 11177 5732 sw
tri 11177 4884 12025 5732 ne
rect 12025 5037 12937 5732
tri 12937 5037 14700 6800 sw
rect 12025 4884 14700 5037
rect -17300 4809 -14700 4884
tri -14700 4809 -14625 4884 nw
tri -13852 4809 -13777 4884 se
rect -13777 4809 -11796 4884
rect -17300 4000 -15300 4809
tri -15300 4209 -14700 4809 nw
tri -14452 4209 -13852 4809 se
rect -13852 4209 -11796 4809
tri -14661 4000 -14452 4209 se
rect -14452 4036 -11796 4209
tri -11796 4036 -10948 4884 nw
tri -10948 4036 -10100 4884 se
rect -10100 4036 -8155 4884
rect -14452 4000 -11832 4036
tri -11832 4000 -11796 4036 nw
tri -10984 4000 -10948 4036 se
rect -10948 4000 -8155 4036
tri -8155 4000 -7271 4884 nw
tri 4671 4000 5555 4884 ne
rect 5555 4036 7500 4884
tri 7500 4036 8348 4884 sw
tri 8348 4036 9196 4884 ne
rect 9196 4809 11177 4884
tri 11177 4809 11252 4884 sw
tri 12025 4809 12100 4884 ne
rect 12100 4809 14700 4884
rect 9196 4209 11252 4809
tri 11252 4209 11852 4809 sw
tri 12100 4209 12700 4809 ne
rect 9196 4036 11852 4209
rect 5555 4000 8348 4036
rect -19300 2000 -15300 4000
tri -14700 3961 -14661 4000 se
rect -14661 3971 -11861 4000
tri -11861 3971 -11832 4000 nw
tri -11013 3971 -10984 4000 se
rect -10984 3971 -8184 4000
tri -8184 3971 -8155 4000 nw
tri 5555 3971 5584 4000 ne
rect 5584 3971 8348 4000
rect -14661 3961 -12100 3971
rect -14700 3732 -12100 3961
tri -12100 3732 -11861 3971 nw
tri -11252 3732 -11013 3971 se
rect -11013 3732 -10100 3971
rect -17900 -2112 -15900 -2000
rect -17900 -3888 -17788 -2112
rect -16012 -3888 -15900 -2112
rect -17900 -4000 -15900 -3888
rect -14700 -5571 -12700 3732
tri -12700 3132 -12100 3732 nw
tri -11852 3132 -11252 3732 se
rect -11252 3132 -10100 3732
tri -12100 2884 -11852 3132 se
rect -11852 2884 -10100 3132
rect -12100 -4494 -10100 2884
tri -10100 2055 -8184 3971 nw
tri 5584 2055 7500 3971 ne
rect 7500 3732 8348 3971
tri 8348 3732 8652 4036 sw
tri 9196 3732 9500 4036 ne
rect 9500 3961 11852 4036
tri 11852 3961 12100 4209 sw
rect 9500 3732 12100 3961
rect 7500 3132 8652 3732
tri 8652 3132 9252 3732 sw
tri 9500 3132 10100 3732 ne
rect 7500 2884 9252 3132
tri 9252 2884 9500 3132 sw
rect -9500 -2112 -7500 -2000
rect -9500 -3888 -9388 -2112
rect -7612 -3888 -7500 -2112
tri -10100 -4494 -9500 -3894 sw
rect -9500 -4000 -7500 -3888
tri -9145 -4494 -8651 -4000 ne
rect -8651 -4494 -7500 -4000
rect -12100 -4722 -9500 -4494
tri -12100 -4971 -11851 -4722 ne
rect -11851 -4796 -9500 -4722
tri -9500 -4796 -9198 -4494 sw
tri -8651 -4796 -8349 -4494 ne
rect -8349 -4796 -7500 -4494
rect -11851 -4971 -9198 -4796
tri -12700 -5571 -12100 -4971 sw
tri -11851 -5571 -11251 -4971 ne
rect -11251 -5571 -9198 -4971
rect -14700 -5645 -12100 -5571
tri -12100 -5645 -12026 -5571 sw
tri -11251 -5645 -11177 -5571 ne
rect -11177 -5645 -9198 -5571
tri -9198 -5645 -8349 -4796 sw
tri -8349 -5645 -7500 -4796 ne
tri -7500 -5645 -4672 -2817 sw
tri 6345 -3972 7500 -2817 se
rect 7500 -3645 9500 2884
rect 7500 -3894 9251 -3645
tri 9251 -3894 9500 -3645 nw
rect 7500 -3972 9173 -3894
tri 9173 -3972 9251 -3894 nw
tri 10022 -3972 10100 -3894 se
rect 10100 -3972 12100 3732
tri 4672 -5645 6345 -3972 se
rect 6345 -4494 8651 -3972
tri 8651 -4494 9173 -3972 nw
tri 9500 -4494 10022 -3972 se
rect 10022 -4494 12100 -3972
rect 6345 -4796 8349 -4494
tri 8349 -4796 8651 -4494 nw
tri 9198 -4796 9500 -4494 se
rect 9500 -4722 12100 -4494
rect 9500 -4796 11851 -4722
rect 6345 -5645 7500 -4796
tri 7500 -5645 8349 -4796 nw
tri 8349 -5645 9198 -4796 se
rect 9198 -4971 11851 -4796
tri 11851 -4971 12100 -4722 nw
rect 9198 -5571 11251 -4971
tri 11251 -5571 11851 -4971 nw
tri 12100 -5571 12700 -4971 se
rect 12700 -5571 14700 4809
rect 9198 -5645 11177 -5571
tri 11177 -5645 11251 -5571 nw
tri 12026 -5645 12100 -5571 se
rect 12100 -5645 14700 -5571
rect -14700 -5799 -12026 -5645
tri -14700 -6800 -13699 -5799 ne
rect -13699 -6494 -12026 -5799
tri -12026 -6494 -11177 -5645 sw
tri -11177 -6494 -10328 -5645 ne
rect -10328 -6494 -8349 -5645
tri -8349 -6494 -7500 -5645 sw
tri -7500 -6494 -6651 -5645 ne
rect -6651 -6494 -4672 -5645
rect -13699 -6800 -11177 -6494
tri -11177 -6800 -10871 -6494 sw
tri -10328 -6800 -10022 -6494 ne
rect -10022 -6800 -7500 -6494
tri -7500 -6800 -7194 -6494 sw
tri -6651 -6800 -6345 -6494 ne
rect -6345 -6800 -4672 -6494
tri -4672 -6800 -3517 -5645 sw
tri 3517 -6800 4672 -5645 se
rect 4672 -6494 6651 -5645
tri 6651 -6494 7500 -5645 nw
tri 7500 -6494 8349 -5645 se
rect 8349 -6494 10328 -5645
tri 10328 -6494 11177 -5645 nw
tri 11177 -6494 12026 -5645 se
rect 12026 -5799 14700 -5645
rect 12026 -6494 12928 -5799
rect 4672 -6800 6345 -6494
tri 6345 -6800 6651 -6494 nw
tri 7194 -6800 7500 -6494 se
rect 7500 -6722 10100 -6494
tri 10100 -6722 10328 -6494 nw
tri 10949 -6722 11177 -6494 se
rect 11177 -6722 12928 -6494
rect 7500 -6800 9251 -6722
tri -13699 -9400 -11099 -6800 ne
rect -11099 -7649 -10871 -6800
tri -10871 -7649 -10022 -6800 sw
tri -10022 -7649 -9173 -6800 ne
rect -9173 -7649 -7194 -6800
tri -7194 -7649 -6345 -6800 sw
tri -6345 -7649 -5496 -6800 ne
rect -5496 -7649 5496 -6800
tri 5496 -7649 6345 -6800 nw
tri 6345 -7649 7194 -6800 se
rect 7194 -7571 9251 -6800
tri 9251 -7571 10100 -6722 nw
tri 10100 -7571 10949 -6722 se
rect 10949 -7571 12928 -6722
tri 12928 -7571 14700 -5799 nw
rect 7194 -7649 9173 -7571
tri 9173 -7649 9251 -7571 nw
tri 10022 -7649 10100 -7571 se
rect 10100 -7649 12700 -7571
rect -11099 -8498 -10022 -7649
tri -10022 -8498 -9173 -7649 sw
tri -9173 -8498 -8324 -7649 ne
rect -8324 -7951 -6345 -7649
tri -6345 -7951 -6043 -7649 sw
tri -5496 -7951 -5194 -7649 ne
rect -5194 -7951 5194 -7649
tri 5194 -7951 5496 -7649 nw
tri 6043 -7951 6345 -7649 se
rect 6345 -7951 8349 -7649
rect -8324 -8498 -6043 -7951
rect -11099 -8551 -9173 -8498
tri -9173 -8551 -9120 -8498 sw
tri -8324 -8551 -8271 -8498 ne
rect -8271 -8551 -6043 -8498
rect -11099 -9400 -9120 -8551
tri -9120 -9400 -8271 -8551 sw
tri -8271 -9400 -7422 -8551 ne
rect -7422 -8800 -6043 -8551
tri -6043 -8800 -5194 -7951 sw
tri -5194 -8800 -4345 -7951 ne
rect -4345 -8800 4345 -7951
tri 4345 -8800 5194 -7951 nw
tri 5194 -8800 6043 -7951 se
rect 6043 -8473 8349 -7951
tri 8349 -8473 9173 -7649 nw
tri 9198 -8473 10022 -7649 se
rect 10022 -7799 12700 -7649
tri 12700 -7799 12928 -7571 nw
rect 10022 -8473 10328 -7799
rect 6043 -8800 7500 -8473
rect -7422 -9400 -5194 -8800
tri -5194 -9400 -4594 -8800 sw
tri 4594 -9400 5194 -8800 se
rect 5194 -9322 7500 -8800
tri 7500 -9322 8349 -8473 nw
tri 8349 -9322 9198 -8473 se
rect 9198 -9322 10328 -8473
rect 5194 -9400 7422 -9322
tri 7422 -9400 7500 -9322 nw
tri 8271 -9400 8349 -9322 se
rect 8349 -9400 10328 -9322
tri -11099 -12000 -8499 -9400 ne
rect -8499 -10249 -8271 -9400
tri -8271 -10249 -7422 -9400 sw
tri -7422 -10249 -6573 -9400 ne
rect -6573 -10171 6651 -9400
tri 6651 -10171 7422 -9400 nw
tri 7500 -10171 8271 -9400 se
rect 8271 -10171 10328 -9400
tri 10328 -10171 12700 -7799 nw
rect -6573 -10249 6345 -10171
rect -8499 -10551 -7422 -10249
tri -7422 -10551 -7120 -10249 sw
tri -6573 -10551 -6271 -10249 ne
rect -6271 -10477 6345 -10249
tri 6345 -10477 6651 -10171 nw
tri 7194 -10477 7500 -10171 se
rect 7500 -10399 10100 -10171
tri 10100 -10399 10328 -10171 nw
rect 7500 -10477 9173 -10399
rect -6271 -10551 5496 -10477
rect -8499 -11400 -7120 -10551
tri -7120 -11400 -6271 -10551 sw
tri -6271 -11400 -5422 -10551 ne
rect -5422 -11326 5496 -10551
tri 5496 -11326 6345 -10477 nw
tri 6345 -11326 7194 -10477 se
rect 7194 -11326 9173 -10477
tri 9173 -11326 10100 -10399 nw
rect -5422 -11400 5422 -11326
tri 5422 -11400 5496 -11326 nw
tri 6271 -11400 6345 -11326 se
rect 6345 -11400 8499 -11326
rect -8499 -12000 -6271 -11400
tri -6271 -12000 -5671 -11400 sw
tri 5671 -12000 6271 -11400 se
rect 6271 -12000 8499 -11400
tri 8499 -12000 9173 -11326 nw
tri -8499 -12999 -7500 -12000 ne
rect -7500 -12999 7500 -12000
tri 7500 -12999 8499 -12000 nw
tri -7500 -14000 -6499 -12999 ne
rect -6499 -14000 6499 -12999
tri 6499 -14000 7500 -12999 nw
<< end >>
