* SPICE3 file created from /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON/captuner_complete_2.ext - technology: sky130A

X0 BOT G0 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_0/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X1 BOT G0 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_0/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X2 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_0/S G0 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_0/S G0 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 BOT G1 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_1/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X5 BOT G1 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_1/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X6 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_1/S G1 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X7 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_1/S G1 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X8 BOT G2 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_2/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X9 BOT G2 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_2/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X10 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_2/S G2 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X11 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_2/S G2 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X12 BOT G3 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X13 BOT G3 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X14 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S G3 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X15 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S G3 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X16 BOT G3 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X17 BOT G3 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X18 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S G3 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X19 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S G3 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X20 BOT G4 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X21 BOT G4 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X22 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S G4 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X23 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S G4 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X24 BOT G4 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X25 BOT G4 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X26 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S G4 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X27 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S G4 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X28 TOP sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=1e+07u
X29 TOP sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_0/S sky130_fd_pr__cap_mim_m3_1 l=1e+06u w=5e+06u
X30 TOP sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S sky130_fd_pr__cap_mim_m3_1 l=8e+06u w=1e+07u
X31 TOP sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_1/S sky130_fd_pr__cap_mim_m3_1 l=1e+06u w=1e+07u
X32 TOP sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_2/S sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=1e+07u
C0 TOP sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S 4.41fF
C1 TOP sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_2/S 2.57fF
C2 BOT sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_1/S 10.32fF
C3 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4/S BOT 20.62fF
C4 BOT sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_2/S 10.36fF
C5 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_0/S BOT 10.34fF
C6 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S TOP 8.02fF
C7 BOT G4 2.52fF
C8 BOT G3 2.53fF
C9 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S BOT 20.72fF
C10 TOP SUB 3.06fF **FLOATING
C11 sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6/S SUB 2.81fF **FLOATING
C12 G4 SUB 3.15fF **FLOATING
C13 BOT SUB 17.11fF **FLOATING
C14 G3 SUB 3.15fF **FLOATING
