magic
tech sky130A
timestamp 1665333164
<< end >>
