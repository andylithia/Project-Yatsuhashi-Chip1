* NGSPICE file created from NMOS_50_0p5_25_4.ext - technology: sky130B

X0 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X1 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X2 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X3 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X4 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X5 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X6 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X7 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X8 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X9 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X10 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X11 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X12 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X13 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X14 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X15 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X16 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X17 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X18 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X19 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X20 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X21 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X22 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X23 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X24 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X25 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X26 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X27 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X28 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X29 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X30 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X31 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X32 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X33 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X34 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X35 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X36 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X37 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X38 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X39 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X40 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X41 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X42 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X43 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X44 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X45 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X46 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X47 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X48 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X49 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X50 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X51 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X52 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X53 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X54 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X55 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X56 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X57 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X58 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X59 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X60 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X61 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X62 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X63 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X64 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X65 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X66 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X67 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X68 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X69 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X70 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X71 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X72 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X73 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X74 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X75 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X76 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X77 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X78 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X79 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X80 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X81 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X82 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X83 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X84 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X85 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X86 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X87 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X88 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X89 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X90 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X91 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X92 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X93 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X94 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X95 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X96 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X97 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X98 SD1 G SD2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
X99 SD2 G SD1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=6e+07u l=500000u
C0 SD2 SD1 1109.22fF
C1 G SD2 86.14fF
C2 G SD1 86.39fF
C3 SD2 SUB 63.86fF $ **FLOATING
C4 SD1 SUB 53.65fF $ **FLOATING
C5 G SUB 66.73fF $ **FLOATING
