magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< error_s >>
rect 79 421 91 424
rect 38 420 91 421
rect 101 420 113 424
rect 151 420 163 424
rect 173 420 185 424
rect 38 412 80 420
rect 38 395 113 412
rect 114 400 125 412
rect 139 400 150 412
rect 42 378 76 395
rect 79 378 113 395
rect -25 262 25 264
rect 0 253 17 255
rect 25 253 27 262
rect 0 246 38 253
rect 71 251 80 279
rect 0 245 34 246
rect 0 229 8 245
rect 17 229 34 245
rect 0 228 34 229
rect 0 221 38 228
rect 25 212 27 221
rect 69 213 80 251
rect 107 207 119 241
rect 129 213 143 241
rect 129 207 141 213
rect 42 94 76 98
rect 42 64 46 94
rect 72 64 76 94
rect 16 55 38 61
rect 80 55 102 61
rect 144 55 148 395
rect 151 378 156 412
rect 180 378 185 412
rect 186 400 197 412
rect 400 395 442 421
rect 806 395 848 421
rect 1063 420 1075 424
rect 1085 420 1097 424
rect 1135 420 1147 424
rect 1157 421 1169 424
rect 1327 421 1339 424
rect 1157 420 1210 421
rect 1168 412 1210 420
rect 1051 400 1062 412
rect 332 341 336 395
rect 400 387 438 395
rect 400 380 408 387
rect 434 380 438 387
rect 810 387 844 395
rect 810 380 814 387
rect 840 380 844 387
rect 388 379 454 380
rect 794 379 860 380
rect 400 371 404 379
rect 454 365 504 367
rect 744 365 794 367
rect 494 361 548 365
rect 700 361 754 365
rect 494 356 514 361
rect 734 356 754 361
rect 504 341 506 356
rect 332 261 336 329
rect 400 305 404 341
rect 498 331 506 341
rect 514 331 515 351
rect 504 315 506 331
rect 525 322 528 356
rect 547 331 548 351
rect 557 331 564 341
rect 684 331 691 341
rect 700 331 701 351
rect 720 322 723 356
rect 733 331 734 351
rect 743 331 750 341
rect 514 315 530 321
rect 532 315 548 321
rect 700 315 716 321
rect 718 315 734 321
rect 794 315 796 365
rect 337 267 373 295
rect 337 261 351 267
rect 174 183 181 207
rect 332 183 336 251
rect 341 233 351 261
rect 361 233 375 267
rect 400 261 411 305
rect 837 267 848 305
rect 875 267 911 295
rect 562 262 612 264
rect 636 262 686 264
rect 400 233 409 261
rect 463 253 497 255
rect 442 246 497 253
rect 463 245 497 246
rect 565 253 596 255
rect 565 245 599 253
rect 400 213 404 233
rect 596 229 599 245
rect 463 228 497 229
rect 442 221 497 228
rect 565 221 599 229
rect 612 212 614 262
rect 652 253 683 255
rect 686 253 688 262
rect 875 261 887 267
rect 652 245 688 253
rect 751 253 785 255
rect 751 246 806 253
rect 751 245 785 246
rect 683 229 688 245
rect 877 233 887 261
rect 897 233 911 267
rect 652 221 688 229
rect 751 228 785 229
rect 751 221 806 228
rect 686 212 688 221
rect 332 103 336 171
rect 400 133 404 183
rect 454 159 504 161
rect 744 159 794 161
rect 504 143 506 159
rect 514 153 530 159
rect 532 153 548 159
rect 700 153 716 159
rect 718 153 734 159
rect 525 143 548 152
rect 700 143 723 152
rect 498 133 506 143
rect 504 109 506 133
rect 514 123 515 143
rect 525 118 528 143
rect 547 123 548 143
rect 557 133 564 143
rect 684 133 691 143
rect 700 123 701 143
rect 720 118 723 143
rect 733 123 734 143
rect 743 133 750 143
rect 514 109 548 113
rect 700 109 734 113
rect 794 109 796 159
rect 400 103 442 104
rect 806 103 848 104
rect 400 96 404 103
rect 295 62 300 96
rect 324 62 329 96
rect 367 62 438 96
rect 810 62 844 96
rect 847 62 881 96
rect 400 61 404 62
rect 378 55 404 61
rect 442 55 464 61
rect 784 55 806 61
rect 848 55 870 61
rect 912 55 916 395
rect 1063 378 1068 412
rect 1092 378 1097 412
rect 1098 400 1109 412
rect 1123 400 1134 412
rect 1135 395 1210 412
rect 1286 420 1339 421
rect 1349 420 1361 424
rect 1399 420 1411 424
rect 1421 420 1433 424
rect 1286 412 1328 420
rect 1286 395 1361 412
rect 1362 400 1373 412
rect 1387 400 1398 412
rect 1100 341 1104 395
rect 1135 378 1206 395
rect 1290 378 1324 395
rect 1327 378 1361 395
rect 1168 371 1172 378
rect 1100 261 1104 329
rect 1168 291 1172 341
rect 1168 251 1177 279
rect 1264 264 1274 291
rect 1223 262 1274 264
rect 1264 261 1275 262
rect 1231 253 1265 255
rect 1273 253 1275 261
rect 1100 183 1104 251
rect 1109 207 1119 241
rect 1129 207 1143 241
rect 1168 207 1179 251
rect 1210 246 1286 253
rect 1319 251 1328 279
rect 1231 228 1265 246
rect 1273 228 1275 246
rect 1210 221 1286 228
rect 1273 213 1275 221
rect 1317 213 1328 251
rect 1264 212 1275 213
rect 1109 183 1116 207
rect 1264 183 1274 212
rect 1355 207 1367 241
rect 1377 213 1391 241
rect 1377 207 1389 213
rect 1100 103 1104 171
rect 1168 133 1172 183
rect 1168 98 1172 103
rect 919 62 924 96
rect 948 62 953 96
rect 1168 94 1206 98
rect 1168 64 1176 94
rect 1202 64 1206 94
rect 1290 94 1324 98
rect 1290 64 1294 94
rect 1320 64 1324 94
rect 1168 61 1172 64
rect 1146 55 1172 61
rect 1210 55 1232 61
rect 1264 55 1286 61
rect 1328 55 1350 61
rect 1392 55 1396 395
rect 1399 378 1404 412
rect 1428 378 1433 412
rect 1434 400 1445 412
rect 1648 395 1690 421
rect 2054 395 2096 421
rect 2311 420 2323 424
rect 2333 420 2345 424
rect 2383 420 2395 424
rect 2405 421 2417 424
rect 2575 421 2587 424
rect 2405 420 2458 421
rect 2416 412 2458 420
rect 2299 400 2310 412
rect 1580 341 1584 395
rect 1648 387 1686 395
rect 1648 380 1656 387
rect 1682 380 1686 387
rect 2058 387 2092 395
rect 2058 380 2062 387
rect 2088 380 2092 387
rect 1636 379 1702 380
rect 2042 379 2108 380
rect 1648 371 1652 379
rect 1702 365 1752 367
rect 1992 365 2042 367
rect 1742 361 1796 365
rect 1948 361 2002 365
rect 1742 356 1762 361
rect 1982 356 2002 361
rect 1752 341 1754 356
rect 1580 261 1584 329
rect 1648 305 1652 341
rect 1746 331 1754 341
rect 1762 331 1763 351
rect 1752 315 1754 331
rect 1773 322 1776 356
rect 1795 331 1796 351
rect 1805 331 1812 341
rect 1932 331 1939 341
rect 1948 331 1949 351
rect 1968 322 1971 356
rect 1981 331 1982 351
rect 1991 331 1998 341
rect 1762 315 1778 321
rect 1780 315 1796 321
rect 1948 315 1964 321
rect 1966 315 1982 321
rect 2042 315 2044 365
rect 1585 267 1621 295
rect 1585 261 1599 267
rect 1422 183 1429 207
rect 1580 183 1584 251
rect 1589 233 1599 261
rect 1609 233 1623 267
rect 1648 261 1659 305
rect 2085 267 2096 305
rect 2123 267 2159 295
rect 1810 262 1860 264
rect 1884 262 1934 264
rect 1648 233 1657 261
rect 1711 253 1745 255
rect 1690 246 1745 253
rect 1711 245 1745 246
rect 1813 253 1844 255
rect 1813 245 1847 253
rect 1648 213 1652 233
rect 1844 229 1847 245
rect 1711 228 1745 229
rect 1690 221 1745 228
rect 1813 221 1847 229
rect 1860 212 1862 262
rect 1900 253 1931 255
rect 1934 253 1936 262
rect 2123 261 2135 267
rect 1900 245 1936 253
rect 1999 253 2033 255
rect 1999 246 2054 253
rect 1999 245 2033 246
rect 1931 229 1936 245
rect 2125 233 2135 261
rect 2145 233 2159 267
rect 1900 221 1936 229
rect 1999 228 2033 229
rect 1999 221 2054 228
rect 1934 212 1936 221
rect 1580 103 1584 171
rect 1648 133 1652 183
rect 1702 159 1752 161
rect 1992 159 2042 161
rect 1752 143 1754 159
rect 1762 153 1778 159
rect 1780 153 1796 159
rect 1948 153 1964 159
rect 1966 153 1982 159
rect 1773 143 1796 152
rect 1948 143 1971 152
rect 1746 133 1754 143
rect 1752 109 1754 133
rect 1762 123 1763 143
rect 1773 118 1776 143
rect 1795 123 1796 143
rect 1805 133 1812 143
rect 1932 133 1939 143
rect 1948 123 1949 143
rect 1968 118 1971 143
rect 1981 123 1982 143
rect 1991 133 1998 143
rect 1762 109 1796 113
rect 1948 109 1982 113
rect 2042 109 2044 159
rect 1648 103 1690 104
rect 2054 103 2096 104
rect 1648 96 1652 103
rect 1543 62 1548 96
rect 1572 62 1577 96
rect 1615 62 1686 96
rect 2058 62 2092 96
rect 2095 62 2129 96
rect 1648 61 1652 62
rect 1626 55 1652 61
rect 1690 55 1712 61
rect 2032 55 2054 61
rect 2096 55 2118 61
rect 2160 55 2164 395
rect 2311 378 2316 412
rect 2340 378 2345 412
rect 2346 400 2357 412
rect 2371 400 2382 412
rect 2383 395 2458 412
rect 2534 420 2587 421
rect 2597 420 2609 424
rect 2647 420 2659 424
rect 2669 420 2681 424
rect 2534 412 2576 420
rect 2534 395 2609 412
rect 2610 400 2621 412
rect 2635 400 2646 412
rect 2348 341 2352 395
rect 2383 378 2454 395
rect 2538 378 2572 395
rect 2575 378 2609 395
rect 2416 371 2420 378
rect 2348 261 2352 329
rect 2416 291 2420 341
rect 2416 251 2425 279
rect 2512 264 2522 291
rect 2471 262 2522 264
rect 2512 261 2523 262
rect 2479 253 2513 255
rect 2521 253 2523 261
rect 2348 183 2352 251
rect 2357 207 2367 241
rect 2377 207 2391 241
rect 2416 207 2427 251
rect 2458 246 2534 253
rect 2567 251 2576 279
rect 2479 228 2513 246
rect 2521 228 2523 246
rect 2458 221 2534 228
rect 2521 213 2523 221
rect 2565 213 2576 251
rect 2512 212 2523 213
rect 2357 183 2364 207
rect 2512 183 2522 212
rect 2603 207 2615 241
rect 2625 213 2639 241
rect 2625 207 2637 213
rect 2348 103 2352 171
rect 2416 133 2420 183
rect 2416 98 2420 103
rect 2167 62 2172 96
rect 2196 62 2201 96
rect 2416 94 2454 98
rect 2416 64 2424 94
rect 2450 64 2454 94
rect 2538 94 2572 98
rect 2538 64 2542 94
rect 2568 64 2572 94
rect 2416 61 2420 64
rect 2394 55 2420 61
rect 2458 55 2480 61
rect 2512 55 2534 61
rect 2576 55 2598 61
rect 2640 55 2644 395
rect 2647 378 2652 412
rect 2676 378 2681 412
rect 2682 400 2693 412
rect 2896 395 2938 421
rect 3302 395 3344 421
rect 3559 420 3571 424
rect 3581 420 3593 424
rect 3631 420 3643 424
rect 3653 421 3665 424
rect 3823 421 3835 424
rect 3653 420 3706 421
rect 3664 412 3706 420
rect 3547 400 3558 412
rect 2828 341 2832 395
rect 2896 387 2934 395
rect 2896 380 2904 387
rect 2930 380 2934 387
rect 3306 387 3340 395
rect 3306 380 3310 387
rect 3336 380 3340 387
rect 2884 379 2950 380
rect 3290 379 3356 380
rect 2896 371 2900 379
rect 2950 365 3000 367
rect 3240 365 3290 367
rect 2990 361 3044 365
rect 3196 361 3250 365
rect 2990 356 3010 361
rect 3230 356 3250 361
rect 3000 341 3002 356
rect 2828 261 2832 329
rect 2896 305 2900 341
rect 2994 331 3002 341
rect 3010 331 3011 351
rect 3000 315 3002 331
rect 3021 322 3024 356
rect 3043 331 3044 351
rect 3053 331 3060 341
rect 3180 331 3187 341
rect 3196 331 3197 351
rect 3216 322 3219 356
rect 3229 331 3230 351
rect 3239 331 3246 341
rect 3010 315 3026 321
rect 3028 315 3044 321
rect 3196 315 3212 321
rect 3214 315 3230 321
rect 3290 315 3292 365
rect 2833 267 2869 295
rect 2833 261 2847 267
rect 2670 183 2677 207
rect 2828 183 2832 251
rect 2837 233 2847 261
rect 2857 233 2871 267
rect 2896 261 2907 305
rect 3333 267 3344 305
rect 3371 267 3407 295
rect 3058 262 3108 264
rect 3132 262 3182 264
rect 2896 233 2905 261
rect 2959 253 2993 255
rect 2938 246 2993 253
rect 2959 245 2993 246
rect 3061 253 3092 255
rect 3061 245 3095 253
rect 2896 213 2900 233
rect 3092 229 3095 245
rect 2959 228 2993 229
rect 2938 221 2993 228
rect 3061 221 3095 229
rect 3108 212 3110 262
rect 3148 253 3179 255
rect 3182 253 3184 262
rect 3371 261 3383 267
rect 3148 245 3184 253
rect 3247 253 3281 255
rect 3247 246 3302 253
rect 3247 245 3281 246
rect 3179 229 3184 245
rect 3373 233 3383 261
rect 3393 233 3407 267
rect 3148 221 3184 229
rect 3247 228 3281 229
rect 3247 221 3302 228
rect 3182 212 3184 221
rect 2828 103 2832 171
rect 2896 133 2900 183
rect 2950 159 3000 161
rect 3240 159 3290 161
rect 3000 143 3002 159
rect 3010 153 3026 159
rect 3028 153 3044 159
rect 3196 153 3212 159
rect 3214 153 3230 159
rect 3021 143 3044 152
rect 3196 143 3219 152
rect 2994 133 3002 143
rect 3000 109 3002 133
rect 3010 123 3011 143
rect 3021 118 3024 143
rect 3043 123 3044 143
rect 3053 133 3060 143
rect 3180 133 3187 143
rect 3196 123 3197 143
rect 3216 118 3219 143
rect 3229 123 3230 143
rect 3239 133 3246 143
rect 3010 109 3044 113
rect 3196 109 3230 113
rect 3290 109 3292 159
rect 2896 103 2938 104
rect 3302 103 3344 104
rect 2896 96 2900 103
rect 2791 62 2796 96
rect 2820 62 2825 96
rect 2863 62 2934 96
rect 3306 62 3340 96
rect 3343 62 3377 96
rect 2896 61 2900 62
rect 2874 55 2900 61
rect 2938 55 2960 61
rect 3280 55 3302 61
rect 3344 55 3366 61
rect 3408 55 3412 395
rect 3559 378 3564 412
rect 3588 378 3593 412
rect 3594 400 3605 412
rect 3619 400 3630 412
rect 3631 395 3706 412
rect 3782 420 3835 421
rect 3845 420 3857 424
rect 3895 420 3907 424
rect 3917 420 3929 424
rect 3782 412 3824 420
rect 3782 395 3857 412
rect 3858 400 3869 412
rect 3883 400 3894 412
rect 3596 341 3600 395
rect 3631 378 3702 395
rect 3786 378 3820 395
rect 3823 378 3857 395
rect 3664 371 3668 378
rect 3596 261 3600 329
rect 3664 291 3668 341
rect 3664 251 3673 279
rect 3760 264 3770 291
rect 3719 262 3770 264
rect 3760 261 3771 262
rect 3727 253 3761 255
rect 3769 253 3771 261
rect 3596 183 3600 251
rect 3605 207 3615 241
rect 3625 207 3639 241
rect 3664 207 3675 251
rect 3706 246 3782 253
rect 3815 251 3824 279
rect 3727 228 3761 246
rect 3769 228 3771 246
rect 3706 221 3782 228
rect 3769 213 3771 221
rect 3813 213 3824 251
rect 3760 212 3771 213
rect 3605 183 3612 207
rect 3760 183 3770 212
rect 3851 207 3863 241
rect 3873 213 3887 241
rect 3873 207 3885 213
rect 3596 103 3600 171
rect 3664 133 3668 183
rect 3664 98 3668 103
rect 3415 62 3420 96
rect 3444 62 3449 96
rect 3664 94 3702 98
rect 3664 64 3672 94
rect 3698 64 3702 94
rect 3786 94 3820 98
rect 3786 64 3790 94
rect 3816 64 3820 94
rect 3664 61 3668 64
rect 3642 55 3668 61
rect 3706 55 3728 61
rect 3760 55 3782 61
rect 3824 55 3846 61
rect 3888 55 3892 395
rect 3895 378 3900 412
rect 3924 378 3929 412
rect 3930 400 3941 412
rect 4144 395 4186 421
rect 4550 395 4592 421
rect 4807 420 4819 424
rect 4829 420 4841 424
rect 4879 420 4891 424
rect 4901 421 4913 424
rect 5071 421 5083 424
rect 4901 420 4954 421
rect 4912 412 4954 420
rect 4795 400 4806 412
rect 4076 341 4080 395
rect 4144 387 4182 395
rect 4144 380 4152 387
rect 4178 380 4182 387
rect 4554 387 4588 395
rect 4554 380 4558 387
rect 4584 380 4588 387
rect 4132 379 4198 380
rect 4538 379 4604 380
rect 4144 371 4148 379
rect 4198 365 4248 367
rect 4488 365 4538 367
rect 4238 361 4292 365
rect 4444 361 4498 365
rect 4238 356 4258 361
rect 4478 356 4498 361
rect 4248 341 4250 356
rect 4076 261 4080 329
rect 4144 305 4148 341
rect 4242 331 4250 341
rect 4258 331 4259 351
rect 4248 315 4250 331
rect 4269 322 4272 356
rect 4291 331 4292 351
rect 4301 331 4308 341
rect 4428 331 4435 341
rect 4444 331 4445 351
rect 4464 322 4467 356
rect 4477 331 4478 351
rect 4487 331 4494 341
rect 4258 315 4274 321
rect 4276 315 4292 321
rect 4444 315 4460 321
rect 4462 315 4478 321
rect 4538 315 4540 365
rect 4081 267 4117 295
rect 4081 261 4095 267
rect 3918 183 3925 207
rect 4076 183 4080 251
rect 4085 233 4095 261
rect 4105 233 4119 267
rect 4144 261 4155 305
rect 4581 267 4592 305
rect 4619 267 4655 295
rect 4306 262 4356 264
rect 4380 262 4430 264
rect 4144 233 4153 261
rect 4207 253 4241 255
rect 4186 246 4241 253
rect 4207 245 4241 246
rect 4309 253 4340 255
rect 4309 245 4343 253
rect 4144 213 4148 233
rect 4340 229 4343 245
rect 4207 228 4241 229
rect 4186 221 4241 228
rect 4309 221 4343 229
rect 4356 212 4358 262
rect 4396 253 4427 255
rect 4430 253 4432 262
rect 4619 261 4631 267
rect 4396 245 4432 253
rect 4495 253 4529 255
rect 4495 246 4550 253
rect 4495 245 4529 246
rect 4427 229 4432 245
rect 4621 233 4631 261
rect 4641 233 4655 267
rect 4396 221 4432 229
rect 4495 228 4529 229
rect 4495 221 4550 228
rect 4430 212 4432 221
rect 4076 103 4080 171
rect 4144 133 4148 183
rect 4198 159 4248 161
rect 4488 159 4538 161
rect 4248 143 4250 159
rect 4258 153 4274 159
rect 4276 153 4292 159
rect 4444 153 4460 159
rect 4462 153 4478 159
rect 4269 143 4292 152
rect 4444 143 4467 152
rect 4242 133 4250 143
rect 4248 109 4250 133
rect 4258 123 4259 143
rect 4269 118 4272 143
rect 4291 123 4292 143
rect 4301 133 4308 143
rect 4428 133 4435 143
rect 4444 123 4445 143
rect 4464 118 4467 143
rect 4477 123 4478 143
rect 4487 133 4494 143
rect 4258 109 4292 113
rect 4444 109 4478 113
rect 4538 109 4540 159
rect 4144 103 4186 104
rect 4550 103 4592 104
rect 4144 96 4148 103
rect 4039 62 4044 96
rect 4068 62 4073 96
rect 4111 62 4182 96
rect 4554 62 4588 96
rect 4591 62 4625 96
rect 4144 61 4148 62
rect 4122 55 4148 61
rect 4186 55 4208 61
rect 4528 55 4550 61
rect 4592 55 4614 61
rect 4656 55 4660 395
rect 4807 378 4812 412
rect 4836 378 4841 412
rect 4842 400 4853 412
rect 4867 400 4878 412
rect 4879 395 4954 412
rect 5030 420 5083 421
rect 5093 420 5105 424
rect 5143 420 5155 424
rect 5165 420 5177 424
rect 5030 412 5072 420
rect 5030 395 5105 412
rect 5106 400 5117 412
rect 5131 400 5142 412
rect 4844 341 4848 395
rect 4879 378 4950 395
rect 5034 378 5068 395
rect 5071 378 5105 395
rect 4912 371 4916 378
rect 4844 261 4848 329
rect 4912 291 4916 341
rect 4912 251 4921 279
rect 5008 264 5018 291
rect 4967 262 5018 264
rect 5008 261 5019 262
rect 4975 253 5009 255
rect 5017 253 5019 261
rect 4844 183 4848 251
rect 4853 207 4863 241
rect 4873 207 4887 241
rect 4912 207 4923 251
rect 4954 246 5030 253
rect 5063 251 5072 279
rect 4975 228 5009 246
rect 5017 228 5019 246
rect 4954 221 5030 228
rect 5017 213 5019 221
rect 5061 213 5072 251
rect 5008 212 5019 213
rect 4853 183 4860 207
rect 5008 183 5018 212
rect 5099 207 5111 241
rect 5121 213 5135 241
rect 5121 207 5133 213
rect 4844 103 4848 171
rect 4912 133 4916 183
rect 4912 98 4916 103
rect 4663 62 4668 96
rect 4692 62 4697 96
rect 4912 94 4950 98
rect 4912 64 4920 94
rect 4946 64 4950 94
rect 5034 94 5068 98
rect 5034 64 5038 94
rect 5064 64 5068 94
rect 4912 61 4916 64
rect 4890 55 4916 61
rect 4954 55 4976 61
rect 5008 55 5030 61
rect 5072 55 5094 61
rect 5136 55 5140 395
rect 5143 378 5148 412
rect 5172 378 5177 412
rect 5178 400 5189 412
rect 5392 395 5434 421
rect 5798 395 5840 421
rect 6055 420 6067 424
rect 6077 420 6089 424
rect 6127 420 6139 424
rect 6149 421 6161 424
rect 6319 421 6331 424
rect 6149 420 6202 421
rect 6160 412 6202 420
rect 6043 400 6054 412
rect 5324 341 5328 395
rect 5392 387 5430 395
rect 5392 380 5400 387
rect 5426 380 5430 387
rect 5802 387 5836 395
rect 5802 380 5806 387
rect 5832 380 5836 387
rect 5380 379 5446 380
rect 5786 379 5852 380
rect 5392 371 5396 379
rect 5446 365 5496 367
rect 5736 365 5786 367
rect 5486 361 5540 365
rect 5692 361 5746 365
rect 5486 356 5506 361
rect 5726 356 5746 361
rect 5496 341 5498 356
rect 5324 261 5328 329
rect 5392 305 5396 341
rect 5490 331 5498 341
rect 5506 331 5507 351
rect 5496 315 5498 331
rect 5517 322 5520 356
rect 5539 331 5540 351
rect 5549 331 5556 341
rect 5676 331 5683 341
rect 5692 331 5693 351
rect 5712 322 5715 356
rect 5725 331 5726 351
rect 5735 331 5742 341
rect 5506 315 5522 321
rect 5524 315 5540 321
rect 5692 315 5708 321
rect 5710 315 5726 321
rect 5786 315 5788 365
rect 5329 267 5365 295
rect 5329 261 5343 267
rect 5166 183 5173 207
rect 5324 183 5328 251
rect 5333 233 5343 261
rect 5353 233 5367 267
rect 5392 261 5403 305
rect 5829 267 5840 305
rect 5867 267 5903 295
rect 5554 262 5604 264
rect 5628 262 5678 264
rect 5392 233 5401 261
rect 5455 253 5489 255
rect 5434 246 5489 253
rect 5455 245 5489 246
rect 5557 253 5588 255
rect 5557 245 5591 253
rect 5392 213 5396 233
rect 5588 229 5591 245
rect 5455 228 5489 229
rect 5434 221 5489 228
rect 5557 221 5591 229
rect 5604 212 5606 262
rect 5644 253 5675 255
rect 5678 253 5680 262
rect 5867 261 5879 267
rect 5644 245 5680 253
rect 5743 253 5777 255
rect 5743 246 5798 253
rect 5743 245 5777 246
rect 5675 229 5680 245
rect 5869 233 5879 261
rect 5889 233 5903 267
rect 5644 221 5680 229
rect 5743 228 5777 229
rect 5743 221 5798 228
rect 5678 212 5680 221
rect 5324 103 5328 171
rect 5392 133 5396 183
rect 5446 159 5496 161
rect 5736 159 5786 161
rect 5496 143 5498 159
rect 5506 153 5522 159
rect 5524 153 5540 159
rect 5692 153 5708 159
rect 5710 153 5726 159
rect 5517 143 5540 152
rect 5692 143 5715 152
rect 5490 133 5498 143
rect 5496 109 5498 133
rect 5506 123 5507 143
rect 5517 118 5520 143
rect 5539 123 5540 143
rect 5549 133 5556 143
rect 5676 133 5683 143
rect 5692 123 5693 143
rect 5712 118 5715 143
rect 5725 123 5726 143
rect 5735 133 5742 143
rect 5506 109 5540 113
rect 5692 109 5726 113
rect 5786 109 5788 159
rect 5392 103 5434 104
rect 5798 103 5840 104
rect 5392 96 5396 103
rect 5287 62 5292 96
rect 5316 62 5321 96
rect 5359 62 5430 96
rect 5802 62 5836 96
rect 5839 62 5873 96
rect 5392 61 5396 62
rect 5370 55 5396 61
rect 5434 55 5456 61
rect 5776 55 5798 61
rect 5840 55 5862 61
rect 5904 55 5908 395
rect 6055 378 6060 412
rect 6084 378 6089 412
rect 6090 400 6101 412
rect 6115 400 6126 412
rect 6127 395 6202 412
rect 6278 420 6331 421
rect 6341 420 6353 424
rect 6391 420 6403 424
rect 6413 420 6425 424
rect 6278 412 6320 420
rect 6278 395 6353 412
rect 6354 400 6365 412
rect 6379 400 6390 412
rect 6092 341 6096 395
rect 6127 378 6198 395
rect 6282 378 6316 395
rect 6319 378 6353 395
rect 6160 371 6164 378
rect 6092 261 6096 329
rect 6160 291 6164 341
rect 6160 251 6169 279
rect 6256 264 6266 291
rect 6215 262 6266 264
rect 6256 261 6267 262
rect 6223 253 6257 255
rect 6265 253 6267 261
rect 6092 183 6096 251
rect 6101 207 6111 241
rect 6121 207 6135 241
rect 6160 207 6171 251
rect 6202 246 6278 253
rect 6311 251 6320 279
rect 6223 228 6257 246
rect 6265 228 6267 246
rect 6202 221 6278 228
rect 6265 213 6267 221
rect 6309 213 6320 251
rect 6256 212 6267 213
rect 6101 183 6108 207
rect 6256 183 6266 212
rect 6347 207 6359 241
rect 6369 213 6383 241
rect 6369 207 6381 213
rect 6092 103 6096 171
rect 6160 133 6164 183
rect 6160 98 6164 103
rect 5911 62 5916 96
rect 5940 62 5945 96
rect 6160 94 6198 98
rect 6160 64 6168 94
rect 6194 64 6198 94
rect 6282 94 6316 98
rect 6282 64 6286 94
rect 6312 64 6316 94
rect 6160 61 6164 64
rect 6138 55 6164 61
rect 6202 55 6224 61
rect 6256 55 6278 61
rect 6320 55 6342 61
rect 6384 55 6388 395
rect 6391 378 6396 412
rect 6420 378 6425 412
rect 6426 400 6437 412
rect 6640 395 6682 421
rect 7046 395 7088 421
rect 7303 420 7315 424
rect 7325 420 7337 424
rect 7375 420 7387 424
rect 7397 421 7409 424
rect 7567 421 7579 424
rect 7397 420 7450 421
rect 7408 412 7450 420
rect 7291 400 7302 412
rect 6572 341 6576 395
rect 6640 387 6678 395
rect 6640 380 6648 387
rect 6674 380 6678 387
rect 7050 387 7084 395
rect 7050 380 7054 387
rect 7080 380 7084 387
rect 6628 379 6694 380
rect 7034 379 7100 380
rect 6640 371 6644 379
rect 6694 365 6744 367
rect 6984 365 7034 367
rect 6734 361 6788 365
rect 6940 361 6994 365
rect 6734 356 6754 361
rect 6974 356 6994 361
rect 6744 341 6746 356
rect 6572 261 6576 329
rect 6640 305 6644 341
rect 6738 331 6746 341
rect 6754 331 6755 351
rect 6744 315 6746 331
rect 6765 322 6768 356
rect 6787 331 6788 351
rect 6797 331 6804 341
rect 6924 331 6931 341
rect 6940 331 6941 351
rect 6960 322 6963 356
rect 6973 331 6974 351
rect 6983 331 6990 341
rect 6754 315 6770 321
rect 6772 315 6788 321
rect 6940 315 6956 321
rect 6958 315 6974 321
rect 7034 315 7036 365
rect 6577 267 6613 295
rect 6577 261 6591 267
rect 6414 183 6421 207
rect 6572 183 6576 251
rect 6581 233 6591 261
rect 6601 233 6615 267
rect 6640 261 6651 305
rect 7077 267 7088 305
rect 7115 267 7151 295
rect 6802 262 6852 264
rect 6876 262 6926 264
rect 6640 233 6649 261
rect 6703 253 6737 255
rect 6682 246 6737 253
rect 6703 245 6737 246
rect 6805 253 6836 255
rect 6805 245 6839 253
rect 6640 213 6644 233
rect 6836 229 6839 245
rect 6703 228 6737 229
rect 6682 221 6737 228
rect 6805 221 6839 229
rect 6852 212 6854 262
rect 6892 253 6923 255
rect 6926 253 6928 262
rect 7115 261 7127 267
rect 6892 245 6928 253
rect 6991 253 7025 255
rect 6991 246 7046 253
rect 6991 245 7025 246
rect 6923 229 6928 245
rect 7117 233 7127 261
rect 7137 233 7151 267
rect 6892 221 6928 229
rect 6991 228 7025 229
rect 6991 221 7046 228
rect 6926 212 6928 221
rect 6572 103 6576 171
rect 6640 133 6644 183
rect 6694 159 6744 161
rect 6984 159 7034 161
rect 6744 143 6746 159
rect 6754 153 6770 159
rect 6772 153 6788 159
rect 6940 153 6956 159
rect 6958 153 6974 159
rect 6765 143 6788 152
rect 6940 143 6963 152
rect 6738 133 6746 143
rect 6744 109 6746 133
rect 6754 123 6755 143
rect 6765 118 6768 143
rect 6787 123 6788 143
rect 6797 133 6804 143
rect 6924 133 6931 143
rect 6940 123 6941 143
rect 6960 118 6963 143
rect 6973 123 6974 143
rect 6983 133 6990 143
rect 6754 109 6788 113
rect 6940 109 6974 113
rect 7034 109 7036 159
rect 6640 103 6682 104
rect 7046 103 7088 104
rect 6640 96 6644 103
rect 6535 62 6540 96
rect 6564 62 6569 96
rect 6607 62 6678 96
rect 7050 62 7084 96
rect 7087 62 7121 96
rect 6640 61 6644 62
rect 6618 55 6644 61
rect 6682 55 6704 61
rect 7024 55 7046 61
rect 7088 55 7110 61
rect 7152 55 7156 395
rect 7303 378 7308 412
rect 7332 378 7337 412
rect 7338 400 7349 412
rect 7363 400 7374 412
rect 7375 395 7450 412
rect 7526 420 7579 421
rect 7589 420 7601 424
rect 7639 420 7651 424
rect 7661 420 7673 424
rect 7526 412 7568 420
rect 7526 395 7601 412
rect 7602 400 7613 412
rect 7627 400 7638 412
rect 7340 341 7344 395
rect 7375 378 7446 395
rect 7530 378 7564 395
rect 7567 378 7601 395
rect 7408 371 7412 378
rect 7340 261 7344 329
rect 7408 291 7412 341
rect 7408 251 7417 279
rect 7504 264 7514 291
rect 7463 262 7514 264
rect 7504 261 7515 262
rect 7471 253 7505 255
rect 7513 253 7515 261
rect 7340 183 7344 251
rect 7349 207 7359 241
rect 7369 207 7383 241
rect 7408 207 7419 251
rect 7450 246 7526 253
rect 7559 251 7568 279
rect 7471 228 7505 246
rect 7513 228 7515 246
rect 7450 221 7526 228
rect 7513 213 7515 221
rect 7557 213 7568 251
rect 7504 212 7515 213
rect 7349 183 7356 207
rect 7504 183 7514 212
rect 7595 207 7607 241
rect 7617 213 7631 241
rect 7617 207 7629 213
rect 7340 103 7344 171
rect 7408 133 7412 183
rect 7408 98 7412 103
rect 7159 62 7164 96
rect 7188 62 7193 96
rect 7408 94 7446 98
rect 7408 64 7416 94
rect 7442 64 7446 94
rect 7530 94 7564 98
rect 7530 64 7534 94
rect 7560 64 7564 94
rect 7408 61 7412 64
rect 7386 55 7412 61
rect 7450 55 7472 61
rect 7504 55 7526 61
rect 7568 55 7590 61
rect 7632 55 7636 395
rect 7639 378 7644 412
rect 7668 378 7673 412
rect 7674 400 7685 412
rect 7888 395 7930 421
rect 8294 395 8336 421
rect 8551 420 8563 424
rect 8573 420 8585 424
rect 8623 420 8635 424
rect 8645 421 8657 424
rect 8815 421 8827 424
rect 8645 420 8698 421
rect 8656 412 8698 420
rect 8539 400 8550 412
rect 7820 341 7824 395
rect 7888 387 7926 395
rect 7888 380 7896 387
rect 7922 380 7926 387
rect 8298 387 8332 395
rect 8298 380 8302 387
rect 8328 380 8332 387
rect 7876 379 7942 380
rect 8282 379 8348 380
rect 7888 371 7892 379
rect 7942 365 7992 367
rect 8232 365 8282 367
rect 7982 361 8036 365
rect 8188 361 8242 365
rect 7982 356 8002 361
rect 8222 356 8242 361
rect 7992 341 7994 356
rect 7820 261 7824 329
rect 7888 305 7892 341
rect 7986 331 7994 341
rect 8002 331 8003 351
rect 7992 315 7994 331
rect 8013 322 8016 356
rect 8035 331 8036 351
rect 8045 331 8052 341
rect 8172 331 8179 341
rect 8188 331 8189 351
rect 8208 322 8211 356
rect 8221 331 8222 351
rect 8231 331 8238 341
rect 8002 315 8018 321
rect 8020 315 8036 321
rect 8188 315 8204 321
rect 8206 315 8222 321
rect 8282 315 8284 365
rect 7825 267 7861 295
rect 7825 261 7839 267
rect 7662 183 7669 207
rect 7820 183 7824 251
rect 7829 233 7839 261
rect 7849 233 7863 267
rect 7888 261 7899 305
rect 8325 267 8336 305
rect 8363 267 8399 295
rect 8050 262 8100 264
rect 8124 262 8174 264
rect 7888 233 7897 261
rect 7951 253 7985 255
rect 7930 246 7985 253
rect 7951 245 7985 246
rect 8053 253 8084 255
rect 8053 245 8087 253
rect 7888 213 7892 233
rect 8084 229 8087 245
rect 7951 228 7985 229
rect 7930 221 7985 228
rect 8053 221 8087 229
rect 8100 212 8102 262
rect 8140 253 8171 255
rect 8174 253 8176 262
rect 8363 261 8375 267
rect 8140 245 8176 253
rect 8239 253 8273 255
rect 8239 246 8294 253
rect 8239 245 8273 246
rect 8171 229 8176 245
rect 8365 233 8375 261
rect 8385 233 8399 267
rect 8140 221 8176 229
rect 8239 228 8273 229
rect 8239 221 8294 228
rect 8174 212 8176 221
rect 7820 103 7824 171
rect 7888 133 7892 183
rect 7942 159 7992 161
rect 8232 159 8282 161
rect 7992 143 7994 159
rect 8002 153 8018 159
rect 8020 153 8036 159
rect 8188 153 8204 159
rect 8206 153 8222 159
rect 8013 143 8036 152
rect 8188 143 8211 152
rect 7986 133 7994 143
rect 7992 109 7994 133
rect 8002 123 8003 143
rect 8013 118 8016 143
rect 8035 123 8036 143
rect 8045 133 8052 143
rect 8172 133 8179 143
rect 8188 123 8189 143
rect 8208 118 8211 143
rect 8221 123 8222 143
rect 8231 133 8238 143
rect 8002 109 8036 113
rect 8188 109 8222 113
rect 8282 109 8284 159
rect 7888 103 7930 104
rect 8294 103 8336 104
rect 7888 96 7892 103
rect 7783 62 7788 96
rect 7812 62 7817 96
rect 7855 62 7926 96
rect 8298 62 8332 96
rect 8335 62 8369 96
rect 7888 61 7892 62
rect 7866 55 7892 61
rect 7930 55 7952 61
rect 8272 55 8294 61
rect 8336 55 8358 61
rect 8400 55 8404 395
rect 8551 378 8556 412
rect 8580 378 8585 412
rect 8586 400 8597 412
rect 8611 400 8622 412
rect 8623 395 8698 412
rect 8774 420 8827 421
rect 8837 420 8849 424
rect 8887 420 8899 424
rect 8909 420 8921 424
rect 8774 412 8816 420
rect 8774 395 8849 412
rect 8850 400 8861 412
rect 8875 400 8886 412
rect 8588 341 8592 395
rect 8623 378 8694 395
rect 8778 378 8812 395
rect 8815 378 8849 395
rect 8656 371 8660 378
rect 8588 261 8592 329
rect 8656 291 8660 341
rect 8656 251 8665 279
rect 8752 264 8762 291
rect 8711 262 8762 264
rect 8752 261 8763 262
rect 8719 253 8753 255
rect 8761 253 8763 261
rect 8588 183 8592 251
rect 8597 207 8607 241
rect 8617 207 8631 241
rect 8656 207 8667 251
rect 8698 246 8774 253
rect 8807 251 8816 279
rect 8719 228 8753 246
rect 8761 228 8763 246
rect 8698 221 8774 228
rect 8761 213 8763 221
rect 8805 213 8816 251
rect 8752 212 8763 213
rect 8597 183 8604 207
rect 8752 183 8762 212
rect 8843 207 8855 241
rect 8865 213 8879 241
rect 8865 207 8877 213
rect 8588 103 8592 171
rect 8656 133 8660 183
rect 8656 98 8660 103
rect 8407 62 8412 96
rect 8436 62 8441 96
rect 8656 94 8694 98
rect 8656 64 8664 94
rect 8690 64 8694 94
rect 8778 94 8812 98
rect 8778 64 8782 94
rect 8808 64 8812 94
rect 8656 61 8660 64
rect 8634 55 8660 61
rect 8698 55 8720 61
rect 8752 55 8774 61
rect 8816 55 8838 61
rect 8880 55 8884 395
rect 8887 378 8892 412
rect 8916 378 8921 412
rect 8922 400 8933 412
rect 9136 395 9178 421
rect 9542 395 9584 421
rect 9799 420 9811 424
rect 9821 420 9833 424
rect 9871 420 9883 424
rect 9893 421 9905 424
rect 10063 421 10075 424
rect 9893 420 9946 421
rect 9904 412 9946 420
rect 9787 400 9798 412
rect 9068 341 9072 395
rect 9136 387 9174 395
rect 9136 380 9144 387
rect 9170 380 9174 387
rect 9546 387 9580 395
rect 9546 380 9550 387
rect 9576 380 9580 387
rect 9124 379 9190 380
rect 9530 379 9596 380
rect 9136 371 9140 379
rect 9190 365 9240 367
rect 9480 365 9530 367
rect 9230 361 9284 365
rect 9436 361 9490 365
rect 9230 356 9250 361
rect 9470 356 9490 361
rect 9240 341 9242 356
rect 9068 261 9072 329
rect 9136 305 9140 341
rect 9234 331 9242 341
rect 9250 331 9251 351
rect 9240 315 9242 331
rect 9261 322 9264 356
rect 9283 331 9284 351
rect 9293 331 9300 341
rect 9420 331 9427 341
rect 9436 331 9437 351
rect 9456 322 9459 356
rect 9469 331 9470 351
rect 9479 331 9486 341
rect 9250 315 9266 321
rect 9268 315 9284 321
rect 9436 315 9452 321
rect 9454 315 9470 321
rect 9530 315 9532 365
rect 9073 267 9109 295
rect 9073 261 9087 267
rect 8910 183 8917 207
rect 9068 183 9072 251
rect 9077 233 9087 261
rect 9097 233 9111 267
rect 9136 261 9147 305
rect 9573 267 9584 305
rect 9611 267 9647 295
rect 9298 262 9348 264
rect 9372 262 9422 264
rect 9136 233 9145 261
rect 9199 253 9233 255
rect 9178 246 9233 253
rect 9199 245 9233 246
rect 9301 253 9332 255
rect 9301 245 9335 253
rect 9136 213 9140 233
rect 9332 229 9335 245
rect 9199 228 9233 229
rect 9178 221 9233 228
rect 9301 221 9335 229
rect 9348 212 9350 262
rect 9388 253 9419 255
rect 9422 253 9424 262
rect 9611 261 9623 267
rect 9388 245 9424 253
rect 9487 253 9521 255
rect 9487 246 9542 253
rect 9487 245 9521 246
rect 9419 229 9424 245
rect 9613 233 9623 261
rect 9633 233 9647 267
rect 9388 221 9424 229
rect 9487 228 9521 229
rect 9487 221 9542 228
rect 9422 212 9424 221
rect 9068 103 9072 171
rect 9136 133 9140 183
rect 9190 159 9240 161
rect 9480 159 9530 161
rect 9240 143 9242 159
rect 9250 153 9266 159
rect 9268 153 9284 159
rect 9436 153 9452 159
rect 9454 153 9470 159
rect 9261 143 9284 152
rect 9436 143 9459 152
rect 9234 133 9242 143
rect 9240 109 9242 133
rect 9250 123 9251 143
rect 9261 118 9264 143
rect 9283 123 9284 143
rect 9293 133 9300 143
rect 9420 133 9427 143
rect 9436 123 9437 143
rect 9456 118 9459 143
rect 9469 123 9470 143
rect 9479 133 9486 143
rect 9250 109 9284 113
rect 9436 109 9470 113
rect 9530 109 9532 159
rect 9136 103 9178 104
rect 9542 103 9584 104
rect 9136 96 9140 103
rect 9031 62 9036 96
rect 9060 62 9065 96
rect 9103 62 9174 96
rect 9546 62 9580 96
rect 9583 62 9617 96
rect 9136 61 9140 62
rect 9114 55 9140 61
rect 9178 55 9200 61
rect 9520 55 9542 61
rect 9584 55 9606 61
rect 9648 55 9652 395
rect 9799 378 9804 412
rect 9828 378 9833 412
rect 9834 400 9845 412
rect 9859 400 9870 412
rect 9871 395 9946 412
rect 10022 420 10075 421
rect 10085 420 10097 424
rect 10135 420 10147 424
rect 10157 420 10169 424
rect 10022 412 10064 420
rect 10022 395 10097 412
rect 10098 400 10109 412
rect 10123 400 10134 412
rect 9836 341 9840 395
rect 9871 378 9942 395
rect 10026 378 10060 395
rect 10063 378 10097 395
rect 9904 371 9908 378
rect 9836 261 9840 329
rect 9904 291 9908 341
rect 9904 251 9913 279
rect 10000 264 10010 291
rect 9959 262 10010 264
rect 10000 261 10011 262
rect 9967 253 10001 255
rect 10009 253 10011 261
rect 9836 183 9840 251
rect 9845 207 9855 241
rect 9865 207 9879 241
rect 9904 207 9915 251
rect 9946 246 10022 253
rect 10055 251 10064 279
rect 9967 228 10001 246
rect 10009 228 10011 246
rect 9946 221 10022 228
rect 10009 213 10011 221
rect 10053 213 10064 251
rect 10000 212 10011 213
rect 9845 183 9852 207
rect 10000 183 10010 212
rect 10091 207 10103 241
rect 10113 213 10127 241
rect 10113 207 10125 213
rect 9836 103 9840 171
rect 9904 133 9908 183
rect 9904 98 9908 103
rect 9655 62 9660 96
rect 9684 62 9689 96
rect 9904 94 9942 98
rect 9904 64 9912 94
rect 9938 64 9942 94
rect 10026 94 10060 98
rect 10026 64 10030 94
rect 10056 64 10060 94
rect 9904 61 9908 64
rect 9882 55 9908 61
rect 9946 55 9968 61
rect 10000 55 10022 61
rect 10064 55 10086 61
rect 10128 55 10132 395
rect 10135 378 10140 412
rect 10164 378 10169 412
rect 10170 400 10181 412
rect 10384 395 10426 421
rect 10790 395 10832 421
rect 11047 420 11059 424
rect 11069 420 11081 424
rect 11119 420 11131 424
rect 11141 421 11153 424
rect 11311 421 11323 424
rect 11141 420 11194 421
rect 11152 412 11194 420
rect 11035 400 11046 412
rect 10316 341 10320 395
rect 10384 387 10422 395
rect 10384 380 10392 387
rect 10418 380 10422 387
rect 10794 387 10828 395
rect 10794 380 10798 387
rect 10824 380 10828 387
rect 10372 379 10438 380
rect 10778 379 10844 380
rect 10384 371 10388 379
rect 10438 365 10488 367
rect 10728 365 10778 367
rect 10478 361 10532 365
rect 10684 361 10738 365
rect 10478 356 10498 361
rect 10718 356 10738 361
rect 10488 341 10490 356
rect 10316 261 10320 329
rect 10384 305 10388 341
rect 10482 331 10490 341
rect 10498 331 10499 351
rect 10488 315 10490 331
rect 10509 322 10512 356
rect 10531 331 10532 351
rect 10541 331 10548 341
rect 10668 331 10675 341
rect 10684 331 10685 351
rect 10704 322 10707 356
rect 10717 331 10718 351
rect 10727 331 10734 341
rect 10498 315 10514 321
rect 10516 315 10532 321
rect 10684 315 10700 321
rect 10702 315 10718 321
rect 10778 315 10780 365
rect 10321 267 10357 295
rect 10321 261 10335 267
rect 10158 183 10165 207
rect 10316 183 10320 251
rect 10325 233 10335 261
rect 10345 233 10359 267
rect 10384 261 10395 305
rect 10821 267 10832 305
rect 10859 267 10895 295
rect 10546 262 10596 264
rect 10620 262 10670 264
rect 10384 233 10393 261
rect 10447 253 10481 255
rect 10426 246 10481 253
rect 10447 245 10481 246
rect 10549 253 10580 255
rect 10549 245 10583 253
rect 10384 213 10388 233
rect 10580 229 10583 245
rect 10447 228 10481 229
rect 10426 221 10481 228
rect 10549 221 10583 229
rect 10596 212 10598 262
rect 10636 253 10667 255
rect 10670 253 10672 262
rect 10859 261 10871 267
rect 10636 245 10672 253
rect 10735 253 10769 255
rect 10735 246 10790 253
rect 10735 245 10769 246
rect 10667 229 10672 245
rect 10861 233 10871 261
rect 10881 233 10895 267
rect 10636 221 10672 229
rect 10735 228 10769 229
rect 10735 221 10790 228
rect 10670 212 10672 221
rect 10316 103 10320 171
rect 10384 133 10388 183
rect 10438 159 10488 161
rect 10728 159 10778 161
rect 10488 143 10490 159
rect 10498 153 10514 159
rect 10516 153 10532 159
rect 10684 153 10700 159
rect 10702 153 10718 159
rect 10509 143 10532 152
rect 10684 143 10707 152
rect 10482 133 10490 143
rect 10488 109 10490 133
rect 10498 123 10499 143
rect 10509 118 10512 143
rect 10531 123 10532 143
rect 10541 133 10548 143
rect 10668 133 10675 143
rect 10684 123 10685 143
rect 10704 118 10707 143
rect 10717 123 10718 143
rect 10727 133 10734 143
rect 10498 109 10532 113
rect 10684 109 10718 113
rect 10778 109 10780 159
rect 10384 103 10426 104
rect 10790 103 10832 104
rect 10384 96 10388 103
rect 10279 62 10284 96
rect 10308 62 10313 96
rect 10351 62 10422 96
rect 10794 62 10828 96
rect 10831 62 10865 96
rect 10384 61 10388 62
rect 10362 55 10388 61
rect 10426 55 10448 61
rect 10768 55 10790 61
rect 10832 55 10854 61
rect 10896 55 10900 395
rect 11047 378 11052 412
rect 11076 378 11081 412
rect 11082 400 11093 412
rect 11107 400 11118 412
rect 11119 395 11194 412
rect 11270 420 11323 421
rect 11333 420 11345 424
rect 11383 420 11395 424
rect 11405 420 11417 424
rect 11270 412 11312 420
rect 11270 395 11345 412
rect 11346 400 11357 412
rect 11371 400 11382 412
rect 11084 341 11088 395
rect 11119 378 11190 395
rect 11274 378 11308 395
rect 11311 378 11345 395
rect 11152 371 11156 378
rect 11084 261 11088 329
rect 11152 291 11156 341
rect 11152 251 11161 279
rect 11248 264 11258 291
rect 11207 262 11258 264
rect 11248 261 11259 262
rect 11215 253 11249 255
rect 11257 253 11259 261
rect 11084 183 11088 251
rect 11093 207 11103 241
rect 11113 207 11127 241
rect 11152 207 11163 251
rect 11194 246 11270 253
rect 11303 251 11312 279
rect 11215 228 11249 246
rect 11257 228 11259 246
rect 11194 221 11270 228
rect 11257 213 11259 221
rect 11301 213 11312 251
rect 11248 212 11259 213
rect 11093 183 11100 207
rect 11248 183 11258 212
rect 11339 207 11351 241
rect 11361 213 11375 241
rect 11361 207 11373 213
rect 11084 103 11088 171
rect 11152 133 11156 183
rect 11152 98 11156 103
rect 10903 62 10908 96
rect 10932 62 10937 96
rect 11152 94 11190 98
rect 11152 64 11160 94
rect 11186 64 11190 94
rect 11274 94 11308 98
rect 11274 64 11278 94
rect 11304 64 11308 94
rect 11152 61 11156 64
rect 11130 55 11156 61
rect 11194 55 11216 61
rect 11248 55 11270 61
rect 11312 55 11334 61
rect 11376 55 11380 395
rect 11383 378 11388 412
rect 11412 378 11417 412
rect 11418 400 11429 412
rect 11632 395 11674 421
rect 12038 395 12080 421
rect 12295 420 12307 424
rect 12317 420 12329 424
rect 12367 420 12379 424
rect 12389 421 12401 424
rect 12559 421 12571 424
rect 12389 420 12442 421
rect 12400 412 12442 420
rect 12283 400 12294 412
rect 11564 341 11568 395
rect 11632 387 11670 395
rect 11632 380 11640 387
rect 11666 380 11670 387
rect 12042 387 12076 395
rect 12042 380 12046 387
rect 12072 380 12076 387
rect 11620 379 11686 380
rect 12026 379 12092 380
rect 11632 371 11636 379
rect 11686 365 11736 367
rect 11976 365 12026 367
rect 11726 361 11780 365
rect 11932 361 11986 365
rect 11726 356 11746 361
rect 11966 356 11986 361
rect 11736 341 11738 356
rect 11564 261 11568 329
rect 11632 305 11636 341
rect 11730 331 11738 341
rect 11746 331 11747 351
rect 11736 315 11738 331
rect 11757 322 11760 356
rect 11779 331 11780 351
rect 11789 331 11796 341
rect 11916 331 11923 341
rect 11932 331 11933 351
rect 11952 322 11955 356
rect 11965 331 11966 351
rect 11975 331 11982 341
rect 11746 315 11762 321
rect 11764 315 11780 321
rect 11932 315 11948 321
rect 11950 315 11966 321
rect 12026 315 12028 365
rect 11569 267 11605 295
rect 11569 261 11583 267
rect 11406 183 11413 207
rect 11564 183 11568 251
rect 11573 233 11583 261
rect 11593 233 11607 267
rect 11632 261 11643 305
rect 12069 267 12080 305
rect 12107 267 12143 295
rect 11794 262 11844 264
rect 11868 262 11918 264
rect 11632 233 11641 261
rect 11695 253 11729 255
rect 11674 246 11729 253
rect 11695 245 11729 246
rect 11797 253 11828 255
rect 11797 245 11831 253
rect 11632 213 11636 233
rect 11828 229 11831 245
rect 11695 228 11729 229
rect 11674 221 11729 228
rect 11797 221 11831 229
rect 11844 212 11846 262
rect 11884 253 11915 255
rect 11918 253 11920 262
rect 12107 261 12119 267
rect 11884 245 11920 253
rect 11983 253 12017 255
rect 11983 246 12038 253
rect 11983 245 12017 246
rect 11915 229 11920 245
rect 12109 233 12119 261
rect 12129 233 12143 267
rect 11884 221 11920 229
rect 11983 228 12017 229
rect 11983 221 12038 228
rect 11918 212 11920 221
rect 11564 103 11568 171
rect 11632 133 11636 183
rect 11686 159 11736 161
rect 11976 159 12026 161
rect 11736 143 11738 159
rect 11746 153 11762 159
rect 11764 153 11780 159
rect 11932 153 11948 159
rect 11950 153 11966 159
rect 11757 143 11780 152
rect 11932 143 11955 152
rect 11730 133 11738 143
rect 11736 109 11738 133
rect 11746 123 11747 143
rect 11757 118 11760 143
rect 11779 123 11780 143
rect 11789 133 11796 143
rect 11916 133 11923 143
rect 11932 123 11933 143
rect 11952 118 11955 143
rect 11965 123 11966 143
rect 11975 133 11982 143
rect 11746 109 11780 113
rect 11932 109 11966 113
rect 12026 109 12028 159
rect 11632 103 11674 104
rect 12038 103 12080 104
rect 11632 96 11636 103
rect 11527 62 11532 96
rect 11556 62 11561 96
rect 11599 62 11670 96
rect 12042 62 12076 96
rect 12079 62 12113 96
rect 11632 61 11636 62
rect 11610 55 11636 61
rect 11674 55 11696 61
rect 12016 55 12038 61
rect 12080 55 12102 61
rect 12144 55 12148 395
rect 12295 378 12300 412
rect 12324 378 12329 412
rect 12330 400 12341 412
rect 12355 400 12366 412
rect 12367 395 12442 412
rect 12518 420 12571 421
rect 12581 420 12593 424
rect 12631 420 12643 424
rect 12653 420 12665 424
rect 12518 412 12560 420
rect 12518 395 12593 412
rect 12594 400 12605 412
rect 12619 400 12630 412
rect 12332 341 12336 395
rect 12367 378 12438 395
rect 12522 378 12556 395
rect 12559 378 12593 395
rect 12400 371 12404 378
rect 12332 261 12336 329
rect 12400 291 12404 341
rect 12400 251 12409 279
rect 12496 264 12506 291
rect 12455 262 12506 264
rect 12496 261 12507 262
rect 12463 253 12497 255
rect 12505 253 12507 261
rect 12332 183 12336 251
rect 12341 207 12351 241
rect 12361 207 12375 241
rect 12400 207 12411 251
rect 12442 246 12518 253
rect 12551 251 12560 279
rect 12463 228 12497 246
rect 12505 228 12507 246
rect 12442 221 12518 228
rect 12505 213 12507 221
rect 12549 213 12560 251
rect 12496 212 12507 213
rect 12341 183 12348 207
rect 12496 183 12506 212
rect 12587 207 12599 241
rect 12609 213 12623 241
rect 12609 207 12621 213
rect 12332 103 12336 171
rect 12400 133 12404 183
rect 12400 98 12404 103
rect 12151 62 12156 96
rect 12180 62 12185 96
rect 12400 94 12438 98
rect 12400 64 12408 94
rect 12434 64 12438 94
rect 12522 94 12556 98
rect 12522 64 12526 94
rect 12552 64 12556 94
rect 12400 61 12404 64
rect 12378 55 12404 61
rect 12442 55 12464 61
rect 12496 55 12518 61
rect 12560 55 12582 61
rect 12624 55 12628 395
rect 12631 378 12636 412
rect 12660 378 12665 412
rect 12666 400 12677 412
rect 12880 395 12922 421
rect 13286 395 13328 421
rect 13543 420 13555 424
rect 13565 420 13577 424
rect 13615 420 13627 424
rect 13637 421 13649 424
rect 13807 421 13819 424
rect 13637 420 13690 421
rect 13648 412 13690 420
rect 13531 400 13542 412
rect 12812 341 12816 395
rect 12880 387 12918 395
rect 12880 380 12888 387
rect 12914 380 12918 387
rect 13290 387 13324 395
rect 13290 380 13294 387
rect 13320 380 13324 387
rect 12868 379 12934 380
rect 13274 379 13340 380
rect 12880 371 12884 379
rect 12934 365 12984 367
rect 13224 365 13274 367
rect 12974 361 13028 365
rect 13180 361 13234 365
rect 12974 356 12994 361
rect 13214 356 13234 361
rect 12984 341 12986 356
rect 12812 261 12816 329
rect 12880 305 12884 341
rect 12978 331 12986 341
rect 12994 331 12995 351
rect 12984 315 12986 331
rect 13005 322 13008 356
rect 13027 331 13028 351
rect 13037 331 13044 341
rect 13164 331 13171 341
rect 13180 331 13181 351
rect 13200 322 13203 356
rect 13213 331 13214 351
rect 13223 331 13230 341
rect 12994 315 13010 321
rect 13012 315 13028 321
rect 13180 315 13196 321
rect 13198 315 13214 321
rect 13274 315 13276 365
rect 12817 267 12853 295
rect 12817 261 12831 267
rect 12654 183 12661 207
rect 12812 183 12816 251
rect 12821 233 12831 261
rect 12841 233 12855 267
rect 12880 261 12891 305
rect 13317 267 13328 305
rect 13355 267 13391 295
rect 13042 262 13092 264
rect 13116 262 13166 264
rect 12880 233 12889 261
rect 12943 253 12977 255
rect 12922 246 12977 253
rect 12943 245 12977 246
rect 13045 253 13076 255
rect 13045 245 13079 253
rect 12880 213 12884 233
rect 13076 229 13079 245
rect 12943 228 12977 229
rect 12922 221 12977 228
rect 13045 221 13079 229
rect 13092 212 13094 262
rect 13132 253 13163 255
rect 13166 253 13168 262
rect 13355 261 13367 267
rect 13132 245 13168 253
rect 13231 253 13265 255
rect 13231 246 13286 253
rect 13231 245 13265 246
rect 13163 229 13168 245
rect 13357 233 13367 261
rect 13377 233 13391 267
rect 13132 221 13168 229
rect 13231 228 13265 229
rect 13231 221 13286 228
rect 13166 212 13168 221
rect 12812 103 12816 171
rect 12880 133 12884 183
rect 12934 159 12984 161
rect 13224 159 13274 161
rect 12984 143 12986 159
rect 12994 153 13010 159
rect 13012 153 13028 159
rect 13180 153 13196 159
rect 13198 153 13214 159
rect 13005 143 13028 152
rect 13180 143 13203 152
rect 12978 133 12986 143
rect 12984 109 12986 133
rect 12994 123 12995 143
rect 13005 118 13008 143
rect 13027 123 13028 143
rect 13037 133 13044 143
rect 13164 133 13171 143
rect 13180 123 13181 143
rect 13200 118 13203 143
rect 13213 123 13214 143
rect 13223 133 13230 143
rect 12994 109 13028 113
rect 13180 109 13214 113
rect 13274 109 13276 159
rect 12880 103 12922 104
rect 13286 103 13328 104
rect 12880 96 12884 103
rect 12775 62 12780 96
rect 12804 62 12809 96
rect 12847 62 12918 96
rect 13290 62 13324 96
rect 13327 62 13361 96
rect 12880 61 12884 62
rect 12858 55 12884 61
rect 12922 55 12944 61
rect 13264 55 13286 61
rect 13328 55 13350 61
rect 13392 55 13396 395
rect 13543 378 13548 412
rect 13572 378 13577 412
rect 13578 400 13589 412
rect 13603 400 13614 412
rect 13615 395 13690 412
rect 13766 420 13819 421
rect 13829 420 13841 424
rect 13879 420 13891 424
rect 13901 420 13913 424
rect 13766 412 13808 420
rect 13766 395 13841 412
rect 13842 400 13853 412
rect 13867 400 13878 412
rect 13580 341 13584 395
rect 13615 378 13686 395
rect 13770 378 13804 395
rect 13807 378 13841 395
rect 13648 371 13652 378
rect 13580 261 13584 329
rect 13648 291 13652 341
rect 13648 251 13657 279
rect 13744 264 13754 291
rect 13703 262 13754 264
rect 13744 261 13755 262
rect 13711 253 13745 255
rect 13753 253 13755 261
rect 13580 183 13584 251
rect 13589 207 13599 241
rect 13609 207 13623 241
rect 13648 207 13659 251
rect 13690 246 13766 253
rect 13799 251 13808 279
rect 13711 228 13745 246
rect 13753 228 13755 246
rect 13690 221 13766 228
rect 13753 213 13755 221
rect 13797 213 13808 251
rect 13744 212 13755 213
rect 13589 183 13596 207
rect 13744 183 13754 212
rect 13835 207 13847 241
rect 13857 213 13871 241
rect 13857 207 13869 213
rect 13580 103 13584 171
rect 13648 133 13652 183
rect 13648 98 13652 103
rect 13399 62 13404 96
rect 13428 62 13433 96
rect 13648 94 13686 98
rect 13648 64 13656 94
rect 13682 64 13686 94
rect 13770 94 13804 98
rect 13770 64 13774 94
rect 13800 64 13804 94
rect 13648 61 13652 64
rect 13626 55 13652 61
rect 13690 55 13712 61
rect 13744 55 13766 61
rect 13808 55 13830 61
rect 13872 55 13876 395
rect 13879 378 13884 412
rect 13908 378 13913 412
rect 13914 400 13925 412
rect 14128 395 14170 421
rect 14534 395 14576 421
rect 14791 420 14803 424
rect 14813 420 14825 424
rect 14863 420 14875 424
rect 14885 421 14897 424
rect 15055 421 15067 424
rect 14885 420 14938 421
rect 14896 412 14938 420
rect 14779 400 14790 412
rect 14060 341 14064 395
rect 14128 387 14166 395
rect 14128 380 14136 387
rect 14162 380 14166 387
rect 14538 387 14572 395
rect 14538 380 14542 387
rect 14568 380 14572 387
rect 14116 379 14182 380
rect 14522 379 14588 380
rect 14128 371 14132 379
rect 14182 365 14232 367
rect 14472 365 14522 367
rect 14222 361 14276 365
rect 14428 361 14482 365
rect 14222 356 14242 361
rect 14462 356 14482 361
rect 14232 341 14234 356
rect 14060 261 14064 329
rect 14128 305 14132 341
rect 14226 331 14234 341
rect 14242 331 14243 351
rect 14232 315 14234 331
rect 14253 322 14256 356
rect 14275 331 14276 351
rect 14285 331 14292 341
rect 14412 331 14419 341
rect 14428 331 14429 351
rect 14448 322 14451 356
rect 14461 331 14462 351
rect 14471 331 14478 341
rect 14242 315 14258 321
rect 14260 315 14276 321
rect 14428 315 14444 321
rect 14446 315 14462 321
rect 14522 315 14524 365
rect 14065 267 14101 295
rect 14065 261 14079 267
rect 13902 183 13909 207
rect 14060 183 14064 251
rect 14069 233 14079 261
rect 14089 233 14103 267
rect 14128 261 14139 305
rect 14565 267 14576 305
rect 14603 267 14639 295
rect 14290 262 14340 264
rect 14364 262 14414 264
rect 14128 233 14137 261
rect 14191 253 14225 255
rect 14170 246 14225 253
rect 14191 245 14225 246
rect 14293 253 14324 255
rect 14293 245 14327 253
rect 14128 213 14132 233
rect 14324 229 14327 245
rect 14191 228 14225 229
rect 14170 221 14225 228
rect 14293 221 14327 229
rect 14340 212 14342 262
rect 14380 253 14411 255
rect 14414 253 14416 262
rect 14603 261 14615 267
rect 14380 245 14416 253
rect 14479 253 14513 255
rect 14479 246 14534 253
rect 14479 245 14513 246
rect 14411 229 14416 245
rect 14605 233 14615 261
rect 14625 233 14639 267
rect 14380 221 14416 229
rect 14479 228 14513 229
rect 14479 221 14534 228
rect 14414 212 14416 221
rect 14060 103 14064 171
rect 14128 133 14132 183
rect 14182 159 14232 161
rect 14472 159 14522 161
rect 14232 143 14234 159
rect 14242 153 14258 159
rect 14260 153 14276 159
rect 14428 153 14444 159
rect 14446 153 14462 159
rect 14253 143 14276 152
rect 14428 143 14451 152
rect 14226 133 14234 143
rect 14232 109 14234 133
rect 14242 123 14243 143
rect 14253 118 14256 143
rect 14275 123 14276 143
rect 14285 133 14292 143
rect 14412 133 14419 143
rect 14428 123 14429 143
rect 14448 118 14451 143
rect 14461 123 14462 143
rect 14471 133 14478 143
rect 14242 109 14276 113
rect 14428 109 14462 113
rect 14522 109 14524 159
rect 14128 103 14170 104
rect 14534 103 14576 104
rect 14128 96 14132 103
rect 14023 62 14028 96
rect 14052 62 14057 96
rect 14095 62 14166 96
rect 14538 62 14572 96
rect 14575 62 14609 96
rect 14128 61 14132 62
rect 14106 55 14132 61
rect 14170 55 14192 61
rect 14512 55 14534 61
rect 14576 55 14598 61
rect 14640 55 14644 395
rect 14791 378 14796 412
rect 14820 378 14825 412
rect 14826 400 14837 412
rect 14851 400 14862 412
rect 14863 395 14938 412
rect 15014 420 15067 421
rect 15077 420 15089 424
rect 15127 420 15139 424
rect 15149 420 15161 424
rect 15014 412 15056 420
rect 15014 395 15089 412
rect 15090 400 15101 412
rect 15115 400 15126 412
rect 14828 341 14832 395
rect 14863 378 14934 395
rect 15018 378 15052 395
rect 15055 378 15089 395
rect 14896 371 14900 378
rect 14828 261 14832 329
rect 14896 291 14900 341
rect 14896 251 14905 279
rect 14992 264 15002 291
rect 14951 262 15002 264
rect 14992 261 15003 262
rect 14959 253 14993 255
rect 15001 253 15003 261
rect 14828 183 14832 251
rect 14837 207 14847 241
rect 14857 207 14871 241
rect 14896 207 14907 251
rect 14938 246 15014 253
rect 15047 251 15056 279
rect 14959 228 14993 246
rect 15001 228 15003 246
rect 14938 221 15014 228
rect 15001 213 15003 221
rect 15045 213 15056 251
rect 14992 212 15003 213
rect 14837 183 14844 207
rect 14992 183 15002 212
rect 15083 207 15095 241
rect 15105 213 15119 241
rect 15105 207 15117 213
rect 14828 103 14832 171
rect 14896 133 14900 183
rect 14896 98 14900 103
rect 14647 62 14652 96
rect 14676 62 14681 96
rect 14896 94 14934 98
rect 14896 64 14904 94
rect 14930 64 14934 94
rect 15018 94 15052 98
rect 15018 64 15022 94
rect 15048 64 15052 94
rect 14896 61 14900 64
rect 14874 55 14900 61
rect 14938 55 14960 61
rect 14992 55 15014 61
rect 15056 55 15078 61
rect 15120 55 15124 395
rect 15127 378 15132 412
rect 15156 378 15161 412
rect 15162 400 15173 412
rect 15376 395 15418 421
rect 15782 395 15824 421
rect 16039 420 16051 424
rect 16061 420 16073 424
rect 16111 420 16123 424
rect 16133 421 16145 424
rect 16303 421 16315 424
rect 16133 420 16186 421
rect 16144 412 16186 420
rect 16027 400 16038 412
rect 15308 341 15312 395
rect 15376 387 15414 395
rect 15376 380 15384 387
rect 15410 380 15414 387
rect 15786 387 15820 395
rect 15786 380 15790 387
rect 15816 380 15820 387
rect 15364 379 15430 380
rect 15770 379 15836 380
rect 15376 371 15380 379
rect 15430 365 15480 367
rect 15720 365 15770 367
rect 15470 361 15524 365
rect 15676 361 15730 365
rect 15470 356 15490 361
rect 15710 356 15730 361
rect 15480 341 15482 356
rect 15308 261 15312 329
rect 15376 305 15380 341
rect 15474 331 15482 341
rect 15490 331 15491 351
rect 15480 315 15482 331
rect 15501 322 15504 356
rect 15523 331 15524 351
rect 15533 331 15540 341
rect 15660 331 15667 341
rect 15676 331 15677 351
rect 15696 322 15699 356
rect 15709 331 15710 351
rect 15719 331 15726 341
rect 15490 315 15506 321
rect 15508 315 15524 321
rect 15676 315 15692 321
rect 15694 315 15710 321
rect 15770 315 15772 365
rect 15313 267 15349 295
rect 15313 261 15327 267
rect 15150 183 15157 207
rect 15308 183 15312 251
rect 15317 233 15327 261
rect 15337 233 15351 267
rect 15376 261 15387 305
rect 15813 267 15824 305
rect 15851 267 15887 295
rect 15538 262 15588 264
rect 15612 262 15662 264
rect 15376 233 15385 261
rect 15439 253 15473 255
rect 15418 246 15473 253
rect 15439 245 15473 246
rect 15541 253 15572 255
rect 15541 245 15575 253
rect 15376 213 15380 233
rect 15572 229 15575 245
rect 15439 228 15473 229
rect 15418 221 15473 228
rect 15541 221 15575 229
rect 15588 212 15590 262
rect 15628 253 15659 255
rect 15662 253 15664 262
rect 15851 261 15863 267
rect 15628 245 15664 253
rect 15727 253 15761 255
rect 15727 246 15782 253
rect 15727 245 15761 246
rect 15659 229 15664 245
rect 15853 233 15863 261
rect 15873 233 15887 267
rect 15628 221 15664 229
rect 15727 228 15761 229
rect 15727 221 15782 228
rect 15662 212 15664 221
rect 15308 103 15312 171
rect 15376 133 15380 183
rect 15430 159 15480 161
rect 15720 159 15770 161
rect 15480 143 15482 159
rect 15490 153 15506 159
rect 15508 153 15524 159
rect 15676 153 15692 159
rect 15694 153 15710 159
rect 15501 143 15524 152
rect 15676 143 15699 152
rect 15474 133 15482 143
rect 15480 109 15482 133
rect 15490 123 15491 143
rect 15501 118 15504 143
rect 15523 123 15524 143
rect 15533 133 15540 143
rect 15660 133 15667 143
rect 15676 123 15677 143
rect 15696 118 15699 143
rect 15709 123 15710 143
rect 15719 133 15726 143
rect 15490 109 15524 113
rect 15676 109 15710 113
rect 15770 109 15772 159
rect 15376 103 15418 104
rect 15782 103 15824 104
rect 15376 96 15380 103
rect 15271 62 15276 96
rect 15300 62 15305 96
rect 15343 62 15414 96
rect 15786 62 15820 96
rect 15823 62 15857 96
rect 15376 61 15380 62
rect 15354 55 15380 61
rect 15418 55 15440 61
rect 15760 55 15782 61
rect 15824 55 15846 61
rect 15888 55 15892 395
rect 16039 378 16044 412
rect 16068 378 16073 412
rect 16074 400 16085 412
rect 16099 400 16110 412
rect 16111 395 16186 412
rect 16262 420 16315 421
rect 16325 420 16337 424
rect 16375 420 16387 424
rect 16397 420 16409 424
rect 16262 412 16304 420
rect 16262 395 16337 412
rect 16338 400 16349 412
rect 16363 400 16374 412
rect 16076 341 16080 395
rect 16111 378 16182 395
rect 16266 378 16300 395
rect 16303 378 16337 395
rect 16144 371 16148 378
rect 16076 261 16080 329
rect 16144 291 16148 341
rect 16144 251 16153 279
rect 16240 264 16250 291
rect 16199 262 16250 264
rect 16240 261 16251 262
rect 16207 253 16241 255
rect 16249 253 16251 261
rect 16076 183 16080 251
rect 16085 207 16095 241
rect 16105 207 16119 241
rect 16144 207 16155 251
rect 16186 246 16262 253
rect 16295 251 16304 279
rect 16207 228 16241 246
rect 16249 228 16251 246
rect 16186 221 16262 228
rect 16249 213 16251 221
rect 16293 213 16304 251
rect 16240 212 16251 213
rect 16085 183 16092 207
rect 16240 183 16250 212
rect 16331 207 16343 241
rect 16353 213 16367 241
rect 16353 207 16365 213
rect 16076 103 16080 171
rect 16144 133 16148 183
rect 16144 98 16148 103
rect 15895 62 15900 96
rect 15924 62 15929 96
rect 16144 94 16182 98
rect 16144 64 16152 94
rect 16178 64 16182 94
rect 16266 94 16300 98
rect 16266 64 16270 94
rect 16296 64 16300 94
rect 16144 61 16148 64
rect 16122 55 16148 61
rect 16186 55 16208 61
rect 16240 55 16262 61
rect 16304 55 16326 61
rect 16368 55 16372 395
rect 16375 378 16380 412
rect 16404 378 16409 412
rect 16410 400 16421 412
rect 16624 395 16666 421
rect 17030 395 17072 421
rect 17287 420 17299 424
rect 17309 420 17321 424
rect 17359 420 17371 424
rect 17381 421 17393 424
rect 17551 421 17563 424
rect 17381 420 17434 421
rect 17392 412 17434 420
rect 17275 400 17286 412
rect 16556 341 16560 395
rect 16624 387 16662 395
rect 16624 380 16632 387
rect 16658 380 16662 387
rect 17034 387 17068 395
rect 17034 380 17038 387
rect 17064 380 17068 387
rect 16612 379 16678 380
rect 17018 379 17084 380
rect 16624 371 16628 379
rect 16678 365 16728 367
rect 16968 365 17018 367
rect 16718 361 16772 365
rect 16924 361 16978 365
rect 16718 356 16738 361
rect 16958 356 16978 361
rect 16728 341 16730 356
rect 16556 261 16560 329
rect 16624 305 16628 341
rect 16722 331 16730 341
rect 16738 331 16739 351
rect 16728 315 16730 331
rect 16749 322 16752 356
rect 16771 331 16772 351
rect 16781 331 16788 341
rect 16908 331 16915 341
rect 16924 331 16925 351
rect 16944 322 16947 356
rect 16957 331 16958 351
rect 16967 331 16974 341
rect 16738 315 16754 321
rect 16756 315 16772 321
rect 16924 315 16940 321
rect 16942 315 16958 321
rect 17018 315 17020 365
rect 16561 267 16597 295
rect 16561 261 16575 267
rect 16398 183 16405 207
rect 16556 183 16560 251
rect 16565 233 16575 261
rect 16585 233 16599 267
rect 16624 261 16635 305
rect 17061 267 17072 305
rect 17099 267 17135 295
rect 16786 262 16836 264
rect 16860 262 16910 264
rect 16624 233 16633 261
rect 16687 253 16721 255
rect 16666 246 16721 253
rect 16687 245 16721 246
rect 16789 253 16820 255
rect 16789 245 16823 253
rect 16624 213 16628 233
rect 16820 229 16823 245
rect 16687 228 16721 229
rect 16666 221 16721 228
rect 16789 221 16823 229
rect 16836 212 16838 262
rect 16876 253 16907 255
rect 16910 253 16912 262
rect 17099 261 17111 267
rect 16876 245 16912 253
rect 16975 253 17009 255
rect 16975 246 17030 253
rect 16975 245 17009 246
rect 16907 229 16912 245
rect 17101 233 17111 261
rect 17121 233 17135 267
rect 16876 221 16912 229
rect 16975 228 17009 229
rect 16975 221 17030 228
rect 16910 212 16912 221
rect 16556 103 16560 171
rect 16624 133 16628 183
rect 16678 159 16728 161
rect 16968 159 17018 161
rect 16728 143 16730 159
rect 16738 153 16754 159
rect 16756 153 16772 159
rect 16924 153 16940 159
rect 16942 153 16958 159
rect 16749 143 16772 152
rect 16924 143 16947 152
rect 16722 133 16730 143
rect 16728 109 16730 133
rect 16738 123 16739 143
rect 16749 118 16752 143
rect 16771 123 16772 143
rect 16781 133 16788 143
rect 16908 133 16915 143
rect 16924 123 16925 143
rect 16944 118 16947 143
rect 16957 123 16958 143
rect 16967 133 16974 143
rect 16738 109 16772 113
rect 16924 109 16958 113
rect 17018 109 17020 159
rect 16624 103 16666 104
rect 17030 103 17072 104
rect 16624 96 16628 103
rect 16519 62 16524 96
rect 16548 62 16553 96
rect 16591 62 16662 96
rect 17034 62 17068 96
rect 17071 62 17105 96
rect 16624 61 16628 62
rect 16602 55 16628 61
rect 16666 55 16688 61
rect 17008 55 17030 61
rect 17072 55 17094 61
rect 17136 55 17140 395
rect 17287 378 17292 412
rect 17316 378 17321 412
rect 17322 400 17333 412
rect 17347 400 17358 412
rect 17359 395 17434 412
rect 17510 420 17563 421
rect 17573 420 17585 424
rect 17623 420 17635 424
rect 17645 420 17657 424
rect 17510 412 17552 420
rect 17510 395 17585 412
rect 17586 400 17597 412
rect 17611 400 17622 412
rect 17324 341 17328 395
rect 17359 378 17430 395
rect 17514 378 17548 395
rect 17551 378 17585 395
rect 17392 371 17396 378
rect 17324 261 17328 329
rect 17392 291 17396 341
rect 17392 251 17401 279
rect 17488 264 17498 291
rect 17447 262 17498 264
rect 17488 261 17499 262
rect 17455 253 17489 255
rect 17497 253 17499 261
rect 17324 183 17328 251
rect 17333 207 17343 241
rect 17353 207 17367 241
rect 17392 207 17403 251
rect 17434 246 17510 253
rect 17543 251 17552 279
rect 17455 228 17489 246
rect 17497 228 17499 246
rect 17434 221 17510 228
rect 17497 213 17499 221
rect 17541 213 17552 251
rect 17488 212 17499 213
rect 17333 183 17340 207
rect 17488 183 17498 212
rect 17579 207 17591 241
rect 17601 213 17615 241
rect 17601 207 17613 213
rect 17324 103 17328 171
rect 17392 133 17396 183
rect 17392 98 17396 103
rect 17143 62 17148 96
rect 17172 62 17177 96
rect 17392 94 17430 98
rect 17392 64 17400 94
rect 17426 64 17430 94
rect 17514 94 17548 98
rect 17514 64 17518 94
rect 17544 64 17548 94
rect 17392 61 17396 64
rect 17370 55 17396 61
rect 17434 55 17456 61
rect 17488 55 17510 61
rect 17552 55 17574 61
rect 17616 55 17620 395
rect 17623 378 17628 412
rect 17652 378 17657 412
rect 17658 400 17669 412
rect 17872 395 17914 421
rect 18278 395 18320 421
rect 18535 420 18547 424
rect 18557 420 18569 424
rect 18607 420 18619 424
rect 18629 421 18641 424
rect 18799 421 18811 424
rect 18629 420 18682 421
rect 18640 412 18682 420
rect 18523 400 18534 412
rect 17804 341 17808 395
rect 17872 387 17910 395
rect 17872 380 17880 387
rect 17906 380 17910 387
rect 18282 387 18316 395
rect 18282 380 18286 387
rect 18312 380 18316 387
rect 17860 379 17926 380
rect 18266 379 18332 380
rect 17872 371 17876 379
rect 17926 365 17976 367
rect 18216 365 18266 367
rect 17966 361 18020 365
rect 18172 361 18226 365
rect 17966 356 17986 361
rect 18206 356 18226 361
rect 17976 341 17978 356
rect 17804 261 17808 329
rect 17872 305 17876 341
rect 17970 331 17978 341
rect 17986 331 17987 351
rect 17976 315 17978 331
rect 17997 322 18000 356
rect 18019 331 18020 351
rect 18029 331 18036 341
rect 18156 331 18163 341
rect 18172 331 18173 351
rect 18192 322 18195 356
rect 18205 331 18206 351
rect 18215 331 18222 341
rect 17986 315 18002 321
rect 18004 315 18020 321
rect 18172 315 18188 321
rect 18190 315 18206 321
rect 18266 315 18268 365
rect 17809 267 17845 295
rect 17809 261 17823 267
rect 17646 183 17653 207
rect 17804 183 17808 251
rect 17813 233 17823 261
rect 17833 233 17847 267
rect 17872 261 17883 305
rect 18309 267 18320 305
rect 18347 267 18383 295
rect 18034 262 18084 264
rect 18108 262 18158 264
rect 17872 233 17881 261
rect 17935 253 17969 255
rect 17914 246 17969 253
rect 17935 245 17969 246
rect 18037 253 18068 255
rect 18037 245 18071 253
rect 17872 213 17876 233
rect 18068 229 18071 245
rect 17935 228 17969 229
rect 17914 221 17969 228
rect 18037 221 18071 229
rect 18084 212 18086 262
rect 18124 253 18155 255
rect 18158 253 18160 262
rect 18347 261 18359 267
rect 18124 245 18160 253
rect 18223 253 18257 255
rect 18223 246 18278 253
rect 18223 245 18257 246
rect 18155 229 18160 245
rect 18349 233 18359 261
rect 18369 233 18383 267
rect 18124 221 18160 229
rect 18223 228 18257 229
rect 18223 221 18278 228
rect 18158 212 18160 221
rect 17804 103 17808 171
rect 17872 133 17876 183
rect 17926 159 17976 161
rect 18216 159 18266 161
rect 17976 143 17978 159
rect 17986 153 18002 159
rect 18004 153 18020 159
rect 18172 153 18188 159
rect 18190 153 18206 159
rect 17997 143 18020 152
rect 18172 143 18195 152
rect 17970 133 17978 143
rect 17976 109 17978 133
rect 17986 123 17987 143
rect 17997 118 18000 143
rect 18019 123 18020 143
rect 18029 133 18036 143
rect 18156 133 18163 143
rect 18172 123 18173 143
rect 18192 118 18195 143
rect 18205 123 18206 143
rect 18215 133 18222 143
rect 17986 109 18020 113
rect 18172 109 18206 113
rect 18266 109 18268 159
rect 17872 103 17914 104
rect 18278 103 18320 104
rect 17872 96 17876 103
rect 17767 62 17772 96
rect 17796 62 17801 96
rect 17839 62 17910 96
rect 18282 62 18316 96
rect 18319 62 18353 96
rect 17872 61 17876 62
rect 17850 55 17876 61
rect 17914 55 17936 61
rect 18256 55 18278 61
rect 18320 55 18342 61
rect 18384 55 18388 395
rect 18535 378 18540 412
rect 18564 378 18569 412
rect 18570 400 18581 412
rect 18595 400 18606 412
rect 18607 395 18682 412
rect 18758 420 18811 421
rect 18821 420 18833 424
rect 18871 420 18883 424
rect 18893 420 18905 424
rect 18758 412 18800 420
rect 18758 395 18833 412
rect 18834 400 18845 412
rect 18859 400 18870 412
rect 18572 341 18576 395
rect 18607 378 18678 395
rect 18762 378 18796 395
rect 18799 378 18833 395
rect 18640 371 18644 378
rect 18572 261 18576 329
rect 18640 291 18644 341
rect 18640 251 18649 279
rect 18736 264 18746 291
rect 18695 262 18746 264
rect 18736 261 18747 262
rect 18703 253 18737 255
rect 18745 253 18747 261
rect 18572 183 18576 251
rect 18581 207 18591 241
rect 18601 207 18615 241
rect 18640 207 18651 251
rect 18682 246 18758 253
rect 18791 251 18800 279
rect 18703 228 18737 246
rect 18745 228 18747 246
rect 18682 221 18758 228
rect 18745 213 18747 221
rect 18789 213 18800 251
rect 18736 212 18747 213
rect 18581 183 18588 207
rect 18736 183 18746 212
rect 18827 207 18839 241
rect 18849 213 18863 241
rect 18849 207 18861 213
rect 18572 103 18576 171
rect 18640 133 18644 183
rect 18640 98 18644 103
rect 18391 62 18396 96
rect 18420 62 18425 96
rect 18640 94 18678 98
rect 18640 64 18648 94
rect 18674 64 18678 94
rect 18762 94 18796 98
rect 18762 64 18766 94
rect 18792 64 18796 94
rect 18640 61 18644 64
rect 18618 55 18644 61
rect 18682 55 18704 61
rect 18736 55 18758 61
rect 18800 55 18822 61
rect 18864 55 18868 395
rect 18871 378 18876 412
rect 18900 378 18905 412
rect 18906 400 18917 412
rect 19120 395 19162 421
rect 19526 395 19568 421
rect 19783 420 19795 424
rect 19805 420 19817 424
rect 19855 420 19867 424
rect 19877 421 19889 424
rect 20047 421 20059 424
rect 19877 420 19930 421
rect 19888 412 19930 420
rect 19771 400 19782 412
rect 19052 341 19056 395
rect 19120 387 19158 395
rect 19120 380 19128 387
rect 19154 380 19158 387
rect 19530 387 19564 395
rect 19530 380 19534 387
rect 19560 380 19564 387
rect 19108 379 19174 380
rect 19514 379 19580 380
rect 19120 371 19124 379
rect 19174 365 19224 367
rect 19464 365 19514 367
rect 19214 361 19268 365
rect 19420 361 19474 365
rect 19214 356 19234 361
rect 19454 356 19474 361
rect 19224 341 19226 356
rect 19052 261 19056 329
rect 19120 305 19124 341
rect 19218 331 19226 341
rect 19234 331 19235 351
rect 19224 315 19226 331
rect 19245 322 19248 356
rect 19267 331 19268 351
rect 19277 331 19284 341
rect 19404 331 19411 341
rect 19420 331 19421 351
rect 19440 322 19443 356
rect 19453 331 19454 351
rect 19463 331 19470 341
rect 19234 315 19250 321
rect 19252 315 19268 321
rect 19420 315 19436 321
rect 19438 315 19454 321
rect 19514 315 19516 365
rect 19057 267 19093 295
rect 19057 261 19071 267
rect 18894 183 18901 207
rect 19052 183 19056 251
rect 19061 233 19071 261
rect 19081 233 19095 267
rect 19120 261 19131 305
rect 19557 267 19568 305
rect 19595 267 19631 295
rect 19282 262 19332 264
rect 19356 262 19406 264
rect 19120 233 19129 261
rect 19183 253 19217 255
rect 19162 246 19217 253
rect 19183 245 19217 246
rect 19285 253 19316 255
rect 19285 245 19319 253
rect 19120 213 19124 233
rect 19316 229 19319 245
rect 19183 228 19217 229
rect 19162 221 19217 228
rect 19285 221 19319 229
rect 19332 212 19334 262
rect 19372 253 19403 255
rect 19406 253 19408 262
rect 19595 261 19607 267
rect 19372 245 19408 253
rect 19471 253 19505 255
rect 19471 246 19526 253
rect 19471 245 19505 246
rect 19403 229 19408 245
rect 19597 233 19607 261
rect 19617 233 19631 267
rect 19372 221 19408 229
rect 19471 228 19505 229
rect 19471 221 19526 228
rect 19406 212 19408 221
rect 19052 103 19056 171
rect 19120 133 19124 183
rect 19174 159 19224 161
rect 19464 159 19514 161
rect 19224 143 19226 159
rect 19234 153 19250 159
rect 19252 153 19268 159
rect 19420 153 19436 159
rect 19438 153 19454 159
rect 19245 143 19268 152
rect 19420 143 19443 152
rect 19218 133 19226 143
rect 19224 109 19226 133
rect 19234 123 19235 143
rect 19245 118 19248 143
rect 19267 123 19268 143
rect 19277 133 19284 143
rect 19404 133 19411 143
rect 19420 123 19421 143
rect 19440 118 19443 143
rect 19453 123 19454 143
rect 19463 133 19470 143
rect 19234 109 19268 113
rect 19420 109 19454 113
rect 19514 109 19516 159
rect 19120 103 19162 104
rect 19526 103 19568 104
rect 19120 96 19124 103
rect 19015 62 19020 96
rect 19044 62 19049 96
rect 19087 62 19158 96
rect 19530 62 19564 96
rect 19567 62 19601 96
rect 19120 61 19124 62
rect 19098 55 19124 61
rect 19162 55 19184 61
rect 19504 55 19526 61
rect 19568 55 19590 61
rect 19632 55 19636 395
rect 19783 378 19788 412
rect 19812 378 19817 412
rect 19818 400 19829 412
rect 19843 400 19854 412
rect 19855 395 19930 412
rect 20006 420 20059 421
rect 20069 420 20081 424
rect 20119 420 20131 424
rect 20141 420 20153 424
rect 20006 412 20048 420
rect 20006 395 20081 412
rect 20082 400 20093 412
rect 20107 400 20118 412
rect 19820 341 19824 395
rect 19855 378 19926 395
rect 20010 378 20044 395
rect 20047 378 20081 395
rect 19888 371 19892 378
rect 19820 261 19824 329
rect 19888 291 19892 341
rect 19888 251 19897 279
rect 19984 264 19994 291
rect 19943 262 19994 264
rect 19984 261 19995 262
rect 19951 253 19985 255
rect 19993 253 19995 261
rect 19820 183 19824 251
rect 19829 207 19839 241
rect 19849 207 19863 241
rect 19888 207 19899 251
rect 19930 246 20006 253
rect 20039 251 20048 279
rect 19951 228 19985 246
rect 19993 228 19995 246
rect 19930 221 20006 228
rect 19993 213 19995 221
rect 20037 213 20048 251
rect 19984 212 19995 213
rect 19829 183 19836 207
rect 19984 183 19994 212
rect 20075 207 20087 241
rect 20097 213 20111 241
rect 20097 207 20109 213
rect 19820 103 19824 171
rect 19888 133 19892 183
rect 19888 98 19892 103
rect 19639 62 19644 96
rect 19668 62 19673 96
rect 19888 94 19926 98
rect 19888 64 19896 94
rect 19922 64 19926 94
rect 20010 94 20044 98
rect 20010 64 20014 94
rect 20040 64 20044 94
rect 19888 61 19892 64
rect 19866 55 19892 61
rect 19930 55 19952 61
rect 19984 55 20006 61
rect 20048 55 20070 61
rect 20112 55 20116 395
rect 20119 378 20124 412
rect 20148 378 20153 412
rect 20154 400 20165 412
rect 20368 395 20410 421
rect 20774 395 20816 421
rect 21031 420 21043 424
rect 21053 420 21065 424
rect 21103 420 21115 424
rect 21125 421 21137 424
rect 21295 421 21307 424
rect 21125 420 21178 421
rect 21136 412 21178 420
rect 21019 400 21030 412
rect 20300 341 20304 395
rect 20368 387 20406 395
rect 20368 380 20376 387
rect 20402 380 20406 387
rect 20778 387 20812 395
rect 20778 380 20782 387
rect 20808 380 20812 387
rect 20356 379 20422 380
rect 20762 379 20828 380
rect 20368 371 20372 379
rect 20422 365 20472 367
rect 20712 365 20762 367
rect 20462 361 20516 365
rect 20668 361 20722 365
rect 20462 356 20482 361
rect 20702 356 20722 361
rect 20472 341 20474 356
rect 20300 261 20304 329
rect 20368 305 20372 341
rect 20466 331 20474 341
rect 20482 331 20483 351
rect 20472 315 20474 331
rect 20493 322 20496 356
rect 20515 331 20516 351
rect 20525 331 20532 341
rect 20652 331 20659 341
rect 20668 331 20669 351
rect 20688 322 20691 356
rect 20701 331 20702 351
rect 20711 331 20718 341
rect 20482 315 20498 321
rect 20500 315 20516 321
rect 20668 315 20684 321
rect 20686 315 20702 321
rect 20762 315 20764 365
rect 20305 267 20341 295
rect 20305 261 20319 267
rect 20142 183 20149 207
rect 20300 183 20304 251
rect 20309 233 20319 261
rect 20329 233 20343 267
rect 20368 261 20379 305
rect 20805 267 20816 305
rect 20843 267 20879 295
rect 20530 262 20580 264
rect 20604 262 20654 264
rect 20368 233 20377 261
rect 20431 253 20465 255
rect 20410 246 20465 253
rect 20431 245 20465 246
rect 20533 253 20564 255
rect 20533 245 20567 253
rect 20368 213 20372 233
rect 20564 229 20567 245
rect 20431 228 20465 229
rect 20410 221 20465 228
rect 20533 221 20567 229
rect 20580 212 20582 262
rect 20620 253 20651 255
rect 20654 253 20656 262
rect 20843 261 20855 267
rect 20620 245 20656 253
rect 20719 253 20753 255
rect 20719 246 20774 253
rect 20719 245 20753 246
rect 20651 229 20656 245
rect 20845 233 20855 261
rect 20865 233 20879 267
rect 20620 221 20656 229
rect 20719 228 20753 229
rect 20719 221 20774 228
rect 20654 212 20656 221
rect 20300 103 20304 171
rect 20368 133 20372 183
rect 20422 159 20472 161
rect 20712 159 20762 161
rect 20472 143 20474 159
rect 20482 153 20498 159
rect 20500 153 20516 159
rect 20668 153 20684 159
rect 20686 153 20702 159
rect 20493 143 20516 152
rect 20668 143 20691 152
rect 20466 133 20474 143
rect 20472 109 20474 133
rect 20482 123 20483 143
rect 20493 118 20496 143
rect 20515 123 20516 143
rect 20525 133 20532 143
rect 20652 133 20659 143
rect 20668 123 20669 143
rect 20688 118 20691 143
rect 20701 123 20702 143
rect 20711 133 20718 143
rect 20482 109 20516 113
rect 20668 109 20702 113
rect 20762 109 20764 159
rect 20368 103 20410 104
rect 20774 103 20816 104
rect 20368 96 20372 103
rect 20263 62 20268 96
rect 20292 62 20297 96
rect 20335 62 20406 96
rect 20778 62 20812 96
rect 20815 62 20849 96
rect 20368 61 20372 62
rect 20346 55 20372 61
rect 20410 55 20432 61
rect 20752 55 20774 61
rect 20816 55 20838 61
rect 20880 55 20884 395
rect 21031 378 21036 412
rect 21060 378 21065 412
rect 21066 400 21077 412
rect 21091 400 21102 412
rect 21103 395 21178 412
rect 21254 420 21307 421
rect 21317 420 21329 424
rect 21367 420 21379 424
rect 21389 420 21401 424
rect 21254 412 21296 420
rect 21254 395 21329 412
rect 21330 400 21341 412
rect 21355 400 21366 412
rect 21068 341 21072 395
rect 21103 378 21174 395
rect 21258 378 21292 395
rect 21295 378 21329 395
rect 21136 371 21140 378
rect 21068 261 21072 329
rect 21136 291 21140 341
rect 21136 251 21145 279
rect 21232 264 21242 291
rect 21191 262 21242 264
rect 21232 261 21243 262
rect 21199 253 21233 255
rect 21241 253 21243 261
rect 21068 183 21072 251
rect 21077 207 21087 241
rect 21097 207 21111 241
rect 21136 207 21147 251
rect 21178 246 21254 253
rect 21287 251 21296 279
rect 21199 228 21233 246
rect 21241 228 21243 246
rect 21178 221 21254 228
rect 21241 213 21243 221
rect 21285 213 21296 251
rect 21232 212 21243 213
rect 21077 183 21084 207
rect 21232 183 21242 212
rect 21323 207 21335 241
rect 21345 213 21359 241
rect 21345 207 21357 213
rect 21068 103 21072 171
rect 21136 133 21140 183
rect 21136 98 21140 103
rect 20887 62 20892 96
rect 20916 62 20921 96
rect 21136 94 21174 98
rect 21136 64 21144 94
rect 21170 64 21174 94
rect 21258 94 21292 98
rect 21258 64 21262 94
rect 21288 64 21292 94
rect 21136 61 21140 64
rect 21114 55 21140 61
rect 21178 55 21200 61
rect 21232 55 21254 61
rect 21296 55 21318 61
rect 21360 55 21364 395
rect 21367 378 21372 412
rect 21396 378 21401 412
rect 21402 400 21413 412
rect 21616 395 21658 421
rect 22022 395 22064 421
rect 22279 420 22291 424
rect 22301 420 22313 424
rect 22351 420 22363 424
rect 22373 421 22385 424
rect 22543 421 22555 424
rect 22373 420 22426 421
rect 22384 412 22426 420
rect 22267 400 22278 412
rect 21548 341 21552 395
rect 21616 387 21654 395
rect 21616 380 21624 387
rect 21650 380 21654 387
rect 22026 387 22060 395
rect 22026 380 22030 387
rect 22056 380 22060 387
rect 21604 379 21670 380
rect 22010 379 22076 380
rect 21616 371 21620 379
rect 21670 365 21720 367
rect 21960 365 22010 367
rect 21710 361 21764 365
rect 21916 361 21970 365
rect 21710 356 21730 361
rect 21950 356 21970 361
rect 21720 341 21722 356
rect 21548 261 21552 329
rect 21616 305 21620 341
rect 21714 331 21722 341
rect 21730 331 21731 351
rect 21720 315 21722 331
rect 21741 322 21744 356
rect 21763 331 21764 351
rect 21773 331 21780 341
rect 21900 331 21907 341
rect 21916 331 21917 351
rect 21936 322 21939 356
rect 21949 331 21950 351
rect 21959 331 21966 341
rect 21730 315 21746 321
rect 21748 315 21764 321
rect 21916 315 21932 321
rect 21934 315 21950 321
rect 22010 315 22012 365
rect 21553 267 21589 295
rect 21553 261 21567 267
rect 21390 183 21397 207
rect 21548 183 21552 251
rect 21557 233 21567 261
rect 21577 233 21591 267
rect 21616 261 21627 305
rect 22053 267 22064 305
rect 22091 267 22127 295
rect 21778 262 21828 264
rect 21852 262 21902 264
rect 21616 233 21625 261
rect 21679 253 21713 255
rect 21658 246 21713 253
rect 21679 245 21713 246
rect 21781 253 21812 255
rect 21781 245 21815 253
rect 21616 213 21620 233
rect 21812 229 21815 245
rect 21679 228 21713 229
rect 21658 221 21713 228
rect 21781 221 21815 229
rect 21828 212 21830 262
rect 21868 253 21899 255
rect 21902 253 21904 262
rect 22091 261 22103 267
rect 21868 245 21904 253
rect 21967 253 22001 255
rect 21967 246 22022 253
rect 21967 245 22001 246
rect 21899 229 21904 245
rect 22093 233 22103 261
rect 22113 233 22127 267
rect 21868 221 21904 229
rect 21967 228 22001 229
rect 21967 221 22022 228
rect 21902 212 21904 221
rect 21548 103 21552 171
rect 21616 133 21620 183
rect 21670 159 21720 161
rect 21960 159 22010 161
rect 21720 143 21722 159
rect 21730 153 21746 159
rect 21748 153 21764 159
rect 21916 153 21932 159
rect 21934 153 21950 159
rect 21741 143 21764 152
rect 21916 143 21939 152
rect 21714 133 21722 143
rect 21720 109 21722 133
rect 21730 123 21731 143
rect 21741 118 21744 143
rect 21763 123 21764 143
rect 21773 133 21780 143
rect 21900 133 21907 143
rect 21916 123 21917 143
rect 21936 118 21939 143
rect 21949 123 21950 143
rect 21959 133 21966 143
rect 21730 109 21764 113
rect 21916 109 21950 113
rect 22010 109 22012 159
rect 21616 103 21658 104
rect 22022 103 22064 104
rect 21616 96 21620 103
rect 21511 62 21516 96
rect 21540 62 21545 96
rect 21583 62 21654 96
rect 22026 62 22060 96
rect 22063 62 22097 96
rect 21616 61 21620 62
rect 21594 55 21620 61
rect 21658 55 21680 61
rect 22000 55 22022 61
rect 22064 55 22086 61
rect 22128 55 22132 395
rect 22279 378 22284 412
rect 22308 378 22313 412
rect 22314 400 22325 412
rect 22339 400 22350 412
rect 22351 395 22426 412
rect 22502 420 22555 421
rect 22565 420 22577 424
rect 22615 420 22627 424
rect 22637 420 22649 424
rect 22502 412 22544 420
rect 22502 395 22577 412
rect 22578 400 22589 412
rect 22603 400 22614 412
rect 22316 341 22320 395
rect 22351 378 22422 395
rect 22506 378 22540 395
rect 22543 378 22577 395
rect 22384 371 22388 378
rect 22316 261 22320 329
rect 22384 291 22388 341
rect 22384 251 22393 279
rect 22480 264 22490 291
rect 22439 262 22490 264
rect 22480 261 22491 262
rect 22447 253 22481 255
rect 22489 253 22491 261
rect 22316 183 22320 251
rect 22325 207 22335 241
rect 22345 207 22359 241
rect 22384 207 22395 251
rect 22426 246 22502 253
rect 22535 251 22544 279
rect 22447 228 22481 246
rect 22489 228 22491 246
rect 22426 221 22502 228
rect 22489 213 22491 221
rect 22533 213 22544 251
rect 22480 212 22491 213
rect 22325 183 22332 207
rect 22480 183 22490 212
rect 22571 207 22583 241
rect 22593 213 22607 241
rect 22593 207 22605 213
rect 22316 103 22320 171
rect 22384 133 22388 183
rect 22384 98 22388 103
rect 22135 62 22140 96
rect 22164 62 22169 96
rect 22384 94 22422 98
rect 22384 64 22392 94
rect 22418 64 22422 94
rect 22506 94 22540 98
rect 22506 64 22510 94
rect 22536 64 22540 94
rect 22384 61 22388 64
rect 22362 55 22388 61
rect 22426 55 22448 61
rect 22480 55 22502 61
rect 22544 55 22566 61
rect 22608 55 22612 395
rect 22615 378 22620 412
rect 22644 378 22649 412
rect 22650 400 22661 412
rect 22864 395 22906 421
rect 23270 395 23312 421
rect 23527 420 23539 424
rect 23549 420 23561 424
rect 23599 420 23611 424
rect 23621 421 23633 424
rect 23791 421 23803 424
rect 23621 420 23674 421
rect 23632 412 23674 420
rect 23515 400 23526 412
rect 22796 341 22800 395
rect 22864 387 22902 395
rect 22864 380 22872 387
rect 22898 380 22902 387
rect 23274 387 23308 395
rect 23274 380 23278 387
rect 23304 380 23308 387
rect 22852 379 22918 380
rect 23258 379 23324 380
rect 22864 371 22868 379
rect 22918 365 22968 367
rect 23208 365 23258 367
rect 22958 361 23012 365
rect 23164 361 23218 365
rect 22958 356 22978 361
rect 23198 356 23218 361
rect 22968 341 22970 356
rect 22796 261 22800 329
rect 22864 305 22868 341
rect 22962 331 22970 341
rect 22978 331 22979 351
rect 22968 315 22970 331
rect 22989 322 22992 356
rect 23011 331 23012 351
rect 23021 331 23028 341
rect 23148 331 23155 341
rect 23164 331 23165 351
rect 23184 322 23187 356
rect 23197 331 23198 351
rect 23207 331 23214 341
rect 22978 315 22994 321
rect 22996 315 23012 321
rect 23164 315 23180 321
rect 23182 315 23198 321
rect 23258 315 23260 365
rect 22801 267 22837 295
rect 22801 261 22815 267
rect 22638 183 22645 207
rect 22796 183 22800 251
rect 22805 233 22815 261
rect 22825 233 22839 267
rect 22864 261 22875 305
rect 23301 267 23312 305
rect 23339 267 23375 295
rect 23026 262 23076 264
rect 23100 262 23150 264
rect 22864 233 22873 261
rect 22927 253 22961 255
rect 22906 246 22961 253
rect 22927 245 22961 246
rect 23029 253 23060 255
rect 23029 245 23063 253
rect 22864 213 22868 233
rect 23060 229 23063 245
rect 22927 228 22961 229
rect 22906 221 22961 228
rect 23029 221 23063 229
rect 23076 212 23078 262
rect 23116 253 23147 255
rect 23150 253 23152 262
rect 23339 261 23351 267
rect 23116 245 23152 253
rect 23215 253 23249 255
rect 23215 246 23270 253
rect 23215 245 23249 246
rect 23147 229 23152 245
rect 23341 233 23351 261
rect 23361 233 23375 267
rect 23116 221 23152 229
rect 23215 228 23249 229
rect 23215 221 23270 228
rect 23150 212 23152 221
rect 22796 103 22800 171
rect 22864 133 22868 183
rect 22918 159 22968 161
rect 23208 159 23258 161
rect 22968 143 22970 159
rect 22978 153 22994 159
rect 22996 153 23012 159
rect 23164 153 23180 159
rect 23182 153 23198 159
rect 22989 143 23012 152
rect 23164 143 23187 152
rect 22962 133 22970 143
rect 22968 109 22970 133
rect 22978 123 22979 143
rect 22989 118 22992 143
rect 23011 123 23012 143
rect 23021 133 23028 143
rect 23148 133 23155 143
rect 23164 123 23165 143
rect 23184 118 23187 143
rect 23197 123 23198 143
rect 23207 133 23214 143
rect 22978 109 23012 113
rect 23164 109 23198 113
rect 23258 109 23260 159
rect 22864 103 22906 104
rect 23270 103 23312 104
rect 22864 96 22868 103
rect 22759 62 22764 96
rect 22788 62 22793 96
rect 22831 62 22902 96
rect 23274 62 23308 96
rect 23311 62 23345 96
rect 22864 61 22868 62
rect 22842 55 22868 61
rect 22906 55 22928 61
rect 23248 55 23270 61
rect 23312 55 23334 61
rect 23376 55 23380 395
rect 23527 378 23532 412
rect 23556 378 23561 412
rect 23562 400 23573 412
rect 23587 400 23598 412
rect 23599 395 23674 412
rect 23750 420 23803 421
rect 23813 420 23825 424
rect 23863 420 23875 424
rect 23885 420 23897 424
rect 23750 412 23792 420
rect 23750 395 23825 412
rect 23826 400 23837 412
rect 23851 400 23862 412
rect 23564 341 23568 395
rect 23599 378 23670 395
rect 23754 378 23788 395
rect 23791 378 23825 395
rect 23632 371 23636 378
rect 23564 261 23568 329
rect 23632 291 23636 341
rect 23632 251 23641 279
rect 23728 264 23738 291
rect 23687 262 23738 264
rect 23728 261 23739 262
rect 23695 253 23729 255
rect 23737 253 23739 261
rect 23564 183 23568 251
rect 23573 207 23583 241
rect 23593 207 23607 241
rect 23632 207 23643 251
rect 23674 246 23750 253
rect 23783 251 23792 279
rect 23695 228 23729 246
rect 23737 228 23739 246
rect 23674 221 23750 228
rect 23737 213 23739 221
rect 23781 213 23792 251
rect 23728 212 23739 213
rect 23573 183 23580 207
rect 23728 183 23738 212
rect 23819 207 23831 241
rect 23841 213 23855 241
rect 23841 207 23853 213
rect 23564 103 23568 171
rect 23632 133 23636 183
rect 23632 98 23636 103
rect 23383 62 23388 96
rect 23412 62 23417 96
rect 23632 94 23670 98
rect 23632 64 23640 94
rect 23666 64 23670 94
rect 23754 94 23788 98
rect 23754 64 23758 94
rect 23784 64 23788 94
rect 23632 61 23636 64
rect 23610 55 23636 61
rect 23674 55 23696 61
rect 23728 55 23750 61
rect 23792 55 23814 61
rect 23856 55 23860 395
rect 23863 378 23868 412
rect 23892 378 23897 412
rect 23898 400 23909 412
rect 24112 395 24154 421
rect 24518 395 24560 421
rect 24775 420 24787 424
rect 24797 420 24809 424
rect 24847 420 24859 424
rect 24869 421 24881 424
rect 25039 421 25051 424
rect 24869 420 24922 421
rect 24880 412 24922 420
rect 24763 400 24774 412
rect 24044 341 24048 395
rect 24112 387 24150 395
rect 24112 380 24120 387
rect 24146 380 24150 387
rect 24522 387 24556 395
rect 24522 380 24526 387
rect 24552 380 24556 387
rect 24100 379 24166 380
rect 24506 379 24572 380
rect 24112 371 24116 379
rect 24166 365 24216 367
rect 24456 365 24506 367
rect 24206 361 24260 365
rect 24412 361 24466 365
rect 24206 356 24226 361
rect 24446 356 24466 361
rect 24216 341 24218 356
rect 24044 261 24048 329
rect 24112 305 24116 341
rect 24210 331 24218 341
rect 24226 331 24227 351
rect 24216 315 24218 331
rect 24237 322 24240 356
rect 24259 331 24260 351
rect 24269 331 24276 341
rect 24396 331 24403 341
rect 24412 331 24413 351
rect 24432 322 24435 356
rect 24445 331 24446 351
rect 24455 331 24462 341
rect 24226 315 24242 321
rect 24244 315 24260 321
rect 24412 315 24428 321
rect 24430 315 24446 321
rect 24506 315 24508 365
rect 24049 267 24085 295
rect 24049 261 24063 267
rect 23886 183 23893 207
rect 24044 183 24048 251
rect 24053 233 24063 261
rect 24073 233 24087 267
rect 24112 261 24123 305
rect 24549 267 24560 305
rect 24587 267 24623 295
rect 24274 262 24324 264
rect 24348 262 24398 264
rect 24112 233 24121 261
rect 24175 253 24209 255
rect 24154 246 24209 253
rect 24175 245 24209 246
rect 24277 253 24308 255
rect 24277 245 24311 253
rect 24112 213 24116 233
rect 24308 229 24311 245
rect 24175 228 24209 229
rect 24154 221 24209 228
rect 24277 221 24311 229
rect 24324 212 24326 262
rect 24364 253 24395 255
rect 24398 253 24400 262
rect 24587 261 24599 267
rect 24364 245 24400 253
rect 24463 253 24497 255
rect 24463 246 24518 253
rect 24463 245 24497 246
rect 24395 229 24400 245
rect 24589 233 24599 261
rect 24609 233 24623 267
rect 24364 221 24400 229
rect 24463 228 24497 229
rect 24463 221 24518 228
rect 24398 212 24400 221
rect 24044 103 24048 171
rect 24112 133 24116 183
rect 24166 159 24216 161
rect 24456 159 24506 161
rect 24216 143 24218 159
rect 24226 153 24242 159
rect 24244 153 24260 159
rect 24412 153 24428 159
rect 24430 153 24446 159
rect 24237 143 24260 152
rect 24412 143 24435 152
rect 24210 133 24218 143
rect 24216 109 24218 133
rect 24226 123 24227 143
rect 24237 118 24240 143
rect 24259 123 24260 143
rect 24269 133 24276 143
rect 24396 133 24403 143
rect 24412 123 24413 143
rect 24432 118 24435 143
rect 24445 123 24446 143
rect 24455 133 24462 143
rect 24226 109 24260 113
rect 24412 109 24446 113
rect 24506 109 24508 159
rect 24112 103 24154 104
rect 24518 103 24560 104
rect 24112 96 24116 103
rect 24007 62 24012 96
rect 24036 62 24041 96
rect 24079 62 24150 96
rect 24522 62 24556 96
rect 24559 62 24593 96
rect 24112 61 24116 62
rect 24090 55 24116 61
rect 24154 55 24176 61
rect 24496 55 24518 61
rect 24560 55 24582 61
rect 24624 55 24628 395
rect 24775 378 24780 412
rect 24804 378 24809 412
rect 24810 400 24821 412
rect 24835 400 24846 412
rect 24847 395 24922 412
rect 24998 420 25051 421
rect 25061 420 25073 424
rect 25111 420 25123 424
rect 25133 420 25145 424
rect 24998 412 25040 420
rect 24998 395 25073 412
rect 25074 400 25085 412
rect 25099 400 25110 412
rect 24812 341 24816 395
rect 24847 378 24918 395
rect 25002 378 25036 395
rect 25039 378 25073 395
rect 24880 371 24884 378
rect 24812 261 24816 329
rect 24880 291 24884 341
rect 24880 251 24889 279
rect 24976 264 24986 291
rect 24935 262 24986 264
rect 24976 261 24987 262
rect 24943 253 24977 255
rect 24985 253 24987 261
rect 24812 183 24816 251
rect 24821 207 24831 241
rect 24841 207 24855 241
rect 24880 207 24891 251
rect 24922 246 24998 253
rect 25031 251 25040 279
rect 24943 228 24977 246
rect 24985 228 24987 246
rect 24922 221 24998 228
rect 24985 213 24987 221
rect 25029 213 25040 251
rect 24976 212 24987 213
rect 24821 183 24828 207
rect 24976 183 24986 212
rect 25067 207 25079 241
rect 25089 213 25103 241
rect 25089 207 25101 213
rect 24812 103 24816 171
rect 24880 133 24884 183
rect 24880 98 24884 103
rect 24631 62 24636 96
rect 24660 62 24665 96
rect 24880 94 24918 98
rect 24880 64 24888 94
rect 24914 64 24918 94
rect 25002 94 25036 98
rect 25002 64 25006 94
rect 25032 64 25036 94
rect 24880 61 24884 64
rect 24858 55 24884 61
rect 24922 55 24944 61
rect 24976 55 24998 61
rect 25040 55 25062 61
rect 25104 55 25108 395
rect 25111 378 25116 412
rect 25140 378 25145 412
rect 25146 400 25157 412
rect 25360 395 25402 421
rect 25766 395 25808 421
rect 26023 420 26035 424
rect 26045 420 26057 424
rect 26095 420 26107 424
rect 26117 421 26129 424
rect 26287 421 26299 424
rect 26117 420 26170 421
rect 26128 412 26170 420
rect 26011 400 26022 412
rect 25292 341 25296 395
rect 25360 387 25398 395
rect 25360 380 25368 387
rect 25394 380 25398 387
rect 25770 387 25804 395
rect 25770 380 25774 387
rect 25800 380 25804 387
rect 25348 379 25414 380
rect 25754 379 25820 380
rect 25360 371 25364 379
rect 25414 365 25464 367
rect 25704 365 25754 367
rect 25454 361 25508 365
rect 25660 361 25714 365
rect 25454 356 25474 361
rect 25694 356 25714 361
rect 25464 341 25466 356
rect 25292 261 25296 329
rect 25360 305 25364 341
rect 25458 331 25466 341
rect 25474 331 25475 351
rect 25464 315 25466 331
rect 25485 322 25488 356
rect 25507 331 25508 351
rect 25517 331 25524 341
rect 25644 331 25651 341
rect 25660 331 25661 351
rect 25680 322 25683 356
rect 25693 331 25694 351
rect 25703 331 25710 341
rect 25474 315 25490 321
rect 25492 315 25508 321
rect 25660 315 25676 321
rect 25678 315 25694 321
rect 25754 315 25756 365
rect 25297 267 25333 295
rect 25297 261 25311 267
rect 25134 183 25141 207
rect 25292 183 25296 251
rect 25301 233 25311 261
rect 25321 233 25335 267
rect 25360 261 25371 305
rect 25797 267 25808 305
rect 25835 267 25871 295
rect 25522 262 25572 264
rect 25596 262 25646 264
rect 25360 233 25369 261
rect 25423 253 25457 255
rect 25402 246 25457 253
rect 25423 245 25457 246
rect 25525 253 25556 255
rect 25525 245 25559 253
rect 25360 213 25364 233
rect 25556 229 25559 245
rect 25423 228 25457 229
rect 25402 221 25457 228
rect 25525 221 25559 229
rect 25572 212 25574 262
rect 25612 253 25643 255
rect 25646 253 25648 262
rect 25835 261 25847 267
rect 25612 245 25648 253
rect 25711 253 25745 255
rect 25711 246 25766 253
rect 25711 245 25745 246
rect 25643 229 25648 245
rect 25837 233 25847 261
rect 25857 233 25871 267
rect 25612 221 25648 229
rect 25711 228 25745 229
rect 25711 221 25766 228
rect 25646 212 25648 221
rect 25292 103 25296 171
rect 25360 133 25364 183
rect 25414 159 25464 161
rect 25704 159 25754 161
rect 25464 143 25466 159
rect 25474 153 25490 159
rect 25492 153 25508 159
rect 25660 153 25676 159
rect 25678 153 25694 159
rect 25485 143 25508 152
rect 25660 143 25683 152
rect 25458 133 25466 143
rect 25464 109 25466 133
rect 25474 123 25475 143
rect 25485 118 25488 143
rect 25507 123 25508 143
rect 25517 133 25524 143
rect 25644 133 25651 143
rect 25660 123 25661 143
rect 25680 118 25683 143
rect 25693 123 25694 143
rect 25703 133 25710 143
rect 25474 109 25508 113
rect 25660 109 25694 113
rect 25754 109 25756 159
rect 25360 103 25402 104
rect 25766 103 25808 104
rect 25360 96 25364 103
rect 25255 62 25260 96
rect 25284 62 25289 96
rect 25327 62 25398 96
rect 25770 62 25804 96
rect 25807 62 25841 96
rect 25360 61 25364 62
rect 25338 55 25364 61
rect 25402 55 25424 61
rect 25744 55 25766 61
rect 25808 55 25830 61
rect 25872 55 25876 395
rect 26023 378 26028 412
rect 26052 378 26057 412
rect 26058 400 26069 412
rect 26083 400 26094 412
rect 26095 395 26170 412
rect 26246 420 26299 421
rect 26309 420 26321 424
rect 26359 420 26371 424
rect 26381 420 26393 424
rect 26246 412 26288 420
rect 26246 395 26321 412
rect 26322 400 26333 412
rect 26347 400 26358 412
rect 26060 341 26064 395
rect 26095 378 26166 395
rect 26250 378 26284 395
rect 26287 378 26321 395
rect 26128 371 26132 378
rect 26060 261 26064 329
rect 26128 291 26132 341
rect 26128 251 26137 279
rect 26224 264 26234 291
rect 26183 262 26234 264
rect 26224 261 26235 262
rect 26191 253 26225 255
rect 26233 253 26235 261
rect 26060 183 26064 251
rect 26069 207 26079 241
rect 26089 207 26103 241
rect 26128 207 26139 251
rect 26170 246 26246 253
rect 26279 251 26288 279
rect 26191 228 26225 246
rect 26233 228 26235 246
rect 26170 221 26246 228
rect 26233 213 26235 221
rect 26277 213 26288 251
rect 26224 212 26235 213
rect 26069 183 26076 207
rect 26224 183 26234 212
rect 26315 207 26327 241
rect 26337 213 26351 241
rect 26337 207 26349 213
rect 26060 103 26064 171
rect 26128 133 26132 183
rect 26128 98 26132 103
rect 25879 62 25884 96
rect 25908 62 25913 96
rect 26128 94 26166 98
rect 26128 64 26136 94
rect 26162 64 26166 94
rect 26250 94 26284 98
rect 26250 64 26254 94
rect 26280 64 26284 94
rect 26128 61 26132 64
rect 26106 55 26132 61
rect 26170 55 26192 61
rect 26224 55 26246 61
rect 26288 55 26310 61
rect 26352 55 26356 395
rect 26359 378 26364 412
rect 26388 378 26393 412
rect 26394 400 26405 412
rect 26608 395 26650 421
rect 27014 395 27056 421
rect 27271 420 27283 424
rect 27293 420 27305 424
rect 27343 420 27355 424
rect 27365 421 27377 424
rect 27535 421 27547 424
rect 27365 420 27418 421
rect 27376 412 27418 420
rect 27259 400 27270 412
rect 26540 341 26544 395
rect 26608 387 26646 395
rect 26608 380 26616 387
rect 26642 380 26646 387
rect 27018 387 27052 395
rect 27018 380 27022 387
rect 27048 380 27052 387
rect 26596 379 26662 380
rect 27002 379 27068 380
rect 26608 371 26612 379
rect 26662 365 26712 367
rect 26952 365 27002 367
rect 26702 361 26756 365
rect 26908 361 26962 365
rect 26702 356 26722 361
rect 26942 356 26962 361
rect 26712 341 26714 356
rect 26540 261 26544 329
rect 26608 305 26612 341
rect 26706 331 26714 341
rect 26722 331 26723 351
rect 26712 315 26714 331
rect 26733 322 26736 356
rect 26755 331 26756 351
rect 26765 331 26772 341
rect 26892 331 26899 341
rect 26908 331 26909 351
rect 26928 322 26931 356
rect 26941 331 26942 351
rect 26951 331 26958 341
rect 26722 315 26738 321
rect 26740 315 26756 321
rect 26908 315 26924 321
rect 26926 315 26942 321
rect 27002 315 27004 365
rect 26545 267 26581 295
rect 26545 261 26559 267
rect 26382 183 26389 207
rect 26540 183 26544 251
rect 26549 233 26559 261
rect 26569 233 26583 267
rect 26608 261 26619 305
rect 27045 267 27056 305
rect 27083 267 27119 295
rect 26770 262 26820 264
rect 26844 262 26894 264
rect 26608 233 26617 261
rect 26671 253 26705 255
rect 26650 246 26705 253
rect 26671 245 26705 246
rect 26773 253 26804 255
rect 26773 245 26807 253
rect 26608 213 26612 233
rect 26804 229 26807 245
rect 26671 228 26705 229
rect 26650 221 26705 228
rect 26773 221 26807 229
rect 26820 212 26822 262
rect 26860 253 26891 255
rect 26894 253 26896 262
rect 27083 261 27095 267
rect 26860 245 26896 253
rect 26959 253 26993 255
rect 26959 246 27014 253
rect 26959 245 26993 246
rect 26891 229 26896 245
rect 27085 233 27095 261
rect 27105 233 27119 267
rect 26860 221 26896 229
rect 26959 228 26993 229
rect 26959 221 27014 228
rect 26894 212 26896 221
rect 26540 103 26544 171
rect 26608 133 26612 183
rect 26662 159 26712 161
rect 26952 159 27002 161
rect 26712 143 26714 159
rect 26722 153 26738 159
rect 26740 153 26756 159
rect 26908 153 26924 159
rect 26926 153 26942 159
rect 26733 143 26756 152
rect 26908 143 26931 152
rect 26706 133 26714 143
rect 26712 109 26714 133
rect 26722 123 26723 143
rect 26733 118 26736 143
rect 26755 123 26756 143
rect 26765 133 26772 143
rect 26892 133 26899 143
rect 26908 123 26909 143
rect 26928 118 26931 143
rect 26941 123 26942 143
rect 26951 133 26958 143
rect 26722 109 26756 113
rect 26908 109 26942 113
rect 27002 109 27004 159
rect 26608 103 26650 104
rect 27014 103 27056 104
rect 26608 96 26612 103
rect 26503 62 26508 96
rect 26532 62 26537 96
rect 26575 62 26646 96
rect 27018 62 27052 96
rect 27055 62 27089 96
rect 26608 61 26612 62
rect 26586 55 26612 61
rect 26650 55 26672 61
rect 26992 55 27014 61
rect 27056 55 27078 61
rect 27120 55 27124 395
rect 27271 378 27276 412
rect 27300 378 27305 412
rect 27306 400 27317 412
rect 27331 400 27342 412
rect 27343 395 27418 412
rect 27494 420 27547 421
rect 27557 420 27569 424
rect 27607 420 27619 424
rect 27629 420 27641 424
rect 27494 412 27536 420
rect 27494 395 27569 412
rect 27570 400 27581 412
rect 27595 400 27606 412
rect 27308 341 27312 395
rect 27343 378 27414 395
rect 27498 378 27532 395
rect 27535 378 27569 395
rect 27376 371 27380 378
rect 27308 261 27312 329
rect 27376 291 27380 341
rect 27376 251 27385 279
rect 27472 264 27482 291
rect 27431 262 27482 264
rect 27472 261 27483 262
rect 27439 253 27473 255
rect 27481 253 27483 261
rect 27308 183 27312 251
rect 27317 207 27327 241
rect 27337 207 27351 241
rect 27376 207 27387 251
rect 27418 246 27494 253
rect 27527 251 27536 279
rect 27439 228 27473 246
rect 27481 228 27483 246
rect 27418 221 27494 228
rect 27481 213 27483 221
rect 27525 213 27536 251
rect 27472 212 27483 213
rect 27317 183 27324 207
rect 27472 183 27482 212
rect 27563 207 27575 241
rect 27585 213 27599 241
rect 27585 207 27597 213
rect 27308 103 27312 171
rect 27376 133 27380 183
rect 27376 98 27380 103
rect 27127 62 27132 96
rect 27156 62 27161 96
rect 27376 94 27414 98
rect 27376 64 27384 94
rect 27410 64 27414 94
rect 27498 94 27532 98
rect 27498 64 27502 94
rect 27528 64 27532 94
rect 27376 61 27380 64
rect 27354 55 27380 61
rect 27418 55 27440 61
rect 27472 55 27494 61
rect 27536 55 27558 61
rect 27600 55 27604 395
rect 27607 378 27612 412
rect 27636 378 27641 412
rect 27642 400 27653 412
rect 27856 395 27898 421
rect 28262 395 28304 421
rect 28519 420 28531 424
rect 28541 420 28553 424
rect 28591 420 28603 424
rect 28613 421 28625 424
rect 28783 421 28795 424
rect 28613 420 28666 421
rect 28624 412 28666 420
rect 28507 400 28518 412
rect 27788 341 27792 395
rect 27856 387 27894 395
rect 27856 380 27864 387
rect 27890 380 27894 387
rect 28266 387 28300 395
rect 28266 380 28270 387
rect 28296 380 28300 387
rect 27844 379 27910 380
rect 28250 379 28316 380
rect 27856 371 27860 379
rect 27910 365 27960 367
rect 28200 365 28250 367
rect 27950 361 28004 365
rect 28156 361 28210 365
rect 27950 356 27970 361
rect 28190 356 28210 361
rect 27960 341 27962 356
rect 27788 261 27792 329
rect 27856 305 27860 341
rect 27954 331 27962 341
rect 27970 331 27971 351
rect 27960 315 27962 331
rect 27981 322 27984 356
rect 28003 331 28004 351
rect 28013 331 28020 341
rect 28140 331 28147 341
rect 28156 331 28157 351
rect 28176 322 28179 356
rect 28189 331 28190 351
rect 28199 331 28206 341
rect 27970 315 27986 321
rect 27988 315 28004 321
rect 28156 315 28172 321
rect 28174 315 28190 321
rect 28250 315 28252 365
rect 27793 267 27829 295
rect 27793 261 27807 267
rect 27630 183 27637 207
rect 27788 183 27792 251
rect 27797 233 27807 261
rect 27817 233 27831 267
rect 27856 261 27867 305
rect 28293 267 28304 305
rect 28331 267 28367 295
rect 28018 262 28068 264
rect 28092 262 28142 264
rect 27856 233 27865 261
rect 27919 253 27953 255
rect 27898 246 27953 253
rect 27919 245 27953 246
rect 28021 253 28052 255
rect 28021 245 28055 253
rect 27856 213 27860 233
rect 28052 229 28055 245
rect 27919 228 27953 229
rect 27898 221 27953 228
rect 28021 221 28055 229
rect 28068 212 28070 262
rect 28108 253 28139 255
rect 28142 253 28144 262
rect 28331 261 28343 267
rect 28108 245 28144 253
rect 28207 253 28241 255
rect 28207 246 28262 253
rect 28207 245 28241 246
rect 28139 229 28144 245
rect 28333 233 28343 261
rect 28353 233 28367 267
rect 28108 221 28144 229
rect 28207 228 28241 229
rect 28207 221 28262 228
rect 28142 212 28144 221
rect 27788 103 27792 171
rect 27856 133 27860 183
rect 27910 159 27960 161
rect 28200 159 28250 161
rect 27960 143 27962 159
rect 27970 153 27986 159
rect 27988 153 28004 159
rect 28156 153 28172 159
rect 28174 153 28190 159
rect 27981 143 28004 152
rect 28156 143 28179 152
rect 27954 133 27962 143
rect 27960 109 27962 133
rect 27970 123 27971 143
rect 27981 118 27984 143
rect 28003 123 28004 143
rect 28013 133 28020 143
rect 28140 133 28147 143
rect 28156 123 28157 143
rect 28176 118 28179 143
rect 28189 123 28190 143
rect 28199 133 28206 143
rect 27970 109 28004 113
rect 28156 109 28190 113
rect 28250 109 28252 159
rect 27856 103 27898 104
rect 28262 103 28304 104
rect 27856 96 27860 103
rect 27751 62 27756 96
rect 27780 62 27785 96
rect 27823 62 27894 96
rect 28266 62 28300 96
rect 28303 62 28337 96
rect 27856 61 27860 62
rect 27834 55 27860 61
rect 27898 55 27920 61
rect 28240 55 28262 61
rect 28304 55 28326 61
rect 28368 55 28372 395
rect 28519 378 28524 412
rect 28548 378 28553 412
rect 28554 400 28565 412
rect 28579 400 28590 412
rect 28591 395 28666 412
rect 28742 420 28795 421
rect 28805 420 28817 424
rect 28855 420 28867 424
rect 28877 420 28889 424
rect 28742 412 28784 420
rect 28742 395 28817 412
rect 28818 400 28829 412
rect 28843 400 28854 412
rect 28556 341 28560 395
rect 28591 378 28662 395
rect 28746 378 28780 395
rect 28783 378 28817 395
rect 28624 371 28628 378
rect 28556 261 28560 329
rect 28624 291 28628 341
rect 28624 251 28633 279
rect 28720 264 28730 291
rect 28679 262 28730 264
rect 28720 261 28731 262
rect 28687 253 28721 255
rect 28729 253 28731 261
rect 28556 183 28560 251
rect 28565 207 28575 241
rect 28585 207 28599 241
rect 28624 207 28635 251
rect 28666 246 28742 253
rect 28775 251 28784 279
rect 28687 228 28721 246
rect 28729 228 28731 246
rect 28666 221 28742 228
rect 28729 213 28731 221
rect 28773 213 28784 251
rect 28720 212 28731 213
rect 28565 183 28572 207
rect 28720 183 28730 212
rect 28811 207 28823 241
rect 28833 213 28847 241
rect 28833 207 28845 213
rect 28556 103 28560 171
rect 28624 133 28628 183
rect 28624 98 28628 103
rect 28375 62 28380 96
rect 28404 62 28409 96
rect 28624 94 28662 98
rect 28624 64 28632 94
rect 28658 64 28662 94
rect 28746 94 28780 98
rect 28746 64 28750 94
rect 28776 64 28780 94
rect 28624 61 28628 64
rect 28602 55 28628 61
rect 28666 55 28688 61
rect 28720 55 28742 61
rect 28784 55 28806 61
rect 28848 55 28852 395
rect 28855 378 28860 412
rect 28884 378 28889 412
rect 28890 400 28901 412
rect 29104 395 29146 421
rect 29510 395 29552 421
rect 29767 420 29779 424
rect 29789 420 29801 424
rect 29839 420 29851 424
rect 29861 421 29873 424
rect 29861 420 29914 421
rect 29872 412 29914 420
rect 29755 400 29766 412
rect 29036 341 29040 395
rect 29104 387 29142 395
rect 29104 380 29112 387
rect 29138 380 29142 387
rect 29514 387 29548 395
rect 29514 380 29518 387
rect 29544 380 29548 387
rect 29092 379 29158 380
rect 29498 379 29564 380
rect 29104 371 29108 379
rect 29158 365 29208 367
rect 29448 365 29498 367
rect 29198 361 29252 365
rect 29404 361 29458 365
rect 29198 356 29218 361
rect 29438 356 29458 361
rect 29208 341 29210 356
rect 29036 261 29040 329
rect 29104 305 29108 341
rect 29202 331 29210 341
rect 29218 331 29219 351
rect 29208 315 29210 331
rect 29229 322 29232 356
rect 29251 331 29252 351
rect 29261 331 29268 341
rect 29388 331 29395 341
rect 29404 331 29405 351
rect 29424 322 29427 356
rect 29437 331 29438 351
rect 29447 331 29454 341
rect 29218 315 29234 321
rect 29236 315 29252 321
rect 29404 315 29420 321
rect 29422 315 29438 321
rect 29498 315 29500 365
rect 29041 267 29077 295
rect 29041 261 29055 267
rect 28878 183 28885 207
rect 29036 183 29040 251
rect 29045 233 29055 261
rect 29065 233 29079 267
rect 29104 261 29115 305
rect 29541 267 29552 305
rect 29579 267 29615 295
rect 29266 262 29316 264
rect 29340 262 29390 264
rect 29104 233 29113 261
rect 29167 253 29201 255
rect 29146 246 29201 253
rect 29167 245 29201 246
rect 29269 253 29300 255
rect 29269 245 29303 253
rect 29104 213 29108 233
rect 29300 229 29303 245
rect 29167 228 29201 229
rect 29146 221 29201 228
rect 29269 221 29303 229
rect 29316 212 29318 262
rect 29356 253 29387 255
rect 29390 253 29392 262
rect 29579 261 29591 267
rect 29356 245 29392 253
rect 29455 253 29489 255
rect 29455 246 29510 253
rect 29455 245 29489 246
rect 29387 229 29392 245
rect 29581 233 29591 261
rect 29601 233 29615 267
rect 29356 221 29392 229
rect 29455 228 29489 229
rect 29455 221 29510 228
rect 29390 212 29392 221
rect 29036 103 29040 171
rect 29104 133 29108 183
rect 29158 159 29208 161
rect 29448 159 29498 161
rect 29208 143 29210 159
rect 29218 153 29234 159
rect 29236 153 29252 159
rect 29404 153 29420 159
rect 29422 153 29438 159
rect 29229 143 29252 152
rect 29404 143 29427 152
rect 29202 133 29210 143
rect 29208 109 29210 133
rect 29218 123 29219 143
rect 29229 118 29232 143
rect 29251 123 29252 143
rect 29261 133 29268 143
rect 29388 133 29395 143
rect 29404 123 29405 143
rect 29424 118 29427 143
rect 29437 123 29438 143
rect 29447 133 29454 143
rect 29218 109 29252 113
rect 29404 109 29438 113
rect 29498 109 29500 159
rect 29104 103 29146 104
rect 29510 103 29552 104
rect 29104 96 29108 103
rect 28999 62 29004 96
rect 29028 62 29033 96
rect 29071 62 29142 96
rect 29514 62 29548 96
rect 29551 62 29585 96
rect 29104 61 29108 62
rect 29082 55 29108 61
rect 29146 55 29168 61
rect 29488 55 29510 61
rect 29552 55 29574 61
rect 29616 55 29620 395
rect 29767 378 29772 412
rect 29796 378 29801 412
rect 29802 400 29813 412
rect 29827 400 29838 412
rect 29839 395 29914 412
rect 29804 341 29808 395
rect 29839 378 29910 395
rect 29872 371 29876 378
rect 29804 261 29808 329
rect 29872 291 29876 341
rect 29872 251 29881 279
rect 29927 262 29977 264
rect 29935 253 29952 255
rect 29804 183 29808 251
rect 29813 207 29823 241
rect 29833 207 29847 241
rect 29872 207 29883 251
rect 29914 246 29969 253
rect 29935 245 29969 246
rect 29944 229 29969 245
rect 29935 228 29969 229
rect 29914 221 29969 228
rect 29977 212 29979 262
rect 29813 183 29820 207
rect 29804 103 29808 171
rect 29872 133 29876 183
rect 29872 98 29876 103
rect 29623 62 29628 96
rect 29652 62 29657 96
rect 29872 94 29910 98
rect 29872 64 29880 94
rect 29906 64 29910 94
rect 29872 61 29876 64
rect 29850 55 29876 61
rect 29914 55 29936 61
rect 38 39 80 55
rect 400 39 442 55
rect 806 39 848 55
rect 1168 39 1210 55
rect 1286 39 1328 55
rect 1648 39 1690 55
rect 2054 39 2096 55
rect 2416 39 2458 55
rect 2534 39 2576 55
rect 2896 39 2938 55
rect 3302 39 3344 55
rect 3664 39 3706 55
rect 3782 39 3824 55
rect 4144 39 4186 55
rect 4550 39 4592 55
rect 4912 39 4954 55
rect 5030 39 5072 55
rect 5392 39 5434 55
rect 5798 39 5840 55
rect 6160 39 6202 55
rect 6278 39 6320 55
rect 6640 39 6682 55
rect 7046 39 7088 55
rect 7408 39 7450 55
rect 7526 39 7568 55
rect 7888 39 7930 55
rect 8294 39 8336 55
rect 8656 39 8698 55
rect 8774 39 8816 55
rect 9136 39 9178 55
rect 9542 39 9584 55
rect 9904 39 9946 55
rect 10022 39 10064 55
rect 10384 39 10426 55
rect 10790 39 10832 55
rect 11152 39 11194 55
rect 11270 39 11312 55
rect 11632 39 11674 55
rect 12038 39 12080 55
rect 12400 39 12442 55
rect 12518 39 12560 55
rect 12880 39 12922 55
rect 13286 39 13328 55
rect 13648 39 13690 55
rect 13766 39 13808 55
rect 14128 39 14170 55
rect 14534 39 14576 55
rect 14896 39 14938 55
rect 15014 39 15056 55
rect 15376 39 15418 55
rect 15782 39 15824 55
rect 16144 39 16186 55
rect 16262 39 16304 55
rect 16624 39 16666 55
rect 17030 39 17072 55
rect 17392 39 17434 55
rect 17510 39 17552 55
rect 17872 39 17914 55
rect 18278 39 18320 55
rect 18640 39 18682 55
rect 18758 39 18800 55
rect 19120 39 19162 55
rect 19526 39 19568 55
rect 19888 39 19930 55
rect 20006 39 20048 55
rect 20368 39 20410 55
rect 20774 39 20816 55
rect 21136 39 21178 55
rect 21254 39 21296 55
rect 21616 39 21658 55
rect 22022 39 22064 55
rect 22384 39 22426 55
rect 22502 39 22544 55
rect 22864 39 22906 55
rect 23270 39 23312 55
rect 23632 39 23674 55
rect 23750 39 23792 55
rect 24112 39 24154 55
rect 24518 39 24560 55
rect 24880 39 24922 55
rect 24998 39 25040 55
rect 25360 39 25402 55
rect 25766 39 25808 55
rect 26128 39 26170 55
rect 26246 39 26288 55
rect 26608 39 26650 55
rect 27014 39 27056 55
rect 27376 39 27418 55
rect 27494 39 27536 55
rect 27856 39 27898 55
rect 28262 39 28304 55
rect 28624 39 28666 55
rect 28742 39 28784 55
rect 29104 39 29146 55
rect 29510 39 29552 55
rect 29872 39 29914 55
rect -25 25 25 27
rect 455 25 505 27
rect 557 25 607 27
rect 641 25 691 27
rect 743 25 793 27
rect 1223 25 1273 27
rect 1703 25 1753 27
rect 1805 25 1855 27
rect 1889 25 1939 27
rect 1991 25 2041 27
rect 2471 25 2521 27
rect 2951 25 3001 27
rect 3053 25 3103 27
rect 3137 25 3187 27
rect 3239 25 3289 27
rect 3719 25 3769 27
rect 4199 25 4249 27
rect 4301 25 4351 27
rect 4385 25 4435 27
rect 4487 25 4537 27
rect 4967 25 5017 27
rect 5447 25 5497 27
rect 5549 25 5599 27
rect 5633 25 5683 27
rect 5735 25 5785 27
rect 6215 25 6265 27
rect 6695 25 6745 27
rect 6797 25 6847 27
rect 6881 25 6931 27
rect 6983 25 7033 27
rect 7463 25 7513 27
rect 7943 25 7993 27
rect 8045 25 8095 27
rect 8129 25 8179 27
rect 8231 25 8281 27
rect 8711 25 8761 27
rect 9191 25 9241 27
rect 9293 25 9343 27
rect 9377 25 9427 27
rect 9479 25 9529 27
rect 9959 25 10009 27
rect 10439 25 10489 27
rect 10541 25 10591 27
rect 10625 25 10675 27
rect 10727 25 10777 27
rect 11207 25 11257 27
rect 11687 25 11737 27
rect 11789 25 11839 27
rect 11873 25 11923 27
rect 11975 25 12025 27
rect 12455 25 12505 27
rect 12935 25 12985 27
rect 13037 25 13087 27
rect 13121 25 13171 27
rect 13223 25 13273 27
rect 13703 25 13753 27
rect 14183 25 14233 27
rect 14285 25 14335 27
rect 14369 25 14419 27
rect 14471 25 14521 27
rect 14951 25 15001 27
rect 15431 25 15481 27
rect 15533 25 15583 27
rect 15617 25 15667 27
rect 15719 25 15769 27
rect 16199 25 16249 27
rect 16679 25 16729 27
rect 16781 25 16831 27
rect 16865 25 16915 27
rect 16967 25 17017 27
rect 17447 25 17497 27
rect 17927 25 17977 27
rect 18029 25 18079 27
rect 18113 25 18163 27
rect 18215 25 18265 27
rect 18695 25 18745 27
rect 19175 25 19225 27
rect 19277 25 19327 27
rect 19361 25 19411 27
rect 19463 25 19513 27
rect 19943 25 19993 27
rect 20423 25 20473 27
rect 20525 25 20575 27
rect 20609 25 20659 27
rect 20711 25 20761 27
rect 21191 25 21241 27
rect 21671 25 21721 27
rect 21773 25 21823 27
rect 21857 25 21907 27
rect 21959 25 22009 27
rect 22439 25 22489 27
rect 22919 25 22969 27
rect 23021 25 23071 27
rect 23105 25 23155 27
rect 23207 25 23257 27
rect 23687 25 23737 27
rect 24167 25 24217 27
rect 24269 25 24319 27
rect 24353 25 24403 27
rect 24455 25 24505 27
rect 24935 25 24985 27
rect 25415 25 25465 27
rect 25517 25 25567 27
rect 25601 25 25651 27
rect 25703 25 25753 27
rect 26183 25 26233 27
rect 26663 25 26713 27
rect 26765 25 26815 27
rect 26849 25 26899 27
rect 26951 25 27001 27
rect 27431 25 27481 27
rect 27911 25 27961 27
rect 28013 25 28063 27
rect 28097 25 28147 27
rect 28199 25 28249 27
rect 28679 25 28729 27
rect 29159 25 29209 27
rect 29261 25 29311 27
rect 29345 25 29395 27
rect 29447 25 29497 27
rect 29927 25 29977 27
rect 16 17 102 25
rect 378 17 464 25
rect 8 -17 17 17
rect 18 15 51 17
rect 80 15 100 17
rect 18 -17 100 15
rect 380 15 404 17
rect 429 15 438 17
rect 442 15 462 17
rect 16 -25 102 -17
rect 42 -41 76 -39
rect 16 -61 38 -55
rect 80 -61 102 -55
rect 144 -79 148 0
rect 332 -55 336 0
rect 380 -17 462 15
rect 463 -17 472 17
rect 480 -17 497 17
rect 378 -25 464 -17
rect 505 -25 507 25
rect 514 -17 548 17
rect 565 -17 582 17
rect 607 -25 609 25
rect 666 -17 683 17
rect 691 -25 693 25
rect 784 17 870 25
rect 1146 17 1232 25
rect 1264 17 1350 25
rect 1626 17 1712 25
rect 700 -17 734 17
rect 751 -17 768 17
rect 776 -17 785 17
rect 786 15 819 17
rect 848 15 868 17
rect 786 -17 868 15
rect 1148 15 1172 17
rect 1197 15 1206 17
rect 1210 15 1230 17
rect 784 -25 870 -17
rect 404 -41 438 -39
rect 810 -41 844 -39
rect 378 -61 404 -55
rect 442 -61 464 -55
rect 784 -61 806 -55
rect 848 -61 870 -55
rect 400 -79 404 -61
rect 912 -79 916 0
rect 1100 -55 1104 0
rect 1148 -17 1230 15
rect 1231 -17 1240 17
rect 1256 -17 1265 17
rect 1266 15 1299 17
rect 1328 15 1348 17
rect 1266 -17 1348 15
rect 1628 15 1652 17
rect 1677 15 1686 17
rect 1690 15 1710 17
rect 1146 -25 1232 -17
rect 1264 -25 1350 -17
rect 1172 -41 1206 -39
rect 1290 -41 1324 -39
rect 1146 -61 1172 -55
rect 1210 -61 1232 -55
rect 1264 -61 1286 -55
rect 1328 -61 1350 -55
rect 1168 -79 1172 -61
rect 1392 -79 1396 0
rect 1580 -55 1584 0
rect 1628 -17 1710 15
rect 1711 -17 1720 17
rect 1728 -17 1745 17
rect 1626 -25 1712 -17
rect 1753 -25 1755 25
rect 1762 -17 1796 17
rect 1813 -17 1830 17
rect 1855 -25 1857 25
rect 1914 -17 1931 17
rect 1939 -25 1941 25
rect 2032 17 2118 25
rect 2394 17 2480 25
rect 2512 17 2598 25
rect 2874 17 2960 25
rect 1948 -17 1982 17
rect 1999 -17 2016 17
rect 2024 -17 2033 17
rect 2034 15 2067 17
rect 2096 15 2116 17
rect 2034 -17 2116 15
rect 2396 15 2420 17
rect 2445 15 2454 17
rect 2458 15 2478 17
rect 2032 -25 2118 -17
rect 1652 -41 1686 -39
rect 2058 -41 2092 -39
rect 1626 -61 1652 -55
rect 1690 -61 1712 -55
rect 2032 -61 2054 -55
rect 2096 -61 2118 -55
rect 1648 -79 1652 -61
rect 2160 -79 2164 0
rect 2348 -55 2352 0
rect 2396 -17 2478 15
rect 2479 -17 2488 17
rect 2504 -17 2513 17
rect 2514 15 2547 17
rect 2576 15 2596 17
rect 2514 -17 2596 15
rect 2876 15 2900 17
rect 2925 15 2934 17
rect 2938 15 2958 17
rect 2394 -25 2480 -17
rect 2512 -25 2598 -17
rect 2420 -41 2454 -39
rect 2538 -41 2572 -39
rect 2394 -61 2420 -55
rect 2458 -61 2480 -55
rect 2512 -61 2534 -55
rect 2576 -61 2598 -55
rect 2416 -79 2420 -61
rect 2640 -79 2644 0
rect 2828 -55 2832 0
rect 2876 -17 2958 15
rect 2959 -17 2968 17
rect 2976 -17 2993 17
rect 2874 -25 2960 -17
rect 3001 -25 3003 25
rect 3010 -17 3044 17
rect 3061 -17 3078 17
rect 3103 -25 3105 25
rect 3162 -17 3179 17
rect 3187 -25 3189 25
rect 3280 17 3366 25
rect 3642 17 3728 25
rect 3760 17 3846 25
rect 4122 17 4208 25
rect 3196 -17 3230 17
rect 3247 -17 3264 17
rect 3272 -17 3281 17
rect 3282 15 3315 17
rect 3344 15 3364 17
rect 3282 -17 3364 15
rect 3644 15 3668 17
rect 3693 15 3702 17
rect 3706 15 3726 17
rect 3280 -25 3366 -17
rect 2900 -41 2934 -39
rect 3306 -41 3340 -39
rect 2874 -61 2900 -55
rect 2938 -61 2960 -55
rect 3280 -61 3302 -55
rect 3344 -61 3366 -55
rect 2896 -79 2900 -61
rect 3408 -79 3412 0
rect 3596 -55 3600 0
rect 3644 -17 3726 15
rect 3727 -17 3736 17
rect 3752 -17 3761 17
rect 3762 15 3795 17
rect 3824 15 3844 17
rect 3762 -17 3844 15
rect 4124 15 4148 17
rect 4173 15 4182 17
rect 4186 15 4206 17
rect 3642 -25 3728 -17
rect 3760 -25 3846 -17
rect 3668 -41 3702 -39
rect 3786 -41 3820 -39
rect 3642 -61 3668 -55
rect 3706 -61 3728 -55
rect 3760 -61 3782 -55
rect 3824 -61 3846 -55
rect 3664 -79 3668 -61
rect 3888 -79 3892 0
rect 4076 -55 4080 0
rect 4124 -17 4206 15
rect 4207 -17 4216 17
rect 4224 -17 4241 17
rect 4122 -25 4208 -17
rect 4249 -25 4251 25
rect 4258 -17 4292 17
rect 4309 -17 4326 17
rect 4351 -25 4353 25
rect 4410 -17 4427 17
rect 4435 -25 4437 25
rect 4528 17 4614 25
rect 4890 17 4976 25
rect 5008 17 5094 25
rect 5370 17 5456 25
rect 4444 -17 4478 17
rect 4495 -17 4512 17
rect 4520 -17 4529 17
rect 4530 15 4563 17
rect 4592 15 4612 17
rect 4530 -17 4612 15
rect 4892 15 4916 17
rect 4941 15 4950 17
rect 4954 15 4974 17
rect 4528 -25 4614 -17
rect 4148 -41 4182 -39
rect 4554 -41 4588 -39
rect 4122 -61 4148 -55
rect 4186 -61 4208 -55
rect 4528 -61 4550 -55
rect 4592 -61 4614 -55
rect 4144 -79 4148 -61
rect 4656 -79 4660 0
rect 4844 -55 4848 0
rect 4892 -17 4974 15
rect 4975 -17 4984 17
rect 5000 -17 5009 17
rect 5010 15 5043 17
rect 5072 15 5092 17
rect 5010 -17 5092 15
rect 5372 15 5396 17
rect 5421 15 5430 17
rect 5434 15 5454 17
rect 4890 -25 4976 -17
rect 5008 -25 5094 -17
rect 4916 -41 4950 -39
rect 5034 -41 5068 -39
rect 4890 -61 4916 -55
rect 4954 -61 4976 -55
rect 5008 -61 5030 -55
rect 5072 -61 5094 -55
rect 4912 -79 4916 -61
rect 5136 -79 5140 0
rect 5324 -55 5328 0
rect 5372 -17 5454 15
rect 5455 -17 5464 17
rect 5472 -17 5489 17
rect 5370 -25 5456 -17
rect 5497 -25 5499 25
rect 5506 -17 5540 17
rect 5557 -17 5574 17
rect 5599 -25 5601 25
rect 5658 -17 5675 17
rect 5683 -25 5685 25
rect 5776 17 5862 25
rect 6138 17 6224 25
rect 6256 17 6342 25
rect 6618 17 6704 25
rect 5692 -17 5726 17
rect 5743 -17 5760 17
rect 5768 -17 5777 17
rect 5778 15 5811 17
rect 5840 15 5860 17
rect 5778 -17 5860 15
rect 6140 15 6164 17
rect 6189 15 6198 17
rect 6202 15 6222 17
rect 5776 -25 5862 -17
rect 5396 -41 5430 -39
rect 5802 -41 5836 -39
rect 5370 -61 5396 -55
rect 5434 -61 5456 -55
rect 5776 -61 5798 -55
rect 5840 -61 5862 -55
rect 5392 -79 5396 -61
rect 5904 -79 5908 0
rect 6092 -55 6096 0
rect 6140 -17 6222 15
rect 6223 -17 6232 17
rect 6248 -17 6257 17
rect 6258 15 6291 17
rect 6320 15 6340 17
rect 6258 -17 6340 15
rect 6620 15 6644 17
rect 6669 15 6678 17
rect 6682 15 6702 17
rect 6138 -25 6224 -17
rect 6256 -25 6342 -17
rect 6164 -41 6198 -39
rect 6282 -41 6316 -39
rect 6138 -61 6164 -55
rect 6202 -61 6224 -55
rect 6256 -61 6278 -55
rect 6320 -61 6342 -55
rect 6160 -79 6164 -61
rect 6384 -79 6388 0
rect 6572 -55 6576 0
rect 6620 -17 6702 15
rect 6703 -17 6712 17
rect 6720 -17 6737 17
rect 6618 -25 6704 -17
rect 6745 -25 6747 25
rect 6754 -17 6788 17
rect 6805 -17 6822 17
rect 6847 -25 6849 25
rect 6906 -17 6923 17
rect 6931 -25 6933 25
rect 7024 17 7110 25
rect 7386 17 7472 25
rect 7504 17 7590 25
rect 7866 17 7952 25
rect 6940 -17 6974 17
rect 6991 -17 7008 17
rect 7016 -17 7025 17
rect 7026 15 7059 17
rect 7088 15 7108 17
rect 7026 -17 7108 15
rect 7388 15 7412 17
rect 7437 15 7446 17
rect 7450 15 7470 17
rect 7024 -25 7110 -17
rect 6644 -41 6678 -39
rect 7050 -41 7084 -39
rect 6618 -61 6644 -55
rect 6682 -61 6704 -55
rect 7024 -61 7046 -55
rect 7088 -61 7110 -55
rect 6640 -79 6644 -61
rect 7152 -79 7156 0
rect 7340 -55 7344 0
rect 7388 -17 7470 15
rect 7471 -17 7480 17
rect 7496 -17 7505 17
rect 7506 15 7539 17
rect 7568 15 7588 17
rect 7506 -17 7588 15
rect 7868 15 7892 17
rect 7917 15 7926 17
rect 7930 15 7950 17
rect 7386 -25 7472 -17
rect 7504 -25 7590 -17
rect 7412 -41 7446 -39
rect 7530 -41 7564 -39
rect 7386 -61 7412 -55
rect 7450 -61 7472 -55
rect 7504 -61 7526 -55
rect 7568 -61 7590 -55
rect 7408 -79 7412 -61
rect 7632 -79 7636 0
rect 7820 -55 7824 0
rect 7868 -17 7950 15
rect 7951 -17 7960 17
rect 7968 -17 7985 17
rect 7866 -25 7952 -17
rect 7993 -25 7995 25
rect 8002 -17 8036 17
rect 8053 -17 8070 17
rect 8095 -25 8097 25
rect 8154 -17 8171 17
rect 8179 -25 8181 25
rect 8272 17 8358 25
rect 8634 17 8720 25
rect 8752 17 8838 25
rect 9114 17 9200 25
rect 8188 -17 8222 17
rect 8239 -17 8256 17
rect 8264 -17 8273 17
rect 8274 15 8307 17
rect 8336 15 8356 17
rect 8274 -17 8356 15
rect 8636 15 8660 17
rect 8685 15 8694 17
rect 8698 15 8718 17
rect 8272 -25 8358 -17
rect 7892 -41 7926 -39
rect 8298 -41 8332 -39
rect 7866 -61 7892 -55
rect 7930 -61 7952 -55
rect 8272 -61 8294 -55
rect 8336 -61 8358 -55
rect 7888 -79 7892 -61
rect 8400 -79 8404 0
rect 8588 -55 8592 0
rect 8636 -17 8718 15
rect 8719 -17 8728 17
rect 8744 -17 8753 17
rect 8754 15 8787 17
rect 8816 15 8836 17
rect 8754 -17 8836 15
rect 9116 15 9140 17
rect 9165 15 9174 17
rect 9178 15 9198 17
rect 8634 -25 8720 -17
rect 8752 -25 8838 -17
rect 8660 -41 8694 -39
rect 8778 -41 8812 -39
rect 8634 -61 8660 -55
rect 8698 -61 8720 -55
rect 8752 -61 8774 -55
rect 8816 -61 8838 -55
rect 8656 -79 8660 -61
rect 8880 -79 8884 0
rect 9068 -55 9072 0
rect 9116 -17 9198 15
rect 9199 -17 9208 17
rect 9216 -17 9233 17
rect 9114 -25 9200 -17
rect 9241 -25 9243 25
rect 9250 -17 9284 17
rect 9301 -17 9318 17
rect 9343 -25 9345 25
rect 9402 -17 9419 17
rect 9427 -25 9429 25
rect 9520 17 9606 25
rect 9882 17 9968 25
rect 10000 17 10086 25
rect 10362 17 10448 25
rect 9436 -17 9470 17
rect 9487 -17 9504 17
rect 9512 -17 9521 17
rect 9522 15 9555 17
rect 9584 15 9604 17
rect 9522 -17 9604 15
rect 9884 15 9908 17
rect 9933 15 9942 17
rect 9946 15 9966 17
rect 9520 -25 9606 -17
rect 9140 -41 9174 -39
rect 9546 -41 9580 -39
rect 9114 -61 9140 -55
rect 9178 -61 9200 -55
rect 9520 -61 9542 -55
rect 9584 -61 9606 -55
rect 9136 -79 9140 -61
rect 9648 -79 9652 0
rect 9836 -55 9840 0
rect 9884 -17 9966 15
rect 9967 -17 9976 17
rect 9992 -17 10001 17
rect 10002 15 10035 17
rect 10064 15 10084 17
rect 10002 -17 10084 15
rect 10364 15 10388 17
rect 10413 15 10422 17
rect 10426 15 10446 17
rect 9882 -25 9968 -17
rect 10000 -25 10086 -17
rect 9908 -41 9942 -39
rect 10026 -41 10060 -39
rect 9882 -61 9908 -55
rect 9946 -61 9968 -55
rect 10000 -61 10022 -55
rect 10064 -61 10086 -55
rect 9904 -79 9908 -61
rect 10128 -79 10132 0
rect 10316 -55 10320 0
rect 10364 -17 10446 15
rect 10447 -17 10456 17
rect 10464 -17 10481 17
rect 10362 -25 10448 -17
rect 10489 -25 10491 25
rect 10498 -17 10532 17
rect 10549 -17 10566 17
rect 10591 -25 10593 25
rect 10650 -17 10667 17
rect 10675 -25 10677 25
rect 10768 17 10854 25
rect 11130 17 11216 25
rect 11248 17 11334 25
rect 11610 17 11696 25
rect 10684 -17 10718 17
rect 10735 -17 10752 17
rect 10760 -17 10769 17
rect 10770 15 10803 17
rect 10832 15 10852 17
rect 10770 -17 10852 15
rect 11132 15 11156 17
rect 11181 15 11190 17
rect 11194 15 11214 17
rect 10768 -25 10854 -17
rect 10388 -41 10422 -39
rect 10794 -41 10828 -39
rect 10362 -61 10388 -55
rect 10426 -61 10448 -55
rect 10768 -61 10790 -55
rect 10832 -61 10854 -55
rect 10384 -79 10388 -61
rect 10896 -79 10900 0
rect 11084 -55 11088 0
rect 11132 -17 11214 15
rect 11215 -17 11224 17
rect 11240 -17 11249 17
rect 11250 15 11283 17
rect 11312 15 11332 17
rect 11250 -17 11332 15
rect 11612 15 11636 17
rect 11661 15 11670 17
rect 11674 15 11694 17
rect 11130 -25 11216 -17
rect 11248 -25 11334 -17
rect 11156 -41 11190 -39
rect 11274 -41 11308 -39
rect 11130 -61 11156 -55
rect 11194 -61 11216 -55
rect 11248 -61 11270 -55
rect 11312 -61 11334 -55
rect 11152 -79 11156 -61
rect 11376 -79 11380 0
rect 11564 -55 11568 0
rect 11612 -17 11694 15
rect 11695 -17 11704 17
rect 11712 -17 11729 17
rect 11610 -25 11696 -17
rect 11737 -25 11739 25
rect 11746 -17 11780 17
rect 11797 -17 11814 17
rect 11839 -25 11841 25
rect 11898 -17 11915 17
rect 11923 -25 11925 25
rect 12016 17 12102 25
rect 12378 17 12464 25
rect 12496 17 12582 25
rect 12858 17 12944 25
rect 11932 -17 11966 17
rect 11983 -17 12000 17
rect 12008 -17 12017 17
rect 12018 15 12051 17
rect 12080 15 12100 17
rect 12018 -17 12100 15
rect 12380 15 12404 17
rect 12429 15 12438 17
rect 12442 15 12462 17
rect 12016 -25 12102 -17
rect 11636 -41 11670 -39
rect 12042 -41 12076 -39
rect 11610 -61 11636 -55
rect 11674 -61 11696 -55
rect 12016 -61 12038 -55
rect 12080 -61 12102 -55
rect 11632 -79 11636 -61
rect 12144 -79 12148 0
rect 12332 -55 12336 0
rect 12380 -17 12462 15
rect 12463 -17 12472 17
rect 12488 -17 12497 17
rect 12498 15 12531 17
rect 12560 15 12580 17
rect 12498 -17 12580 15
rect 12860 15 12884 17
rect 12909 15 12918 17
rect 12922 15 12942 17
rect 12378 -25 12464 -17
rect 12496 -25 12582 -17
rect 12404 -41 12438 -39
rect 12522 -41 12556 -39
rect 12378 -61 12404 -55
rect 12442 -61 12464 -55
rect 12496 -61 12518 -55
rect 12560 -61 12582 -55
rect 12400 -79 12404 -61
rect 12624 -79 12628 0
rect 12812 -55 12816 0
rect 12860 -17 12942 15
rect 12943 -17 12952 17
rect 12960 -17 12977 17
rect 12858 -25 12944 -17
rect 12985 -25 12987 25
rect 12994 -17 13028 17
rect 13045 -17 13062 17
rect 13087 -25 13089 25
rect 13146 -17 13163 17
rect 13171 -25 13173 25
rect 13264 17 13350 25
rect 13626 17 13712 25
rect 13744 17 13830 25
rect 14106 17 14192 25
rect 13180 -17 13214 17
rect 13231 -17 13248 17
rect 13256 -17 13265 17
rect 13266 15 13299 17
rect 13328 15 13348 17
rect 13266 -17 13348 15
rect 13628 15 13652 17
rect 13677 15 13686 17
rect 13690 15 13710 17
rect 13264 -25 13350 -17
rect 12884 -41 12918 -39
rect 13290 -41 13324 -39
rect 12858 -61 12884 -55
rect 12922 -61 12944 -55
rect 13264 -61 13286 -55
rect 13328 -61 13350 -55
rect 12880 -79 12884 -61
rect 13392 -79 13396 0
rect 13580 -55 13584 0
rect 13628 -17 13710 15
rect 13711 -17 13720 17
rect 13736 -17 13745 17
rect 13746 15 13779 17
rect 13808 15 13828 17
rect 13746 -17 13828 15
rect 14108 15 14132 17
rect 14157 15 14166 17
rect 14170 15 14190 17
rect 13626 -25 13712 -17
rect 13744 -25 13830 -17
rect 13652 -41 13686 -39
rect 13770 -41 13804 -39
rect 13626 -61 13652 -55
rect 13690 -61 13712 -55
rect 13744 -61 13766 -55
rect 13808 -61 13830 -55
rect 13648 -79 13652 -61
rect 13872 -79 13876 0
rect 14060 -55 14064 0
rect 14108 -17 14190 15
rect 14191 -17 14200 17
rect 14208 -17 14225 17
rect 14106 -25 14192 -17
rect 14233 -25 14235 25
rect 14242 -17 14276 17
rect 14293 -17 14310 17
rect 14335 -25 14337 25
rect 14394 -17 14411 17
rect 14419 -25 14421 25
rect 14512 17 14598 25
rect 14874 17 14960 25
rect 14992 17 15078 25
rect 15354 17 15440 25
rect 14428 -17 14462 17
rect 14479 -17 14496 17
rect 14504 -17 14513 17
rect 14514 15 14547 17
rect 14576 15 14596 17
rect 14514 -17 14596 15
rect 14876 15 14900 17
rect 14925 15 14934 17
rect 14938 15 14958 17
rect 14512 -25 14598 -17
rect 14132 -41 14166 -39
rect 14538 -41 14572 -39
rect 14106 -61 14132 -55
rect 14170 -61 14192 -55
rect 14512 -61 14534 -55
rect 14576 -61 14598 -55
rect 14128 -79 14132 -61
rect 14640 -79 14644 0
rect 14828 -55 14832 0
rect 14876 -17 14958 15
rect 14959 -17 14968 17
rect 14984 -17 14993 17
rect 14994 15 15027 17
rect 15056 15 15076 17
rect 14994 -17 15076 15
rect 15356 15 15380 17
rect 15405 15 15414 17
rect 15418 15 15438 17
rect 14874 -25 14960 -17
rect 14992 -25 15078 -17
rect 14900 -41 14934 -39
rect 15018 -41 15052 -39
rect 14874 -61 14900 -55
rect 14938 -61 14960 -55
rect 14992 -61 15014 -55
rect 15056 -61 15078 -55
rect 14896 -79 14900 -61
rect 15120 -79 15124 0
rect 15308 -55 15312 0
rect 15356 -17 15438 15
rect 15439 -17 15448 17
rect 15456 -17 15473 17
rect 15354 -25 15440 -17
rect 15481 -25 15483 25
rect 15490 -17 15524 17
rect 15541 -17 15558 17
rect 15583 -25 15585 25
rect 15642 -17 15659 17
rect 15667 -25 15669 25
rect 15760 17 15846 25
rect 16122 17 16208 25
rect 16240 17 16326 25
rect 16602 17 16688 25
rect 15676 -17 15710 17
rect 15727 -17 15744 17
rect 15752 -17 15761 17
rect 15762 15 15795 17
rect 15824 15 15844 17
rect 15762 -17 15844 15
rect 16124 15 16148 17
rect 16173 15 16182 17
rect 16186 15 16206 17
rect 15760 -25 15846 -17
rect 15380 -41 15414 -39
rect 15786 -41 15820 -39
rect 15354 -61 15380 -55
rect 15418 -61 15440 -55
rect 15760 -61 15782 -55
rect 15824 -61 15846 -55
rect 15376 -79 15380 -61
rect 15888 -79 15892 0
rect 16076 -55 16080 0
rect 16124 -17 16206 15
rect 16207 -17 16216 17
rect 16232 -17 16241 17
rect 16242 15 16275 17
rect 16304 15 16324 17
rect 16242 -17 16324 15
rect 16604 15 16628 17
rect 16653 15 16662 17
rect 16666 15 16686 17
rect 16122 -25 16208 -17
rect 16240 -25 16326 -17
rect 16148 -41 16182 -39
rect 16266 -41 16300 -39
rect 16122 -61 16148 -55
rect 16186 -61 16208 -55
rect 16240 -61 16262 -55
rect 16304 -61 16326 -55
rect 16144 -79 16148 -61
rect 16368 -79 16372 0
rect 16556 -55 16560 0
rect 16604 -17 16686 15
rect 16687 -17 16696 17
rect 16704 -17 16721 17
rect 16602 -25 16688 -17
rect 16729 -25 16731 25
rect 16738 -17 16772 17
rect 16789 -17 16806 17
rect 16831 -25 16833 25
rect 16890 -17 16907 17
rect 16915 -25 16917 25
rect 17008 17 17094 25
rect 17370 17 17456 25
rect 17488 17 17574 25
rect 17850 17 17936 25
rect 16924 -17 16958 17
rect 16975 -17 16992 17
rect 17000 -17 17009 17
rect 17010 15 17043 17
rect 17072 15 17092 17
rect 17010 -17 17092 15
rect 17372 15 17396 17
rect 17421 15 17430 17
rect 17434 15 17454 17
rect 17008 -25 17094 -17
rect 16628 -41 16662 -39
rect 17034 -41 17068 -39
rect 16602 -61 16628 -55
rect 16666 -61 16688 -55
rect 17008 -61 17030 -55
rect 17072 -61 17094 -55
rect 16624 -79 16628 -61
rect 17136 -79 17140 0
rect 17324 -55 17328 0
rect 17372 -17 17454 15
rect 17455 -17 17464 17
rect 17480 -17 17489 17
rect 17490 15 17523 17
rect 17552 15 17572 17
rect 17490 -17 17572 15
rect 17852 15 17876 17
rect 17901 15 17910 17
rect 17914 15 17934 17
rect 17370 -25 17456 -17
rect 17488 -25 17574 -17
rect 17396 -41 17430 -39
rect 17514 -41 17548 -39
rect 17370 -61 17396 -55
rect 17434 -61 17456 -55
rect 17488 -61 17510 -55
rect 17552 -61 17574 -55
rect 17392 -79 17396 -61
rect 17616 -79 17620 0
rect 17804 -55 17808 0
rect 17852 -17 17934 15
rect 17935 -17 17944 17
rect 17952 -17 17969 17
rect 17850 -25 17936 -17
rect 17977 -25 17979 25
rect 17986 -17 18020 17
rect 18037 -17 18054 17
rect 18079 -25 18081 25
rect 18138 -17 18155 17
rect 18163 -25 18165 25
rect 18256 17 18342 25
rect 18618 17 18704 25
rect 18736 17 18822 25
rect 19098 17 19184 25
rect 18172 -17 18206 17
rect 18223 -17 18240 17
rect 18248 -17 18257 17
rect 18258 15 18291 17
rect 18320 15 18340 17
rect 18258 -17 18340 15
rect 18620 15 18644 17
rect 18669 15 18678 17
rect 18682 15 18702 17
rect 18256 -25 18342 -17
rect 17876 -41 17910 -39
rect 18282 -41 18316 -39
rect 17850 -61 17876 -55
rect 17914 -61 17936 -55
rect 18256 -61 18278 -55
rect 18320 -61 18342 -55
rect 17872 -79 17876 -61
rect 18384 -79 18388 0
rect 18572 -55 18576 0
rect 18620 -17 18702 15
rect 18703 -17 18712 17
rect 18728 -17 18737 17
rect 18738 15 18771 17
rect 18800 15 18820 17
rect 18738 -17 18820 15
rect 19100 15 19124 17
rect 19149 15 19158 17
rect 19162 15 19182 17
rect 18618 -25 18704 -17
rect 18736 -25 18822 -17
rect 18644 -41 18678 -39
rect 18762 -41 18796 -39
rect 18618 -61 18644 -55
rect 18682 -61 18704 -55
rect 18736 -61 18758 -55
rect 18800 -61 18822 -55
rect 18640 -79 18644 -61
rect 18864 -79 18868 0
rect 19052 -55 19056 0
rect 19100 -17 19182 15
rect 19183 -17 19192 17
rect 19200 -17 19217 17
rect 19098 -25 19184 -17
rect 19225 -25 19227 25
rect 19234 -17 19268 17
rect 19285 -17 19302 17
rect 19327 -25 19329 25
rect 19386 -17 19403 17
rect 19411 -25 19413 25
rect 19504 17 19590 25
rect 19866 17 19952 25
rect 19984 17 20070 25
rect 20346 17 20432 25
rect 19420 -17 19454 17
rect 19471 -17 19488 17
rect 19496 -17 19505 17
rect 19506 15 19539 17
rect 19568 15 19588 17
rect 19506 -17 19588 15
rect 19868 15 19892 17
rect 19917 15 19926 17
rect 19930 15 19950 17
rect 19504 -25 19590 -17
rect 19124 -41 19158 -39
rect 19530 -41 19564 -39
rect 19098 -61 19124 -55
rect 19162 -61 19184 -55
rect 19504 -61 19526 -55
rect 19568 -61 19590 -55
rect 19120 -79 19124 -61
rect 19632 -79 19636 0
rect 19820 -55 19824 0
rect 19868 -17 19950 15
rect 19951 -17 19960 17
rect 19976 -17 19985 17
rect 19986 15 20019 17
rect 20048 15 20068 17
rect 19986 -17 20068 15
rect 20348 15 20372 17
rect 20397 15 20406 17
rect 20410 15 20430 17
rect 19866 -25 19952 -17
rect 19984 -25 20070 -17
rect 19892 -41 19926 -39
rect 20010 -41 20044 -39
rect 19866 -61 19892 -55
rect 19930 -61 19952 -55
rect 19984 -61 20006 -55
rect 20048 -61 20070 -55
rect 19888 -79 19892 -61
rect 20112 -79 20116 0
rect 20300 -55 20304 0
rect 20348 -17 20430 15
rect 20431 -17 20440 17
rect 20448 -17 20465 17
rect 20346 -25 20432 -17
rect 20473 -25 20475 25
rect 20482 -17 20516 17
rect 20533 -17 20550 17
rect 20575 -25 20577 25
rect 20634 -17 20651 17
rect 20659 -25 20661 25
rect 20752 17 20838 25
rect 21114 17 21200 25
rect 21232 17 21318 25
rect 21594 17 21680 25
rect 20668 -17 20702 17
rect 20719 -17 20736 17
rect 20744 -17 20753 17
rect 20754 15 20787 17
rect 20816 15 20836 17
rect 20754 -17 20836 15
rect 21116 15 21140 17
rect 21165 15 21174 17
rect 21178 15 21198 17
rect 20752 -25 20838 -17
rect 20372 -41 20406 -39
rect 20778 -41 20812 -39
rect 20346 -61 20372 -55
rect 20410 -61 20432 -55
rect 20752 -61 20774 -55
rect 20816 -61 20838 -55
rect 20368 -79 20372 -61
rect 20880 -79 20884 0
rect 21068 -55 21072 0
rect 21116 -17 21198 15
rect 21199 -17 21208 17
rect 21224 -17 21233 17
rect 21234 15 21267 17
rect 21296 15 21316 17
rect 21234 -17 21316 15
rect 21596 15 21620 17
rect 21645 15 21654 17
rect 21658 15 21678 17
rect 21114 -25 21200 -17
rect 21232 -25 21318 -17
rect 21140 -41 21174 -39
rect 21258 -41 21292 -39
rect 21114 -61 21140 -55
rect 21178 -61 21200 -55
rect 21232 -61 21254 -55
rect 21296 -61 21318 -55
rect 21136 -79 21140 -61
rect 21360 -79 21364 0
rect 21548 -55 21552 0
rect 21596 -17 21678 15
rect 21679 -17 21688 17
rect 21696 -17 21713 17
rect 21594 -25 21680 -17
rect 21721 -25 21723 25
rect 21730 -17 21764 17
rect 21781 -17 21798 17
rect 21823 -25 21825 25
rect 21882 -17 21899 17
rect 21907 -25 21909 25
rect 22000 17 22086 25
rect 22362 17 22448 25
rect 22480 17 22566 25
rect 22842 17 22928 25
rect 21916 -17 21950 17
rect 21967 -17 21984 17
rect 21992 -17 22001 17
rect 22002 15 22035 17
rect 22064 15 22084 17
rect 22002 -17 22084 15
rect 22364 15 22388 17
rect 22413 15 22422 17
rect 22426 15 22446 17
rect 22000 -25 22086 -17
rect 21620 -41 21654 -39
rect 22026 -41 22060 -39
rect 21594 -61 21620 -55
rect 21658 -61 21680 -55
rect 22000 -61 22022 -55
rect 22064 -61 22086 -55
rect 21616 -79 21620 -61
rect 22128 -79 22132 0
rect 22316 -55 22320 0
rect 22364 -17 22446 15
rect 22447 -17 22456 17
rect 22472 -17 22481 17
rect 22482 15 22515 17
rect 22544 15 22564 17
rect 22482 -17 22564 15
rect 22844 15 22868 17
rect 22893 15 22902 17
rect 22906 15 22926 17
rect 22362 -25 22448 -17
rect 22480 -25 22566 -17
rect 22388 -41 22422 -39
rect 22506 -41 22540 -39
rect 22362 -61 22388 -55
rect 22426 -61 22448 -55
rect 22480 -61 22502 -55
rect 22544 -61 22566 -55
rect 22384 -79 22388 -61
rect 22608 -79 22612 0
rect 22796 -55 22800 0
rect 22844 -17 22926 15
rect 22927 -17 22936 17
rect 22944 -17 22961 17
rect 22842 -25 22928 -17
rect 22969 -25 22971 25
rect 22978 -17 23012 17
rect 23029 -17 23046 17
rect 23071 -25 23073 25
rect 23130 -17 23147 17
rect 23155 -25 23157 25
rect 23248 17 23334 25
rect 23610 17 23696 25
rect 23728 17 23814 25
rect 24090 17 24176 25
rect 23164 -17 23198 17
rect 23215 -17 23232 17
rect 23240 -17 23249 17
rect 23250 15 23283 17
rect 23312 15 23332 17
rect 23250 -17 23332 15
rect 23612 15 23636 17
rect 23661 15 23670 17
rect 23674 15 23694 17
rect 23248 -25 23334 -17
rect 22868 -41 22902 -39
rect 23274 -41 23308 -39
rect 22842 -61 22868 -55
rect 22906 -61 22928 -55
rect 23248 -61 23270 -55
rect 23312 -61 23334 -55
rect 22864 -79 22868 -61
rect 23376 -79 23380 0
rect 23564 -55 23568 0
rect 23612 -17 23694 15
rect 23695 -17 23704 17
rect 23720 -17 23729 17
rect 23730 15 23763 17
rect 23792 15 23812 17
rect 23730 -17 23812 15
rect 24092 15 24116 17
rect 24141 15 24150 17
rect 24154 15 24174 17
rect 23610 -25 23696 -17
rect 23728 -25 23814 -17
rect 23636 -41 23670 -39
rect 23754 -41 23788 -39
rect 23610 -61 23636 -55
rect 23674 -61 23696 -55
rect 23728 -61 23750 -55
rect 23792 -61 23814 -55
rect 23632 -79 23636 -61
rect 23856 -79 23860 0
rect 24044 -55 24048 0
rect 24092 -17 24174 15
rect 24175 -17 24184 17
rect 24192 -17 24209 17
rect 24090 -25 24176 -17
rect 24217 -25 24219 25
rect 24226 -17 24260 17
rect 24277 -17 24294 17
rect 24319 -25 24321 25
rect 24378 -17 24395 17
rect 24403 -25 24405 25
rect 24496 17 24582 25
rect 24858 17 24944 25
rect 24976 17 25062 25
rect 25338 17 25424 25
rect 24412 -17 24446 17
rect 24463 -17 24480 17
rect 24488 -17 24497 17
rect 24498 15 24531 17
rect 24560 15 24580 17
rect 24498 -17 24580 15
rect 24860 15 24884 17
rect 24909 15 24918 17
rect 24922 15 24942 17
rect 24496 -25 24582 -17
rect 24116 -41 24150 -39
rect 24522 -41 24556 -39
rect 24090 -61 24116 -55
rect 24154 -61 24176 -55
rect 24496 -61 24518 -55
rect 24560 -61 24582 -55
rect 24112 -79 24116 -61
rect 24624 -79 24628 0
rect 24812 -55 24816 0
rect 24860 -17 24942 15
rect 24943 -17 24952 17
rect 24968 -17 24977 17
rect 24978 15 25011 17
rect 25040 15 25060 17
rect 24978 -17 25060 15
rect 25340 15 25364 17
rect 25389 15 25398 17
rect 25402 15 25422 17
rect 24858 -25 24944 -17
rect 24976 -25 25062 -17
rect 24884 -41 24918 -39
rect 25002 -41 25036 -39
rect 24858 -61 24884 -55
rect 24922 -61 24944 -55
rect 24976 -61 24998 -55
rect 25040 -61 25062 -55
rect 24880 -79 24884 -61
rect 25104 -79 25108 0
rect 25292 -55 25296 0
rect 25340 -17 25422 15
rect 25423 -17 25432 17
rect 25440 -17 25457 17
rect 25338 -25 25424 -17
rect 25465 -25 25467 25
rect 25474 -17 25508 17
rect 25525 -17 25542 17
rect 25567 -25 25569 25
rect 25626 -17 25643 17
rect 25651 -25 25653 25
rect 25744 17 25830 25
rect 26106 17 26192 25
rect 26224 17 26310 25
rect 26586 17 26672 25
rect 25660 -17 25694 17
rect 25711 -17 25728 17
rect 25736 -17 25745 17
rect 25746 15 25779 17
rect 25808 15 25828 17
rect 25746 -17 25828 15
rect 26108 15 26132 17
rect 26157 15 26166 17
rect 26170 15 26190 17
rect 25744 -25 25830 -17
rect 25364 -41 25398 -39
rect 25770 -41 25804 -39
rect 25338 -61 25364 -55
rect 25402 -61 25424 -55
rect 25744 -61 25766 -55
rect 25808 -61 25830 -55
rect 25360 -79 25364 -61
rect 25872 -79 25876 0
rect 26060 -55 26064 0
rect 26108 -17 26190 15
rect 26191 -17 26200 17
rect 26216 -17 26225 17
rect 26226 15 26259 17
rect 26288 15 26308 17
rect 26226 -17 26308 15
rect 26588 15 26612 17
rect 26637 15 26646 17
rect 26650 15 26670 17
rect 26106 -25 26192 -17
rect 26224 -25 26310 -17
rect 26132 -41 26166 -39
rect 26250 -41 26284 -39
rect 26106 -61 26132 -55
rect 26170 -61 26192 -55
rect 26224 -61 26246 -55
rect 26288 -61 26310 -55
rect 26128 -79 26132 -61
rect 26352 -79 26356 0
rect 26540 -55 26544 0
rect 26588 -17 26670 15
rect 26671 -17 26680 17
rect 26688 -17 26705 17
rect 26586 -25 26672 -17
rect 26713 -25 26715 25
rect 26722 -17 26756 17
rect 26773 -17 26790 17
rect 26815 -25 26817 25
rect 26874 -17 26891 17
rect 26899 -25 26901 25
rect 26992 17 27078 25
rect 27354 17 27440 25
rect 27472 17 27558 25
rect 27834 17 27920 25
rect 26908 -17 26942 17
rect 26959 -17 26976 17
rect 26984 -17 26993 17
rect 26994 15 27027 17
rect 27056 15 27076 17
rect 26994 -17 27076 15
rect 27356 15 27380 17
rect 27405 15 27414 17
rect 27418 15 27438 17
rect 26992 -25 27078 -17
rect 26612 -41 26646 -39
rect 27018 -41 27052 -39
rect 26586 -61 26612 -55
rect 26650 -61 26672 -55
rect 26992 -61 27014 -55
rect 27056 -61 27078 -55
rect 26608 -79 26612 -61
rect 27120 -79 27124 0
rect 27308 -55 27312 0
rect 27356 -17 27438 15
rect 27439 -17 27448 17
rect 27464 -17 27473 17
rect 27474 15 27507 17
rect 27536 15 27556 17
rect 27474 -17 27556 15
rect 27836 15 27860 17
rect 27885 15 27894 17
rect 27898 15 27918 17
rect 27354 -25 27440 -17
rect 27472 -25 27558 -17
rect 27380 -41 27414 -39
rect 27498 -41 27532 -39
rect 27354 -61 27380 -55
rect 27418 -61 27440 -55
rect 27472 -61 27494 -55
rect 27536 -61 27558 -55
rect 27376 -79 27380 -61
rect 27600 -79 27604 0
rect 27788 -55 27792 0
rect 27836 -17 27918 15
rect 27919 -17 27928 17
rect 27936 -17 27953 17
rect 27834 -25 27920 -17
rect 27961 -25 27963 25
rect 27970 -17 28004 17
rect 28021 -17 28038 17
rect 28063 -25 28065 25
rect 28122 -17 28139 17
rect 28147 -25 28149 25
rect 28240 17 28326 25
rect 28602 17 28688 25
rect 28720 17 28806 25
rect 29082 17 29168 25
rect 28156 -17 28190 17
rect 28207 -17 28224 17
rect 28232 -17 28241 17
rect 28242 15 28275 17
rect 28304 15 28324 17
rect 28242 -17 28324 15
rect 28604 15 28628 17
rect 28653 15 28662 17
rect 28666 15 28686 17
rect 28240 -25 28326 -17
rect 27860 -41 27894 -39
rect 28266 -41 28300 -39
rect 27834 -61 27860 -55
rect 27898 -61 27920 -55
rect 28240 -61 28262 -55
rect 28304 -61 28326 -55
rect 27856 -79 27860 -61
rect 28368 -79 28372 0
rect 28556 -55 28560 0
rect 28604 -17 28686 15
rect 28687 -17 28696 17
rect 28712 -17 28721 17
rect 28722 15 28755 17
rect 28784 15 28804 17
rect 28722 -17 28804 15
rect 29084 15 29108 17
rect 29133 15 29142 17
rect 29146 15 29166 17
rect 28602 -25 28688 -17
rect 28720 -25 28806 -17
rect 28628 -41 28662 -39
rect 28746 -41 28780 -39
rect 28602 -61 28628 -55
rect 28666 -61 28688 -55
rect 28720 -61 28742 -55
rect 28784 -61 28806 -55
rect 28624 -79 28628 -61
rect 28848 -79 28852 0
rect 29036 -55 29040 0
rect 29084 -17 29166 15
rect 29167 -17 29176 17
rect 29184 -17 29201 17
rect 29082 -25 29168 -17
rect 29209 -25 29211 25
rect 29218 -17 29252 17
rect 29269 -17 29286 17
rect 29311 -25 29313 25
rect 29370 -17 29387 17
rect 29395 -25 29397 25
rect 29488 17 29574 25
rect 29850 17 29936 25
rect 29404 -17 29438 17
rect 29455 -17 29472 17
rect 29480 -17 29489 17
rect 29490 15 29523 17
rect 29552 15 29572 17
rect 29490 -17 29572 15
rect 29852 15 29876 17
rect 29901 15 29910 17
rect 29914 15 29934 17
rect 29488 -25 29574 -17
rect 29108 -41 29142 -39
rect 29514 -41 29548 -39
rect 29082 -61 29108 -55
rect 29146 -61 29168 -55
rect 29488 -61 29510 -55
rect 29552 -61 29574 -55
rect 29104 -79 29108 -61
rect 29616 -79 29620 0
rect 29804 -55 29808 0
rect 29852 -17 29934 15
rect 29935 -17 29944 17
rect 29850 -25 29936 -17
rect 29977 -25 29979 25
rect 29876 -41 29910 -39
rect 29850 -61 29876 -55
rect 29914 -61 29936 -55
rect 29872 -79 29876 -61
rect 38 -105 80 -79
rect 400 -105 442 -79
rect 806 -105 848 -79
rect 1168 -105 1210 -79
rect 1286 -105 1328 -79
rect 1648 -105 1690 -79
rect 2054 -105 2096 -79
rect 2416 -105 2458 -79
rect 2534 -105 2576 -79
rect 2896 -105 2938 -79
rect 3302 -105 3344 -79
rect 3664 -105 3706 -79
rect 3782 -105 3824 -79
rect 4144 -105 4186 -79
rect 4550 -105 4592 -79
rect 4912 -105 4954 -79
rect 5030 -105 5072 -79
rect 5392 -105 5434 -79
rect 5798 -105 5840 -79
rect 6160 -105 6202 -79
rect 6278 -105 6320 -79
rect 6640 -105 6682 -79
rect 7046 -105 7088 -79
rect 7408 -105 7450 -79
rect 7526 -105 7568 -79
rect 7888 -105 7930 -79
rect 8294 -105 8336 -79
rect 8656 -105 8698 -79
rect 8774 -105 8816 -79
rect 9136 -105 9178 -79
rect 9542 -105 9584 -79
rect 9904 -105 9946 -79
rect 10022 -105 10064 -79
rect 10384 -105 10426 -79
rect 10790 -105 10832 -79
rect 11152 -105 11194 -79
rect 11270 -105 11312 -79
rect 11632 -105 11674 -79
rect 12038 -105 12080 -79
rect 12400 -105 12442 -79
rect 12518 -105 12560 -79
rect 12880 -105 12922 -79
rect 13286 -105 13328 -79
rect 13648 -105 13690 -79
rect 13766 -105 13808 -79
rect 14128 -105 14170 -79
rect 14534 -105 14576 -79
rect 14896 -105 14938 -79
rect 15014 -105 15056 -79
rect 15376 -105 15418 -79
rect 15782 -105 15824 -79
rect 16144 -105 16186 -79
rect 16262 -105 16304 -79
rect 16624 -105 16666 -79
rect 17030 -105 17072 -79
rect 17392 -105 17434 -79
rect 17510 -105 17552 -79
rect 17872 -105 17914 -79
rect 18278 -105 18320 -79
rect 18640 -105 18682 -79
rect 18758 -105 18800 -79
rect 19120 -105 19162 -79
rect 19526 -105 19568 -79
rect 19888 -105 19930 -79
rect 20006 -105 20048 -79
rect 20368 -105 20410 -79
rect 20774 -105 20816 -79
rect 21136 -105 21178 -79
rect 21254 -105 21296 -79
rect 21616 -105 21658 -79
rect 22022 -105 22064 -79
rect 22384 -105 22426 -79
rect 22502 -105 22544 -79
rect 22864 -105 22906 -79
rect 23270 -105 23312 -79
rect 23632 -105 23674 -79
rect 23750 -105 23792 -79
rect 24112 -105 24154 -79
rect 24518 -105 24560 -79
rect 24880 -105 24922 -79
rect 24998 -105 25040 -79
rect 25360 -105 25402 -79
rect 25766 -105 25808 -79
rect 26128 -105 26170 -79
rect 26246 -105 26288 -79
rect 26608 -105 26650 -79
rect 27014 -105 27056 -79
rect 27376 -105 27418 -79
rect 27494 -105 27536 -79
rect 27856 -105 27898 -79
rect 28262 -105 28304 -79
rect 28624 -105 28666 -79
rect 28742 -105 28784 -79
rect 29104 -105 29146 -79
rect 29510 -105 29552 -79
rect 29872 -105 29914 -79
<< metal1 >>
rect 78 0 114 395
rect 150 0 186 395
rect 222 79 258 420
rect 294 0 330 395
rect 366 0 402 395
rect 846 0 882 395
rect 918 0 954 395
rect 990 79 1026 420
rect 1062 0 1098 395
rect 1134 0 1170 395
rect 1326 0 1362 395
rect 1398 0 1434 395
rect 1470 79 1506 420
rect 1542 0 1578 395
rect 1614 0 1650 395
rect 2094 0 2130 395
rect 2166 0 2202 395
rect 2238 79 2274 420
rect 2310 0 2346 395
rect 2382 0 2418 395
rect 2574 0 2610 395
rect 2646 0 2682 395
rect 2718 79 2754 420
rect 2790 0 2826 395
rect 2862 0 2898 395
rect 3342 0 3378 395
rect 3414 0 3450 395
rect 3486 79 3522 420
rect 3558 0 3594 395
rect 3630 0 3666 395
rect 3822 0 3858 395
rect 3894 0 3930 395
rect 3966 79 4002 420
rect 4038 0 4074 395
rect 4110 0 4146 395
rect 4590 0 4626 395
rect 4662 0 4698 395
rect 4734 79 4770 420
rect 4806 0 4842 395
rect 4878 0 4914 395
rect 5070 0 5106 395
rect 5142 0 5178 395
rect 5214 79 5250 420
rect 5286 0 5322 395
rect 5358 0 5394 395
rect 5838 0 5874 395
rect 5910 0 5946 395
rect 5982 79 6018 420
rect 6054 0 6090 395
rect 6126 0 6162 395
rect 6318 0 6354 395
rect 6390 0 6426 395
rect 6462 79 6498 420
rect 6534 0 6570 395
rect 6606 0 6642 395
rect 7086 0 7122 395
rect 7158 0 7194 395
rect 7230 79 7266 420
rect 7302 0 7338 395
rect 7374 0 7410 395
rect 7566 0 7602 395
rect 7638 0 7674 395
rect 7710 79 7746 420
rect 7782 0 7818 395
rect 7854 0 7890 395
rect 8334 0 8370 395
rect 8406 0 8442 395
rect 8478 79 8514 420
rect 8550 0 8586 395
rect 8622 0 8658 395
rect 8814 0 8850 395
rect 8886 0 8922 395
rect 8958 79 8994 420
rect 9030 0 9066 395
rect 9102 0 9138 395
rect 9582 0 9618 395
rect 9654 0 9690 395
rect 9726 79 9762 420
rect 9798 0 9834 395
rect 9870 0 9906 395
rect 10062 0 10098 395
rect 10134 0 10170 395
rect 10206 79 10242 420
rect 10278 0 10314 395
rect 10350 0 10386 395
rect 10830 0 10866 395
rect 10902 0 10938 395
rect 10974 79 11010 420
rect 11046 0 11082 395
rect 11118 0 11154 395
rect 11310 0 11346 395
rect 11382 0 11418 395
rect 11454 79 11490 420
rect 11526 0 11562 395
rect 11598 0 11634 395
rect 12078 0 12114 395
rect 12150 0 12186 395
rect 12222 79 12258 420
rect 12294 0 12330 395
rect 12366 0 12402 395
rect 12558 0 12594 395
rect 12630 0 12666 395
rect 12702 79 12738 420
rect 12774 0 12810 395
rect 12846 0 12882 395
rect 13326 0 13362 395
rect 13398 0 13434 395
rect 13470 79 13506 420
rect 13542 0 13578 395
rect 13614 0 13650 395
rect 13806 0 13842 395
rect 13878 0 13914 395
rect 13950 79 13986 420
rect 14022 0 14058 395
rect 14094 0 14130 395
rect 14574 0 14610 395
rect 14646 0 14682 395
rect 14718 79 14754 420
rect 14790 0 14826 395
rect 14862 0 14898 395
rect 15054 0 15090 395
rect 15126 0 15162 395
rect 15198 79 15234 420
rect 15270 0 15306 395
rect 15342 0 15378 395
rect 15822 0 15858 395
rect 15894 0 15930 395
rect 15966 79 16002 420
rect 16038 0 16074 395
rect 16110 0 16146 395
rect 16302 0 16338 395
rect 16374 0 16410 395
rect 16446 79 16482 420
rect 16518 0 16554 395
rect 16590 0 16626 395
rect 17070 0 17106 395
rect 17142 0 17178 395
rect 17214 79 17250 420
rect 17286 0 17322 395
rect 17358 0 17394 395
rect 17550 0 17586 395
rect 17622 0 17658 395
rect 17694 79 17730 420
rect 17766 0 17802 395
rect 17838 0 17874 395
rect 18318 0 18354 395
rect 18390 0 18426 395
rect 18462 79 18498 420
rect 18534 0 18570 395
rect 18606 0 18642 395
rect 18798 0 18834 395
rect 18870 0 18906 395
rect 18942 79 18978 420
rect 19014 0 19050 395
rect 19086 0 19122 395
rect 19566 0 19602 395
rect 19638 0 19674 395
rect 19710 79 19746 420
rect 19782 0 19818 395
rect 19854 0 19890 395
rect 20046 0 20082 395
rect 20118 0 20154 395
rect 20190 79 20226 420
rect 20262 0 20298 395
rect 20334 0 20370 395
rect 20814 0 20850 395
rect 20886 0 20922 395
rect 20958 79 20994 420
rect 21030 0 21066 395
rect 21102 0 21138 395
rect 21294 0 21330 395
rect 21366 0 21402 395
rect 21438 79 21474 420
rect 21510 0 21546 395
rect 21582 0 21618 395
rect 22062 0 22098 395
rect 22134 0 22170 395
rect 22206 79 22242 420
rect 22278 0 22314 395
rect 22350 0 22386 395
rect 22542 0 22578 395
rect 22614 0 22650 395
rect 22686 79 22722 420
rect 22758 0 22794 395
rect 22830 0 22866 395
rect 23310 0 23346 395
rect 23382 0 23418 395
rect 23454 79 23490 420
rect 23526 0 23562 395
rect 23598 0 23634 395
rect 23790 0 23826 395
rect 23862 0 23898 395
rect 23934 79 23970 420
rect 24006 0 24042 395
rect 24078 0 24114 395
rect 24558 0 24594 395
rect 24630 0 24666 395
rect 24702 79 24738 420
rect 24774 0 24810 395
rect 24846 0 24882 395
rect 25038 0 25074 395
rect 25110 0 25146 395
rect 25182 79 25218 420
rect 25254 0 25290 395
rect 25326 0 25362 395
rect 25806 0 25842 395
rect 25878 0 25914 395
rect 25950 79 25986 420
rect 26022 0 26058 395
rect 26094 0 26130 395
rect 26286 0 26322 395
rect 26358 0 26394 395
rect 26430 79 26466 420
rect 26502 0 26538 395
rect 26574 0 26610 395
rect 27054 0 27090 395
rect 27126 0 27162 395
rect 27198 79 27234 420
rect 27270 0 27306 395
rect 27342 0 27378 395
rect 27534 0 27570 395
rect 27606 0 27642 395
rect 27678 79 27714 420
rect 27750 0 27786 395
rect 27822 0 27858 395
rect 28302 0 28338 395
rect 28374 0 28410 395
rect 28446 79 28482 420
rect 28518 0 28554 395
rect 28590 0 28626 395
rect 28782 0 28818 395
rect 28854 0 28890 395
rect 28926 79 28962 420
rect 28998 0 29034 395
rect 29070 0 29106 395
rect 29550 0 29586 395
rect 29622 0 29658 395
rect 29694 79 29730 420
rect 29766 0 29802 395
rect 29838 0 29874 395
<< metal2 >>
rect 0 323 29952 371
rect 186 199 294 275
rect 954 199 1062 275
rect 1434 199 1542 275
rect 2202 199 2310 275
rect 2682 199 2790 275
rect 3450 199 3558 275
rect 3930 199 4038 275
rect 4698 199 4806 275
rect 5178 199 5286 275
rect 5946 199 6054 275
rect 6426 199 6534 275
rect 7194 199 7302 275
rect 7674 199 7782 275
rect 8442 199 8550 275
rect 8922 199 9030 275
rect 9690 199 9798 275
rect 10170 199 10278 275
rect 10938 199 11046 275
rect 11418 199 11526 275
rect 12186 199 12294 275
rect 12666 199 12774 275
rect 13434 199 13542 275
rect 13914 199 14022 275
rect 14682 199 14790 275
rect 15162 199 15270 275
rect 15930 199 16038 275
rect 16410 199 16518 275
rect 17178 199 17286 275
rect 17658 199 17766 275
rect 18426 199 18534 275
rect 18906 199 19014 275
rect 19674 199 19782 275
rect 20154 199 20262 275
rect 20922 199 21030 275
rect 21402 199 21510 275
rect 22170 199 22278 275
rect 22650 199 22758 275
rect 23418 199 23526 275
rect 23898 199 24006 275
rect 24666 199 24774 275
rect 25146 199 25254 275
rect 25914 199 26022 275
rect 26394 199 26502 275
rect 27162 199 27270 275
rect 27642 199 27750 275
rect 28410 199 28518 275
rect 28890 199 28998 275
rect 29658 199 29766 275
rect 0 103 29952 151
rect 186 -55 294 55
rect 954 -55 1062 55
rect 1434 -55 1542 55
rect 2202 -55 2310 55
rect 2682 -55 2790 55
rect 3450 -55 3558 55
rect 3930 -55 4038 55
rect 4698 -55 4806 55
rect 5178 -55 5286 55
rect 5946 -55 6054 55
rect 6426 -55 6534 55
rect 7194 -55 7302 55
rect 7674 -55 7782 55
rect 8442 -55 8550 55
rect 8922 -55 9030 55
rect 9690 -55 9798 55
rect 10170 -55 10278 55
rect 10938 -55 11046 55
rect 11418 -55 11526 55
rect 12186 -55 12294 55
rect 12666 -55 12774 55
rect 13434 -55 13542 55
rect 13914 -55 14022 55
rect 14682 -55 14790 55
rect 15162 -55 15270 55
rect 15930 -55 16038 55
rect 16410 -55 16518 55
rect 17178 -55 17286 55
rect 17658 -55 17766 55
rect 18426 -55 18534 55
rect 18906 -55 19014 55
rect 19674 -55 19782 55
rect 20154 -55 20262 55
rect 20922 -55 21030 55
rect 21402 -55 21510 55
rect 22170 -55 22278 55
rect 22650 -55 22758 55
rect 23418 -55 23526 55
rect 23898 -55 24006 55
rect 24666 -55 24774 55
rect 25146 -55 25254 55
rect 25914 -55 26022 55
rect 26394 -55 26502 55
rect 27162 -55 27270 55
rect 27642 -55 27750 55
rect 28410 -55 28518 55
rect 28890 -55 28998 55
rect 29658 -55 29766 55
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1661296025
transform -1 0 29952 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_1
timestamp 1661296025
transform 1 0 28704 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_2
timestamp 1661296025
transform -1 0 28704 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_3
timestamp 1661296025
transform 1 0 27456 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_4
timestamp 1661296025
transform -1 0 27456 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_5
timestamp 1661296025
transform 1 0 26208 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_6
timestamp 1661296025
transform -1 0 26208 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_7
timestamp 1661296025
transform 1 0 24960 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_8
timestamp 1661296025
transform -1 0 24960 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_9
timestamp 1661296025
transform 1 0 23712 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_10
timestamp 1661296025
transform -1 0 23712 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_11
timestamp 1661296025
transform 1 0 22464 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_12
timestamp 1661296025
transform -1 0 22464 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_13
timestamp 1661296025
transform 1 0 21216 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_14
timestamp 1661296025
transform -1 0 21216 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_15
timestamp 1661296025
transform 1 0 19968 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_16
timestamp 1661296025
transform -1 0 19968 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_17
timestamp 1661296025
transform 1 0 18720 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_18
timestamp 1661296025
transform -1 0 18720 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_19
timestamp 1661296025
transform 1 0 17472 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_20
timestamp 1661296025
transform -1 0 17472 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_21
timestamp 1661296025
transform 1 0 16224 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_22
timestamp 1661296025
transform -1 0 16224 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_23
timestamp 1661296025
transform 1 0 14976 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_24
timestamp 1661296025
transform -1 0 14976 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_25
timestamp 1661296025
transform 1 0 13728 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_26
timestamp 1661296025
transform -1 0 13728 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_27
timestamp 1661296025
transform 1 0 12480 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_28
timestamp 1661296025
transform -1 0 12480 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_29
timestamp 1661296025
transform 1 0 11232 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_30
timestamp 1661296025
transform -1 0 11232 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_31
timestamp 1661296025
transform 1 0 9984 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_32
timestamp 1661296025
transform -1 0 9984 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_33
timestamp 1661296025
transform 1 0 8736 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_34
timestamp 1661296025
transform -1 0 8736 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_35
timestamp 1661296025
transform 1 0 7488 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_36
timestamp 1661296025
transform -1 0 7488 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_37
timestamp 1661296025
transform 1 0 6240 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_38
timestamp 1661296025
transform -1 0 6240 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_39
timestamp 1661296025
transform 1 0 4992 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_40
timestamp 1661296025
transform -1 0 4992 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_41
timestamp 1661296025
transform 1 0 3744 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_42
timestamp 1661296025
transform -1 0 3744 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_43
timestamp 1661296025
transform 1 0 2496 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_44
timestamp 1661296025
transform -1 0 2496 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_45
timestamp 1661296025
transform 1 0 1248 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_46
timestamp 1661296025
transform -1 0 1248 0 1 0
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_47
timestamp 1661296025
transform 1 0 0 0 1 0
box -42 -105 650 424
<< labels >>
rlabel metal1 s 78 0 114 395 4 bl_0_0
port 1 nsew
rlabel metal1 s 150 0 186 395 4 br_0_0
port 2 nsew
rlabel metal1 s 294 0 330 395 4 bl_1_0
port 3 nsew
rlabel metal1 s 366 0 402 395 4 br_1_0
port 4 nsew
rlabel metal1 s 1134 0 1170 395 4 bl_0_1
port 5 nsew
rlabel metal1 s 1062 0 1098 395 4 br_0_1
port 6 nsew
rlabel metal1 s 918 0 954 395 4 bl_1_1
port 7 nsew
rlabel metal1 s 846 0 882 395 4 br_1_1
port 8 nsew
rlabel metal1 s 1326 0 1362 395 4 bl_0_2
port 9 nsew
rlabel metal1 s 1398 0 1434 395 4 br_0_2
port 10 nsew
rlabel metal1 s 1542 0 1578 395 4 bl_1_2
port 11 nsew
rlabel metal1 s 1614 0 1650 395 4 br_1_2
port 12 nsew
rlabel metal1 s 2382 0 2418 395 4 bl_0_3
port 13 nsew
rlabel metal1 s 2310 0 2346 395 4 br_0_3
port 14 nsew
rlabel metal1 s 2166 0 2202 395 4 bl_1_3
port 15 nsew
rlabel metal1 s 2094 0 2130 395 4 br_1_3
port 16 nsew
rlabel metal1 s 2574 0 2610 395 4 bl_0_4
port 17 nsew
rlabel metal1 s 2646 0 2682 395 4 br_0_4
port 18 nsew
rlabel metal1 s 2790 0 2826 395 4 bl_1_4
port 19 nsew
rlabel metal1 s 2862 0 2898 395 4 br_1_4
port 20 nsew
rlabel metal1 s 3630 0 3666 395 4 bl_0_5
port 21 nsew
rlabel metal1 s 3558 0 3594 395 4 br_0_5
port 22 nsew
rlabel metal1 s 3414 0 3450 395 4 bl_1_5
port 23 nsew
rlabel metal1 s 3342 0 3378 395 4 br_1_5
port 24 nsew
rlabel metal1 s 3822 0 3858 395 4 bl_0_6
port 25 nsew
rlabel metal1 s 3894 0 3930 395 4 br_0_6
port 26 nsew
rlabel metal1 s 4038 0 4074 395 4 bl_1_6
port 27 nsew
rlabel metal1 s 4110 0 4146 395 4 br_1_6
port 28 nsew
rlabel metal1 s 4878 0 4914 395 4 bl_0_7
port 29 nsew
rlabel metal1 s 4806 0 4842 395 4 br_0_7
port 30 nsew
rlabel metal1 s 4662 0 4698 395 4 bl_1_7
port 31 nsew
rlabel metal1 s 4590 0 4626 395 4 br_1_7
port 32 nsew
rlabel metal1 s 5070 0 5106 395 4 bl_0_8
port 33 nsew
rlabel metal1 s 5142 0 5178 395 4 br_0_8
port 34 nsew
rlabel metal1 s 5286 0 5322 395 4 bl_1_8
port 35 nsew
rlabel metal1 s 5358 0 5394 395 4 br_1_8
port 36 nsew
rlabel metal1 s 6126 0 6162 395 4 bl_0_9
port 37 nsew
rlabel metal1 s 6054 0 6090 395 4 br_0_9
port 38 nsew
rlabel metal1 s 5910 0 5946 395 4 bl_1_9
port 39 nsew
rlabel metal1 s 5838 0 5874 395 4 br_1_9
port 40 nsew
rlabel metal1 s 6318 0 6354 395 4 bl_0_10
port 41 nsew
rlabel metal1 s 6390 0 6426 395 4 br_0_10
port 42 nsew
rlabel metal1 s 6534 0 6570 395 4 bl_1_10
port 43 nsew
rlabel metal1 s 6606 0 6642 395 4 br_1_10
port 44 nsew
rlabel metal1 s 7374 0 7410 395 4 bl_0_11
port 45 nsew
rlabel metal1 s 7302 0 7338 395 4 br_0_11
port 46 nsew
rlabel metal1 s 7158 0 7194 395 4 bl_1_11
port 47 nsew
rlabel metal1 s 7086 0 7122 395 4 br_1_11
port 48 nsew
rlabel metal1 s 7566 0 7602 395 4 bl_0_12
port 49 nsew
rlabel metal1 s 7638 0 7674 395 4 br_0_12
port 50 nsew
rlabel metal1 s 7782 0 7818 395 4 bl_1_12
port 51 nsew
rlabel metal1 s 7854 0 7890 395 4 br_1_12
port 52 nsew
rlabel metal1 s 8622 0 8658 395 4 bl_0_13
port 53 nsew
rlabel metal1 s 8550 0 8586 395 4 br_0_13
port 54 nsew
rlabel metal1 s 8406 0 8442 395 4 bl_1_13
port 55 nsew
rlabel metal1 s 8334 0 8370 395 4 br_1_13
port 56 nsew
rlabel metal1 s 8814 0 8850 395 4 bl_0_14
port 57 nsew
rlabel metal1 s 8886 0 8922 395 4 br_0_14
port 58 nsew
rlabel metal1 s 9030 0 9066 395 4 bl_1_14
port 59 nsew
rlabel metal1 s 9102 0 9138 395 4 br_1_14
port 60 nsew
rlabel metal1 s 9870 0 9906 395 4 bl_0_15
port 61 nsew
rlabel metal1 s 9798 0 9834 395 4 br_0_15
port 62 nsew
rlabel metal1 s 9654 0 9690 395 4 bl_1_15
port 63 nsew
rlabel metal1 s 9582 0 9618 395 4 br_1_15
port 64 nsew
rlabel metal1 s 10062 0 10098 395 4 bl_0_16
port 65 nsew
rlabel metal1 s 10134 0 10170 395 4 br_0_16
port 66 nsew
rlabel metal1 s 10278 0 10314 395 4 bl_1_16
port 67 nsew
rlabel metal1 s 10350 0 10386 395 4 br_1_16
port 68 nsew
rlabel metal1 s 11118 0 11154 395 4 bl_0_17
port 69 nsew
rlabel metal1 s 11046 0 11082 395 4 br_0_17
port 70 nsew
rlabel metal1 s 10902 0 10938 395 4 bl_1_17
port 71 nsew
rlabel metal1 s 10830 0 10866 395 4 br_1_17
port 72 nsew
rlabel metal1 s 11310 0 11346 395 4 bl_0_18
port 73 nsew
rlabel metal1 s 11382 0 11418 395 4 br_0_18
port 74 nsew
rlabel metal1 s 11526 0 11562 395 4 bl_1_18
port 75 nsew
rlabel metal1 s 11598 0 11634 395 4 br_1_18
port 76 nsew
rlabel metal1 s 12366 0 12402 395 4 bl_0_19
port 77 nsew
rlabel metal1 s 12294 0 12330 395 4 br_0_19
port 78 nsew
rlabel metal1 s 12150 0 12186 395 4 bl_1_19
port 79 nsew
rlabel metal1 s 12078 0 12114 395 4 br_1_19
port 80 nsew
rlabel metal1 s 12558 0 12594 395 4 bl_0_20
port 81 nsew
rlabel metal1 s 12630 0 12666 395 4 br_0_20
port 82 nsew
rlabel metal1 s 12774 0 12810 395 4 bl_1_20
port 83 nsew
rlabel metal1 s 12846 0 12882 395 4 br_1_20
port 84 nsew
rlabel metal1 s 13614 0 13650 395 4 bl_0_21
port 85 nsew
rlabel metal1 s 13542 0 13578 395 4 br_0_21
port 86 nsew
rlabel metal1 s 13398 0 13434 395 4 bl_1_21
port 87 nsew
rlabel metal1 s 13326 0 13362 395 4 br_1_21
port 88 nsew
rlabel metal1 s 13806 0 13842 395 4 bl_0_22
port 89 nsew
rlabel metal1 s 13878 0 13914 395 4 br_0_22
port 90 nsew
rlabel metal1 s 14022 0 14058 395 4 bl_1_22
port 91 nsew
rlabel metal1 s 14094 0 14130 395 4 br_1_22
port 92 nsew
rlabel metal1 s 14862 0 14898 395 4 bl_0_23
port 93 nsew
rlabel metal1 s 14790 0 14826 395 4 br_0_23
port 94 nsew
rlabel metal1 s 14646 0 14682 395 4 bl_1_23
port 95 nsew
rlabel metal1 s 14574 0 14610 395 4 br_1_23
port 96 nsew
rlabel metal1 s 15054 0 15090 395 4 bl_0_24
port 97 nsew
rlabel metal1 s 15126 0 15162 395 4 br_0_24
port 98 nsew
rlabel metal1 s 15270 0 15306 395 4 bl_1_24
port 99 nsew
rlabel metal1 s 15342 0 15378 395 4 br_1_24
port 100 nsew
rlabel metal1 s 16110 0 16146 395 4 bl_0_25
port 101 nsew
rlabel metal1 s 16038 0 16074 395 4 br_0_25
port 102 nsew
rlabel metal1 s 15894 0 15930 395 4 bl_1_25
port 103 nsew
rlabel metal1 s 15822 0 15858 395 4 br_1_25
port 104 nsew
rlabel metal1 s 16302 0 16338 395 4 bl_0_26
port 105 nsew
rlabel metal1 s 16374 0 16410 395 4 br_0_26
port 106 nsew
rlabel metal1 s 16518 0 16554 395 4 bl_1_26
port 107 nsew
rlabel metal1 s 16590 0 16626 395 4 br_1_26
port 108 nsew
rlabel metal1 s 17358 0 17394 395 4 bl_0_27
port 109 nsew
rlabel metal1 s 17286 0 17322 395 4 br_0_27
port 110 nsew
rlabel metal1 s 17142 0 17178 395 4 bl_1_27
port 111 nsew
rlabel metal1 s 17070 0 17106 395 4 br_1_27
port 112 nsew
rlabel metal1 s 17550 0 17586 395 4 bl_0_28
port 113 nsew
rlabel metal1 s 17622 0 17658 395 4 br_0_28
port 114 nsew
rlabel metal1 s 17766 0 17802 395 4 bl_1_28
port 115 nsew
rlabel metal1 s 17838 0 17874 395 4 br_1_28
port 116 nsew
rlabel metal1 s 18606 0 18642 395 4 bl_0_29
port 117 nsew
rlabel metal1 s 18534 0 18570 395 4 br_0_29
port 118 nsew
rlabel metal1 s 18390 0 18426 395 4 bl_1_29
port 119 nsew
rlabel metal1 s 18318 0 18354 395 4 br_1_29
port 120 nsew
rlabel metal1 s 18798 0 18834 395 4 bl_0_30
port 121 nsew
rlabel metal1 s 18870 0 18906 395 4 br_0_30
port 122 nsew
rlabel metal1 s 19014 0 19050 395 4 bl_1_30
port 123 nsew
rlabel metal1 s 19086 0 19122 395 4 br_1_30
port 124 nsew
rlabel metal1 s 19854 0 19890 395 4 bl_0_31
port 125 nsew
rlabel metal1 s 19782 0 19818 395 4 br_0_31
port 126 nsew
rlabel metal1 s 19638 0 19674 395 4 bl_1_31
port 127 nsew
rlabel metal1 s 19566 0 19602 395 4 br_1_31
port 128 nsew
rlabel metal1 s 20046 0 20082 395 4 bl_0_32
port 129 nsew
rlabel metal1 s 20118 0 20154 395 4 br_0_32
port 130 nsew
rlabel metal1 s 20262 0 20298 395 4 bl_1_32
port 131 nsew
rlabel metal1 s 20334 0 20370 395 4 br_1_32
port 132 nsew
rlabel metal1 s 21102 0 21138 395 4 bl_0_33
port 133 nsew
rlabel metal1 s 21030 0 21066 395 4 br_0_33
port 134 nsew
rlabel metal1 s 20886 0 20922 395 4 bl_1_33
port 135 nsew
rlabel metal1 s 20814 0 20850 395 4 br_1_33
port 136 nsew
rlabel metal1 s 21294 0 21330 395 4 bl_0_34
port 137 nsew
rlabel metal1 s 21366 0 21402 395 4 br_0_34
port 138 nsew
rlabel metal1 s 21510 0 21546 395 4 bl_1_34
port 139 nsew
rlabel metal1 s 21582 0 21618 395 4 br_1_34
port 140 nsew
rlabel metal1 s 22350 0 22386 395 4 bl_0_35
port 141 nsew
rlabel metal1 s 22278 0 22314 395 4 br_0_35
port 142 nsew
rlabel metal1 s 22134 0 22170 395 4 bl_1_35
port 143 nsew
rlabel metal1 s 22062 0 22098 395 4 br_1_35
port 144 nsew
rlabel metal1 s 22542 0 22578 395 4 bl_0_36
port 145 nsew
rlabel metal1 s 22614 0 22650 395 4 br_0_36
port 146 nsew
rlabel metal1 s 22758 0 22794 395 4 bl_1_36
port 147 nsew
rlabel metal1 s 22830 0 22866 395 4 br_1_36
port 148 nsew
rlabel metal1 s 23598 0 23634 395 4 bl_0_37
port 149 nsew
rlabel metal1 s 23526 0 23562 395 4 br_0_37
port 150 nsew
rlabel metal1 s 23382 0 23418 395 4 bl_1_37
port 151 nsew
rlabel metal1 s 23310 0 23346 395 4 br_1_37
port 152 nsew
rlabel metal1 s 23790 0 23826 395 4 bl_0_38
port 153 nsew
rlabel metal1 s 23862 0 23898 395 4 br_0_38
port 154 nsew
rlabel metal1 s 24006 0 24042 395 4 bl_1_38
port 155 nsew
rlabel metal1 s 24078 0 24114 395 4 br_1_38
port 156 nsew
rlabel metal1 s 24846 0 24882 395 4 bl_0_39
port 157 nsew
rlabel metal1 s 24774 0 24810 395 4 br_0_39
port 158 nsew
rlabel metal1 s 24630 0 24666 395 4 bl_1_39
port 159 nsew
rlabel metal1 s 24558 0 24594 395 4 br_1_39
port 160 nsew
rlabel metal1 s 25038 0 25074 395 4 bl_0_40
port 161 nsew
rlabel metal1 s 25110 0 25146 395 4 br_0_40
port 162 nsew
rlabel metal1 s 25254 0 25290 395 4 bl_1_40
port 163 nsew
rlabel metal1 s 25326 0 25362 395 4 br_1_40
port 164 nsew
rlabel metal1 s 26094 0 26130 395 4 bl_0_41
port 165 nsew
rlabel metal1 s 26022 0 26058 395 4 br_0_41
port 166 nsew
rlabel metal1 s 25878 0 25914 395 4 bl_1_41
port 167 nsew
rlabel metal1 s 25806 0 25842 395 4 br_1_41
port 168 nsew
rlabel metal1 s 26286 0 26322 395 4 bl_0_42
port 169 nsew
rlabel metal1 s 26358 0 26394 395 4 br_0_42
port 170 nsew
rlabel metal1 s 26502 0 26538 395 4 bl_1_42
port 171 nsew
rlabel metal1 s 26574 0 26610 395 4 br_1_42
port 172 nsew
rlabel metal1 s 27342 0 27378 395 4 bl_0_43
port 173 nsew
rlabel metal1 s 27270 0 27306 395 4 br_0_43
port 174 nsew
rlabel metal1 s 27126 0 27162 395 4 bl_1_43
port 175 nsew
rlabel metal1 s 27054 0 27090 395 4 br_1_43
port 176 nsew
rlabel metal1 s 27534 0 27570 395 4 bl_0_44
port 177 nsew
rlabel metal1 s 27606 0 27642 395 4 br_0_44
port 178 nsew
rlabel metal1 s 27750 0 27786 395 4 bl_1_44
port 179 nsew
rlabel metal1 s 27822 0 27858 395 4 br_1_44
port 180 nsew
rlabel metal1 s 28590 0 28626 395 4 bl_0_45
port 181 nsew
rlabel metal1 s 28518 0 28554 395 4 br_0_45
port 182 nsew
rlabel metal1 s 28374 0 28410 395 4 bl_1_45
port 183 nsew
rlabel metal1 s 28302 0 28338 395 4 br_1_45
port 184 nsew
rlabel metal1 s 28782 0 28818 395 4 bl_0_46
port 185 nsew
rlabel metal1 s 28854 0 28890 395 4 br_0_46
port 186 nsew
rlabel metal1 s 28998 0 29034 395 4 bl_1_46
port 187 nsew
rlabel metal1 s 29070 0 29106 395 4 br_1_46
port 188 nsew
rlabel metal1 s 29838 0 29874 395 4 bl_0_47
port 189 nsew
rlabel metal1 s 29766 0 29802 395 4 br_0_47
port 190 nsew
rlabel metal1 s 29622 0 29658 395 4 bl_1_47
port 191 nsew
rlabel metal1 s 29550 0 29586 395 4 br_1_47
port 192 nsew
rlabel metal2 s 0 323 29952 371 4 wl_0_0
port 193 nsew
rlabel metal2 s 0 103 29952 151 4 wl_1_0
port 194 nsew
rlabel metal1 s 3966 79 4002 420 4 vdd
port 195 nsew
rlabel metal1 s 11454 79 11490 420 4 vdd
port 195 nsew
rlabel metal1 s 19710 79 19746 420 4 vdd
port 195 nsew
rlabel metal1 s 15198 79 15234 420 4 vdd
port 195 nsew
rlabel metal1 s 15966 79 16002 420 4 vdd
port 195 nsew
rlabel metal1 s 5982 79 6018 420 4 vdd
port 195 nsew
rlabel metal1 s 12222 79 12258 420 4 vdd
port 195 nsew
rlabel metal1 s 10206 79 10242 420 4 vdd
port 195 nsew
rlabel metal1 s 17214 79 17250 420 4 vdd
port 195 nsew
rlabel metal1 s 25182 79 25218 420 4 vdd
port 195 nsew
rlabel metal1 s 22206 79 22242 420 4 vdd
port 195 nsew
rlabel metal1 s 28446 79 28482 420 4 vdd
port 195 nsew
rlabel metal1 s 24702 79 24738 420 4 vdd
port 195 nsew
rlabel metal1 s 18942 79 18978 420 4 vdd
port 195 nsew
rlabel metal1 s 2238 79 2274 420 4 vdd
port 195 nsew
rlabel metal1 s 10974 79 11010 420 4 vdd
port 195 nsew
rlabel metal1 s 12702 79 12738 420 4 vdd
port 195 nsew
rlabel metal1 s 9726 79 9762 420 4 vdd
port 195 nsew
rlabel metal1 s 13950 79 13986 420 4 vdd
port 195 nsew
rlabel metal1 s 23934 79 23970 420 4 vdd
port 195 nsew
rlabel metal1 s 8478 79 8514 420 4 vdd
port 195 nsew
rlabel metal1 s 20958 79 20994 420 4 vdd
port 195 nsew
rlabel metal1 s 990 79 1026 420 4 vdd
port 195 nsew
rlabel metal1 s 13470 79 13506 420 4 vdd
port 195 nsew
rlabel metal1 s 27678 79 27714 420 4 vdd
port 195 nsew
rlabel metal1 s 2718 79 2754 420 4 vdd
port 195 nsew
rlabel metal1 s 222 79 258 420 4 vdd
port 195 nsew
rlabel metal1 s 28926 79 28962 420 4 vdd
port 195 nsew
rlabel metal1 s 7230 79 7266 420 4 vdd
port 195 nsew
rlabel metal1 s 3486 79 3522 420 4 vdd
port 195 nsew
rlabel metal1 s 25950 79 25986 420 4 vdd
port 195 nsew
rlabel metal1 s 29694 79 29730 420 4 vdd
port 195 nsew
rlabel metal1 s 1470 79 1506 420 4 vdd
port 195 nsew
rlabel metal1 s 6462 79 6498 420 4 vdd
port 195 nsew
rlabel metal1 s 26430 79 26466 420 4 vdd
port 195 nsew
rlabel metal1 s 14718 79 14754 420 4 vdd
port 195 nsew
rlabel metal1 s 23454 79 23490 420 4 vdd
port 195 nsew
rlabel metal1 s 21438 79 21474 420 4 vdd
port 195 nsew
rlabel metal1 s 18462 79 18498 420 4 vdd
port 195 nsew
rlabel metal1 s 20190 79 20226 420 4 vdd
port 195 nsew
rlabel metal1 s 4734 79 4770 420 4 vdd
port 195 nsew
rlabel metal1 s 5214 79 5250 420 4 vdd
port 195 nsew
rlabel metal1 s 22686 79 22722 420 4 vdd
port 195 nsew
rlabel metal1 s 16446 79 16482 420 4 vdd
port 195 nsew
rlabel metal1 s 17694 79 17730 420 4 vdd
port 195 nsew
rlabel metal1 s 27198 79 27234 420 4 vdd
port 195 nsew
rlabel metal1 s 7710 79 7746 420 4 vdd
port 195 nsew
rlabel metal1 s 8958 79 8994 420 4 vdd
port 195 nsew
rlabel metal2 s 27162 199 27270 275 4 gnd
port 196 nsew
rlabel metal2 s 25914 -55 26022 55 4 gnd
port 196 nsew
rlabel metal2 s 9690 -55 9798 55 4 gnd
port 196 nsew
rlabel metal2 s 17658 199 17766 275 4 gnd
port 196 nsew
rlabel metal2 s 10938 199 11046 275 4 gnd
port 196 nsew
rlabel metal2 s 12666 -55 12774 55 4 gnd
port 196 nsew
rlabel metal2 s 8922 -55 9030 55 4 gnd
port 196 nsew
rlabel metal2 s 13434 -55 13542 55 4 gnd
port 196 nsew
rlabel metal2 s 10170 -55 10278 55 4 gnd
port 196 nsew
rlabel metal2 s 13434 199 13542 275 4 gnd
port 196 nsew
rlabel metal2 s 3450 -55 3558 55 4 gnd
port 196 nsew
rlabel metal2 s 4698 -55 4806 55 4 gnd
port 196 nsew
rlabel metal2 s 2682 199 2790 275 4 gnd
port 196 nsew
rlabel metal2 s 15930 199 16038 275 4 gnd
port 196 nsew
rlabel metal2 s 27642 -55 27750 55 4 gnd
port 196 nsew
rlabel metal2 s 28410 199 28518 275 4 gnd
port 196 nsew
rlabel metal2 s 23418 199 23526 275 4 gnd
port 196 nsew
rlabel metal2 s 29658 199 29766 275 4 gnd
port 196 nsew
rlabel metal2 s 15930 -55 16038 55 4 gnd
port 196 nsew
rlabel metal2 s 6426 199 6534 275 4 gnd
port 196 nsew
rlabel metal2 s 12666 199 12774 275 4 gnd
port 196 nsew
rlabel metal2 s 22170 -55 22278 55 4 gnd
port 196 nsew
rlabel metal2 s 28890 -55 28998 55 4 gnd
port 196 nsew
rlabel metal2 s 21402 199 21510 275 4 gnd
port 196 nsew
rlabel metal2 s 12186 -55 12294 55 4 gnd
port 196 nsew
rlabel metal2 s 8442 199 8550 275 4 gnd
port 196 nsew
rlabel metal2 s 954 199 1062 275 4 gnd
port 196 nsew
rlabel metal2 s 16410 199 16518 275 4 gnd
port 196 nsew
rlabel metal2 s 22650 -55 22758 55 4 gnd
port 196 nsew
rlabel metal2 s 186 199 294 275 4 gnd
port 196 nsew
rlabel metal2 s 12186 199 12294 275 4 gnd
port 196 nsew
rlabel metal2 s 13914 -55 14022 55 4 gnd
port 196 nsew
rlabel metal2 s 24666 199 24774 275 4 gnd
port 196 nsew
rlabel metal2 s 28890 199 28998 275 4 gnd
port 196 nsew
rlabel metal2 s 25146 -55 25254 55 4 gnd
port 196 nsew
rlabel metal2 s 23898 199 24006 275 4 gnd
port 196 nsew
rlabel metal2 s 11418 -55 11526 55 4 gnd
port 196 nsew
rlabel metal2 s 5178 -55 5286 55 4 gnd
port 196 nsew
rlabel metal2 s 26394 199 26502 275 4 gnd
port 196 nsew
rlabel metal2 s 8442 -55 8550 55 4 gnd
port 196 nsew
rlabel metal2 s 186 -55 294 55 4 gnd
port 196 nsew
rlabel metal2 s 3930 -55 4038 55 4 gnd
port 196 nsew
rlabel metal2 s 2202 -55 2310 55 4 gnd
port 196 nsew
rlabel metal2 s 3450 199 3558 275 4 gnd
port 196 nsew
rlabel metal2 s 17178 -55 17286 55 4 gnd
port 196 nsew
rlabel metal2 s 2682 -55 2790 55 4 gnd
port 196 nsew
rlabel metal2 s 17178 199 17286 275 4 gnd
port 196 nsew
rlabel metal2 s 7194 199 7302 275 4 gnd
port 196 nsew
rlabel metal2 s 20922 199 21030 275 4 gnd
port 196 nsew
rlabel metal2 s 2202 199 2310 275 4 gnd
port 196 nsew
rlabel metal2 s 18906 199 19014 275 4 gnd
port 196 nsew
rlabel metal2 s 1434 199 1542 275 4 gnd
port 196 nsew
rlabel metal2 s 20154 -55 20262 55 4 gnd
port 196 nsew
rlabel metal2 s 27162 -55 27270 55 4 gnd
port 196 nsew
rlabel metal2 s 20154 199 20262 275 4 gnd
port 196 nsew
rlabel metal2 s 5946 199 6054 275 4 gnd
port 196 nsew
rlabel metal2 s 15162 199 15270 275 4 gnd
port 196 nsew
rlabel metal2 s 10170 199 10278 275 4 gnd
port 196 nsew
rlabel metal2 s 18906 -55 19014 55 4 gnd
port 196 nsew
rlabel metal2 s 6426 -55 6534 55 4 gnd
port 196 nsew
rlabel metal2 s 20922 -55 21030 55 4 gnd
port 196 nsew
rlabel metal2 s 1434 -55 1542 55 4 gnd
port 196 nsew
rlabel metal2 s 24666 -55 24774 55 4 gnd
port 196 nsew
rlabel metal2 s 8922 199 9030 275 4 gnd
port 196 nsew
rlabel metal2 s 7674 199 7782 275 4 gnd
port 196 nsew
rlabel metal2 s 29658 -55 29766 55 4 gnd
port 196 nsew
rlabel metal2 s 21402 -55 21510 55 4 gnd
port 196 nsew
rlabel metal2 s 7194 -55 7302 55 4 gnd
port 196 nsew
rlabel metal2 s 18426 199 18534 275 4 gnd
port 196 nsew
rlabel metal2 s 4698 199 4806 275 4 gnd
port 196 nsew
rlabel metal2 s 17658 -55 17766 55 4 gnd
port 196 nsew
rlabel metal2 s 14682 199 14790 275 4 gnd
port 196 nsew
rlabel metal2 s 28410 -55 28518 55 4 gnd
port 196 nsew
rlabel metal2 s 19674 199 19782 275 4 gnd
port 196 nsew
rlabel metal2 s 9690 199 9798 275 4 gnd
port 196 nsew
rlabel metal2 s 15162 -55 15270 55 4 gnd
port 196 nsew
rlabel metal2 s 13914 199 14022 275 4 gnd
port 196 nsew
rlabel metal2 s 25914 199 26022 275 4 gnd
port 196 nsew
rlabel metal2 s 3930 199 4038 275 4 gnd
port 196 nsew
rlabel metal2 s 22170 199 22278 275 4 gnd
port 196 nsew
rlabel metal2 s 26394 -55 26502 55 4 gnd
port 196 nsew
rlabel metal2 s 23898 -55 24006 55 4 gnd
port 196 nsew
rlabel metal2 s 7674 -55 7782 55 4 gnd
port 196 nsew
rlabel metal2 s 23418 -55 23526 55 4 gnd
port 196 nsew
rlabel metal2 s 18426 -55 18534 55 4 gnd
port 196 nsew
rlabel metal2 s 25146 199 25254 275 4 gnd
port 196 nsew
rlabel metal2 s 19674 -55 19782 55 4 gnd
port 196 nsew
rlabel metal2 s 5946 -55 6054 55 4 gnd
port 196 nsew
rlabel metal2 s 27642 199 27750 275 4 gnd
port 196 nsew
rlabel metal2 s 22650 199 22758 275 4 gnd
port 196 nsew
rlabel metal2 s 11418 199 11526 275 4 gnd
port 196 nsew
rlabel metal2 s 5178 199 5286 275 4 gnd
port 196 nsew
rlabel metal2 s 10938 -55 11046 55 4 gnd
port 196 nsew
rlabel metal2 s 16410 -55 16518 55 4 gnd
port 196 nsew
rlabel metal2 s 954 -55 1062 55 4 gnd
port 196 nsew
rlabel metal2 s 14682 -55 14790 55 4 gnd
port 196 nsew
<< properties >>
string FIXED_BBOX 0 0 29952 395
<< end >>
