magic
tech sky130B
magscale 1 2
timestamp 1661277727
<< pwell >>
rect -510 2220 520 3420
<< psubdiff >>
rect -500 3354 -430 3390
rect -500 3320 -480 3354
rect -446 3320 -430 3354
rect -500 3284 -430 3320
rect -500 3250 -480 3284
rect -446 3250 -430 3284
rect -500 3214 -430 3250
rect -500 3180 -480 3214
rect -446 3180 -430 3214
rect -500 3144 -430 3180
rect -500 3110 -480 3144
rect -446 3110 -430 3144
rect -500 3074 -430 3110
rect -500 3040 -480 3074
rect -446 3040 -430 3074
rect -500 3004 -430 3040
rect -500 2970 -480 3004
rect -446 2970 -430 3004
rect -500 2934 -430 2970
rect -500 2900 -480 2934
rect -446 2900 -430 2934
rect -500 2864 -430 2900
rect -500 2830 -480 2864
rect -446 2830 -430 2864
rect -500 2794 -430 2830
rect -500 2760 -480 2794
rect -446 2760 -430 2794
rect -500 2724 -430 2760
rect -500 2690 -480 2724
rect -446 2690 -430 2724
rect -500 2654 -430 2690
rect -500 2620 -480 2654
rect -446 2620 -430 2654
rect -500 2584 -430 2620
rect -500 2550 -480 2584
rect -446 2550 -430 2584
rect -500 2514 -430 2550
rect -500 2480 -480 2514
rect -446 2480 -430 2514
rect -500 2444 -430 2480
rect -500 2410 -480 2444
rect -446 2410 -430 2444
rect -500 2374 -430 2410
rect -500 2340 -480 2374
rect -446 2340 -430 2374
rect -500 2310 -430 2340
rect 437 3354 517 3390
rect 437 3320 457 3354
rect 491 3320 517 3354
rect 437 3284 517 3320
rect 437 3250 457 3284
rect 491 3250 517 3284
rect 437 3214 517 3250
rect 437 3180 457 3214
rect 491 3180 517 3214
rect 437 3144 517 3180
rect 437 3110 457 3144
rect 491 3110 517 3144
rect 437 3074 517 3110
rect 437 3040 457 3074
rect 491 3040 517 3074
rect 437 3004 517 3040
rect 437 2970 457 3004
rect 491 2970 517 3004
rect 437 2934 517 2970
rect 437 2900 457 2934
rect 491 2900 517 2934
rect 437 2864 517 2900
rect 437 2830 457 2864
rect 491 2830 517 2864
rect 437 2794 517 2830
rect 437 2760 457 2794
rect 491 2760 517 2794
rect 437 2724 517 2760
rect 437 2690 457 2724
rect 491 2690 517 2724
rect 437 2654 517 2690
rect 437 2620 457 2654
rect 491 2620 517 2654
rect 437 2584 517 2620
rect 437 2550 457 2584
rect 491 2550 517 2584
rect 437 2514 517 2550
rect 437 2480 457 2514
rect 491 2480 517 2514
rect 437 2444 517 2480
rect 437 2410 457 2444
rect 491 2410 517 2444
rect 437 2374 517 2410
rect 437 2340 457 2374
rect 491 2340 517 2374
rect 437 2310 517 2340
rect -500 2290 520 2310
rect -500 2250 -460 2290
rect 480 2250 520 2290
rect -500 2230 520 2250
<< psubdiffcont >>
rect -480 3320 -446 3354
rect -480 3250 -446 3284
rect -480 3180 -446 3214
rect -480 3110 -446 3144
rect -480 3040 -446 3074
rect -480 2970 -446 3004
rect -480 2900 -446 2934
rect -480 2830 -446 2864
rect -480 2760 -446 2794
rect -480 2690 -446 2724
rect -480 2620 -446 2654
rect -480 2550 -446 2584
rect -480 2480 -446 2514
rect -480 2410 -446 2444
rect -480 2340 -446 2374
rect 457 3320 491 3354
rect 457 3250 491 3284
rect 457 3180 491 3214
rect 457 3110 491 3144
rect 457 3040 491 3074
rect 457 2970 491 3004
rect 457 2900 491 2934
rect 457 2830 491 2864
rect 457 2760 491 2794
rect 457 2690 491 2724
rect 457 2620 491 2654
rect 457 2550 491 2584
rect 457 2480 491 2514
rect 457 2410 491 2444
rect 457 2340 491 2374
rect -460 2250 480 2290
<< poly >>
rect -5 3479 17 3483
rect -5 3417 24 3479
rect 2 3413 24 3417
<< polycont >>
rect -316 3429 -282 3463
rect -44 3429 -10 3463
rect 24 3429 58 3463
rect 300 3429 334 3463
<< locali >>
rect -332 3429 -316 3463
rect -282 3429 -44 3463
rect -10 3429 24 3463
rect 58 3429 300 3463
rect 334 3429 361 3463
rect -490 3354 -440 3370
rect -490 3320 -480 3354
rect -446 3320 -440 3354
rect -490 3284 -440 3320
rect -490 3240 -480 3284
rect -446 3240 -440 3284
rect -490 3214 -440 3240
rect -490 3160 -480 3214
rect -446 3160 -440 3214
rect -490 3144 -440 3160
rect -490 3080 -480 3144
rect -446 3080 -440 3144
rect -490 3074 -440 3080
rect -490 3040 -480 3074
rect -446 3040 -440 3074
rect -490 3034 -440 3040
rect -490 2970 -480 3034
rect -446 2970 -440 3034
rect -490 2954 -440 2970
rect -490 2900 -480 2954
rect -446 2900 -440 2954
rect -490 2874 -440 2900
rect -490 2830 -480 2874
rect -446 2830 -440 2874
rect -490 2794 -440 2830
rect -490 2760 -480 2794
rect -446 2760 -440 2794
rect -490 2724 -440 2760
rect -490 2680 -480 2724
rect -446 2680 -440 2724
rect -490 2654 -440 2680
rect -490 2600 -480 2654
rect -446 2600 -440 2654
rect -490 2584 -440 2600
rect -490 2520 -480 2584
rect -446 2520 -440 2584
rect -490 2514 -440 2520
rect -490 2480 -480 2514
rect -446 2480 -440 2514
rect -490 2474 -440 2480
rect -490 2410 -480 2474
rect -446 2410 -440 2474
rect -490 2394 -440 2410
rect -490 2340 -480 2394
rect -446 2340 -440 2394
rect -490 2300 -440 2340
rect 447 3354 507 3370
rect 447 3320 457 3354
rect 491 3320 507 3354
rect 447 3284 507 3320
rect 447 3240 457 3284
rect 491 3240 507 3284
rect 447 3214 507 3240
rect 447 3160 457 3214
rect 491 3160 507 3214
rect 447 3144 507 3160
rect 447 3080 457 3144
rect 491 3080 507 3144
rect 447 3074 507 3080
rect 447 3040 457 3074
rect 491 3040 507 3074
rect 447 3034 507 3040
rect 447 2970 457 3034
rect 491 2970 507 3034
rect 447 2954 507 2970
rect 447 2900 457 2954
rect 491 2900 507 2954
rect 447 2874 507 2900
rect 447 2830 457 2874
rect 491 2830 507 2874
rect 447 2794 507 2830
rect 447 2760 457 2794
rect 491 2760 507 2794
rect 447 2724 507 2760
rect 447 2680 457 2724
rect 491 2680 507 2724
rect 447 2654 507 2680
rect 447 2600 457 2654
rect 491 2600 507 2654
rect 447 2584 507 2600
rect 447 2520 457 2584
rect 491 2520 507 2584
rect 447 2514 507 2520
rect 447 2480 457 2514
rect 491 2480 507 2514
rect 447 2474 507 2480
rect 447 2410 457 2474
rect 491 2410 507 2474
rect 447 2394 507 2410
rect 447 2340 457 2394
rect 491 2340 507 2394
rect 447 2300 507 2340
rect -490 2290 507 2300
rect -490 2250 -460 2290
rect 480 2250 507 2290
rect -490 2240 507 2250
<< viali >>
rect -480 3320 -446 3354
rect -480 3250 -446 3274
rect -480 3240 -446 3250
rect -480 3180 -446 3194
rect -480 3160 -446 3180
rect -480 3110 -446 3114
rect -480 3080 -446 3110
rect -480 3004 -446 3034
rect -480 3000 -446 3004
rect -480 2934 -446 2954
rect -480 2920 -446 2934
rect -480 2864 -446 2874
rect -480 2840 -446 2864
rect -480 2760 -446 2794
rect -480 2690 -446 2714
rect -480 2680 -446 2690
rect -480 2620 -446 2634
rect -480 2600 -446 2620
rect -480 2550 -446 2554
rect -480 2520 -446 2550
rect -480 2444 -446 2474
rect -480 2440 -446 2444
rect -480 2374 -446 2394
rect -480 2360 -446 2374
rect 457 3320 491 3354
rect 457 3250 491 3274
rect 457 3240 491 3250
rect 457 3180 491 3194
rect 457 3160 491 3180
rect 457 3110 491 3114
rect 457 3080 491 3110
rect 457 3004 491 3034
rect 457 3000 491 3004
rect 457 2934 491 2954
rect 457 2920 491 2934
rect 457 2864 491 2874
rect 457 2840 491 2864
rect 457 2760 491 2794
rect 457 2690 491 2714
rect 457 2680 491 2690
rect 457 2620 491 2634
rect 457 2600 491 2620
rect 457 2550 491 2554
rect 457 2520 491 2550
rect 457 2444 491 2474
rect 457 2440 491 2444
rect 457 2374 491 2394
rect 457 2360 491 2374
<< metal1 >>
rect -340 3520 357 3580
rect -5 3417 17 3483
rect -500 3354 -430 3390
rect -500 3320 -480 3354
rect -446 3320 -430 3354
rect -500 3274 -430 3320
rect -500 3240 -480 3274
rect -446 3240 -430 3274
rect -500 3194 -430 3240
rect -500 3160 -480 3194
rect -446 3160 -430 3194
rect -500 3114 -430 3160
rect -500 3080 -480 3114
rect -446 3080 -430 3114
rect -500 3034 -430 3080
rect -500 3000 -480 3034
rect -446 3000 -430 3034
rect -500 2954 -430 3000
rect -500 2920 -480 2954
rect -446 2920 -430 2954
rect -500 2874 -430 2920
rect -500 2840 -480 2874
rect -446 2840 -430 2874
rect -500 2794 -430 2840
rect -500 2760 -480 2794
rect -446 2760 -430 2794
rect -500 2714 -430 2760
rect -500 2680 -480 2714
rect -446 2680 -430 2714
rect -500 2634 -430 2680
rect -500 2600 -480 2634
rect -446 2600 -430 2634
rect -500 2554 -430 2600
rect -500 2520 -480 2554
rect -446 2520 -430 2554
rect -500 2474 -430 2520
rect -500 2440 -480 2474
rect -446 2440 -430 2474
rect -500 2394 -430 2440
rect -500 2360 -480 2394
rect -446 2360 -430 2394
rect -500 2230 -430 2360
rect -363 2310 -310 3380
rect 327 2310 381 3380
rect -360 2300 381 2310
rect -360 2220 -340 2300
rect 360 2230 381 2300
rect 437 3354 507 3390
rect 437 3320 457 3354
rect 491 3320 507 3354
rect 437 3274 507 3320
rect 437 3240 457 3274
rect 491 3240 507 3274
rect 437 3194 507 3240
rect 437 3160 457 3194
rect 491 3160 507 3194
rect 437 3114 507 3160
rect 437 3080 457 3114
rect 491 3080 507 3114
rect 437 3034 507 3080
rect 437 3000 457 3034
rect 491 3000 507 3034
rect 437 2954 507 3000
rect 437 2920 457 2954
rect 491 2920 507 2954
rect 437 2874 507 2920
rect 437 2840 457 2874
rect 491 2840 507 2874
rect 437 2794 507 2840
rect 437 2760 457 2794
rect 491 2760 507 2794
rect 437 2714 507 2760
rect 437 2680 457 2714
rect 491 2680 507 2714
rect 437 2634 507 2680
rect 437 2600 457 2634
rect 491 2600 507 2634
rect 437 2554 507 2600
rect 437 2520 457 2554
rect 491 2520 507 2554
rect 437 2474 507 2520
rect 437 2440 457 2474
rect 491 2440 507 2474
rect 437 2394 507 2440
rect 437 2360 457 2394
rect 491 2360 507 2394
rect 437 2290 507 2360
rect 437 2230 510 2290
rect 360 2220 380 2230
<< via1 >>
rect -340 2220 360 2300
<< metal2 >>
rect -340 3420 377 3500
rect -360 2220 -340 2300
rect 360 2220 380 2300
use sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap  sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0
timestamp 1659107442
transform 1 0 -501 0 1 2289
box 100 -41 576 1290
use sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap  sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_1
timestamp 1659107442
transform 1 0 -157 0 1 2289
box 100 -41 576 1290
<< labels >>
rlabel space -490 2210 -370 2230 1 S
rlabel metal1 -340 3520 -310 3580 1 G
rlabel metal2 -340 3420 -300 3500 1 SD
<< end >>
