** sch_path: /home/al/openmpw/Project-Yatsuhashi-Chip1/xschem/nfet_impedance_test.sch
**.subckt nfet_impedance_test
XM1 vd net1 vs GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
V1 net1 GND 1.8
V2 __UNCONNECTED_PIN__0 GND 0.9
R1 GND vd 0.001 m=1
vsweep vs GND 0
**** begin user architecture code
.lib /home/al/openmpw/pdk_1/sky130B/libs.tech/ngspice/sky130.lib.spice tt
* .include /home/al/openmpw/pdk_1/sky130B/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice



.dc vsweep 0 1.8 0.02
* .ac dec 1000 0.01e9 100e9
.control
run
display
plot abs((v(vs)-v(vd))/@R1[I])
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
