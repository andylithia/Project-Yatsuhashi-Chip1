magic
tech sky130B
magscale 1 2
timestamp 1661649517
<< metal4 >>
rect 13700 8424 17700 8536
rect 13700 4648 13812 8424
rect 17588 4648 17700 8424
tri 12042 1471 13700 3129 se
rect 13700 1471 17700 4648
tri 9100 -1471 12042 1471 se
rect 12042 -1471 13100 1471
rect 9100 -4648 13100 -1471
tri 13100 -3129 17700 1471 nw
rect 9100 -8424 9212 -4648
rect 12988 -8424 13100 -4648
rect 9100 -8536 13100 -8424
<< via4 >>
rect 13812 4648 17588 8424
rect 9212 -8424 12988 -4648
<< metal5 >>
tri -14584 23500 -10584 27500 se
rect -10584 23500 5984 27500
tri 5984 23500 9984 27500 sw
tri -18300 19784 -14584 23500 se
rect -14584 22900 -9527 23500
tri -9527 22900 -8927 23500 nw
tri 4327 22900 4927 23500 ne
rect 4927 22900 9984 23500
rect -14584 22052 -10375 22900
tri -10375 22052 -9527 22900 nw
tri -9527 22052 -8679 22900 se
rect -8679 22052 4079 22900
tri 4079 22052 4927 22900 sw
tri 4927 22052 5775 22900 ne
rect 5775 22052 9984 22900
rect -14584 21204 -11223 22052
tri -11223 21204 -10375 22052 nw
tri -10375 21204 -9527 22052 se
rect -9527 21204 4927 22052
tri 4927 21204 5775 22052 sw
tri 5775 21204 6623 22052 ne
rect 6623 21204 9984 22052
rect -14584 20632 -11795 21204
tri -11795 20632 -11223 21204 nw
tri -10947 20632 -10375 21204 se
rect -10375 20632 5775 21204
tri 5775 20632 6347 21204 sw
tri 6623 20632 7195 21204 ne
rect 7195 20632 9984 21204
rect -14584 19784 -12643 20632
tri -12643 19784 -11795 20632 nw
tri -11795 19784 -10947 20632 se
rect -10947 19784 6347 20632
tri 6347 19784 7195 20632 sw
tri 7195 19784 8043 20632 ne
rect 8043 19784 9984 20632
tri 9984 19784 13700 23500 sw
tri -20241 17843 -18300 19784 se
rect -18300 19748 -12679 19784
tri -12679 19748 -12643 19784 nw
tri -11831 19748 -11795 19784 se
rect -11795 19748 7195 19784
rect -18300 18900 -13527 19748
tri -13527 18900 -12679 19748 nw
tri -12679 18900 -11831 19748 se
rect -11831 18936 7195 19748
tri 7195 18936 8043 19784 sw
tri 8043 18936 8891 19784 ne
rect 8891 18936 13700 19784
rect -11831 18900 8043 18936
tri 8043 18900 8079 18936 sw
tri 8891 18900 8927 18936 ne
rect 8927 18900 13700 18936
rect -18300 18052 -14375 18900
tri -14375 18052 -13527 18900 nw
tri -13527 18052 -12679 18900 se
rect -12679 18052 -8043 18900
rect -18300 17843 -14584 18052
tri -14584 17843 -14375 18052 nw
tri -13736 17843 -13527 18052 se
rect -13527 17879 -8043 18052
tri -8043 17879 -7022 18900 nw
tri 2422 17879 3443 18900 ne
rect 3443 18727 8079 18900
tri 8079 18727 8252 18900 sw
tri 8927 18727 9100 18900 ne
rect 9100 18727 13700 18900
rect 3443 17879 8252 18727
tri 8252 17879 9100 18727 sw
tri 9100 17879 9948 18727 ne
rect 9948 17879 13700 18727
rect -13527 17843 -8079 17879
tri -8079 17843 -8043 17879 nw
tri 3443 17843 3479 17879 ne
rect 3479 17843 9100 17879
tri -22300 15784 -20241 17843 se
rect -20241 16995 -15432 17843
tri -15432 16995 -14584 17843 nw
tri -14584 16995 -13736 17843 se
rect -13736 16995 -11795 17843
rect -20241 16147 -16280 16995
tri -16280 16147 -15432 16995 nw
tri -15432 16147 -14584 16995 se
rect -14584 16147 -11795 16995
rect -20241 15784 -16852 16147
rect -22300 15575 -16852 15784
tri -16852 15575 -16280 16147 nw
tri -16004 15575 -15432 16147 se
rect -15432 15575 -11795 16147
rect -22300 14727 -17700 15575
tri -17700 14727 -16852 15575 nw
tri -16852 14727 -16004 15575 se
rect -16004 14727 -11795 15575
rect -22300 8536 -18300 14727
tri -18300 14127 -17700 14727 nw
tri -17452 14127 -16852 14727 se
rect -16852 14127 -11795 14727
tri -11795 14127 -8079 17843 nw
tri 3479 14127 7195 17843 ne
rect 7195 17031 9100 17843
tri 9100 17031 9948 17879 sw
tri 9948 17031 10796 17879 ne
rect 10796 17031 13700 17879
rect 7195 16183 9948 17031
tri 9948 16183 10796 17031 sw
tri 10796 16183 11644 17031 ne
rect 11644 16183 13700 17031
rect 7195 15575 10796 16183
tri 10796 15575 11404 16183 sw
tri 11644 15575 12252 16183 ne
rect 12252 15784 13700 16183
tri 13700 15784 17700 19784 sw
rect 12252 15575 17700 15784
rect 7195 14727 11404 15575
tri 11404 14727 12252 15575 sw
tri 12252 14727 13100 15575 ne
rect 13100 14727 17700 15575
rect 7195 14127 12252 14727
tri 12252 14127 12852 14727 sw
tri 13100 14127 13700 14727 ne
rect -23322 4536 -18300 8536
tri -17700 13879 -17452 14127 se
rect -17452 13879 -12679 14127
rect -17700 13243 -12679 13879
tri -12679 13243 -11795 14127 nw
tri 7195 13243 8079 14127 ne
rect 8079 13879 12852 14127
tri 12852 13879 13100 14127 sw
rect 8079 13243 13100 13879
rect -23322 -8536 -18300 -4536
rect -22300 -14727 -18300 -8536
rect -17700 -13243 -13700 13243
tri -13700 12222 -12679 13243 nw
tri 8079 12222 9100 13243 ne
rect 9100 1471 13100 13243
rect 13700 8424 17700 14727
rect 13700 4648 13812 8424
rect 17588 4648 17700 8424
rect 13700 4536 17700 4648
tri 9100 -1471 12042 1471 ne
rect 12042 -1471 13100 1471
tri 13100 -1471 17700 3129 sw
tri 12042 -2529 13100 -1471 ne
rect 13100 -2529 17700 -1471
tri 13100 -3129 13700 -2529 ne
rect 9100 -4648 13100 -4536
rect 9100 -8424 9212 -4648
rect 12988 -8424 13100 -4648
tri -13700 -13243 -12679 -12222 sw
tri 8079 -13243 9100 -12222 se
rect 9100 -13243 13100 -8424
rect -17700 -13879 -12679 -13243
tri -17700 -14127 -17452 -13879 ne
rect -17452 -14127 -12679 -13879
tri -12679 -14127 -11795 -13243 sw
tri 7195 -14127 8079 -13243 se
rect 8079 -13879 13100 -13243
rect 8079 -14127 12852 -13879
tri 12852 -14127 13100 -13879 nw
tri -18300 -14727 -17700 -14127 sw
tri -17452 -14727 -16852 -14127 ne
rect -16852 -14727 -11795 -14127
rect -22300 -15575 -17700 -14727
tri -17700 -15575 -16852 -14727 sw
tri -16852 -15575 -16004 -14727 ne
rect -16004 -15575 -11795 -14727
rect -22300 -15784 -16852 -15575
tri -22300 -17843 -20241 -15784 ne
rect -20241 -16147 -16852 -15784
tri -16852 -16147 -16280 -15575 sw
tri -16004 -16147 -15432 -15575 ne
rect -15432 -16147 -11795 -15575
rect -20241 -16995 -16280 -16147
tri -16280 -16995 -15432 -16147 sw
tri -15432 -16995 -14584 -16147 ne
rect -14584 -16995 -11795 -16147
rect -20241 -17843 -15432 -16995
tri -15432 -17843 -14584 -16995 sw
tri -14584 -17843 -13736 -16995 ne
rect -13736 -17843 -11795 -16995
tri -11795 -17843 -8079 -14127 sw
tri 3479 -17843 7195 -14127 se
rect 7195 -14727 12252 -14127
tri 12252 -14727 12852 -14127 nw
tri 13100 -14727 13700 -14127 se
rect 13700 -14727 17700 -2529
rect 7195 -15575 11404 -14727
tri 11404 -15575 12252 -14727 nw
tri 12252 -15575 13100 -14727 se
rect 13100 -15575 17700 -14727
rect 7195 -16183 10796 -15575
tri 10796 -16183 11404 -15575 nw
tri 11644 -16183 12252 -15575 se
rect 12252 -15784 17700 -15575
rect 12252 -16183 13700 -15784
rect 7195 -17031 9948 -16183
tri 9948 -17031 10796 -16183 nw
tri 10796 -17031 11644 -16183 se
rect 11644 -17031 13700 -16183
rect 7195 -17843 9100 -17031
tri -20241 -19784 -18300 -17843 ne
rect -18300 -18052 -14584 -17843
tri -14584 -18052 -14375 -17843 sw
tri -13736 -18052 -13527 -17843 ne
rect -13527 -17879 -8079 -17843
tri -8079 -17879 -8043 -17843 sw
tri 3443 -17879 3479 -17843 se
rect 3479 -17879 9100 -17843
tri 9100 -17879 9948 -17031 nw
tri 9948 -17879 10796 -17031 se
rect 10796 -17879 13700 -17031
rect -13527 -18052 -8043 -17879
rect -18300 -18900 -14375 -18052
tri -14375 -18900 -13527 -18052 sw
tri -13527 -18900 -12679 -18052 ne
rect -12679 -18900 -8043 -18052
tri -8043 -18900 -7022 -17879 sw
tri 2422 -18900 3443 -17879 se
rect 3443 -18727 8252 -17879
tri 8252 -18727 9100 -17879 nw
tri 9100 -18727 9948 -17879 se
rect 9948 -18727 13700 -17879
rect 3443 -18900 8079 -18727
tri 8079 -18900 8252 -18727 nw
tri 8927 -18900 9100 -18727 se
rect 9100 -18900 13700 -18727
rect -18300 -19748 -13527 -18900
tri -13527 -19748 -12679 -18900 sw
tri -12679 -19748 -11831 -18900 ne
rect -11831 -18936 8043 -18900
tri 8043 -18936 8079 -18900 nw
tri 8891 -18936 8927 -18900 se
rect 8927 -18936 13700 -18900
rect -11831 -19748 7195 -18936
rect -18300 -19784 -12679 -19748
tri -12679 -19784 -12643 -19748 sw
tri -11831 -19784 -11795 -19748 ne
rect -11795 -19784 7195 -19748
tri 7195 -19784 8043 -18936 nw
tri 8043 -19784 8891 -18936 se
rect 8891 -19784 13700 -18936
tri 13700 -19784 17700 -15784 nw
tri -18300 -23500 -14584 -19784 ne
rect -14584 -20632 -12643 -19784
tri -12643 -20632 -11795 -19784 sw
tri -11795 -20632 -10947 -19784 ne
rect -10947 -20632 6347 -19784
tri 6347 -20632 7195 -19784 nw
tri 7195 -20632 8043 -19784 se
rect 8043 -20632 9984 -19784
rect -14584 -21204 -11795 -20632
tri -11795 -21204 -11223 -20632 sw
tri -10947 -21204 -10375 -20632 ne
rect -10375 -21204 5775 -20632
tri 5775 -21204 6347 -20632 nw
tri 6623 -21204 7195 -20632 se
rect 7195 -21204 9984 -20632
rect -14584 -22052 -11223 -21204
tri -11223 -22052 -10375 -21204 sw
tri -10375 -22052 -9527 -21204 ne
rect -9527 -22052 4927 -21204
tri 4927 -22052 5775 -21204 nw
tri 5775 -22052 6623 -21204 se
rect 6623 -22052 9984 -21204
rect -14584 -22900 -10375 -22052
tri -10375 -22900 -9527 -22052 sw
tri -9527 -22900 -8679 -22052 ne
rect -8679 -22900 4079 -22052
tri 4079 -22900 4927 -22052 nw
tri 4927 -22900 5775 -22052 se
rect 5775 -22900 9984 -22052
rect -14584 -23500 -9527 -22900
tri -9527 -23500 -8927 -22900 sw
tri 4327 -23500 4927 -22900 se
rect 4927 -23500 9984 -22900
tri 9984 -23500 13700 -19784 nw
tri -14584 -27500 -10584 -23500 ne
rect -10584 -27500 5984 -23500
tri 5984 -27500 9984 -23500 nw
<< end >>
