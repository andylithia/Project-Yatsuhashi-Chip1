magic
tech sky130A
magscale 1 2
timestamp 1665269856
<< metal4 >>
rect -77600 -27112 -53600 -27000
rect -77600 -33888 -60488 -27112
rect -53712 -33888 -53600 -27112
rect -77600 -34000 -53600 -33888
<< via4 >>
rect -60488 -33888 -53712 -27112
<< metal5 >>
tri -57962 25500 -50962 32500 se
rect -50962 25500 2962 32500
tri 2962 25500 9962 32500 sw
tri -61400 22062 -57962 25500 se
rect -57962 24700 -48862 25500
tri -48862 24700 -48062 25500 nw
tri 62 24700 862 25500 ne
rect 862 24700 9962 25500
rect -57962 23569 -49993 24700
tri -49993 23569 -48862 24700 nw
tri -48862 23569 -47731 24700 se
rect -47731 23569 -269 24700
tri -269 23569 862 24700 sw
tri 862 23569 1993 24700 ne
rect 1993 23569 9962 24700
rect -57962 23193 -50369 23569
tri -50369 23193 -49993 23569 nw
tri -49238 23193 -48862 23569 se
rect -48862 23193 862 23569
rect -57962 22062 -51500 23193
tri -51500 22062 -50369 23193 nw
tri -50369 22062 -49238 23193 se
rect -49238 22438 862 23193
tri 862 22438 1993 23569 sw
tri 1993 22438 3124 23569 ne
rect 3124 22438 9962 23569
rect -49238 22062 1993 22438
tri -69200 14262 -61400 22062 se
rect -61400 20931 -52631 22062
tri -52631 20931 -51500 22062 nw
tri -51500 20931 -50369 22062 se
rect -50369 21307 1993 22062
tri 1993 21307 3124 22438 sw
tri 3124 21307 4255 22438 ne
rect 4255 21307 9962 22438
rect -50369 20931 3124 21307
tri 3124 20931 3500 21307 sw
tri 4255 20931 4631 21307 ne
rect 4631 20931 9962 21307
rect -61400 19800 -53762 20931
tri -53762 19800 -52631 20931 nw
tri -52631 19800 -51500 20931 se
rect -51500 19962 3500 20931
tri 3500 19962 4469 20931 sw
tri 4631 19962 5600 20931 ne
rect 5600 19962 9962 20931
rect -51500 19800 4469 19962
rect -61400 18831 -54731 19800
tri -54731 18831 -53762 19800 nw
tri -53600 18831 -52631 19800 se
rect -52631 18831 4469 19800
tri 4469 18831 5600 19962 sw
tri 5600 18831 6731 19962 ne
rect 6731 18831 9962 19962
rect -61400 17700 -55862 18831
tri -55862 17700 -54731 18831 nw
tri -54731 17700 -53600 18831 se
rect -53600 17700 5600 18831
tri 5600 17700 6731 18831 sw
tri 6731 17700 7862 18831 ne
rect 7862 17700 9962 18831
tri 9962 17700 17762 25500 sw
rect -61400 16569 -56993 17700
tri -56993 16569 -55862 17700 nw
tri -55862 16569 -54731 17700 se
rect -54731 16900 -45631 17700
tri -45631 16900 -44831 17700 nw
tri -3169 16900 -2369 17700 ne
rect -2369 16900 6731 17700
rect -54731 16569 -46762 16900
rect -61400 15438 -58124 16569
tri -58124 15438 -56993 16569 nw
tri -56993 15438 -55862 16569 se
rect -55862 15769 -46762 16569
tri -46762 15769 -45631 16900 nw
tri -45631 15769 -44500 16900 se
rect -44500 15769 -3500 16900
tri -3500 15769 -2369 16900 sw
tri -2369 15769 -1238 16900 ne
rect -1238 16569 6731 16900
tri 6731 16569 7862 17700 sw
tri 7862 16569 8993 17700 ne
rect 8993 16569 17762 17700
rect -1238 15769 7862 16569
rect -55862 15438 -47893 15769
rect -61400 14424 -59138 15438
tri -59138 14424 -58124 15438 nw
tri -58007 14424 -56993 15438 se
rect -56993 14638 -47893 15438
tri -47893 14638 -46762 15769 nw
tri -46762 14638 -45631 15769 se
rect -45631 14638 -2369 15769
tri -2369 14638 -1238 15769 sw
tri -1238 14638 -107 15769 ne
rect -107 15438 7862 15769
tri 7862 15438 8993 16569 sw
tri 8993 15438 10124 16569 ne
rect 10124 15438 17762 16569
rect -107 14638 8993 15438
rect -56993 14424 -49024 14638
rect -61400 14262 -60269 14424
tri -71300 12162 -69200 14262 se
rect -69200 13293 -60269 14262
tri -60269 13293 -59138 14424 nw
tri -59138 13293 -58007 14424 se
rect -58007 13507 -49024 14424
tri -49024 13507 -47893 14638 nw
tri -47893 13507 -46762 14638 se
rect -46762 13507 -1238 14638
tri -1238 13507 -107 14638 sw
tri -107 13507 1024 14638 ne
rect 1024 14307 8993 14638
tri 8993 14307 10124 15438 sw
tri 10124 14307 11255 15438 ne
rect 11255 14307 17762 15438
rect 1024 13507 10124 14307
rect -58007 13293 -49238 13507
tri -49238 13293 -49024 13507 nw
tri -48107 13293 -47893 13507 se
rect -47893 13293 -107 13507
tri -107 13293 107 13507 sw
tri 1024 13293 1238 13507 ne
rect 1238 13293 10124 13507
tri 10124 13293 11138 14307 sw
tri 11255 13293 12269 14307 ne
rect 12269 13293 17762 14307
rect -69200 12162 -61400 13293
tri -61400 12162 -60269 13293 nw
tri -60269 12162 -59138 13293 se
rect -59138 12162 -50369 13293
tri -50369 12162 -49238 13293 nw
tri -49238 12162 -48107 13293 se
rect -48107 12162 107 13293
tri 107 12162 1238 13293 sw
tri 1238 12162 2369 13293 ne
rect 2369 12162 11138 13293
tri 11138 12162 12269 13293 sw
tri 12269 12162 13400 13293 ne
rect 13400 12162 17762 13293
tri -77000 6462 -71300 12162 se
rect -71300 11031 -62531 12162
tri -62531 11031 -61400 12162 nw
tri -61400 11031 -60269 12162 se
rect -60269 11031 -51500 12162
tri -51500 11031 -50369 12162 nw
tri -50369 11031 -49238 12162 se
rect -49238 11031 1238 12162
tri 1238 11031 2369 12162 sw
tri 2369 11031 3500 12162 ne
rect 3500 11031 12269 12162
tri 12269 11031 13400 12162 sw
tri 13400 11031 14531 12162 ne
rect 14531 11031 17762 12162
rect -71300 9900 -63662 11031
tri -63662 9900 -62531 11031 nw
tri -62531 9900 -61400 11031 se
rect -61400 9900 -52631 11031
tri -52631 9900 -51500 11031 nw
tri -51500 9900 -50369 11031 se
rect -50369 9900 2369 11031
tri 2369 9900 3500 11031 sw
tri 3500 9900 4631 11031 ne
rect 4631 9900 13400 11031
tri 13400 9900 14531 11031 sw
tri 14531 9900 15662 11031 ne
rect 15662 9900 17762 11031
tri 17762 9900 25562 17700 sw
rect -71300 8769 -64793 9900
tri -64793 8769 -63662 9900 nw
tri -63662 8769 -62531 9900 se
rect -62531 8769 -53762 9900
tri -53762 8769 -52631 9900 nw
tri -52631 8769 -51500 9900 se
rect -71300 7638 -65924 8769
tri -65924 7638 -64793 8769 nw
tri -64793 7638 -63662 8769 se
rect -63662 7638 -54893 8769
tri -54893 7638 -53762 8769 nw
tri -53762 7638 -52631 8769 se
rect -52631 7638 -51500 8769
rect -71300 6624 -66938 7638
tri -66938 6624 -65924 7638 nw
tri -65807 6624 -64793 7638 se
rect -64793 6624 -56024 7638
rect -71300 6462 -68069 6624
tri -79100 4362 -77000 6462 se
rect -77000 5493 -68069 6462
tri -68069 5493 -66938 6624 nw
tri -66938 5493 -65807 6624 se
rect -65807 6507 -56024 6624
tri -56024 6507 -54893 7638 nw
tri -54893 6507 -53762 7638 se
rect -53762 6507 -51500 7638
rect -65807 5493 -57155 6507
rect -77000 4362 -69200 5493
tri -69200 4362 -68069 5493 nw
tri -68069 4362 -66938 5493 se
rect -66938 5376 -57155 5493
tri -57155 5376 -56024 6507 nw
tri -56024 5376 -54893 6507 se
rect -54893 5376 -51500 6507
rect -66938 4524 -58007 5376
tri -58007 4524 -57155 5376 nw
tri -56876 4524 -56024 5376 se
rect -56024 4524 -51500 5376
rect -66938 4362 -59138 4524
tri -84000 -538 -79100 4362 se
rect -79100 3231 -70331 4362
tri -70331 3231 -69200 4362 nw
tri -69200 3231 -68069 4362 se
rect -68069 3393 -59138 4362
tri -59138 3393 -58007 4524 nw
tri -58007 3393 -56876 4524 se
rect -56876 3393 -51500 4524
rect -68069 3231 -60269 3393
rect -79100 2100 -71462 3231
tri -71462 2100 -70331 3231 nw
tri -70331 2100 -69200 3231 se
rect -69200 2262 -60269 3231
tri -60269 2262 -59138 3393 nw
tri -59138 2262 -58007 3393 se
rect -58007 2262 -51500 3393
rect -69200 2100 -61400 2262
rect -79100 1131 -72431 2100
tri -72431 1131 -71462 2100 nw
tri -71300 1131 -70331 2100 se
rect -70331 1131 -61400 2100
tri -61400 1131 -60269 2262 nw
tri -60269 1131 -59138 2262 se
rect -59138 1131 -51500 2262
rect -79100 0 -73562 1131
tri -73562 0 -72431 1131 nw
tri -72431 0 -71300 1131 se
rect -71300 0 -62531 1131
tri -62531 0 -61400 1131 nw
tri -61400 0 -60269 1131 se
rect -60269 0 -51500 1131
tri -51500 0 -41600 9900 nw
tri -6400 0 3500 9900 ne
tri 3500 8769 4631 9900 sw
tri 4631 8769 5762 9900 ne
rect 5762 8769 14531 9900
tri 14531 8769 15662 9900 sw
tri 15662 8769 16793 9900 ne
rect 16793 8769 25562 9900
rect 3500 7638 4631 8769
tri 4631 7638 5762 8769 sw
tri 5762 7638 6893 8769 ne
rect 6893 7638 15662 8769
tri 15662 7638 16793 8769 sw
tri 16793 7638 17924 8769 ne
rect 17924 7638 25562 8769
rect 3500 6507 5762 7638
tri 5762 6507 6893 7638 sw
tri 6893 6507 8024 7638 ne
rect 8024 6507 16793 7638
tri 16793 6507 17924 7638 sw
tri 17924 6507 19055 7638 ne
rect 19055 6507 25562 7638
rect 3500 5376 6893 6507
tri 6893 5376 8024 6507 sw
tri 8024 5376 9155 6507 ne
rect 9155 5376 17924 6507
tri 17924 5376 19055 6507 sw
tri 19055 5376 20186 6507 ne
rect 20186 5376 25562 6507
rect 3500 4524 8024 5376
tri 8024 4524 8876 5376 sw
tri 9155 4524 10007 5376 ne
rect 10007 4524 19055 5376
tri 19055 4524 19907 5376 sw
tri 20186 4524 21038 5376 ne
rect 21038 4524 25562 5376
rect 3500 3393 8876 4524
tri 8876 3393 10007 4524 sw
tri 10007 3393 11138 4524 ne
rect 11138 3393 19907 4524
tri 19907 3393 21038 4524 sw
tri 21038 3393 22169 4524 ne
rect 22169 3393 25562 4524
rect 3500 2262 10007 3393
tri 10007 2262 11138 3393 sw
tri 11138 2262 12269 3393 ne
rect 12269 2262 21038 3393
tri 21038 2262 22169 3393 sw
tri 22169 2262 23300 3393 ne
rect 23300 2262 25562 3393
rect 3500 1131 11138 2262
tri 11138 1131 12269 2262 sw
tri 12269 1131 13400 2262 ne
rect 13400 1131 22169 2262
tri 22169 1131 23300 2262 sw
tri 23300 1131 24431 2262 ne
rect 24431 1131 25562 2262
rect 3500 0 12269 1131
tri 12269 0 13400 1131 sw
tri 13400 0 14531 1131 ne
rect 14531 0 23300 1131
tri 23300 0 24431 1131 sw
tri 24431 0 25562 1131 ne
tri 25562 0 35462 9900 sw
rect -79100 -538 -74693 0
rect -84000 -1131 -74693 -538
tri -74693 -1131 -73562 0 nw
tri -73562 -1131 -72431 0 se
rect -72431 -1131 -63662 0
tri -63662 -1131 -62531 0 nw
tri -62531 -1131 -61400 0 se
rect -84000 -1507 -75069 -1131
tri -75069 -1507 -74693 -1131 nw
tri -73938 -1507 -73562 -1131 se
rect -73562 -1507 -64793 -1131
rect -84000 -2638 -76200 -1507
tri -76200 -2638 -75069 -1507 nw
tri -75069 -2638 -73938 -1507 se
rect -73938 -2262 -64793 -1507
tri -64793 -2262 -63662 -1131 nw
tri -63662 -2262 -62531 -1131 se
rect -62531 -2262 -61400 -1131
rect -73938 -2638 -65924 -2262
rect -84000 -13000 -77000 -2638
tri -77000 -3438 -76200 -2638 nw
tri -75869 -3438 -75069 -2638 se
rect -75069 -3393 -65924 -2638
tri -65924 -3393 -64793 -2262 nw
tri -64793 -3393 -63662 -2262 se
rect -63662 -3393 -61400 -2262
rect -75069 -3438 -66138 -3393
tri -76200 -3769 -75869 -3438 se
rect -75869 -3607 -66138 -3438
tri -66138 -3607 -65924 -3393 nw
tri -65007 -3607 -64793 -3393 se
rect -64793 -3607 -61400 -3393
rect -75869 -3769 -67269 -3607
rect -76200 -4738 -67269 -3769
tri -67269 -4738 -66138 -3607 nw
tri -66138 -4738 -65007 -3607 se
rect -65007 -4738 -61400 -3607
rect -76200 -5869 -68400 -4738
tri -68400 -5869 -67269 -4738 nw
tri -67269 -5869 -66138 -4738 se
rect -66138 -5869 -61400 -4738
rect -76200 -39647 -69200 -5869
tri -69200 -6669 -68400 -5869 nw
tri -68400 -7000 -67269 -5869 se
rect -67269 -7000 -61400 -5869
rect -68400 -36416 -61400 -7000
tri -61400 -9900 -51500 0 nw
tri 3500 -9900 13400 0 ne
tri 13400 -1131 14531 0 sw
tri 14531 -1131 15662 0 ne
rect 15662 -1131 24431 0
tri 24431 -1131 25562 0 sw
tri 25562 -1131 26693 0 ne
rect 26693 -538 35462 0
tri 35462 -538 36000 0 sw
rect 26693 -1131 36000 -538
rect 13400 -2262 14531 -1131
tri 14531 -2262 15662 -1131 sw
tri 15662 -2262 16793 -1131 ne
rect 16793 -1507 25562 -1131
tri 25562 -1507 25938 -1131 sw
tri 26693 -1507 27069 -1131 ne
rect 27069 -1507 36000 -1131
rect 16793 -2262 25938 -1507
rect 13400 -3393 15662 -2262
tri 15662 -3393 16793 -2262 sw
tri 16793 -3393 17924 -2262 ne
rect 17924 -2638 25938 -2262
tri 25938 -2638 27069 -1507 sw
tri 27069 -2638 28200 -1507 ne
rect 28200 -2638 36000 -1507
rect 17924 -3393 27069 -2638
rect 13400 -3607 16793 -3393
tri 16793 -3607 17007 -3393 sw
tri 17924 -3607 18138 -3393 ne
rect 18138 -3607 27069 -3393
rect 13400 -4738 17007 -3607
tri 17007 -4738 18138 -3607 sw
tri 18138 -4738 19269 -3607 ne
rect 19269 -3769 27069 -3607
tri 27069 -3769 28200 -2638 sw
tri 28200 -3438 29000 -2638 ne
rect 19269 -4738 28200 -3769
rect 13400 -5869 18138 -4738
tri 18138 -5869 19269 -4738 sw
tri 19269 -5869 20400 -4738 ne
rect 20400 -5869 28200 -4738
rect 13400 -7000 19269 -5869
tri 19269 -7000 20400 -5869 sw
tri 20400 -6669 21200 -5869 ne
rect -60600 -27112 -53600 -27000
rect -60600 -33888 -60488 -27112
rect -53712 -33888 -53600 -27112
rect -60600 -35284 -53600 -33888
tri -61400 -36416 -60600 -35616 sw
tri -60600 -36416 -59468 -35284 ne
rect -59468 -36416 -53600 -35284
rect -68400 -37548 -60600 -36416
tri -60600 -37548 -59468 -36416 sw
tri -59468 -37548 -58336 -36416 ne
rect -58336 -37548 -53600 -36416
rect -68400 -38515 -59468 -37548
tri -69200 -39647 -68400 -38847 sw
tri -68400 -39647 -67268 -38515 ne
rect -67268 -38680 -59468 -38515
tri -59468 -38680 -58336 -37548 sw
tri -58336 -38680 -57204 -37548 ne
rect -57204 -38680 -53600 -37548
rect -67268 -38888 -58336 -38680
tri -58336 -38888 -58128 -38680 sw
tri -57204 -38888 -56996 -38680 ne
rect -56996 -38888 -53600 -38680
rect -67268 -39647 -58128 -38888
rect -76200 -40779 -68400 -39647
tri -68400 -40779 -67268 -39647 sw
tri -67268 -40779 -66136 -39647 ne
rect -66136 -40020 -58128 -39647
tri -58128 -40020 -56996 -38888 sw
tri -56996 -40020 -55864 -38888 ne
rect -55864 -40020 -53600 -38888
rect -66136 -40779 -56996 -40020
rect -76200 -41152 -67268 -40779
tri -67268 -41152 -66895 -40779 sw
tri -66136 -41152 -65763 -40779 ne
rect -65763 -41152 -56996 -40779
tri -56996 -41152 -55864 -40020 sw
tri -55864 -41152 -54732 -40020 ne
rect -54732 -41152 -53600 -40020
rect -76200 -41746 -66895 -41152
tri -76200 -49900 -68046 -41746 ne
rect -68046 -42284 -66895 -41746
tri -66895 -42284 -65763 -41152 sw
tri -65763 -42284 -64631 -41152 ne
rect -64631 -42284 -55864 -41152
tri -55864 -42284 -54732 -41152 sw
tri -54732 -42284 -53600 -41152 ne
tri -53600 -42284 -43701 -32385 sw
tri 5784 -40001 13400 -32385 se
rect 13400 -35284 20400 -7000
rect 13400 -36416 19268 -35284
tri 19268 -36416 20400 -35284 nw
tri 20400 -36416 21200 -35616 se
rect 21200 -36416 28200 -5869
rect 13400 -37548 18136 -36416
tri 18136 -37548 19268 -36416 nw
tri 19268 -37548 20400 -36416 se
rect 20400 -37548 28200 -36416
rect 13400 -37737 17947 -37548
tri 17947 -37737 18136 -37548 nw
tri 19079 -37737 19268 -37548 se
rect 19268 -37737 28200 -37548
rect 13400 -38869 16815 -37737
tri 16815 -38869 17947 -37737 nw
tri 17947 -38869 19079 -37737 se
rect 19079 -38515 28200 -37737
rect 19079 -38869 27068 -38515
rect 13400 -40001 15683 -38869
tri 15683 -40001 16815 -38869 nw
tri 16815 -40001 17947 -38869 se
rect 17947 -39647 27068 -38869
tri 27068 -39647 28200 -38515 nw
tri 28200 -39647 29000 -38847 se
rect 29000 -39647 36000 -2638
rect 17947 -40001 25936 -39647
tri 3501 -42284 5784 -40001 se
rect 5784 -41133 14551 -40001
tri 14551 -41133 15683 -40001 nw
tri 15683 -41133 16815 -40001 se
rect 16815 -40779 25936 -40001
tri 25936 -40779 27068 -39647 nw
tri 27068 -40779 28200 -39647 se
rect 28200 -40779 36000 -39647
rect 16815 -41133 25563 -40779
rect 5784 -41152 14532 -41133
tri 14532 -41152 14551 -41133 nw
tri 15664 -41152 15683 -41133 se
rect 15683 -41152 25563 -41133
tri 25563 -41152 25936 -40779 nw
tri 26695 -41152 27068 -40779 se
rect 27068 -41152 36000 -40779
rect 5784 -42284 13400 -41152
tri 13400 -42284 14532 -41152 nw
tri 14532 -42284 15664 -41152 se
rect 15664 -42284 24431 -41152
tri 24431 -42284 25563 -41152 nw
tri 25563 -42284 26695 -41152 se
rect 26695 -41746 36000 -41152
rect 26695 -42284 29000 -41746
rect -68046 -43416 -65763 -42284
tri -65763 -43416 -64631 -42284 sw
tri -64631 -43416 -63499 -42284 ne
rect -63499 -43416 -54732 -42284
tri -54732 -43416 -53600 -42284 sw
tri -53600 -43416 -52468 -42284 ne
rect -52468 -43416 -43701 -42284
rect -68046 -44548 -64631 -43416
tri -64631 -44548 -63499 -43416 sw
tri -63499 -44548 -62367 -43416 ne
rect -62367 -44548 -53600 -43416
tri -53600 -44548 -52468 -43416 sw
tri -52468 -44548 -51336 -43416 ne
rect -51336 -44548 -43701 -43416
rect -68046 -45680 -63499 -44548
tri -63499 -45680 -62367 -44548 sw
tri -62367 -45680 -61235 -44548 ne
rect -61235 -45680 -52468 -44548
tri -52468 -45680 -51336 -44548 sw
tri -51336 -45680 -50204 -44548 ne
rect -50204 -45680 -43701 -44548
rect -68046 -46504 -62367 -45680
tri -62367 -46504 -61543 -45680 sw
tri -61235 -46504 -60411 -45680 ne
rect -60411 -46504 -51336 -45680
tri -51336 -46504 -50512 -45680 sw
tri -50204 -46504 -49380 -45680 ne
rect -49380 -46504 -43701 -45680
rect -68046 -47636 -61543 -46504
tri -61543 -47636 -60411 -46504 sw
tri -60411 -47636 -59279 -46504 ne
rect -59279 -47636 -50512 -46504
tri -50512 -47636 -49380 -46504 sw
tri -49380 -47636 -48248 -46504 ne
rect -48248 -47636 -43701 -46504
rect -68046 -48768 -60411 -47636
tri -60411 -48768 -59279 -47636 sw
tri -59279 -48768 -58147 -47636 ne
rect -58147 -48768 -49380 -47636
tri -49380 -48768 -48248 -47636 sw
tri -48248 -48768 -47116 -47636 ne
rect -47116 -48768 -43701 -47636
rect -68046 -49900 -59279 -48768
tri -59279 -49900 -58147 -48768 sw
tri -58147 -49900 -57015 -48768 ne
rect -57015 -49900 -48248 -48768
tri -48248 -49900 -47116 -48768 sw
tri -47116 -49900 -45984 -48768 ne
rect -45984 -49900 -43701 -48768
tri -43701 -49900 -36085 -42284 sw
tri -4115 -49900 3501 -42284 se
rect 3501 -43416 12268 -42284
tri 12268 -43416 13400 -42284 nw
tri 13400 -43416 14532 -42284 se
rect 14532 -43416 23299 -42284
tri 23299 -43416 24431 -42284 nw
tri 24431 -43416 25563 -42284 se
rect 25563 -43416 29000 -42284
rect 3501 -44548 11136 -43416
tri 11136 -44548 12268 -43416 nw
tri 12268 -44548 13400 -43416 se
rect 13400 -44383 22332 -43416
tri 22332 -44383 23299 -43416 nw
tri 23464 -44383 24431 -43416 se
rect 24431 -44383 29000 -43416
rect 13400 -44548 21200 -44383
rect 3501 -45680 10004 -44548
tri 10004 -45680 11136 -44548 nw
tri 11136 -45680 12268 -44548 se
rect 12268 -45515 21200 -44548
tri 21200 -45515 22332 -44383 nw
tri 22332 -45515 23464 -44383 se
rect 23464 -45515 29000 -44383
rect 12268 -45680 20068 -45515
rect 3501 -46504 9180 -45680
tri 9180 -46504 10004 -45680 nw
tri 10312 -46504 11136 -45680 se
rect 11136 -46504 20068 -45680
rect 3501 -47636 8048 -46504
tri 8048 -47636 9180 -46504 nw
tri 9180 -47636 10312 -46504 se
rect 10312 -46647 20068 -46504
tri 20068 -46647 21200 -45515 nw
tri 21200 -46647 22332 -45515 se
rect 22332 -46647 29000 -45515
rect 10312 -47636 18936 -46647
rect 3501 -48768 6916 -47636
tri 6916 -48768 8048 -47636 nw
tri 8048 -48768 9180 -47636 se
rect 9180 -47779 18936 -47636
tri 18936 -47779 20068 -46647 nw
tri 20068 -47779 21200 -46647 se
rect 21200 -47779 29000 -46647
rect 9180 -48768 17947 -47779
tri 17947 -48768 18936 -47779 nw
tri 19079 -48768 20068 -47779 se
rect 20068 -48746 29000 -47779
tri 29000 -48746 36000 -41746 nw
rect 20068 -48768 21200 -48746
rect 3501 -49900 5784 -48768
tri 5784 -49900 6916 -48768 nw
tri 6916 -49900 8048 -48768 se
rect 8048 -49900 16815 -48768
tri 16815 -49900 17947 -48768 nw
tri 17947 -49900 19079 -48768 se
rect 19079 -49900 21200 -48768
tri -68046 -57700 -60246 -49900 ne
rect -60246 -51032 -58147 -49900
tri -58147 -51032 -57015 -49900 sw
tri -57015 -51032 -55883 -49900 ne
rect -55883 -51032 -47116 -49900
tri -47116 -51032 -45984 -49900 sw
tri -45984 -51032 -44852 -49900 ne
rect -44852 -51032 4652 -49900
tri 4652 -51032 5784 -49900 nw
tri 5784 -51032 6916 -49900 se
rect 6916 -51032 15683 -49900
tri 15683 -51032 16815 -49900 nw
tri 16815 -51032 17947 -49900 se
rect 17947 -51032 21200 -49900
rect -60246 -52164 -57015 -51032
tri -57015 -52164 -55883 -51032 sw
tri -55883 -52164 -54751 -51032 ne
rect -54751 -52164 -45984 -51032
tri -45984 -52164 -44852 -51032 sw
tri -44852 -52164 -43720 -51032 ne
rect -43720 -52164 3520 -51032
tri 3520 -52164 4652 -51032 nw
tri 4652 -52164 5784 -51032 se
rect 5784 -52164 14551 -51032
tri 14551 -52164 15683 -51032 nw
tri 15683 -52164 16815 -51032 se
rect 16815 -52164 21200 -51032
rect -60246 -53296 -55883 -52164
tri -55883 -53296 -54751 -52164 sw
tri -54751 -53296 -53619 -52164 ne
rect -53619 -53296 -44852 -52164
tri -44852 -53296 -43720 -52164 sw
tri -43720 -53296 -42588 -52164 ne
rect -42588 -53296 2388 -52164
tri 2388 -53296 3520 -52164 nw
tri 3520 -53296 4652 -52164 se
rect 4652 -52183 14532 -52164
tri 14532 -52183 14551 -52164 nw
tri 15664 -52183 15683 -52164 se
rect 15683 -52183 21200 -52164
rect 4652 -53296 13400 -52183
rect -60246 -54304 -54751 -53296
tri -54751 -54304 -53743 -53296 sw
tri -53619 -54304 -52611 -53296 ne
rect -52611 -53504 -43720 -53296
tri -43720 -53504 -43512 -53296 sw
tri -42588 -53504 -42380 -53296 ne
rect -42380 -53504 2180 -53296
tri 2180 -53504 2388 -53296 nw
tri 3312 -53504 3520 -53296 se
rect 3520 -53315 13400 -53296
tri 13400 -53315 14532 -52183 nw
tri 14532 -53315 15664 -52183 se
rect 15664 -53315 21200 -52183
rect 3520 -53504 12268 -53315
rect -52611 -54304 -43512 -53504
rect -60246 -55436 -53743 -54304
tri -53743 -55436 -52611 -54304 sw
tri -52611 -55436 -51479 -54304 ne
rect -51479 -54636 -43512 -54304
tri -43512 -54636 -42380 -53504 sw
tri -42380 -54636 -41248 -53504 ne
rect -41248 -54636 1048 -53504
tri 1048 -54636 2180 -53504 nw
tri 2180 -54636 3312 -53504 se
rect 3312 -54447 12268 -53504
tri 12268 -54447 13400 -53315 nw
tri 13400 -54447 14532 -53315 se
rect 14532 -54447 21200 -53315
rect 3312 -54636 11136 -54447
rect -51479 -55436 -42380 -54636
rect -60246 -56568 -52611 -55436
tri -52611 -56568 -51479 -55436 sw
tri -51479 -56568 -50347 -55436 ne
rect -50347 -55768 -42380 -55436
tri -42380 -55768 -41248 -54636 sw
tri -41248 -55768 -40116 -54636 ne
rect -40116 -55768 -84 -54636
tri -84 -55768 1048 -54636 nw
tri 1048 -55768 2180 -54636 se
rect 2180 -55579 11136 -54636
tri 11136 -55579 12268 -54447 nw
tri 12268 -55579 13400 -54447 se
rect 13400 -55579 21200 -54447
rect 2180 -55768 10147 -55579
rect -50347 -56568 -41248 -55768
rect -60246 -57700 -51479 -56568
tri -51479 -57700 -50347 -56568 sw
tri -50347 -57700 -49215 -56568 ne
rect -49215 -56900 -41248 -56568
tri -41248 -56900 -40116 -55768 sw
tri -40116 -56900 -38984 -55768 ne
rect -38984 -56900 -1216 -55768
tri -1216 -56900 -84 -55768 nw
tri -84 -56900 1048 -55768 se
rect 1048 -56568 10147 -55768
tri 10147 -56568 11136 -55579 nw
tri 11279 -56568 12268 -55579 se
rect 12268 -56546 21200 -55579
tri 21200 -56546 29000 -48746 nw
rect 12268 -56568 13400 -56546
rect 1048 -56900 9015 -56568
rect -49215 -57700 -40116 -56900
tri -40116 -57700 -39316 -56900 sw
tri -884 -57700 -84 -56900 se
rect -84 -57700 9015 -56900
tri 9015 -57700 10147 -56568 nw
tri 10147 -57700 11279 -56568 se
rect 11279 -57700 13400 -56568
tri -60246 -65500 -52446 -57700 ne
rect -52446 -58832 -50347 -57700
tri -50347 -58832 -49215 -57700 sw
tri -49215 -58832 -48083 -57700 ne
rect -48083 -58832 7883 -57700
tri 7883 -58832 9015 -57700 nw
tri 9015 -58832 10147 -57700 se
rect 10147 -58832 13400 -57700
rect -52446 -59964 -49215 -58832
tri -49215 -59964 -48083 -58832 sw
tri -48083 -59964 -46951 -58832 ne
rect -46951 -59799 6916 -58832
tri 6916 -59799 7883 -58832 nw
tri 8048 -59799 9015 -58832 se
rect 9015 -59799 13400 -58832
rect -46951 -59964 5784 -59799
rect -52446 -61096 -48083 -59964
tri -48083 -61096 -46951 -59964 sw
tri -46951 -61096 -45819 -59964 ne
rect -45819 -60931 5784 -59964
tri 5784 -60931 6916 -59799 nw
tri 6916 -60931 8048 -59799 se
rect 8048 -60931 13400 -59799
rect -45819 -61096 4652 -60931
rect -52446 -61304 -46951 -61096
tri -46951 -61304 -46743 -61096 sw
tri -45819 -61304 -45611 -61096 ne
rect -45611 -61304 4652 -61096
rect -52446 -62436 -46743 -61304
tri -46743 -62436 -45611 -61304 sw
tri -45611 -62436 -44479 -61304 ne
rect -44479 -62063 4652 -61304
tri 4652 -62063 5784 -60931 nw
tri 5784 -62063 6916 -60931 se
rect 6916 -62063 13400 -60931
rect -44479 -62436 3520 -62063
rect -52446 -63568 -45611 -62436
tri -45611 -63568 -44479 -62436 sw
tri -44479 -63568 -43347 -62436 ne
rect -43347 -63195 3520 -62436
tri 3520 -63195 4652 -62063 nw
tri 4652 -63195 5784 -62063 se
rect 5784 -63195 13400 -62063
rect -43347 -63568 3147 -63195
tri 3147 -63568 3520 -63195 nw
tri 4279 -63568 4652 -63195 se
rect 4652 -63568 13400 -63195
rect -52446 -64700 -44479 -63568
tri -44479 -64700 -43347 -63568 sw
tri -43347 -64700 -42215 -63568 ne
rect -42215 -64700 2015 -63568
tri 2015 -64700 3147 -63568 nw
tri 3147 -64700 4279 -63568 se
rect 4279 -64346 13400 -63568
tri 13400 -64346 21200 -56546 nw
rect 4279 -64700 5246 -64346
rect -52446 -65500 -43347 -64700
tri -43347 -65500 -42547 -64700 sw
tri 2347 -65500 3147 -64700 se
rect 3147 -65500 5246 -64700
tri -52446 -72500 -45446 -65500 ne
rect -45446 -72500 5246 -65500
tri 5246 -72500 13400 -64346 nw
<< end >>
