magic
tech sky130A
magscale 1 2
timestamp 1664327021
<< metal2 >>
rect 6500 6100 7800 6500
rect 12800 6100 14100 6500
rect 19100 6100 20400 6500
rect 6500 5500 7800 5900
rect 12800 5500 14100 5900
rect 19100 5500 20400 5900
rect 6500 4900 7800 5300
rect 12800 4900 14100 5300
rect 19100 4900 20400 5300
rect 6500 4300 7800 4700
rect 12800 4300 14100 4700
rect 19100 4300 20400 4700
rect 6500 3700 7800 4100
rect 12800 3700 14100 4100
rect 19100 3700 20400 4100
rect 6500 3100 7800 3500
rect 12800 3100 14100 3500
rect 19100 3100 20400 3500
rect 6500 2500 7800 2900
rect 12800 2500 14100 2900
rect 19100 2500 20400 2900
rect 6500 1900 7800 2300
rect 12800 1900 14100 2300
rect 19100 1900 20400 2300
rect 6500 1300 7800 1700
rect 12800 1300 14100 1700
rect 19100 1300 20400 1700
rect 6500 700 7800 1100
rect 12800 700 14100 1100
rect 19100 700 20400 1100
rect 6500 100 7800 500
rect 12800 100 14100 500
rect 19100 100 20400 500
rect 6900 -500 7400 100
rect 13200 -500 13700 100
rect 19500 -500 20000 100
rect 6500 -900 7800 -500
rect 12800 -900 14100 -500
rect 19100 -900 20400 -500
rect 6500 -1500 7800 -1100
rect 12800 -1500 14100 -1100
rect 19100 -1500 20400 -1100
rect 6500 -2100 7800 -1700
rect 12800 -2100 14100 -1700
rect 19100 -2100 20400 -1700
rect 6500 -2700 7800 -2300
rect 12800 -2700 14100 -2300
rect 19100 -2700 20400 -2300
rect 6500 -3300 7800 -2900
rect 12800 -3300 14100 -2900
rect 19100 -3300 20400 -2900
rect 6500 -3900 7800 -3500
rect 12800 -3900 14100 -3500
rect 19100 -3900 20400 -3500
rect 6500 -4500 7800 -4100
rect 12800 -4500 14100 -4100
rect 19100 -4500 20400 -4100
rect 6500 -5100 7800 -4700
rect 12800 -5100 14100 -4700
rect 19100 -5100 20400 -4700
rect 6500 -5700 7800 -5300
rect 12800 -5700 14100 -5300
rect 19100 -5700 20400 -5300
rect 6500 -6300 7800 -5900
rect 12800 -6300 14100 -5900
rect 19100 -6300 20400 -5900
rect 6500 -6900 7800 -6500
rect 12800 -6900 14100 -6500
rect 19100 -6900 20400 -6500
<< metal3 >>
rect 1560 6560 6380 6589
rect 1560 6220 1620 6560
rect 5020 6220 6380 6560
rect 1560 6189 6380 6220
rect 7860 6560 12680 6589
rect 7860 6220 7880 6560
rect 9260 6220 12680 6560
rect 7860 6189 12680 6220
rect 1560 1100 6380 1140
rect 1560 780 1700 1100
rect 4900 780 6380 1100
rect 1560 740 6380 780
rect 7860 1100 12680 1140
rect 7860 780 11440 1100
rect 12660 780 12680 1100
rect 7860 740 12680 780
rect 3100 400 5000 500
rect 3100 300 3300 400
rect 1400 100 3300 300
rect 4800 300 5000 400
rect 7800 300 12800 500
rect 14100 400 19100 500
rect 14100 300 15900 400
rect 4800 180 7400 300
rect 4800 100 7020 180
rect 1400 20 7020 100
rect 7380 20 7400 180
rect 1400 0 7400 20
rect 7600 180 13700 300
rect 7600 20 13320 180
rect 13680 20 13700 180
rect 7600 0 13700 20
rect 13900 100 15900 300
rect 17400 300 19100 400
rect 20400 300 25400 500
rect 17400 180 20000 300
rect 17400 100 19620 180
rect 13900 20 19620 100
rect 19980 20 20000 180
rect 13900 0 20000 20
rect 20200 0 25400 300
rect 7600 -200 7900 0
rect 9400 -100 12000 0
rect 13900 -100 14100 0
rect 20200 -100 20500 0
rect 22000 -100 24600 0
rect 6500 -400 7900 -200
rect 12800 -300 14100 -100
rect 19100 -300 20500 -100
rect 3100 -500 5000 -400
rect 6500 -500 6800 -400
rect 9400 -500 12000 -400
rect 12800 -500 13100 -300
rect 15700 -500 17600 -400
rect 19100 -500 19400 -300
rect 22000 -500 24600 -400
rect 1400 -800 3300 -500
rect 4800 -800 6800 -500
rect 7000 -520 13100 -500
rect 7000 -680 7020 -520
rect 7380 -680 13100 -520
rect 7000 -800 13100 -680
rect 13300 -520 15900 -500
rect 13300 -680 13320 -520
rect 13680 -680 15900 -520
rect 13300 -800 15900 -680
rect 17400 -800 19400 -500
rect 19600 -520 25400 -500
rect 19600 -680 19620 -520
rect 19980 -680 25400 -520
rect 19600 -800 25400 -680
rect 3100 -900 5000 -800
rect 15700 -900 17600 -800
rect 1560 -1060 6380 -1011
rect 1560 -1360 3260 -1060
rect 4840 -1360 6380 -1060
rect 1560 -1411 6380 -1360
rect 7860 -1040 12680 -1011
rect 7860 -1380 7900 -1040
rect 9260 -1380 12680 -1040
rect 7860 -1411 12680 -1380
rect 1560 -6500 6380 -6460
rect 1560 -6820 5140 -6500
rect 6360 -6820 6380 -6500
rect 1560 -6860 6380 -6820
rect 7860 -6480 12680 -6460
rect 7860 -6840 9640 -6480
rect 11060 -6840 12680 -6480
rect 7860 -6860 12680 -6840
<< via3 >>
rect 1620 6220 5020 6560
rect 7880 6220 9260 6560
rect 14220 6220 17620 6560
rect 20480 6220 21860 6560
rect 1700 780 4900 1100
rect 11440 780 12660 1100
rect 14300 780 17500 1100
rect 24040 780 25260 1100
rect 3300 100 4800 400
rect 7020 20 7380 180
rect 13320 20 13680 180
rect 15900 100 17400 400
rect 19620 20 19980 180
rect 3300 -800 4800 -500
rect 7020 -680 7380 -520
rect 13320 -680 13680 -520
rect 15900 -800 17400 -500
rect 19620 -680 19980 -520
rect 3260 -1360 4840 -1060
rect 7900 -1380 9260 -1040
rect 15860 -1360 17440 -1060
rect 20500 -1380 21860 -1040
rect 5140 -6820 6360 -6500
rect 9640 -6840 11060 -6480
rect 17740 -6820 18960 -6500
rect 22240 -6840 23660 -6480
<< metal4 >>
rect 5200 11100 6700 11200
rect 5200 9500 5300 11100
rect 6600 9500 6700 11100
rect 1400 8000 2900 8200
rect 1400 6600 1600 8000
rect 2800 6600 2900 8000
rect 1400 6560 5100 6600
rect 1400 6220 1620 6560
rect 5020 6220 5100 6560
rect 1400 6180 5100 6220
rect 1400 1100 5000 1140
rect 1400 780 1700 1100
rect 4900 780 5000 1100
rect 1400 700 5000 780
rect 1400 -9900 2900 700
rect 3200 400 4900 500
rect 3200 100 3300 400
rect 4800 100 4900 400
rect 3200 0 4900 100
rect 3200 -500 4900 -400
rect 3200 -800 3300 -500
rect 4800 -800 4900 -500
rect 3200 -900 4900 -800
rect 3220 -1060 4880 -1020
rect 3220 -1360 3260 -1060
rect 4840 -1360 4880 -1060
rect 3220 -1400 4880 -1360
rect 3300 -6900 4800 -1400
rect 5200 -6460 6700 9500
rect 7700 11100 9200 11200
rect 7700 9500 7800 11100
rect 9100 9500 9200 11100
rect 7700 6600 9200 9500
rect 17800 11100 19300 11200
rect 17800 9500 17900 11100
rect 19200 9500 19300 11100
rect 9600 8100 11100 8200
rect 7700 6560 9300 6600
rect 7700 6220 7880 6560
rect 9260 6220 9300 6560
rect 7700 6180 9300 6220
rect 9600 6500 9800 8100
rect 11000 6500 11100 8100
rect 7000 180 7400 200
rect 7000 20 7020 180
rect 7380 20 7400 180
rect 7000 -520 7400 20
rect 7000 -680 7020 -520
rect 7380 -680 7400 -520
rect 7000 -700 7400 -680
rect 5100 -6500 6700 -6460
rect 5100 -6820 5140 -6500
rect 6360 -6820 6700 -6500
rect 5100 -6860 6700 -6820
rect 7700 -1040 9300 -1000
rect 7700 -1380 7900 -1040
rect 9260 -1380 9300 -1040
rect 7700 -1420 9300 -1380
rect 3300 -8500 3400 -6900
rect 4700 -8500 4800 -6900
rect 3300 -8600 4800 -8500
rect 1400 -11500 1500 -9900
rect 2800 -11500 2900 -9900
rect 1400 -11600 2900 -11500
rect 7700 -9900 9200 -1420
rect 9600 -6480 11100 6500
rect 14000 8000 15500 8200
rect 14000 6600 14200 8000
rect 15400 6600 15500 8000
rect 14000 6560 17700 6600
rect 14000 6220 14220 6560
rect 17620 6220 17700 6560
rect 14000 6180 17700 6220
rect 14000 6080 15500 6180
rect 11400 1100 13000 1140
rect 11400 780 11440 1100
rect 12660 780 13000 1100
rect 11400 740 13000 780
rect 9600 -6840 9640 -6480
rect 11060 -6840 11100 -6480
rect 9600 -6860 11100 -6840
rect 11500 -6900 13000 740
rect 14000 1100 17600 1140
rect 14000 780 14300 1100
rect 17500 780 17600 1100
rect 14000 700 17600 780
rect 13300 180 13700 200
rect 13300 20 13320 180
rect 13680 20 13700 180
rect 13300 -520 13700 20
rect 13300 -680 13320 -520
rect 13680 -680 13700 -520
rect 13300 -700 13700 -680
rect 11500 -8500 11600 -6900
rect 12900 -8500 13000 -6900
rect 11500 -8600 13000 -8500
rect 7700 -11500 7800 -9900
rect 9100 -11500 9200 -9900
rect 7700 -11600 9200 -11500
rect 14000 -9900 15500 700
rect 15800 400 17500 500
rect 15800 100 15900 400
rect 17400 100 17500 400
rect 15800 0 17500 100
rect 15800 -500 17500 -400
rect 15800 -800 15900 -500
rect 17400 -800 17500 -500
rect 15800 -900 17500 -800
rect 15820 -1060 17480 -1020
rect 15820 -1360 15860 -1060
rect 17440 -1360 17480 -1060
rect 15820 -1400 17480 -1360
rect 15900 -6900 17400 -1400
rect 17800 -6460 19300 9500
rect 20300 11100 21800 11200
rect 20300 9500 20400 11100
rect 21700 9500 21800 11100
rect 20300 8200 21800 9500
rect 20300 6560 21900 8200
rect 20300 6220 20480 6560
rect 21860 6220 21900 6560
rect 20300 6180 21900 6220
rect 22200 8100 23700 8200
rect 22200 6500 22400 8100
rect 23600 6500 23700 8100
rect 20300 6040 21800 6180
rect 19600 180 20000 200
rect 19600 20 19620 180
rect 19980 20 20000 180
rect 19600 -520 20000 20
rect 19600 -680 19620 -520
rect 19980 -680 20000 -520
rect 19600 -700 20000 -680
rect 17700 -6500 19300 -6460
rect 17700 -6820 17740 -6500
rect 18960 -6820 19300 -6500
rect 17700 -6860 19300 -6820
rect 20300 -1040 21900 -1000
rect 20300 -1380 20500 -1040
rect 21860 -1380 21900 -1040
rect 20300 -1420 21900 -1380
rect 15900 -8500 16000 -6900
rect 17300 -8500 17400 -6900
rect 15900 -8600 17400 -8500
rect 14000 -11500 14100 -9900
rect 15400 -11500 15500 -9900
rect 14000 -11600 15500 -11500
rect 20300 -9900 21800 -1420
rect 22200 -6480 23700 6500
rect 24000 1100 25340 1140
rect 24000 780 24040 1100
rect 25260 780 25340 1100
rect 24000 740 25340 780
rect 22200 -6840 22240 -6480
rect 23660 -6840 23700 -6480
rect 22200 -6860 23700 -6840
rect 24100 700 25340 740
rect 24100 -6900 25600 700
rect 24100 -8500 24200 -6900
rect 25500 -8500 25600 -6900
rect 24100 -8600 25600 -8500
rect 20300 -11500 20400 -9900
rect 21700 -11500 21800 -9900
rect 20300 -11600 21800 -11500
<< via4 >>
rect 5300 9500 6600 11100
rect 1600 6600 2800 8000
rect 3300 100 4800 400
rect 3300 -800 4800 -500
rect 7800 9500 9100 11100
rect 17900 9500 19200 11100
rect 9800 6500 11000 8100
rect 3400 -8500 4700 -6900
rect 1500 -11500 2800 -9900
rect 14200 6600 15400 8000
rect 11600 -8500 12900 -6900
rect 7800 -11500 9100 -9900
rect 15900 100 17400 400
rect 15900 -800 17400 -500
rect 20400 9500 21700 11100
rect 22400 6500 23600 8100
rect 16000 -8500 17300 -6900
rect 14100 -11500 15400 -9900
rect 24200 -8500 25500 -6900
rect 20400 -11500 21700 -9900
<< metal5 >>
rect 1400 8200 4200 11400
rect 22800 11200 25600 11400
rect 5200 11100 25600 11200
rect 5200 9500 5300 11100
rect 6600 9500 7800 11100
rect 9100 9500 17900 11100
rect 19200 9500 20400 11100
rect 21700 9500 25600 11100
rect 5200 9400 25600 9500
rect 1400 8100 23700 8200
rect 1400 8000 9800 8100
rect 1400 6600 1600 8000
rect 2800 6600 9800 8000
rect 1400 6500 9800 6600
rect 11000 8000 22400 8100
rect 11000 6600 14200 8000
rect 15400 6600 22400 8000
rect 11000 6500 22400 6600
rect 23600 6500 23700 8100
rect 1400 6400 23700 6500
rect 1300 400 25500 500
rect 1300 100 3300 400
rect 4800 100 15900 400
rect 17400 100 25500 400
rect 1300 0 25500 100
rect 1300 -500 25500 -400
rect 1300 -800 3300 -500
rect 4800 -800 15900 -500
rect 17400 -800 25500 -500
rect 1300 -900 25500 -800
rect 3300 -6900 25600 -6800
rect 3300 -8500 3400 -6900
rect 4700 -8500 11600 -6900
rect 12900 -8500 16000 -6900
rect 17300 -8500 24200 -6900
rect 25500 -8500 25600 -6900
rect 3300 -8600 25600 -8500
rect 1400 -9900 21800 -9800
rect 1400 -11500 1500 -9900
rect 2800 -11500 7800 -9900
rect 9100 -11500 14100 -9900
rect 15400 -11500 20400 -9900
rect 21700 -11500 21800 -9900
rect 1400 -11600 21800 -11500
rect 1400 -11800 4200 -11600
rect 22800 -11800 25600 -8600
use ./CLASSE/NMOS_30_0p5_30_3  NMOS_30_0p5_30_1_0 ./CLASSE
timestamp 1664325575
transform 1 0 1400 0 1 400
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_3  NMOS_30_0p5_30_1_1
timestamp 1664325575
transform 1 0 7700 0 1 400
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_3  NMOS_30_0p5_30_1_2
timestamp 1664325575
transform 1 0 14000 0 1 400
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_3  NMOS_30_0p5_30_1_3
timestamp 1664325575
transform 1 0 20300 0 1 400
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_3  NMOS_30_0p5_30_1_4
timestamp 1664325575
transform 1 0 20300 0 1 -7200
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_3  NMOS_30_0p5_30_1_5
timestamp 1664325575
transform 1 0 14000 0 1 -7200
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_3  NMOS_30_0p5_30_1_6
timestamp 1664325575
transform 1 0 7700 0 1 -7200
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_3  NMOS_30_0p5_30_1_7
timestamp 1664325575
transform 1 0 1400 0 1 -7200
box 0 0 5138 6516
<< labels >>
rlabel metal5 1300 0 1400 500 1 GL
rlabel metal5 1300 -900 1400 -400 1 GR
rlabel metal5 1400 -11800 4200 -11600 1 SD2L
rlabel metal5 22800 -11800 25600 -11600 1 SD2R
rlabel metal5 22800 11200 25600 11400 1 SD1R
rlabel metal5 1400 11200 4200 11400 1 SD1L
rlabel metal2 13300 1400 13600 1500 1 SUB
<< end >>
