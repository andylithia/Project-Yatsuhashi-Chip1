** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/LNA5_with_output_buf.sch
**.subckt LNA5_with_output_buf
V1 VDD GND 1.8
V2 net10 GND dc 0.9 ac 1 portnum 1 z0 50
Ldeg3 net1 GNDI 0.6n m=1
C2 vgate1 net1 100f m=1
R1 net8 net15 1k m=1
Ldeg1 vgate1 net2 0.5n m=1
I0 GNDI vbias1 0.5m
Ldeg2 VDDI net3 3n m=1
XM5 n_ds1 vgate1 net1 GNDI sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=6
XM1 vbias1 vbias1 GNDI GNDI sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=1
XM2 net3 VDDI n_ds1 GNDI sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=6
XC7 vbias1 GNDI sky130_fd_pr__cap_mim_m3_1 W=20 L=30 MF=1 m=1
Ldeg5 net4 VDDI 2n m=1
R3 net4 VDD 3 m=1
Ldeg6 net5 GND 2n m=1
R4 net5 GNDI 3 m=1
XM12 net6 net9 net16 GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=3
V4 net14 GND DC 0.9 AC 0 portnum 2 z0 50
L1 net11 GND 1n m=1
C17 net14 net6 200f m=1
L2 net7 net6 1.4n m=1
C12 __UNCONNECTED_PIN__0 net3 80f m=1
XC3 net17 GNDI sky130_fd_pr__cap_mim_m3_1 W=20 L=120 MF=1 m=1
C8 GNDI GND 200f m=1
C19 VDD VDDI 200f m=1
R2 net17 VDDI 5 m=1
C5 net8 __UNCONNECTED_PIN__1 1n m=1
C4 VDDI net3 150f m=1
Ldeg4 net2 net8 1n m=1
Ldeg7 vbias1 net15 1n m=1
Ldeg8 net9 net13 3n m=1
R5 net13 net12 2k m=1
V3 net7 GND 0.9
XM4 net16 net9 net11 GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=3
V5 net12 GND 1.2
C1 net13 net10 1n m=1
C6 net6 net7 500f m=1
R6 net13 net6 1k m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice



.subckt sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=2.828e+12p pd=2.132e+07u as=4.242e+12p
+ ps=3.198e+07u w=5.05e+06u l=150000u
X1 SOURCE SUBSTRATE SUBSTRATE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.03e+12p
+ ps=2.14e+07u w=5.05e+06u l=150000u
X2 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X5 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends
.sp dec 1000 0.1e9 10e9 1
* .ac dec 1000 0.01e9 100e9
.control
run
display
let z11=50*(1+s_1_1)/(1-s_1_1)
let z22=50*(1+s_2_2)/(1-s_2_2)
let S11 = S_1_1
let S21 = S_2_1
let S12 = S_1_2
let S22 = S_2_2

* Stability
let delta=S11*S22-S12*S21
let K    = (1-mag(S11)^2-mag(S22)^2+mag(delta)^2)/(2*mag(S12*S21))
let mu   = (1-mag(S11)^2)/(mag(S22-conj(S11)*delta)+mag(S21*S12))
* plot real(z11) real(z22)
* plot imag(z11) imag(z22)
plot db(S_1_1) db(S_2_2) db(S_2_1)

plot K
plot mag(delta)
plot mu
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL GNDI
.end
