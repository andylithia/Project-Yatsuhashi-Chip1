magic
tech sky130B
magscale 1 2
timestamp 1662234432
<< nwell >>
rect -4811 -684 4811 684
<< pmos >>
rect -4615 -464 -4415 536
rect -4357 -464 -4157 536
rect -4099 -464 -3899 536
rect -3841 -464 -3641 536
rect -3583 -464 -3383 536
rect -3325 -464 -3125 536
rect -3067 -464 -2867 536
rect -2809 -464 -2609 536
rect -2551 -464 -2351 536
rect -2293 -464 -2093 536
rect -2035 -464 -1835 536
rect -1777 -464 -1577 536
rect -1519 -464 -1319 536
rect -1261 -464 -1061 536
rect -1003 -464 -803 536
rect -745 -464 -545 536
rect -487 -464 -287 536
rect -229 -464 -29 536
rect 29 -464 229 536
rect 287 -464 487 536
rect 545 -464 745 536
rect 803 -464 1003 536
rect 1061 -464 1261 536
rect 1319 -464 1519 536
rect 1577 -464 1777 536
rect 1835 -464 2035 536
rect 2093 -464 2293 536
rect 2351 -464 2551 536
rect 2609 -464 2809 536
rect 2867 -464 3067 536
rect 3125 -464 3325 536
rect 3383 -464 3583 536
rect 3641 -464 3841 536
rect 3899 -464 4099 536
rect 4157 -464 4357 536
rect 4415 -464 4615 536
<< pdiff >>
rect -4673 524 -4615 536
rect -4673 -452 -4661 524
rect -4627 -452 -4615 524
rect -4673 -464 -4615 -452
rect -4415 524 -4357 536
rect -4415 -452 -4403 524
rect -4369 -452 -4357 524
rect -4415 -464 -4357 -452
rect -4157 524 -4099 536
rect -4157 -452 -4145 524
rect -4111 -452 -4099 524
rect -4157 -464 -4099 -452
rect -3899 524 -3841 536
rect -3899 -452 -3887 524
rect -3853 -452 -3841 524
rect -3899 -464 -3841 -452
rect -3641 524 -3583 536
rect -3641 -452 -3629 524
rect -3595 -452 -3583 524
rect -3641 -464 -3583 -452
rect -3383 524 -3325 536
rect -3383 -452 -3371 524
rect -3337 -452 -3325 524
rect -3383 -464 -3325 -452
rect -3125 524 -3067 536
rect -3125 -452 -3113 524
rect -3079 -452 -3067 524
rect -3125 -464 -3067 -452
rect -2867 524 -2809 536
rect -2867 -452 -2855 524
rect -2821 -452 -2809 524
rect -2867 -464 -2809 -452
rect -2609 524 -2551 536
rect -2609 -452 -2597 524
rect -2563 -452 -2551 524
rect -2609 -464 -2551 -452
rect -2351 524 -2293 536
rect -2351 -452 -2339 524
rect -2305 -452 -2293 524
rect -2351 -464 -2293 -452
rect -2093 524 -2035 536
rect -2093 -452 -2081 524
rect -2047 -452 -2035 524
rect -2093 -464 -2035 -452
rect -1835 524 -1777 536
rect -1835 -452 -1823 524
rect -1789 -452 -1777 524
rect -1835 -464 -1777 -452
rect -1577 524 -1519 536
rect -1577 -452 -1565 524
rect -1531 -452 -1519 524
rect -1577 -464 -1519 -452
rect -1319 524 -1261 536
rect -1319 -452 -1307 524
rect -1273 -452 -1261 524
rect -1319 -464 -1261 -452
rect -1061 524 -1003 536
rect -1061 -452 -1049 524
rect -1015 -452 -1003 524
rect -1061 -464 -1003 -452
rect -803 524 -745 536
rect -803 -452 -791 524
rect -757 -452 -745 524
rect -803 -464 -745 -452
rect -545 524 -487 536
rect -545 -452 -533 524
rect -499 -452 -487 524
rect -545 -464 -487 -452
rect -287 524 -229 536
rect -287 -452 -275 524
rect -241 -452 -229 524
rect -287 -464 -229 -452
rect -29 524 29 536
rect -29 -452 -17 524
rect 17 -452 29 524
rect -29 -464 29 -452
rect 229 524 287 536
rect 229 -452 241 524
rect 275 -452 287 524
rect 229 -464 287 -452
rect 487 524 545 536
rect 487 -452 499 524
rect 533 -452 545 524
rect 487 -464 545 -452
rect 745 524 803 536
rect 745 -452 757 524
rect 791 -452 803 524
rect 745 -464 803 -452
rect 1003 524 1061 536
rect 1003 -452 1015 524
rect 1049 -452 1061 524
rect 1003 -464 1061 -452
rect 1261 524 1319 536
rect 1261 -452 1273 524
rect 1307 -452 1319 524
rect 1261 -464 1319 -452
rect 1519 524 1577 536
rect 1519 -452 1531 524
rect 1565 -452 1577 524
rect 1519 -464 1577 -452
rect 1777 524 1835 536
rect 1777 -452 1789 524
rect 1823 -452 1835 524
rect 1777 -464 1835 -452
rect 2035 524 2093 536
rect 2035 -452 2047 524
rect 2081 -452 2093 524
rect 2035 -464 2093 -452
rect 2293 524 2351 536
rect 2293 -452 2305 524
rect 2339 -452 2351 524
rect 2293 -464 2351 -452
rect 2551 524 2609 536
rect 2551 -452 2563 524
rect 2597 -452 2609 524
rect 2551 -464 2609 -452
rect 2809 524 2867 536
rect 2809 -452 2821 524
rect 2855 -452 2867 524
rect 2809 -464 2867 -452
rect 3067 524 3125 536
rect 3067 -452 3079 524
rect 3113 -452 3125 524
rect 3067 -464 3125 -452
rect 3325 524 3383 536
rect 3325 -452 3337 524
rect 3371 -452 3383 524
rect 3325 -464 3383 -452
rect 3583 524 3641 536
rect 3583 -452 3595 524
rect 3629 -452 3641 524
rect 3583 -464 3641 -452
rect 3841 524 3899 536
rect 3841 -452 3853 524
rect 3887 -452 3899 524
rect 3841 -464 3899 -452
rect 4099 524 4157 536
rect 4099 -452 4111 524
rect 4145 -452 4157 524
rect 4099 -464 4157 -452
rect 4357 524 4415 536
rect 4357 -452 4369 524
rect 4403 -452 4415 524
rect 4357 -464 4415 -452
rect 4615 524 4673 536
rect 4615 -452 4627 524
rect 4661 -452 4673 524
rect 4615 -464 4673 -452
<< pdiffc >>
rect -4661 -452 -4627 524
rect -4403 -452 -4369 524
rect -4145 -452 -4111 524
rect -3887 -452 -3853 524
rect -3629 -452 -3595 524
rect -3371 -452 -3337 524
rect -3113 -452 -3079 524
rect -2855 -452 -2821 524
rect -2597 -452 -2563 524
rect -2339 -452 -2305 524
rect -2081 -452 -2047 524
rect -1823 -452 -1789 524
rect -1565 -452 -1531 524
rect -1307 -452 -1273 524
rect -1049 -452 -1015 524
rect -791 -452 -757 524
rect -533 -452 -499 524
rect -275 -452 -241 524
rect -17 -452 17 524
rect 241 -452 275 524
rect 499 -452 533 524
rect 757 -452 791 524
rect 1015 -452 1049 524
rect 1273 -452 1307 524
rect 1531 -452 1565 524
rect 1789 -452 1823 524
rect 2047 -452 2081 524
rect 2305 -452 2339 524
rect 2563 -452 2597 524
rect 2821 -452 2855 524
rect 3079 -452 3113 524
rect 3337 -452 3371 524
rect 3595 -452 3629 524
rect 3853 -452 3887 524
rect 4111 -452 4145 524
rect 4369 -452 4403 524
rect 4627 -452 4661 524
<< nsubdiff >>
rect -4775 614 -4679 648
rect 4679 614 4775 648
rect -4775 551 -4741 614
rect 4741 551 4775 614
rect -4775 -614 -4741 -551
rect 4741 -614 4775 -551
rect -4775 -648 -4679 -614
rect 4679 -648 4775 -614
<< nsubdiffcont >>
rect -4679 614 4679 648
rect -4775 -551 -4741 551
rect 4741 -551 4775 551
rect -4679 -648 4679 -614
<< poly >>
rect -4615 536 -4415 562
rect -4357 536 -4157 562
rect -4099 536 -3899 562
rect -3841 536 -3641 562
rect -3583 536 -3383 562
rect -3325 536 -3125 562
rect -3067 536 -2867 562
rect -2809 536 -2609 562
rect -2551 536 -2351 562
rect -2293 536 -2093 562
rect -2035 536 -1835 562
rect -1777 536 -1577 562
rect -1519 536 -1319 562
rect -1261 536 -1061 562
rect -1003 536 -803 562
rect -745 536 -545 562
rect -487 536 -287 562
rect -229 536 -29 562
rect 29 536 229 562
rect 287 536 487 562
rect 545 536 745 562
rect 803 536 1003 562
rect 1061 536 1261 562
rect 1319 536 1519 562
rect 1577 536 1777 562
rect 1835 536 2035 562
rect 2093 536 2293 562
rect 2351 536 2551 562
rect 2609 536 2809 562
rect 2867 536 3067 562
rect 3125 536 3325 562
rect 3383 536 3583 562
rect 3641 536 3841 562
rect 3899 536 4099 562
rect 4157 536 4357 562
rect 4415 536 4615 562
rect -4615 -511 -4415 -464
rect -4615 -545 -4599 -511
rect -4431 -545 -4415 -511
rect -4615 -561 -4415 -545
rect -4357 -511 -4157 -464
rect -4357 -545 -4341 -511
rect -4173 -545 -4157 -511
rect -4357 -561 -4157 -545
rect -4099 -511 -3899 -464
rect -4099 -545 -4083 -511
rect -3915 -545 -3899 -511
rect -4099 -561 -3899 -545
rect -3841 -511 -3641 -464
rect -3841 -545 -3825 -511
rect -3657 -545 -3641 -511
rect -3841 -561 -3641 -545
rect -3583 -511 -3383 -464
rect -3583 -545 -3567 -511
rect -3399 -545 -3383 -511
rect -3583 -561 -3383 -545
rect -3325 -511 -3125 -464
rect -3325 -545 -3309 -511
rect -3141 -545 -3125 -511
rect -3325 -561 -3125 -545
rect -3067 -511 -2867 -464
rect -3067 -545 -3051 -511
rect -2883 -545 -2867 -511
rect -3067 -561 -2867 -545
rect -2809 -511 -2609 -464
rect -2809 -545 -2793 -511
rect -2625 -545 -2609 -511
rect -2809 -561 -2609 -545
rect -2551 -511 -2351 -464
rect -2551 -545 -2535 -511
rect -2367 -545 -2351 -511
rect -2551 -561 -2351 -545
rect -2293 -511 -2093 -464
rect -2293 -545 -2277 -511
rect -2109 -545 -2093 -511
rect -2293 -561 -2093 -545
rect -2035 -511 -1835 -464
rect -2035 -545 -2019 -511
rect -1851 -545 -1835 -511
rect -2035 -561 -1835 -545
rect -1777 -511 -1577 -464
rect -1777 -545 -1761 -511
rect -1593 -545 -1577 -511
rect -1777 -561 -1577 -545
rect -1519 -511 -1319 -464
rect -1519 -545 -1503 -511
rect -1335 -545 -1319 -511
rect -1519 -561 -1319 -545
rect -1261 -511 -1061 -464
rect -1261 -545 -1245 -511
rect -1077 -545 -1061 -511
rect -1261 -561 -1061 -545
rect -1003 -511 -803 -464
rect -1003 -545 -987 -511
rect -819 -545 -803 -511
rect -1003 -561 -803 -545
rect -745 -511 -545 -464
rect -745 -545 -729 -511
rect -561 -545 -545 -511
rect -745 -561 -545 -545
rect -487 -511 -287 -464
rect -487 -545 -471 -511
rect -303 -545 -287 -511
rect -487 -561 -287 -545
rect -229 -511 -29 -464
rect -229 -545 -213 -511
rect -45 -545 -29 -511
rect -229 -561 -29 -545
rect 29 -511 229 -464
rect 29 -545 45 -511
rect 213 -545 229 -511
rect 29 -561 229 -545
rect 287 -511 487 -464
rect 287 -545 303 -511
rect 471 -545 487 -511
rect 287 -561 487 -545
rect 545 -511 745 -464
rect 545 -545 561 -511
rect 729 -545 745 -511
rect 545 -561 745 -545
rect 803 -511 1003 -464
rect 803 -545 819 -511
rect 987 -545 1003 -511
rect 803 -561 1003 -545
rect 1061 -511 1261 -464
rect 1061 -545 1077 -511
rect 1245 -545 1261 -511
rect 1061 -561 1261 -545
rect 1319 -511 1519 -464
rect 1319 -545 1335 -511
rect 1503 -545 1519 -511
rect 1319 -561 1519 -545
rect 1577 -511 1777 -464
rect 1577 -545 1593 -511
rect 1761 -545 1777 -511
rect 1577 -561 1777 -545
rect 1835 -511 2035 -464
rect 1835 -545 1851 -511
rect 2019 -545 2035 -511
rect 1835 -561 2035 -545
rect 2093 -511 2293 -464
rect 2093 -545 2109 -511
rect 2277 -545 2293 -511
rect 2093 -561 2293 -545
rect 2351 -511 2551 -464
rect 2351 -545 2367 -511
rect 2535 -545 2551 -511
rect 2351 -561 2551 -545
rect 2609 -511 2809 -464
rect 2609 -545 2625 -511
rect 2793 -545 2809 -511
rect 2609 -561 2809 -545
rect 2867 -511 3067 -464
rect 2867 -545 2883 -511
rect 3051 -545 3067 -511
rect 2867 -561 3067 -545
rect 3125 -511 3325 -464
rect 3125 -545 3141 -511
rect 3309 -545 3325 -511
rect 3125 -561 3325 -545
rect 3383 -511 3583 -464
rect 3383 -545 3399 -511
rect 3567 -545 3583 -511
rect 3383 -561 3583 -545
rect 3641 -511 3841 -464
rect 3641 -545 3657 -511
rect 3825 -545 3841 -511
rect 3641 -561 3841 -545
rect 3899 -511 4099 -464
rect 3899 -545 3915 -511
rect 4083 -545 4099 -511
rect 3899 -561 4099 -545
rect 4157 -511 4357 -464
rect 4157 -545 4173 -511
rect 4341 -545 4357 -511
rect 4157 -561 4357 -545
rect 4415 -511 4615 -464
rect 4415 -545 4431 -511
rect 4599 -545 4615 -511
rect 4415 -561 4615 -545
<< polycont >>
rect -4599 -545 -4431 -511
rect -4341 -545 -4173 -511
rect -4083 -545 -3915 -511
rect -3825 -545 -3657 -511
rect -3567 -545 -3399 -511
rect -3309 -545 -3141 -511
rect -3051 -545 -2883 -511
rect -2793 -545 -2625 -511
rect -2535 -545 -2367 -511
rect -2277 -545 -2109 -511
rect -2019 -545 -1851 -511
rect -1761 -545 -1593 -511
rect -1503 -545 -1335 -511
rect -1245 -545 -1077 -511
rect -987 -545 -819 -511
rect -729 -545 -561 -511
rect -471 -545 -303 -511
rect -213 -545 -45 -511
rect 45 -545 213 -511
rect 303 -545 471 -511
rect 561 -545 729 -511
rect 819 -545 987 -511
rect 1077 -545 1245 -511
rect 1335 -545 1503 -511
rect 1593 -545 1761 -511
rect 1851 -545 2019 -511
rect 2109 -545 2277 -511
rect 2367 -545 2535 -511
rect 2625 -545 2793 -511
rect 2883 -545 3051 -511
rect 3141 -545 3309 -511
rect 3399 -545 3567 -511
rect 3657 -545 3825 -511
rect 3915 -545 4083 -511
rect 4173 -545 4341 -511
rect 4431 -545 4599 -511
<< locali >>
rect -4775 614 -4679 648
rect 4679 614 4775 648
rect -4775 551 -4741 614
rect 4741 551 4775 614
rect -4661 524 -4627 540
rect -4661 -468 -4627 -452
rect -4403 524 -4369 540
rect -4403 -468 -4369 -452
rect -4145 524 -4111 540
rect -4145 -468 -4111 -452
rect -3887 524 -3853 540
rect -3887 -468 -3853 -452
rect -3629 524 -3595 540
rect -3629 -468 -3595 -452
rect -3371 524 -3337 540
rect -3371 -468 -3337 -452
rect -3113 524 -3079 540
rect -3113 -468 -3079 -452
rect -2855 524 -2821 540
rect -2855 -468 -2821 -452
rect -2597 524 -2563 540
rect -2597 -468 -2563 -452
rect -2339 524 -2305 540
rect -2339 -468 -2305 -452
rect -2081 524 -2047 540
rect -2081 -468 -2047 -452
rect -1823 524 -1789 540
rect -1823 -468 -1789 -452
rect -1565 524 -1531 540
rect -1565 -468 -1531 -452
rect -1307 524 -1273 540
rect -1307 -468 -1273 -452
rect -1049 524 -1015 540
rect -1049 -468 -1015 -452
rect -791 524 -757 540
rect -791 -468 -757 -452
rect -533 524 -499 540
rect -533 -468 -499 -452
rect -275 524 -241 540
rect -275 -468 -241 -452
rect -17 524 17 540
rect -17 -468 17 -452
rect 241 524 275 540
rect 241 -468 275 -452
rect 499 524 533 540
rect 499 -468 533 -452
rect 757 524 791 540
rect 757 -468 791 -452
rect 1015 524 1049 540
rect 1015 -468 1049 -452
rect 1273 524 1307 540
rect 1273 -468 1307 -452
rect 1531 524 1565 540
rect 1531 -468 1565 -452
rect 1789 524 1823 540
rect 1789 -468 1823 -452
rect 2047 524 2081 540
rect 2047 -468 2081 -452
rect 2305 524 2339 540
rect 2305 -468 2339 -452
rect 2563 524 2597 540
rect 2563 -468 2597 -452
rect 2821 524 2855 540
rect 2821 -468 2855 -452
rect 3079 524 3113 540
rect 3079 -468 3113 -452
rect 3337 524 3371 540
rect 3337 -468 3371 -452
rect 3595 524 3629 540
rect 3595 -468 3629 -452
rect 3853 524 3887 540
rect 3853 -468 3887 -452
rect 4111 524 4145 540
rect 4111 -468 4145 -452
rect 4369 524 4403 540
rect 4369 -468 4403 -452
rect 4627 524 4661 540
rect 4627 -468 4661 -452
rect -4615 -545 -4599 -511
rect -4431 -545 -4415 -511
rect -4357 -545 -4341 -511
rect -4173 -545 -4157 -511
rect -4099 -545 -4083 -511
rect -3915 -545 -3899 -511
rect -3841 -545 -3825 -511
rect -3657 -545 -3641 -511
rect -3583 -545 -3567 -511
rect -3399 -545 -3383 -511
rect -3325 -545 -3309 -511
rect -3141 -545 -3125 -511
rect -3067 -545 -3051 -511
rect -2883 -545 -2867 -511
rect -2809 -545 -2793 -511
rect -2625 -545 -2609 -511
rect -2551 -545 -2535 -511
rect -2367 -545 -2351 -511
rect -2293 -545 -2277 -511
rect -2109 -545 -2093 -511
rect -2035 -545 -2019 -511
rect -1851 -545 -1835 -511
rect -1777 -545 -1761 -511
rect -1593 -545 -1577 -511
rect -1519 -545 -1503 -511
rect -1335 -545 -1319 -511
rect -1261 -545 -1245 -511
rect -1077 -545 -1061 -511
rect -1003 -545 -987 -511
rect -819 -545 -803 -511
rect -745 -545 -729 -511
rect -561 -545 -545 -511
rect -487 -545 -471 -511
rect -303 -545 -287 -511
rect -229 -545 -213 -511
rect -45 -545 -29 -511
rect 29 -545 45 -511
rect 213 -545 229 -511
rect 287 -545 303 -511
rect 471 -545 487 -511
rect 545 -545 561 -511
rect 729 -545 745 -511
rect 803 -545 819 -511
rect 987 -545 1003 -511
rect 1061 -545 1077 -511
rect 1245 -545 1261 -511
rect 1319 -545 1335 -511
rect 1503 -545 1519 -511
rect 1577 -545 1593 -511
rect 1761 -545 1777 -511
rect 1835 -545 1851 -511
rect 2019 -545 2035 -511
rect 2093 -545 2109 -511
rect 2277 -545 2293 -511
rect 2351 -545 2367 -511
rect 2535 -545 2551 -511
rect 2609 -545 2625 -511
rect 2793 -545 2809 -511
rect 2867 -545 2883 -511
rect 3051 -545 3067 -511
rect 3125 -545 3141 -511
rect 3309 -545 3325 -511
rect 3383 -545 3399 -511
rect 3567 -545 3583 -511
rect 3641 -545 3657 -511
rect 3825 -545 3841 -511
rect 3899 -545 3915 -511
rect 4083 -545 4099 -511
rect 4157 -545 4173 -511
rect 4341 -545 4357 -511
rect 4415 -545 4431 -511
rect 4599 -545 4615 -511
rect -4775 -614 -4741 -551
rect 4741 -614 4775 -551
rect -4775 -648 -4679 -614
rect 4679 -648 4775 -614
<< viali >>
rect -4661 -452 -4627 524
rect -4403 -452 -4369 524
rect -4145 -452 -4111 524
rect -3887 -452 -3853 524
rect -3629 -452 -3595 524
rect -3371 -452 -3337 524
rect -3113 -452 -3079 524
rect -2855 -452 -2821 524
rect -2597 -452 -2563 524
rect -2339 -452 -2305 524
rect -2081 -452 -2047 524
rect -1823 -452 -1789 524
rect -1565 -452 -1531 524
rect -1307 -452 -1273 524
rect -1049 -452 -1015 524
rect -791 -452 -757 524
rect -533 -452 -499 524
rect -275 -452 -241 524
rect -17 -452 17 524
rect 241 -452 275 524
rect 499 -452 533 524
rect 757 -452 791 524
rect 1015 -452 1049 524
rect 1273 -452 1307 524
rect 1531 -452 1565 524
rect 1789 -452 1823 524
rect 2047 -452 2081 524
rect 2305 -452 2339 524
rect 2563 -452 2597 524
rect 2821 -452 2855 524
rect 3079 -452 3113 524
rect 3337 -452 3371 524
rect 3595 -452 3629 524
rect 3853 -452 3887 524
rect 4111 -452 4145 524
rect 4369 -452 4403 524
rect 4627 -452 4661 524
rect -4599 -545 -4431 -511
rect -4341 -545 -4173 -511
rect -4083 -545 -3915 -511
rect -3825 -545 -3657 -511
rect -3567 -545 -3399 -511
rect -3309 -545 -3141 -511
rect -3051 -545 -2883 -511
rect -2793 -545 -2625 -511
rect -2535 -545 -2367 -511
rect -2277 -545 -2109 -511
rect -2019 -545 -1851 -511
rect -1761 -545 -1593 -511
rect -1503 -545 -1335 -511
rect -1245 -545 -1077 -511
rect -987 -545 -819 -511
rect -729 -545 -561 -511
rect -471 -545 -303 -511
rect -213 -545 -45 -511
rect 45 -545 213 -511
rect 303 -545 471 -511
rect 561 -545 729 -511
rect 819 -545 987 -511
rect 1077 -545 1245 -511
rect 1335 -545 1503 -511
rect 1593 -545 1761 -511
rect 1851 -545 2019 -511
rect 2109 -545 2277 -511
rect 2367 -545 2535 -511
rect 2625 -545 2793 -511
rect 2883 -545 3051 -511
rect 3141 -545 3309 -511
rect 3399 -545 3567 -511
rect 3657 -545 3825 -511
rect 3915 -545 4083 -511
rect 4173 -545 4341 -511
rect 4431 -545 4599 -511
<< metal1 >>
rect -4667 524 -4621 536
rect -4667 -452 -4661 524
rect -4627 -452 -4621 524
rect -4667 -464 -4621 -452
rect -4409 524 -4363 536
rect -4409 -452 -4403 524
rect -4369 -452 -4363 524
rect -4409 -464 -4363 -452
rect -4151 524 -4105 536
rect -4151 -452 -4145 524
rect -4111 -452 -4105 524
rect -4151 -464 -4105 -452
rect -3893 524 -3847 536
rect -3893 -452 -3887 524
rect -3853 -452 -3847 524
rect -3893 -464 -3847 -452
rect -3635 524 -3589 536
rect -3635 -452 -3629 524
rect -3595 -452 -3589 524
rect -3635 -464 -3589 -452
rect -3377 524 -3331 536
rect -3377 -452 -3371 524
rect -3337 -452 -3331 524
rect -3377 -464 -3331 -452
rect -3119 524 -3073 536
rect -3119 -452 -3113 524
rect -3079 -452 -3073 524
rect -3119 -464 -3073 -452
rect -2861 524 -2815 536
rect -2861 -452 -2855 524
rect -2821 -452 -2815 524
rect -2861 -464 -2815 -452
rect -2603 524 -2557 536
rect -2603 -452 -2597 524
rect -2563 -452 -2557 524
rect -2603 -464 -2557 -452
rect -2345 524 -2299 536
rect -2345 -452 -2339 524
rect -2305 -452 -2299 524
rect -2345 -464 -2299 -452
rect -2087 524 -2041 536
rect -2087 -452 -2081 524
rect -2047 -452 -2041 524
rect -2087 -464 -2041 -452
rect -1829 524 -1783 536
rect -1829 -452 -1823 524
rect -1789 -452 -1783 524
rect -1829 -464 -1783 -452
rect -1571 524 -1525 536
rect -1571 -452 -1565 524
rect -1531 -452 -1525 524
rect -1571 -464 -1525 -452
rect -1313 524 -1267 536
rect -1313 -452 -1307 524
rect -1273 -452 -1267 524
rect -1313 -464 -1267 -452
rect -1055 524 -1009 536
rect -1055 -452 -1049 524
rect -1015 -452 -1009 524
rect -1055 -464 -1009 -452
rect -797 524 -751 536
rect -797 -452 -791 524
rect -757 -452 -751 524
rect -797 -464 -751 -452
rect -539 524 -493 536
rect -539 -452 -533 524
rect -499 -452 -493 524
rect -539 -464 -493 -452
rect -281 524 -235 536
rect -281 -452 -275 524
rect -241 -452 -235 524
rect -281 -464 -235 -452
rect -23 524 23 536
rect -23 -452 -17 524
rect 17 -452 23 524
rect -23 -464 23 -452
rect 235 524 281 536
rect 235 -452 241 524
rect 275 -452 281 524
rect 235 -464 281 -452
rect 493 524 539 536
rect 493 -452 499 524
rect 533 -452 539 524
rect 493 -464 539 -452
rect 751 524 797 536
rect 751 -452 757 524
rect 791 -452 797 524
rect 751 -464 797 -452
rect 1009 524 1055 536
rect 1009 -452 1015 524
rect 1049 -452 1055 524
rect 1009 -464 1055 -452
rect 1267 524 1313 536
rect 1267 -452 1273 524
rect 1307 -452 1313 524
rect 1267 -464 1313 -452
rect 1525 524 1571 536
rect 1525 -452 1531 524
rect 1565 -452 1571 524
rect 1525 -464 1571 -452
rect 1783 524 1829 536
rect 1783 -452 1789 524
rect 1823 -452 1829 524
rect 1783 -464 1829 -452
rect 2041 524 2087 536
rect 2041 -452 2047 524
rect 2081 -452 2087 524
rect 2041 -464 2087 -452
rect 2299 524 2345 536
rect 2299 -452 2305 524
rect 2339 -452 2345 524
rect 2299 -464 2345 -452
rect 2557 524 2603 536
rect 2557 -452 2563 524
rect 2597 -452 2603 524
rect 2557 -464 2603 -452
rect 2815 524 2861 536
rect 2815 -452 2821 524
rect 2855 -452 2861 524
rect 2815 -464 2861 -452
rect 3073 524 3119 536
rect 3073 -452 3079 524
rect 3113 -452 3119 524
rect 3073 -464 3119 -452
rect 3331 524 3377 536
rect 3331 -452 3337 524
rect 3371 -452 3377 524
rect 3331 -464 3377 -452
rect 3589 524 3635 536
rect 3589 -452 3595 524
rect 3629 -452 3635 524
rect 3589 -464 3635 -452
rect 3847 524 3893 536
rect 3847 -452 3853 524
rect 3887 -452 3893 524
rect 3847 -464 3893 -452
rect 4105 524 4151 536
rect 4105 -452 4111 524
rect 4145 -452 4151 524
rect 4105 -464 4151 -452
rect 4363 524 4409 536
rect 4363 -452 4369 524
rect 4403 -452 4409 524
rect 4363 -464 4409 -452
rect 4621 524 4667 536
rect 4621 -452 4627 524
rect 4661 -452 4667 524
rect 4621 -464 4667 -452
rect -4611 -511 -4419 -505
rect -4611 -545 -4599 -511
rect -4431 -545 -4419 -511
rect -4611 -551 -4419 -545
rect -4353 -511 -4161 -505
rect -4353 -545 -4341 -511
rect -4173 -545 -4161 -511
rect -4353 -551 -4161 -545
rect -4095 -511 -3903 -505
rect -4095 -545 -4083 -511
rect -3915 -545 -3903 -511
rect -4095 -551 -3903 -545
rect -3837 -511 -3645 -505
rect -3837 -545 -3825 -511
rect -3657 -545 -3645 -511
rect -3837 -551 -3645 -545
rect -3579 -511 -3387 -505
rect -3579 -545 -3567 -511
rect -3399 -545 -3387 -511
rect -3579 -551 -3387 -545
rect -3321 -511 -3129 -505
rect -3321 -545 -3309 -511
rect -3141 -545 -3129 -511
rect -3321 -551 -3129 -545
rect -3063 -511 -2871 -505
rect -3063 -545 -3051 -511
rect -2883 -545 -2871 -511
rect -3063 -551 -2871 -545
rect -2805 -511 -2613 -505
rect -2805 -545 -2793 -511
rect -2625 -545 -2613 -511
rect -2805 -551 -2613 -545
rect -2547 -511 -2355 -505
rect -2547 -545 -2535 -511
rect -2367 -545 -2355 -511
rect -2547 -551 -2355 -545
rect -2289 -511 -2097 -505
rect -2289 -545 -2277 -511
rect -2109 -545 -2097 -511
rect -2289 -551 -2097 -545
rect -2031 -511 -1839 -505
rect -2031 -545 -2019 -511
rect -1851 -545 -1839 -511
rect -2031 -551 -1839 -545
rect -1773 -511 -1581 -505
rect -1773 -545 -1761 -511
rect -1593 -545 -1581 -511
rect -1773 -551 -1581 -545
rect -1515 -511 -1323 -505
rect -1515 -545 -1503 -511
rect -1335 -545 -1323 -511
rect -1515 -551 -1323 -545
rect -1257 -511 -1065 -505
rect -1257 -545 -1245 -511
rect -1077 -545 -1065 -511
rect -1257 -551 -1065 -545
rect -999 -511 -807 -505
rect -999 -545 -987 -511
rect -819 -545 -807 -511
rect -999 -551 -807 -545
rect -741 -511 -549 -505
rect -741 -545 -729 -511
rect -561 -545 -549 -511
rect -741 -551 -549 -545
rect -483 -511 -291 -505
rect -483 -545 -471 -511
rect -303 -545 -291 -511
rect -483 -551 -291 -545
rect -225 -511 -33 -505
rect -225 -545 -213 -511
rect -45 -545 -33 -511
rect -225 -551 -33 -545
rect 33 -511 225 -505
rect 33 -545 45 -511
rect 213 -545 225 -511
rect 33 -551 225 -545
rect 291 -511 483 -505
rect 291 -545 303 -511
rect 471 -545 483 -511
rect 291 -551 483 -545
rect 549 -511 741 -505
rect 549 -545 561 -511
rect 729 -545 741 -511
rect 549 -551 741 -545
rect 807 -511 999 -505
rect 807 -545 819 -511
rect 987 -545 999 -511
rect 807 -551 999 -545
rect 1065 -511 1257 -505
rect 1065 -545 1077 -511
rect 1245 -545 1257 -511
rect 1065 -551 1257 -545
rect 1323 -511 1515 -505
rect 1323 -545 1335 -511
rect 1503 -545 1515 -511
rect 1323 -551 1515 -545
rect 1581 -511 1773 -505
rect 1581 -545 1593 -511
rect 1761 -545 1773 -511
rect 1581 -551 1773 -545
rect 1839 -511 2031 -505
rect 1839 -545 1851 -511
rect 2019 -545 2031 -511
rect 1839 -551 2031 -545
rect 2097 -511 2289 -505
rect 2097 -545 2109 -511
rect 2277 -545 2289 -511
rect 2097 -551 2289 -545
rect 2355 -511 2547 -505
rect 2355 -545 2367 -511
rect 2535 -545 2547 -511
rect 2355 -551 2547 -545
rect 2613 -511 2805 -505
rect 2613 -545 2625 -511
rect 2793 -545 2805 -511
rect 2613 -551 2805 -545
rect 2871 -511 3063 -505
rect 2871 -545 2883 -511
rect 3051 -545 3063 -511
rect 2871 -551 3063 -545
rect 3129 -511 3321 -505
rect 3129 -545 3141 -511
rect 3309 -545 3321 -511
rect 3129 -551 3321 -545
rect 3387 -511 3579 -505
rect 3387 -545 3399 -511
rect 3567 -545 3579 -511
rect 3387 -551 3579 -545
rect 3645 -511 3837 -505
rect 3645 -545 3657 -511
rect 3825 -545 3837 -511
rect 3645 -551 3837 -545
rect 3903 -511 4095 -505
rect 3903 -545 3915 -511
rect 4083 -545 4095 -511
rect 3903 -551 4095 -545
rect 4161 -511 4353 -505
rect 4161 -545 4173 -511
rect 4341 -545 4353 -511
rect 4161 -551 4353 -545
rect 4419 -511 4611 -505
rect 4419 -545 4431 -511
rect 4599 -545 4611 -511
rect 4419 -551 4611 -545
<< properties >>
string FIXED_BBOX -4758 -631 4758 631
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 1 m 1 nf 36 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
