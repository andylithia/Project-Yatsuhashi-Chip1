magic
tech sky130B
magscale 1 2
timestamp 1662234432
<< nwell >>
rect -296 -21071 296 21071
<< pmos >>
rect -100 19923 100 20923
rect -100 18758 100 19758
rect -100 17593 100 18593
rect -100 16428 100 17428
rect -100 15263 100 16263
rect -100 14098 100 15098
rect -100 12933 100 13933
rect -100 11768 100 12768
rect -100 10603 100 11603
rect -100 9438 100 10438
rect -100 8273 100 9273
rect -100 7108 100 8108
rect -100 5943 100 6943
rect -100 4778 100 5778
rect -100 3613 100 4613
rect -100 2448 100 3448
rect -100 1283 100 2283
rect -100 118 100 1118
rect -100 -1047 100 -47
rect -100 -2212 100 -1212
rect -100 -3377 100 -2377
rect -100 -4542 100 -3542
rect -100 -5707 100 -4707
rect -100 -6872 100 -5872
rect -100 -8037 100 -7037
rect -100 -9202 100 -8202
rect -100 -10367 100 -9367
rect -100 -11532 100 -10532
rect -100 -12697 100 -11697
rect -100 -13862 100 -12862
rect -100 -15027 100 -14027
rect -100 -16192 100 -15192
rect -100 -17357 100 -16357
rect -100 -18522 100 -17522
rect -100 -19687 100 -18687
rect -100 -20852 100 -19852
<< pdiff >>
rect -158 20911 -100 20923
rect -158 19935 -146 20911
rect -112 19935 -100 20911
rect -158 19923 -100 19935
rect 100 20911 158 20923
rect 100 19935 112 20911
rect 146 19935 158 20911
rect 100 19923 158 19935
rect -158 19746 -100 19758
rect -158 18770 -146 19746
rect -112 18770 -100 19746
rect -158 18758 -100 18770
rect 100 19746 158 19758
rect 100 18770 112 19746
rect 146 18770 158 19746
rect 100 18758 158 18770
rect -158 18581 -100 18593
rect -158 17605 -146 18581
rect -112 17605 -100 18581
rect -158 17593 -100 17605
rect 100 18581 158 18593
rect 100 17605 112 18581
rect 146 17605 158 18581
rect 100 17593 158 17605
rect -158 17416 -100 17428
rect -158 16440 -146 17416
rect -112 16440 -100 17416
rect -158 16428 -100 16440
rect 100 17416 158 17428
rect 100 16440 112 17416
rect 146 16440 158 17416
rect 100 16428 158 16440
rect -158 16251 -100 16263
rect -158 15275 -146 16251
rect -112 15275 -100 16251
rect -158 15263 -100 15275
rect 100 16251 158 16263
rect 100 15275 112 16251
rect 146 15275 158 16251
rect 100 15263 158 15275
rect -158 15086 -100 15098
rect -158 14110 -146 15086
rect -112 14110 -100 15086
rect -158 14098 -100 14110
rect 100 15086 158 15098
rect 100 14110 112 15086
rect 146 14110 158 15086
rect 100 14098 158 14110
rect -158 13921 -100 13933
rect -158 12945 -146 13921
rect -112 12945 -100 13921
rect -158 12933 -100 12945
rect 100 13921 158 13933
rect 100 12945 112 13921
rect 146 12945 158 13921
rect 100 12933 158 12945
rect -158 12756 -100 12768
rect -158 11780 -146 12756
rect -112 11780 -100 12756
rect -158 11768 -100 11780
rect 100 12756 158 12768
rect 100 11780 112 12756
rect 146 11780 158 12756
rect 100 11768 158 11780
rect -158 11591 -100 11603
rect -158 10615 -146 11591
rect -112 10615 -100 11591
rect -158 10603 -100 10615
rect 100 11591 158 11603
rect 100 10615 112 11591
rect 146 10615 158 11591
rect 100 10603 158 10615
rect -158 10426 -100 10438
rect -158 9450 -146 10426
rect -112 9450 -100 10426
rect -158 9438 -100 9450
rect 100 10426 158 10438
rect 100 9450 112 10426
rect 146 9450 158 10426
rect 100 9438 158 9450
rect -158 9261 -100 9273
rect -158 8285 -146 9261
rect -112 8285 -100 9261
rect -158 8273 -100 8285
rect 100 9261 158 9273
rect 100 8285 112 9261
rect 146 8285 158 9261
rect 100 8273 158 8285
rect -158 8096 -100 8108
rect -158 7120 -146 8096
rect -112 7120 -100 8096
rect -158 7108 -100 7120
rect 100 8096 158 8108
rect 100 7120 112 8096
rect 146 7120 158 8096
rect 100 7108 158 7120
rect -158 6931 -100 6943
rect -158 5955 -146 6931
rect -112 5955 -100 6931
rect -158 5943 -100 5955
rect 100 6931 158 6943
rect 100 5955 112 6931
rect 146 5955 158 6931
rect 100 5943 158 5955
rect -158 5766 -100 5778
rect -158 4790 -146 5766
rect -112 4790 -100 5766
rect -158 4778 -100 4790
rect 100 5766 158 5778
rect 100 4790 112 5766
rect 146 4790 158 5766
rect 100 4778 158 4790
rect -158 4601 -100 4613
rect -158 3625 -146 4601
rect -112 3625 -100 4601
rect -158 3613 -100 3625
rect 100 4601 158 4613
rect 100 3625 112 4601
rect 146 3625 158 4601
rect 100 3613 158 3625
rect -158 3436 -100 3448
rect -158 2460 -146 3436
rect -112 2460 -100 3436
rect -158 2448 -100 2460
rect 100 3436 158 3448
rect 100 2460 112 3436
rect 146 2460 158 3436
rect 100 2448 158 2460
rect -158 2271 -100 2283
rect -158 1295 -146 2271
rect -112 1295 -100 2271
rect -158 1283 -100 1295
rect 100 2271 158 2283
rect 100 1295 112 2271
rect 146 1295 158 2271
rect 100 1283 158 1295
rect -158 1106 -100 1118
rect -158 130 -146 1106
rect -112 130 -100 1106
rect -158 118 -100 130
rect 100 1106 158 1118
rect 100 130 112 1106
rect 146 130 158 1106
rect 100 118 158 130
rect -158 -59 -100 -47
rect -158 -1035 -146 -59
rect -112 -1035 -100 -59
rect -158 -1047 -100 -1035
rect 100 -59 158 -47
rect 100 -1035 112 -59
rect 146 -1035 158 -59
rect 100 -1047 158 -1035
rect -158 -1224 -100 -1212
rect -158 -2200 -146 -1224
rect -112 -2200 -100 -1224
rect -158 -2212 -100 -2200
rect 100 -1224 158 -1212
rect 100 -2200 112 -1224
rect 146 -2200 158 -1224
rect 100 -2212 158 -2200
rect -158 -2389 -100 -2377
rect -158 -3365 -146 -2389
rect -112 -3365 -100 -2389
rect -158 -3377 -100 -3365
rect 100 -2389 158 -2377
rect 100 -3365 112 -2389
rect 146 -3365 158 -2389
rect 100 -3377 158 -3365
rect -158 -3554 -100 -3542
rect -158 -4530 -146 -3554
rect -112 -4530 -100 -3554
rect -158 -4542 -100 -4530
rect 100 -3554 158 -3542
rect 100 -4530 112 -3554
rect 146 -4530 158 -3554
rect 100 -4542 158 -4530
rect -158 -4719 -100 -4707
rect -158 -5695 -146 -4719
rect -112 -5695 -100 -4719
rect -158 -5707 -100 -5695
rect 100 -4719 158 -4707
rect 100 -5695 112 -4719
rect 146 -5695 158 -4719
rect 100 -5707 158 -5695
rect -158 -5884 -100 -5872
rect -158 -6860 -146 -5884
rect -112 -6860 -100 -5884
rect -158 -6872 -100 -6860
rect 100 -5884 158 -5872
rect 100 -6860 112 -5884
rect 146 -6860 158 -5884
rect 100 -6872 158 -6860
rect -158 -7049 -100 -7037
rect -158 -8025 -146 -7049
rect -112 -8025 -100 -7049
rect -158 -8037 -100 -8025
rect 100 -7049 158 -7037
rect 100 -8025 112 -7049
rect 146 -8025 158 -7049
rect 100 -8037 158 -8025
rect -158 -8214 -100 -8202
rect -158 -9190 -146 -8214
rect -112 -9190 -100 -8214
rect -158 -9202 -100 -9190
rect 100 -8214 158 -8202
rect 100 -9190 112 -8214
rect 146 -9190 158 -8214
rect 100 -9202 158 -9190
rect -158 -9379 -100 -9367
rect -158 -10355 -146 -9379
rect -112 -10355 -100 -9379
rect -158 -10367 -100 -10355
rect 100 -9379 158 -9367
rect 100 -10355 112 -9379
rect 146 -10355 158 -9379
rect 100 -10367 158 -10355
rect -158 -10544 -100 -10532
rect -158 -11520 -146 -10544
rect -112 -11520 -100 -10544
rect -158 -11532 -100 -11520
rect 100 -10544 158 -10532
rect 100 -11520 112 -10544
rect 146 -11520 158 -10544
rect 100 -11532 158 -11520
rect -158 -11709 -100 -11697
rect -158 -12685 -146 -11709
rect -112 -12685 -100 -11709
rect -158 -12697 -100 -12685
rect 100 -11709 158 -11697
rect 100 -12685 112 -11709
rect 146 -12685 158 -11709
rect 100 -12697 158 -12685
rect -158 -12874 -100 -12862
rect -158 -13850 -146 -12874
rect -112 -13850 -100 -12874
rect -158 -13862 -100 -13850
rect 100 -12874 158 -12862
rect 100 -13850 112 -12874
rect 146 -13850 158 -12874
rect 100 -13862 158 -13850
rect -158 -14039 -100 -14027
rect -158 -15015 -146 -14039
rect -112 -15015 -100 -14039
rect -158 -15027 -100 -15015
rect 100 -14039 158 -14027
rect 100 -15015 112 -14039
rect 146 -15015 158 -14039
rect 100 -15027 158 -15015
rect -158 -15204 -100 -15192
rect -158 -16180 -146 -15204
rect -112 -16180 -100 -15204
rect -158 -16192 -100 -16180
rect 100 -15204 158 -15192
rect 100 -16180 112 -15204
rect 146 -16180 158 -15204
rect 100 -16192 158 -16180
rect -158 -16369 -100 -16357
rect -158 -17345 -146 -16369
rect -112 -17345 -100 -16369
rect -158 -17357 -100 -17345
rect 100 -16369 158 -16357
rect 100 -17345 112 -16369
rect 146 -17345 158 -16369
rect 100 -17357 158 -17345
rect -158 -17534 -100 -17522
rect -158 -18510 -146 -17534
rect -112 -18510 -100 -17534
rect -158 -18522 -100 -18510
rect 100 -17534 158 -17522
rect 100 -18510 112 -17534
rect 146 -18510 158 -17534
rect 100 -18522 158 -18510
rect -158 -18699 -100 -18687
rect -158 -19675 -146 -18699
rect -112 -19675 -100 -18699
rect -158 -19687 -100 -19675
rect 100 -18699 158 -18687
rect 100 -19675 112 -18699
rect 146 -19675 158 -18699
rect 100 -19687 158 -19675
rect -158 -19864 -100 -19852
rect -158 -20840 -146 -19864
rect -112 -20840 -100 -19864
rect -158 -20852 -100 -20840
rect 100 -19864 158 -19852
rect 100 -20840 112 -19864
rect 146 -20840 158 -19864
rect 100 -20852 158 -20840
<< pdiffc >>
rect -146 19935 -112 20911
rect 112 19935 146 20911
rect -146 18770 -112 19746
rect 112 18770 146 19746
rect -146 17605 -112 18581
rect 112 17605 146 18581
rect -146 16440 -112 17416
rect 112 16440 146 17416
rect -146 15275 -112 16251
rect 112 15275 146 16251
rect -146 14110 -112 15086
rect 112 14110 146 15086
rect -146 12945 -112 13921
rect 112 12945 146 13921
rect -146 11780 -112 12756
rect 112 11780 146 12756
rect -146 10615 -112 11591
rect 112 10615 146 11591
rect -146 9450 -112 10426
rect 112 9450 146 10426
rect -146 8285 -112 9261
rect 112 8285 146 9261
rect -146 7120 -112 8096
rect 112 7120 146 8096
rect -146 5955 -112 6931
rect 112 5955 146 6931
rect -146 4790 -112 5766
rect 112 4790 146 5766
rect -146 3625 -112 4601
rect 112 3625 146 4601
rect -146 2460 -112 3436
rect 112 2460 146 3436
rect -146 1295 -112 2271
rect 112 1295 146 2271
rect -146 130 -112 1106
rect 112 130 146 1106
rect -146 -1035 -112 -59
rect 112 -1035 146 -59
rect -146 -2200 -112 -1224
rect 112 -2200 146 -1224
rect -146 -3365 -112 -2389
rect 112 -3365 146 -2389
rect -146 -4530 -112 -3554
rect 112 -4530 146 -3554
rect -146 -5695 -112 -4719
rect 112 -5695 146 -4719
rect -146 -6860 -112 -5884
rect 112 -6860 146 -5884
rect -146 -8025 -112 -7049
rect 112 -8025 146 -7049
rect -146 -9190 -112 -8214
rect 112 -9190 146 -8214
rect -146 -10355 -112 -9379
rect 112 -10355 146 -9379
rect -146 -11520 -112 -10544
rect 112 -11520 146 -10544
rect -146 -12685 -112 -11709
rect 112 -12685 146 -11709
rect -146 -13850 -112 -12874
rect 112 -13850 146 -12874
rect -146 -15015 -112 -14039
rect 112 -15015 146 -14039
rect -146 -16180 -112 -15204
rect 112 -16180 146 -15204
rect -146 -17345 -112 -16369
rect 112 -17345 146 -16369
rect -146 -18510 -112 -17534
rect 112 -18510 146 -17534
rect -146 -19675 -112 -18699
rect 112 -19675 146 -18699
rect -146 -20840 -112 -19864
rect 112 -20840 146 -19864
<< nsubdiff >>
rect -260 21001 -164 21035
rect 164 21001 260 21035
rect -260 20939 -226 21001
rect 226 20939 260 21001
rect -260 -21001 -226 -20939
rect 226 -21001 260 -20939
rect -260 -21035 -164 -21001
rect 164 -21035 260 -21001
<< nsubdiffcont >>
rect -164 21001 164 21035
rect -260 -20939 -226 20939
rect 226 -20939 260 20939
rect -164 -21035 164 -21001
<< poly >>
rect -100 20923 100 20949
rect -100 19876 100 19923
rect -100 19842 -84 19876
rect 84 19842 100 19876
rect -100 19826 100 19842
rect -100 19758 100 19784
rect -100 18711 100 18758
rect -100 18677 -84 18711
rect 84 18677 100 18711
rect -100 18661 100 18677
rect -100 18593 100 18619
rect -100 17546 100 17593
rect -100 17512 -84 17546
rect 84 17512 100 17546
rect -100 17496 100 17512
rect -100 17428 100 17454
rect -100 16381 100 16428
rect -100 16347 -84 16381
rect 84 16347 100 16381
rect -100 16331 100 16347
rect -100 16263 100 16289
rect -100 15216 100 15263
rect -100 15182 -84 15216
rect 84 15182 100 15216
rect -100 15166 100 15182
rect -100 15098 100 15124
rect -100 14051 100 14098
rect -100 14017 -84 14051
rect 84 14017 100 14051
rect -100 14001 100 14017
rect -100 13933 100 13959
rect -100 12886 100 12933
rect -100 12852 -84 12886
rect 84 12852 100 12886
rect -100 12836 100 12852
rect -100 12768 100 12794
rect -100 11721 100 11768
rect -100 11687 -84 11721
rect 84 11687 100 11721
rect -100 11671 100 11687
rect -100 11603 100 11629
rect -100 10556 100 10603
rect -100 10522 -84 10556
rect 84 10522 100 10556
rect -100 10506 100 10522
rect -100 10438 100 10464
rect -100 9391 100 9438
rect -100 9357 -84 9391
rect 84 9357 100 9391
rect -100 9341 100 9357
rect -100 9273 100 9299
rect -100 8226 100 8273
rect -100 8192 -84 8226
rect 84 8192 100 8226
rect -100 8176 100 8192
rect -100 8108 100 8134
rect -100 7061 100 7108
rect -100 7027 -84 7061
rect 84 7027 100 7061
rect -100 7011 100 7027
rect -100 6943 100 6969
rect -100 5896 100 5943
rect -100 5862 -84 5896
rect 84 5862 100 5896
rect -100 5846 100 5862
rect -100 5778 100 5804
rect -100 4731 100 4778
rect -100 4697 -84 4731
rect 84 4697 100 4731
rect -100 4681 100 4697
rect -100 4613 100 4639
rect -100 3566 100 3613
rect -100 3532 -84 3566
rect 84 3532 100 3566
rect -100 3516 100 3532
rect -100 3448 100 3474
rect -100 2401 100 2448
rect -100 2367 -84 2401
rect 84 2367 100 2401
rect -100 2351 100 2367
rect -100 2283 100 2309
rect -100 1236 100 1283
rect -100 1202 -84 1236
rect 84 1202 100 1236
rect -100 1186 100 1202
rect -100 1118 100 1144
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -47 100 -21
rect -100 -1094 100 -1047
rect -100 -1128 -84 -1094
rect 84 -1128 100 -1094
rect -100 -1144 100 -1128
rect -100 -1212 100 -1186
rect -100 -2259 100 -2212
rect -100 -2293 -84 -2259
rect 84 -2293 100 -2259
rect -100 -2309 100 -2293
rect -100 -2377 100 -2351
rect -100 -3424 100 -3377
rect -100 -3458 -84 -3424
rect 84 -3458 100 -3424
rect -100 -3474 100 -3458
rect -100 -3542 100 -3516
rect -100 -4589 100 -4542
rect -100 -4623 -84 -4589
rect 84 -4623 100 -4589
rect -100 -4639 100 -4623
rect -100 -4707 100 -4681
rect -100 -5754 100 -5707
rect -100 -5788 -84 -5754
rect 84 -5788 100 -5754
rect -100 -5804 100 -5788
rect -100 -5872 100 -5846
rect -100 -6919 100 -6872
rect -100 -6953 -84 -6919
rect 84 -6953 100 -6919
rect -100 -6969 100 -6953
rect -100 -7037 100 -7011
rect -100 -8084 100 -8037
rect -100 -8118 -84 -8084
rect 84 -8118 100 -8084
rect -100 -8134 100 -8118
rect -100 -8202 100 -8176
rect -100 -9249 100 -9202
rect -100 -9283 -84 -9249
rect 84 -9283 100 -9249
rect -100 -9299 100 -9283
rect -100 -9367 100 -9341
rect -100 -10414 100 -10367
rect -100 -10448 -84 -10414
rect 84 -10448 100 -10414
rect -100 -10464 100 -10448
rect -100 -10532 100 -10506
rect -100 -11579 100 -11532
rect -100 -11613 -84 -11579
rect 84 -11613 100 -11579
rect -100 -11629 100 -11613
rect -100 -11697 100 -11671
rect -100 -12744 100 -12697
rect -100 -12778 -84 -12744
rect 84 -12778 100 -12744
rect -100 -12794 100 -12778
rect -100 -12862 100 -12836
rect -100 -13909 100 -13862
rect -100 -13943 -84 -13909
rect 84 -13943 100 -13909
rect -100 -13959 100 -13943
rect -100 -14027 100 -14001
rect -100 -15074 100 -15027
rect -100 -15108 -84 -15074
rect 84 -15108 100 -15074
rect -100 -15124 100 -15108
rect -100 -15192 100 -15166
rect -100 -16239 100 -16192
rect -100 -16273 -84 -16239
rect 84 -16273 100 -16239
rect -100 -16289 100 -16273
rect -100 -16357 100 -16331
rect -100 -17404 100 -17357
rect -100 -17438 -84 -17404
rect 84 -17438 100 -17404
rect -100 -17454 100 -17438
rect -100 -17522 100 -17496
rect -100 -18569 100 -18522
rect -100 -18603 -84 -18569
rect 84 -18603 100 -18569
rect -100 -18619 100 -18603
rect -100 -18687 100 -18661
rect -100 -19734 100 -19687
rect -100 -19768 -84 -19734
rect 84 -19768 100 -19734
rect -100 -19784 100 -19768
rect -100 -19852 100 -19826
rect -100 -20899 100 -20852
rect -100 -20933 -84 -20899
rect 84 -20933 100 -20899
rect -100 -20949 100 -20933
<< polycont >>
rect -84 19842 84 19876
rect -84 18677 84 18711
rect -84 17512 84 17546
rect -84 16347 84 16381
rect -84 15182 84 15216
rect -84 14017 84 14051
rect -84 12852 84 12886
rect -84 11687 84 11721
rect -84 10522 84 10556
rect -84 9357 84 9391
rect -84 8192 84 8226
rect -84 7027 84 7061
rect -84 5862 84 5896
rect -84 4697 84 4731
rect -84 3532 84 3566
rect -84 2367 84 2401
rect -84 1202 84 1236
rect -84 37 84 71
rect -84 -1128 84 -1094
rect -84 -2293 84 -2259
rect -84 -3458 84 -3424
rect -84 -4623 84 -4589
rect -84 -5788 84 -5754
rect -84 -6953 84 -6919
rect -84 -8118 84 -8084
rect -84 -9283 84 -9249
rect -84 -10448 84 -10414
rect -84 -11613 84 -11579
rect -84 -12778 84 -12744
rect -84 -13943 84 -13909
rect -84 -15108 84 -15074
rect -84 -16273 84 -16239
rect -84 -17438 84 -17404
rect -84 -18603 84 -18569
rect -84 -19768 84 -19734
rect -84 -20933 84 -20899
<< locali >>
rect -260 21001 -164 21035
rect 164 21001 260 21035
rect -260 20939 -226 21001
rect 226 20939 260 21001
rect -146 20911 -112 20927
rect -146 19919 -112 19935
rect 112 20911 146 20927
rect 112 19919 146 19935
rect -100 19842 -84 19876
rect 84 19842 100 19876
rect -146 19746 -112 19762
rect -146 18754 -112 18770
rect 112 19746 146 19762
rect 112 18754 146 18770
rect -100 18677 -84 18711
rect 84 18677 100 18711
rect -146 18581 -112 18597
rect -146 17589 -112 17605
rect 112 18581 146 18597
rect 112 17589 146 17605
rect -100 17512 -84 17546
rect 84 17512 100 17546
rect -146 17416 -112 17432
rect -146 16424 -112 16440
rect 112 17416 146 17432
rect 112 16424 146 16440
rect -100 16347 -84 16381
rect 84 16347 100 16381
rect -146 16251 -112 16267
rect -146 15259 -112 15275
rect 112 16251 146 16267
rect 112 15259 146 15275
rect -100 15182 -84 15216
rect 84 15182 100 15216
rect -146 15086 -112 15102
rect -146 14094 -112 14110
rect 112 15086 146 15102
rect 112 14094 146 14110
rect -100 14017 -84 14051
rect 84 14017 100 14051
rect -146 13921 -112 13937
rect -146 12929 -112 12945
rect 112 13921 146 13937
rect 112 12929 146 12945
rect -100 12852 -84 12886
rect 84 12852 100 12886
rect -146 12756 -112 12772
rect -146 11764 -112 11780
rect 112 12756 146 12772
rect 112 11764 146 11780
rect -100 11687 -84 11721
rect 84 11687 100 11721
rect -146 11591 -112 11607
rect -146 10599 -112 10615
rect 112 11591 146 11607
rect 112 10599 146 10615
rect -100 10522 -84 10556
rect 84 10522 100 10556
rect -146 10426 -112 10442
rect -146 9434 -112 9450
rect 112 10426 146 10442
rect 112 9434 146 9450
rect -100 9357 -84 9391
rect 84 9357 100 9391
rect -146 9261 -112 9277
rect -146 8269 -112 8285
rect 112 9261 146 9277
rect 112 8269 146 8285
rect -100 8192 -84 8226
rect 84 8192 100 8226
rect -146 8096 -112 8112
rect -146 7104 -112 7120
rect 112 8096 146 8112
rect 112 7104 146 7120
rect -100 7027 -84 7061
rect 84 7027 100 7061
rect -146 6931 -112 6947
rect -146 5939 -112 5955
rect 112 6931 146 6947
rect 112 5939 146 5955
rect -100 5862 -84 5896
rect 84 5862 100 5896
rect -146 5766 -112 5782
rect -146 4774 -112 4790
rect 112 5766 146 5782
rect 112 4774 146 4790
rect -100 4697 -84 4731
rect 84 4697 100 4731
rect -146 4601 -112 4617
rect -146 3609 -112 3625
rect 112 4601 146 4617
rect 112 3609 146 3625
rect -100 3532 -84 3566
rect 84 3532 100 3566
rect -146 3436 -112 3452
rect -146 2444 -112 2460
rect 112 3436 146 3452
rect 112 2444 146 2460
rect -100 2367 -84 2401
rect 84 2367 100 2401
rect -146 2271 -112 2287
rect -146 1279 -112 1295
rect 112 2271 146 2287
rect 112 1279 146 1295
rect -100 1202 -84 1236
rect 84 1202 100 1236
rect -146 1106 -112 1122
rect -146 114 -112 130
rect 112 1106 146 1122
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -146 -59 -112 -43
rect -146 -1051 -112 -1035
rect 112 -59 146 -43
rect 112 -1051 146 -1035
rect -100 -1128 -84 -1094
rect 84 -1128 100 -1094
rect -146 -1224 -112 -1208
rect -146 -2216 -112 -2200
rect 112 -1224 146 -1208
rect 112 -2216 146 -2200
rect -100 -2293 -84 -2259
rect 84 -2293 100 -2259
rect -146 -2389 -112 -2373
rect -146 -3381 -112 -3365
rect 112 -2389 146 -2373
rect 112 -3381 146 -3365
rect -100 -3458 -84 -3424
rect 84 -3458 100 -3424
rect -146 -3554 -112 -3538
rect -146 -4546 -112 -4530
rect 112 -3554 146 -3538
rect 112 -4546 146 -4530
rect -100 -4623 -84 -4589
rect 84 -4623 100 -4589
rect -146 -4719 -112 -4703
rect -146 -5711 -112 -5695
rect 112 -4719 146 -4703
rect 112 -5711 146 -5695
rect -100 -5788 -84 -5754
rect 84 -5788 100 -5754
rect -146 -5884 -112 -5868
rect -146 -6876 -112 -6860
rect 112 -5884 146 -5868
rect 112 -6876 146 -6860
rect -100 -6953 -84 -6919
rect 84 -6953 100 -6919
rect -146 -7049 -112 -7033
rect -146 -8041 -112 -8025
rect 112 -7049 146 -7033
rect 112 -8041 146 -8025
rect -100 -8118 -84 -8084
rect 84 -8118 100 -8084
rect -146 -8214 -112 -8198
rect -146 -9206 -112 -9190
rect 112 -8214 146 -8198
rect 112 -9206 146 -9190
rect -100 -9283 -84 -9249
rect 84 -9283 100 -9249
rect -146 -9379 -112 -9363
rect -146 -10371 -112 -10355
rect 112 -9379 146 -9363
rect 112 -10371 146 -10355
rect -100 -10448 -84 -10414
rect 84 -10448 100 -10414
rect -146 -10544 -112 -10528
rect -146 -11536 -112 -11520
rect 112 -10544 146 -10528
rect 112 -11536 146 -11520
rect -100 -11613 -84 -11579
rect 84 -11613 100 -11579
rect -146 -11709 -112 -11693
rect -146 -12701 -112 -12685
rect 112 -11709 146 -11693
rect 112 -12701 146 -12685
rect -100 -12778 -84 -12744
rect 84 -12778 100 -12744
rect -146 -12874 -112 -12858
rect -146 -13866 -112 -13850
rect 112 -12874 146 -12858
rect 112 -13866 146 -13850
rect -100 -13943 -84 -13909
rect 84 -13943 100 -13909
rect -146 -14039 -112 -14023
rect -146 -15031 -112 -15015
rect 112 -14039 146 -14023
rect 112 -15031 146 -15015
rect -100 -15108 -84 -15074
rect 84 -15108 100 -15074
rect -146 -15204 -112 -15188
rect -146 -16196 -112 -16180
rect 112 -15204 146 -15188
rect 112 -16196 146 -16180
rect -100 -16273 -84 -16239
rect 84 -16273 100 -16239
rect -146 -16369 -112 -16353
rect -146 -17361 -112 -17345
rect 112 -16369 146 -16353
rect 112 -17361 146 -17345
rect -100 -17438 -84 -17404
rect 84 -17438 100 -17404
rect -146 -17534 -112 -17518
rect -146 -18526 -112 -18510
rect 112 -17534 146 -17518
rect 112 -18526 146 -18510
rect -100 -18603 -84 -18569
rect 84 -18603 100 -18569
rect -146 -18699 -112 -18683
rect -146 -19691 -112 -19675
rect 112 -18699 146 -18683
rect 112 -19691 146 -19675
rect -100 -19768 -84 -19734
rect 84 -19768 100 -19734
rect -146 -19864 -112 -19848
rect -146 -20856 -112 -20840
rect 112 -19864 146 -19848
rect 112 -20856 146 -20840
rect -100 -20933 -84 -20899
rect 84 -20933 100 -20899
rect -260 -21001 -226 -20939
rect 226 -21001 260 -20939
rect -260 -21035 -164 -21001
rect 164 -21035 260 -21001
<< viali >>
rect -146 19935 -112 20911
rect 112 19935 146 20911
rect -84 19842 84 19876
rect -146 18770 -112 19746
rect 112 18770 146 19746
rect -84 18677 84 18711
rect -146 17605 -112 18581
rect 112 17605 146 18581
rect -84 17512 84 17546
rect -146 16440 -112 17416
rect 112 16440 146 17416
rect -84 16347 84 16381
rect -146 15275 -112 16251
rect 112 15275 146 16251
rect -84 15182 84 15216
rect -146 14110 -112 15086
rect 112 14110 146 15086
rect -84 14017 84 14051
rect -146 12945 -112 13921
rect 112 12945 146 13921
rect -84 12852 84 12886
rect -146 11780 -112 12756
rect 112 11780 146 12756
rect -84 11687 84 11721
rect -146 10615 -112 11591
rect 112 10615 146 11591
rect -84 10522 84 10556
rect -146 9450 -112 10426
rect 112 9450 146 10426
rect -84 9357 84 9391
rect -146 8285 -112 9261
rect 112 8285 146 9261
rect -84 8192 84 8226
rect -146 7120 -112 8096
rect 112 7120 146 8096
rect -84 7027 84 7061
rect -146 5955 -112 6931
rect 112 5955 146 6931
rect -84 5862 84 5896
rect -146 4790 -112 5766
rect 112 4790 146 5766
rect -84 4697 84 4731
rect -146 3625 -112 4601
rect 112 3625 146 4601
rect -84 3532 84 3566
rect -146 2460 -112 3436
rect 112 2460 146 3436
rect -84 2367 84 2401
rect -146 1295 -112 2271
rect 112 1295 146 2271
rect -84 1202 84 1236
rect -146 130 -112 1106
rect 112 130 146 1106
rect -84 37 84 71
rect -146 -1035 -112 -59
rect 112 -1035 146 -59
rect -84 -1128 84 -1094
rect -146 -2200 -112 -1224
rect 112 -2200 146 -1224
rect -84 -2293 84 -2259
rect -146 -3365 -112 -2389
rect 112 -3365 146 -2389
rect -84 -3458 84 -3424
rect -146 -4530 -112 -3554
rect 112 -4530 146 -3554
rect -84 -4623 84 -4589
rect -146 -5695 -112 -4719
rect 112 -5695 146 -4719
rect -84 -5788 84 -5754
rect -146 -6860 -112 -5884
rect 112 -6860 146 -5884
rect -84 -6953 84 -6919
rect -146 -8025 -112 -7049
rect 112 -8025 146 -7049
rect -84 -8118 84 -8084
rect -146 -9190 -112 -8214
rect 112 -9190 146 -8214
rect -84 -9283 84 -9249
rect -146 -10355 -112 -9379
rect 112 -10355 146 -9379
rect -84 -10448 84 -10414
rect -146 -11520 -112 -10544
rect 112 -11520 146 -10544
rect -84 -11613 84 -11579
rect -146 -12685 -112 -11709
rect 112 -12685 146 -11709
rect -84 -12778 84 -12744
rect -146 -13850 -112 -12874
rect 112 -13850 146 -12874
rect -84 -13943 84 -13909
rect -146 -15015 -112 -14039
rect 112 -15015 146 -14039
rect -84 -15108 84 -15074
rect -146 -16180 -112 -15204
rect 112 -16180 146 -15204
rect -84 -16273 84 -16239
rect -146 -17345 -112 -16369
rect 112 -17345 146 -16369
rect -84 -17438 84 -17404
rect -146 -18510 -112 -17534
rect 112 -18510 146 -17534
rect -84 -18603 84 -18569
rect -146 -19675 -112 -18699
rect 112 -19675 146 -18699
rect -84 -19768 84 -19734
rect -146 -20840 -112 -19864
rect 112 -20840 146 -19864
rect -84 -20933 84 -20899
<< metal1 >>
rect -152 20911 -106 20923
rect -152 19935 -146 20911
rect -112 19935 -106 20911
rect -152 19923 -106 19935
rect 106 20911 152 20923
rect 106 19935 112 20911
rect 146 19935 152 20911
rect 106 19923 152 19935
rect -96 19876 96 19882
rect -96 19842 -84 19876
rect 84 19842 96 19876
rect -96 19836 96 19842
rect -152 19746 -106 19758
rect -152 18770 -146 19746
rect -112 18770 -106 19746
rect -152 18758 -106 18770
rect 106 19746 152 19758
rect 106 18770 112 19746
rect 146 18770 152 19746
rect 106 18758 152 18770
rect -96 18711 96 18717
rect -96 18677 -84 18711
rect 84 18677 96 18711
rect -96 18671 96 18677
rect -152 18581 -106 18593
rect -152 17605 -146 18581
rect -112 17605 -106 18581
rect -152 17593 -106 17605
rect 106 18581 152 18593
rect 106 17605 112 18581
rect 146 17605 152 18581
rect 106 17593 152 17605
rect -96 17546 96 17552
rect -96 17512 -84 17546
rect 84 17512 96 17546
rect -96 17506 96 17512
rect -152 17416 -106 17428
rect -152 16440 -146 17416
rect -112 16440 -106 17416
rect -152 16428 -106 16440
rect 106 17416 152 17428
rect 106 16440 112 17416
rect 146 16440 152 17416
rect 106 16428 152 16440
rect -96 16381 96 16387
rect -96 16347 -84 16381
rect 84 16347 96 16381
rect -96 16341 96 16347
rect -152 16251 -106 16263
rect -152 15275 -146 16251
rect -112 15275 -106 16251
rect -152 15263 -106 15275
rect 106 16251 152 16263
rect 106 15275 112 16251
rect 146 15275 152 16251
rect 106 15263 152 15275
rect -96 15216 96 15222
rect -96 15182 -84 15216
rect 84 15182 96 15216
rect -96 15176 96 15182
rect -152 15086 -106 15098
rect -152 14110 -146 15086
rect -112 14110 -106 15086
rect -152 14098 -106 14110
rect 106 15086 152 15098
rect 106 14110 112 15086
rect 146 14110 152 15086
rect 106 14098 152 14110
rect -96 14051 96 14057
rect -96 14017 -84 14051
rect 84 14017 96 14051
rect -96 14011 96 14017
rect -152 13921 -106 13933
rect -152 12945 -146 13921
rect -112 12945 -106 13921
rect -152 12933 -106 12945
rect 106 13921 152 13933
rect 106 12945 112 13921
rect 146 12945 152 13921
rect 106 12933 152 12945
rect -96 12886 96 12892
rect -96 12852 -84 12886
rect 84 12852 96 12886
rect -96 12846 96 12852
rect -152 12756 -106 12768
rect -152 11780 -146 12756
rect -112 11780 -106 12756
rect -152 11768 -106 11780
rect 106 12756 152 12768
rect 106 11780 112 12756
rect 146 11780 152 12756
rect 106 11768 152 11780
rect -96 11721 96 11727
rect -96 11687 -84 11721
rect 84 11687 96 11721
rect -96 11681 96 11687
rect -152 11591 -106 11603
rect -152 10615 -146 11591
rect -112 10615 -106 11591
rect -152 10603 -106 10615
rect 106 11591 152 11603
rect 106 10615 112 11591
rect 146 10615 152 11591
rect 106 10603 152 10615
rect -96 10556 96 10562
rect -96 10522 -84 10556
rect 84 10522 96 10556
rect -96 10516 96 10522
rect -152 10426 -106 10438
rect -152 9450 -146 10426
rect -112 9450 -106 10426
rect -152 9438 -106 9450
rect 106 10426 152 10438
rect 106 9450 112 10426
rect 146 9450 152 10426
rect 106 9438 152 9450
rect -96 9391 96 9397
rect -96 9357 -84 9391
rect 84 9357 96 9391
rect -96 9351 96 9357
rect -152 9261 -106 9273
rect -152 8285 -146 9261
rect -112 8285 -106 9261
rect -152 8273 -106 8285
rect 106 9261 152 9273
rect 106 8285 112 9261
rect 146 8285 152 9261
rect 106 8273 152 8285
rect -96 8226 96 8232
rect -96 8192 -84 8226
rect 84 8192 96 8226
rect -96 8186 96 8192
rect -152 8096 -106 8108
rect -152 7120 -146 8096
rect -112 7120 -106 8096
rect -152 7108 -106 7120
rect 106 8096 152 8108
rect 106 7120 112 8096
rect 146 7120 152 8096
rect 106 7108 152 7120
rect -96 7061 96 7067
rect -96 7027 -84 7061
rect 84 7027 96 7061
rect -96 7021 96 7027
rect -152 6931 -106 6943
rect -152 5955 -146 6931
rect -112 5955 -106 6931
rect -152 5943 -106 5955
rect 106 6931 152 6943
rect 106 5955 112 6931
rect 146 5955 152 6931
rect 106 5943 152 5955
rect -96 5896 96 5902
rect -96 5862 -84 5896
rect 84 5862 96 5896
rect -96 5856 96 5862
rect -152 5766 -106 5778
rect -152 4790 -146 5766
rect -112 4790 -106 5766
rect -152 4778 -106 4790
rect 106 5766 152 5778
rect 106 4790 112 5766
rect 146 4790 152 5766
rect 106 4778 152 4790
rect -96 4731 96 4737
rect -96 4697 -84 4731
rect 84 4697 96 4731
rect -96 4691 96 4697
rect -152 4601 -106 4613
rect -152 3625 -146 4601
rect -112 3625 -106 4601
rect -152 3613 -106 3625
rect 106 4601 152 4613
rect 106 3625 112 4601
rect 146 3625 152 4601
rect 106 3613 152 3625
rect -96 3566 96 3572
rect -96 3532 -84 3566
rect 84 3532 96 3566
rect -96 3526 96 3532
rect -152 3436 -106 3448
rect -152 2460 -146 3436
rect -112 2460 -106 3436
rect -152 2448 -106 2460
rect 106 3436 152 3448
rect 106 2460 112 3436
rect 146 2460 152 3436
rect 106 2448 152 2460
rect -96 2401 96 2407
rect -96 2367 -84 2401
rect 84 2367 96 2401
rect -96 2361 96 2367
rect -152 2271 -106 2283
rect -152 1295 -146 2271
rect -112 1295 -106 2271
rect -152 1283 -106 1295
rect 106 2271 152 2283
rect 106 1295 112 2271
rect 146 1295 152 2271
rect 106 1283 152 1295
rect -96 1236 96 1242
rect -96 1202 -84 1236
rect 84 1202 96 1236
rect -96 1196 96 1202
rect -152 1106 -106 1118
rect -152 130 -146 1106
rect -112 130 -106 1106
rect -152 118 -106 130
rect 106 1106 152 1118
rect 106 130 112 1106
rect 146 130 152 1106
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -152 -59 -106 -47
rect -152 -1035 -146 -59
rect -112 -1035 -106 -59
rect -152 -1047 -106 -1035
rect 106 -59 152 -47
rect 106 -1035 112 -59
rect 146 -1035 152 -59
rect 106 -1047 152 -1035
rect -96 -1094 96 -1088
rect -96 -1128 -84 -1094
rect 84 -1128 96 -1094
rect -96 -1134 96 -1128
rect -152 -1224 -106 -1212
rect -152 -2200 -146 -1224
rect -112 -2200 -106 -1224
rect -152 -2212 -106 -2200
rect 106 -1224 152 -1212
rect 106 -2200 112 -1224
rect 146 -2200 152 -1224
rect 106 -2212 152 -2200
rect -96 -2259 96 -2253
rect -96 -2293 -84 -2259
rect 84 -2293 96 -2259
rect -96 -2299 96 -2293
rect -152 -2389 -106 -2377
rect -152 -3365 -146 -2389
rect -112 -3365 -106 -2389
rect -152 -3377 -106 -3365
rect 106 -2389 152 -2377
rect 106 -3365 112 -2389
rect 146 -3365 152 -2389
rect 106 -3377 152 -3365
rect -96 -3424 96 -3418
rect -96 -3458 -84 -3424
rect 84 -3458 96 -3424
rect -96 -3464 96 -3458
rect -152 -3554 -106 -3542
rect -152 -4530 -146 -3554
rect -112 -4530 -106 -3554
rect -152 -4542 -106 -4530
rect 106 -3554 152 -3542
rect 106 -4530 112 -3554
rect 146 -4530 152 -3554
rect 106 -4542 152 -4530
rect -96 -4589 96 -4583
rect -96 -4623 -84 -4589
rect 84 -4623 96 -4589
rect -96 -4629 96 -4623
rect -152 -4719 -106 -4707
rect -152 -5695 -146 -4719
rect -112 -5695 -106 -4719
rect -152 -5707 -106 -5695
rect 106 -4719 152 -4707
rect 106 -5695 112 -4719
rect 146 -5695 152 -4719
rect 106 -5707 152 -5695
rect -96 -5754 96 -5748
rect -96 -5788 -84 -5754
rect 84 -5788 96 -5754
rect -96 -5794 96 -5788
rect -152 -5884 -106 -5872
rect -152 -6860 -146 -5884
rect -112 -6860 -106 -5884
rect -152 -6872 -106 -6860
rect 106 -5884 152 -5872
rect 106 -6860 112 -5884
rect 146 -6860 152 -5884
rect 106 -6872 152 -6860
rect -96 -6919 96 -6913
rect -96 -6953 -84 -6919
rect 84 -6953 96 -6919
rect -96 -6959 96 -6953
rect -152 -7049 -106 -7037
rect -152 -8025 -146 -7049
rect -112 -8025 -106 -7049
rect -152 -8037 -106 -8025
rect 106 -7049 152 -7037
rect 106 -8025 112 -7049
rect 146 -8025 152 -7049
rect 106 -8037 152 -8025
rect -96 -8084 96 -8078
rect -96 -8118 -84 -8084
rect 84 -8118 96 -8084
rect -96 -8124 96 -8118
rect -152 -8214 -106 -8202
rect -152 -9190 -146 -8214
rect -112 -9190 -106 -8214
rect -152 -9202 -106 -9190
rect 106 -8214 152 -8202
rect 106 -9190 112 -8214
rect 146 -9190 152 -8214
rect 106 -9202 152 -9190
rect -96 -9249 96 -9243
rect -96 -9283 -84 -9249
rect 84 -9283 96 -9249
rect -96 -9289 96 -9283
rect -152 -9379 -106 -9367
rect -152 -10355 -146 -9379
rect -112 -10355 -106 -9379
rect -152 -10367 -106 -10355
rect 106 -9379 152 -9367
rect 106 -10355 112 -9379
rect 146 -10355 152 -9379
rect 106 -10367 152 -10355
rect -96 -10414 96 -10408
rect -96 -10448 -84 -10414
rect 84 -10448 96 -10414
rect -96 -10454 96 -10448
rect -152 -10544 -106 -10532
rect -152 -11520 -146 -10544
rect -112 -11520 -106 -10544
rect -152 -11532 -106 -11520
rect 106 -10544 152 -10532
rect 106 -11520 112 -10544
rect 146 -11520 152 -10544
rect 106 -11532 152 -11520
rect -96 -11579 96 -11573
rect -96 -11613 -84 -11579
rect 84 -11613 96 -11579
rect -96 -11619 96 -11613
rect -152 -11709 -106 -11697
rect -152 -12685 -146 -11709
rect -112 -12685 -106 -11709
rect -152 -12697 -106 -12685
rect 106 -11709 152 -11697
rect 106 -12685 112 -11709
rect 146 -12685 152 -11709
rect 106 -12697 152 -12685
rect -96 -12744 96 -12738
rect -96 -12778 -84 -12744
rect 84 -12778 96 -12744
rect -96 -12784 96 -12778
rect -152 -12874 -106 -12862
rect -152 -13850 -146 -12874
rect -112 -13850 -106 -12874
rect -152 -13862 -106 -13850
rect 106 -12874 152 -12862
rect 106 -13850 112 -12874
rect 146 -13850 152 -12874
rect 106 -13862 152 -13850
rect -96 -13909 96 -13903
rect -96 -13943 -84 -13909
rect 84 -13943 96 -13909
rect -96 -13949 96 -13943
rect -152 -14039 -106 -14027
rect -152 -15015 -146 -14039
rect -112 -15015 -106 -14039
rect -152 -15027 -106 -15015
rect 106 -14039 152 -14027
rect 106 -15015 112 -14039
rect 146 -15015 152 -14039
rect 106 -15027 152 -15015
rect -96 -15074 96 -15068
rect -96 -15108 -84 -15074
rect 84 -15108 96 -15074
rect -96 -15114 96 -15108
rect -152 -15204 -106 -15192
rect -152 -16180 -146 -15204
rect -112 -16180 -106 -15204
rect -152 -16192 -106 -16180
rect 106 -15204 152 -15192
rect 106 -16180 112 -15204
rect 146 -16180 152 -15204
rect 106 -16192 152 -16180
rect -96 -16239 96 -16233
rect -96 -16273 -84 -16239
rect 84 -16273 96 -16239
rect -96 -16279 96 -16273
rect -152 -16369 -106 -16357
rect -152 -17345 -146 -16369
rect -112 -17345 -106 -16369
rect -152 -17357 -106 -17345
rect 106 -16369 152 -16357
rect 106 -17345 112 -16369
rect 146 -17345 152 -16369
rect 106 -17357 152 -17345
rect -96 -17404 96 -17398
rect -96 -17438 -84 -17404
rect 84 -17438 96 -17404
rect -96 -17444 96 -17438
rect -152 -17534 -106 -17522
rect -152 -18510 -146 -17534
rect -112 -18510 -106 -17534
rect -152 -18522 -106 -18510
rect 106 -17534 152 -17522
rect 106 -18510 112 -17534
rect 146 -18510 152 -17534
rect 106 -18522 152 -18510
rect -96 -18569 96 -18563
rect -96 -18603 -84 -18569
rect 84 -18603 96 -18569
rect -96 -18609 96 -18603
rect -152 -18699 -106 -18687
rect -152 -19675 -146 -18699
rect -112 -19675 -106 -18699
rect -152 -19687 -106 -19675
rect 106 -18699 152 -18687
rect 106 -19675 112 -18699
rect 146 -19675 152 -18699
rect 106 -19687 152 -19675
rect -96 -19734 96 -19728
rect -96 -19768 -84 -19734
rect 84 -19768 96 -19734
rect -96 -19774 96 -19768
rect -152 -19864 -106 -19852
rect -152 -20840 -146 -19864
rect -112 -20840 -106 -19864
rect -152 -20852 -106 -20840
rect 106 -19864 152 -19852
rect 106 -20840 112 -19864
rect 146 -20840 152 -19864
rect 106 -20852 152 -20840
rect -96 -20899 96 -20893
rect -96 -20933 -84 -20899
rect 84 -20933 96 -20899
rect -96 -20939 96 -20933
<< properties >>
string FIXED_BBOX -243 -21018 243 21018
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 1 m 36 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
