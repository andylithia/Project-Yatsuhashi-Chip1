magic
tech sky130A
magscale 1 2
timestamp 1659107442
<< error_p >>
rect 138 92 194 1102
rect 224 92 280 1102
rect 310 92 366 1102
rect 396 92 452 1102
rect 482 92 538 1102
<< pwell >>
rect 100 66 576 1128
<< nmos >>
rect 194 92 224 1102
rect 280 92 310 1102
rect 366 92 396 1102
rect 452 92 482 1102
<< ndiff >>
rect 138 1090 194 1102
rect 138 1056 149 1090
rect 183 1056 194 1090
rect 138 1022 194 1056
rect 138 988 149 1022
rect 183 988 194 1022
rect 138 954 194 988
rect 138 920 149 954
rect 183 920 194 954
rect 138 886 194 920
rect 138 852 149 886
rect 183 852 194 886
rect 138 818 194 852
rect 138 784 149 818
rect 183 784 194 818
rect 138 750 194 784
rect 138 716 149 750
rect 183 716 194 750
rect 138 682 194 716
rect 138 648 149 682
rect 183 648 194 682
rect 138 614 194 648
rect 138 580 149 614
rect 183 580 194 614
rect 138 546 194 580
rect 138 512 149 546
rect 183 512 194 546
rect 138 478 194 512
rect 138 444 149 478
rect 183 444 194 478
rect 138 410 194 444
rect 138 376 149 410
rect 183 376 194 410
rect 138 342 194 376
rect 138 308 149 342
rect 183 308 194 342
rect 138 274 194 308
rect 138 240 149 274
rect 183 240 194 274
rect 138 206 194 240
rect 138 172 149 206
rect 183 172 194 206
rect 138 138 194 172
rect 138 104 149 138
rect 183 104 194 138
rect 138 92 194 104
rect 224 1090 280 1102
rect 224 1056 235 1090
rect 269 1056 280 1090
rect 224 1022 280 1056
rect 224 988 235 1022
rect 269 988 280 1022
rect 224 954 280 988
rect 224 920 235 954
rect 269 920 280 954
rect 224 886 280 920
rect 224 852 235 886
rect 269 852 280 886
rect 224 818 280 852
rect 224 784 235 818
rect 269 784 280 818
rect 224 750 280 784
rect 224 716 235 750
rect 269 716 280 750
rect 224 682 280 716
rect 224 648 235 682
rect 269 648 280 682
rect 224 614 280 648
rect 224 580 235 614
rect 269 580 280 614
rect 224 546 280 580
rect 224 512 235 546
rect 269 512 280 546
rect 224 478 280 512
rect 224 444 235 478
rect 269 444 280 478
rect 224 410 280 444
rect 224 376 235 410
rect 269 376 280 410
rect 224 342 280 376
rect 224 308 235 342
rect 269 308 280 342
rect 224 274 280 308
rect 224 240 235 274
rect 269 240 280 274
rect 224 206 280 240
rect 224 172 235 206
rect 269 172 280 206
rect 224 138 280 172
rect 224 104 235 138
rect 269 104 280 138
rect 224 92 280 104
rect 310 1090 366 1102
rect 310 1056 321 1090
rect 355 1056 366 1090
rect 310 1022 366 1056
rect 310 988 321 1022
rect 355 988 366 1022
rect 310 954 366 988
rect 310 920 321 954
rect 355 920 366 954
rect 310 886 366 920
rect 310 852 321 886
rect 355 852 366 886
rect 310 818 366 852
rect 310 784 321 818
rect 355 784 366 818
rect 310 750 366 784
rect 310 716 321 750
rect 355 716 366 750
rect 310 682 366 716
rect 310 648 321 682
rect 355 648 366 682
rect 310 614 366 648
rect 310 580 321 614
rect 355 580 366 614
rect 310 546 366 580
rect 310 512 321 546
rect 355 512 366 546
rect 310 478 366 512
rect 310 444 321 478
rect 355 444 366 478
rect 310 410 366 444
rect 310 376 321 410
rect 355 376 366 410
rect 310 342 366 376
rect 310 308 321 342
rect 355 308 366 342
rect 310 274 366 308
rect 310 240 321 274
rect 355 240 366 274
rect 310 206 366 240
rect 310 172 321 206
rect 355 172 366 206
rect 310 138 366 172
rect 310 104 321 138
rect 355 104 366 138
rect 310 92 366 104
rect 396 1090 452 1102
rect 396 1056 407 1090
rect 441 1056 452 1090
rect 396 1022 452 1056
rect 396 988 407 1022
rect 441 988 452 1022
rect 396 954 452 988
rect 396 920 407 954
rect 441 920 452 954
rect 396 886 452 920
rect 396 852 407 886
rect 441 852 452 886
rect 396 818 452 852
rect 396 784 407 818
rect 441 784 452 818
rect 396 750 452 784
rect 396 716 407 750
rect 441 716 452 750
rect 396 682 452 716
rect 396 648 407 682
rect 441 648 452 682
rect 396 614 452 648
rect 396 580 407 614
rect 441 580 452 614
rect 396 546 452 580
rect 396 512 407 546
rect 441 512 452 546
rect 396 478 452 512
rect 396 444 407 478
rect 441 444 452 478
rect 396 410 452 444
rect 396 376 407 410
rect 441 376 452 410
rect 396 342 452 376
rect 396 308 407 342
rect 441 308 452 342
rect 396 274 452 308
rect 396 240 407 274
rect 441 240 452 274
rect 396 206 452 240
rect 396 172 407 206
rect 441 172 452 206
rect 396 138 452 172
rect 396 104 407 138
rect 441 104 452 138
rect 396 92 452 104
rect 482 1090 538 1102
rect 482 1056 493 1090
rect 527 1056 538 1090
rect 482 1022 538 1056
rect 482 988 493 1022
rect 527 988 538 1022
rect 482 954 538 988
rect 482 920 493 954
rect 527 920 538 954
rect 482 886 538 920
rect 482 852 493 886
rect 527 852 538 886
rect 482 818 538 852
rect 482 784 493 818
rect 527 784 538 818
rect 482 750 538 784
rect 482 716 493 750
rect 527 716 538 750
rect 482 682 538 716
rect 482 648 493 682
rect 527 648 538 682
rect 482 614 538 648
rect 482 580 493 614
rect 527 580 538 614
rect 482 546 538 580
rect 482 512 493 546
rect 527 512 538 546
rect 482 478 538 512
rect 482 444 493 478
rect 527 444 538 478
rect 482 410 538 444
rect 482 376 493 410
rect 527 376 538 410
rect 482 342 538 376
rect 482 308 493 342
rect 527 308 538 342
rect 482 274 538 308
rect 482 240 493 274
rect 527 240 538 274
rect 482 206 538 240
rect 482 172 493 206
rect 527 172 538 206
rect 482 138 538 172
rect 482 104 493 138
rect 527 104 538 138
rect 482 92 538 104
<< ndiffc >>
rect 149 1056 183 1090
rect 149 988 183 1022
rect 149 920 183 954
rect 149 852 183 886
rect 149 784 183 818
rect 149 716 183 750
rect 149 648 183 682
rect 149 580 183 614
rect 149 512 183 546
rect 149 444 183 478
rect 149 376 183 410
rect 149 308 183 342
rect 149 240 183 274
rect 149 172 183 206
rect 149 104 183 138
rect 235 1056 269 1090
rect 235 988 269 1022
rect 235 920 269 954
rect 235 852 269 886
rect 235 784 269 818
rect 235 716 269 750
rect 235 648 269 682
rect 235 580 269 614
rect 235 512 269 546
rect 235 444 269 478
rect 235 376 269 410
rect 235 308 269 342
rect 235 240 269 274
rect 235 172 269 206
rect 235 104 269 138
rect 321 1056 355 1090
rect 321 988 355 1022
rect 321 920 355 954
rect 321 852 355 886
rect 321 784 355 818
rect 321 716 355 750
rect 321 648 355 682
rect 321 580 355 614
rect 321 512 355 546
rect 321 444 355 478
rect 321 376 355 410
rect 321 308 355 342
rect 321 240 355 274
rect 321 172 355 206
rect 321 104 355 138
rect 407 1056 441 1090
rect 407 988 441 1022
rect 407 920 441 954
rect 407 852 441 886
rect 407 784 441 818
rect 407 716 441 750
rect 407 648 441 682
rect 407 580 441 614
rect 407 512 441 546
rect 407 444 441 478
rect 407 376 441 410
rect 407 308 441 342
rect 407 240 441 274
rect 407 172 441 206
rect 407 104 441 138
rect 493 1056 527 1090
rect 493 988 527 1022
rect 493 920 527 954
rect 493 852 527 886
rect 493 784 527 818
rect 493 716 527 750
rect 493 648 527 682
rect 493 580 527 614
rect 493 512 527 546
rect 493 444 527 478
rect 493 376 527 410
rect 493 308 527 342
rect 493 240 527 274
rect 493 172 527 206
rect 493 104 527 138
<< poly >>
rect 169 1174 528 1194
rect 169 1140 253 1174
rect 287 1140 321 1174
rect 355 1140 389 1174
rect 423 1140 528 1174
rect 169 1124 528 1140
rect 194 1102 224 1124
rect 280 1102 310 1124
rect 366 1102 396 1124
rect 452 1102 482 1124
rect 194 66 224 92
rect 280 66 310 92
rect 366 66 396 92
rect 452 66 482 92
rect 194 36 482 66
<< polycont >>
rect 253 1140 287 1174
rect 321 1140 355 1174
rect 389 1140 423 1174
<< locali >>
rect 169 1140 249 1174
rect 287 1140 321 1174
rect 355 1140 389 1174
rect 427 1140 457 1174
rect 149 1090 183 1106
rect 149 1022 183 1048
rect 149 954 183 976
rect 149 886 183 904
rect 149 818 183 832
rect 149 750 183 760
rect 149 682 183 688
rect 149 614 183 616
rect 149 578 183 580
rect 149 506 183 512
rect 149 434 183 444
rect 149 362 183 376
rect 149 290 183 308
rect 149 218 183 240
rect 149 146 183 172
rect 149 88 183 104
rect 235 1090 269 1106
rect 235 1022 269 1048
rect 235 954 269 976
rect 235 886 269 904
rect 235 818 269 832
rect 235 750 269 760
rect 235 682 269 688
rect 235 614 269 616
rect 235 578 269 580
rect 235 506 269 512
rect 235 434 269 444
rect 235 362 269 376
rect 235 290 269 308
rect 235 218 269 240
rect 235 146 269 172
rect 235 88 269 104
rect 321 1090 355 1106
rect 321 1022 355 1048
rect 321 954 355 976
rect 321 886 355 904
rect 321 818 355 832
rect 321 750 355 760
rect 321 682 355 688
rect 321 614 355 616
rect 321 578 355 580
rect 321 506 355 512
rect 321 434 355 444
rect 321 362 355 376
rect 321 290 355 308
rect 321 218 355 240
rect 321 146 355 172
rect 321 88 355 104
rect 407 1090 441 1106
rect 407 1022 441 1048
rect 407 954 441 976
rect 407 886 441 904
rect 407 818 441 832
rect 407 750 441 760
rect 407 682 441 688
rect 407 614 441 616
rect 407 578 441 580
rect 407 506 441 512
rect 407 434 441 444
rect 407 362 441 376
rect 407 290 441 308
rect 407 218 441 240
rect 407 146 441 172
rect 407 88 441 104
rect 493 1090 527 1106
rect 493 1022 527 1048
rect 493 954 527 976
rect 493 886 527 904
rect 493 818 527 832
rect 493 750 527 760
rect 493 682 527 688
rect 493 614 527 616
rect 493 578 527 580
rect 493 506 527 512
rect 493 434 527 444
rect 493 362 527 376
rect 493 290 527 308
rect 493 218 527 240
rect 493 146 527 172
rect 493 88 527 104
<< viali >>
rect 249 1140 253 1174
rect 253 1140 283 1174
rect 321 1140 355 1174
rect 393 1140 423 1174
rect 423 1140 427 1174
rect 149 1056 183 1082
rect 149 1048 183 1056
rect 149 988 183 1010
rect 149 976 183 988
rect 149 920 183 938
rect 149 904 183 920
rect 149 852 183 866
rect 149 832 183 852
rect 149 784 183 794
rect 149 760 183 784
rect 149 716 183 722
rect 149 688 183 716
rect 149 648 183 650
rect 149 616 183 648
rect 149 546 183 578
rect 149 544 183 546
rect 149 478 183 506
rect 149 472 183 478
rect 149 410 183 434
rect 149 400 183 410
rect 149 342 183 362
rect 149 328 183 342
rect 149 274 183 290
rect 149 256 183 274
rect 149 206 183 218
rect 149 184 183 206
rect 149 138 183 146
rect 149 112 183 138
rect 235 1056 269 1082
rect 235 1048 269 1056
rect 235 988 269 1010
rect 235 976 269 988
rect 235 920 269 938
rect 235 904 269 920
rect 235 852 269 866
rect 235 832 269 852
rect 235 784 269 794
rect 235 760 269 784
rect 235 716 269 722
rect 235 688 269 716
rect 235 648 269 650
rect 235 616 269 648
rect 235 546 269 578
rect 235 544 269 546
rect 235 478 269 506
rect 235 472 269 478
rect 235 410 269 434
rect 235 400 269 410
rect 235 342 269 362
rect 235 328 269 342
rect 235 274 269 290
rect 235 256 269 274
rect 235 206 269 218
rect 235 184 269 206
rect 235 138 269 146
rect 235 112 269 138
rect 321 1056 355 1082
rect 321 1048 355 1056
rect 321 988 355 1010
rect 321 976 355 988
rect 321 920 355 938
rect 321 904 355 920
rect 321 852 355 866
rect 321 832 355 852
rect 321 784 355 794
rect 321 760 355 784
rect 321 716 355 722
rect 321 688 355 716
rect 321 648 355 650
rect 321 616 355 648
rect 321 546 355 578
rect 321 544 355 546
rect 321 478 355 506
rect 321 472 355 478
rect 321 410 355 434
rect 321 400 355 410
rect 321 342 355 362
rect 321 328 355 342
rect 321 274 355 290
rect 321 256 355 274
rect 321 206 355 218
rect 321 184 355 206
rect 321 138 355 146
rect 321 112 355 138
rect 407 1056 441 1082
rect 407 1048 441 1056
rect 407 988 441 1010
rect 407 976 441 988
rect 407 920 441 938
rect 407 904 441 920
rect 407 852 441 866
rect 407 832 441 852
rect 407 784 441 794
rect 407 760 441 784
rect 407 716 441 722
rect 407 688 441 716
rect 407 648 441 650
rect 407 616 441 648
rect 407 546 441 578
rect 407 544 441 546
rect 407 478 441 506
rect 407 472 441 478
rect 407 410 441 434
rect 407 400 441 410
rect 407 342 441 362
rect 407 328 441 342
rect 407 274 441 290
rect 407 256 441 274
rect 407 206 441 218
rect 407 184 441 206
rect 407 138 441 146
rect 407 112 441 138
rect 493 1056 527 1082
rect 493 1048 527 1056
rect 493 988 527 1010
rect 493 976 527 988
rect 493 920 527 938
rect 493 904 527 920
rect 493 852 527 866
rect 493 832 527 852
rect 493 784 527 794
rect 493 760 527 784
rect 493 716 527 722
rect 493 688 527 716
rect 493 648 527 650
rect 493 616 527 648
rect 493 546 527 578
rect 493 544 527 546
rect 493 478 527 506
rect 493 472 527 478
rect 493 410 527 434
rect 493 400 527 410
rect 493 342 527 362
rect 493 328 527 342
rect 493 274 527 290
rect 493 256 527 274
rect 493 206 527 218
rect 493 184 527 206
rect 493 138 527 146
rect 493 112 527 138
<< metal1 >>
rect 165 1174 511 1290
rect 165 1140 249 1174
rect 283 1140 321 1174
rect 355 1140 393 1174
rect 427 1140 511 1174
rect 165 1128 511 1140
rect 140 1082 192 1094
rect 140 1048 149 1082
rect 183 1048 192 1082
rect 140 1010 192 1048
rect 140 976 149 1010
rect 183 976 192 1010
rect 140 938 192 976
rect 140 904 149 938
rect 183 904 192 938
rect 140 866 192 904
rect 140 832 149 866
rect 183 832 192 866
rect 140 794 192 832
rect 140 760 149 794
rect 183 760 192 794
rect 140 722 192 760
rect 140 688 149 722
rect 183 688 192 722
rect 140 650 192 688
rect 140 616 149 650
rect 183 616 192 650
rect 140 578 192 616
rect 140 544 149 578
rect 183 544 192 578
rect 140 506 192 544
rect 140 472 149 506
rect 183 472 192 506
rect 140 434 192 472
rect 140 400 149 434
rect 183 400 192 434
rect 140 362 192 400
rect 140 328 149 362
rect 183 328 192 362
rect 140 290 192 328
rect 140 256 149 290
rect 183 256 192 290
rect 140 218 192 256
rect 140 184 149 218
rect 183 184 192 218
rect 140 146 192 184
rect 140 112 149 146
rect 183 112 192 146
rect 140 10 192 112
rect 226 1082 278 1094
rect 226 1048 235 1082
rect 269 1048 278 1082
rect 226 1022 278 1048
rect 226 942 278 970
rect 226 866 278 890
rect 226 862 235 866
rect 269 862 278 866
rect 226 794 278 810
rect 226 782 235 794
rect 269 782 278 794
rect 226 722 278 730
rect 226 702 235 722
rect 269 702 278 722
rect 226 622 235 650
rect 269 622 278 650
rect 226 544 235 570
rect 269 544 278 570
rect 226 542 278 544
rect 226 472 235 490
rect 269 472 278 490
rect 226 462 278 472
rect 226 400 235 410
rect 269 400 278 410
rect 226 382 278 400
rect 226 328 235 330
rect 269 328 278 330
rect 226 302 278 328
rect 226 222 278 250
rect 226 146 278 170
rect 226 112 235 146
rect 269 112 278 146
rect 226 100 278 112
rect 312 1082 364 1094
rect 312 1048 321 1082
rect 355 1048 364 1082
rect 312 1010 364 1048
rect 312 976 321 1010
rect 355 976 364 1010
rect 312 938 364 976
rect 312 904 321 938
rect 355 904 364 938
rect 312 866 364 904
rect 312 832 321 866
rect 355 832 364 866
rect 312 794 364 832
rect 312 760 321 794
rect 355 760 364 794
rect 312 722 364 760
rect 312 688 321 722
rect 355 688 364 722
rect 312 650 364 688
rect 312 616 321 650
rect 355 616 364 650
rect 312 578 364 616
rect 312 544 321 578
rect 355 544 364 578
rect 312 506 364 544
rect 312 472 321 506
rect 355 472 364 506
rect 312 434 364 472
rect 312 400 321 434
rect 355 400 364 434
rect 312 362 364 400
rect 312 328 321 362
rect 355 328 364 362
rect 312 290 364 328
rect 312 256 321 290
rect 355 256 364 290
rect 312 218 364 256
rect 312 184 321 218
rect 355 184 364 218
rect 312 146 364 184
rect 312 112 321 146
rect 355 112 364 146
rect 312 10 364 112
rect 398 1082 450 1094
rect 398 1048 407 1082
rect 441 1048 450 1082
rect 398 1022 450 1048
rect 398 942 450 970
rect 398 866 450 890
rect 398 862 407 866
rect 441 862 450 866
rect 398 794 450 810
rect 398 782 407 794
rect 441 782 450 794
rect 398 722 450 730
rect 398 702 407 722
rect 441 702 450 722
rect 398 622 407 650
rect 441 622 450 650
rect 398 544 407 570
rect 441 544 450 570
rect 398 542 450 544
rect 398 472 407 490
rect 441 472 450 490
rect 398 462 450 472
rect 398 400 407 410
rect 441 400 450 410
rect 398 382 450 400
rect 398 328 407 330
rect 441 328 450 330
rect 398 302 450 328
rect 398 222 450 250
rect 398 146 450 170
rect 398 112 407 146
rect 441 112 450 146
rect 398 100 450 112
rect 484 1082 536 1094
rect 484 1048 493 1082
rect 527 1048 536 1082
rect 484 1010 536 1048
rect 484 976 493 1010
rect 527 976 536 1010
rect 484 938 536 976
rect 484 904 493 938
rect 527 904 536 938
rect 484 866 536 904
rect 484 832 493 866
rect 527 832 536 866
rect 484 794 536 832
rect 484 760 493 794
rect 527 760 536 794
rect 484 722 536 760
rect 484 688 493 722
rect 527 688 536 722
rect 484 650 536 688
rect 484 616 493 650
rect 527 616 536 650
rect 484 578 536 616
rect 484 544 493 578
rect 527 544 536 578
rect 484 506 536 544
rect 484 472 493 506
rect 527 472 536 506
rect 484 434 536 472
rect 484 400 493 434
rect 527 400 536 434
rect 484 362 536 400
rect 484 328 493 362
rect 527 328 536 362
rect 484 290 536 328
rect 484 256 493 290
rect 527 256 536 290
rect 484 218 536 256
rect 484 184 493 218
rect 527 184 536 218
rect 484 146 536 184
rect 484 112 493 146
rect 527 112 536 146
rect 484 10 536 112
rect 140 -40 536 10
<< via1 >>
rect 226 1010 278 1022
rect 226 976 235 1010
rect 235 976 269 1010
rect 269 976 278 1010
rect 226 970 278 976
rect 226 938 278 942
rect 226 904 235 938
rect 235 904 269 938
rect 269 904 278 938
rect 226 890 278 904
rect 226 832 235 862
rect 235 832 269 862
rect 269 832 278 862
rect 226 810 278 832
rect 226 760 235 782
rect 235 760 269 782
rect 269 760 278 782
rect 226 730 278 760
rect 226 688 235 702
rect 235 688 269 702
rect 269 688 278 702
rect 226 650 278 688
rect 226 616 235 622
rect 235 616 269 622
rect 269 616 278 622
rect 226 578 278 616
rect 226 570 235 578
rect 235 570 269 578
rect 269 570 278 578
rect 226 506 278 542
rect 226 490 235 506
rect 235 490 269 506
rect 269 490 278 506
rect 226 434 278 462
rect 226 410 235 434
rect 235 410 269 434
rect 269 410 278 434
rect 226 362 278 382
rect 226 330 235 362
rect 235 330 269 362
rect 269 330 278 362
rect 226 290 278 302
rect 226 256 235 290
rect 235 256 269 290
rect 269 256 278 290
rect 226 250 278 256
rect 226 218 278 222
rect 226 184 235 218
rect 235 184 269 218
rect 269 184 278 218
rect 226 170 278 184
rect 398 1010 450 1022
rect 398 976 407 1010
rect 407 976 441 1010
rect 441 976 450 1010
rect 398 970 450 976
rect 398 938 450 942
rect 398 904 407 938
rect 407 904 441 938
rect 441 904 450 938
rect 398 890 450 904
rect 398 832 407 862
rect 407 832 441 862
rect 441 832 450 862
rect 398 810 450 832
rect 398 760 407 782
rect 407 760 441 782
rect 441 760 450 782
rect 398 730 450 760
rect 398 688 407 702
rect 407 688 441 702
rect 441 688 450 702
rect 398 650 450 688
rect 398 616 407 622
rect 407 616 441 622
rect 441 616 450 622
rect 398 578 450 616
rect 398 570 407 578
rect 407 570 441 578
rect 441 570 450 578
rect 398 506 450 542
rect 398 490 407 506
rect 407 490 441 506
rect 441 490 450 506
rect 398 434 450 462
rect 398 410 407 434
rect 407 410 441 434
rect 441 410 450 434
rect 398 362 450 382
rect 398 330 407 362
rect 407 330 441 362
rect 441 330 450 362
rect 398 290 450 302
rect 398 256 407 290
rect 407 256 441 290
rect 441 256 450 290
rect 398 250 450 256
rect 398 218 450 222
rect 398 184 407 218
rect 407 184 441 218
rect 441 184 450 218
rect 398 170 450 184
<< metal2 >>
rect 160 1130 540 1210
rect 226 1022 278 1130
rect 226 942 278 970
rect 226 862 278 890
rect 226 782 278 810
rect 226 702 278 730
rect 226 622 278 650
rect 226 542 278 570
rect 226 462 278 490
rect 226 382 278 410
rect 226 302 278 330
rect 226 222 278 250
rect 226 100 278 170
rect 398 1022 450 1130
rect 398 942 450 970
rect 398 862 450 890
rect 398 782 450 810
rect 398 702 450 730
rect 398 622 450 650
rect 398 542 450 570
rect 398 462 450 490
rect 398 382 450 410
rect 398 302 450 330
rect 398 222 450 250
rect 398 100 450 170
<< labels >>
rlabel metal1 165 1260 511 1290 1 G
rlabel metal1 139 -41 536 11 1 D
rlabel metal2 160 1130 190 1210 1 S
<< end >>
