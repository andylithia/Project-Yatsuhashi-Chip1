magic
tech sky130A
magscale 1 2
timestamp 1658692977
<< metal1 >>
rect -2771 3169 -1406 3228
rect -2771 2834 -2575 3169
rect -1350 2950 -1250 3050
rect -2771 2620 -1406 2834
rect -2771 2284 -2575 2620
rect -1350 2400 -1250 2500
rect -2771 2070 -1306 2284
rect -2771 1734 -2476 2070
rect -1250 1850 -1150 1950
rect -2771 1520 -1306 1734
rect -2771 1184 -2575 1520
rect -1350 1300 -1250 1400
rect -2771 1126 -2358 1184
rect -2771 1125 -2575 1126
rect -2771 1124 -2631 1125
<< metal2 >>
rect -1850 2200 -1450 3250
rect -1750 1600 -1350 2200
rect -1850 1000 -1450 1600
<< via2 >>
rect -2050 2950 -1950 3200
rect -2050 2250 -1950 2600
rect -1950 1750 -1850 2050
rect -2050 1150 -1950 1450
<< metal3 >>
rect -3300 3250 -2100 3300
rect -3300 3200 -1900 3250
rect -3300 2950 -2050 3200
rect -1950 2950 -1900 3200
rect -3300 2900 -1900 2950
rect -3300 2650 -2100 2800
rect -3300 2600 -1900 2650
rect -1500 2600 -300 3300
rect -3300 2250 -2050 2600
rect -1950 2250 -1900 2600
rect -3300 2200 -1900 2250
rect -1750 2300 -300 2600
rect -1750 2100 -1500 2300
rect -3300 1500 -2100 2100
rect -2000 2050 -300 2100
rect -2000 1750 -1950 2050
rect -1850 1750 -300 2050
rect -2000 1700 -300 1750
rect -3300 1450 -1900 1500
rect -3300 1150 -2050 1450
rect -1950 1150 -1900 1450
rect -3300 1100 -1900 1150
rect -1500 1100 -300 1700
<< mimcap >>
rect -3200 3160 -2200 3200
rect -3200 3040 -3160 3160
rect -2240 3040 -2200 3160
rect -3200 3000 -2200 3040
rect -1400 3160 -400 3200
rect -3200 2660 -2200 2700
rect -3200 2340 -3160 2660
rect -2240 2340 -2200 2660
rect -1400 2440 -1360 3160
rect -440 2440 -400 3160
rect -1400 2400 -400 2440
rect -3200 2300 -2200 2340
rect -3200 1960 -2200 2000
rect -3200 1240 -3160 1960
rect -2240 1240 -2200 1960
rect -3200 1200 -2200 1240
rect -1400 1960 -400 2000
rect -1400 1240 -1360 1960
rect -440 1240 -400 1960
rect -1400 1200 -400 1240
<< mimcapcontact >>
rect -3160 3040 -2240 3160
rect -3160 2340 -2240 2660
rect -1360 2440 -440 3160
rect -3160 1240 -2240 1960
rect -1360 1240 -440 1960
<< metal4 >>
rect -3300 3200 -2100 3300
rect -2000 3250 -1600 3400
rect -2000 3200 -1850 3250
rect -3300 3160 -1850 3200
rect -3300 3040 -3160 3160
rect -2240 3040 -1850 3160
rect -3300 3000 -1850 3040
rect -3300 2900 -2100 3000
rect -3200 2800 -3050 2900
rect -3300 2700 -2100 2800
rect -2000 2700 -1850 3000
rect -3300 2660 -1850 2700
rect -3300 2340 -3160 2660
rect -2240 2340 -1850 2660
rect -3300 2300 -1850 2340
rect -3300 2200 -2100 2300
rect -3200 2100 -3050 2200
rect -3300 2000 -2100 2100
rect -2000 2000 -1850 2300
rect -3300 1960 -1850 2000
rect -3300 1240 -3160 1960
rect -2240 1600 -1850 1960
rect -1750 3100 -1600 3250
rect -1500 3160 -300 3300
rect -1500 3100 -1360 3160
rect -1750 2500 -1360 3100
rect -1750 2000 -1600 2500
rect -1500 2440 -1360 2500
rect -440 2440 -300 3160
rect -1500 2300 -300 2440
rect -550 2100 -400 2300
rect -1500 2000 -300 2100
rect -1750 1960 -300 2000
rect -1750 1600 -1360 1960
rect -2240 1240 -2100 1600
rect -3300 1100 -2100 1240
rect -1500 1240 -1360 1600
rect -440 1240 -300 1960
rect -1500 1100 -300 1240
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1649977179
transform 0 1 -2510 -1 0 3264
box 10 10 514 1204
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1
timestamp 1649977179
transform 0 1 -2510 -1 0 2714
box 10 10 514 1204
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2
timestamp 1649977179
transform 0 1 -2410 -1 0 2164
box 10 10 514 1204
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3
timestamp 1649977179
transform 0 1 -2510 -1 0 1614
box 10 10 514 1204
<< labels >>
rlabel metal2 -1850 1000 -1450 1100 1 bot
rlabel metal4 -2000 3300 -1600 3400 1 top
rlabel metal1 -2771 1124 -2631 3228 1 sub
rlabel mimcapcontact -1350 2950 -1250 3050 1 D0
rlabel metal3 -1350 2400 -1250 2500 1 D1
rlabel mimcapcontact -1250 1850 -1150 1950 1 D3
rlabel mimcapcontact -1350 1300 -1250 1400 1 D2
<< end >>
