magic
tech sky130B
magscale 1 2
timestamp 1659838778
<< error_p >>
rect -3864 181 -3806 187
rect -3746 181 -3688 187
rect -3628 181 -3570 187
rect -3510 181 -3452 187
rect -3392 181 -3334 187
rect -3274 181 -3216 187
rect -3156 181 -3098 187
rect -3038 181 -2980 187
rect -2920 181 -2862 187
rect -2802 181 -2744 187
rect -2684 181 -2626 187
rect -2566 181 -2508 187
rect -2448 181 -2390 187
rect -2330 181 -2272 187
rect -2212 181 -2154 187
rect -2094 181 -2036 187
rect -1976 181 -1918 187
rect -1858 181 -1800 187
rect -1740 181 -1682 187
rect -1622 181 -1564 187
rect -1504 181 -1446 187
rect -1386 181 -1328 187
rect -1268 181 -1210 187
rect -1150 181 -1092 187
rect -1032 181 -974 187
rect -914 181 -856 187
rect -796 181 -738 187
rect -678 181 -620 187
rect -560 181 -502 187
rect -442 181 -384 187
rect -324 181 -266 187
rect -206 181 -148 187
rect -88 181 -30 187
rect 30 181 88 187
rect 148 181 206 187
rect 266 181 324 187
rect 384 181 442 187
rect 502 181 560 187
rect 620 181 678 187
rect 738 181 796 187
rect 856 181 914 187
rect 974 181 1032 187
rect 1092 181 1150 187
rect 1210 181 1268 187
rect 1328 181 1386 187
rect 1446 181 1504 187
rect 1564 181 1622 187
rect 1682 181 1740 187
rect 1800 181 1858 187
rect 1918 181 1976 187
rect 2036 181 2094 187
rect 2154 181 2212 187
rect 2272 181 2330 187
rect 2390 181 2448 187
rect 2508 181 2566 187
rect 2626 181 2684 187
rect 2744 181 2802 187
rect 2862 181 2920 187
rect 2980 181 3038 187
rect 3098 181 3156 187
rect 3216 181 3274 187
rect 3334 181 3392 187
rect 3452 181 3510 187
rect 3570 181 3628 187
rect 3688 181 3746 187
rect 3806 181 3864 187
rect -3864 147 -3852 181
rect -3746 147 -3734 181
rect -3628 147 -3616 181
rect -3510 147 -3498 181
rect -3392 147 -3380 181
rect -3274 147 -3262 181
rect -3156 147 -3144 181
rect -3038 147 -3026 181
rect -2920 147 -2908 181
rect -2802 147 -2790 181
rect -2684 147 -2672 181
rect -2566 147 -2554 181
rect -2448 147 -2436 181
rect -2330 147 -2318 181
rect -2212 147 -2200 181
rect -2094 147 -2082 181
rect -1976 147 -1964 181
rect -1858 147 -1846 181
rect -1740 147 -1728 181
rect -1622 147 -1610 181
rect -1504 147 -1492 181
rect -1386 147 -1374 181
rect -1268 147 -1256 181
rect -1150 147 -1138 181
rect -1032 147 -1020 181
rect -914 147 -902 181
rect -796 147 -784 181
rect -678 147 -666 181
rect -560 147 -548 181
rect -442 147 -430 181
rect -324 147 -312 181
rect -206 147 -194 181
rect -88 147 -76 181
rect 30 147 42 181
rect 148 147 160 181
rect 266 147 278 181
rect 384 147 396 181
rect 502 147 514 181
rect 620 147 632 181
rect 738 147 750 181
rect 856 147 868 181
rect 974 147 986 181
rect 1092 147 1104 181
rect 1210 147 1222 181
rect 1328 147 1340 181
rect 1446 147 1458 181
rect 1564 147 1576 181
rect 1682 147 1694 181
rect 1800 147 1812 181
rect 1918 147 1930 181
rect 2036 147 2048 181
rect 2154 147 2166 181
rect 2272 147 2284 181
rect 2390 147 2402 181
rect 2508 147 2520 181
rect 2626 147 2638 181
rect 2744 147 2756 181
rect 2862 147 2874 181
rect 2980 147 2992 181
rect 3098 147 3110 181
rect 3216 147 3228 181
rect 3334 147 3346 181
rect 3452 147 3464 181
rect 3570 147 3582 181
rect 3688 147 3700 181
rect 3806 147 3818 181
rect -3864 141 -3806 147
rect -3746 141 -3688 147
rect -3628 141 -3570 147
rect -3510 141 -3452 147
rect -3392 141 -3334 147
rect -3274 141 -3216 147
rect -3156 141 -3098 147
rect -3038 141 -2980 147
rect -2920 141 -2862 147
rect -2802 141 -2744 147
rect -2684 141 -2626 147
rect -2566 141 -2508 147
rect -2448 141 -2390 147
rect -2330 141 -2272 147
rect -2212 141 -2154 147
rect -2094 141 -2036 147
rect -1976 141 -1918 147
rect -1858 141 -1800 147
rect -1740 141 -1682 147
rect -1622 141 -1564 147
rect -1504 141 -1446 147
rect -1386 141 -1328 147
rect -1268 141 -1210 147
rect -1150 141 -1092 147
rect -1032 141 -974 147
rect -914 141 -856 147
rect -796 141 -738 147
rect -678 141 -620 147
rect -560 141 -502 147
rect -442 141 -384 147
rect -324 141 -266 147
rect -206 141 -148 147
rect -88 141 -30 147
rect 30 141 88 147
rect 148 141 206 147
rect 266 141 324 147
rect 384 141 442 147
rect 502 141 560 147
rect 620 141 678 147
rect 738 141 796 147
rect 856 141 914 147
rect 974 141 1032 147
rect 1092 141 1150 147
rect 1210 141 1268 147
rect 1328 141 1386 147
rect 1446 141 1504 147
rect 1564 141 1622 147
rect 1682 141 1740 147
rect 1800 141 1858 147
rect 1918 141 1976 147
rect 2036 141 2094 147
rect 2154 141 2212 147
rect 2272 141 2330 147
rect 2390 141 2448 147
rect 2508 141 2566 147
rect 2626 141 2684 147
rect 2744 141 2802 147
rect 2862 141 2920 147
rect 2980 141 3038 147
rect 3098 141 3156 147
rect 3216 141 3274 147
rect 3334 141 3392 147
rect 3452 141 3510 147
rect 3570 141 3628 147
rect 3688 141 3746 147
rect 3806 141 3864 147
rect -3864 -147 -3806 -141
rect -3746 -147 -3688 -141
rect -3628 -147 -3570 -141
rect -3510 -147 -3452 -141
rect -3392 -147 -3334 -141
rect -3274 -147 -3216 -141
rect -3156 -147 -3098 -141
rect -3038 -147 -2980 -141
rect -2920 -147 -2862 -141
rect -2802 -147 -2744 -141
rect -2684 -147 -2626 -141
rect -2566 -147 -2508 -141
rect -2448 -147 -2390 -141
rect -2330 -147 -2272 -141
rect -2212 -147 -2154 -141
rect -2094 -147 -2036 -141
rect -1976 -147 -1918 -141
rect -1858 -147 -1800 -141
rect -1740 -147 -1682 -141
rect -1622 -147 -1564 -141
rect -1504 -147 -1446 -141
rect -1386 -147 -1328 -141
rect -1268 -147 -1210 -141
rect -1150 -147 -1092 -141
rect -1032 -147 -974 -141
rect -914 -147 -856 -141
rect -796 -147 -738 -141
rect -678 -147 -620 -141
rect -560 -147 -502 -141
rect -442 -147 -384 -141
rect -324 -147 -266 -141
rect -206 -147 -148 -141
rect -88 -147 -30 -141
rect 30 -147 88 -141
rect 148 -147 206 -141
rect 266 -147 324 -141
rect 384 -147 442 -141
rect 502 -147 560 -141
rect 620 -147 678 -141
rect 738 -147 796 -141
rect 856 -147 914 -141
rect 974 -147 1032 -141
rect 1092 -147 1150 -141
rect 1210 -147 1268 -141
rect 1328 -147 1386 -141
rect 1446 -147 1504 -141
rect 1564 -147 1622 -141
rect 1682 -147 1740 -141
rect 1800 -147 1858 -141
rect 1918 -147 1976 -141
rect 2036 -147 2094 -141
rect 2154 -147 2212 -141
rect 2272 -147 2330 -141
rect 2390 -147 2448 -141
rect 2508 -147 2566 -141
rect 2626 -147 2684 -141
rect 2744 -147 2802 -141
rect 2862 -147 2920 -141
rect 2980 -147 3038 -141
rect 3098 -147 3156 -141
rect 3216 -147 3274 -141
rect 3334 -147 3392 -141
rect 3452 -147 3510 -141
rect 3570 -147 3628 -141
rect 3688 -147 3746 -141
rect 3806 -147 3864 -141
rect -3864 -181 -3852 -147
rect -3746 -181 -3734 -147
rect -3628 -181 -3616 -147
rect -3510 -181 -3498 -147
rect -3392 -181 -3380 -147
rect -3274 -181 -3262 -147
rect -3156 -181 -3144 -147
rect -3038 -181 -3026 -147
rect -2920 -181 -2908 -147
rect -2802 -181 -2790 -147
rect -2684 -181 -2672 -147
rect -2566 -181 -2554 -147
rect -2448 -181 -2436 -147
rect -2330 -181 -2318 -147
rect -2212 -181 -2200 -147
rect -2094 -181 -2082 -147
rect -1976 -181 -1964 -147
rect -1858 -181 -1846 -147
rect -1740 -181 -1728 -147
rect -1622 -181 -1610 -147
rect -1504 -181 -1492 -147
rect -1386 -181 -1374 -147
rect -1268 -181 -1256 -147
rect -1150 -181 -1138 -147
rect -1032 -181 -1020 -147
rect -914 -181 -902 -147
rect -796 -181 -784 -147
rect -678 -181 -666 -147
rect -560 -181 -548 -147
rect -442 -181 -430 -147
rect -324 -181 -312 -147
rect -206 -181 -194 -147
rect -88 -181 -76 -147
rect 30 -181 42 -147
rect 148 -181 160 -147
rect 266 -181 278 -147
rect 384 -181 396 -147
rect 502 -181 514 -147
rect 620 -181 632 -147
rect 738 -181 750 -147
rect 856 -181 868 -147
rect 974 -181 986 -147
rect 1092 -181 1104 -147
rect 1210 -181 1222 -147
rect 1328 -181 1340 -147
rect 1446 -181 1458 -147
rect 1564 -181 1576 -147
rect 1682 -181 1694 -147
rect 1800 -181 1812 -147
rect 1918 -181 1930 -147
rect 2036 -181 2048 -147
rect 2154 -181 2166 -147
rect 2272 -181 2284 -147
rect 2390 -181 2402 -147
rect 2508 -181 2520 -147
rect 2626 -181 2638 -147
rect 2744 -181 2756 -147
rect 2862 -181 2874 -147
rect 2980 -181 2992 -147
rect 3098 -181 3110 -147
rect 3216 -181 3228 -147
rect 3334 -181 3346 -147
rect 3452 -181 3464 -147
rect 3570 -181 3582 -147
rect 3688 -181 3700 -147
rect 3806 -181 3818 -147
rect -3864 -187 -3806 -181
rect -3746 -187 -3688 -181
rect -3628 -187 -3570 -181
rect -3510 -187 -3452 -181
rect -3392 -187 -3334 -181
rect -3274 -187 -3216 -181
rect -3156 -187 -3098 -181
rect -3038 -187 -2980 -181
rect -2920 -187 -2862 -181
rect -2802 -187 -2744 -181
rect -2684 -187 -2626 -181
rect -2566 -187 -2508 -181
rect -2448 -187 -2390 -181
rect -2330 -187 -2272 -181
rect -2212 -187 -2154 -181
rect -2094 -187 -2036 -181
rect -1976 -187 -1918 -181
rect -1858 -187 -1800 -181
rect -1740 -187 -1682 -181
rect -1622 -187 -1564 -181
rect -1504 -187 -1446 -181
rect -1386 -187 -1328 -181
rect -1268 -187 -1210 -181
rect -1150 -187 -1092 -181
rect -1032 -187 -974 -181
rect -914 -187 -856 -181
rect -796 -187 -738 -181
rect -678 -187 -620 -181
rect -560 -187 -502 -181
rect -442 -187 -384 -181
rect -324 -187 -266 -181
rect -206 -187 -148 -181
rect -88 -187 -30 -181
rect 30 -187 88 -181
rect 148 -187 206 -181
rect 266 -187 324 -181
rect 384 -187 442 -181
rect 502 -187 560 -181
rect 620 -187 678 -181
rect 738 -187 796 -181
rect 856 -187 914 -181
rect 974 -187 1032 -181
rect 1092 -187 1150 -181
rect 1210 -187 1268 -181
rect 1328 -187 1386 -181
rect 1446 -187 1504 -181
rect 1564 -187 1622 -181
rect 1682 -187 1740 -181
rect 1800 -187 1858 -181
rect 1918 -187 1976 -181
rect 2036 -187 2094 -181
rect 2154 -187 2212 -181
rect 2272 -187 2330 -181
rect 2390 -187 2448 -181
rect 2508 -187 2566 -181
rect 2626 -187 2684 -181
rect 2744 -187 2802 -181
rect 2862 -187 2920 -181
rect 2980 -187 3038 -181
rect 3098 -187 3156 -181
rect 3216 -187 3274 -181
rect 3334 -187 3392 -181
rect 3452 -187 3510 -181
rect 3570 -187 3628 -181
rect 3688 -187 3746 -181
rect 3806 -187 3864 -181
<< nwell >>
rect -4061 -319 4061 319
<< pmos >>
rect -3865 -100 -3805 100
rect -3747 -100 -3687 100
rect -3629 -100 -3569 100
rect -3511 -100 -3451 100
rect -3393 -100 -3333 100
rect -3275 -100 -3215 100
rect -3157 -100 -3097 100
rect -3039 -100 -2979 100
rect -2921 -100 -2861 100
rect -2803 -100 -2743 100
rect -2685 -100 -2625 100
rect -2567 -100 -2507 100
rect -2449 -100 -2389 100
rect -2331 -100 -2271 100
rect -2213 -100 -2153 100
rect -2095 -100 -2035 100
rect -1977 -100 -1917 100
rect -1859 -100 -1799 100
rect -1741 -100 -1681 100
rect -1623 -100 -1563 100
rect -1505 -100 -1445 100
rect -1387 -100 -1327 100
rect -1269 -100 -1209 100
rect -1151 -100 -1091 100
rect -1033 -100 -973 100
rect -915 -100 -855 100
rect -797 -100 -737 100
rect -679 -100 -619 100
rect -561 -100 -501 100
rect -443 -100 -383 100
rect -325 -100 -265 100
rect -207 -100 -147 100
rect -89 -100 -29 100
rect 29 -100 89 100
rect 147 -100 207 100
rect 265 -100 325 100
rect 383 -100 443 100
rect 501 -100 561 100
rect 619 -100 679 100
rect 737 -100 797 100
rect 855 -100 915 100
rect 973 -100 1033 100
rect 1091 -100 1151 100
rect 1209 -100 1269 100
rect 1327 -100 1387 100
rect 1445 -100 1505 100
rect 1563 -100 1623 100
rect 1681 -100 1741 100
rect 1799 -100 1859 100
rect 1917 -100 1977 100
rect 2035 -100 2095 100
rect 2153 -100 2213 100
rect 2271 -100 2331 100
rect 2389 -100 2449 100
rect 2507 -100 2567 100
rect 2625 -100 2685 100
rect 2743 -100 2803 100
rect 2861 -100 2921 100
rect 2979 -100 3039 100
rect 3097 -100 3157 100
rect 3215 -100 3275 100
rect 3333 -100 3393 100
rect 3451 -100 3511 100
rect 3569 -100 3629 100
rect 3687 -100 3747 100
rect 3805 -100 3865 100
<< pdiff >>
rect -3923 88 -3865 100
rect -3923 -88 -3911 88
rect -3877 -88 -3865 88
rect -3923 -100 -3865 -88
rect -3805 88 -3747 100
rect -3805 -88 -3793 88
rect -3759 -88 -3747 88
rect -3805 -100 -3747 -88
rect -3687 88 -3629 100
rect -3687 -88 -3675 88
rect -3641 -88 -3629 88
rect -3687 -100 -3629 -88
rect -3569 88 -3511 100
rect -3569 -88 -3557 88
rect -3523 -88 -3511 88
rect -3569 -100 -3511 -88
rect -3451 88 -3393 100
rect -3451 -88 -3439 88
rect -3405 -88 -3393 88
rect -3451 -100 -3393 -88
rect -3333 88 -3275 100
rect -3333 -88 -3321 88
rect -3287 -88 -3275 88
rect -3333 -100 -3275 -88
rect -3215 88 -3157 100
rect -3215 -88 -3203 88
rect -3169 -88 -3157 88
rect -3215 -100 -3157 -88
rect -3097 88 -3039 100
rect -3097 -88 -3085 88
rect -3051 -88 -3039 88
rect -3097 -100 -3039 -88
rect -2979 88 -2921 100
rect -2979 -88 -2967 88
rect -2933 -88 -2921 88
rect -2979 -100 -2921 -88
rect -2861 88 -2803 100
rect -2861 -88 -2849 88
rect -2815 -88 -2803 88
rect -2861 -100 -2803 -88
rect -2743 88 -2685 100
rect -2743 -88 -2731 88
rect -2697 -88 -2685 88
rect -2743 -100 -2685 -88
rect -2625 88 -2567 100
rect -2625 -88 -2613 88
rect -2579 -88 -2567 88
rect -2625 -100 -2567 -88
rect -2507 88 -2449 100
rect -2507 -88 -2495 88
rect -2461 -88 -2449 88
rect -2507 -100 -2449 -88
rect -2389 88 -2331 100
rect -2389 -88 -2377 88
rect -2343 -88 -2331 88
rect -2389 -100 -2331 -88
rect -2271 88 -2213 100
rect -2271 -88 -2259 88
rect -2225 -88 -2213 88
rect -2271 -100 -2213 -88
rect -2153 88 -2095 100
rect -2153 -88 -2141 88
rect -2107 -88 -2095 88
rect -2153 -100 -2095 -88
rect -2035 88 -1977 100
rect -2035 -88 -2023 88
rect -1989 -88 -1977 88
rect -2035 -100 -1977 -88
rect -1917 88 -1859 100
rect -1917 -88 -1905 88
rect -1871 -88 -1859 88
rect -1917 -100 -1859 -88
rect -1799 88 -1741 100
rect -1799 -88 -1787 88
rect -1753 -88 -1741 88
rect -1799 -100 -1741 -88
rect -1681 88 -1623 100
rect -1681 -88 -1669 88
rect -1635 -88 -1623 88
rect -1681 -100 -1623 -88
rect -1563 88 -1505 100
rect -1563 -88 -1551 88
rect -1517 -88 -1505 88
rect -1563 -100 -1505 -88
rect -1445 88 -1387 100
rect -1445 -88 -1433 88
rect -1399 -88 -1387 88
rect -1445 -100 -1387 -88
rect -1327 88 -1269 100
rect -1327 -88 -1315 88
rect -1281 -88 -1269 88
rect -1327 -100 -1269 -88
rect -1209 88 -1151 100
rect -1209 -88 -1197 88
rect -1163 -88 -1151 88
rect -1209 -100 -1151 -88
rect -1091 88 -1033 100
rect -1091 -88 -1079 88
rect -1045 -88 -1033 88
rect -1091 -100 -1033 -88
rect -973 88 -915 100
rect -973 -88 -961 88
rect -927 -88 -915 88
rect -973 -100 -915 -88
rect -855 88 -797 100
rect -855 -88 -843 88
rect -809 -88 -797 88
rect -855 -100 -797 -88
rect -737 88 -679 100
rect -737 -88 -725 88
rect -691 -88 -679 88
rect -737 -100 -679 -88
rect -619 88 -561 100
rect -619 -88 -607 88
rect -573 -88 -561 88
rect -619 -100 -561 -88
rect -501 88 -443 100
rect -501 -88 -489 88
rect -455 -88 -443 88
rect -501 -100 -443 -88
rect -383 88 -325 100
rect -383 -88 -371 88
rect -337 -88 -325 88
rect -383 -100 -325 -88
rect -265 88 -207 100
rect -265 -88 -253 88
rect -219 -88 -207 88
rect -265 -100 -207 -88
rect -147 88 -89 100
rect -147 -88 -135 88
rect -101 -88 -89 88
rect -147 -100 -89 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 89 88 147 100
rect 89 -88 101 88
rect 135 -88 147 88
rect 89 -100 147 -88
rect 207 88 265 100
rect 207 -88 219 88
rect 253 -88 265 88
rect 207 -100 265 -88
rect 325 88 383 100
rect 325 -88 337 88
rect 371 -88 383 88
rect 325 -100 383 -88
rect 443 88 501 100
rect 443 -88 455 88
rect 489 -88 501 88
rect 443 -100 501 -88
rect 561 88 619 100
rect 561 -88 573 88
rect 607 -88 619 88
rect 561 -100 619 -88
rect 679 88 737 100
rect 679 -88 691 88
rect 725 -88 737 88
rect 679 -100 737 -88
rect 797 88 855 100
rect 797 -88 809 88
rect 843 -88 855 88
rect 797 -100 855 -88
rect 915 88 973 100
rect 915 -88 927 88
rect 961 -88 973 88
rect 915 -100 973 -88
rect 1033 88 1091 100
rect 1033 -88 1045 88
rect 1079 -88 1091 88
rect 1033 -100 1091 -88
rect 1151 88 1209 100
rect 1151 -88 1163 88
rect 1197 -88 1209 88
rect 1151 -100 1209 -88
rect 1269 88 1327 100
rect 1269 -88 1281 88
rect 1315 -88 1327 88
rect 1269 -100 1327 -88
rect 1387 88 1445 100
rect 1387 -88 1399 88
rect 1433 -88 1445 88
rect 1387 -100 1445 -88
rect 1505 88 1563 100
rect 1505 -88 1517 88
rect 1551 -88 1563 88
rect 1505 -100 1563 -88
rect 1623 88 1681 100
rect 1623 -88 1635 88
rect 1669 -88 1681 88
rect 1623 -100 1681 -88
rect 1741 88 1799 100
rect 1741 -88 1753 88
rect 1787 -88 1799 88
rect 1741 -100 1799 -88
rect 1859 88 1917 100
rect 1859 -88 1871 88
rect 1905 -88 1917 88
rect 1859 -100 1917 -88
rect 1977 88 2035 100
rect 1977 -88 1989 88
rect 2023 -88 2035 88
rect 1977 -100 2035 -88
rect 2095 88 2153 100
rect 2095 -88 2107 88
rect 2141 -88 2153 88
rect 2095 -100 2153 -88
rect 2213 88 2271 100
rect 2213 -88 2225 88
rect 2259 -88 2271 88
rect 2213 -100 2271 -88
rect 2331 88 2389 100
rect 2331 -88 2343 88
rect 2377 -88 2389 88
rect 2331 -100 2389 -88
rect 2449 88 2507 100
rect 2449 -88 2461 88
rect 2495 -88 2507 88
rect 2449 -100 2507 -88
rect 2567 88 2625 100
rect 2567 -88 2579 88
rect 2613 -88 2625 88
rect 2567 -100 2625 -88
rect 2685 88 2743 100
rect 2685 -88 2697 88
rect 2731 -88 2743 88
rect 2685 -100 2743 -88
rect 2803 88 2861 100
rect 2803 -88 2815 88
rect 2849 -88 2861 88
rect 2803 -100 2861 -88
rect 2921 88 2979 100
rect 2921 -88 2933 88
rect 2967 -88 2979 88
rect 2921 -100 2979 -88
rect 3039 88 3097 100
rect 3039 -88 3051 88
rect 3085 -88 3097 88
rect 3039 -100 3097 -88
rect 3157 88 3215 100
rect 3157 -88 3169 88
rect 3203 -88 3215 88
rect 3157 -100 3215 -88
rect 3275 88 3333 100
rect 3275 -88 3287 88
rect 3321 -88 3333 88
rect 3275 -100 3333 -88
rect 3393 88 3451 100
rect 3393 -88 3405 88
rect 3439 -88 3451 88
rect 3393 -100 3451 -88
rect 3511 88 3569 100
rect 3511 -88 3523 88
rect 3557 -88 3569 88
rect 3511 -100 3569 -88
rect 3629 88 3687 100
rect 3629 -88 3641 88
rect 3675 -88 3687 88
rect 3629 -100 3687 -88
rect 3747 88 3805 100
rect 3747 -88 3759 88
rect 3793 -88 3805 88
rect 3747 -100 3805 -88
rect 3865 88 3923 100
rect 3865 -88 3877 88
rect 3911 -88 3923 88
rect 3865 -100 3923 -88
<< pdiffc >>
rect -3911 -88 -3877 88
rect -3793 -88 -3759 88
rect -3675 -88 -3641 88
rect -3557 -88 -3523 88
rect -3439 -88 -3405 88
rect -3321 -88 -3287 88
rect -3203 -88 -3169 88
rect -3085 -88 -3051 88
rect -2967 -88 -2933 88
rect -2849 -88 -2815 88
rect -2731 -88 -2697 88
rect -2613 -88 -2579 88
rect -2495 -88 -2461 88
rect -2377 -88 -2343 88
rect -2259 -88 -2225 88
rect -2141 -88 -2107 88
rect -2023 -88 -1989 88
rect -1905 -88 -1871 88
rect -1787 -88 -1753 88
rect -1669 -88 -1635 88
rect -1551 -88 -1517 88
rect -1433 -88 -1399 88
rect -1315 -88 -1281 88
rect -1197 -88 -1163 88
rect -1079 -88 -1045 88
rect -961 -88 -927 88
rect -843 -88 -809 88
rect -725 -88 -691 88
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
rect 691 -88 725 88
rect 809 -88 843 88
rect 927 -88 961 88
rect 1045 -88 1079 88
rect 1163 -88 1197 88
rect 1281 -88 1315 88
rect 1399 -88 1433 88
rect 1517 -88 1551 88
rect 1635 -88 1669 88
rect 1753 -88 1787 88
rect 1871 -88 1905 88
rect 1989 -88 2023 88
rect 2107 -88 2141 88
rect 2225 -88 2259 88
rect 2343 -88 2377 88
rect 2461 -88 2495 88
rect 2579 -88 2613 88
rect 2697 -88 2731 88
rect 2815 -88 2849 88
rect 2933 -88 2967 88
rect 3051 -88 3085 88
rect 3169 -88 3203 88
rect 3287 -88 3321 88
rect 3405 -88 3439 88
rect 3523 -88 3557 88
rect 3641 -88 3675 88
rect 3759 -88 3793 88
rect 3877 -88 3911 88
<< nsubdiff >>
rect -4025 249 -3929 283
rect 3929 249 4025 283
rect -4025 187 -3991 249
rect 3991 187 4025 249
rect -4025 -249 -3991 -187
rect 3991 -249 4025 -187
rect -4025 -283 -3929 -249
rect 3929 -283 4025 -249
<< nsubdiffcont >>
rect -3929 249 3929 283
rect -4025 -187 -3991 187
rect 3991 -187 4025 187
rect -3929 -283 3929 -249
<< poly >>
rect -3868 181 -3802 197
rect -3868 147 -3852 181
rect -3818 147 -3802 181
rect -3868 131 -3802 147
rect -3750 181 -3684 197
rect -3750 147 -3734 181
rect -3700 147 -3684 181
rect -3750 131 -3684 147
rect -3632 181 -3566 197
rect -3632 147 -3616 181
rect -3582 147 -3566 181
rect -3632 131 -3566 147
rect -3514 181 -3448 197
rect -3514 147 -3498 181
rect -3464 147 -3448 181
rect -3514 131 -3448 147
rect -3396 181 -3330 197
rect -3396 147 -3380 181
rect -3346 147 -3330 181
rect -3396 131 -3330 147
rect -3278 181 -3212 197
rect -3278 147 -3262 181
rect -3228 147 -3212 181
rect -3278 131 -3212 147
rect -3160 181 -3094 197
rect -3160 147 -3144 181
rect -3110 147 -3094 181
rect -3160 131 -3094 147
rect -3042 181 -2976 197
rect -3042 147 -3026 181
rect -2992 147 -2976 181
rect -3042 131 -2976 147
rect -2924 181 -2858 197
rect -2924 147 -2908 181
rect -2874 147 -2858 181
rect -2924 131 -2858 147
rect -2806 181 -2740 197
rect -2806 147 -2790 181
rect -2756 147 -2740 181
rect -2806 131 -2740 147
rect -2688 181 -2622 197
rect -2688 147 -2672 181
rect -2638 147 -2622 181
rect -2688 131 -2622 147
rect -2570 181 -2504 197
rect -2570 147 -2554 181
rect -2520 147 -2504 181
rect -2570 131 -2504 147
rect -2452 181 -2386 197
rect -2452 147 -2436 181
rect -2402 147 -2386 181
rect -2452 131 -2386 147
rect -2334 181 -2268 197
rect -2334 147 -2318 181
rect -2284 147 -2268 181
rect -2334 131 -2268 147
rect -2216 181 -2150 197
rect -2216 147 -2200 181
rect -2166 147 -2150 181
rect -2216 131 -2150 147
rect -2098 181 -2032 197
rect -2098 147 -2082 181
rect -2048 147 -2032 181
rect -2098 131 -2032 147
rect -1980 181 -1914 197
rect -1980 147 -1964 181
rect -1930 147 -1914 181
rect -1980 131 -1914 147
rect -1862 181 -1796 197
rect -1862 147 -1846 181
rect -1812 147 -1796 181
rect -1862 131 -1796 147
rect -1744 181 -1678 197
rect -1744 147 -1728 181
rect -1694 147 -1678 181
rect -1744 131 -1678 147
rect -1626 181 -1560 197
rect -1626 147 -1610 181
rect -1576 147 -1560 181
rect -1626 131 -1560 147
rect -1508 181 -1442 197
rect -1508 147 -1492 181
rect -1458 147 -1442 181
rect -1508 131 -1442 147
rect -1390 181 -1324 197
rect -1390 147 -1374 181
rect -1340 147 -1324 181
rect -1390 131 -1324 147
rect -1272 181 -1206 197
rect -1272 147 -1256 181
rect -1222 147 -1206 181
rect -1272 131 -1206 147
rect -1154 181 -1088 197
rect -1154 147 -1138 181
rect -1104 147 -1088 181
rect -1154 131 -1088 147
rect -1036 181 -970 197
rect -1036 147 -1020 181
rect -986 147 -970 181
rect -1036 131 -970 147
rect -918 181 -852 197
rect -918 147 -902 181
rect -868 147 -852 181
rect -918 131 -852 147
rect -800 181 -734 197
rect -800 147 -784 181
rect -750 147 -734 181
rect -800 131 -734 147
rect -682 181 -616 197
rect -682 147 -666 181
rect -632 147 -616 181
rect -682 131 -616 147
rect -564 181 -498 197
rect -564 147 -548 181
rect -514 147 -498 181
rect -564 131 -498 147
rect -446 181 -380 197
rect -446 147 -430 181
rect -396 147 -380 181
rect -446 131 -380 147
rect -328 181 -262 197
rect -328 147 -312 181
rect -278 147 -262 181
rect -328 131 -262 147
rect -210 181 -144 197
rect -210 147 -194 181
rect -160 147 -144 181
rect -210 131 -144 147
rect -92 181 -26 197
rect -92 147 -76 181
rect -42 147 -26 181
rect -92 131 -26 147
rect 26 181 92 197
rect 26 147 42 181
rect 76 147 92 181
rect 26 131 92 147
rect 144 181 210 197
rect 144 147 160 181
rect 194 147 210 181
rect 144 131 210 147
rect 262 181 328 197
rect 262 147 278 181
rect 312 147 328 181
rect 262 131 328 147
rect 380 181 446 197
rect 380 147 396 181
rect 430 147 446 181
rect 380 131 446 147
rect 498 181 564 197
rect 498 147 514 181
rect 548 147 564 181
rect 498 131 564 147
rect 616 181 682 197
rect 616 147 632 181
rect 666 147 682 181
rect 616 131 682 147
rect 734 181 800 197
rect 734 147 750 181
rect 784 147 800 181
rect 734 131 800 147
rect 852 181 918 197
rect 852 147 868 181
rect 902 147 918 181
rect 852 131 918 147
rect 970 181 1036 197
rect 970 147 986 181
rect 1020 147 1036 181
rect 970 131 1036 147
rect 1088 181 1154 197
rect 1088 147 1104 181
rect 1138 147 1154 181
rect 1088 131 1154 147
rect 1206 181 1272 197
rect 1206 147 1222 181
rect 1256 147 1272 181
rect 1206 131 1272 147
rect 1324 181 1390 197
rect 1324 147 1340 181
rect 1374 147 1390 181
rect 1324 131 1390 147
rect 1442 181 1508 197
rect 1442 147 1458 181
rect 1492 147 1508 181
rect 1442 131 1508 147
rect 1560 181 1626 197
rect 1560 147 1576 181
rect 1610 147 1626 181
rect 1560 131 1626 147
rect 1678 181 1744 197
rect 1678 147 1694 181
rect 1728 147 1744 181
rect 1678 131 1744 147
rect 1796 181 1862 197
rect 1796 147 1812 181
rect 1846 147 1862 181
rect 1796 131 1862 147
rect 1914 181 1980 197
rect 1914 147 1930 181
rect 1964 147 1980 181
rect 1914 131 1980 147
rect 2032 181 2098 197
rect 2032 147 2048 181
rect 2082 147 2098 181
rect 2032 131 2098 147
rect 2150 181 2216 197
rect 2150 147 2166 181
rect 2200 147 2216 181
rect 2150 131 2216 147
rect 2268 181 2334 197
rect 2268 147 2284 181
rect 2318 147 2334 181
rect 2268 131 2334 147
rect 2386 181 2452 197
rect 2386 147 2402 181
rect 2436 147 2452 181
rect 2386 131 2452 147
rect 2504 181 2570 197
rect 2504 147 2520 181
rect 2554 147 2570 181
rect 2504 131 2570 147
rect 2622 181 2688 197
rect 2622 147 2638 181
rect 2672 147 2688 181
rect 2622 131 2688 147
rect 2740 181 2806 197
rect 2740 147 2756 181
rect 2790 147 2806 181
rect 2740 131 2806 147
rect 2858 181 2924 197
rect 2858 147 2874 181
rect 2908 147 2924 181
rect 2858 131 2924 147
rect 2976 181 3042 197
rect 2976 147 2992 181
rect 3026 147 3042 181
rect 2976 131 3042 147
rect 3094 181 3160 197
rect 3094 147 3110 181
rect 3144 147 3160 181
rect 3094 131 3160 147
rect 3212 181 3278 197
rect 3212 147 3228 181
rect 3262 147 3278 181
rect 3212 131 3278 147
rect 3330 181 3396 197
rect 3330 147 3346 181
rect 3380 147 3396 181
rect 3330 131 3396 147
rect 3448 181 3514 197
rect 3448 147 3464 181
rect 3498 147 3514 181
rect 3448 131 3514 147
rect 3566 181 3632 197
rect 3566 147 3582 181
rect 3616 147 3632 181
rect 3566 131 3632 147
rect 3684 181 3750 197
rect 3684 147 3700 181
rect 3734 147 3750 181
rect 3684 131 3750 147
rect 3802 181 3868 197
rect 3802 147 3818 181
rect 3852 147 3868 181
rect 3802 131 3868 147
rect -3865 100 -3805 131
rect -3747 100 -3687 131
rect -3629 100 -3569 131
rect -3511 100 -3451 131
rect -3393 100 -3333 131
rect -3275 100 -3215 131
rect -3157 100 -3097 131
rect -3039 100 -2979 131
rect -2921 100 -2861 131
rect -2803 100 -2743 131
rect -2685 100 -2625 131
rect -2567 100 -2507 131
rect -2449 100 -2389 131
rect -2331 100 -2271 131
rect -2213 100 -2153 131
rect -2095 100 -2035 131
rect -1977 100 -1917 131
rect -1859 100 -1799 131
rect -1741 100 -1681 131
rect -1623 100 -1563 131
rect -1505 100 -1445 131
rect -1387 100 -1327 131
rect -1269 100 -1209 131
rect -1151 100 -1091 131
rect -1033 100 -973 131
rect -915 100 -855 131
rect -797 100 -737 131
rect -679 100 -619 131
rect -561 100 -501 131
rect -443 100 -383 131
rect -325 100 -265 131
rect -207 100 -147 131
rect -89 100 -29 131
rect 29 100 89 131
rect 147 100 207 131
rect 265 100 325 131
rect 383 100 443 131
rect 501 100 561 131
rect 619 100 679 131
rect 737 100 797 131
rect 855 100 915 131
rect 973 100 1033 131
rect 1091 100 1151 131
rect 1209 100 1269 131
rect 1327 100 1387 131
rect 1445 100 1505 131
rect 1563 100 1623 131
rect 1681 100 1741 131
rect 1799 100 1859 131
rect 1917 100 1977 131
rect 2035 100 2095 131
rect 2153 100 2213 131
rect 2271 100 2331 131
rect 2389 100 2449 131
rect 2507 100 2567 131
rect 2625 100 2685 131
rect 2743 100 2803 131
rect 2861 100 2921 131
rect 2979 100 3039 131
rect 3097 100 3157 131
rect 3215 100 3275 131
rect 3333 100 3393 131
rect 3451 100 3511 131
rect 3569 100 3629 131
rect 3687 100 3747 131
rect 3805 100 3865 131
rect -3865 -131 -3805 -100
rect -3747 -131 -3687 -100
rect -3629 -131 -3569 -100
rect -3511 -131 -3451 -100
rect -3393 -131 -3333 -100
rect -3275 -131 -3215 -100
rect -3157 -131 -3097 -100
rect -3039 -131 -2979 -100
rect -2921 -131 -2861 -100
rect -2803 -131 -2743 -100
rect -2685 -131 -2625 -100
rect -2567 -131 -2507 -100
rect -2449 -131 -2389 -100
rect -2331 -131 -2271 -100
rect -2213 -131 -2153 -100
rect -2095 -131 -2035 -100
rect -1977 -131 -1917 -100
rect -1859 -131 -1799 -100
rect -1741 -131 -1681 -100
rect -1623 -131 -1563 -100
rect -1505 -131 -1445 -100
rect -1387 -131 -1327 -100
rect -1269 -131 -1209 -100
rect -1151 -131 -1091 -100
rect -1033 -131 -973 -100
rect -915 -131 -855 -100
rect -797 -131 -737 -100
rect -679 -131 -619 -100
rect -561 -131 -501 -100
rect -443 -131 -383 -100
rect -325 -131 -265 -100
rect -207 -131 -147 -100
rect -89 -131 -29 -100
rect 29 -131 89 -100
rect 147 -131 207 -100
rect 265 -131 325 -100
rect 383 -131 443 -100
rect 501 -131 561 -100
rect 619 -131 679 -100
rect 737 -131 797 -100
rect 855 -131 915 -100
rect 973 -131 1033 -100
rect 1091 -131 1151 -100
rect 1209 -131 1269 -100
rect 1327 -131 1387 -100
rect 1445 -131 1505 -100
rect 1563 -131 1623 -100
rect 1681 -131 1741 -100
rect 1799 -131 1859 -100
rect 1917 -131 1977 -100
rect 2035 -131 2095 -100
rect 2153 -131 2213 -100
rect 2271 -131 2331 -100
rect 2389 -131 2449 -100
rect 2507 -131 2567 -100
rect 2625 -131 2685 -100
rect 2743 -131 2803 -100
rect 2861 -131 2921 -100
rect 2979 -131 3039 -100
rect 3097 -131 3157 -100
rect 3215 -131 3275 -100
rect 3333 -131 3393 -100
rect 3451 -131 3511 -100
rect 3569 -131 3629 -100
rect 3687 -131 3747 -100
rect 3805 -131 3865 -100
rect -3868 -147 -3802 -131
rect -3868 -181 -3852 -147
rect -3818 -181 -3802 -147
rect -3868 -197 -3802 -181
rect -3750 -147 -3684 -131
rect -3750 -181 -3734 -147
rect -3700 -181 -3684 -147
rect -3750 -197 -3684 -181
rect -3632 -147 -3566 -131
rect -3632 -181 -3616 -147
rect -3582 -181 -3566 -147
rect -3632 -197 -3566 -181
rect -3514 -147 -3448 -131
rect -3514 -181 -3498 -147
rect -3464 -181 -3448 -147
rect -3514 -197 -3448 -181
rect -3396 -147 -3330 -131
rect -3396 -181 -3380 -147
rect -3346 -181 -3330 -147
rect -3396 -197 -3330 -181
rect -3278 -147 -3212 -131
rect -3278 -181 -3262 -147
rect -3228 -181 -3212 -147
rect -3278 -197 -3212 -181
rect -3160 -147 -3094 -131
rect -3160 -181 -3144 -147
rect -3110 -181 -3094 -147
rect -3160 -197 -3094 -181
rect -3042 -147 -2976 -131
rect -3042 -181 -3026 -147
rect -2992 -181 -2976 -147
rect -3042 -197 -2976 -181
rect -2924 -147 -2858 -131
rect -2924 -181 -2908 -147
rect -2874 -181 -2858 -147
rect -2924 -197 -2858 -181
rect -2806 -147 -2740 -131
rect -2806 -181 -2790 -147
rect -2756 -181 -2740 -147
rect -2806 -197 -2740 -181
rect -2688 -147 -2622 -131
rect -2688 -181 -2672 -147
rect -2638 -181 -2622 -147
rect -2688 -197 -2622 -181
rect -2570 -147 -2504 -131
rect -2570 -181 -2554 -147
rect -2520 -181 -2504 -147
rect -2570 -197 -2504 -181
rect -2452 -147 -2386 -131
rect -2452 -181 -2436 -147
rect -2402 -181 -2386 -147
rect -2452 -197 -2386 -181
rect -2334 -147 -2268 -131
rect -2334 -181 -2318 -147
rect -2284 -181 -2268 -147
rect -2334 -197 -2268 -181
rect -2216 -147 -2150 -131
rect -2216 -181 -2200 -147
rect -2166 -181 -2150 -147
rect -2216 -197 -2150 -181
rect -2098 -147 -2032 -131
rect -2098 -181 -2082 -147
rect -2048 -181 -2032 -147
rect -2098 -197 -2032 -181
rect -1980 -147 -1914 -131
rect -1980 -181 -1964 -147
rect -1930 -181 -1914 -147
rect -1980 -197 -1914 -181
rect -1862 -147 -1796 -131
rect -1862 -181 -1846 -147
rect -1812 -181 -1796 -147
rect -1862 -197 -1796 -181
rect -1744 -147 -1678 -131
rect -1744 -181 -1728 -147
rect -1694 -181 -1678 -147
rect -1744 -197 -1678 -181
rect -1626 -147 -1560 -131
rect -1626 -181 -1610 -147
rect -1576 -181 -1560 -147
rect -1626 -197 -1560 -181
rect -1508 -147 -1442 -131
rect -1508 -181 -1492 -147
rect -1458 -181 -1442 -147
rect -1508 -197 -1442 -181
rect -1390 -147 -1324 -131
rect -1390 -181 -1374 -147
rect -1340 -181 -1324 -147
rect -1390 -197 -1324 -181
rect -1272 -147 -1206 -131
rect -1272 -181 -1256 -147
rect -1222 -181 -1206 -147
rect -1272 -197 -1206 -181
rect -1154 -147 -1088 -131
rect -1154 -181 -1138 -147
rect -1104 -181 -1088 -147
rect -1154 -197 -1088 -181
rect -1036 -147 -970 -131
rect -1036 -181 -1020 -147
rect -986 -181 -970 -147
rect -1036 -197 -970 -181
rect -918 -147 -852 -131
rect -918 -181 -902 -147
rect -868 -181 -852 -147
rect -918 -197 -852 -181
rect -800 -147 -734 -131
rect -800 -181 -784 -147
rect -750 -181 -734 -147
rect -800 -197 -734 -181
rect -682 -147 -616 -131
rect -682 -181 -666 -147
rect -632 -181 -616 -147
rect -682 -197 -616 -181
rect -564 -147 -498 -131
rect -564 -181 -548 -147
rect -514 -181 -498 -147
rect -564 -197 -498 -181
rect -446 -147 -380 -131
rect -446 -181 -430 -147
rect -396 -181 -380 -147
rect -446 -197 -380 -181
rect -328 -147 -262 -131
rect -328 -181 -312 -147
rect -278 -181 -262 -147
rect -328 -197 -262 -181
rect -210 -147 -144 -131
rect -210 -181 -194 -147
rect -160 -181 -144 -147
rect -210 -197 -144 -181
rect -92 -147 -26 -131
rect -92 -181 -76 -147
rect -42 -181 -26 -147
rect -92 -197 -26 -181
rect 26 -147 92 -131
rect 26 -181 42 -147
rect 76 -181 92 -147
rect 26 -197 92 -181
rect 144 -147 210 -131
rect 144 -181 160 -147
rect 194 -181 210 -147
rect 144 -197 210 -181
rect 262 -147 328 -131
rect 262 -181 278 -147
rect 312 -181 328 -147
rect 262 -197 328 -181
rect 380 -147 446 -131
rect 380 -181 396 -147
rect 430 -181 446 -147
rect 380 -197 446 -181
rect 498 -147 564 -131
rect 498 -181 514 -147
rect 548 -181 564 -147
rect 498 -197 564 -181
rect 616 -147 682 -131
rect 616 -181 632 -147
rect 666 -181 682 -147
rect 616 -197 682 -181
rect 734 -147 800 -131
rect 734 -181 750 -147
rect 784 -181 800 -147
rect 734 -197 800 -181
rect 852 -147 918 -131
rect 852 -181 868 -147
rect 902 -181 918 -147
rect 852 -197 918 -181
rect 970 -147 1036 -131
rect 970 -181 986 -147
rect 1020 -181 1036 -147
rect 970 -197 1036 -181
rect 1088 -147 1154 -131
rect 1088 -181 1104 -147
rect 1138 -181 1154 -147
rect 1088 -197 1154 -181
rect 1206 -147 1272 -131
rect 1206 -181 1222 -147
rect 1256 -181 1272 -147
rect 1206 -197 1272 -181
rect 1324 -147 1390 -131
rect 1324 -181 1340 -147
rect 1374 -181 1390 -147
rect 1324 -197 1390 -181
rect 1442 -147 1508 -131
rect 1442 -181 1458 -147
rect 1492 -181 1508 -147
rect 1442 -197 1508 -181
rect 1560 -147 1626 -131
rect 1560 -181 1576 -147
rect 1610 -181 1626 -147
rect 1560 -197 1626 -181
rect 1678 -147 1744 -131
rect 1678 -181 1694 -147
rect 1728 -181 1744 -147
rect 1678 -197 1744 -181
rect 1796 -147 1862 -131
rect 1796 -181 1812 -147
rect 1846 -181 1862 -147
rect 1796 -197 1862 -181
rect 1914 -147 1980 -131
rect 1914 -181 1930 -147
rect 1964 -181 1980 -147
rect 1914 -197 1980 -181
rect 2032 -147 2098 -131
rect 2032 -181 2048 -147
rect 2082 -181 2098 -147
rect 2032 -197 2098 -181
rect 2150 -147 2216 -131
rect 2150 -181 2166 -147
rect 2200 -181 2216 -147
rect 2150 -197 2216 -181
rect 2268 -147 2334 -131
rect 2268 -181 2284 -147
rect 2318 -181 2334 -147
rect 2268 -197 2334 -181
rect 2386 -147 2452 -131
rect 2386 -181 2402 -147
rect 2436 -181 2452 -147
rect 2386 -197 2452 -181
rect 2504 -147 2570 -131
rect 2504 -181 2520 -147
rect 2554 -181 2570 -147
rect 2504 -197 2570 -181
rect 2622 -147 2688 -131
rect 2622 -181 2638 -147
rect 2672 -181 2688 -147
rect 2622 -197 2688 -181
rect 2740 -147 2806 -131
rect 2740 -181 2756 -147
rect 2790 -181 2806 -147
rect 2740 -197 2806 -181
rect 2858 -147 2924 -131
rect 2858 -181 2874 -147
rect 2908 -181 2924 -147
rect 2858 -197 2924 -181
rect 2976 -147 3042 -131
rect 2976 -181 2992 -147
rect 3026 -181 3042 -147
rect 2976 -197 3042 -181
rect 3094 -147 3160 -131
rect 3094 -181 3110 -147
rect 3144 -181 3160 -147
rect 3094 -197 3160 -181
rect 3212 -147 3278 -131
rect 3212 -181 3228 -147
rect 3262 -181 3278 -147
rect 3212 -197 3278 -181
rect 3330 -147 3396 -131
rect 3330 -181 3346 -147
rect 3380 -181 3396 -147
rect 3330 -197 3396 -181
rect 3448 -147 3514 -131
rect 3448 -181 3464 -147
rect 3498 -181 3514 -147
rect 3448 -197 3514 -181
rect 3566 -147 3632 -131
rect 3566 -181 3582 -147
rect 3616 -181 3632 -147
rect 3566 -197 3632 -181
rect 3684 -147 3750 -131
rect 3684 -181 3700 -147
rect 3734 -181 3750 -147
rect 3684 -197 3750 -181
rect 3802 -147 3868 -131
rect 3802 -181 3818 -147
rect 3852 -181 3868 -147
rect 3802 -197 3868 -181
<< polycont >>
rect -3852 147 -3818 181
rect -3734 147 -3700 181
rect -3616 147 -3582 181
rect -3498 147 -3464 181
rect -3380 147 -3346 181
rect -3262 147 -3228 181
rect -3144 147 -3110 181
rect -3026 147 -2992 181
rect -2908 147 -2874 181
rect -2790 147 -2756 181
rect -2672 147 -2638 181
rect -2554 147 -2520 181
rect -2436 147 -2402 181
rect -2318 147 -2284 181
rect -2200 147 -2166 181
rect -2082 147 -2048 181
rect -1964 147 -1930 181
rect -1846 147 -1812 181
rect -1728 147 -1694 181
rect -1610 147 -1576 181
rect -1492 147 -1458 181
rect -1374 147 -1340 181
rect -1256 147 -1222 181
rect -1138 147 -1104 181
rect -1020 147 -986 181
rect -902 147 -868 181
rect -784 147 -750 181
rect -666 147 -632 181
rect -548 147 -514 181
rect -430 147 -396 181
rect -312 147 -278 181
rect -194 147 -160 181
rect -76 147 -42 181
rect 42 147 76 181
rect 160 147 194 181
rect 278 147 312 181
rect 396 147 430 181
rect 514 147 548 181
rect 632 147 666 181
rect 750 147 784 181
rect 868 147 902 181
rect 986 147 1020 181
rect 1104 147 1138 181
rect 1222 147 1256 181
rect 1340 147 1374 181
rect 1458 147 1492 181
rect 1576 147 1610 181
rect 1694 147 1728 181
rect 1812 147 1846 181
rect 1930 147 1964 181
rect 2048 147 2082 181
rect 2166 147 2200 181
rect 2284 147 2318 181
rect 2402 147 2436 181
rect 2520 147 2554 181
rect 2638 147 2672 181
rect 2756 147 2790 181
rect 2874 147 2908 181
rect 2992 147 3026 181
rect 3110 147 3144 181
rect 3228 147 3262 181
rect 3346 147 3380 181
rect 3464 147 3498 181
rect 3582 147 3616 181
rect 3700 147 3734 181
rect 3818 147 3852 181
rect -3852 -181 -3818 -147
rect -3734 -181 -3700 -147
rect -3616 -181 -3582 -147
rect -3498 -181 -3464 -147
rect -3380 -181 -3346 -147
rect -3262 -181 -3228 -147
rect -3144 -181 -3110 -147
rect -3026 -181 -2992 -147
rect -2908 -181 -2874 -147
rect -2790 -181 -2756 -147
rect -2672 -181 -2638 -147
rect -2554 -181 -2520 -147
rect -2436 -181 -2402 -147
rect -2318 -181 -2284 -147
rect -2200 -181 -2166 -147
rect -2082 -181 -2048 -147
rect -1964 -181 -1930 -147
rect -1846 -181 -1812 -147
rect -1728 -181 -1694 -147
rect -1610 -181 -1576 -147
rect -1492 -181 -1458 -147
rect -1374 -181 -1340 -147
rect -1256 -181 -1222 -147
rect -1138 -181 -1104 -147
rect -1020 -181 -986 -147
rect -902 -181 -868 -147
rect -784 -181 -750 -147
rect -666 -181 -632 -147
rect -548 -181 -514 -147
rect -430 -181 -396 -147
rect -312 -181 -278 -147
rect -194 -181 -160 -147
rect -76 -181 -42 -147
rect 42 -181 76 -147
rect 160 -181 194 -147
rect 278 -181 312 -147
rect 396 -181 430 -147
rect 514 -181 548 -147
rect 632 -181 666 -147
rect 750 -181 784 -147
rect 868 -181 902 -147
rect 986 -181 1020 -147
rect 1104 -181 1138 -147
rect 1222 -181 1256 -147
rect 1340 -181 1374 -147
rect 1458 -181 1492 -147
rect 1576 -181 1610 -147
rect 1694 -181 1728 -147
rect 1812 -181 1846 -147
rect 1930 -181 1964 -147
rect 2048 -181 2082 -147
rect 2166 -181 2200 -147
rect 2284 -181 2318 -147
rect 2402 -181 2436 -147
rect 2520 -181 2554 -147
rect 2638 -181 2672 -147
rect 2756 -181 2790 -147
rect 2874 -181 2908 -147
rect 2992 -181 3026 -147
rect 3110 -181 3144 -147
rect 3228 -181 3262 -147
rect 3346 -181 3380 -147
rect 3464 -181 3498 -147
rect 3582 -181 3616 -147
rect 3700 -181 3734 -147
rect 3818 -181 3852 -147
<< locali >>
rect -4025 249 -3929 283
rect 3929 249 4025 283
rect -4025 187 -3991 249
rect 3991 187 4025 249
rect -3868 147 -3852 181
rect -3818 147 -3802 181
rect -3750 147 -3734 181
rect -3700 147 -3684 181
rect -3632 147 -3616 181
rect -3582 147 -3566 181
rect -3514 147 -3498 181
rect -3464 147 -3448 181
rect -3396 147 -3380 181
rect -3346 147 -3330 181
rect -3278 147 -3262 181
rect -3228 147 -3212 181
rect -3160 147 -3144 181
rect -3110 147 -3094 181
rect -3042 147 -3026 181
rect -2992 147 -2976 181
rect -2924 147 -2908 181
rect -2874 147 -2858 181
rect -2806 147 -2790 181
rect -2756 147 -2740 181
rect -2688 147 -2672 181
rect -2638 147 -2622 181
rect -2570 147 -2554 181
rect -2520 147 -2504 181
rect -2452 147 -2436 181
rect -2402 147 -2386 181
rect -2334 147 -2318 181
rect -2284 147 -2268 181
rect -2216 147 -2200 181
rect -2166 147 -2150 181
rect -2098 147 -2082 181
rect -2048 147 -2032 181
rect -1980 147 -1964 181
rect -1930 147 -1914 181
rect -1862 147 -1846 181
rect -1812 147 -1796 181
rect -1744 147 -1728 181
rect -1694 147 -1678 181
rect -1626 147 -1610 181
rect -1576 147 -1560 181
rect -1508 147 -1492 181
rect -1458 147 -1442 181
rect -1390 147 -1374 181
rect -1340 147 -1324 181
rect -1272 147 -1256 181
rect -1222 147 -1206 181
rect -1154 147 -1138 181
rect -1104 147 -1088 181
rect -1036 147 -1020 181
rect -986 147 -970 181
rect -918 147 -902 181
rect -868 147 -852 181
rect -800 147 -784 181
rect -750 147 -734 181
rect -682 147 -666 181
rect -632 147 -616 181
rect -564 147 -548 181
rect -514 147 -498 181
rect -446 147 -430 181
rect -396 147 -380 181
rect -328 147 -312 181
rect -278 147 -262 181
rect -210 147 -194 181
rect -160 147 -144 181
rect -92 147 -76 181
rect -42 147 -26 181
rect 26 147 42 181
rect 76 147 92 181
rect 144 147 160 181
rect 194 147 210 181
rect 262 147 278 181
rect 312 147 328 181
rect 380 147 396 181
rect 430 147 446 181
rect 498 147 514 181
rect 548 147 564 181
rect 616 147 632 181
rect 666 147 682 181
rect 734 147 750 181
rect 784 147 800 181
rect 852 147 868 181
rect 902 147 918 181
rect 970 147 986 181
rect 1020 147 1036 181
rect 1088 147 1104 181
rect 1138 147 1154 181
rect 1206 147 1222 181
rect 1256 147 1272 181
rect 1324 147 1340 181
rect 1374 147 1390 181
rect 1442 147 1458 181
rect 1492 147 1508 181
rect 1560 147 1576 181
rect 1610 147 1626 181
rect 1678 147 1694 181
rect 1728 147 1744 181
rect 1796 147 1812 181
rect 1846 147 1862 181
rect 1914 147 1930 181
rect 1964 147 1980 181
rect 2032 147 2048 181
rect 2082 147 2098 181
rect 2150 147 2166 181
rect 2200 147 2216 181
rect 2268 147 2284 181
rect 2318 147 2334 181
rect 2386 147 2402 181
rect 2436 147 2452 181
rect 2504 147 2520 181
rect 2554 147 2570 181
rect 2622 147 2638 181
rect 2672 147 2688 181
rect 2740 147 2756 181
rect 2790 147 2806 181
rect 2858 147 2874 181
rect 2908 147 2924 181
rect 2976 147 2992 181
rect 3026 147 3042 181
rect 3094 147 3110 181
rect 3144 147 3160 181
rect 3212 147 3228 181
rect 3262 147 3278 181
rect 3330 147 3346 181
rect 3380 147 3396 181
rect 3448 147 3464 181
rect 3498 147 3514 181
rect 3566 147 3582 181
rect 3616 147 3632 181
rect 3684 147 3700 181
rect 3734 147 3750 181
rect 3802 147 3818 181
rect 3852 147 3868 181
rect -3911 88 -3877 104
rect -3911 -104 -3877 -88
rect -3793 88 -3759 104
rect -3793 -104 -3759 -88
rect -3675 88 -3641 104
rect -3675 -104 -3641 -88
rect -3557 88 -3523 104
rect -3557 -104 -3523 -88
rect -3439 88 -3405 104
rect -3439 -104 -3405 -88
rect -3321 88 -3287 104
rect -3321 -104 -3287 -88
rect -3203 88 -3169 104
rect -3203 -104 -3169 -88
rect -3085 88 -3051 104
rect -3085 -104 -3051 -88
rect -2967 88 -2933 104
rect -2967 -104 -2933 -88
rect -2849 88 -2815 104
rect -2849 -104 -2815 -88
rect -2731 88 -2697 104
rect -2731 -104 -2697 -88
rect -2613 88 -2579 104
rect -2613 -104 -2579 -88
rect -2495 88 -2461 104
rect -2495 -104 -2461 -88
rect -2377 88 -2343 104
rect -2377 -104 -2343 -88
rect -2259 88 -2225 104
rect -2259 -104 -2225 -88
rect -2141 88 -2107 104
rect -2141 -104 -2107 -88
rect -2023 88 -1989 104
rect -2023 -104 -1989 -88
rect -1905 88 -1871 104
rect -1905 -104 -1871 -88
rect -1787 88 -1753 104
rect -1787 -104 -1753 -88
rect -1669 88 -1635 104
rect -1669 -104 -1635 -88
rect -1551 88 -1517 104
rect -1551 -104 -1517 -88
rect -1433 88 -1399 104
rect -1433 -104 -1399 -88
rect -1315 88 -1281 104
rect -1315 -104 -1281 -88
rect -1197 88 -1163 104
rect -1197 -104 -1163 -88
rect -1079 88 -1045 104
rect -1079 -104 -1045 -88
rect -961 88 -927 104
rect -961 -104 -927 -88
rect -843 88 -809 104
rect -843 -104 -809 -88
rect -725 88 -691 104
rect -725 -104 -691 -88
rect -607 88 -573 104
rect -607 -104 -573 -88
rect -489 88 -455 104
rect -489 -104 -455 -88
rect -371 88 -337 104
rect -371 -104 -337 -88
rect -253 88 -219 104
rect -253 -104 -219 -88
rect -135 88 -101 104
rect -135 -104 -101 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 101 88 135 104
rect 101 -104 135 -88
rect 219 88 253 104
rect 219 -104 253 -88
rect 337 88 371 104
rect 337 -104 371 -88
rect 455 88 489 104
rect 455 -104 489 -88
rect 573 88 607 104
rect 573 -104 607 -88
rect 691 88 725 104
rect 691 -104 725 -88
rect 809 88 843 104
rect 809 -104 843 -88
rect 927 88 961 104
rect 927 -104 961 -88
rect 1045 88 1079 104
rect 1045 -104 1079 -88
rect 1163 88 1197 104
rect 1163 -104 1197 -88
rect 1281 88 1315 104
rect 1281 -104 1315 -88
rect 1399 88 1433 104
rect 1399 -104 1433 -88
rect 1517 88 1551 104
rect 1517 -104 1551 -88
rect 1635 88 1669 104
rect 1635 -104 1669 -88
rect 1753 88 1787 104
rect 1753 -104 1787 -88
rect 1871 88 1905 104
rect 1871 -104 1905 -88
rect 1989 88 2023 104
rect 1989 -104 2023 -88
rect 2107 88 2141 104
rect 2107 -104 2141 -88
rect 2225 88 2259 104
rect 2225 -104 2259 -88
rect 2343 88 2377 104
rect 2343 -104 2377 -88
rect 2461 88 2495 104
rect 2461 -104 2495 -88
rect 2579 88 2613 104
rect 2579 -104 2613 -88
rect 2697 88 2731 104
rect 2697 -104 2731 -88
rect 2815 88 2849 104
rect 2815 -104 2849 -88
rect 2933 88 2967 104
rect 2933 -104 2967 -88
rect 3051 88 3085 104
rect 3051 -104 3085 -88
rect 3169 88 3203 104
rect 3169 -104 3203 -88
rect 3287 88 3321 104
rect 3287 -104 3321 -88
rect 3405 88 3439 104
rect 3405 -104 3439 -88
rect 3523 88 3557 104
rect 3523 -104 3557 -88
rect 3641 88 3675 104
rect 3641 -104 3675 -88
rect 3759 88 3793 104
rect 3759 -104 3793 -88
rect 3877 88 3911 104
rect 3877 -104 3911 -88
rect -3868 -181 -3852 -147
rect -3818 -181 -3802 -147
rect -3750 -181 -3734 -147
rect -3700 -181 -3684 -147
rect -3632 -181 -3616 -147
rect -3582 -181 -3566 -147
rect -3514 -181 -3498 -147
rect -3464 -181 -3448 -147
rect -3396 -181 -3380 -147
rect -3346 -181 -3330 -147
rect -3278 -181 -3262 -147
rect -3228 -181 -3212 -147
rect -3160 -181 -3144 -147
rect -3110 -181 -3094 -147
rect -3042 -181 -3026 -147
rect -2992 -181 -2976 -147
rect -2924 -181 -2908 -147
rect -2874 -181 -2858 -147
rect -2806 -181 -2790 -147
rect -2756 -181 -2740 -147
rect -2688 -181 -2672 -147
rect -2638 -181 -2622 -147
rect -2570 -181 -2554 -147
rect -2520 -181 -2504 -147
rect -2452 -181 -2436 -147
rect -2402 -181 -2386 -147
rect -2334 -181 -2318 -147
rect -2284 -181 -2268 -147
rect -2216 -181 -2200 -147
rect -2166 -181 -2150 -147
rect -2098 -181 -2082 -147
rect -2048 -181 -2032 -147
rect -1980 -181 -1964 -147
rect -1930 -181 -1914 -147
rect -1862 -181 -1846 -147
rect -1812 -181 -1796 -147
rect -1744 -181 -1728 -147
rect -1694 -181 -1678 -147
rect -1626 -181 -1610 -147
rect -1576 -181 -1560 -147
rect -1508 -181 -1492 -147
rect -1458 -181 -1442 -147
rect -1390 -181 -1374 -147
rect -1340 -181 -1324 -147
rect -1272 -181 -1256 -147
rect -1222 -181 -1206 -147
rect -1154 -181 -1138 -147
rect -1104 -181 -1088 -147
rect -1036 -181 -1020 -147
rect -986 -181 -970 -147
rect -918 -181 -902 -147
rect -868 -181 -852 -147
rect -800 -181 -784 -147
rect -750 -181 -734 -147
rect -682 -181 -666 -147
rect -632 -181 -616 -147
rect -564 -181 -548 -147
rect -514 -181 -498 -147
rect -446 -181 -430 -147
rect -396 -181 -380 -147
rect -328 -181 -312 -147
rect -278 -181 -262 -147
rect -210 -181 -194 -147
rect -160 -181 -144 -147
rect -92 -181 -76 -147
rect -42 -181 -26 -147
rect 26 -181 42 -147
rect 76 -181 92 -147
rect 144 -181 160 -147
rect 194 -181 210 -147
rect 262 -181 278 -147
rect 312 -181 328 -147
rect 380 -181 396 -147
rect 430 -181 446 -147
rect 498 -181 514 -147
rect 548 -181 564 -147
rect 616 -181 632 -147
rect 666 -181 682 -147
rect 734 -181 750 -147
rect 784 -181 800 -147
rect 852 -181 868 -147
rect 902 -181 918 -147
rect 970 -181 986 -147
rect 1020 -181 1036 -147
rect 1088 -181 1104 -147
rect 1138 -181 1154 -147
rect 1206 -181 1222 -147
rect 1256 -181 1272 -147
rect 1324 -181 1340 -147
rect 1374 -181 1390 -147
rect 1442 -181 1458 -147
rect 1492 -181 1508 -147
rect 1560 -181 1576 -147
rect 1610 -181 1626 -147
rect 1678 -181 1694 -147
rect 1728 -181 1744 -147
rect 1796 -181 1812 -147
rect 1846 -181 1862 -147
rect 1914 -181 1930 -147
rect 1964 -181 1980 -147
rect 2032 -181 2048 -147
rect 2082 -181 2098 -147
rect 2150 -181 2166 -147
rect 2200 -181 2216 -147
rect 2268 -181 2284 -147
rect 2318 -181 2334 -147
rect 2386 -181 2402 -147
rect 2436 -181 2452 -147
rect 2504 -181 2520 -147
rect 2554 -181 2570 -147
rect 2622 -181 2638 -147
rect 2672 -181 2688 -147
rect 2740 -181 2756 -147
rect 2790 -181 2806 -147
rect 2858 -181 2874 -147
rect 2908 -181 2924 -147
rect 2976 -181 2992 -147
rect 3026 -181 3042 -147
rect 3094 -181 3110 -147
rect 3144 -181 3160 -147
rect 3212 -181 3228 -147
rect 3262 -181 3278 -147
rect 3330 -181 3346 -147
rect 3380 -181 3396 -147
rect 3448 -181 3464 -147
rect 3498 -181 3514 -147
rect 3566 -181 3582 -147
rect 3616 -181 3632 -147
rect 3684 -181 3700 -147
rect 3734 -181 3750 -147
rect 3802 -181 3818 -147
rect 3852 -181 3868 -147
rect -4025 -249 -3991 -187
rect 3991 -249 4025 -187
rect -4025 -283 -3929 -249
rect 3929 -283 4025 -249
<< viali >>
rect -3852 147 -3818 181
rect -3734 147 -3700 181
rect -3616 147 -3582 181
rect -3498 147 -3464 181
rect -3380 147 -3346 181
rect -3262 147 -3228 181
rect -3144 147 -3110 181
rect -3026 147 -2992 181
rect -2908 147 -2874 181
rect -2790 147 -2756 181
rect -2672 147 -2638 181
rect -2554 147 -2520 181
rect -2436 147 -2402 181
rect -2318 147 -2284 181
rect -2200 147 -2166 181
rect -2082 147 -2048 181
rect -1964 147 -1930 181
rect -1846 147 -1812 181
rect -1728 147 -1694 181
rect -1610 147 -1576 181
rect -1492 147 -1458 181
rect -1374 147 -1340 181
rect -1256 147 -1222 181
rect -1138 147 -1104 181
rect -1020 147 -986 181
rect -902 147 -868 181
rect -784 147 -750 181
rect -666 147 -632 181
rect -548 147 -514 181
rect -430 147 -396 181
rect -312 147 -278 181
rect -194 147 -160 181
rect -76 147 -42 181
rect 42 147 76 181
rect 160 147 194 181
rect 278 147 312 181
rect 396 147 430 181
rect 514 147 548 181
rect 632 147 666 181
rect 750 147 784 181
rect 868 147 902 181
rect 986 147 1020 181
rect 1104 147 1138 181
rect 1222 147 1256 181
rect 1340 147 1374 181
rect 1458 147 1492 181
rect 1576 147 1610 181
rect 1694 147 1728 181
rect 1812 147 1846 181
rect 1930 147 1964 181
rect 2048 147 2082 181
rect 2166 147 2200 181
rect 2284 147 2318 181
rect 2402 147 2436 181
rect 2520 147 2554 181
rect 2638 147 2672 181
rect 2756 147 2790 181
rect 2874 147 2908 181
rect 2992 147 3026 181
rect 3110 147 3144 181
rect 3228 147 3262 181
rect 3346 147 3380 181
rect 3464 147 3498 181
rect 3582 147 3616 181
rect 3700 147 3734 181
rect 3818 147 3852 181
rect -3911 -88 -3877 88
rect -3793 -88 -3759 88
rect -3675 -88 -3641 88
rect -3557 -88 -3523 88
rect -3439 -88 -3405 88
rect -3321 -88 -3287 88
rect -3203 -88 -3169 88
rect -3085 -88 -3051 88
rect -2967 -88 -2933 88
rect -2849 -88 -2815 88
rect -2731 -88 -2697 88
rect -2613 -88 -2579 88
rect -2495 -88 -2461 88
rect -2377 -88 -2343 88
rect -2259 -88 -2225 88
rect -2141 -88 -2107 88
rect -2023 -88 -1989 88
rect -1905 -88 -1871 88
rect -1787 -88 -1753 88
rect -1669 -88 -1635 88
rect -1551 -88 -1517 88
rect -1433 -88 -1399 88
rect -1315 -88 -1281 88
rect -1197 -88 -1163 88
rect -1079 -88 -1045 88
rect -961 -88 -927 88
rect -843 -88 -809 88
rect -725 -88 -691 88
rect -607 -88 -573 88
rect -489 -88 -455 88
rect -371 -88 -337 88
rect -253 -88 -219 88
rect -135 -88 -101 88
rect -17 -88 17 88
rect 101 -88 135 88
rect 219 -88 253 88
rect 337 -88 371 88
rect 455 -88 489 88
rect 573 -88 607 88
rect 691 -88 725 88
rect 809 -88 843 88
rect 927 -88 961 88
rect 1045 -88 1079 88
rect 1163 -88 1197 88
rect 1281 -88 1315 88
rect 1399 -88 1433 88
rect 1517 -88 1551 88
rect 1635 -88 1669 88
rect 1753 -88 1787 88
rect 1871 -88 1905 88
rect 1989 -88 2023 88
rect 2107 -88 2141 88
rect 2225 -88 2259 88
rect 2343 -88 2377 88
rect 2461 -88 2495 88
rect 2579 -88 2613 88
rect 2697 -88 2731 88
rect 2815 -88 2849 88
rect 2933 -88 2967 88
rect 3051 -88 3085 88
rect 3169 -88 3203 88
rect 3287 -88 3321 88
rect 3405 -88 3439 88
rect 3523 -88 3557 88
rect 3641 -88 3675 88
rect 3759 -88 3793 88
rect 3877 -88 3911 88
rect -3852 -181 -3818 -147
rect -3734 -181 -3700 -147
rect -3616 -181 -3582 -147
rect -3498 -181 -3464 -147
rect -3380 -181 -3346 -147
rect -3262 -181 -3228 -147
rect -3144 -181 -3110 -147
rect -3026 -181 -2992 -147
rect -2908 -181 -2874 -147
rect -2790 -181 -2756 -147
rect -2672 -181 -2638 -147
rect -2554 -181 -2520 -147
rect -2436 -181 -2402 -147
rect -2318 -181 -2284 -147
rect -2200 -181 -2166 -147
rect -2082 -181 -2048 -147
rect -1964 -181 -1930 -147
rect -1846 -181 -1812 -147
rect -1728 -181 -1694 -147
rect -1610 -181 -1576 -147
rect -1492 -181 -1458 -147
rect -1374 -181 -1340 -147
rect -1256 -181 -1222 -147
rect -1138 -181 -1104 -147
rect -1020 -181 -986 -147
rect -902 -181 -868 -147
rect -784 -181 -750 -147
rect -666 -181 -632 -147
rect -548 -181 -514 -147
rect -430 -181 -396 -147
rect -312 -181 -278 -147
rect -194 -181 -160 -147
rect -76 -181 -42 -147
rect 42 -181 76 -147
rect 160 -181 194 -147
rect 278 -181 312 -147
rect 396 -181 430 -147
rect 514 -181 548 -147
rect 632 -181 666 -147
rect 750 -181 784 -147
rect 868 -181 902 -147
rect 986 -181 1020 -147
rect 1104 -181 1138 -147
rect 1222 -181 1256 -147
rect 1340 -181 1374 -147
rect 1458 -181 1492 -147
rect 1576 -181 1610 -147
rect 1694 -181 1728 -147
rect 1812 -181 1846 -147
rect 1930 -181 1964 -147
rect 2048 -181 2082 -147
rect 2166 -181 2200 -147
rect 2284 -181 2318 -147
rect 2402 -181 2436 -147
rect 2520 -181 2554 -147
rect 2638 -181 2672 -147
rect 2756 -181 2790 -147
rect 2874 -181 2908 -147
rect 2992 -181 3026 -147
rect 3110 -181 3144 -147
rect 3228 -181 3262 -147
rect 3346 -181 3380 -147
rect 3464 -181 3498 -147
rect 3582 -181 3616 -147
rect 3700 -181 3734 -147
rect 3818 -181 3852 -147
<< metal1 >>
rect -3864 181 -3806 187
rect -3864 147 -3852 181
rect -3818 147 -3806 181
rect -3864 141 -3806 147
rect -3746 181 -3688 187
rect -3746 147 -3734 181
rect -3700 147 -3688 181
rect -3746 141 -3688 147
rect -3628 181 -3570 187
rect -3628 147 -3616 181
rect -3582 147 -3570 181
rect -3628 141 -3570 147
rect -3510 181 -3452 187
rect -3510 147 -3498 181
rect -3464 147 -3452 181
rect -3510 141 -3452 147
rect -3392 181 -3334 187
rect -3392 147 -3380 181
rect -3346 147 -3334 181
rect -3392 141 -3334 147
rect -3274 181 -3216 187
rect -3274 147 -3262 181
rect -3228 147 -3216 181
rect -3274 141 -3216 147
rect -3156 181 -3098 187
rect -3156 147 -3144 181
rect -3110 147 -3098 181
rect -3156 141 -3098 147
rect -3038 181 -2980 187
rect -3038 147 -3026 181
rect -2992 147 -2980 181
rect -3038 141 -2980 147
rect -2920 181 -2862 187
rect -2920 147 -2908 181
rect -2874 147 -2862 181
rect -2920 141 -2862 147
rect -2802 181 -2744 187
rect -2802 147 -2790 181
rect -2756 147 -2744 181
rect -2802 141 -2744 147
rect -2684 181 -2626 187
rect -2684 147 -2672 181
rect -2638 147 -2626 181
rect -2684 141 -2626 147
rect -2566 181 -2508 187
rect -2566 147 -2554 181
rect -2520 147 -2508 181
rect -2566 141 -2508 147
rect -2448 181 -2390 187
rect -2448 147 -2436 181
rect -2402 147 -2390 181
rect -2448 141 -2390 147
rect -2330 181 -2272 187
rect -2330 147 -2318 181
rect -2284 147 -2272 181
rect -2330 141 -2272 147
rect -2212 181 -2154 187
rect -2212 147 -2200 181
rect -2166 147 -2154 181
rect -2212 141 -2154 147
rect -2094 181 -2036 187
rect -2094 147 -2082 181
rect -2048 147 -2036 181
rect -2094 141 -2036 147
rect -1976 181 -1918 187
rect -1976 147 -1964 181
rect -1930 147 -1918 181
rect -1976 141 -1918 147
rect -1858 181 -1800 187
rect -1858 147 -1846 181
rect -1812 147 -1800 181
rect -1858 141 -1800 147
rect -1740 181 -1682 187
rect -1740 147 -1728 181
rect -1694 147 -1682 181
rect -1740 141 -1682 147
rect -1622 181 -1564 187
rect -1622 147 -1610 181
rect -1576 147 -1564 181
rect -1622 141 -1564 147
rect -1504 181 -1446 187
rect -1504 147 -1492 181
rect -1458 147 -1446 181
rect -1504 141 -1446 147
rect -1386 181 -1328 187
rect -1386 147 -1374 181
rect -1340 147 -1328 181
rect -1386 141 -1328 147
rect -1268 181 -1210 187
rect -1268 147 -1256 181
rect -1222 147 -1210 181
rect -1268 141 -1210 147
rect -1150 181 -1092 187
rect -1150 147 -1138 181
rect -1104 147 -1092 181
rect -1150 141 -1092 147
rect -1032 181 -974 187
rect -1032 147 -1020 181
rect -986 147 -974 181
rect -1032 141 -974 147
rect -914 181 -856 187
rect -914 147 -902 181
rect -868 147 -856 181
rect -914 141 -856 147
rect -796 181 -738 187
rect -796 147 -784 181
rect -750 147 -738 181
rect -796 141 -738 147
rect -678 181 -620 187
rect -678 147 -666 181
rect -632 147 -620 181
rect -678 141 -620 147
rect -560 181 -502 187
rect -560 147 -548 181
rect -514 147 -502 181
rect -560 141 -502 147
rect -442 181 -384 187
rect -442 147 -430 181
rect -396 147 -384 181
rect -442 141 -384 147
rect -324 181 -266 187
rect -324 147 -312 181
rect -278 147 -266 181
rect -324 141 -266 147
rect -206 181 -148 187
rect -206 147 -194 181
rect -160 147 -148 181
rect -206 141 -148 147
rect -88 181 -30 187
rect -88 147 -76 181
rect -42 147 -30 181
rect -88 141 -30 147
rect 30 181 88 187
rect 30 147 42 181
rect 76 147 88 181
rect 30 141 88 147
rect 148 181 206 187
rect 148 147 160 181
rect 194 147 206 181
rect 148 141 206 147
rect 266 181 324 187
rect 266 147 278 181
rect 312 147 324 181
rect 266 141 324 147
rect 384 181 442 187
rect 384 147 396 181
rect 430 147 442 181
rect 384 141 442 147
rect 502 181 560 187
rect 502 147 514 181
rect 548 147 560 181
rect 502 141 560 147
rect 620 181 678 187
rect 620 147 632 181
rect 666 147 678 181
rect 620 141 678 147
rect 738 181 796 187
rect 738 147 750 181
rect 784 147 796 181
rect 738 141 796 147
rect 856 181 914 187
rect 856 147 868 181
rect 902 147 914 181
rect 856 141 914 147
rect 974 181 1032 187
rect 974 147 986 181
rect 1020 147 1032 181
rect 974 141 1032 147
rect 1092 181 1150 187
rect 1092 147 1104 181
rect 1138 147 1150 181
rect 1092 141 1150 147
rect 1210 181 1268 187
rect 1210 147 1222 181
rect 1256 147 1268 181
rect 1210 141 1268 147
rect 1328 181 1386 187
rect 1328 147 1340 181
rect 1374 147 1386 181
rect 1328 141 1386 147
rect 1446 181 1504 187
rect 1446 147 1458 181
rect 1492 147 1504 181
rect 1446 141 1504 147
rect 1564 181 1622 187
rect 1564 147 1576 181
rect 1610 147 1622 181
rect 1564 141 1622 147
rect 1682 181 1740 187
rect 1682 147 1694 181
rect 1728 147 1740 181
rect 1682 141 1740 147
rect 1800 181 1858 187
rect 1800 147 1812 181
rect 1846 147 1858 181
rect 1800 141 1858 147
rect 1918 181 1976 187
rect 1918 147 1930 181
rect 1964 147 1976 181
rect 1918 141 1976 147
rect 2036 181 2094 187
rect 2036 147 2048 181
rect 2082 147 2094 181
rect 2036 141 2094 147
rect 2154 181 2212 187
rect 2154 147 2166 181
rect 2200 147 2212 181
rect 2154 141 2212 147
rect 2272 181 2330 187
rect 2272 147 2284 181
rect 2318 147 2330 181
rect 2272 141 2330 147
rect 2390 181 2448 187
rect 2390 147 2402 181
rect 2436 147 2448 181
rect 2390 141 2448 147
rect 2508 181 2566 187
rect 2508 147 2520 181
rect 2554 147 2566 181
rect 2508 141 2566 147
rect 2626 181 2684 187
rect 2626 147 2638 181
rect 2672 147 2684 181
rect 2626 141 2684 147
rect 2744 181 2802 187
rect 2744 147 2756 181
rect 2790 147 2802 181
rect 2744 141 2802 147
rect 2862 181 2920 187
rect 2862 147 2874 181
rect 2908 147 2920 181
rect 2862 141 2920 147
rect 2980 181 3038 187
rect 2980 147 2992 181
rect 3026 147 3038 181
rect 2980 141 3038 147
rect 3098 181 3156 187
rect 3098 147 3110 181
rect 3144 147 3156 181
rect 3098 141 3156 147
rect 3216 181 3274 187
rect 3216 147 3228 181
rect 3262 147 3274 181
rect 3216 141 3274 147
rect 3334 181 3392 187
rect 3334 147 3346 181
rect 3380 147 3392 181
rect 3334 141 3392 147
rect 3452 181 3510 187
rect 3452 147 3464 181
rect 3498 147 3510 181
rect 3452 141 3510 147
rect 3570 181 3628 187
rect 3570 147 3582 181
rect 3616 147 3628 181
rect 3570 141 3628 147
rect 3688 181 3746 187
rect 3688 147 3700 181
rect 3734 147 3746 181
rect 3688 141 3746 147
rect 3806 181 3864 187
rect 3806 147 3818 181
rect 3852 147 3864 181
rect 3806 141 3864 147
rect -3917 88 -3871 100
rect -3917 -88 -3911 88
rect -3877 -88 -3871 88
rect -3917 -100 -3871 -88
rect -3799 88 -3753 100
rect -3799 -88 -3793 88
rect -3759 -88 -3753 88
rect -3799 -100 -3753 -88
rect -3681 88 -3635 100
rect -3681 -88 -3675 88
rect -3641 -88 -3635 88
rect -3681 -100 -3635 -88
rect -3563 88 -3517 100
rect -3563 -88 -3557 88
rect -3523 -88 -3517 88
rect -3563 -100 -3517 -88
rect -3445 88 -3399 100
rect -3445 -88 -3439 88
rect -3405 -88 -3399 88
rect -3445 -100 -3399 -88
rect -3327 88 -3281 100
rect -3327 -88 -3321 88
rect -3287 -88 -3281 88
rect -3327 -100 -3281 -88
rect -3209 88 -3163 100
rect -3209 -88 -3203 88
rect -3169 -88 -3163 88
rect -3209 -100 -3163 -88
rect -3091 88 -3045 100
rect -3091 -88 -3085 88
rect -3051 -88 -3045 88
rect -3091 -100 -3045 -88
rect -2973 88 -2927 100
rect -2973 -88 -2967 88
rect -2933 -88 -2927 88
rect -2973 -100 -2927 -88
rect -2855 88 -2809 100
rect -2855 -88 -2849 88
rect -2815 -88 -2809 88
rect -2855 -100 -2809 -88
rect -2737 88 -2691 100
rect -2737 -88 -2731 88
rect -2697 -88 -2691 88
rect -2737 -100 -2691 -88
rect -2619 88 -2573 100
rect -2619 -88 -2613 88
rect -2579 -88 -2573 88
rect -2619 -100 -2573 -88
rect -2501 88 -2455 100
rect -2501 -88 -2495 88
rect -2461 -88 -2455 88
rect -2501 -100 -2455 -88
rect -2383 88 -2337 100
rect -2383 -88 -2377 88
rect -2343 -88 -2337 88
rect -2383 -100 -2337 -88
rect -2265 88 -2219 100
rect -2265 -88 -2259 88
rect -2225 -88 -2219 88
rect -2265 -100 -2219 -88
rect -2147 88 -2101 100
rect -2147 -88 -2141 88
rect -2107 -88 -2101 88
rect -2147 -100 -2101 -88
rect -2029 88 -1983 100
rect -2029 -88 -2023 88
rect -1989 -88 -1983 88
rect -2029 -100 -1983 -88
rect -1911 88 -1865 100
rect -1911 -88 -1905 88
rect -1871 -88 -1865 88
rect -1911 -100 -1865 -88
rect -1793 88 -1747 100
rect -1793 -88 -1787 88
rect -1753 -88 -1747 88
rect -1793 -100 -1747 -88
rect -1675 88 -1629 100
rect -1675 -88 -1669 88
rect -1635 -88 -1629 88
rect -1675 -100 -1629 -88
rect -1557 88 -1511 100
rect -1557 -88 -1551 88
rect -1517 -88 -1511 88
rect -1557 -100 -1511 -88
rect -1439 88 -1393 100
rect -1439 -88 -1433 88
rect -1399 -88 -1393 88
rect -1439 -100 -1393 -88
rect -1321 88 -1275 100
rect -1321 -88 -1315 88
rect -1281 -88 -1275 88
rect -1321 -100 -1275 -88
rect -1203 88 -1157 100
rect -1203 -88 -1197 88
rect -1163 -88 -1157 88
rect -1203 -100 -1157 -88
rect -1085 88 -1039 100
rect -1085 -88 -1079 88
rect -1045 -88 -1039 88
rect -1085 -100 -1039 -88
rect -967 88 -921 100
rect -967 -88 -961 88
rect -927 -88 -921 88
rect -967 -100 -921 -88
rect -849 88 -803 100
rect -849 -88 -843 88
rect -809 -88 -803 88
rect -849 -100 -803 -88
rect -731 88 -685 100
rect -731 -88 -725 88
rect -691 -88 -685 88
rect -731 -100 -685 -88
rect -613 88 -567 100
rect -613 -88 -607 88
rect -573 -88 -567 88
rect -613 -100 -567 -88
rect -495 88 -449 100
rect -495 -88 -489 88
rect -455 -88 -449 88
rect -495 -100 -449 -88
rect -377 88 -331 100
rect -377 -88 -371 88
rect -337 -88 -331 88
rect -377 -100 -331 -88
rect -259 88 -213 100
rect -259 -88 -253 88
rect -219 -88 -213 88
rect -259 -100 -213 -88
rect -141 88 -95 100
rect -141 -88 -135 88
rect -101 -88 -95 88
rect -141 -100 -95 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 95 88 141 100
rect 95 -88 101 88
rect 135 -88 141 88
rect 95 -100 141 -88
rect 213 88 259 100
rect 213 -88 219 88
rect 253 -88 259 88
rect 213 -100 259 -88
rect 331 88 377 100
rect 331 -88 337 88
rect 371 -88 377 88
rect 331 -100 377 -88
rect 449 88 495 100
rect 449 -88 455 88
rect 489 -88 495 88
rect 449 -100 495 -88
rect 567 88 613 100
rect 567 -88 573 88
rect 607 -88 613 88
rect 567 -100 613 -88
rect 685 88 731 100
rect 685 -88 691 88
rect 725 -88 731 88
rect 685 -100 731 -88
rect 803 88 849 100
rect 803 -88 809 88
rect 843 -88 849 88
rect 803 -100 849 -88
rect 921 88 967 100
rect 921 -88 927 88
rect 961 -88 967 88
rect 921 -100 967 -88
rect 1039 88 1085 100
rect 1039 -88 1045 88
rect 1079 -88 1085 88
rect 1039 -100 1085 -88
rect 1157 88 1203 100
rect 1157 -88 1163 88
rect 1197 -88 1203 88
rect 1157 -100 1203 -88
rect 1275 88 1321 100
rect 1275 -88 1281 88
rect 1315 -88 1321 88
rect 1275 -100 1321 -88
rect 1393 88 1439 100
rect 1393 -88 1399 88
rect 1433 -88 1439 88
rect 1393 -100 1439 -88
rect 1511 88 1557 100
rect 1511 -88 1517 88
rect 1551 -88 1557 88
rect 1511 -100 1557 -88
rect 1629 88 1675 100
rect 1629 -88 1635 88
rect 1669 -88 1675 88
rect 1629 -100 1675 -88
rect 1747 88 1793 100
rect 1747 -88 1753 88
rect 1787 -88 1793 88
rect 1747 -100 1793 -88
rect 1865 88 1911 100
rect 1865 -88 1871 88
rect 1905 -88 1911 88
rect 1865 -100 1911 -88
rect 1983 88 2029 100
rect 1983 -88 1989 88
rect 2023 -88 2029 88
rect 1983 -100 2029 -88
rect 2101 88 2147 100
rect 2101 -88 2107 88
rect 2141 -88 2147 88
rect 2101 -100 2147 -88
rect 2219 88 2265 100
rect 2219 -88 2225 88
rect 2259 -88 2265 88
rect 2219 -100 2265 -88
rect 2337 88 2383 100
rect 2337 -88 2343 88
rect 2377 -88 2383 88
rect 2337 -100 2383 -88
rect 2455 88 2501 100
rect 2455 -88 2461 88
rect 2495 -88 2501 88
rect 2455 -100 2501 -88
rect 2573 88 2619 100
rect 2573 -88 2579 88
rect 2613 -88 2619 88
rect 2573 -100 2619 -88
rect 2691 88 2737 100
rect 2691 -88 2697 88
rect 2731 -88 2737 88
rect 2691 -100 2737 -88
rect 2809 88 2855 100
rect 2809 -88 2815 88
rect 2849 -88 2855 88
rect 2809 -100 2855 -88
rect 2927 88 2973 100
rect 2927 -88 2933 88
rect 2967 -88 2973 88
rect 2927 -100 2973 -88
rect 3045 88 3091 100
rect 3045 -88 3051 88
rect 3085 -88 3091 88
rect 3045 -100 3091 -88
rect 3163 88 3209 100
rect 3163 -88 3169 88
rect 3203 -88 3209 88
rect 3163 -100 3209 -88
rect 3281 88 3327 100
rect 3281 -88 3287 88
rect 3321 -88 3327 88
rect 3281 -100 3327 -88
rect 3399 88 3445 100
rect 3399 -88 3405 88
rect 3439 -88 3445 88
rect 3399 -100 3445 -88
rect 3517 88 3563 100
rect 3517 -88 3523 88
rect 3557 -88 3563 88
rect 3517 -100 3563 -88
rect 3635 88 3681 100
rect 3635 -88 3641 88
rect 3675 -88 3681 88
rect 3635 -100 3681 -88
rect 3753 88 3799 100
rect 3753 -88 3759 88
rect 3793 -88 3799 88
rect 3753 -100 3799 -88
rect 3871 88 3917 100
rect 3871 -88 3877 88
rect 3911 -88 3917 88
rect 3871 -100 3917 -88
rect -3864 -147 -3806 -141
rect -3864 -181 -3852 -147
rect -3818 -181 -3806 -147
rect -3864 -187 -3806 -181
rect -3746 -147 -3688 -141
rect -3746 -181 -3734 -147
rect -3700 -181 -3688 -147
rect -3746 -187 -3688 -181
rect -3628 -147 -3570 -141
rect -3628 -181 -3616 -147
rect -3582 -181 -3570 -147
rect -3628 -187 -3570 -181
rect -3510 -147 -3452 -141
rect -3510 -181 -3498 -147
rect -3464 -181 -3452 -147
rect -3510 -187 -3452 -181
rect -3392 -147 -3334 -141
rect -3392 -181 -3380 -147
rect -3346 -181 -3334 -147
rect -3392 -187 -3334 -181
rect -3274 -147 -3216 -141
rect -3274 -181 -3262 -147
rect -3228 -181 -3216 -147
rect -3274 -187 -3216 -181
rect -3156 -147 -3098 -141
rect -3156 -181 -3144 -147
rect -3110 -181 -3098 -147
rect -3156 -187 -3098 -181
rect -3038 -147 -2980 -141
rect -3038 -181 -3026 -147
rect -2992 -181 -2980 -147
rect -3038 -187 -2980 -181
rect -2920 -147 -2862 -141
rect -2920 -181 -2908 -147
rect -2874 -181 -2862 -147
rect -2920 -187 -2862 -181
rect -2802 -147 -2744 -141
rect -2802 -181 -2790 -147
rect -2756 -181 -2744 -147
rect -2802 -187 -2744 -181
rect -2684 -147 -2626 -141
rect -2684 -181 -2672 -147
rect -2638 -181 -2626 -147
rect -2684 -187 -2626 -181
rect -2566 -147 -2508 -141
rect -2566 -181 -2554 -147
rect -2520 -181 -2508 -147
rect -2566 -187 -2508 -181
rect -2448 -147 -2390 -141
rect -2448 -181 -2436 -147
rect -2402 -181 -2390 -147
rect -2448 -187 -2390 -181
rect -2330 -147 -2272 -141
rect -2330 -181 -2318 -147
rect -2284 -181 -2272 -147
rect -2330 -187 -2272 -181
rect -2212 -147 -2154 -141
rect -2212 -181 -2200 -147
rect -2166 -181 -2154 -147
rect -2212 -187 -2154 -181
rect -2094 -147 -2036 -141
rect -2094 -181 -2082 -147
rect -2048 -181 -2036 -147
rect -2094 -187 -2036 -181
rect -1976 -147 -1918 -141
rect -1976 -181 -1964 -147
rect -1930 -181 -1918 -147
rect -1976 -187 -1918 -181
rect -1858 -147 -1800 -141
rect -1858 -181 -1846 -147
rect -1812 -181 -1800 -147
rect -1858 -187 -1800 -181
rect -1740 -147 -1682 -141
rect -1740 -181 -1728 -147
rect -1694 -181 -1682 -147
rect -1740 -187 -1682 -181
rect -1622 -147 -1564 -141
rect -1622 -181 -1610 -147
rect -1576 -181 -1564 -147
rect -1622 -187 -1564 -181
rect -1504 -147 -1446 -141
rect -1504 -181 -1492 -147
rect -1458 -181 -1446 -147
rect -1504 -187 -1446 -181
rect -1386 -147 -1328 -141
rect -1386 -181 -1374 -147
rect -1340 -181 -1328 -147
rect -1386 -187 -1328 -181
rect -1268 -147 -1210 -141
rect -1268 -181 -1256 -147
rect -1222 -181 -1210 -147
rect -1268 -187 -1210 -181
rect -1150 -147 -1092 -141
rect -1150 -181 -1138 -147
rect -1104 -181 -1092 -147
rect -1150 -187 -1092 -181
rect -1032 -147 -974 -141
rect -1032 -181 -1020 -147
rect -986 -181 -974 -147
rect -1032 -187 -974 -181
rect -914 -147 -856 -141
rect -914 -181 -902 -147
rect -868 -181 -856 -147
rect -914 -187 -856 -181
rect -796 -147 -738 -141
rect -796 -181 -784 -147
rect -750 -181 -738 -147
rect -796 -187 -738 -181
rect -678 -147 -620 -141
rect -678 -181 -666 -147
rect -632 -181 -620 -147
rect -678 -187 -620 -181
rect -560 -147 -502 -141
rect -560 -181 -548 -147
rect -514 -181 -502 -147
rect -560 -187 -502 -181
rect -442 -147 -384 -141
rect -442 -181 -430 -147
rect -396 -181 -384 -147
rect -442 -187 -384 -181
rect -324 -147 -266 -141
rect -324 -181 -312 -147
rect -278 -181 -266 -147
rect -324 -187 -266 -181
rect -206 -147 -148 -141
rect -206 -181 -194 -147
rect -160 -181 -148 -147
rect -206 -187 -148 -181
rect -88 -147 -30 -141
rect -88 -181 -76 -147
rect -42 -181 -30 -147
rect -88 -187 -30 -181
rect 30 -147 88 -141
rect 30 -181 42 -147
rect 76 -181 88 -147
rect 30 -187 88 -181
rect 148 -147 206 -141
rect 148 -181 160 -147
rect 194 -181 206 -147
rect 148 -187 206 -181
rect 266 -147 324 -141
rect 266 -181 278 -147
rect 312 -181 324 -147
rect 266 -187 324 -181
rect 384 -147 442 -141
rect 384 -181 396 -147
rect 430 -181 442 -147
rect 384 -187 442 -181
rect 502 -147 560 -141
rect 502 -181 514 -147
rect 548 -181 560 -147
rect 502 -187 560 -181
rect 620 -147 678 -141
rect 620 -181 632 -147
rect 666 -181 678 -147
rect 620 -187 678 -181
rect 738 -147 796 -141
rect 738 -181 750 -147
rect 784 -181 796 -147
rect 738 -187 796 -181
rect 856 -147 914 -141
rect 856 -181 868 -147
rect 902 -181 914 -147
rect 856 -187 914 -181
rect 974 -147 1032 -141
rect 974 -181 986 -147
rect 1020 -181 1032 -147
rect 974 -187 1032 -181
rect 1092 -147 1150 -141
rect 1092 -181 1104 -147
rect 1138 -181 1150 -147
rect 1092 -187 1150 -181
rect 1210 -147 1268 -141
rect 1210 -181 1222 -147
rect 1256 -181 1268 -147
rect 1210 -187 1268 -181
rect 1328 -147 1386 -141
rect 1328 -181 1340 -147
rect 1374 -181 1386 -147
rect 1328 -187 1386 -181
rect 1446 -147 1504 -141
rect 1446 -181 1458 -147
rect 1492 -181 1504 -147
rect 1446 -187 1504 -181
rect 1564 -147 1622 -141
rect 1564 -181 1576 -147
rect 1610 -181 1622 -147
rect 1564 -187 1622 -181
rect 1682 -147 1740 -141
rect 1682 -181 1694 -147
rect 1728 -181 1740 -147
rect 1682 -187 1740 -181
rect 1800 -147 1858 -141
rect 1800 -181 1812 -147
rect 1846 -181 1858 -147
rect 1800 -187 1858 -181
rect 1918 -147 1976 -141
rect 1918 -181 1930 -147
rect 1964 -181 1976 -147
rect 1918 -187 1976 -181
rect 2036 -147 2094 -141
rect 2036 -181 2048 -147
rect 2082 -181 2094 -147
rect 2036 -187 2094 -181
rect 2154 -147 2212 -141
rect 2154 -181 2166 -147
rect 2200 -181 2212 -147
rect 2154 -187 2212 -181
rect 2272 -147 2330 -141
rect 2272 -181 2284 -147
rect 2318 -181 2330 -147
rect 2272 -187 2330 -181
rect 2390 -147 2448 -141
rect 2390 -181 2402 -147
rect 2436 -181 2448 -147
rect 2390 -187 2448 -181
rect 2508 -147 2566 -141
rect 2508 -181 2520 -147
rect 2554 -181 2566 -147
rect 2508 -187 2566 -181
rect 2626 -147 2684 -141
rect 2626 -181 2638 -147
rect 2672 -181 2684 -147
rect 2626 -187 2684 -181
rect 2744 -147 2802 -141
rect 2744 -181 2756 -147
rect 2790 -181 2802 -147
rect 2744 -187 2802 -181
rect 2862 -147 2920 -141
rect 2862 -181 2874 -147
rect 2908 -181 2920 -147
rect 2862 -187 2920 -181
rect 2980 -147 3038 -141
rect 2980 -181 2992 -147
rect 3026 -181 3038 -147
rect 2980 -187 3038 -181
rect 3098 -147 3156 -141
rect 3098 -181 3110 -147
rect 3144 -181 3156 -147
rect 3098 -187 3156 -181
rect 3216 -147 3274 -141
rect 3216 -181 3228 -147
rect 3262 -181 3274 -147
rect 3216 -187 3274 -181
rect 3334 -147 3392 -141
rect 3334 -181 3346 -147
rect 3380 -181 3392 -147
rect 3334 -187 3392 -181
rect 3452 -147 3510 -141
rect 3452 -181 3464 -147
rect 3498 -181 3510 -147
rect 3452 -187 3510 -181
rect 3570 -147 3628 -141
rect 3570 -181 3582 -147
rect 3616 -181 3628 -147
rect 3570 -187 3628 -181
rect 3688 -147 3746 -141
rect 3688 -181 3700 -147
rect 3734 -181 3746 -147
rect 3688 -187 3746 -181
rect 3806 -147 3864 -141
rect 3806 -181 3818 -147
rect 3852 -181 3864 -147
rect 3806 -187 3864 -181
<< properties >>
string FIXED_BBOX -4008 -266 4008 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.3 m 1 nf 66 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
