magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< nwell >>
rect 428 0 760 490
<< poly >>
rect 77 155 136 185
rect 260 155 456 185
<< locali >>
rect 60 137 94 203
rect 165 103 742 137
<< metal1 >>
rect 184 0 212 395
rect 580 0 608 395
use sky130_sram_1r1w_24x128_8_contact_12  sky130_sram_1r1w_24x128_8_contact_12_0
timestamp 1661296025
transform 1 0 569 0 1 354
box -59 -43 109 125
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_0
timestamp 1661296025
transform 1 0 565 0 1 187
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_1
timestamp 1661296025
transform 1 0 169 0 1 187
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_2
timestamp 1661296025
transform 1 0 169 0 1 362
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_3
timestamp 1661296025
transform 1 0 565 0 1 362
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_14  sky130_sram_1r1w_24x128_8_contact_14_0
timestamp 1661296025
transform 1 0 173 0 1 354
box -26 -26 76 108
use sky130_sram_1r1w_24x128_8_contact_15  sky130_sram_1r1w_24x128_8_contact_15_0
timestamp 1661296025
transform 1 0 44 0 1 137
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_nmos_m1_w0_360_sli_dli_da_p  sky130_sram_1r1w_24x128_8_nmos_m1_w0_360_sli_dli_da_p_0
timestamp 1661296025
transform 0 1 162 -1 0 245
box -26 -26 176 98
use sky130_sram_1r1w_24x128_8_pmos_m1_w1_120_sli_dli_da_p  sky130_sram_1r1w_24x128_8_pmos_m1_w1_120_sli_dli_da_p_0
timestamp 1661296025
transform 0 1 482 -1 0 245
box -59 -54 209 278
<< labels >>
rlabel locali s 77 170 77 170 4 A
port 1 nsew
rlabel locali s 453 120 453 120 4 Z
port 2 nsew
rlabel metal1 s 184 0 212 395 4 gnd
port 3 nsew
rlabel metal1 s 580 0 608 395 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 742 395
<< end >>
