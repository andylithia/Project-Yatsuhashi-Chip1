magic
tech sky130A
magscale 1 2
timestamp 1664545297
<< pwell >>
rect -13400 43400 -8262 49916
rect -7100 43400 -1962 49916
rect -800 43400 4338 49916
rect 5500 43400 10638 49916
rect -13400 36400 -8262 42916
rect -7100 36400 -1962 42916
rect -800 36400 4338 42916
rect 5500 36400 10638 42916
rect -13400 28100 -8262 34616
rect -7100 28100 -1962 34616
rect -800 28100 4338 34616
rect 5500 28100 10638 34616
rect -13400 21100 -8262 27616
rect -7100 21100 -1962 27616
rect -800 21100 4338 27616
rect 5500 21100 10638 27616
rect -13400 12800 -8262 19316
rect -7100 12800 -1962 19316
rect -800 12800 4338 19316
rect 5500 12800 10638 19316
rect -13400 5800 -8262 12316
rect -7100 5800 -1962 12316
rect -800 5800 4338 12316
rect 5500 5800 10638 12316
<< mvnmos >>
rect -13172 43658 -13072 49658
rect -13014 43658 -12914 49658
rect -12856 43658 -12756 49658
rect -12698 43658 -12598 49658
rect -12540 43658 -12440 49658
rect -12382 43658 -12282 49658
rect -12224 43658 -12124 49658
rect -12066 43658 -11966 49658
rect -11908 43658 -11808 49658
rect -11750 43658 -11650 49658
rect -11592 43658 -11492 49658
rect -11434 43658 -11334 49658
rect -11276 43658 -11176 49658
rect -11118 43658 -11018 49658
rect -10960 43658 -10860 49658
rect -10802 43658 -10702 49658
rect -10644 43658 -10544 49658
rect -10486 43658 -10386 49658
rect -10328 43658 -10228 49658
rect -10170 43658 -10070 49658
rect -10012 43658 -9912 49658
rect -9854 43658 -9754 49658
rect -9696 43658 -9596 49658
rect -9538 43658 -9438 49658
rect -9380 43658 -9280 49658
rect -9222 43658 -9122 49658
rect -9064 43658 -8964 49658
rect -8906 43658 -8806 49658
rect -8748 43658 -8648 49658
rect -8590 43658 -8490 49658
rect -6872 43658 -6772 49658
rect -6714 43658 -6614 49658
rect -6556 43658 -6456 49658
rect -6398 43658 -6298 49658
rect -6240 43658 -6140 49658
rect -6082 43658 -5982 49658
rect -5924 43658 -5824 49658
rect -5766 43658 -5666 49658
rect -5608 43658 -5508 49658
rect -5450 43658 -5350 49658
rect -5292 43658 -5192 49658
rect -5134 43658 -5034 49658
rect -4976 43658 -4876 49658
rect -4818 43658 -4718 49658
rect -4660 43658 -4560 49658
rect -4502 43658 -4402 49658
rect -4344 43658 -4244 49658
rect -4186 43658 -4086 49658
rect -4028 43658 -3928 49658
rect -3870 43658 -3770 49658
rect -3712 43658 -3612 49658
rect -3554 43658 -3454 49658
rect -3396 43658 -3296 49658
rect -3238 43658 -3138 49658
rect -3080 43658 -2980 49658
rect -2922 43658 -2822 49658
rect -2764 43658 -2664 49658
rect -2606 43658 -2506 49658
rect -2448 43658 -2348 49658
rect -2290 43658 -2190 49658
rect -572 43658 -472 49658
rect -414 43658 -314 49658
rect -256 43658 -156 49658
rect -98 43658 2 49658
rect 60 43658 160 49658
rect 218 43658 318 49658
rect 376 43658 476 49658
rect 534 43658 634 49658
rect 692 43658 792 49658
rect 850 43658 950 49658
rect 1008 43658 1108 49658
rect 1166 43658 1266 49658
rect 1324 43658 1424 49658
rect 1482 43658 1582 49658
rect 1640 43658 1740 49658
rect 1798 43658 1898 49658
rect 1956 43658 2056 49658
rect 2114 43658 2214 49658
rect 2272 43658 2372 49658
rect 2430 43658 2530 49658
rect 2588 43658 2688 49658
rect 2746 43658 2846 49658
rect 2904 43658 3004 49658
rect 3062 43658 3162 49658
rect 3220 43658 3320 49658
rect 3378 43658 3478 49658
rect 3536 43658 3636 49658
rect 3694 43658 3794 49658
rect 3852 43658 3952 49658
rect 4010 43658 4110 49658
rect 5728 43658 5828 49658
rect 5886 43658 5986 49658
rect 6044 43658 6144 49658
rect 6202 43658 6302 49658
rect 6360 43658 6460 49658
rect 6518 43658 6618 49658
rect 6676 43658 6776 49658
rect 6834 43658 6934 49658
rect 6992 43658 7092 49658
rect 7150 43658 7250 49658
rect 7308 43658 7408 49658
rect 7466 43658 7566 49658
rect 7624 43658 7724 49658
rect 7782 43658 7882 49658
rect 7940 43658 8040 49658
rect 8098 43658 8198 49658
rect 8256 43658 8356 49658
rect 8414 43658 8514 49658
rect 8572 43658 8672 49658
rect 8730 43658 8830 49658
rect 8888 43658 8988 49658
rect 9046 43658 9146 49658
rect 9204 43658 9304 49658
rect 9362 43658 9462 49658
rect 9520 43658 9620 49658
rect 9678 43658 9778 49658
rect 9836 43658 9936 49658
rect 9994 43658 10094 49658
rect 10152 43658 10252 49658
rect 10310 43658 10410 49658
rect -13172 36658 -13072 42658
rect -13014 36658 -12914 42658
rect -12856 36658 -12756 42658
rect -12698 36658 -12598 42658
rect -12540 36658 -12440 42658
rect -12382 36658 -12282 42658
rect -12224 36658 -12124 42658
rect -12066 36658 -11966 42658
rect -11908 36658 -11808 42658
rect -11750 36658 -11650 42658
rect -11592 36658 -11492 42658
rect -11434 36658 -11334 42658
rect -11276 36658 -11176 42658
rect -11118 36658 -11018 42658
rect -10960 36658 -10860 42658
rect -10802 36658 -10702 42658
rect -10644 36658 -10544 42658
rect -10486 36658 -10386 42658
rect -10328 36658 -10228 42658
rect -10170 36658 -10070 42658
rect -10012 36658 -9912 42658
rect -9854 36658 -9754 42658
rect -9696 36658 -9596 42658
rect -9538 36658 -9438 42658
rect -9380 36658 -9280 42658
rect -9222 36658 -9122 42658
rect -9064 36658 -8964 42658
rect -8906 36658 -8806 42658
rect -8748 36658 -8648 42658
rect -8590 36658 -8490 42658
rect -6872 36658 -6772 42658
rect -6714 36658 -6614 42658
rect -6556 36658 -6456 42658
rect -6398 36658 -6298 42658
rect -6240 36658 -6140 42658
rect -6082 36658 -5982 42658
rect -5924 36658 -5824 42658
rect -5766 36658 -5666 42658
rect -5608 36658 -5508 42658
rect -5450 36658 -5350 42658
rect -5292 36658 -5192 42658
rect -5134 36658 -5034 42658
rect -4976 36658 -4876 42658
rect -4818 36658 -4718 42658
rect -4660 36658 -4560 42658
rect -4502 36658 -4402 42658
rect -4344 36658 -4244 42658
rect -4186 36658 -4086 42658
rect -4028 36658 -3928 42658
rect -3870 36658 -3770 42658
rect -3712 36658 -3612 42658
rect -3554 36658 -3454 42658
rect -3396 36658 -3296 42658
rect -3238 36658 -3138 42658
rect -3080 36658 -2980 42658
rect -2922 36658 -2822 42658
rect -2764 36658 -2664 42658
rect -2606 36658 -2506 42658
rect -2448 36658 -2348 42658
rect -2290 36658 -2190 42658
rect -572 36658 -472 42658
rect -414 36658 -314 42658
rect -256 36658 -156 42658
rect -98 36658 2 42658
rect 60 36658 160 42658
rect 218 36658 318 42658
rect 376 36658 476 42658
rect 534 36658 634 42658
rect 692 36658 792 42658
rect 850 36658 950 42658
rect 1008 36658 1108 42658
rect 1166 36658 1266 42658
rect 1324 36658 1424 42658
rect 1482 36658 1582 42658
rect 1640 36658 1740 42658
rect 1798 36658 1898 42658
rect 1956 36658 2056 42658
rect 2114 36658 2214 42658
rect 2272 36658 2372 42658
rect 2430 36658 2530 42658
rect 2588 36658 2688 42658
rect 2746 36658 2846 42658
rect 2904 36658 3004 42658
rect 3062 36658 3162 42658
rect 3220 36658 3320 42658
rect 3378 36658 3478 42658
rect 3536 36658 3636 42658
rect 3694 36658 3794 42658
rect 3852 36658 3952 42658
rect 4010 36658 4110 42658
rect 5728 36658 5828 42658
rect 5886 36658 5986 42658
rect 6044 36658 6144 42658
rect 6202 36658 6302 42658
rect 6360 36658 6460 42658
rect 6518 36658 6618 42658
rect 6676 36658 6776 42658
rect 6834 36658 6934 42658
rect 6992 36658 7092 42658
rect 7150 36658 7250 42658
rect 7308 36658 7408 42658
rect 7466 36658 7566 42658
rect 7624 36658 7724 42658
rect 7782 36658 7882 42658
rect 7940 36658 8040 42658
rect 8098 36658 8198 42658
rect 8256 36658 8356 42658
rect 8414 36658 8514 42658
rect 8572 36658 8672 42658
rect 8730 36658 8830 42658
rect 8888 36658 8988 42658
rect 9046 36658 9146 42658
rect 9204 36658 9304 42658
rect 9362 36658 9462 42658
rect 9520 36658 9620 42658
rect 9678 36658 9778 42658
rect 9836 36658 9936 42658
rect 9994 36658 10094 42658
rect 10152 36658 10252 42658
rect 10310 36658 10410 42658
rect -13172 28358 -13072 34358
rect -13014 28358 -12914 34358
rect -12856 28358 -12756 34358
rect -12698 28358 -12598 34358
rect -12540 28358 -12440 34358
rect -12382 28358 -12282 34358
rect -12224 28358 -12124 34358
rect -12066 28358 -11966 34358
rect -11908 28358 -11808 34358
rect -11750 28358 -11650 34358
rect -11592 28358 -11492 34358
rect -11434 28358 -11334 34358
rect -11276 28358 -11176 34358
rect -11118 28358 -11018 34358
rect -10960 28358 -10860 34358
rect -10802 28358 -10702 34358
rect -10644 28358 -10544 34358
rect -10486 28358 -10386 34358
rect -10328 28358 -10228 34358
rect -10170 28358 -10070 34358
rect -10012 28358 -9912 34358
rect -9854 28358 -9754 34358
rect -9696 28358 -9596 34358
rect -9538 28358 -9438 34358
rect -9380 28358 -9280 34358
rect -9222 28358 -9122 34358
rect -9064 28358 -8964 34358
rect -8906 28358 -8806 34358
rect -8748 28358 -8648 34358
rect -8590 28358 -8490 34358
rect -6872 28358 -6772 34358
rect -6714 28358 -6614 34358
rect -6556 28358 -6456 34358
rect -6398 28358 -6298 34358
rect -6240 28358 -6140 34358
rect -6082 28358 -5982 34358
rect -5924 28358 -5824 34358
rect -5766 28358 -5666 34358
rect -5608 28358 -5508 34358
rect -5450 28358 -5350 34358
rect -5292 28358 -5192 34358
rect -5134 28358 -5034 34358
rect -4976 28358 -4876 34358
rect -4818 28358 -4718 34358
rect -4660 28358 -4560 34358
rect -4502 28358 -4402 34358
rect -4344 28358 -4244 34358
rect -4186 28358 -4086 34358
rect -4028 28358 -3928 34358
rect -3870 28358 -3770 34358
rect -3712 28358 -3612 34358
rect -3554 28358 -3454 34358
rect -3396 28358 -3296 34358
rect -3238 28358 -3138 34358
rect -3080 28358 -2980 34358
rect -2922 28358 -2822 34358
rect -2764 28358 -2664 34358
rect -2606 28358 -2506 34358
rect -2448 28358 -2348 34358
rect -2290 28358 -2190 34358
rect -572 28358 -472 34358
rect -414 28358 -314 34358
rect -256 28358 -156 34358
rect -98 28358 2 34358
rect 60 28358 160 34358
rect 218 28358 318 34358
rect 376 28358 476 34358
rect 534 28358 634 34358
rect 692 28358 792 34358
rect 850 28358 950 34358
rect 1008 28358 1108 34358
rect 1166 28358 1266 34358
rect 1324 28358 1424 34358
rect 1482 28358 1582 34358
rect 1640 28358 1740 34358
rect 1798 28358 1898 34358
rect 1956 28358 2056 34358
rect 2114 28358 2214 34358
rect 2272 28358 2372 34358
rect 2430 28358 2530 34358
rect 2588 28358 2688 34358
rect 2746 28358 2846 34358
rect 2904 28358 3004 34358
rect 3062 28358 3162 34358
rect 3220 28358 3320 34358
rect 3378 28358 3478 34358
rect 3536 28358 3636 34358
rect 3694 28358 3794 34358
rect 3852 28358 3952 34358
rect 4010 28358 4110 34358
rect 5728 28358 5828 34358
rect 5886 28358 5986 34358
rect 6044 28358 6144 34358
rect 6202 28358 6302 34358
rect 6360 28358 6460 34358
rect 6518 28358 6618 34358
rect 6676 28358 6776 34358
rect 6834 28358 6934 34358
rect 6992 28358 7092 34358
rect 7150 28358 7250 34358
rect 7308 28358 7408 34358
rect 7466 28358 7566 34358
rect 7624 28358 7724 34358
rect 7782 28358 7882 34358
rect 7940 28358 8040 34358
rect 8098 28358 8198 34358
rect 8256 28358 8356 34358
rect 8414 28358 8514 34358
rect 8572 28358 8672 34358
rect 8730 28358 8830 34358
rect 8888 28358 8988 34358
rect 9046 28358 9146 34358
rect 9204 28358 9304 34358
rect 9362 28358 9462 34358
rect 9520 28358 9620 34358
rect 9678 28358 9778 34358
rect 9836 28358 9936 34358
rect 9994 28358 10094 34358
rect 10152 28358 10252 34358
rect 10310 28358 10410 34358
rect -13172 21358 -13072 27358
rect -13014 21358 -12914 27358
rect -12856 21358 -12756 27358
rect -12698 21358 -12598 27358
rect -12540 21358 -12440 27358
rect -12382 21358 -12282 27358
rect -12224 21358 -12124 27358
rect -12066 21358 -11966 27358
rect -11908 21358 -11808 27358
rect -11750 21358 -11650 27358
rect -11592 21358 -11492 27358
rect -11434 21358 -11334 27358
rect -11276 21358 -11176 27358
rect -11118 21358 -11018 27358
rect -10960 21358 -10860 27358
rect -10802 21358 -10702 27358
rect -10644 21358 -10544 27358
rect -10486 21358 -10386 27358
rect -10328 21358 -10228 27358
rect -10170 21358 -10070 27358
rect -10012 21358 -9912 27358
rect -9854 21358 -9754 27358
rect -9696 21358 -9596 27358
rect -9538 21358 -9438 27358
rect -9380 21358 -9280 27358
rect -9222 21358 -9122 27358
rect -9064 21358 -8964 27358
rect -8906 21358 -8806 27358
rect -8748 21358 -8648 27358
rect -8590 21358 -8490 27358
rect -6872 21358 -6772 27358
rect -6714 21358 -6614 27358
rect -6556 21358 -6456 27358
rect -6398 21358 -6298 27358
rect -6240 21358 -6140 27358
rect -6082 21358 -5982 27358
rect -5924 21358 -5824 27358
rect -5766 21358 -5666 27358
rect -5608 21358 -5508 27358
rect -5450 21358 -5350 27358
rect -5292 21358 -5192 27358
rect -5134 21358 -5034 27358
rect -4976 21358 -4876 27358
rect -4818 21358 -4718 27358
rect -4660 21358 -4560 27358
rect -4502 21358 -4402 27358
rect -4344 21358 -4244 27358
rect -4186 21358 -4086 27358
rect -4028 21358 -3928 27358
rect -3870 21358 -3770 27358
rect -3712 21358 -3612 27358
rect -3554 21358 -3454 27358
rect -3396 21358 -3296 27358
rect -3238 21358 -3138 27358
rect -3080 21358 -2980 27358
rect -2922 21358 -2822 27358
rect -2764 21358 -2664 27358
rect -2606 21358 -2506 27358
rect -2448 21358 -2348 27358
rect -2290 21358 -2190 27358
rect -572 21358 -472 27358
rect -414 21358 -314 27358
rect -256 21358 -156 27358
rect -98 21358 2 27358
rect 60 21358 160 27358
rect 218 21358 318 27358
rect 376 21358 476 27358
rect 534 21358 634 27358
rect 692 21358 792 27358
rect 850 21358 950 27358
rect 1008 21358 1108 27358
rect 1166 21358 1266 27358
rect 1324 21358 1424 27358
rect 1482 21358 1582 27358
rect 1640 21358 1740 27358
rect 1798 21358 1898 27358
rect 1956 21358 2056 27358
rect 2114 21358 2214 27358
rect 2272 21358 2372 27358
rect 2430 21358 2530 27358
rect 2588 21358 2688 27358
rect 2746 21358 2846 27358
rect 2904 21358 3004 27358
rect 3062 21358 3162 27358
rect 3220 21358 3320 27358
rect 3378 21358 3478 27358
rect 3536 21358 3636 27358
rect 3694 21358 3794 27358
rect 3852 21358 3952 27358
rect 4010 21358 4110 27358
rect 5728 21358 5828 27358
rect 5886 21358 5986 27358
rect 6044 21358 6144 27358
rect 6202 21358 6302 27358
rect 6360 21358 6460 27358
rect 6518 21358 6618 27358
rect 6676 21358 6776 27358
rect 6834 21358 6934 27358
rect 6992 21358 7092 27358
rect 7150 21358 7250 27358
rect 7308 21358 7408 27358
rect 7466 21358 7566 27358
rect 7624 21358 7724 27358
rect 7782 21358 7882 27358
rect 7940 21358 8040 27358
rect 8098 21358 8198 27358
rect 8256 21358 8356 27358
rect 8414 21358 8514 27358
rect 8572 21358 8672 27358
rect 8730 21358 8830 27358
rect 8888 21358 8988 27358
rect 9046 21358 9146 27358
rect 9204 21358 9304 27358
rect 9362 21358 9462 27358
rect 9520 21358 9620 27358
rect 9678 21358 9778 27358
rect 9836 21358 9936 27358
rect 9994 21358 10094 27358
rect 10152 21358 10252 27358
rect 10310 21358 10410 27358
rect -13172 13058 -13072 19058
rect -13014 13058 -12914 19058
rect -12856 13058 -12756 19058
rect -12698 13058 -12598 19058
rect -12540 13058 -12440 19058
rect -12382 13058 -12282 19058
rect -12224 13058 -12124 19058
rect -12066 13058 -11966 19058
rect -11908 13058 -11808 19058
rect -11750 13058 -11650 19058
rect -11592 13058 -11492 19058
rect -11434 13058 -11334 19058
rect -11276 13058 -11176 19058
rect -11118 13058 -11018 19058
rect -10960 13058 -10860 19058
rect -10802 13058 -10702 19058
rect -10644 13058 -10544 19058
rect -10486 13058 -10386 19058
rect -10328 13058 -10228 19058
rect -10170 13058 -10070 19058
rect -10012 13058 -9912 19058
rect -9854 13058 -9754 19058
rect -9696 13058 -9596 19058
rect -9538 13058 -9438 19058
rect -9380 13058 -9280 19058
rect -9222 13058 -9122 19058
rect -9064 13058 -8964 19058
rect -8906 13058 -8806 19058
rect -8748 13058 -8648 19058
rect -8590 13058 -8490 19058
rect -6872 13058 -6772 19058
rect -6714 13058 -6614 19058
rect -6556 13058 -6456 19058
rect -6398 13058 -6298 19058
rect -6240 13058 -6140 19058
rect -6082 13058 -5982 19058
rect -5924 13058 -5824 19058
rect -5766 13058 -5666 19058
rect -5608 13058 -5508 19058
rect -5450 13058 -5350 19058
rect -5292 13058 -5192 19058
rect -5134 13058 -5034 19058
rect -4976 13058 -4876 19058
rect -4818 13058 -4718 19058
rect -4660 13058 -4560 19058
rect -4502 13058 -4402 19058
rect -4344 13058 -4244 19058
rect -4186 13058 -4086 19058
rect -4028 13058 -3928 19058
rect -3870 13058 -3770 19058
rect -3712 13058 -3612 19058
rect -3554 13058 -3454 19058
rect -3396 13058 -3296 19058
rect -3238 13058 -3138 19058
rect -3080 13058 -2980 19058
rect -2922 13058 -2822 19058
rect -2764 13058 -2664 19058
rect -2606 13058 -2506 19058
rect -2448 13058 -2348 19058
rect -2290 13058 -2190 19058
rect -572 13058 -472 19058
rect -414 13058 -314 19058
rect -256 13058 -156 19058
rect -98 13058 2 19058
rect 60 13058 160 19058
rect 218 13058 318 19058
rect 376 13058 476 19058
rect 534 13058 634 19058
rect 692 13058 792 19058
rect 850 13058 950 19058
rect 1008 13058 1108 19058
rect 1166 13058 1266 19058
rect 1324 13058 1424 19058
rect 1482 13058 1582 19058
rect 1640 13058 1740 19058
rect 1798 13058 1898 19058
rect 1956 13058 2056 19058
rect 2114 13058 2214 19058
rect 2272 13058 2372 19058
rect 2430 13058 2530 19058
rect 2588 13058 2688 19058
rect 2746 13058 2846 19058
rect 2904 13058 3004 19058
rect 3062 13058 3162 19058
rect 3220 13058 3320 19058
rect 3378 13058 3478 19058
rect 3536 13058 3636 19058
rect 3694 13058 3794 19058
rect 3852 13058 3952 19058
rect 4010 13058 4110 19058
rect 5728 13058 5828 19058
rect 5886 13058 5986 19058
rect 6044 13058 6144 19058
rect 6202 13058 6302 19058
rect 6360 13058 6460 19058
rect 6518 13058 6618 19058
rect 6676 13058 6776 19058
rect 6834 13058 6934 19058
rect 6992 13058 7092 19058
rect 7150 13058 7250 19058
rect 7308 13058 7408 19058
rect 7466 13058 7566 19058
rect 7624 13058 7724 19058
rect 7782 13058 7882 19058
rect 7940 13058 8040 19058
rect 8098 13058 8198 19058
rect 8256 13058 8356 19058
rect 8414 13058 8514 19058
rect 8572 13058 8672 19058
rect 8730 13058 8830 19058
rect 8888 13058 8988 19058
rect 9046 13058 9146 19058
rect 9204 13058 9304 19058
rect 9362 13058 9462 19058
rect 9520 13058 9620 19058
rect 9678 13058 9778 19058
rect 9836 13058 9936 19058
rect 9994 13058 10094 19058
rect 10152 13058 10252 19058
rect 10310 13058 10410 19058
rect -13172 6058 -13072 12058
rect -13014 6058 -12914 12058
rect -12856 6058 -12756 12058
rect -12698 6058 -12598 12058
rect -12540 6058 -12440 12058
rect -12382 6058 -12282 12058
rect -12224 6058 -12124 12058
rect -12066 6058 -11966 12058
rect -11908 6058 -11808 12058
rect -11750 6058 -11650 12058
rect -11592 6058 -11492 12058
rect -11434 6058 -11334 12058
rect -11276 6058 -11176 12058
rect -11118 6058 -11018 12058
rect -10960 6058 -10860 12058
rect -10802 6058 -10702 12058
rect -10644 6058 -10544 12058
rect -10486 6058 -10386 12058
rect -10328 6058 -10228 12058
rect -10170 6058 -10070 12058
rect -10012 6058 -9912 12058
rect -9854 6058 -9754 12058
rect -9696 6058 -9596 12058
rect -9538 6058 -9438 12058
rect -9380 6058 -9280 12058
rect -9222 6058 -9122 12058
rect -9064 6058 -8964 12058
rect -8906 6058 -8806 12058
rect -8748 6058 -8648 12058
rect -8590 6058 -8490 12058
rect -6872 6058 -6772 12058
rect -6714 6058 -6614 12058
rect -6556 6058 -6456 12058
rect -6398 6058 -6298 12058
rect -6240 6058 -6140 12058
rect -6082 6058 -5982 12058
rect -5924 6058 -5824 12058
rect -5766 6058 -5666 12058
rect -5608 6058 -5508 12058
rect -5450 6058 -5350 12058
rect -5292 6058 -5192 12058
rect -5134 6058 -5034 12058
rect -4976 6058 -4876 12058
rect -4818 6058 -4718 12058
rect -4660 6058 -4560 12058
rect -4502 6058 -4402 12058
rect -4344 6058 -4244 12058
rect -4186 6058 -4086 12058
rect -4028 6058 -3928 12058
rect -3870 6058 -3770 12058
rect -3712 6058 -3612 12058
rect -3554 6058 -3454 12058
rect -3396 6058 -3296 12058
rect -3238 6058 -3138 12058
rect -3080 6058 -2980 12058
rect -2922 6058 -2822 12058
rect -2764 6058 -2664 12058
rect -2606 6058 -2506 12058
rect -2448 6058 -2348 12058
rect -2290 6058 -2190 12058
rect -572 6058 -472 12058
rect -414 6058 -314 12058
rect -256 6058 -156 12058
rect -98 6058 2 12058
rect 60 6058 160 12058
rect 218 6058 318 12058
rect 376 6058 476 12058
rect 534 6058 634 12058
rect 692 6058 792 12058
rect 850 6058 950 12058
rect 1008 6058 1108 12058
rect 1166 6058 1266 12058
rect 1324 6058 1424 12058
rect 1482 6058 1582 12058
rect 1640 6058 1740 12058
rect 1798 6058 1898 12058
rect 1956 6058 2056 12058
rect 2114 6058 2214 12058
rect 2272 6058 2372 12058
rect 2430 6058 2530 12058
rect 2588 6058 2688 12058
rect 2746 6058 2846 12058
rect 2904 6058 3004 12058
rect 3062 6058 3162 12058
rect 3220 6058 3320 12058
rect 3378 6058 3478 12058
rect 3536 6058 3636 12058
rect 3694 6058 3794 12058
rect 3852 6058 3952 12058
rect 4010 6058 4110 12058
rect 5728 6058 5828 12058
rect 5886 6058 5986 12058
rect 6044 6058 6144 12058
rect 6202 6058 6302 12058
rect 6360 6058 6460 12058
rect 6518 6058 6618 12058
rect 6676 6058 6776 12058
rect 6834 6058 6934 12058
rect 6992 6058 7092 12058
rect 7150 6058 7250 12058
rect 7308 6058 7408 12058
rect 7466 6058 7566 12058
rect 7624 6058 7724 12058
rect 7782 6058 7882 12058
rect 7940 6058 8040 12058
rect 8098 6058 8198 12058
rect 8256 6058 8356 12058
rect 8414 6058 8514 12058
rect 8572 6058 8672 12058
rect 8730 6058 8830 12058
rect 8888 6058 8988 12058
rect 9046 6058 9146 12058
rect 9204 6058 9304 12058
rect 9362 6058 9462 12058
rect 9520 6058 9620 12058
rect 9678 6058 9778 12058
rect 9836 6058 9936 12058
rect 9994 6058 10094 12058
rect 10152 6058 10252 12058
rect 10310 6058 10410 12058
<< mvndiff >>
rect -13230 49646 -13172 49658
rect -13230 43670 -13218 49646
rect -13184 43670 -13172 49646
rect -13230 43658 -13172 43670
rect -13072 49646 -13014 49658
rect -13072 43670 -13060 49646
rect -13026 43670 -13014 49646
rect -13072 43658 -13014 43670
rect -12914 49646 -12856 49658
rect -12914 43670 -12902 49646
rect -12868 43670 -12856 49646
rect -12914 43658 -12856 43670
rect -12756 49646 -12698 49658
rect -12756 43670 -12744 49646
rect -12710 43670 -12698 49646
rect -12756 43658 -12698 43670
rect -12598 49646 -12540 49658
rect -12598 43670 -12586 49646
rect -12552 43670 -12540 49646
rect -12598 43658 -12540 43670
rect -12440 49646 -12382 49658
rect -12440 43670 -12428 49646
rect -12394 43670 -12382 49646
rect -12440 43658 -12382 43670
rect -12282 49646 -12224 49658
rect -12282 43670 -12270 49646
rect -12236 43670 -12224 49646
rect -12282 43658 -12224 43670
rect -12124 49646 -12066 49658
rect -12124 43670 -12112 49646
rect -12078 43670 -12066 49646
rect -12124 43658 -12066 43670
rect -11966 49646 -11908 49658
rect -11966 43670 -11954 49646
rect -11920 43670 -11908 49646
rect -11966 43658 -11908 43670
rect -11808 49646 -11750 49658
rect -11808 43670 -11796 49646
rect -11762 43670 -11750 49646
rect -11808 43658 -11750 43670
rect -11650 49646 -11592 49658
rect -11650 43670 -11638 49646
rect -11604 43670 -11592 49646
rect -11650 43658 -11592 43670
rect -11492 49646 -11434 49658
rect -11492 43670 -11480 49646
rect -11446 43670 -11434 49646
rect -11492 43658 -11434 43670
rect -11334 49646 -11276 49658
rect -11334 43670 -11322 49646
rect -11288 43670 -11276 49646
rect -11334 43658 -11276 43670
rect -11176 49646 -11118 49658
rect -11176 43670 -11164 49646
rect -11130 43670 -11118 49646
rect -11176 43658 -11118 43670
rect -11018 49646 -10960 49658
rect -11018 43670 -11006 49646
rect -10972 43670 -10960 49646
rect -11018 43658 -10960 43670
rect -10860 49646 -10802 49658
rect -10860 43670 -10848 49646
rect -10814 43670 -10802 49646
rect -10860 43658 -10802 43670
rect -10702 49646 -10644 49658
rect -10702 43670 -10690 49646
rect -10656 43670 -10644 49646
rect -10702 43658 -10644 43670
rect -10544 49646 -10486 49658
rect -10544 43670 -10532 49646
rect -10498 43670 -10486 49646
rect -10544 43658 -10486 43670
rect -10386 49646 -10328 49658
rect -10386 43670 -10374 49646
rect -10340 43670 -10328 49646
rect -10386 43658 -10328 43670
rect -10228 49646 -10170 49658
rect -10228 43670 -10216 49646
rect -10182 43670 -10170 49646
rect -10228 43658 -10170 43670
rect -10070 49646 -10012 49658
rect -10070 43670 -10058 49646
rect -10024 43670 -10012 49646
rect -10070 43658 -10012 43670
rect -9912 49646 -9854 49658
rect -9912 43670 -9900 49646
rect -9866 43670 -9854 49646
rect -9912 43658 -9854 43670
rect -9754 49646 -9696 49658
rect -9754 43670 -9742 49646
rect -9708 43670 -9696 49646
rect -9754 43658 -9696 43670
rect -9596 49646 -9538 49658
rect -9596 43670 -9584 49646
rect -9550 43670 -9538 49646
rect -9596 43658 -9538 43670
rect -9438 49646 -9380 49658
rect -9438 43670 -9426 49646
rect -9392 43670 -9380 49646
rect -9438 43658 -9380 43670
rect -9280 49646 -9222 49658
rect -9280 43670 -9268 49646
rect -9234 43670 -9222 49646
rect -9280 43658 -9222 43670
rect -9122 49646 -9064 49658
rect -9122 43670 -9110 49646
rect -9076 43670 -9064 49646
rect -9122 43658 -9064 43670
rect -8964 49646 -8906 49658
rect -8964 43670 -8952 49646
rect -8918 43670 -8906 49646
rect -8964 43658 -8906 43670
rect -8806 49646 -8748 49658
rect -8806 43670 -8794 49646
rect -8760 43670 -8748 49646
rect -8806 43658 -8748 43670
rect -8648 49646 -8590 49658
rect -8648 43670 -8636 49646
rect -8602 43670 -8590 49646
rect -8648 43658 -8590 43670
rect -8490 49646 -8432 49658
rect -8490 43670 -8478 49646
rect -8444 43670 -8432 49646
rect -8490 43658 -8432 43670
rect -6930 49646 -6872 49658
rect -6930 43670 -6918 49646
rect -6884 43670 -6872 49646
rect -6930 43658 -6872 43670
rect -6772 49646 -6714 49658
rect -6772 43670 -6760 49646
rect -6726 43670 -6714 49646
rect -6772 43658 -6714 43670
rect -6614 49646 -6556 49658
rect -6614 43670 -6602 49646
rect -6568 43670 -6556 49646
rect -6614 43658 -6556 43670
rect -6456 49646 -6398 49658
rect -6456 43670 -6444 49646
rect -6410 43670 -6398 49646
rect -6456 43658 -6398 43670
rect -6298 49646 -6240 49658
rect -6298 43670 -6286 49646
rect -6252 43670 -6240 49646
rect -6298 43658 -6240 43670
rect -6140 49646 -6082 49658
rect -6140 43670 -6128 49646
rect -6094 43670 -6082 49646
rect -6140 43658 -6082 43670
rect -5982 49646 -5924 49658
rect -5982 43670 -5970 49646
rect -5936 43670 -5924 49646
rect -5982 43658 -5924 43670
rect -5824 49646 -5766 49658
rect -5824 43670 -5812 49646
rect -5778 43670 -5766 49646
rect -5824 43658 -5766 43670
rect -5666 49646 -5608 49658
rect -5666 43670 -5654 49646
rect -5620 43670 -5608 49646
rect -5666 43658 -5608 43670
rect -5508 49646 -5450 49658
rect -5508 43670 -5496 49646
rect -5462 43670 -5450 49646
rect -5508 43658 -5450 43670
rect -5350 49646 -5292 49658
rect -5350 43670 -5338 49646
rect -5304 43670 -5292 49646
rect -5350 43658 -5292 43670
rect -5192 49646 -5134 49658
rect -5192 43670 -5180 49646
rect -5146 43670 -5134 49646
rect -5192 43658 -5134 43670
rect -5034 49646 -4976 49658
rect -5034 43670 -5022 49646
rect -4988 43670 -4976 49646
rect -5034 43658 -4976 43670
rect -4876 49646 -4818 49658
rect -4876 43670 -4864 49646
rect -4830 43670 -4818 49646
rect -4876 43658 -4818 43670
rect -4718 49646 -4660 49658
rect -4718 43670 -4706 49646
rect -4672 43670 -4660 49646
rect -4718 43658 -4660 43670
rect -4560 49646 -4502 49658
rect -4560 43670 -4548 49646
rect -4514 43670 -4502 49646
rect -4560 43658 -4502 43670
rect -4402 49646 -4344 49658
rect -4402 43670 -4390 49646
rect -4356 43670 -4344 49646
rect -4402 43658 -4344 43670
rect -4244 49646 -4186 49658
rect -4244 43670 -4232 49646
rect -4198 43670 -4186 49646
rect -4244 43658 -4186 43670
rect -4086 49646 -4028 49658
rect -4086 43670 -4074 49646
rect -4040 43670 -4028 49646
rect -4086 43658 -4028 43670
rect -3928 49646 -3870 49658
rect -3928 43670 -3916 49646
rect -3882 43670 -3870 49646
rect -3928 43658 -3870 43670
rect -3770 49646 -3712 49658
rect -3770 43670 -3758 49646
rect -3724 43670 -3712 49646
rect -3770 43658 -3712 43670
rect -3612 49646 -3554 49658
rect -3612 43670 -3600 49646
rect -3566 43670 -3554 49646
rect -3612 43658 -3554 43670
rect -3454 49646 -3396 49658
rect -3454 43670 -3442 49646
rect -3408 43670 -3396 49646
rect -3454 43658 -3396 43670
rect -3296 49646 -3238 49658
rect -3296 43670 -3284 49646
rect -3250 43670 -3238 49646
rect -3296 43658 -3238 43670
rect -3138 49646 -3080 49658
rect -3138 43670 -3126 49646
rect -3092 43670 -3080 49646
rect -3138 43658 -3080 43670
rect -2980 49646 -2922 49658
rect -2980 43670 -2968 49646
rect -2934 43670 -2922 49646
rect -2980 43658 -2922 43670
rect -2822 49646 -2764 49658
rect -2822 43670 -2810 49646
rect -2776 43670 -2764 49646
rect -2822 43658 -2764 43670
rect -2664 49646 -2606 49658
rect -2664 43670 -2652 49646
rect -2618 43670 -2606 49646
rect -2664 43658 -2606 43670
rect -2506 49646 -2448 49658
rect -2506 43670 -2494 49646
rect -2460 43670 -2448 49646
rect -2506 43658 -2448 43670
rect -2348 49646 -2290 49658
rect -2348 43670 -2336 49646
rect -2302 43670 -2290 49646
rect -2348 43658 -2290 43670
rect -2190 49646 -2132 49658
rect -2190 43670 -2178 49646
rect -2144 43670 -2132 49646
rect -2190 43658 -2132 43670
rect -630 49646 -572 49658
rect -630 43670 -618 49646
rect -584 43670 -572 49646
rect -630 43658 -572 43670
rect -472 49646 -414 49658
rect -472 43670 -460 49646
rect -426 43670 -414 49646
rect -472 43658 -414 43670
rect -314 49646 -256 49658
rect -314 43670 -302 49646
rect -268 43670 -256 49646
rect -314 43658 -256 43670
rect -156 49646 -98 49658
rect -156 43670 -144 49646
rect -110 43670 -98 49646
rect -156 43658 -98 43670
rect 2 49646 60 49658
rect 2 43670 14 49646
rect 48 43670 60 49646
rect 2 43658 60 43670
rect 160 49646 218 49658
rect 160 43670 172 49646
rect 206 43670 218 49646
rect 160 43658 218 43670
rect 318 49646 376 49658
rect 318 43670 330 49646
rect 364 43670 376 49646
rect 318 43658 376 43670
rect 476 49646 534 49658
rect 476 43670 488 49646
rect 522 43670 534 49646
rect 476 43658 534 43670
rect 634 49646 692 49658
rect 634 43670 646 49646
rect 680 43670 692 49646
rect 634 43658 692 43670
rect 792 49646 850 49658
rect 792 43670 804 49646
rect 838 43670 850 49646
rect 792 43658 850 43670
rect 950 49646 1008 49658
rect 950 43670 962 49646
rect 996 43670 1008 49646
rect 950 43658 1008 43670
rect 1108 49646 1166 49658
rect 1108 43670 1120 49646
rect 1154 43670 1166 49646
rect 1108 43658 1166 43670
rect 1266 49646 1324 49658
rect 1266 43670 1278 49646
rect 1312 43670 1324 49646
rect 1266 43658 1324 43670
rect 1424 49646 1482 49658
rect 1424 43670 1436 49646
rect 1470 43670 1482 49646
rect 1424 43658 1482 43670
rect 1582 49646 1640 49658
rect 1582 43670 1594 49646
rect 1628 43670 1640 49646
rect 1582 43658 1640 43670
rect 1740 49646 1798 49658
rect 1740 43670 1752 49646
rect 1786 43670 1798 49646
rect 1740 43658 1798 43670
rect 1898 49646 1956 49658
rect 1898 43670 1910 49646
rect 1944 43670 1956 49646
rect 1898 43658 1956 43670
rect 2056 49646 2114 49658
rect 2056 43670 2068 49646
rect 2102 43670 2114 49646
rect 2056 43658 2114 43670
rect 2214 49646 2272 49658
rect 2214 43670 2226 49646
rect 2260 43670 2272 49646
rect 2214 43658 2272 43670
rect 2372 49646 2430 49658
rect 2372 43670 2384 49646
rect 2418 43670 2430 49646
rect 2372 43658 2430 43670
rect 2530 49646 2588 49658
rect 2530 43670 2542 49646
rect 2576 43670 2588 49646
rect 2530 43658 2588 43670
rect 2688 49646 2746 49658
rect 2688 43670 2700 49646
rect 2734 43670 2746 49646
rect 2688 43658 2746 43670
rect 2846 49646 2904 49658
rect 2846 43670 2858 49646
rect 2892 43670 2904 49646
rect 2846 43658 2904 43670
rect 3004 49646 3062 49658
rect 3004 43670 3016 49646
rect 3050 43670 3062 49646
rect 3004 43658 3062 43670
rect 3162 49646 3220 49658
rect 3162 43670 3174 49646
rect 3208 43670 3220 49646
rect 3162 43658 3220 43670
rect 3320 49646 3378 49658
rect 3320 43670 3332 49646
rect 3366 43670 3378 49646
rect 3320 43658 3378 43670
rect 3478 49646 3536 49658
rect 3478 43670 3490 49646
rect 3524 43670 3536 49646
rect 3478 43658 3536 43670
rect 3636 49646 3694 49658
rect 3636 43670 3648 49646
rect 3682 43670 3694 49646
rect 3636 43658 3694 43670
rect 3794 49646 3852 49658
rect 3794 43670 3806 49646
rect 3840 43670 3852 49646
rect 3794 43658 3852 43670
rect 3952 49646 4010 49658
rect 3952 43670 3964 49646
rect 3998 43670 4010 49646
rect 3952 43658 4010 43670
rect 4110 49646 4168 49658
rect 4110 43670 4122 49646
rect 4156 43670 4168 49646
rect 4110 43658 4168 43670
rect 5670 49646 5728 49658
rect 5670 43670 5682 49646
rect 5716 43670 5728 49646
rect 5670 43658 5728 43670
rect 5828 49646 5886 49658
rect 5828 43670 5840 49646
rect 5874 43670 5886 49646
rect 5828 43658 5886 43670
rect 5986 49646 6044 49658
rect 5986 43670 5998 49646
rect 6032 43670 6044 49646
rect 5986 43658 6044 43670
rect 6144 49646 6202 49658
rect 6144 43670 6156 49646
rect 6190 43670 6202 49646
rect 6144 43658 6202 43670
rect 6302 49646 6360 49658
rect 6302 43670 6314 49646
rect 6348 43670 6360 49646
rect 6302 43658 6360 43670
rect 6460 49646 6518 49658
rect 6460 43670 6472 49646
rect 6506 43670 6518 49646
rect 6460 43658 6518 43670
rect 6618 49646 6676 49658
rect 6618 43670 6630 49646
rect 6664 43670 6676 49646
rect 6618 43658 6676 43670
rect 6776 49646 6834 49658
rect 6776 43670 6788 49646
rect 6822 43670 6834 49646
rect 6776 43658 6834 43670
rect 6934 49646 6992 49658
rect 6934 43670 6946 49646
rect 6980 43670 6992 49646
rect 6934 43658 6992 43670
rect 7092 49646 7150 49658
rect 7092 43670 7104 49646
rect 7138 43670 7150 49646
rect 7092 43658 7150 43670
rect 7250 49646 7308 49658
rect 7250 43670 7262 49646
rect 7296 43670 7308 49646
rect 7250 43658 7308 43670
rect 7408 49646 7466 49658
rect 7408 43670 7420 49646
rect 7454 43670 7466 49646
rect 7408 43658 7466 43670
rect 7566 49646 7624 49658
rect 7566 43670 7578 49646
rect 7612 43670 7624 49646
rect 7566 43658 7624 43670
rect 7724 49646 7782 49658
rect 7724 43670 7736 49646
rect 7770 43670 7782 49646
rect 7724 43658 7782 43670
rect 7882 49646 7940 49658
rect 7882 43670 7894 49646
rect 7928 43670 7940 49646
rect 7882 43658 7940 43670
rect 8040 49646 8098 49658
rect 8040 43670 8052 49646
rect 8086 43670 8098 49646
rect 8040 43658 8098 43670
rect 8198 49646 8256 49658
rect 8198 43670 8210 49646
rect 8244 43670 8256 49646
rect 8198 43658 8256 43670
rect 8356 49646 8414 49658
rect 8356 43670 8368 49646
rect 8402 43670 8414 49646
rect 8356 43658 8414 43670
rect 8514 49646 8572 49658
rect 8514 43670 8526 49646
rect 8560 43670 8572 49646
rect 8514 43658 8572 43670
rect 8672 49646 8730 49658
rect 8672 43670 8684 49646
rect 8718 43670 8730 49646
rect 8672 43658 8730 43670
rect 8830 49646 8888 49658
rect 8830 43670 8842 49646
rect 8876 43670 8888 49646
rect 8830 43658 8888 43670
rect 8988 49646 9046 49658
rect 8988 43670 9000 49646
rect 9034 43670 9046 49646
rect 8988 43658 9046 43670
rect 9146 49646 9204 49658
rect 9146 43670 9158 49646
rect 9192 43670 9204 49646
rect 9146 43658 9204 43670
rect 9304 49646 9362 49658
rect 9304 43670 9316 49646
rect 9350 43670 9362 49646
rect 9304 43658 9362 43670
rect 9462 49646 9520 49658
rect 9462 43670 9474 49646
rect 9508 43670 9520 49646
rect 9462 43658 9520 43670
rect 9620 49646 9678 49658
rect 9620 43670 9632 49646
rect 9666 43670 9678 49646
rect 9620 43658 9678 43670
rect 9778 49646 9836 49658
rect 9778 43670 9790 49646
rect 9824 43670 9836 49646
rect 9778 43658 9836 43670
rect 9936 49646 9994 49658
rect 9936 43670 9948 49646
rect 9982 43670 9994 49646
rect 9936 43658 9994 43670
rect 10094 49646 10152 49658
rect 10094 43670 10106 49646
rect 10140 43670 10152 49646
rect 10094 43658 10152 43670
rect 10252 49646 10310 49658
rect 10252 43670 10264 49646
rect 10298 43670 10310 49646
rect 10252 43658 10310 43670
rect 10410 49646 10468 49658
rect 10410 43670 10422 49646
rect 10456 43670 10468 49646
rect 10410 43658 10468 43670
rect -13230 42646 -13172 42658
rect -13230 36670 -13218 42646
rect -13184 36670 -13172 42646
rect -13230 36658 -13172 36670
rect -13072 42646 -13014 42658
rect -13072 36670 -13060 42646
rect -13026 36670 -13014 42646
rect -13072 36658 -13014 36670
rect -12914 42646 -12856 42658
rect -12914 36670 -12902 42646
rect -12868 36670 -12856 42646
rect -12914 36658 -12856 36670
rect -12756 42646 -12698 42658
rect -12756 36670 -12744 42646
rect -12710 36670 -12698 42646
rect -12756 36658 -12698 36670
rect -12598 42646 -12540 42658
rect -12598 36670 -12586 42646
rect -12552 36670 -12540 42646
rect -12598 36658 -12540 36670
rect -12440 42646 -12382 42658
rect -12440 36670 -12428 42646
rect -12394 36670 -12382 42646
rect -12440 36658 -12382 36670
rect -12282 42646 -12224 42658
rect -12282 36670 -12270 42646
rect -12236 36670 -12224 42646
rect -12282 36658 -12224 36670
rect -12124 42646 -12066 42658
rect -12124 36670 -12112 42646
rect -12078 36670 -12066 42646
rect -12124 36658 -12066 36670
rect -11966 42646 -11908 42658
rect -11966 36670 -11954 42646
rect -11920 36670 -11908 42646
rect -11966 36658 -11908 36670
rect -11808 42646 -11750 42658
rect -11808 36670 -11796 42646
rect -11762 36670 -11750 42646
rect -11808 36658 -11750 36670
rect -11650 42646 -11592 42658
rect -11650 36670 -11638 42646
rect -11604 36670 -11592 42646
rect -11650 36658 -11592 36670
rect -11492 42646 -11434 42658
rect -11492 36670 -11480 42646
rect -11446 36670 -11434 42646
rect -11492 36658 -11434 36670
rect -11334 42646 -11276 42658
rect -11334 36670 -11322 42646
rect -11288 36670 -11276 42646
rect -11334 36658 -11276 36670
rect -11176 42646 -11118 42658
rect -11176 36670 -11164 42646
rect -11130 36670 -11118 42646
rect -11176 36658 -11118 36670
rect -11018 42646 -10960 42658
rect -11018 36670 -11006 42646
rect -10972 36670 -10960 42646
rect -11018 36658 -10960 36670
rect -10860 42646 -10802 42658
rect -10860 36670 -10848 42646
rect -10814 36670 -10802 42646
rect -10860 36658 -10802 36670
rect -10702 42646 -10644 42658
rect -10702 36670 -10690 42646
rect -10656 36670 -10644 42646
rect -10702 36658 -10644 36670
rect -10544 42646 -10486 42658
rect -10544 36670 -10532 42646
rect -10498 36670 -10486 42646
rect -10544 36658 -10486 36670
rect -10386 42646 -10328 42658
rect -10386 36670 -10374 42646
rect -10340 36670 -10328 42646
rect -10386 36658 -10328 36670
rect -10228 42646 -10170 42658
rect -10228 36670 -10216 42646
rect -10182 36670 -10170 42646
rect -10228 36658 -10170 36670
rect -10070 42646 -10012 42658
rect -10070 36670 -10058 42646
rect -10024 36670 -10012 42646
rect -10070 36658 -10012 36670
rect -9912 42646 -9854 42658
rect -9912 36670 -9900 42646
rect -9866 36670 -9854 42646
rect -9912 36658 -9854 36670
rect -9754 42646 -9696 42658
rect -9754 36670 -9742 42646
rect -9708 36670 -9696 42646
rect -9754 36658 -9696 36670
rect -9596 42646 -9538 42658
rect -9596 36670 -9584 42646
rect -9550 36670 -9538 42646
rect -9596 36658 -9538 36670
rect -9438 42646 -9380 42658
rect -9438 36670 -9426 42646
rect -9392 36670 -9380 42646
rect -9438 36658 -9380 36670
rect -9280 42646 -9222 42658
rect -9280 36670 -9268 42646
rect -9234 36670 -9222 42646
rect -9280 36658 -9222 36670
rect -9122 42646 -9064 42658
rect -9122 36670 -9110 42646
rect -9076 36670 -9064 42646
rect -9122 36658 -9064 36670
rect -8964 42646 -8906 42658
rect -8964 36670 -8952 42646
rect -8918 36670 -8906 42646
rect -8964 36658 -8906 36670
rect -8806 42646 -8748 42658
rect -8806 36670 -8794 42646
rect -8760 36670 -8748 42646
rect -8806 36658 -8748 36670
rect -8648 42646 -8590 42658
rect -8648 36670 -8636 42646
rect -8602 36670 -8590 42646
rect -8648 36658 -8590 36670
rect -8490 42646 -8432 42658
rect -8490 36670 -8478 42646
rect -8444 36670 -8432 42646
rect -8490 36658 -8432 36670
rect -6930 42646 -6872 42658
rect -6930 36670 -6918 42646
rect -6884 36670 -6872 42646
rect -6930 36658 -6872 36670
rect -6772 42646 -6714 42658
rect -6772 36670 -6760 42646
rect -6726 36670 -6714 42646
rect -6772 36658 -6714 36670
rect -6614 42646 -6556 42658
rect -6614 36670 -6602 42646
rect -6568 36670 -6556 42646
rect -6614 36658 -6556 36670
rect -6456 42646 -6398 42658
rect -6456 36670 -6444 42646
rect -6410 36670 -6398 42646
rect -6456 36658 -6398 36670
rect -6298 42646 -6240 42658
rect -6298 36670 -6286 42646
rect -6252 36670 -6240 42646
rect -6298 36658 -6240 36670
rect -6140 42646 -6082 42658
rect -6140 36670 -6128 42646
rect -6094 36670 -6082 42646
rect -6140 36658 -6082 36670
rect -5982 42646 -5924 42658
rect -5982 36670 -5970 42646
rect -5936 36670 -5924 42646
rect -5982 36658 -5924 36670
rect -5824 42646 -5766 42658
rect -5824 36670 -5812 42646
rect -5778 36670 -5766 42646
rect -5824 36658 -5766 36670
rect -5666 42646 -5608 42658
rect -5666 36670 -5654 42646
rect -5620 36670 -5608 42646
rect -5666 36658 -5608 36670
rect -5508 42646 -5450 42658
rect -5508 36670 -5496 42646
rect -5462 36670 -5450 42646
rect -5508 36658 -5450 36670
rect -5350 42646 -5292 42658
rect -5350 36670 -5338 42646
rect -5304 36670 -5292 42646
rect -5350 36658 -5292 36670
rect -5192 42646 -5134 42658
rect -5192 36670 -5180 42646
rect -5146 36670 -5134 42646
rect -5192 36658 -5134 36670
rect -5034 42646 -4976 42658
rect -5034 36670 -5022 42646
rect -4988 36670 -4976 42646
rect -5034 36658 -4976 36670
rect -4876 42646 -4818 42658
rect -4876 36670 -4864 42646
rect -4830 36670 -4818 42646
rect -4876 36658 -4818 36670
rect -4718 42646 -4660 42658
rect -4718 36670 -4706 42646
rect -4672 36670 -4660 42646
rect -4718 36658 -4660 36670
rect -4560 42646 -4502 42658
rect -4560 36670 -4548 42646
rect -4514 36670 -4502 42646
rect -4560 36658 -4502 36670
rect -4402 42646 -4344 42658
rect -4402 36670 -4390 42646
rect -4356 36670 -4344 42646
rect -4402 36658 -4344 36670
rect -4244 42646 -4186 42658
rect -4244 36670 -4232 42646
rect -4198 36670 -4186 42646
rect -4244 36658 -4186 36670
rect -4086 42646 -4028 42658
rect -4086 36670 -4074 42646
rect -4040 36670 -4028 42646
rect -4086 36658 -4028 36670
rect -3928 42646 -3870 42658
rect -3928 36670 -3916 42646
rect -3882 36670 -3870 42646
rect -3928 36658 -3870 36670
rect -3770 42646 -3712 42658
rect -3770 36670 -3758 42646
rect -3724 36670 -3712 42646
rect -3770 36658 -3712 36670
rect -3612 42646 -3554 42658
rect -3612 36670 -3600 42646
rect -3566 36670 -3554 42646
rect -3612 36658 -3554 36670
rect -3454 42646 -3396 42658
rect -3454 36670 -3442 42646
rect -3408 36670 -3396 42646
rect -3454 36658 -3396 36670
rect -3296 42646 -3238 42658
rect -3296 36670 -3284 42646
rect -3250 36670 -3238 42646
rect -3296 36658 -3238 36670
rect -3138 42646 -3080 42658
rect -3138 36670 -3126 42646
rect -3092 36670 -3080 42646
rect -3138 36658 -3080 36670
rect -2980 42646 -2922 42658
rect -2980 36670 -2968 42646
rect -2934 36670 -2922 42646
rect -2980 36658 -2922 36670
rect -2822 42646 -2764 42658
rect -2822 36670 -2810 42646
rect -2776 36670 -2764 42646
rect -2822 36658 -2764 36670
rect -2664 42646 -2606 42658
rect -2664 36670 -2652 42646
rect -2618 36670 -2606 42646
rect -2664 36658 -2606 36670
rect -2506 42646 -2448 42658
rect -2506 36670 -2494 42646
rect -2460 36670 -2448 42646
rect -2506 36658 -2448 36670
rect -2348 42646 -2290 42658
rect -2348 36670 -2336 42646
rect -2302 36670 -2290 42646
rect -2348 36658 -2290 36670
rect -2190 42646 -2132 42658
rect -2190 36670 -2178 42646
rect -2144 36670 -2132 42646
rect -2190 36658 -2132 36670
rect -630 42646 -572 42658
rect -630 36670 -618 42646
rect -584 36670 -572 42646
rect -630 36658 -572 36670
rect -472 42646 -414 42658
rect -472 36670 -460 42646
rect -426 36670 -414 42646
rect -472 36658 -414 36670
rect -314 42646 -256 42658
rect -314 36670 -302 42646
rect -268 36670 -256 42646
rect -314 36658 -256 36670
rect -156 42646 -98 42658
rect -156 36670 -144 42646
rect -110 36670 -98 42646
rect -156 36658 -98 36670
rect 2 42646 60 42658
rect 2 36670 14 42646
rect 48 36670 60 42646
rect 2 36658 60 36670
rect 160 42646 218 42658
rect 160 36670 172 42646
rect 206 36670 218 42646
rect 160 36658 218 36670
rect 318 42646 376 42658
rect 318 36670 330 42646
rect 364 36670 376 42646
rect 318 36658 376 36670
rect 476 42646 534 42658
rect 476 36670 488 42646
rect 522 36670 534 42646
rect 476 36658 534 36670
rect 634 42646 692 42658
rect 634 36670 646 42646
rect 680 36670 692 42646
rect 634 36658 692 36670
rect 792 42646 850 42658
rect 792 36670 804 42646
rect 838 36670 850 42646
rect 792 36658 850 36670
rect 950 42646 1008 42658
rect 950 36670 962 42646
rect 996 36670 1008 42646
rect 950 36658 1008 36670
rect 1108 42646 1166 42658
rect 1108 36670 1120 42646
rect 1154 36670 1166 42646
rect 1108 36658 1166 36670
rect 1266 42646 1324 42658
rect 1266 36670 1278 42646
rect 1312 36670 1324 42646
rect 1266 36658 1324 36670
rect 1424 42646 1482 42658
rect 1424 36670 1436 42646
rect 1470 36670 1482 42646
rect 1424 36658 1482 36670
rect 1582 42646 1640 42658
rect 1582 36670 1594 42646
rect 1628 36670 1640 42646
rect 1582 36658 1640 36670
rect 1740 42646 1798 42658
rect 1740 36670 1752 42646
rect 1786 36670 1798 42646
rect 1740 36658 1798 36670
rect 1898 42646 1956 42658
rect 1898 36670 1910 42646
rect 1944 36670 1956 42646
rect 1898 36658 1956 36670
rect 2056 42646 2114 42658
rect 2056 36670 2068 42646
rect 2102 36670 2114 42646
rect 2056 36658 2114 36670
rect 2214 42646 2272 42658
rect 2214 36670 2226 42646
rect 2260 36670 2272 42646
rect 2214 36658 2272 36670
rect 2372 42646 2430 42658
rect 2372 36670 2384 42646
rect 2418 36670 2430 42646
rect 2372 36658 2430 36670
rect 2530 42646 2588 42658
rect 2530 36670 2542 42646
rect 2576 36670 2588 42646
rect 2530 36658 2588 36670
rect 2688 42646 2746 42658
rect 2688 36670 2700 42646
rect 2734 36670 2746 42646
rect 2688 36658 2746 36670
rect 2846 42646 2904 42658
rect 2846 36670 2858 42646
rect 2892 36670 2904 42646
rect 2846 36658 2904 36670
rect 3004 42646 3062 42658
rect 3004 36670 3016 42646
rect 3050 36670 3062 42646
rect 3004 36658 3062 36670
rect 3162 42646 3220 42658
rect 3162 36670 3174 42646
rect 3208 36670 3220 42646
rect 3162 36658 3220 36670
rect 3320 42646 3378 42658
rect 3320 36670 3332 42646
rect 3366 36670 3378 42646
rect 3320 36658 3378 36670
rect 3478 42646 3536 42658
rect 3478 36670 3490 42646
rect 3524 36670 3536 42646
rect 3478 36658 3536 36670
rect 3636 42646 3694 42658
rect 3636 36670 3648 42646
rect 3682 36670 3694 42646
rect 3636 36658 3694 36670
rect 3794 42646 3852 42658
rect 3794 36670 3806 42646
rect 3840 36670 3852 42646
rect 3794 36658 3852 36670
rect 3952 42646 4010 42658
rect 3952 36670 3964 42646
rect 3998 36670 4010 42646
rect 3952 36658 4010 36670
rect 4110 42646 4168 42658
rect 4110 36670 4122 42646
rect 4156 36670 4168 42646
rect 4110 36658 4168 36670
rect 5670 42646 5728 42658
rect 5670 36670 5682 42646
rect 5716 36670 5728 42646
rect 5670 36658 5728 36670
rect 5828 42646 5886 42658
rect 5828 36670 5840 42646
rect 5874 36670 5886 42646
rect 5828 36658 5886 36670
rect 5986 42646 6044 42658
rect 5986 36670 5998 42646
rect 6032 36670 6044 42646
rect 5986 36658 6044 36670
rect 6144 42646 6202 42658
rect 6144 36670 6156 42646
rect 6190 36670 6202 42646
rect 6144 36658 6202 36670
rect 6302 42646 6360 42658
rect 6302 36670 6314 42646
rect 6348 36670 6360 42646
rect 6302 36658 6360 36670
rect 6460 42646 6518 42658
rect 6460 36670 6472 42646
rect 6506 36670 6518 42646
rect 6460 36658 6518 36670
rect 6618 42646 6676 42658
rect 6618 36670 6630 42646
rect 6664 36670 6676 42646
rect 6618 36658 6676 36670
rect 6776 42646 6834 42658
rect 6776 36670 6788 42646
rect 6822 36670 6834 42646
rect 6776 36658 6834 36670
rect 6934 42646 6992 42658
rect 6934 36670 6946 42646
rect 6980 36670 6992 42646
rect 6934 36658 6992 36670
rect 7092 42646 7150 42658
rect 7092 36670 7104 42646
rect 7138 36670 7150 42646
rect 7092 36658 7150 36670
rect 7250 42646 7308 42658
rect 7250 36670 7262 42646
rect 7296 36670 7308 42646
rect 7250 36658 7308 36670
rect 7408 42646 7466 42658
rect 7408 36670 7420 42646
rect 7454 36670 7466 42646
rect 7408 36658 7466 36670
rect 7566 42646 7624 42658
rect 7566 36670 7578 42646
rect 7612 36670 7624 42646
rect 7566 36658 7624 36670
rect 7724 42646 7782 42658
rect 7724 36670 7736 42646
rect 7770 36670 7782 42646
rect 7724 36658 7782 36670
rect 7882 42646 7940 42658
rect 7882 36670 7894 42646
rect 7928 36670 7940 42646
rect 7882 36658 7940 36670
rect 8040 42646 8098 42658
rect 8040 36670 8052 42646
rect 8086 36670 8098 42646
rect 8040 36658 8098 36670
rect 8198 42646 8256 42658
rect 8198 36670 8210 42646
rect 8244 36670 8256 42646
rect 8198 36658 8256 36670
rect 8356 42646 8414 42658
rect 8356 36670 8368 42646
rect 8402 36670 8414 42646
rect 8356 36658 8414 36670
rect 8514 42646 8572 42658
rect 8514 36670 8526 42646
rect 8560 36670 8572 42646
rect 8514 36658 8572 36670
rect 8672 42646 8730 42658
rect 8672 36670 8684 42646
rect 8718 36670 8730 42646
rect 8672 36658 8730 36670
rect 8830 42646 8888 42658
rect 8830 36670 8842 42646
rect 8876 36670 8888 42646
rect 8830 36658 8888 36670
rect 8988 42646 9046 42658
rect 8988 36670 9000 42646
rect 9034 36670 9046 42646
rect 8988 36658 9046 36670
rect 9146 42646 9204 42658
rect 9146 36670 9158 42646
rect 9192 36670 9204 42646
rect 9146 36658 9204 36670
rect 9304 42646 9362 42658
rect 9304 36670 9316 42646
rect 9350 36670 9362 42646
rect 9304 36658 9362 36670
rect 9462 42646 9520 42658
rect 9462 36670 9474 42646
rect 9508 36670 9520 42646
rect 9462 36658 9520 36670
rect 9620 42646 9678 42658
rect 9620 36670 9632 42646
rect 9666 36670 9678 42646
rect 9620 36658 9678 36670
rect 9778 42646 9836 42658
rect 9778 36670 9790 42646
rect 9824 36670 9836 42646
rect 9778 36658 9836 36670
rect 9936 42646 9994 42658
rect 9936 36670 9948 42646
rect 9982 36670 9994 42646
rect 9936 36658 9994 36670
rect 10094 42646 10152 42658
rect 10094 36670 10106 42646
rect 10140 36670 10152 42646
rect 10094 36658 10152 36670
rect 10252 42646 10310 42658
rect 10252 36670 10264 42646
rect 10298 36670 10310 42646
rect 10252 36658 10310 36670
rect 10410 42646 10468 42658
rect 10410 36670 10422 42646
rect 10456 36670 10468 42646
rect 10410 36658 10468 36670
rect -13230 34346 -13172 34358
rect -13230 28370 -13218 34346
rect -13184 28370 -13172 34346
rect -13230 28358 -13172 28370
rect -13072 34346 -13014 34358
rect -13072 28370 -13060 34346
rect -13026 28370 -13014 34346
rect -13072 28358 -13014 28370
rect -12914 34346 -12856 34358
rect -12914 28370 -12902 34346
rect -12868 28370 -12856 34346
rect -12914 28358 -12856 28370
rect -12756 34346 -12698 34358
rect -12756 28370 -12744 34346
rect -12710 28370 -12698 34346
rect -12756 28358 -12698 28370
rect -12598 34346 -12540 34358
rect -12598 28370 -12586 34346
rect -12552 28370 -12540 34346
rect -12598 28358 -12540 28370
rect -12440 34346 -12382 34358
rect -12440 28370 -12428 34346
rect -12394 28370 -12382 34346
rect -12440 28358 -12382 28370
rect -12282 34346 -12224 34358
rect -12282 28370 -12270 34346
rect -12236 28370 -12224 34346
rect -12282 28358 -12224 28370
rect -12124 34346 -12066 34358
rect -12124 28370 -12112 34346
rect -12078 28370 -12066 34346
rect -12124 28358 -12066 28370
rect -11966 34346 -11908 34358
rect -11966 28370 -11954 34346
rect -11920 28370 -11908 34346
rect -11966 28358 -11908 28370
rect -11808 34346 -11750 34358
rect -11808 28370 -11796 34346
rect -11762 28370 -11750 34346
rect -11808 28358 -11750 28370
rect -11650 34346 -11592 34358
rect -11650 28370 -11638 34346
rect -11604 28370 -11592 34346
rect -11650 28358 -11592 28370
rect -11492 34346 -11434 34358
rect -11492 28370 -11480 34346
rect -11446 28370 -11434 34346
rect -11492 28358 -11434 28370
rect -11334 34346 -11276 34358
rect -11334 28370 -11322 34346
rect -11288 28370 -11276 34346
rect -11334 28358 -11276 28370
rect -11176 34346 -11118 34358
rect -11176 28370 -11164 34346
rect -11130 28370 -11118 34346
rect -11176 28358 -11118 28370
rect -11018 34346 -10960 34358
rect -11018 28370 -11006 34346
rect -10972 28370 -10960 34346
rect -11018 28358 -10960 28370
rect -10860 34346 -10802 34358
rect -10860 28370 -10848 34346
rect -10814 28370 -10802 34346
rect -10860 28358 -10802 28370
rect -10702 34346 -10644 34358
rect -10702 28370 -10690 34346
rect -10656 28370 -10644 34346
rect -10702 28358 -10644 28370
rect -10544 34346 -10486 34358
rect -10544 28370 -10532 34346
rect -10498 28370 -10486 34346
rect -10544 28358 -10486 28370
rect -10386 34346 -10328 34358
rect -10386 28370 -10374 34346
rect -10340 28370 -10328 34346
rect -10386 28358 -10328 28370
rect -10228 34346 -10170 34358
rect -10228 28370 -10216 34346
rect -10182 28370 -10170 34346
rect -10228 28358 -10170 28370
rect -10070 34346 -10012 34358
rect -10070 28370 -10058 34346
rect -10024 28370 -10012 34346
rect -10070 28358 -10012 28370
rect -9912 34346 -9854 34358
rect -9912 28370 -9900 34346
rect -9866 28370 -9854 34346
rect -9912 28358 -9854 28370
rect -9754 34346 -9696 34358
rect -9754 28370 -9742 34346
rect -9708 28370 -9696 34346
rect -9754 28358 -9696 28370
rect -9596 34346 -9538 34358
rect -9596 28370 -9584 34346
rect -9550 28370 -9538 34346
rect -9596 28358 -9538 28370
rect -9438 34346 -9380 34358
rect -9438 28370 -9426 34346
rect -9392 28370 -9380 34346
rect -9438 28358 -9380 28370
rect -9280 34346 -9222 34358
rect -9280 28370 -9268 34346
rect -9234 28370 -9222 34346
rect -9280 28358 -9222 28370
rect -9122 34346 -9064 34358
rect -9122 28370 -9110 34346
rect -9076 28370 -9064 34346
rect -9122 28358 -9064 28370
rect -8964 34346 -8906 34358
rect -8964 28370 -8952 34346
rect -8918 28370 -8906 34346
rect -8964 28358 -8906 28370
rect -8806 34346 -8748 34358
rect -8806 28370 -8794 34346
rect -8760 28370 -8748 34346
rect -8806 28358 -8748 28370
rect -8648 34346 -8590 34358
rect -8648 28370 -8636 34346
rect -8602 28370 -8590 34346
rect -8648 28358 -8590 28370
rect -8490 34346 -8432 34358
rect -8490 28370 -8478 34346
rect -8444 28370 -8432 34346
rect -8490 28358 -8432 28370
rect -6930 34346 -6872 34358
rect -6930 28370 -6918 34346
rect -6884 28370 -6872 34346
rect -6930 28358 -6872 28370
rect -6772 34346 -6714 34358
rect -6772 28370 -6760 34346
rect -6726 28370 -6714 34346
rect -6772 28358 -6714 28370
rect -6614 34346 -6556 34358
rect -6614 28370 -6602 34346
rect -6568 28370 -6556 34346
rect -6614 28358 -6556 28370
rect -6456 34346 -6398 34358
rect -6456 28370 -6444 34346
rect -6410 28370 -6398 34346
rect -6456 28358 -6398 28370
rect -6298 34346 -6240 34358
rect -6298 28370 -6286 34346
rect -6252 28370 -6240 34346
rect -6298 28358 -6240 28370
rect -6140 34346 -6082 34358
rect -6140 28370 -6128 34346
rect -6094 28370 -6082 34346
rect -6140 28358 -6082 28370
rect -5982 34346 -5924 34358
rect -5982 28370 -5970 34346
rect -5936 28370 -5924 34346
rect -5982 28358 -5924 28370
rect -5824 34346 -5766 34358
rect -5824 28370 -5812 34346
rect -5778 28370 -5766 34346
rect -5824 28358 -5766 28370
rect -5666 34346 -5608 34358
rect -5666 28370 -5654 34346
rect -5620 28370 -5608 34346
rect -5666 28358 -5608 28370
rect -5508 34346 -5450 34358
rect -5508 28370 -5496 34346
rect -5462 28370 -5450 34346
rect -5508 28358 -5450 28370
rect -5350 34346 -5292 34358
rect -5350 28370 -5338 34346
rect -5304 28370 -5292 34346
rect -5350 28358 -5292 28370
rect -5192 34346 -5134 34358
rect -5192 28370 -5180 34346
rect -5146 28370 -5134 34346
rect -5192 28358 -5134 28370
rect -5034 34346 -4976 34358
rect -5034 28370 -5022 34346
rect -4988 28370 -4976 34346
rect -5034 28358 -4976 28370
rect -4876 34346 -4818 34358
rect -4876 28370 -4864 34346
rect -4830 28370 -4818 34346
rect -4876 28358 -4818 28370
rect -4718 34346 -4660 34358
rect -4718 28370 -4706 34346
rect -4672 28370 -4660 34346
rect -4718 28358 -4660 28370
rect -4560 34346 -4502 34358
rect -4560 28370 -4548 34346
rect -4514 28370 -4502 34346
rect -4560 28358 -4502 28370
rect -4402 34346 -4344 34358
rect -4402 28370 -4390 34346
rect -4356 28370 -4344 34346
rect -4402 28358 -4344 28370
rect -4244 34346 -4186 34358
rect -4244 28370 -4232 34346
rect -4198 28370 -4186 34346
rect -4244 28358 -4186 28370
rect -4086 34346 -4028 34358
rect -4086 28370 -4074 34346
rect -4040 28370 -4028 34346
rect -4086 28358 -4028 28370
rect -3928 34346 -3870 34358
rect -3928 28370 -3916 34346
rect -3882 28370 -3870 34346
rect -3928 28358 -3870 28370
rect -3770 34346 -3712 34358
rect -3770 28370 -3758 34346
rect -3724 28370 -3712 34346
rect -3770 28358 -3712 28370
rect -3612 34346 -3554 34358
rect -3612 28370 -3600 34346
rect -3566 28370 -3554 34346
rect -3612 28358 -3554 28370
rect -3454 34346 -3396 34358
rect -3454 28370 -3442 34346
rect -3408 28370 -3396 34346
rect -3454 28358 -3396 28370
rect -3296 34346 -3238 34358
rect -3296 28370 -3284 34346
rect -3250 28370 -3238 34346
rect -3296 28358 -3238 28370
rect -3138 34346 -3080 34358
rect -3138 28370 -3126 34346
rect -3092 28370 -3080 34346
rect -3138 28358 -3080 28370
rect -2980 34346 -2922 34358
rect -2980 28370 -2968 34346
rect -2934 28370 -2922 34346
rect -2980 28358 -2922 28370
rect -2822 34346 -2764 34358
rect -2822 28370 -2810 34346
rect -2776 28370 -2764 34346
rect -2822 28358 -2764 28370
rect -2664 34346 -2606 34358
rect -2664 28370 -2652 34346
rect -2618 28370 -2606 34346
rect -2664 28358 -2606 28370
rect -2506 34346 -2448 34358
rect -2506 28370 -2494 34346
rect -2460 28370 -2448 34346
rect -2506 28358 -2448 28370
rect -2348 34346 -2290 34358
rect -2348 28370 -2336 34346
rect -2302 28370 -2290 34346
rect -2348 28358 -2290 28370
rect -2190 34346 -2132 34358
rect -2190 28370 -2178 34346
rect -2144 28370 -2132 34346
rect -2190 28358 -2132 28370
rect -630 34346 -572 34358
rect -630 28370 -618 34346
rect -584 28370 -572 34346
rect -630 28358 -572 28370
rect -472 34346 -414 34358
rect -472 28370 -460 34346
rect -426 28370 -414 34346
rect -472 28358 -414 28370
rect -314 34346 -256 34358
rect -314 28370 -302 34346
rect -268 28370 -256 34346
rect -314 28358 -256 28370
rect -156 34346 -98 34358
rect -156 28370 -144 34346
rect -110 28370 -98 34346
rect -156 28358 -98 28370
rect 2 34346 60 34358
rect 2 28370 14 34346
rect 48 28370 60 34346
rect 2 28358 60 28370
rect 160 34346 218 34358
rect 160 28370 172 34346
rect 206 28370 218 34346
rect 160 28358 218 28370
rect 318 34346 376 34358
rect 318 28370 330 34346
rect 364 28370 376 34346
rect 318 28358 376 28370
rect 476 34346 534 34358
rect 476 28370 488 34346
rect 522 28370 534 34346
rect 476 28358 534 28370
rect 634 34346 692 34358
rect 634 28370 646 34346
rect 680 28370 692 34346
rect 634 28358 692 28370
rect 792 34346 850 34358
rect 792 28370 804 34346
rect 838 28370 850 34346
rect 792 28358 850 28370
rect 950 34346 1008 34358
rect 950 28370 962 34346
rect 996 28370 1008 34346
rect 950 28358 1008 28370
rect 1108 34346 1166 34358
rect 1108 28370 1120 34346
rect 1154 28370 1166 34346
rect 1108 28358 1166 28370
rect 1266 34346 1324 34358
rect 1266 28370 1278 34346
rect 1312 28370 1324 34346
rect 1266 28358 1324 28370
rect 1424 34346 1482 34358
rect 1424 28370 1436 34346
rect 1470 28370 1482 34346
rect 1424 28358 1482 28370
rect 1582 34346 1640 34358
rect 1582 28370 1594 34346
rect 1628 28370 1640 34346
rect 1582 28358 1640 28370
rect 1740 34346 1798 34358
rect 1740 28370 1752 34346
rect 1786 28370 1798 34346
rect 1740 28358 1798 28370
rect 1898 34346 1956 34358
rect 1898 28370 1910 34346
rect 1944 28370 1956 34346
rect 1898 28358 1956 28370
rect 2056 34346 2114 34358
rect 2056 28370 2068 34346
rect 2102 28370 2114 34346
rect 2056 28358 2114 28370
rect 2214 34346 2272 34358
rect 2214 28370 2226 34346
rect 2260 28370 2272 34346
rect 2214 28358 2272 28370
rect 2372 34346 2430 34358
rect 2372 28370 2384 34346
rect 2418 28370 2430 34346
rect 2372 28358 2430 28370
rect 2530 34346 2588 34358
rect 2530 28370 2542 34346
rect 2576 28370 2588 34346
rect 2530 28358 2588 28370
rect 2688 34346 2746 34358
rect 2688 28370 2700 34346
rect 2734 28370 2746 34346
rect 2688 28358 2746 28370
rect 2846 34346 2904 34358
rect 2846 28370 2858 34346
rect 2892 28370 2904 34346
rect 2846 28358 2904 28370
rect 3004 34346 3062 34358
rect 3004 28370 3016 34346
rect 3050 28370 3062 34346
rect 3004 28358 3062 28370
rect 3162 34346 3220 34358
rect 3162 28370 3174 34346
rect 3208 28370 3220 34346
rect 3162 28358 3220 28370
rect 3320 34346 3378 34358
rect 3320 28370 3332 34346
rect 3366 28370 3378 34346
rect 3320 28358 3378 28370
rect 3478 34346 3536 34358
rect 3478 28370 3490 34346
rect 3524 28370 3536 34346
rect 3478 28358 3536 28370
rect 3636 34346 3694 34358
rect 3636 28370 3648 34346
rect 3682 28370 3694 34346
rect 3636 28358 3694 28370
rect 3794 34346 3852 34358
rect 3794 28370 3806 34346
rect 3840 28370 3852 34346
rect 3794 28358 3852 28370
rect 3952 34346 4010 34358
rect 3952 28370 3964 34346
rect 3998 28370 4010 34346
rect 3952 28358 4010 28370
rect 4110 34346 4168 34358
rect 4110 28370 4122 34346
rect 4156 28370 4168 34346
rect 4110 28358 4168 28370
rect 5670 34346 5728 34358
rect 5670 28370 5682 34346
rect 5716 28370 5728 34346
rect 5670 28358 5728 28370
rect 5828 34346 5886 34358
rect 5828 28370 5840 34346
rect 5874 28370 5886 34346
rect 5828 28358 5886 28370
rect 5986 34346 6044 34358
rect 5986 28370 5998 34346
rect 6032 28370 6044 34346
rect 5986 28358 6044 28370
rect 6144 34346 6202 34358
rect 6144 28370 6156 34346
rect 6190 28370 6202 34346
rect 6144 28358 6202 28370
rect 6302 34346 6360 34358
rect 6302 28370 6314 34346
rect 6348 28370 6360 34346
rect 6302 28358 6360 28370
rect 6460 34346 6518 34358
rect 6460 28370 6472 34346
rect 6506 28370 6518 34346
rect 6460 28358 6518 28370
rect 6618 34346 6676 34358
rect 6618 28370 6630 34346
rect 6664 28370 6676 34346
rect 6618 28358 6676 28370
rect 6776 34346 6834 34358
rect 6776 28370 6788 34346
rect 6822 28370 6834 34346
rect 6776 28358 6834 28370
rect 6934 34346 6992 34358
rect 6934 28370 6946 34346
rect 6980 28370 6992 34346
rect 6934 28358 6992 28370
rect 7092 34346 7150 34358
rect 7092 28370 7104 34346
rect 7138 28370 7150 34346
rect 7092 28358 7150 28370
rect 7250 34346 7308 34358
rect 7250 28370 7262 34346
rect 7296 28370 7308 34346
rect 7250 28358 7308 28370
rect 7408 34346 7466 34358
rect 7408 28370 7420 34346
rect 7454 28370 7466 34346
rect 7408 28358 7466 28370
rect 7566 34346 7624 34358
rect 7566 28370 7578 34346
rect 7612 28370 7624 34346
rect 7566 28358 7624 28370
rect 7724 34346 7782 34358
rect 7724 28370 7736 34346
rect 7770 28370 7782 34346
rect 7724 28358 7782 28370
rect 7882 34346 7940 34358
rect 7882 28370 7894 34346
rect 7928 28370 7940 34346
rect 7882 28358 7940 28370
rect 8040 34346 8098 34358
rect 8040 28370 8052 34346
rect 8086 28370 8098 34346
rect 8040 28358 8098 28370
rect 8198 34346 8256 34358
rect 8198 28370 8210 34346
rect 8244 28370 8256 34346
rect 8198 28358 8256 28370
rect 8356 34346 8414 34358
rect 8356 28370 8368 34346
rect 8402 28370 8414 34346
rect 8356 28358 8414 28370
rect 8514 34346 8572 34358
rect 8514 28370 8526 34346
rect 8560 28370 8572 34346
rect 8514 28358 8572 28370
rect 8672 34346 8730 34358
rect 8672 28370 8684 34346
rect 8718 28370 8730 34346
rect 8672 28358 8730 28370
rect 8830 34346 8888 34358
rect 8830 28370 8842 34346
rect 8876 28370 8888 34346
rect 8830 28358 8888 28370
rect 8988 34346 9046 34358
rect 8988 28370 9000 34346
rect 9034 28370 9046 34346
rect 8988 28358 9046 28370
rect 9146 34346 9204 34358
rect 9146 28370 9158 34346
rect 9192 28370 9204 34346
rect 9146 28358 9204 28370
rect 9304 34346 9362 34358
rect 9304 28370 9316 34346
rect 9350 28370 9362 34346
rect 9304 28358 9362 28370
rect 9462 34346 9520 34358
rect 9462 28370 9474 34346
rect 9508 28370 9520 34346
rect 9462 28358 9520 28370
rect 9620 34346 9678 34358
rect 9620 28370 9632 34346
rect 9666 28370 9678 34346
rect 9620 28358 9678 28370
rect 9778 34346 9836 34358
rect 9778 28370 9790 34346
rect 9824 28370 9836 34346
rect 9778 28358 9836 28370
rect 9936 34346 9994 34358
rect 9936 28370 9948 34346
rect 9982 28370 9994 34346
rect 9936 28358 9994 28370
rect 10094 34346 10152 34358
rect 10094 28370 10106 34346
rect 10140 28370 10152 34346
rect 10094 28358 10152 28370
rect 10252 34346 10310 34358
rect 10252 28370 10264 34346
rect 10298 28370 10310 34346
rect 10252 28358 10310 28370
rect 10410 34346 10468 34358
rect 10410 28370 10422 34346
rect 10456 28370 10468 34346
rect 10410 28358 10468 28370
rect -13230 27346 -13172 27358
rect -13230 21370 -13218 27346
rect -13184 21370 -13172 27346
rect -13230 21358 -13172 21370
rect -13072 27346 -13014 27358
rect -13072 21370 -13060 27346
rect -13026 21370 -13014 27346
rect -13072 21358 -13014 21370
rect -12914 27346 -12856 27358
rect -12914 21370 -12902 27346
rect -12868 21370 -12856 27346
rect -12914 21358 -12856 21370
rect -12756 27346 -12698 27358
rect -12756 21370 -12744 27346
rect -12710 21370 -12698 27346
rect -12756 21358 -12698 21370
rect -12598 27346 -12540 27358
rect -12598 21370 -12586 27346
rect -12552 21370 -12540 27346
rect -12598 21358 -12540 21370
rect -12440 27346 -12382 27358
rect -12440 21370 -12428 27346
rect -12394 21370 -12382 27346
rect -12440 21358 -12382 21370
rect -12282 27346 -12224 27358
rect -12282 21370 -12270 27346
rect -12236 21370 -12224 27346
rect -12282 21358 -12224 21370
rect -12124 27346 -12066 27358
rect -12124 21370 -12112 27346
rect -12078 21370 -12066 27346
rect -12124 21358 -12066 21370
rect -11966 27346 -11908 27358
rect -11966 21370 -11954 27346
rect -11920 21370 -11908 27346
rect -11966 21358 -11908 21370
rect -11808 27346 -11750 27358
rect -11808 21370 -11796 27346
rect -11762 21370 -11750 27346
rect -11808 21358 -11750 21370
rect -11650 27346 -11592 27358
rect -11650 21370 -11638 27346
rect -11604 21370 -11592 27346
rect -11650 21358 -11592 21370
rect -11492 27346 -11434 27358
rect -11492 21370 -11480 27346
rect -11446 21370 -11434 27346
rect -11492 21358 -11434 21370
rect -11334 27346 -11276 27358
rect -11334 21370 -11322 27346
rect -11288 21370 -11276 27346
rect -11334 21358 -11276 21370
rect -11176 27346 -11118 27358
rect -11176 21370 -11164 27346
rect -11130 21370 -11118 27346
rect -11176 21358 -11118 21370
rect -11018 27346 -10960 27358
rect -11018 21370 -11006 27346
rect -10972 21370 -10960 27346
rect -11018 21358 -10960 21370
rect -10860 27346 -10802 27358
rect -10860 21370 -10848 27346
rect -10814 21370 -10802 27346
rect -10860 21358 -10802 21370
rect -10702 27346 -10644 27358
rect -10702 21370 -10690 27346
rect -10656 21370 -10644 27346
rect -10702 21358 -10644 21370
rect -10544 27346 -10486 27358
rect -10544 21370 -10532 27346
rect -10498 21370 -10486 27346
rect -10544 21358 -10486 21370
rect -10386 27346 -10328 27358
rect -10386 21370 -10374 27346
rect -10340 21370 -10328 27346
rect -10386 21358 -10328 21370
rect -10228 27346 -10170 27358
rect -10228 21370 -10216 27346
rect -10182 21370 -10170 27346
rect -10228 21358 -10170 21370
rect -10070 27346 -10012 27358
rect -10070 21370 -10058 27346
rect -10024 21370 -10012 27346
rect -10070 21358 -10012 21370
rect -9912 27346 -9854 27358
rect -9912 21370 -9900 27346
rect -9866 21370 -9854 27346
rect -9912 21358 -9854 21370
rect -9754 27346 -9696 27358
rect -9754 21370 -9742 27346
rect -9708 21370 -9696 27346
rect -9754 21358 -9696 21370
rect -9596 27346 -9538 27358
rect -9596 21370 -9584 27346
rect -9550 21370 -9538 27346
rect -9596 21358 -9538 21370
rect -9438 27346 -9380 27358
rect -9438 21370 -9426 27346
rect -9392 21370 -9380 27346
rect -9438 21358 -9380 21370
rect -9280 27346 -9222 27358
rect -9280 21370 -9268 27346
rect -9234 21370 -9222 27346
rect -9280 21358 -9222 21370
rect -9122 27346 -9064 27358
rect -9122 21370 -9110 27346
rect -9076 21370 -9064 27346
rect -9122 21358 -9064 21370
rect -8964 27346 -8906 27358
rect -8964 21370 -8952 27346
rect -8918 21370 -8906 27346
rect -8964 21358 -8906 21370
rect -8806 27346 -8748 27358
rect -8806 21370 -8794 27346
rect -8760 21370 -8748 27346
rect -8806 21358 -8748 21370
rect -8648 27346 -8590 27358
rect -8648 21370 -8636 27346
rect -8602 21370 -8590 27346
rect -8648 21358 -8590 21370
rect -8490 27346 -8432 27358
rect -8490 21370 -8478 27346
rect -8444 21370 -8432 27346
rect -8490 21358 -8432 21370
rect -6930 27346 -6872 27358
rect -6930 21370 -6918 27346
rect -6884 21370 -6872 27346
rect -6930 21358 -6872 21370
rect -6772 27346 -6714 27358
rect -6772 21370 -6760 27346
rect -6726 21370 -6714 27346
rect -6772 21358 -6714 21370
rect -6614 27346 -6556 27358
rect -6614 21370 -6602 27346
rect -6568 21370 -6556 27346
rect -6614 21358 -6556 21370
rect -6456 27346 -6398 27358
rect -6456 21370 -6444 27346
rect -6410 21370 -6398 27346
rect -6456 21358 -6398 21370
rect -6298 27346 -6240 27358
rect -6298 21370 -6286 27346
rect -6252 21370 -6240 27346
rect -6298 21358 -6240 21370
rect -6140 27346 -6082 27358
rect -6140 21370 -6128 27346
rect -6094 21370 -6082 27346
rect -6140 21358 -6082 21370
rect -5982 27346 -5924 27358
rect -5982 21370 -5970 27346
rect -5936 21370 -5924 27346
rect -5982 21358 -5924 21370
rect -5824 27346 -5766 27358
rect -5824 21370 -5812 27346
rect -5778 21370 -5766 27346
rect -5824 21358 -5766 21370
rect -5666 27346 -5608 27358
rect -5666 21370 -5654 27346
rect -5620 21370 -5608 27346
rect -5666 21358 -5608 21370
rect -5508 27346 -5450 27358
rect -5508 21370 -5496 27346
rect -5462 21370 -5450 27346
rect -5508 21358 -5450 21370
rect -5350 27346 -5292 27358
rect -5350 21370 -5338 27346
rect -5304 21370 -5292 27346
rect -5350 21358 -5292 21370
rect -5192 27346 -5134 27358
rect -5192 21370 -5180 27346
rect -5146 21370 -5134 27346
rect -5192 21358 -5134 21370
rect -5034 27346 -4976 27358
rect -5034 21370 -5022 27346
rect -4988 21370 -4976 27346
rect -5034 21358 -4976 21370
rect -4876 27346 -4818 27358
rect -4876 21370 -4864 27346
rect -4830 21370 -4818 27346
rect -4876 21358 -4818 21370
rect -4718 27346 -4660 27358
rect -4718 21370 -4706 27346
rect -4672 21370 -4660 27346
rect -4718 21358 -4660 21370
rect -4560 27346 -4502 27358
rect -4560 21370 -4548 27346
rect -4514 21370 -4502 27346
rect -4560 21358 -4502 21370
rect -4402 27346 -4344 27358
rect -4402 21370 -4390 27346
rect -4356 21370 -4344 27346
rect -4402 21358 -4344 21370
rect -4244 27346 -4186 27358
rect -4244 21370 -4232 27346
rect -4198 21370 -4186 27346
rect -4244 21358 -4186 21370
rect -4086 27346 -4028 27358
rect -4086 21370 -4074 27346
rect -4040 21370 -4028 27346
rect -4086 21358 -4028 21370
rect -3928 27346 -3870 27358
rect -3928 21370 -3916 27346
rect -3882 21370 -3870 27346
rect -3928 21358 -3870 21370
rect -3770 27346 -3712 27358
rect -3770 21370 -3758 27346
rect -3724 21370 -3712 27346
rect -3770 21358 -3712 21370
rect -3612 27346 -3554 27358
rect -3612 21370 -3600 27346
rect -3566 21370 -3554 27346
rect -3612 21358 -3554 21370
rect -3454 27346 -3396 27358
rect -3454 21370 -3442 27346
rect -3408 21370 -3396 27346
rect -3454 21358 -3396 21370
rect -3296 27346 -3238 27358
rect -3296 21370 -3284 27346
rect -3250 21370 -3238 27346
rect -3296 21358 -3238 21370
rect -3138 27346 -3080 27358
rect -3138 21370 -3126 27346
rect -3092 21370 -3080 27346
rect -3138 21358 -3080 21370
rect -2980 27346 -2922 27358
rect -2980 21370 -2968 27346
rect -2934 21370 -2922 27346
rect -2980 21358 -2922 21370
rect -2822 27346 -2764 27358
rect -2822 21370 -2810 27346
rect -2776 21370 -2764 27346
rect -2822 21358 -2764 21370
rect -2664 27346 -2606 27358
rect -2664 21370 -2652 27346
rect -2618 21370 -2606 27346
rect -2664 21358 -2606 21370
rect -2506 27346 -2448 27358
rect -2506 21370 -2494 27346
rect -2460 21370 -2448 27346
rect -2506 21358 -2448 21370
rect -2348 27346 -2290 27358
rect -2348 21370 -2336 27346
rect -2302 21370 -2290 27346
rect -2348 21358 -2290 21370
rect -2190 27346 -2132 27358
rect -2190 21370 -2178 27346
rect -2144 21370 -2132 27346
rect -2190 21358 -2132 21370
rect -630 27346 -572 27358
rect -630 21370 -618 27346
rect -584 21370 -572 27346
rect -630 21358 -572 21370
rect -472 27346 -414 27358
rect -472 21370 -460 27346
rect -426 21370 -414 27346
rect -472 21358 -414 21370
rect -314 27346 -256 27358
rect -314 21370 -302 27346
rect -268 21370 -256 27346
rect -314 21358 -256 21370
rect -156 27346 -98 27358
rect -156 21370 -144 27346
rect -110 21370 -98 27346
rect -156 21358 -98 21370
rect 2 27346 60 27358
rect 2 21370 14 27346
rect 48 21370 60 27346
rect 2 21358 60 21370
rect 160 27346 218 27358
rect 160 21370 172 27346
rect 206 21370 218 27346
rect 160 21358 218 21370
rect 318 27346 376 27358
rect 318 21370 330 27346
rect 364 21370 376 27346
rect 318 21358 376 21370
rect 476 27346 534 27358
rect 476 21370 488 27346
rect 522 21370 534 27346
rect 476 21358 534 21370
rect 634 27346 692 27358
rect 634 21370 646 27346
rect 680 21370 692 27346
rect 634 21358 692 21370
rect 792 27346 850 27358
rect 792 21370 804 27346
rect 838 21370 850 27346
rect 792 21358 850 21370
rect 950 27346 1008 27358
rect 950 21370 962 27346
rect 996 21370 1008 27346
rect 950 21358 1008 21370
rect 1108 27346 1166 27358
rect 1108 21370 1120 27346
rect 1154 21370 1166 27346
rect 1108 21358 1166 21370
rect 1266 27346 1324 27358
rect 1266 21370 1278 27346
rect 1312 21370 1324 27346
rect 1266 21358 1324 21370
rect 1424 27346 1482 27358
rect 1424 21370 1436 27346
rect 1470 21370 1482 27346
rect 1424 21358 1482 21370
rect 1582 27346 1640 27358
rect 1582 21370 1594 27346
rect 1628 21370 1640 27346
rect 1582 21358 1640 21370
rect 1740 27346 1798 27358
rect 1740 21370 1752 27346
rect 1786 21370 1798 27346
rect 1740 21358 1798 21370
rect 1898 27346 1956 27358
rect 1898 21370 1910 27346
rect 1944 21370 1956 27346
rect 1898 21358 1956 21370
rect 2056 27346 2114 27358
rect 2056 21370 2068 27346
rect 2102 21370 2114 27346
rect 2056 21358 2114 21370
rect 2214 27346 2272 27358
rect 2214 21370 2226 27346
rect 2260 21370 2272 27346
rect 2214 21358 2272 21370
rect 2372 27346 2430 27358
rect 2372 21370 2384 27346
rect 2418 21370 2430 27346
rect 2372 21358 2430 21370
rect 2530 27346 2588 27358
rect 2530 21370 2542 27346
rect 2576 21370 2588 27346
rect 2530 21358 2588 21370
rect 2688 27346 2746 27358
rect 2688 21370 2700 27346
rect 2734 21370 2746 27346
rect 2688 21358 2746 21370
rect 2846 27346 2904 27358
rect 2846 21370 2858 27346
rect 2892 21370 2904 27346
rect 2846 21358 2904 21370
rect 3004 27346 3062 27358
rect 3004 21370 3016 27346
rect 3050 21370 3062 27346
rect 3004 21358 3062 21370
rect 3162 27346 3220 27358
rect 3162 21370 3174 27346
rect 3208 21370 3220 27346
rect 3162 21358 3220 21370
rect 3320 27346 3378 27358
rect 3320 21370 3332 27346
rect 3366 21370 3378 27346
rect 3320 21358 3378 21370
rect 3478 27346 3536 27358
rect 3478 21370 3490 27346
rect 3524 21370 3536 27346
rect 3478 21358 3536 21370
rect 3636 27346 3694 27358
rect 3636 21370 3648 27346
rect 3682 21370 3694 27346
rect 3636 21358 3694 21370
rect 3794 27346 3852 27358
rect 3794 21370 3806 27346
rect 3840 21370 3852 27346
rect 3794 21358 3852 21370
rect 3952 27346 4010 27358
rect 3952 21370 3964 27346
rect 3998 21370 4010 27346
rect 3952 21358 4010 21370
rect 4110 27346 4168 27358
rect 4110 21370 4122 27346
rect 4156 21370 4168 27346
rect 4110 21358 4168 21370
rect 5670 27346 5728 27358
rect 5670 21370 5682 27346
rect 5716 21370 5728 27346
rect 5670 21358 5728 21370
rect 5828 27346 5886 27358
rect 5828 21370 5840 27346
rect 5874 21370 5886 27346
rect 5828 21358 5886 21370
rect 5986 27346 6044 27358
rect 5986 21370 5998 27346
rect 6032 21370 6044 27346
rect 5986 21358 6044 21370
rect 6144 27346 6202 27358
rect 6144 21370 6156 27346
rect 6190 21370 6202 27346
rect 6144 21358 6202 21370
rect 6302 27346 6360 27358
rect 6302 21370 6314 27346
rect 6348 21370 6360 27346
rect 6302 21358 6360 21370
rect 6460 27346 6518 27358
rect 6460 21370 6472 27346
rect 6506 21370 6518 27346
rect 6460 21358 6518 21370
rect 6618 27346 6676 27358
rect 6618 21370 6630 27346
rect 6664 21370 6676 27346
rect 6618 21358 6676 21370
rect 6776 27346 6834 27358
rect 6776 21370 6788 27346
rect 6822 21370 6834 27346
rect 6776 21358 6834 21370
rect 6934 27346 6992 27358
rect 6934 21370 6946 27346
rect 6980 21370 6992 27346
rect 6934 21358 6992 21370
rect 7092 27346 7150 27358
rect 7092 21370 7104 27346
rect 7138 21370 7150 27346
rect 7092 21358 7150 21370
rect 7250 27346 7308 27358
rect 7250 21370 7262 27346
rect 7296 21370 7308 27346
rect 7250 21358 7308 21370
rect 7408 27346 7466 27358
rect 7408 21370 7420 27346
rect 7454 21370 7466 27346
rect 7408 21358 7466 21370
rect 7566 27346 7624 27358
rect 7566 21370 7578 27346
rect 7612 21370 7624 27346
rect 7566 21358 7624 21370
rect 7724 27346 7782 27358
rect 7724 21370 7736 27346
rect 7770 21370 7782 27346
rect 7724 21358 7782 21370
rect 7882 27346 7940 27358
rect 7882 21370 7894 27346
rect 7928 21370 7940 27346
rect 7882 21358 7940 21370
rect 8040 27346 8098 27358
rect 8040 21370 8052 27346
rect 8086 21370 8098 27346
rect 8040 21358 8098 21370
rect 8198 27346 8256 27358
rect 8198 21370 8210 27346
rect 8244 21370 8256 27346
rect 8198 21358 8256 21370
rect 8356 27346 8414 27358
rect 8356 21370 8368 27346
rect 8402 21370 8414 27346
rect 8356 21358 8414 21370
rect 8514 27346 8572 27358
rect 8514 21370 8526 27346
rect 8560 21370 8572 27346
rect 8514 21358 8572 21370
rect 8672 27346 8730 27358
rect 8672 21370 8684 27346
rect 8718 21370 8730 27346
rect 8672 21358 8730 21370
rect 8830 27346 8888 27358
rect 8830 21370 8842 27346
rect 8876 21370 8888 27346
rect 8830 21358 8888 21370
rect 8988 27346 9046 27358
rect 8988 21370 9000 27346
rect 9034 21370 9046 27346
rect 8988 21358 9046 21370
rect 9146 27346 9204 27358
rect 9146 21370 9158 27346
rect 9192 21370 9204 27346
rect 9146 21358 9204 21370
rect 9304 27346 9362 27358
rect 9304 21370 9316 27346
rect 9350 21370 9362 27346
rect 9304 21358 9362 21370
rect 9462 27346 9520 27358
rect 9462 21370 9474 27346
rect 9508 21370 9520 27346
rect 9462 21358 9520 21370
rect 9620 27346 9678 27358
rect 9620 21370 9632 27346
rect 9666 21370 9678 27346
rect 9620 21358 9678 21370
rect 9778 27346 9836 27358
rect 9778 21370 9790 27346
rect 9824 21370 9836 27346
rect 9778 21358 9836 21370
rect 9936 27346 9994 27358
rect 9936 21370 9948 27346
rect 9982 21370 9994 27346
rect 9936 21358 9994 21370
rect 10094 27346 10152 27358
rect 10094 21370 10106 27346
rect 10140 21370 10152 27346
rect 10094 21358 10152 21370
rect 10252 27346 10310 27358
rect 10252 21370 10264 27346
rect 10298 21370 10310 27346
rect 10252 21358 10310 21370
rect 10410 27346 10468 27358
rect 10410 21370 10422 27346
rect 10456 21370 10468 27346
rect 10410 21358 10468 21370
rect -13230 19046 -13172 19058
rect -13230 13070 -13218 19046
rect -13184 13070 -13172 19046
rect -13230 13058 -13172 13070
rect -13072 19046 -13014 19058
rect -13072 13070 -13060 19046
rect -13026 13070 -13014 19046
rect -13072 13058 -13014 13070
rect -12914 19046 -12856 19058
rect -12914 13070 -12902 19046
rect -12868 13070 -12856 19046
rect -12914 13058 -12856 13070
rect -12756 19046 -12698 19058
rect -12756 13070 -12744 19046
rect -12710 13070 -12698 19046
rect -12756 13058 -12698 13070
rect -12598 19046 -12540 19058
rect -12598 13070 -12586 19046
rect -12552 13070 -12540 19046
rect -12598 13058 -12540 13070
rect -12440 19046 -12382 19058
rect -12440 13070 -12428 19046
rect -12394 13070 -12382 19046
rect -12440 13058 -12382 13070
rect -12282 19046 -12224 19058
rect -12282 13070 -12270 19046
rect -12236 13070 -12224 19046
rect -12282 13058 -12224 13070
rect -12124 19046 -12066 19058
rect -12124 13070 -12112 19046
rect -12078 13070 -12066 19046
rect -12124 13058 -12066 13070
rect -11966 19046 -11908 19058
rect -11966 13070 -11954 19046
rect -11920 13070 -11908 19046
rect -11966 13058 -11908 13070
rect -11808 19046 -11750 19058
rect -11808 13070 -11796 19046
rect -11762 13070 -11750 19046
rect -11808 13058 -11750 13070
rect -11650 19046 -11592 19058
rect -11650 13070 -11638 19046
rect -11604 13070 -11592 19046
rect -11650 13058 -11592 13070
rect -11492 19046 -11434 19058
rect -11492 13070 -11480 19046
rect -11446 13070 -11434 19046
rect -11492 13058 -11434 13070
rect -11334 19046 -11276 19058
rect -11334 13070 -11322 19046
rect -11288 13070 -11276 19046
rect -11334 13058 -11276 13070
rect -11176 19046 -11118 19058
rect -11176 13070 -11164 19046
rect -11130 13070 -11118 19046
rect -11176 13058 -11118 13070
rect -11018 19046 -10960 19058
rect -11018 13070 -11006 19046
rect -10972 13070 -10960 19046
rect -11018 13058 -10960 13070
rect -10860 19046 -10802 19058
rect -10860 13070 -10848 19046
rect -10814 13070 -10802 19046
rect -10860 13058 -10802 13070
rect -10702 19046 -10644 19058
rect -10702 13070 -10690 19046
rect -10656 13070 -10644 19046
rect -10702 13058 -10644 13070
rect -10544 19046 -10486 19058
rect -10544 13070 -10532 19046
rect -10498 13070 -10486 19046
rect -10544 13058 -10486 13070
rect -10386 19046 -10328 19058
rect -10386 13070 -10374 19046
rect -10340 13070 -10328 19046
rect -10386 13058 -10328 13070
rect -10228 19046 -10170 19058
rect -10228 13070 -10216 19046
rect -10182 13070 -10170 19046
rect -10228 13058 -10170 13070
rect -10070 19046 -10012 19058
rect -10070 13070 -10058 19046
rect -10024 13070 -10012 19046
rect -10070 13058 -10012 13070
rect -9912 19046 -9854 19058
rect -9912 13070 -9900 19046
rect -9866 13070 -9854 19046
rect -9912 13058 -9854 13070
rect -9754 19046 -9696 19058
rect -9754 13070 -9742 19046
rect -9708 13070 -9696 19046
rect -9754 13058 -9696 13070
rect -9596 19046 -9538 19058
rect -9596 13070 -9584 19046
rect -9550 13070 -9538 19046
rect -9596 13058 -9538 13070
rect -9438 19046 -9380 19058
rect -9438 13070 -9426 19046
rect -9392 13070 -9380 19046
rect -9438 13058 -9380 13070
rect -9280 19046 -9222 19058
rect -9280 13070 -9268 19046
rect -9234 13070 -9222 19046
rect -9280 13058 -9222 13070
rect -9122 19046 -9064 19058
rect -9122 13070 -9110 19046
rect -9076 13070 -9064 19046
rect -9122 13058 -9064 13070
rect -8964 19046 -8906 19058
rect -8964 13070 -8952 19046
rect -8918 13070 -8906 19046
rect -8964 13058 -8906 13070
rect -8806 19046 -8748 19058
rect -8806 13070 -8794 19046
rect -8760 13070 -8748 19046
rect -8806 13058 -8748 13070
rect -8648 19046 -8590 19058
rect -8648 13070 -8636 19046
rect -8602 13070 -8590 19046
rect -8648 13058 -8590 13070
rect -8490 19046 -8432 19058
rect -8490 13070 -8478 19046
rect -8444 13070 -8432 19046
rect -8490 13058 -8432 13070
rect -6930 19046 -6872 19058
rect -6930 13070 -6918 19046
rect -6884 13070 -6872 19046
rect -6930 13058 -6872 13070
rect -6772 19046 -6714 19058
rect -6772 13070 -6760 19046
rect -6726 13070 -6714 19046
rect -6772 13058 -6714 13070
rect -6614 19046 -6556 19058
rect -6614 13070 -6602 19046
rect -6568 13070 -6556 19046
rect -6614 13058 -6556 13070
rect -6456 19046 -6398 19058
rect -6456 13070 -6444 19046
rect -6410 13070 -6398 19046
rect -6456 13058 -6398 13070
rect -6298 19046 -6240 19058
rect -6298 13070 -6286 19046
rect -6252 13070 -6240 19046
rect -6298 13058 -6240 13070
rect -6140 19046 -6082 19058
rect -6140 13070 -6128 19046
rect -6094 13070 -6082 19046
rect -6140 13058 -6082 13070
rect -5982 19046 -5924 19058
rect -5982 13070 -5970 19046
rect -5936 13070 -5924 19046
rect -5982 13058 -5924 13070
rect -5824 19046 -5766 19058
rect -5824 13070 -5812 19046
rect -5778 13070 -5766 19046
rect -5824 13058 -5766 13070
rect -5666 19046 -5608 19058
rect -5666 13070 -5654 19046
rect -5620 13070 -5608 19046
rect -5666 13058 -5608 13070
rect -5508 19046 -5450 19058
rect -5508 13070 -5496 19046
rect -5462 13070 -5450 19046
rect -5508 13058 -5450 13070
rect -5350 19046 -5292 19058
rect -5350 13070 -5338 19046
rect -5304 13070 -5292 19046
rect -5350 13058 -5292 13070
rect -5192 19046 -5134 19058
rect -5192 13070 -5180 19046
rect -5146 13070 -5134 19046
rect -5192 13058 -5134 13070
rect -5034 19046 -4976 19058
rect -5034 13070 -5022 19046
rect -4988 13070 -4976 19046
rect -5034 13058 -4976 13070
rect -4876 19046 -4818 19058
rect -4876 13070 -4864 19046
rect -4830 13070 -4818 19046
rect -4876 13058 -4818 13070
rect -4718 19046 -4660 19058
rect -4718 13070 -4706 19046
rect -4672 13070 -4660 19046
rect -4718 13058 -4660 13070
rect -4560 19046 -4502 19058
rect -4560 13070 -4548 19046
rect -4514 13070 -4502 19046
rect -4560 13058 -4502 13070
rect -4402 19046 -4344 19058
rect -4402 13070 -4390 19046
rect -4356 13070 -4344 19046
rect -4402 13058 -4344 13070
rect -4244 19046 -4186 19058
rect -4244 13070 -4232 19046
rect -4198 13070 -4186 19046
rect -4244 13058 -4186 13070
rect -4086 19046 -4028 19058
rect -4086 13070 -4074 19046
rect -4040 13070 -4028 19046
rect -4086 13058 -4028 13070
rect -3928 19046 -3870 19058
rect -3928 13070 -3916 19046
rect -3882 13070 -3870 19046
rect -3928 13058 -3870 13070
rect -3770 19046 -3712 19058
rect -3770 13070 -3758 19046
rect -3724 13070 -3712 19046
rect -3770 13058 -3712 13070
rect -3612 19046 -3554 19058
rect -3612 13070 -3600 19046
rect -3566 13070 -3554 19046
rect -3612 13058 -3554 13070
rect -3454 19046 -3396 19058
rect -3454 13070 -3442 19046
rect -3408 13070 -3396 19046
rect -3454 13058 -3396 13070
rect -3296 19046 -3238 19058
rect -3296 13070 -3284 19046
rect -3250 13070 -3238 19046
rect -3296 13058 -3238 13070
rect -3138 19046 -3080 19058
rect -3138 13070 -3126 19046
rect -3092 13070 -3080 19046
rect -3138 13058 -3080 13070
rect -2980 19046 -2922 19058
rect -2980 13070 -2968 19046
rect -2934 13070 -2922 19046
rect -2980 13058 -2922 13070
rect -2822 19046 -2764 19058
rect -2822 13070 -2810 19046
rect -2776 13070 -2764 19046
rect -2822 13058 -2764 13070
rect -2664 19046 -2606 19058
rect -2664 13070 -2652 19046
rect -2618 13070 -2606 19046
rect -2664 13058 -2606 13070
rect -2506 19046 -2448 19058
rect -2506 13070 -2494 19046
rect -2460 13070 -2448 19046
rect -2506 13058 -2448 13070
rect -2348 19046 -2290 19058
rect -2348 13070 -2336 19046
rect -2302 13070 -2290 19046
rect -2348 13058 -2290 13070
rect -2190 19046 -2132 19058
rect -2190 13070 -2178 19046
rect -2144 13070 -2132 19046
rect -2190 13058 -2132 13070
rect -630 19046 -572 19058
rect -630 13070 -618 19046
rect -584 13070 -572 19046
rect -630 13058 -572 13070
rect -472 19046 -414 19058
rect -472 13070 -460 19046
rect -426 13070 -414 19046
rect -472 13058 -414 13070
rect -314 19046 -256 19058
rect -314 13070 -302 19046
rect -268 13070 -256 19046
rect -314 13058 -256 13070
rect -156 19046 -98 19058
rect -156 13070 -144 19046
rect -110 13070 -98 19046
rect -156 13058 -98 13070
rect 2 19046 60 19058
rect 2 13070 14 19046
rect 48 13070 60 19046
rect 2 13058 60 13070
rect 160 19046 218 19058
rect 160 13070 172 19046
rect 206 13070 218 19046
rect 160 13058 218 13070
rect 318 19046 376 19058
rect 318 13070 330 19046
rect 364 13070 376 19046
rect 318 13058 376 13070
rect 476 19046 534 19058
rect 476 13070 488 19046
rect 522 13070 534 19046
rect 476 13058 534 13070
rect 634 19046 692 19058
rect 634 13070 646 19046
rect 680 13070 692 19046
rect 634 13058 692 13070
rect 792 19046 850 19058
rect 792 13070 804 19046
rect 838 13070 850 19046
rect 792 13058 850 13070
rect 950 19046 1008 19058
rect 950 13070 962 19046
rect 996 13070 1008 19046
rect 950 13058 1008 13070
rect 1108 19046 1166 19058
rect 1108 13070 1120 19046
rect 1154 13070 1166 19046
rect 1108 13058 1166 13070
rect 1266 19046 1324 19058
rect 1266 13070 1278 19046
rect 1312 13070 1324 19046
rect 1266 13058 1324 13070
rect 1424 19046 1482 19058
rect 1424 13070 1436 19046
rect 1470 13070 1482 19046
rect 1424 13058 1482 13070
rect 1582 19046 1640 19058
rect 1582 13070 1594 19046
rect 1628 13070 1640 19046
rect 1582 13058 1640 13070
rect 1740 19046 1798 19058
rect 1740 13070 1752 19046
rect 1786 13070 1798 19046
rect 1740 13058 1798 13070
rect 1898 19046 1956 19058
rect 1898 13070 1910 19046
rect 1944 13070 1956 19046
rect 1898 13058 1956 13070
rect 2056 19046 2114 19058
rect 2056 13070 2068 19046
rect 2102 13070 2114 19046
rect 2056 13058 2114 13070
rect 2214 19046 2272 19058
rect 2214 13070 2226 19046
rect 2260 13070 2272 19046
rect 2214 13058 2272 13070
rect 2372 19046 2430 19058
rect 2372 13070 2384 19046
rect 2418 13070 2430 19046
rect 2372 13058 2430 13070
rect 2530 19046 2588 19058
rect 2530 13070 2542 19046
rect 2576 13070 2588 19046
rect 2530 13058 2588 13070
rect 2688 19046 2746 19058
rect 2688 13070 2700 19046
rect 2734 13070 2746 19046
rect 2688 13058 2746 13070
rect 2846 19046 2904 19058
rect 2846 13070 2858 19046
rect 2892 13070 2904 19046
rect 2846 13058 2904 13070
rect 3004 19046 3062 19058
rect 3004 13070 3016 19046
rect 3050 13070 3062 19046
rect 3004 13058 3062 13070
rect 3162 19046 3220 19058
rect 3162 13070 3174 19046
rect 3208 13070 3220 19046
rect 3162 13058 3220 13070
rect 3320 19046 3378 19058
rect 3320 13070 3332 19046
rect 3366 13070 3378 19046
rect 3320 13058 3378 13070
rect 3478 19046 3536 19058
rect 3478 13070 3490 19046
rect 3524 13070 3536 19046
rect 3478 13058 3536 13070
rect 3636 19046 3694 19058
rect 3636 13070 3648 19046
rect 3682 13070 3694 19046
rect 3636 13058 3694 13070
rect 3794 19046 3852 19058
rect 3794 13070 3806 19046
rect 3840 13070 3852 19046
rect 3794 13058 3852 13070
rect 3952 19046 4010 19058
rect 3952 13070 3964 19046
rect 3998 13070 4010 19046
rect 3952 13058 4010 13070
rect 4110 19046 4168 19058
rect 4110 13070 4122 19046
rect 4156 13070 4168 19046
rect 4110 13058 4168 13070
rect 5670 19046 5728 19058
rect 5670 13070 5682 19046
rect 5716 13070 5728 19046
rect 5670 13058 5728 13070
rect 5828 19046 5886 19058
rect 5828 13070 5840 19046
rect 5874 13070 5886 19046
rect 5828 13058 5886 13070
rect 5986 19046 6044 19058
rect 5986 13070 5998 19046
rect 6032 13070 6044 19046
rect 5986 13058 6044 13070
rect 6144 19046 6202 19058
rect 6144 13070 6156 19046
rect 6190 13070 6202 19046
rect 6144 13058 6202 13070
rect 6302 19046 6360 19058
rect 6302 13070 6314 19046
rect 6348 13070 6360 19046
rect 6302 13058 6360 13070
rect 6460 19046 6518 19058
rect 6460 13070 6472 19046
rect 6506 13070 6518 19046
rect 6460 13058 6518 13070
rect 6618 19046 6676 19058
rect 6618 13070 6630 19046
rect 6664 13070 6676 19046
rect 6618 13058 6676 13070
rect 6776 19046 6834 19058
rect 6776 13070 6788 19046
rect 6822 13070 6834 19046
rect 6776 13058 6834 13070
rect 6934 19046 6992 19058
rect 6934 13070 6946 19046
rect 6980 13070 6992 19046
rect 6934 13058 6992 13070
rect 7092 19046 7150 19058
rect 7092 13070 7104 19046
rect 7138 13070 7150 19046
rect 7092 13058 7150 13070
rect 7250 19046 7308 19058
rect 7250 13070 7262 19046
rect 7296 13070 7308 19046
rect 7250 13058 7308 13070
rect 7408 19046 7466 19058
rect 7408 13070 7420 19046
rect 7454 13070 7466 19046
rect 7408 13058 7466 13070
rect 7566 19046 7624 19058
rect 7566 13070 7578 19046
rect 7612 13070 7624 19046
rect 7566 13058 7624 13070
rect 7724 19046 7782 19058
rect 7724 13070 7736 19046
rect 7770 13070 7782 19046
rect 7724 13058 7782 13070
rect 7882 19046 7940 19058
rect 7882 13070 7894 19046
rect 7928 13070 7940 19046
rect 7882 13058 7940 13070
rect 8040 19046 8098 19058
rect 8040 13070 8052 19046
rect 8086 13070 8098 19046
rect 8040 13058 8098 13070
rect 8198 19046 8256 19058
rect 8198 13070 8210 19046
rect 8244 13070 8256 19046
rect 8198 13058 8256 13070
rect 8356 19046 8414 19058
rect 8356 13070 8368 19046
rect 8402 13070 8414 19046
rect 8356 13058 8414 13070
rect 8514 19046 8572 19058
rect 8514 13070 8526 19046
rect 8560 13070 8572 19046
rect 8514 13058 8572 13070
rect 8672 19046 8730 19058
rect 8672 13070 8684 19046
rect 8718 13070 8730 19046
rect 8672 13058 8730 13070
rect 8830 19046 8888 19058
rect 8830 13070 8842 19046
rect 8876 13070 8888 19046
rect 8830 13058 8888 13070
rect 8988 19046 9046 19058
rect 8988 13070 9000 19046
rect 9034 13070 9046 19046
rect 8988 13058 9046 13070
rect 9146 19046 9204 19058
rect 9146 13070 9158 19046
rect 9192 13070 9204 19046
rect 9146 13058 9204 13070
rect 9304 19046 9362 19058
rect 9304 13070 9316 19046
rect 9350 13070 9362 19046
rect 9304 13058 9362 13070
rect 9462 19046 9520 19058
rect 9462 13070 9474 19046
rect 9508 13070 9520 19046
rect 9462 13058 9520 13070
rect 9620 19046 9678 19058
rect 9620 13070 9632 19046
rect 9666 13070 9678 19046
rect 9620 13058 9678 13070
rect 9778 19046 9836 19058
rect 9778 13070 9790 19046
rect 9824 13070 9836 19046
rect 9778 13058 9836 13070
rect 9936 19046 9994 19058
rect 9936 13070 9948 19046
rect 9982 13070 9994 19046
rect 9936 13058 9994 13070
rect 10094 19046 10152 19058
rect 10094 13070 10106 19046
rect 10140 13070 10152 19046
rect 10094 13058 10152 13070
rect 10252 19046 10310 19058
rect 10252 13070 10264 19046
rect 10298 13070 10310 19046
rect 10252 13058 10310 13070
rect 10410 19046 10468 19058
rect 10410 13070 10422 19046
rect 10456 13070 10468 19046
rect 10410 13058 10468 13070
rect -13230 12046 -13172 12058
rect -13230 6070 -13218 12046
rect -13184 6070 -13172 12046
rect -13230 6058 -13172 6070
rect -13072 12046 -13014 12058
rect -13072 6070 -13060 12046
rect -13026 6070 -13014 12046
rect -13072 6058 -13014 6070
rect -12914 12046 -12856 12058
rect -12914 6070 -12902 12046
rect -12868 6070 -12856 12046
rect -12914 6058 -12856 6070
rect -12756 12046 -12698 12058
rect -12756 6070 -12744 12046
rect -12710 6070 -12698 12046
rect -12756 6058 -12698 6070
rect -12598 12046 -12540 12058
rect -12598 6070 -12586 12046
rect -12552 6070 -12540 12046
rect -12598 6058 -12540 6070
rect -12440 12046 -12382 12058
rect -12440 6070 -12428 12046
rect -12394 6070 -12382 12046
rect -12440 6058 -12382 6070
rect -12282 12046 -12224 12058
rect -12282 6070 -12270 12046
rect -12236 6070 -12224 12046
rect -12282 6058 -12224 6070
rect -12124 12046 -12066 12058
rect -12124 6070 -12112 12046
rect -12078 6070 -12066 12046
rect -12124 6058 -12066 6070
rect -11966 12046 -11908 12058
rect -11966 6070 -11954 12046
rect -11920 6070 -11908 12046
rect -11966 6058 -11908 6070
rect -11808 12046 -11750 12058
rect -11808 6070 -11796 12046
rect -11762 6070 -11750 12046
rect -11808 6058 -11750 6070
rect -11650 12046 -11592 12058
rect -11650 6070 -11638 12046
rect -11604 6070 -11592 12046
rect -11650 6058 -11592 6070
rect -11492 12046 -11434 12058
rect -11492 6070 -11480 12046
rect -11446 6070 -11434 12046
rect -11492 6058 -11434 6070
rect -11334 12046 -11276 12058
rect -11334 6070 -11322 12046
rect -11288 6070 -11276 12046
rect -11334 6058 -11276 6070
rect -11176 12046 -11118 12058
rect -11176 6070 -11164 12046
rect -11130 6070 -11118 12046
rect -11176 6058 -11118 6070
rect -11018 12046 -10960 12058
rect -11018 6070 -11006 12046
rect -10972 6070 -10960 12046
rect -11018 6058 -10960 6070
rect -10860 12046 -10802 12058
rect -10860 6070 -10848 12046
rect -10814 6070 -10802 12046
rect -10860 6058 -10802 6070
rect -10702 12046 -10644 12058
rect -10702 6070 -10690 12046
rect -10656 6070 -10644 12046
rect -10702 6058 -10644 6070
rect -10544 12046 -10486 12058
rect -10544 6070 -10532 12046
rect -10498 6070 -10486 12046
rect -10544 6058 -10486 6070
rect -10386 12046 -10328 12058
rect -10386 6070 -10374 12046
rect -10340 6070 -10328 12046
rect -10386 6058 -10328 6070
rect -10228 12046 -10170 12058
rect -10228 6070 -10216 12046
rect -10182 6070 -10170 12046
rect -10228 6058 -10170 6070
rect -10070 12046 -10012 12058
rect -10070 6070 -10058 12046
rect -10024 6070 -10012 12046
rect -10070 6058 -10012 6070
rect -9912 12046 -9854 12058
rect -9912 6070 -9900 12046
rect -9866 6070 -9854 12046
rect -9912 6058 -9854 6070
rect -9754 12046 -9696 12058
rect -9754 6070 -9742 12046
rect -9708 6070 -9696 12046
rect -9754 6058 -9696 6070
rect -9596 12046 -9538 12058
rect -9596 6070 -9584 12046
rect -9550 6070 -9538 12046
rect -9596 6058 -9538 6070
rect -9438 12046 -9380 12058
rect -9438 6070 -9426 12046
rect -9392 6070 -9380 12046
rect -9438 6058 -9380 6070
rect -9280 12046 -9222 12058
rect -9280 6070 -9268 12046
rect -9234 6070 -9222 12046
rect -9280 6058 -9222 6070
rect -9122 12046 -9064 12058
rect -9122 6070 -9110 12046
rect -9076 6070 -9064 12046
rect -9122 6058 -9064 6070
rect -8964 12046 -8906 12058
rect -8964 6070 -8952 12046
rect -8918 6070 -8906 12046
rect -8964 6058 -8906 6070
rect -8806 12046 -8748 12058
rect -8806 6070 -8794 12046
rect -8760 6070 -8748 12046
rect -8806 6058 -8748 6070
rect -8648 12046 -8590 12058
rect -8648 6070 -8636 12046
rect -8602 6070 -8590 12046
rect -8648 6058 -8590 6070
rect -8490 12046 -8432 12058
rect -8490 6070 -8478 12046
rect -8444 6070 -8432 12046
rect -8490 6058 -8432 6070
rect -6930 12046 -6872 12058
rect -6930 6070 -6918 12046
rect -6884 6070 -6872 12046
rect -6930 6058 -6872 6070
rect -6772 12046 -6714 12058
rect -6772 6070 -6760 12046
rect -6726 6070 -6714 12046
rect -6772 6058 -6714 6070
rect -6614 12046 -6556 12058
rect -6614 6070 -6602 12046
rect -6568 6070 -6556 12046
rect -6614 6058 -6556 6070
rect -6456 12046 -6398 12058
rect -6456 6070 -6444 12046
rect -6410 6070 -6398 12046
rect -6456 6058 -6398 6070
rect -6298 12046 -6240 12058
rect -6298 6070 -6286 12046
rect -6252 6070 -6240 12046
rect -6298 6058 -6240 6070
rect -6140 12046 -6082 12058
rect -6140 6070 -6128 12046
rect -6094 6070 -6082 12046
rect -6140 6058 -6082 6070
rect -5982 12046 -5924 12058
rect -5982 6070 -5970 12046
rect -5936 6070 -5924 12046
rect -5982 6058 -5924 6070
rect -5824 12046 -5766 12058
rect -5824 6070 -5812 12046
rect -5778 6070 -5766 12046
rect -5824 6058 -5766 6070
rect -5666 12046 -5608 12058
rect -5666 6070 -5654 12046
rect -5620 6070 -5608 12046
rect -5666 6058 -5608 6070
rect -5508 12046 -5450 12058
rect -5508 6070 -5496 12046
rect -5462 6070 -5450 12046
rect -5508 6058 -5450 6070
rect -5350 12046 -5292 12058
rect -5350 6070 -5338 12046
rect -5304 6070 -5292 12046
rect -5350 6058 -5292 6070
rect -5192 12046 -5134 12058
rect -5192 6070 -5180 12046
rect -5146 6070 -5134 12046
rect -5192 6058 -5134 6070
rect -5034 12046 -4976 12058
rect -5034 6070 -5022 12046
rect -4988 6070 -4976 12046
rect -5034 6058 -4976 6070
rect -4876 12046 -4818 12058
rect -4876 6070 -4864 12046
rect -4830 6070 -4818 12046
rect -4876 6058 -4818 6070
rect -4718 12046 -4660 12058
rect -4718 6070 -4706 12046
rect -4672 6070 -4660 12046
rect -4718 6058 -4660 6070
rect -4560 12046 -4502 12058
rect -4560 6070 -4548 12046
rect -4514 6070 -4502 12046
rect -4560 6058 -4502 6070
rect -4402 12046 -4344 12058
rect -4402 6070 -4390 12046
rect -4356 6070 -4344 12046
rect -4402 6058 -4344 6070
rect -4244 12046 -4186 12058
rect -4244 6070 -4232 12046
rect -4198 6070 -4186 12046
rect -4244 6058 -4186 6070
rect -4086 12046 -4028 12058
rect -4086 6070 -4074 12046
rect -4040 6070 -4028 12046
rect -4086 6058 -4028 6070
rect -3928 12046 -3870 12058
rect -3928 6070 -3916 12046
rect -3882 6070 -3870 12046
rect -3928 6058 -3870 6070
rect -3770 12046 -3712 12058
rect -3770 6070 -3758 12046
rect -3724 6070 -3712 12046
rect -3770 6058 -3712 6070
rect -3612 12046 -3554 12058
rect -3612 6070 -3600 12046
rect -3566 6070 -3554 12046
rect -3612 6058 -3554 6070
rect -3454 12046 -3396 12058
rect -3454 6070 -3442 12046
rect -3408 6070 -3396 12046
rect -3454 6058 -3396 6070
rect -3296 12046 -3238 12058
rect -3296 6070 -3284 12046
rect -3250 6070 -3238 12046
rect -3296 6058 -3238 6070
rect -3138 12046 -3080 12058
rect -3138 6070 -3126 12046
rect -3092 6070 -3080 12046
rect -3138 6058 -3080 6070
rect -2980 12046 -2922 12058
rect -2980 6070 -2968 12046
rect -2934 6070 -2922 12046
rect -2980 6058 -2922 6070
rect -2822 12046 -2764 12058
rect -2822 6070 -2810 12046
rect -2776 6070 -2764 12046
rect -2822 6058 -2764 6070
rect -2664 12046 -2606 12058
rect -2664 6070 -2652 12046
rect -2618 6070 -2606 12046
rect -2664 6058 -2606 6070
rect -2506 12046 -2448 12058
rect -2506 6070 -2494 12046
rect -2460 6070 -2448 12046
rect -2506 6058 -2448 6070
rect -2348 12046 -2290 12058
rect -2348 6070 -2336 12046
rect -2302 6070 -2290 12046
rect -2348 6058 -2290 6070
rect -2190 12046 -2132 12058
rect -2190 6070 -2178 12046
rect -2144 6070 -2132 12046
rect -2190 6058 -2132 6070
rect -630 12046 -572 12058
rect -630 6070 -618 12046
rect -584 6070 -572 12046
rect -630 6058 -572 6070
rect -472 12046 -414 12058
rect -472 6070 -460 12046
rect -426 6070 -414 12046
rect -472 6058 -414 6070
rect -314 12046 -256 12058
rect -314 6070 -302 12046
rect -268 6070 -256 12046
rect -314 6058 -256 6070
rect -156 12046 -98 12058
rect -156 6070 -144 12046
rect -110 6070 -98 12046
rect -156 6058 -98 6070
rect 2 12046 60 12058
rect 2 6070 14 12046
rect 48 6070 60 12046
rect 2 6058 60 6070
rect 160 12046 218 12058
rect 160 6070 172 12046
rect 206 6070 218 12046
rect 160 6058 218 6070
rect 318 12046 376 12058
rect 318 6070 330 12046
rect 364 6070 376 12046
rect 318 6058 376 6070
rect 476 12046 534 12058
rect 476 6070 488 12046
rect 522 6070 534 12046
rect 476 6058 534 6070
rect 634 12046 692 12058
rect 634 6070 646 12046
rect 680 6070 692 12046
rect 634 6058 692 6070
rect 792 12046 850 12058
rect 792 6070 804 12046
rect 838 6070 850 12046
rect 792 6058 850 6070
rect 950 12046 1008 12058
rect 950 6070 962 12046
rect 996 6070 1008 12046
rect 950 6058 1008 6070
rect 1108 12046 1166 12058
rect 1108 6070 1120 12046
rect 1154 6070 1166 12046
rect 1108 6058 1166 6070
rect 1266 12046 1324 12058
rect 1266 6070 1278 12046
rect 1312 6070 1324 12046
rect 1266 6058 1324 6070
rect 1424 12046 1482 12058
rect 1424 6070 1436 12046
rect 1470 6070 1482 12046
rect 1424 6058 1482 6070
rect 1582 12046 1640 12058
rect 1582 6070 1594 12046
rect 1628 6070 1640 12046
rect 1582 6058 1640 6070
rect 1740 12046 1798 12058
rect 1740 6070 1752 12046
rect 1786 6070 1798 12046
rect 1740 6058 1798 6070
rect 1898 12046 1956 12058
rect 1898 6070 1910 12046
rect 1944 6070 1956 12046
rect 1898 6058 1956 6070
rect 2056 12046 2114 12058
rect 2056 6070 2068 12046
rect 2102 6070 2114 12046
rect 2056 6058 2114 6070
rect 2214 12046 2272 12058
rect 2214 6070 2226 12046
rect 2260 6070 2272 12046
rect 2214 6058 2272 6070
rect 2372 12046 2430 12058
rect 2372 6070 2384 12046
rect 2418 6070 2430 12046
rect 2372 6058 2430 6070
rect 2530 12046 2588 12058
rect 2530 6070 2542 12046
rect 2576 6070 2588 12046
rect 2530 6058 2588 6070
rect 2688 12046 2746 12058
rect 2688 6070 2700 12046
rect 2734 6070 2746 12046
rect 2688 6058 2746 6070
rect 2846 12046 2904 12058
rect 2846 6070 2858 12046
rect 2892 6070 2904 12046
rect 2846 6058 2904 6070
rect 3004 12046 3062 12058
rect 3004 6070 3016 12046
rect 3050 6070 3062 12046
rect 3004 6058 3062 6070
rect 3162 12046 3220 12058
rect 3162 6070 3174 12046
rect 3208 6070 3220 12046
rect 3162 6058 3220 6070
rect 3320 12046 3378 12058
rect 3320 6070 3332 12046
rect 3366 6070 3378 12046
rect 3320 6058 3378 6070
rect 3478 12046 3536 12058
rect 3478 6070 3490 12046
rect 3524 6070 3536 12046
rect 3478 6058 3536 6070
rect 3636 12046 3694 12058
rect 3636 6070 3648 12046
rect 3682 6070 3694 12046
rect 3636 6058 3694 6070
rect 3794 12046 3852 12058
rect 3794 6070 3806 12046
rect 3840 6070 3852 12046
rect 3794 6058 3852 6070
rect 3952 12046 4010 12058
rect 3952 6070 3964 12046
rect 3998 6070 4010 12046
rect 3952 6058 4010 6070
rect 4110 12046 4168 12058
rect 4110 6070 4122 12046
rect 4156 6070 4168 12046
rect 4110 6058 4168 6070
rect 5670 12046 5728 12058
rect 5670 6070 5682 12046
rect 5716 6070 5728 12046
rect 5670 6058 5728 6070
rect 5828 12046 5886 12058
rect 5828 6070 5840 12046
rect 5874 6070 5886 12046
rect 5828 6058 5886 6070
rect 5986 12046 6044 12058
rect 5986 6070 5998 12046
rect 6032 6070 6044 12046
rect 5986 6058 6044 6070
rect 6144 12046 6202 12058
rect 6144 6070 6156 12046
rect 6190 6070 6202 12046
rect 6144 6058 6202 6070
rect 6302 12046 6360 12058
rect 6302 6070 6314 12046
rect 6348 6070 6360 12046
rect 6302 6058 6360 6070
rect 6460 12046 6518 12058
rect 6460 6070 6472 12046
rect 6506 6070 6518 12046
rect 6460 6058 6518 6070
rect 6618 12046 6676 12058
rect 6618 6070 6630 12046
rect 6664 6070 6676 12046
rect 6618 6058 6676 6070
rect 6776 12046 6834 12058
rect 6776 6070 6788 12046
rect 6822 6070 6834 12046
rect 6776 6058 6834 6070
rect 6934 12046 6992 12058
rect 6934 6070 6946 12046
rect 6980 6070 6992 12046
rect 6934 6058 6992 6070
rect 7092 12046 7150 12058
rect 7092 6070 7104 12046
rect 7138 6070 7150 12046
rect 7092 6058 7150 6070
rect 7250 12046 7308 12058
rect 7250 6070 7262 12046
rect 7296 6070 7308 12046
rect 7250 6058 7308 6070
rect 7408 12046 7466 12058
rect 7408 6070 7420 12046
rect 7454 6070 7466 12046
rect 7408 6058 7466 6070
rect 7566 12046 7624 12058
rect 7566 6070 7578 12046
rect 7612 6070 7624 12046
rect 7566 6058 7624 6070
rect 7724 12046 7782 12058
rect 7724 6070 7736 12046
rect 7770 6070 7782 12046
rect 7724 6058 7782 6070
rect 7882 12046 7940 12058
rect 7882 6070 7894 12046
rect 7928 6070 7940 12046
rect 7882 6058 7940 6070
rect 8040 12046 8098 12058
rect 8040 6070 8052 12046
rect 8086 6070 8098 12046
rect 8040 6058 8098 6070
rect 8198 12046 8256 12058
rect 8198 6070 8210 12046
rect 8244 6070 8256 12046
rect 8198 6058 8256 6070
rect 8356 12046 8414 12058
rect 8356 6070 8368 12046
rect 8402 6070 8414 12046
rect 8356 6058 8414 6070
rect 8514 12046 8572 12058
rect 8514 6070 8526 12046
rect 8560 6070 8572 12046
rect 8514 6058 8572 6070
rect 8672 12046 8730 12058
rect 8672 6070 8684 12046
rect 8718 6070 8730 12046
rect 8672 6058 8730 6070
rect 8830 12046 8888 12058
rect 8830 6070 8842 12046
rect 8876 6070 8888 12046
rect 8830 6058 8888 6070
rect 8988 12046 9046 12058
rect 8988 6070 9000 12046
rect 9034 6070 9046 12046
rect 8988 6058 9046 6070
rect 9146 12046 9204 12058
rect 9146 6070 9158 12046
rect 9192 6070 9204 12046
rect 9146 6058 9204 6070
rect 9304 12046 9362 12058
rect 9304 6070 9316 12046
rect 9350 6070 9362 12046
rect 9304 6058 9362 6070
rect 9462 12046 9520 12058
rect 9462 6070 9474 12046
rect 9508 6070 9520 12046
rect 9462 6058 9520 6070
rect 9620 12046 9678 12058
rect 9620 6070 9632 12046
rect 9666 6070 9678 12046
rect 9620 6058 9678 6070
rect 9778 12046 9836 12058
rect 9778 6070 9790 12046
rect 9824 6070 9836 12046
rect 9778 6058 9836 6070
rect 9936 12046 9994 12058
rect 9936 6070 9948 12046
rect 9982 6070 9994 12046
rect 9936 6058 9994 6070
rect 10094 12046 10152 12058
rect 10094 6070 10106 12046
rect 10140 6070 10152 12046
rect 10094 6058 10152 6070
rect 10252 12046 10310 12058
rect 10252 6070 10264 12046
rect 10298 6070 10310 12046
rect 10252 6058 10310 6070
rect 10410 12046 10468 12058
rect 10410 6070 10422 12046
rect 10456 6070 10468 12046
rect 10410 6058 10468 6070
<< mvndiffc >>
rect -13218 43670 -13184 49646
rect -13060 43670 -13026 49646
rect -12902 43670 -12868 49646
rect -12744 43670 -12710 49646
rect -12586 43670 -12552 49646
rect -12428 43670 -12394 49646
rect -12270 43670 -12236 49646
rect -12112 43670 -12078 49646
rect -11954 43670 -11920 49646
rect -11796 43670 -11762 49646
rect -11638 43670 -11604 49646
rect -11480 43670 -11446 49646
rect -11322 43670 -11288 49646
rect -11164 43670 -11130 49646
rect -11006 43670 -10972 49646
rect -10848 43670 -10814 49646
rect -10690 43670 -10656 49646
rect -10532 43670 -10498 49646
rect -10374 43670 -10340 49646
rect -10216 43670 -10182 49646
rect -10058 43670 -10024 49646
rect -9900 43670 -9866 49646
rect -9742 43670 -9708 49646
rect -9584 43670 -9550 49646
rect -9426 43670 -9392 49646
rect -9268 43670 -9234 49646
rect -9110 43670 -9076 49646
rect -8952 43670 -8918 49646
rect -8794 43670 -8760 49646
rect -8636 43670 -8602 49646
rect -8478 43670 -8444 49646
rect -6918 43670 -6884 49646
rect -6760 43670 -6726 49646
rect -6602 43670 -6568 49646
rect -6444 43670 -6410 49646
rect -6286 43670 -6252 49646
rect -6128 43670 -6094 49646
rect -5970 43670 -5936 49646
rect -5812 43670 -5778 49646
rect -5654 43670 -5620 49646
rect -5496 43670 -5462 49646
rect -5338 43670 -5304 49646
rect -5180 43670 -5146 49646
rect -5022 43670 -4988 49646
rect -4864 43670 -4830 49646
rect -4706 43670 -4672 49646
rect -4548 43670 -4514 49646
rect -4390 43670 -4356 49646
rect -4232 43670 -4198 49646
rect -4074 43670 -4040 49646
rect -3916 43670 -3882 49646
rect -3758 43670 -3724 49646
rect -3600 43670 -3566 49646
rect -3442 43670 -3408 49646
rect -3284 43670 -3250 49646
rect -3126 43670 -3092 49646
rect -2968 43670 -2934 49646
rect -2810 43670 -2776 49646
rect -2652 43670 -2618 49646
rect -2494 43670 -2460 49646
rect -2336 43670 -2302 49646
rect -2178 43670 -2144 49646
rect -618 43670 -584 49646
rect -460 43670 -426 49646
rect -302 43670 -268 49646
rect -144 43670 -110 49646
rect 14 43670 48 49646
rect 172 43670 206 49646
rect 330 43670 364 49646
rect 488 43670 522 49646
rect 646 43670 680 49646
rect 804 43670 838 49646
rect 962 43670 996 49646
rect 1120 43670 1154 49646
rect 1278 43670 1312 49646
rect 1436 43670 1470 49646
rect 1594 43670 1628 49646
rect 1752 43670 1786 49646
rect 1910 43670 1944 49646
rect 2068 43670 2102 49646
rect 2226 43670 2260 49646
rect 2384 43670 2418 49646
rect 2542 43670 2576 49646
rect 2700 43670 2734 49646
rect 2858 43670 2892 49646
rect 3016 43670 3050 49646
rect 3174 43670 3208 49646
rect 3332 43670 3366 49646
rect 3490 43670 3524 49646
rect 3648 43670 3682 49646
rect 3806 43670 3840 49646
rect 3964 43670 3998 49646
rect 4122 43670 4156 49646
rect 5682 43670 5716 49646
rect 5840 43670 5874 49646
rect 5998 43670 6032 49646
rect 6156 43670 6190 49646
rect 6314 43670 6348 49646
rect 6472 43670 6506 49646
rect 6630 43670 6664 49646
rect 6788 43670 6822 49646
rect 6946 43670 6980 49646
rect 7104 43670 7138 49646
rect 7262 43670 7296 49646
rect 7420 43670 7454 49646
rect 7578 43670 7612 49646
rect 7736 43670 7770 49646
rect 7894 43670 7928 49646
rect 8052 43670 8086 49646
rect 8210 43670 8244 49646
rect 8368 43670 8402 49646
rect 8526 43670 8560 49646
rect 8684 43670 8718 49646
rect 8842 43670 8876 49646
rect 9000 43670 9034 49646
rect 9158 43670 9192 49646
rect 9316 43670 9350 49646
rect 9474 43670 9508 49646
rect 9632 43670 9666 49646
rect 9790 43670 9824 49646
rect 9948 43670 9982 49646
rect 10106 43670 10140 49646
rect 10264 43670 10298 49646
rect 10422 43670 10456 49646
rect -13218 36670 -13184 42646
rect -13060 36670 -13026 42646
rect -12902 36670 -12868 42646
rect -12744 36670 -12710 42646
rect -12586 36670 -12552 42646
rect -12428 36670 -12394 42646
rect -12270 36670 -12236 42646
rect -12112 36670 -12078 42646
rect -11954 36670 -11920 42646
rect -11796 36670 -11762 42646
rect -11638 36670 -11604 42646
rect -11480 36670 -11446 42646
rect -11322 36670 -11288 42646
rect -11164 36670 -11130 42646
rect -11006 36670 -10972 42646
rect -10848 36670 -10814 42646
rect -10690 36670 -10656 42646
rect -10532 36670 -10498 42646
rect -10374 36670 -10340 42646
rect -10216 36670 -10182 42646
rect -10058 36670 -10024 42646
rect -9900 36670 -9866 42646
rect -9742 36670 -9708 42646
rect -9584 36670 -9550 42646
rect -9426 36670 -9392 42646
rect -9268 36670 -9234 42646
rect -9110 36670 -9076 42646
rect -8952 36670 -8918 42646
rect -8794 36670 -8760 42646
rect -8636 36670 -8602 42646
rect -8478 36670 -8444 42646
rect -6918 36670 -6884 42646
rect -6760 36670 -6726 42646
rect -6602 36670 -6568 42646
rect -6444 36670 -6410 42646
rect -6286 36670 -6252 42646
rect -6128 36670 -6094 42646
rect -5970 36670 -5936 42646
rect -5812 36670 -5778 42646
rect -5654 36670 -5620 42646
rect -5496 36670 -5462 42646
rect -5338 36670 -5304 42646
rect -5180 36670 -5146 42646
rect -5022 36670 -4988 42646
rect -4864 36670 -4830 42646
rect -4706 36670 -4672 42646
rect -4548 36670 -4514 42646
rect -4390 36670 -4356 42646
rect -4232 36670 -4198 42646
rect -4074 36670 -4040 42646
rect -3916 36670 -3882 42646
rect -3758 36670 -3724 42646
rect -3600 36670 -3566 42646
rect -3442 36670 -3408 42646
rect -3284 36670 -3250 42646
rect -3126 36670 -3092 42646
rect -2968 36670 -2934 42646
rect -2810 36670 -2776 42646
rect -2652 36670 -2618 42646
rect -2494 36670 -2460 42646
rect -2336 36670 -2302 42646
rect -2178 36670 -2144 42646
rect -618 36670 -584 42646
rect -460 36670 -426 42646
rect -302 36670 -268 42646
rect -144 36670 -110 42646
rect 14 36670 48 42646
rect 172 36670 206 42646
rect 330 36670 364 42646
rect 488 36670 522 42646
rect 646 36670 680 42646
rect 804 36670 838 42646
rect 962 36670 996 42646
rect 1120 36670 1154 42646
rect 1278 36670 1312 42646
rect 1436 36670 1470 42646
rect 1594 36670 1628 42646
rect 1752 36670 1786 42646
rect 1910 36670 1944 42646
rect 2068 36670 2102 42646
rect 2226 36670 2260 42646
rect 2384 36670 2418 42646
rect 2542 36670 2576 42646
rect 2700 36670 2734 42646
rect 2858 36670 2892 42646
rect 3016 36670 3050 42646
rect 3174 36670 3208 42646
rect 3332 36670 3366 42646
rect 3490 36670 3524 42646
rect 3648 36670 3682 42646
rect 3806 36670 3840 42646
rect 3964 36670 3998 42646
rect 4122 36670 4156 42646
rect 5682 36670 5716 42646
rect 5840 36670 5874 42646
rect 5998 36670 6032 42646
rect 6156 36670 6190 42646
rect 6314 36670 6348 42646
rect 6472 36670 6506 42646
rect 6630 36670 6664 42646
rect 6788 36670 6822 42646
rect 6946 36670 6980 42646
rect 7104 36670 7138 42646
rect 7262 36670 7296 42646
rect 7420 36670 7454 42646
rect 7578 36670 7612 42646
rect 7736 36670 7770 42646
rect 7894 36670 7928 42646
rect 8052 36670 8086 42646
rect 8210 36670 8244 42646
rect 8368 36670 8402 42646
rect 8526 36670 8560 42646
rect 8684 36670 8718 42646
rect 8842 36670 8876 42646
rect 9000 36670 9034 42646
rect 9158 36670 9192 42646
rect 9316 36670 9350 42646
rect 9474 36670 9508 42646
rect 9632 36670 9666 42646
rect 9790 36670 9824 42646
rect 9948 36670 9982 42646
rect 10106 36670 10140 42646
rect 10264 36670 10298 42646
rect 10422 36670 10456 42646
rect -13218 28370 -13184 34346
rect -13060 28370 -13026 34346
rect -12902 28370 -12868 34346
rect -12744 28370 -12710 34346
rect -12586 28370 -12552 34346
rect -12428 28370 -12394 34346
rect -12270 28370 -12236 34346
rect -12112 28370 -12078 34346
rect -11954 28370 -11920 34346
rect -11796 28370 -11762 34346
rect -11638 28370 -11604 34346
rect -11480 28370 -11446 34346
rect -11322 28370 -11288 34346
rect -11164 28370 -11130 34346
rect -11006 28370 -10972 34346
rect -10848 28370 -10814 34346
rect -10690 28370 -10656 34346
rect -10532 28370 -10498 34346
rect -10374 28370 -10340 34346
rect -10216 28370 -10182 34346
rect -10058 28370 -10024 34346
rect -9900 28370 -9866 34346
rect -9742 28370 -9708 34346
rect -9584 28370 -9550 34346
rect -9426 28370 -9392 34346
rect -9268 28370 -9234 34346
rect -9110 28370 -9076 34346
rect -8952 28370 -8918 34346
rect -8794 28370 -8760 34346
rect -8636 28370 -8602 34346
rect -8478 28370 -8444 34346
rect -6918 28370 -6884 34346
rect -6760 28370 -6726 34346
rect -6602 28370 -6568 34346
rect -6444 28370 -6410 34346
rect -6286 28370 -6252 34346
rect -6128 28370 -6094 34346
rect -5970 28370 -5936 34346
rect -5812 28370 -5778 34346
rect -5654 28370 -5620 34346
rect -5496 28370 -5462 34346
rect -5338 28370 -5304 34346
rect -5180 28370 -5146 34346
rect -5022 28370 -4988 34346
rect -4864 28370 -4830 34346
rect -4706 28370 -4672 34346
rect -4548 28370 -4514 34346
rect -4390 28370 -4356 34346
rect -4232 28370 -4198 34346
rect -4074 28370 -4040 34346
rect -3916 28370 -3882 34346
rect -3758 28370 -3724 34346
rect -3600 28370 -3566 34346
rect -3442 28370 -3408 34346
rect -3284 28370 -3250 34346
rect -3126 28370 -3092 34346
rect -2968 28370 -2934 34346
rect -2810 28370 -2776 34346
rect -2652 28370 -2618 34346
rect -2494 28370 -2460 34346
rect -2336 28370 -2302 34346
rect -2178 28370 -2144 34346
rect -618 28370 -584 34346
rect -460 28370 -426 34346
rect -302 28370 -268 34346
rect -144 28370 -110 34346
rect 14 28370 48 34346
rect 172 28370 206 34346
rect 330 28370 364 34346
rect 488 28370 522 34346
rect 646 28370 680 34346
rect 804 28370 838 34346
rect 962 28370 996 34346
rect 1120 28370 1154 34346
rect 1278 28370 1312 34346
rect 1436 28370 1470 34346
rect 1594 28370 1628 34346
rect 1752 28370 1786 34346
rect 1910 28370 1944 34346
rect 2068 28370 2102 34346
rect 2226 28370 2260 34346
rect 2384 28370 2418 34346
rect 2542 28370 2576 34346
rect 2700 28370 2734 34346
rect 2858 28370 2892 34346
rect 3016 28370 3050 34346
rect 3174 28370 3208 34346
rect 3332 28370 3366 34346
rect 3490 28370 3524 34346
rect 3648 28370 3682 34346
rect 3806 28370 3840 34346
rect 3964 28370 3998 34346
rect 4122 28370 4156 34346
rect 5682 28370 5716 34346
rect 5840 28370 5874 34346
rect 5998 28370 6032 34346
rect 6156 28370 6190 34346
rect 6314 28370 6348 34346
rect 6472 28370 6506 34346
rect 6630 28370 6664 34346
rect 6788 28370 6822 34346
rect 6946 28370 6980 34346
rect 7104 28370 7138 34346
rect 7262 28370 7296 34346
rect 7420 28370 7454 34346
rect 7578 28370 7612 34346
rect 7736 28370 7770 34346
rect 7894 28370 7928 34346
rect 8052 28370 8086 34346
rect 8210 28370 8244 34346
rect 8368 28370 8402 34346
rect 8526 28370 8560 34346
rect 8684 28370 8718 34346
rect 8842 28370 8876 34346
rect 9000 28370 9034 34346
rect 9158 28370 9192 34346
rect 9316 28370 9350 34346
rect 9474 28370 9508 34346
rect 9632 28370 9666 34346
rect 9790 28370 9824 34346
rect 9948 28370 9982 34346
rect 10106 28370 10140 34346
rect 10264 28370 10298 34346
rect 10422 28370 10456 34346
rect -13218 21370 -13184 27346
rect -13060 21370 -13026 27346
rect -12902 21370 -12868 27346
rect -12744 21370 -12710 27346
rect -12586 21370 -12552 27346
rect -12428 21370 -12394 27346
rect -12270 21370 -12236 27346
rect -12112 21370 -12078 27346
rect -11954 21370 -11920 27346
rect -11796 21370 -11762 27346
rect -11638 21370 -11604 27346
rect -11480 21370 -11446 27346
rect -11322 21370 -11288 27346
rect -11164 21370 -11130 27346
rect -11006 21370 -10972 27346
rect -10848 21370 -10814 27346
rect -10690 21370 -10656 27346
rect -10532 21370 -10498 27346
rect -10374 21370 -10340 27346
rect -10216 21370 -10182 27346
rect -10058 21370 -10024 27346
rect -9900 21370 -9866 27346
rect -9742 21370 -9708 27346
rect -9584 21370 -9550 27346
rect -9426 21370 -9392 27346
rect -9268 21370 -9234 27346
rect -9110 21370 -9076 27346
rect -8952 21370 -8918 27346
rect -8794 21370 -8760 27346
rect -8636 21370 -8602 27346
rect -8478 21370 -8444 27346
rect -6918 21370 -6884 27346
rect -6760 21370 -6726 27346
rect -6602 21370 -6568 27346
rect -6444 21370 -6410 27346
rect -6286 21370 -6252 27346
rect -6128 21370 -6094 27346
rect -5970 21370 -5936 27346
rect -5812 21370 -5778 27346
rect -5654 21370 -5620 27346
rect -5496 21370 -5462 27346
rect -5338 21370 -5304 27346
rect -5180 21370 -5146 27346
rect -5022 21370 -4988 27346
rect -4864 21370 -4830 27346
rect -4706 21370 -4672 27346
rect -4548 21370 -4514 27346
rect -4390 21370 -4356 27346
rect -4232 21370 -4198 27346
rect -4074 21370 -4040 27346
rect -3916 21370 -3882 27346
rect -3758 21370 -3724 27346
rect -3600 21370 -3566 27346
rect -3442 21370 -3408 27346
rect -3284 21370 -3250 27346
rect -3126 21370 -3092 27346
rect -2968 21370 -2934 27346
rect -2810 21370 -2776 27346
rect -2652 21370 -2618 27346
rect -2494 21370 -2460 27346
rect -2336 21370 -2302 27346
rect -2178 21370 -2144 27346
rect -618 21370 -584 27346
rect -460 21370 -426 27346
rect -302 21370 -268 27346
rect -144 21370 -110 27346
rect 14 21370 48 27346
rect 172 21370 206 27346
rect 330 21370 364 27346
rect 488 21370 522 27346
rect 646 21370 680 27346
rect 804 21370 838 27346
rect 962 21370 996 27346
rect 1120 21370 1154 27346
rect 1278 21370 1312 27346
rect 1436 21370 1470 27346
rect 1594 21370 1628 27346
rect 1752 21370 1786 27346
rect 1910 21370 1944 27346
rect 2068 21370 2102 27346
rect 2226 21370 2260 27346
rect 2384 21370 2418 27346
rect 2542 21370 2576 27346
rect 2700 21370 2734 27346
rect 2858 21370 2892 27346
rect 3016 21370 3050 27346
rect 3174 21370 3208 27346
rect 3332 21370 3366 27346
rect 3490 21370 3524 27346
rect 3648 21370 3682 27346
rect 3806 21370 3840 27346
rect 3964 21370 3998 27346
rect 4122 21370 4156 27346
rect 5682 21370 5716 27346
rect 5840 21370 5874 27346
rect 5998 21370 6032 27346
rect 6156 21370 6190 27346
rect 6314 21370 6348 27346
rect 6472 21370 6506 27346
rect 6630 21370 6664 27346
rect 6788 21370 6822 27346
rect 6946 21370 6980 27346
rect 7104 21370 7138 27346
rect 7262 21370 7296 27346
rect 7420 21370 7454 27346
rect 7578 21370 7612 27346
rect 7736 21370 7770 27346
rect 7894 21370 7928 27346
rect 8052 21370 8086 27346
rect 8210 21370 8244 27346
rect 8368 21370 8402 27346
rect 8526 21370 8560 27346
rect 8684 21370 8718 27346
rect 8842 21370 8876 27346
rect 9000 21370 9034 27346
rect 9158 21370 9192 27346
rect 9316 21370 9350 27346
rect 9474 21370 9508 27346
rect 9632 21370 9666 27346
rect 9790 21370 9824 27346
rect 9948 21370 9982 27346
rect 10106 21370 10140 27346
rect 10264 21370 10298 27346
rect 10422 21370 10456 27346
rect -13218 13070 -13184 19046
rect -13060 13070 -13026 19046
rect -12902 13070 -12868 19046
rect -12744 13070 -12710 19046
rect -12586 13070 -12552 19046
rect -12428 13070 -12394 19046
rect -12270 13070 -12236 19046
rect -12112 13070 -12078 19046
rect -11954 13070 -11920 19046
rect -11796 13070 -11762 19046
rect -11638 13070 -11604 19046
rect -11480 13070 -11446 19046
rect -11322 13070 -11288 19046
rect -11164 13070 -11130 19046
rect -11006 13070 -10972 19046
rect -10848 13070 -10814 19046
rect -10690 13070 -10656 19046
rect -10532 13070 -10498 19046
rect -10374 13070 -10340 19046
rect -10216 13070 -10182 19046
rect -10058 13070 -10024 19046
rect -9900 13070 -9866 19046
rect -9742 13070 -9708 19046
rect -9584 13070 -9550 19046
rect -9426 13070 -9392 19046
rect -9268 13070 -9234 19046
rect -9110 13070 -9076 19046
rect -8952 13070 -8918 19046
rect -8794 13070 -8760 19046
rect -8636 13070 -8602 19046
rect -8478 13070 -8444 19046
rect -6918 13070 -6884 19046
rect -6760 13070 -6726 19046
rect -6602 13070 -6568 19046
rect -6444 13070 -6410 19046
rect -6286 13070 -6252 19046
rect -6128 13070 -6094 19046
rect -5970 13070 -5936 19046
rect -5812 13070 -5778 19046
rect -5654 13070 -5620 19046
rect -5496 13070 -5462 19046
rect -5338 13070 -5304 19046
rect -5180 13070 -5146 19046
rect -5022 13070 -4988 19046
rect -4864 13070 -4830 19046
rect -4706 13070 -4672 19046
rect -4548 13070 -4514 19046
rect -4390 13070 -4356 19046
rect -4232 13070 -4198 19046
rect -4074 13070 -4040 19046
rect -3916 13070 -3882 19046
rect -3758 13070 -3724 19046
rect -3600 13070 -3566 19046
rect -3442 13070 -3408 19046
rect -3284 13070 -3250 19046
rect -3126 13070 -3092 19046
rect -2968 13070 -2934 19046
rect -2810 13070 -2776 19046
rect -2652 13070 -2618 19046
rect -2494 13070 -2460 19046
rect -2336 13070 -2302 19046
rect -2178 13070 -2144 19046
rect -618 13070 -584 19046
rect -460 13070 -426 19046
rect -302 13070 -268 19046
rect -144 13070 -110 19046
rect 14 13070 48 19046
rect 172 13070 206 19046
rect 330 13070 364 19046
rect 488 13070 522 19046
rect 646 13070 680 19046
rect 804 13070 838 19046
rect 962 13070 996 19046
rect 1120 13070 1154 19046
rect 1278 13070 1312 19046
rect 1436 13070 1470 19046
rect 1594 13070 1628 19046
rect 1752 13070 1786 19046
rect 1910 13070 1944 19046
rect 2068 13070 2102 19046
rect 2226 13070 2260 19046
rect 2384 13070 2418 19046
rect 2542 13070 2576 19046
rect 2700 13070 2734 19046
rect 2858 13070 2892 19046
rect 3016 13070 3050 19046
rect 3174 13070 3208 19046
rect 3332 13070 3366 19046
rect 3490 13070 3524 19046
rect 3648 13070 3682 19046
rect 3806 13070 3840 19046
rect 3964 13070 3998 19046
rect 4122 13070 4156 19046
rect 5682 13070 5716 19046
rect 5840 13070 5874 19046
rect 5998 13070 6032 19046
rect 6156 13070 6190 19046
rect 6314 13070 6348 19046
rect 6472 13070 6506 19046
rect 6630 13070 6664 19046
rect 6788 13070 6822 19046
rect 6946 13070 6980 19046
rect 7104 13070 7138 19046
rect 7262 13070 7296 19046
rect 7420 13070 7454 19046
rect 7578 13070 7612 19046
rect 7736 13070 7770 19046
rect 7894 13070 7928 19046
rect 8052 13070 8086 19046
rect 8210 13070 8244 19046
rect 8368 13070 8402 19046
rect 8526 13070 8560 19046
rect 8684 13070 8718 19046
rect 8842 13070 8876 19046
rect 9000 13070 9034 19046
rect 9158 13070 9192 19046
rect 9316 13070 9350 19046
rect 9474 13070 9508 19046
rect 9632 13070 9666 19046
rect 9790 13070 9824 19046
rect 9948 13070 9982 19046
rect 10106 13070 10140 19046
rect 10264 13070 10298 19046
rect 10422 13070 10456 19046
rect -13218 6070 -13184 12046
rect -13060 6070 -13026 12046
rect -12902 6070 -12868 12046
rect -12744 6070 -12710 12046
rect -12586 6070 -12552 12046
rect -12428 6070 -12394 12046
rect -12270 6070 -12236 12046
rect -12112 6070 -12078 12046
rect -11954 6070 -11920 12046
rect -11796 6070 -11762 12046
rect -11638 6070 -11604 12046
rect -11480 6070 -11446 12046
rect -11322 6070 -11288 12046
rect -11164 6070 -11130 12046
rect -11006 6070 -10972 12046
rect -10848 6070 -10814 12046
rect -10690 6070 -10656 12046
rect -10532 6070 -10498 12046
rect -10374 6070 -10340 12046
rect -10216 6070 -10182 12046
rect -10058 6070 -10024 12046
rect -9900 6070 -9866 12046
rect -9742 6070 -9708 12046
rect -9584 6070 -9550 12046
rect -9426 6070 -9392 12046
rect -9268 6070 -9234 12046
rect -9110 6070 -9076 12046
rect -8952 6070 -8918 12046
rect -8794 6070 -8760 12046
rect -8636 6070 -8602 12046
rect -8478 6070 -8444 12046
rect -6918 6070 -6884 12046
rect -6760 6070 -6726 12046
rect -6602 6070 -6568 12046
rect -6444 6070 -6410 12046
rect -6286 6070 -6252 12046
rect -6128 6070 -6094 12046
rect -5970 6070 -5936 12046
rect -5812 6070 -5778 12046
rect -5654 6070 -5620 12046
rect -5496 6070 -5462 12046
rect -5338 6070 -5304 12046
rect -5180 6070 -5146 12046
rect -5022 6070 -4988 12046
rect -4864 6070 -4830 12046
rect -4706 6070 -4672 12046
rect -4548 6070 -4514 12046
rect -4390 6070 -4356 12046
rect -4232 6070 -4198 12046
rect -4074 6070 -4040 12046
rect -3916 6070 -3882 12046
rect -3758 6070 -3724 12046
rect -3600 6070 -3566 12046
rect -3442 6070 -3408 12046
rect -3284 6070 -3250 12046
rect -3126 6070 -3092 12046
rect -2968 6070 -2934 12046
rect -2810 6070 -2776 12046
rect -2652 6070 -2618 12046
rect -2494 6070 -2460 12046
rect -2336 6070 -2302 12046
rect -2178 6070 -2144 12046
rect -618 6070 -584 12046
rect -460 6070 -426 12046
rect -302 6070 -268 12046
rect -144 6070 -110 12046
rect 14 6070 48 12046
rect 172 6070 206 12046
rect 330 6070 364 12046
rect 488 6070 522 12046
rect 646 6070 680 12046
rect 804 6070 838 12046
rect 962 6070 996 12046
rect 1120 6070 1154 12046
rect 1278 6070 1312 12046
rect 1436 6070 1470 12046
rect 1594 6070 1628 12046
rect 1752 6070 1786 12046
rect 1910 6070 1944 12046
rect 2068 6070 2102 12046
rect 2226 6070 2260 12046
rect 2384 6070 2418 12046
rect 2542 6070 2576 12046
rect 2700 6070 2734 12046
rect 2858 6070 2892 12046
rect 3016 6070 3050 12046
rect 3174 6070 3208 12046
rect 3332 6070 3366 12046
rect 3490 6070 3524 12046
rect 3648 6070 3682 12046
rect 3806 6070 3840 12046
rect 3964 6070 3998 12046
rect 4122 6070 4156 12046
rect 5682 6070 5716 12046
rect 5840 6070 5874 12046
rect 5998 6070 6032 12046
rect 6156 6070 6190 12046
rect 6314 6070 6348 12046
rect 6472 6070 6506 12046
rect 6630 6070 6664 12046
rect 6788 6070 6822 12046
rect 6946 6070 6980 12046
rect 7104 6070 7138 12046
rect 7262 6070 7296 12046
rect 7420 6070 7454 12046
rect 7578 6070 7612 12046
rect 7736 6070 7770 12046
rect 7894 6070 7928 12046
rect 8052 6070 8086 12046
rect 8210 6070 8244 12046
rect 8368 6070 8402 12046
rect 8526 6070 8560 12046
rect 8684 6070 8718 12046
rect 8842 6070 8876 12046
rect 9000 6070 9034 12046
rect 9158 6070 9192 12046
rect 9316 6070 9350 12046
rect 9474 6070 9508 12046
rect 9632 6070 9666 12046
rect 9790 6070 9824 12046
rect 9948 6070 9982 12046
rect 10106 6070 10140 12046
rect 10264 6070 10298 12046
rect 10422 6070 10456 12046
<< mvpsubdiff >>
rect -13364 49868 -8298 49880
rect -13364 49834 -13256 49868
rect -8406 49834 -8298 49868
rect -13364 49822 -8298 49834
rect -13364 49772 -13306 49822
rect -13364 43544 -13352 49772
rect -13318 43544 -13306 49772
rect -8356 49772 -8298 49822
rect -13364 43494 -13306 43544
rect -8356 43544 -8344 49772
rect -8310 43544 -8298 49772
rect -8356 43494 -8298 43544
rect -13364 43482 -8298 43494
rect -13364 43448 -13256 43482
rect -8406 43448 -8298 43482
rect -13364 43436 -8298 43448
rect -7064 49868 -1998 49880
rect -7064 49834 -6956 49868
rect -2106 49834 -1998 49868
rect -7064 49822 -1998 49834
rect -7064 49772 -7006 49822
rect -7064 43544 -7052 49772
rect -7018 43544 -7006 49772
rect -2056 49772 -1998 49822
rect -7064 43494 -7006 43544
rect -2056 43544 -2044 49772
rect -2010 43544 -1998 49772
rect -2056 43494 -1998 43544
rect -7064 43482 -1998 43494
rect -7064 43448 -6956 43482
rect -2106 43448 -1998 43482
rect -7064 43436 -1998 43448
rect -764 49868 4302 49880
rect -764 49834 -656 49868
rect 4194 49834 4302 49868
rect -764 49822 4302 49834
rect -764 49772 -706 49822
rect -764 43544 -752 49772
rect -718 43544 -706 49772
rect 4244 49772 4302 49822
rect -764 43494 -706 43544
rect 4244 43544 4256 49772
rect 4290 43544 4302 49772
rect 4244 43494 4302 43544
rect -764 43482 4302 43494
rect -764 43448 -656 43482
rect 4194 43448 4302 43482
rect -764 43436 4302 43448
rect 5536 49868 10602 49880
rect 5536 49834 5644 49868
rect 10494 49834 10602 49868
rect 5536 49822 10602 49834
rect 5536 49772 5594 49822
rect 5536 43544 5548 49772
rect 5582 43544 5594 49772
rect 10544 49772 10602 49822
rect 5536 43494 5594 43544
rect 10544 43544 10556 49772
rect 10590 43544 10602 49772
rect 10544 43494 10602 43544
rect 5536 43482 10602 43494
rect 5536 43448 5644 43482
rect 10494 43448 10602 43482
rect 5536 43436 10602 43448
rect -13364 42868 -8298 42880
rect -13364 42834 -13256 42868
rect -8406 42834 -8298 42868
rect -13364 42822 -8298 42834
rect -13364 42772 -13306 42822
rect -13364 36544 -13352 42772
rect -13318 36544 -13306 42772
rect -8356 42772 -8298 42822
rect -13364 36494 -13306 36544
rect -8356 36544 -8344 42772
rect -8310 36544 -8298 42772
rect -8356 36494 -8298 36544
rect -13364 36482 -8298 36494
rect -13364 36448 -13256 36482
rect -8406 36448 -8298 36482
rect -13364 36436 -8298 36448
rect -7064 42868 -1998 42880
rect -7064 42834 -6956 42868
rect -2106 42834 -1998 42868
rect -7064 42822 -1998 42834
rect -7064 42772 -7006 42822
rect -7064 36544 -7052 42772
rect -7018 36544 -7006 42772
rect -2056 42772 -1998 42822
rect -7064 36494 -7006 36544
rect -2056 36544 -2044 42772
rect -2010 36544 -1998 42772
rect -2056 36494 -1998 36544
rect -7064 36482 -1998 36494
rect -7064 36448 -6956 36482
rect -2106 36448 -1998 36482
rect -7064 36436 -1998 36448
rect -764 42868 4302 42880
rect -764 42834 -656 42868
rect 4194 42834 4302 42868
rect -764 42822 4302 42834
rect -764 42772 -706 42822
rect -764 36544 -752 42772
rect -718 36544 -706 42772
rect 4244 42772 4302 42822
rect -764 36494 -706 36544
rect 4244 36544 4256 42772
rect 4290 36544 4302 42772
rect 4244 36494 4302 36544
rect -764 36482 4302 36494
rect -764 36448 -656 36482
rect 4194 36448 4302 36482
rect -764 36436 4302 36448
rect 5536 42868 10602 42880
rect 5536 42834 5644 42868
rect 10494 42834 10602 42868
rect 5536 42822 10602 42834
rect 5536 42772 5594 42822
rect 5536 36544 5548 42772
rect 5582 36544 5594 42772
rect 10544 42772 10602 42822
rect 5536 36494 5594 36544
rect 10544 36544 10556 42772
rect 10590 36544 10602 42772
rect 10544 36494 10602 36544
rect 5536 36482 10602 36494
rect 5536 36448 5644 36482
rect 10494 36448 10602 36482
rect 5536 36436 10602 36448
rect -13364 34568 -8298 34580
rect -13364 34534 -13256 34568
rect -8406 34534 -8298 34568
rect -13364 34522 -8298 34534
rect -13364 34472 -13306 34522
rect -13364 28244 -13352 34472
rect -13318 28244 -13306 34472
rect -8356 34472 -8298 34522
rect -13364 28194 -13306 28244
rect -8356 28244 -8344 34472
rect -8310 28244 -8298 34472
rect -8356 28194 -8298 28244
rect -13364 28182 -8298 28194
rect -13364 28148 -13256 28182
rect -8406 28148 -8298 28182
rect -13364 28136 -8298 28148
rect -7064 34568 -1998 34580
rect -7064 34534 -6956 34568
rect -2106 34534 -1998 34568
rect -7064 34522 -1998 34534
rect -7064 34472 -7006 34522
rect -7064 28244 -7052 34472
rect -7018 28244 -7006 34472
rect -2056 34472 -1998 34522
rect -7064 28194 -7006 28244
rect -2056 28244 -2044 34472
rect -2010 28244 -1998 34472
rect -2056 28194 -1998 28244
rect -7064 28182 -1998 28194
rect -7064 28148 -6956 28182
rect -2106 28148 -1998 28182
rect -7064 28136 -1998 28148
rect -764 34568 4302 34580
rect -764 34534 -656 34568
rect 4194 34534 4302 34568
rect -764 34522 4302 34534
rect -764 34472 -706 34522
rect -764 28244 -752 34472
rect -718 28244 -706 34472
rect 4244 34472 4302 34522
rect -764 28194 -706 28244
rect 4244 28244 4256 34472
rect 4290 28244 4302 34472
rect 4244 28194 4302 28244
rect -764 28182 4302 28194
rect -764 28148 -656 28182
rect 4194 28148 4302 28182
rect -764 28136 4302 28148
rect 5536 34568 10602 34580
rect 5536 34534 5644 34568
rect 10494 34534 10602 34568
rect 5536 34522 10602 34534
rect 5536 34472 5594 34522
rect 5536 28244 5548 34472
rect 5582 28244 5594 34472
rect 10544 34472 10602 34522
rect 5536 28194 5594 28244
rect 10544 28244 10556 34472
rect 10590 28244 10602 34472
rect 10544 28194 10602 28244
rect 5536 28182 10602 28194
rect 5536 28148 5644 28182
rect 10494 28148 10602 28182
rect 5536 28136 10602 28148
rect -13364 27568 -8298 27580
rect -13364 27534 -13256 27568
rect -8406 27534 -8298 27568
rect -13364 27522 -8298 27534
rect -13364 27472 -13306 27522
rect -13364 21244 -13352 27472
rect -13318 21244 -13306 27472
rect -8356 27472 -8298 27522
rect -13364 21194 -13306 21244
rect -8356 21244 -8344 27472
rect -8310 21244 -8298 27472
rect -8356 21194 -8298 21244
rect -13364 21182 -8298 21194
rect -13364 21148 -13256 21182
rect -8406 21148 -8298 21182
rect -13364 21136 -8298 21148
rect -7064 27568 -1998 27580
rect -7064 27534 -6956 27568
rect -2106 27534 -1998 27568
rect -7064 27522 -1998 27534
rect -7064 27472 -7006 27522
rect -7064 21244 -7052 27472
rect -7018 21244 -7006 27472
rect -2056 27472 -1998 27522
rect -7064 21194 -7006 21244
rect -2056 21244 -2044 27472
rect -2010 21244 -1998 27472
rect -2056 21194 -1998 21244
rect -7064 21182 -1998 21194
rect -7064 21148 -6956 21182
rect -2106 21148 -1998 21182
rect -7064 21136 -1998 21148
rect -764 27568 4302 27580
rect -764 27534 -656 27568
rect 4194 27534 4302 27568
rect -764 27522 4302 27534
rect -764 27472 -706 27522
rect -764 21244 -752 27472
rect -718 21244 -706 27472
rect 4244 27472 4302 27522
rect -764 21194 -706 21244
rect 4244 21244 4256 27472
rect 4290 21244 4302 27472
rect 4244 21194 4302 21244
rect -764 21182 4302 21194
rect -764 21148 -656 21182
rect 4194 21148 4302 21182
rect -764 21136 4302 21148
rect 5536 27568 10602 27580
rect 5536 27534 5644 27568
rect 10494 27534 10602 27568
rect 5536 27522 10602 27534
rect 5536 27472 5594 27522
rect 5536 21244 5548 27472
rect 5582 21244 5594 27472
rect 10544 27472 10602 27522
rect 5536 21194 5594 21244
rect 10544 21244 10556 27472
rect 10590 21244 10602 27472
rect 10544 21194 10602 21244
rect 5536 21182 10602 21194
rect 5536 21148 5644 21182
rect 10494 21148 10602 21182
rect 5536 21136 10602 21148
rect -13364 19268 -8298 19280
rect -13364 19234 -13256 19268
rect -8406 19234 -8298 19268
rect -13364 19222 -8298 19234
rect -13364 19172 -13306 19222
rect -13364 12944 -13352 19172
rect -13318 12944 -13306 19172
rect -8356 19172 -8298 19222
rect -13364 12894 -13306 12944
rect -8356 12944 -8344 19172
rect -8310 12944 -8298 19172
rect -8356 12894 -8298 12944
rect -13364 12882 -8298 12894
rect -13364 12848 -13256 12882
rect -8406 12848 -8298 12882
rect -13364 12836 -8298 12848
rect -7064 19268 -1998 19280
rect -7064 19234 -6956 19268
rect -2106 19234 -1998 19268
rect -7064 19222 -1998 19234
rect -7064 19172 -7006 19222
rect -7064 12944 -7052 19172
rect -7018 12944 -7006 19172
rect -2056 19172 -1998 19222
rect -7064 12894 -7006 12944
rect -2056 12944 -2044 19172
rect -2010 12944 -1998 19172
rect -2056 12894 -1998 12944
rect -7064 12882 -1998 12894
rect -7064 12848 -6956 12882
rect -2106 12848 -1998 12882
rect -7064 12836 -1998 12848
rect -764 19268 4302 19280
rect -764 19234 -656 19268
rect 4194 19234 4302 19268
rect -764 19222 4302 19234
rect -764 19172 -706 19222
rect -764 12944 -752 19172
rect -718 12944 -706 19172
rect 4244 19172 4302 19222
rect -764 12894 -706 12944
rect 4244 12944 4256 19172
rect 4290 12944 4302 19172
rect 4244 12894 4302 12944
rect -764 12882 4302 12894
rect -764 12848 -656 12882
rect 4194 12848 4302 12882
rect -764 12836 4302 12848
rect 5536 19268 10602 19280
rect 5536 19234 5644 19268
rect 10494 19234 10602 19268
rect 5536 19222 10602 19234
rect 5536 19172 5594 19222
rect 5536 12944 5548 19172
rect 5582 12944 5594 19172
rect 10544 19172 10602 19222
rect 5536 12894 5594 12944
rect 10544 12944 10556 19172
rect 10590 12944 10602 19172
rect 10544 12894 10602 12944
rect 5536 12882 10602 12894
rect 5536 12848 5644 12882
rect 10494 12848 10602 12882
rect 5536 12836 10602 12848
rect -13364 12268 -8298 12280
rect -13364 12234 -13256 12268
rect -8406 12234 -8298 12268
rect -13364 12222 -8298 12234
rect -13364 12172 -13306 12222
rect -13364 5944 -13352 12172
rect -13318 5944 -13306 12172
rect -8356 12172 -8298 12222
rect -13364 5894 -13306 5944
rect -8356 5944 -8344 12172
rect -8310 5944 -8298 12172
rect -8356 5894 -8298 5944
rect -13364 5882 -8298 5894
rect -13364 5848 -13256 5882
rect -8406 5848 -8298 5882
rect -13364 5836 -8298 5848
rect -7064 12268 -1998 12280
rect -7064 12234 -6956 12268
rect -2106 12234 -1998 12268
rect -7064 12222 -1998 12234
rect -7064 12172 -7006 12222
rect -7064 5944 -7052 12172
rect -7018 5944 -7006 12172
rect -2056 12172 -1998 12222
rect -7064 5894 -7006 5944
rect -2056 5944 -2044 12172
rect -2010 5944 -1998 12172
rect -2056 5894 -1998 5944
rect -7064 5882 -1998 5894
rect -7064 5848 -6956 5882
rect -2106 5848 -1998 5882
rect -7064 5836 -1998 5848
rect -764 12268 4302 12280
rect -764 12234 -656 12268
rect 4194 12234 4302 12268
rect -764 12222 4302 12234
rect -764 12172 -706 12222
rect -764 5944 -752 12172
rect -718 5944 -706 12172
rect 4244 12172 4302 12222
rect -764 5894 -706 5944
rect 4244 5944 4256 12172
rect 4290 5944 4302 12172
rect 4244 5894 4302 5944
rect -764 5882 4302 5894
rect -764 5848 -656 5882
rect 4194 5848 4302 5882
rect -764 5836 4302 5848
rect 5536 12268 10602 12280
rect 5536 12234 5644 12268
rect 10494 12234 10602 12268
rect 5536 12222 10602 12234
rect 5536 12172 5594 12222
rect 5536 5944 5548 12172
rect 5582 5944 5594 12172
rect 10544 12172 10602 12222
rect 5536 5894 5594 5944
rect 10544 5944 10556 12172
rect 10590 5944 10602 12172
rect 10544 5894 10602 5944
rect 5536 5882 10602 5894
rect 5536 5848 5644 5882
rect 10494 5848 10602 5882
rect 5536 5836 10602 5848
<< mvpsubdiffcont >>
rect -13256 49834 -8406 49868
rect -13352 43544 -13318 49772
rect -8344 43544 -8310 49772
rect -13256 43448 -8406 43482
rect -6956 49834 -2106 49868
rect -7052 43544 -7018 49772
rect -2044 43544 -2010 49772
rect -6956 43448 -2106 43482
rect -656 49834 4194 49868
rect -752 43544 -718 49772
rect 4256 43544 4290 49772
rect -656 43448 4194 43482
rect 5644 49834 10494 49868
rect 5548 43544 5582 49772
rect 10556 43544 10590 49772
rect 5644 43448 10494 43482
rect -13256 42834 -8406 42868
rect -13352 36544 -13318 42772
rect -8344 36544 -8310 42772
rect -13256 36448 -8406 36482
rect -6956 42834 -2106 42868
rect -7052 36544 -7018 42772
rect -2044 36544 -2010 42772
rect -6956 36448 -2106 36482
rect -656 42834 4194 42868
rect -752 36544 -718 42772
rect 4256 36544 4290 42772
rect -656 36448 4194 36482
rect 5644 42834 10494 42868
rect 5548 36544 5582 42772
rect 10556 36544 10590 42772
rect 5644 36448 10494 36482
rect -13256 34534 -8406 34568
rect -13352 28244 -13318 34472
rect -8344 28244 -8310 34472
rect -13256 28148 -8406 28182
rect -6956 34534 -2106 34568
rect -7052 28244 -7018 34472
rect -2044 28244 -2010 34472
rect -6956 28148 -2106 28182
rect -656 34534 4194 34568
rect -752 28244 -718 34472
rect 4256 28244 4290 34472
rect -656 28148 4194 28182
rect 5644 34534 10494 34568
rect 5548 28244 5582 34472
rect 10556 28244 10590 34472
rect 5644 28148 10494 28182
rect -13256 27534 -8406 27568
rect -13352 21244 -13318 27472
rect -8344 21244 -8310 27472
rect -13256 21148 -8406 21182
rect -6956 27534 -2106 27568
rect -7052 21244 -7018 27472
rect -2044 21244 -2010 27472
rect -6956 21148 -2106 21182
rect -656 27534 4194 27568
rect -752 21244 -718 27472
rect 4256 21244 4290 27472
rect -656 21148 4194 21182
rect 5644 27534 10494 27568
rect 5548 21244 5582 27472
rect 10556 21244 10590 27472
rect 5644 21148 10494 21182
rect -13256 19234 -8406 19268
rect -13352 12944 -13318 19172
rect -8344 12944 -8310 19172
rect -13256 12848 -8406 12882
rect -6956 19234 -2106 19268
rect -7052 12944 -7018 19172
rect -2044 12944 -2010 19172
rect -6956 12848 -2106 12882
rect -656 19234 4194 19268
rect -752 12944 -718 19172
rect 4256 12944 4290 19172
rect -656 12848 4194 12882
rect 5644 19234 10494 19268
rect 5548 12944 5582 19172
rect 10556 12944 10590 19172
rect 5644 12848 10494 12882
rect -13256 12234 -8406 12268
rect -13352 5944 -13318 12172
rect -8344 5944 -8310 12172
rect -13256 5848 -8406 5882
rect -6956 12234 -2106 12268
rect -7052 5944 -7018 12172
rect -2044 5944 -2010 12172
rect -6956 5848 -2106 5882
rect -656 12234 4194 12268
rect -752 5944 -718 12172
rect 4256 5944 4290 12172
rect -656 5848 4194 5882
rect 5644 12234 10494 12268
rect 5548 5944 5582 12172
rect 10556 5944 10590 12172
rect 5644 5848 10494 5882
<< poly >>
rect -13172 49730 -13072 49746
rect -13172 49696 -13156 49730
rect -13088 49696 -13072 49730
rect -13172 49658 -13072 49696
rect -13014 49730 -12914 49746
rect -13014 49696 -12998 49730
rect -12930 49696 -12914 49730
rect -13014 49658 -12914 49696
rect -12856 49730 -12756 49746
rect -12856 49696 -12840 49730
rect -12772 49696 -12756 49730
rect -12856 49658 -12756 49696
rect -12698 49730 -12598 49746
rect -12698 49696 -12682 49730
rect -12614 49696 -12598 49730
rect -12698 49658 -12598 49696
rect -12540 49730 -12440 49746
rect -12540 49696 -12524 49730
rect -12456 49696 -12440 49730
rect -12540 49658 -12440 49696
rect -12382 49730 -12282 49746
rect -12382 49696 -12366 49730
rect -12298 49696 -12282 49730
rect -12382 49658 -12282 49696
rect -12224 49730 -12124 49746
rect -12224 49696 -12208 49730
rect -12140 49696 -12124 49730
rect -12224 49658 -12124 49696
rect -12066 49730 -11966 49746
rect -12066 49696 -12050 49730
rect -11982 49696 -11966 49730
rect -12066 49658 -11966 49696
rect -11908 49730 -11808 49746
rect -11908 49696 -11892 49730
rect -11824 49696 -11808 49730
rect -11908 49658 -11808 49696
rect -11750 49730 -11650 49746
rect -11750 49696 -11734 49730
rect -11666 49696 -11650 49730
rect -11750 49658 -11650 49696
rect -11592 49730 -11492 49746
rect -11592 49696 -11576 49730
rect -11508 49696 -11492 49730
rect -11592 49658 -11492 49696
rect -11434 49730 -11334 49746
rect -11434 49696 -11418 49730
rect -11350 49696 -11334 49730
rect -11434 49658 -11334 49696
rect -11276 49730 -11176 49746
rect -11276 49696 -11260 49730
rect -11192 49696 -11176 49730
rect -11276 49658 -11176 49696
rect -11118 49730 -11018 49746
rect -11118 49696 -11102 49730
rect -11034 49696 -11018 49730
rect -11118 49658 -11018 49696
rect -10960 49730 -10860 49746
rect -10960 49696 -10944 49730
rect -10876 49696 -10860 49730
rect -10960 49658 -10860 49696
rect -10802 49730 -10702 49746
rect -10802 49696 -10786 49730
rect -10718 49696 -10702 49730
rect -10802 49658 -10702 49696
rect -10644 49730 -10544 49746
rect -10644 49696 -10628 49730
rect -10560 49696 -10544 49730
rect -10644 49658 -10544 49696
rect -10486 49730 -10386 49746
rect -10486 49696 -10470 49730
rect -10402 49696 -10386 49730
rect -10486 49658 -10386 49696
rect -10328 49730 -10228 49746
rect -10328 49696 -10312 49730
rect -10244 49696 -10228 49730
rect -10328 49658 -10228 49696
rect -10170 49730 -10070 49746
rect -10170 49696 -10154 49730
rect -10086 49696 -10070 49730
rect -10170 49658 -10070 49696
rect -10012 49730 -9912 49746
rect -10012 49696 -9996 49730
rect -9928 49696 -9912 49730
rect -10012 49658 -9912 49696
rect -9854 49730 -9754 49746
rect -9854 49696 -9838 49730
rect -9770 49696 -9754 49730
rect -9854 49658 -9754 49696
rect -9696 49730 -9596 49746
rect -9696 49696 -9680 49730
rect -9612 49696 -9596 49730
rect -9696 49658 -9596 49696
rect -9538 49730 -9438 49746
rect -9538 49696 -9522 49730
rect -9454 49696 -9438 49730
rect -9538 49658 -9438 49696
rect -9380 49730 -9280 49746
rect -9380 49696 -9364 49730
rect -9296 49696 -9280 49730
rect -9380 49658 -9280 49696
rect -9222 49730 -9122 49746
rect -9222 49696 -9206 49730
rect -9138 49696 -9122 49730
rect -9222 49658 -9122 49696
rect -9064 49730 -8964 49746
rect -9064 49696 -9048 49730
rect -8980 49696 -8964 49730
rect -9064 49658 -8964 49696
rect -8906 49730 -8806 49746
rect -8906 49696 -8890 49730
rect -8822 49696 -8806 49730
rect -8906 49658 -8806 49696
rect -8748 49730 -8648 49746
rect -8748 49696 -8732 49730
rect -8664 49696 -8648 49730
rect -8748 49658 -8648 49696
rect -8590 49730 -8490 49746
rect -8590 49696 -8574 49730
rect -8506 49696 -8490 49730
rect -8590 49658 -8490 49696
rect -13172 43620 -13072 43658
rect -13172 43586 -13156 43620
rect -13088 43586 -13072 43620
rect -13172 43570 -13072 43586
rect -13014 43620 -12914 43658
rect -13014 43586 -12998 43620
rect -12930 43586 -12914 43620
rect -13014 43570 -12914 43586
rect -12856 43620 -12756 43658
rect -12856 43586 -12840 43620
rect -12772 43586 -12756 43620
rect -12856 43570 -12756 43586
rect -12698 43620 -12598 43658
rect -12698 43586 -12682 43620
rect -12614 43586 -12598 43620
rect -12698 43570 -12598 43586
rect -12540 43620 -12440 43658
rect -12540 43586 -12524 43620
rect -12456 43586 -12440 43620
rect -12540 43570 -12440 43586
rect -12382 43620 -12282 43658
rect -12382 43586 -12366 43620
rect -12298 43586 -12282 43620
rect -12382 43570 -12282 43586
rect -12224 43620 -12124 43658
rect -12224 43586 -12208 43620
rect -12140 43586 -12124 43620
rect -12224 43570 -12124 43586
rect -12066 43620 -11966 43658
rect -12066 43586 -12050 43620
rect -11982 43586 -11966 43620
rect -12066 43570 -11966 43586
rect -11908 43620 -11808 43658
rect -11908 43586 -11892 43620
rect -11824 43586 -11808 43620
rect -11908 43570 -11808 43586
rect -11750 43620 -11650 43658
rect -11750 43586 -11734 43620
rect -11666 43586 -11650 43620
rect -11750 43570 -11650 43586
rect -11592 43620 -11492 43658
rect -11592 43586 -11576 43620
rect -11508 43586 -11492 43620
rect -11592 43570 -11492 43586
rect -11434 43620 -11334 43658
rect -11434 43586 -11418 43620
rect -11350 43586 -11334 43620
rect -11434 43570 -11334 43586
rect -11276 43620 -11176 43658
rect -11276 43586 -11260 43620
rect -11192 43586 -11176 43620
rect -11276 43570 -11176 43586
rect -11118 43620 -11018 43658
rect -11118 43586 -11102 43620
rect -11034 43586 -11018 43620
rect -11118 43570 -11018 43586
rect -10960 43620 -10860 43658
rect -10960 43586 -10944 43620
rect -10876 43586 -10860 43620
rect -10960 43570 -10860 43586
rect -10802 43620 -10702 43658
rect -10802 43586 -10786 43620
rect -10718 43586 -10702 43620
rect -10802 43570 -10702 43586
rect -10644 43620 -10544 43658
rect -10644 43586 -10628 43620
rect -10560 43586 -10544 43620
rect -10644 43570 -10544 43586
rect -10486 43620 -10386 43658
rect -10486 43586 -10470 43620
rect -10402 43586 -10386 43620
rect -10486 43570 -10386 43586
rect -10328 43620 -10228 43658
rect -10328 43586 -10312 43620
rect -10244 43586 -10228 43620
rect -10328 43570 -10228 43586
rect -10170 43620 -10070 43658
rect -10170 43586 -10154 43620
rect -10086 43586 -10070 43620
rect -10170 43570 -10070 43586
rect -10012 43620 -9912 43658
rect -10012 43586 -9996 43620
rect -9928 43586 -9912 43620
rect -10012 43570 -9912 43586
rect -9854 43620 -9754 43658
rect -9854 43586 -9838 43620
rect -9770 43586 -9754 43620
rect -9854 43570 -9754 43586
rect -9696 43620 -9596 43658
rect -9696 43586 -9680 43620
rect -9612 43586 -9596 43620
rect -9696 43570 -9596 43586
rect -9538 43620 -9438 43658
rect -9538 43586 -9522 43620
rect -9454 43586 -9438 43620
rect -9538 43570 -9438 43586
rect -9380 43620 -9280 43658
rect -9380 43586 -9364 43620
rect -9296 43586 -9280 43620
rect -9380 43570 -9280 43586
rect -9222 43620 -9122 43658
rect -9222 43586 -9206 43620
rect -9138 43586 -9122 43620
rect -9222 43570 -9122 43586
rect -9064 43620 -8964 43658
rect -9064 43586 -9048 43620
rect -8980 43586 -8964 43620
rect -9064 43570 -8964 43586
rect -8906 43620 -8806 43658
rect -8906 43586 -8890 43620
rect -8822 43586 -8806 43620
rect -8906 43570 -8806 43586
rect -8748 43620 -8648 43658
rect -8748 43586 -8732 43620
rect -8664 43586 -8648 43620
rect -8748 43570 -8648 43586
rect -8590 43620 -8490 43658
rect -8590 43586 -8574 43620
rect -8506 43586 -8490 43620
rect -8590 43570 -8490 43586
rect -6872 49730 -6772 49746
rect -6872 49696 -6856 49730
rect -6788 49696 -6772 49730
rect -6872 49658 -6772 49696
rect -6714 49730 -6614 49746
rect -6714 49696 -6698 49730
rect -6630 49696 -6614 49730
rect -6714 49658 -6614 49696
rect -6556 49730 -6456 49746
rect -6556 49696 -6540 49730
rect -6472 49696 -6456 49730
rect -6556 49658 -6456 49696
rect -6398 49730 -6298 49746
rect -6398 49696 -6382 49730
rect -6314 49696 -6298 49730
rect -6398 49658 -6298 49696
rect -6240 49730 -6140 49746
rect -6240 49696 -6224 49730
rect -6156 49696 -6140 49730
rect -6240 49658 -6140 49696
rect -6082 49730 -5982 49746
rect -6082 49696 -6066 49730
rect -5998 49696 -5982 49730
rect -6082 49658 -5982 49696
rect -5924 49730 -5824 49746
rect -5924 49696 -5908 49730
rect -5840 49696 -5824 49730
rect -5924 49658 -5824 49696
rect -5766 49730 -5666 49746
rect -5766 49696 -5750 49730
rect -5682 49696 -5666 49730
rect -5766 49658 -5666 49696
rect -5608 49730 -5508 49746
rect -5608 49696 -5592 49730
rect -5524 49696 -5508 49730
rect -5608 49658 -5508 49696
rect -5450 49730 -5350 49746
rect -5450 49696 -5434 49730
rect -5366 49696 -5350 49730
rect -5450 49658 -5350 49696
rect -5292 49730 -5192 49746
rect -5292 49696 -5276 49730
rect -5208 49696 -5192 49730
rect -5292 49658 -5192 49696
rect -5134 49730 -5034 49746
rect -5134 49696 -5118 49730
rect -5050 49696 -5034 49730
rect -5134 49658 -5034 49696
rect -4976 49730 -4876 49746
rect -4976 49696 -4960 49730
rect -4892 49696 -4876 49730
rect -4976 49658 -4876 49696
rect -4818 49730 -4718 49746
rect -4818 49696 -4802 49730
rect -4734 49696 -4718 49730
rect -4818 49658 -4718 49696
rect -4660 49730 -4560 49746
rect -4660 49696 -4644 49730
rect -4576 49696 -4560 49730
rect -4660 49658 -4560 49696
rect -4502 49730 -4402 49746
rect -4502 49696 -4486 49730
rect -4418 49696 -4402 49730
rect -4502 49658 -4402 49696
rect -4344 49730 -4244 49746
rect -4344 49696 -4328 49730
rect -4260 49696 -4244 49730
rect -4344 49658 -4244 49696
rect -4186 49730 -4086 49746
rect -4186 49696 -4170 49730
rect -4102 49696 -4086 49730
rect -4186 49658 -4086 49696
rect -4028 49730 -3928 49746
rect -4028 49696 -4012 49730
rect -3944 49696 -3928 49730
rect -4028 49658 -3928 49696
rect -3870 49730 -3770 49746
rect -3870 49696 -3854 49730
rect -3786 49696 -3770 49730
rect -3870 49658 -3770 49696
rect -3712 49730 -3612 49746
rect -3712 49696 -3696 49730
rect -3628 49696 -3612 49730
rect -3712 49658 -3612 49696
rect -3554 49730 -3454 49746
rect -3554 49696 -3538 49730
rect -3470 49696 -3454 49730
rect -3554 49658 -3454 49696
rect -3396 49730 -3296 49746
rect -3396 49696 -3380 49730
rect -3312 49696 -3296 49730
rect -3396 49658 -3296 49696
rect -3238 49730 -3138 49746
rect -3238 49696 -3222 49730
rect -3154 49696 -3138 49730
rect -3238 49658 -3138 49696
rect -3080 49730 -2980 49746
rect -3080 49696 -3064 49730
rect -2996 49696 -2980 49730
rect -3080 49658 -2980 49696
rect -2922 49730 -2822 49746
rect -2922 49696 -2906 49730
rect -2838 49696 -2822 49730
rect -2922 49658 -2822 49696
rect -2764 49730 -2664 49746
rect -2764 49696 -2748 49730
rect -2680 49696 -2664 49730
rect -2764 49658 -2664 49696
rect -2606 49730 -2506 49746
rect -2606 49696 -2590 49730
rect -2522 49696 -2506 49730
rect -2606 49658 -2506 49696
rect -2448 49730 -2348 49746
rect -2448 49696 -2432 49730
rect -2364 49696 -2348 49730
rect -2448 49658 -2348 49696
rect -2290 49730 -2190 49746
rect -2290 49696 -2274 49730
rect -2206 49696 -2190 49730
rect -2290 49658 -2190 49696
rect -6872 43620 -6772 43658
rect -6872 43586 -6856 43620
rect -6788 43586 -6772 43620
rect -6872 43570 -6772 43586
rect -6714 43620 -6614 43658
rect -6714 43586 -6698 43620
rect -6630 43586 -6614 43620
rect -6714 43570 -6614 43586
rect -6556 43620 -6456 43658
rect -6556 43586 -6540 43620
rect -6472 43586 -6456 43620
rect -6556 43570 -6456 43586
rect -6398 43620 -6298 43658
rect -6398 43586 -6382 43620
rect -6314 43586 -6298 43620
rect -6398 43570 -6298 43586
rect -6240 43620 -6140 43658
rect -6240 43586 -6224 43620
rect -6156 43586 -6140 43620
rect -6240 43570 -6140 43586
rect -6082 43620 -5982 43658
rect -6082 43586 -6066 43620
rect -5998 43586 -5982 43620
rect -6082 43570 -5982 43586
rect -5924 43620 -5824 43658
rect -5924 43586 -5908 43620
rect -5840 43586 -5824 43620
rect -5924 43570 -5824 43586
rect -5766 43620 -5666 43658
rect -5766 43586 -5750 43620
rect -5682 43586 -5666 43620
rect -5766 43570 -5666 43586
rect -5608 43620 -5508 43658
rect -5608 43586 -5592 43620
rect -5524 43586 -5508 43620
rect -5608 43570 -5508 43586
rect -5450 43620 -5350 43658
rect -5450 43586 -5434 43620
rect -5366 43586 -5350 43620
rect -5450 43570 -5350 43586
rect -5292 43620 -5192 43658
rect -5292 43586 -5276 43620
rect -5208 43586 -5192 43620
rect -5292 43570 -5192 43586
rect -5134 43620 -5034 43658
rect -5134 43586 -5118 43620
rect -5050 43586 -5034 43620
rect -5134 43570 -5034 43586
rect -4976 43620 -4876 43658
rect -4976 43586 -4960 43620
rect -4892 43586 -4876 43620
rect -4976 43570 -4876 43586
rect -4818 43620 -4718 43658
rect -4818 43586 -4802 43620
rect -4734 43586 -4718 43620
rect -4818 43570 -4718 43586
rect -4660 43620 -4560 43658
rect -4660 43586 -4644 43620
rect -4576 43586 -4560 43620
rect -4660 43570 -4560 43586
rect -4502 43620 -4402 43658
rect -4502 43586 -4486 43620
rect -4418 43586 -4402 43620
rect -4502 43570 -4402 43586
rect -4344 43620 -4244 43658
rect -4344 43586 -4328 43620
rect -4260 43586 -4244 43620
rect -4344 43570 -4244 43586
rect -4186 43620 -4086 43658
rect -4186 43586 -4170 43620
rect -4102 43586 -4086 43620
rect -4186 43570 -4086 43586
rect -4028 43620 -3928 43658
rect -4028 43586 -4012 43620
rect -3944 43586 -3928 43620
rect -4028 43570 -3928 43586
rect -3870 43620 -3770 43658
rect -3870 43586 -3854 43620
rect -3786 43586 -3770 43620
rect -3870 43570 -3770 43586
rect -3712 43620 -3612 43658
rect -3712 43586 -3696 43620
rect -3628 43586 -3612 43620
rect -3712 43570 -3612 43586
rect -3554 43620 -3454 43658
rect -3554 43586 -3538 43620
rect -3470 43586 -3454 43620
rect -3554 43570 -3454 43586
rect -3396 43620 -3296 43658
rect -3396 43586 -3380 43620
rect -3312 43586 -3296 43620
rect -3396 43570 -3296 43586
rect -3238 43620 -3138 43658
rect -3238 43586 -3222 43620
rect -3154 43586 -3138 43620
rect -3238 43570 -3138 43586
rect -3080 43620 -2980 43658
rect -3080 43586 -3064 43620
rect -2996 43586 -2980 43620
rect -3080 43570 -2980 43586
rect -2922 43620 -2822 43658
rect -2922 43586 -2906 43620
rect -2838 43586 -2822 43620
rect -2922 43570 -2822 43586
rect -2764 43620 -2664 43658
rect -2764 43586 -2748 43620
rect -2680 43586 -2664 43620
rect -2764 43570 -2664 43586
rect -2606 43620 -2506 43658
rect -2606 43586 -2590 43620
rect -2522 43586 -2506 43620
rect -2606 43570 -2506 43586
rect -2448 43620 -2348 43658
rect -2448 43586 -2432 43620
rect -2364 43586 -2348 43620
rect -2448 43570 -2348 43586
rect -2290 43620 -2190 43658
rect -2290 43586 -2274 43620
rect -2206 43586 -2190 43620
rect -2290 43570 -2190 43586
rect -572 49730 -472 49746
rect -572 49696 -556 49730
rect -488 49696 -472 49730
rect -572 49658 -472 49696
rect -414 49730 -314 49746
rect -414 49696 -398 49730
rect -330 49696 -314 49730
rect -414 49658 -314 49696
rect -256 49730 -156 49746
rect -256 49696 -240 49730
rect -172 49696 -156 49730
rect -256 49658 -156 49696
rect -98 49730 2 49746
rect -98 49696 -82 49730
rect -14 49696 2 49730
rect -98 49658 2 49696
rect 60 49730 160 49746
rect 60 49696 76 49730
rect 144 49696 160 49730
rect 60 49658 160 49696
rect 218 49730 318 49746
rect 218 49696 234 49730
rect 302 49696 318 49730
rect 218 49658 318 49696
rect 376 49730 476 49746
rect 376 49696 392 49730
rect 460 49696 476 49730
rect 376 49658 476 49696
rect 534 49730 634 49746
rect 534 49696 550 49730
rect 618 49696 634 49730
rect 534 49658 634 49696
rect 692 49730 792 49746
rect 692 49696 708 49730
rect 776 49696 792 49730
rect 692 49658 792 49696
rect 850 49730 950 49746
rect 850 49696 866 49730
rect 934 49696 950 49730
rect 850 49658 950 49696
rect 1008 49730 1108 49746
rect 1008 49696 1024 49730
rect 1092 49696 1108 49730
rect 1008 49658 1108 49696
rect 1166 49730 1266 49746
rect 1166 49696 1182 49730
rect 1250 49696 1266 49730
rect 1166 49658 1266 49696
rect 1324 49730 1424 49746
rect 1324 49696 1340 49730
rect 1408 49696 1424 49730
rect 1324 49658 1424 49696
rect 1482 49730 1582 49746
rect 1482 49696 1498 49730
rect 1566 49696 1582 49730
rect 1482 49658 1582 49696
rect 1640 49730 1740 49746
rect 1640 49696 1656 49730
rect 1724 49696 1740 49730
rect 1640 49658 1740 49696
rect 1798 49730 1898 49746
rect 1798 49696 1814 49730
rect 1882 49696 1898 49730
rect 1798 49658 1898 49696
rect 1956 49730 2056 49746
rect 1956 49696 1972 49730
rect 2040 49696 2056 49730
rect 1956 49658 2056 49696
rect 2114 49730 2214 49746
rect 2114 49696 2130 49730
rect 2198 49696 2214 49730
rect 2114 49658 2214 49696
rect 2272 49730 2372 49746
rect 2272 49696 2288 49730
rect 2356 49696 2372 49730
rect 2272 49658 2372 49696
rect 2430 49730 2530 49746
rect 2430 49696 2446 49730
rect 2514 49696 2530 49730
rect 2430 49658 2530 49696
rect 2588 49730 2688 49746
rect 2588 49696 2604 49730
rect 2672 49696 2688 49730
rect 2588 49658 2688 49696
rect 2746 49730 2846 49746
rect 2746 49696 2762 49730
rect 2830 49696 2846 49730
rect 2746 49658 2846 49696
rect 2904 49730 3004 49746
rect 2904 49696 2920 49730
rect 2988 49696 3004 49730
rect 2904 49658 3004 49696
rect 3062 49730 3162 49746
rect 3062 49696 3078 49730
rect 3146 49696 3162 49730
rect 3062 49658 3162 49696
rect 3220 49730 3320 49746
rect 3220 49696 3236 49730
rect 3304 49696 3320 49730
rect 3220 49658 3320 49696
rect 3378 49730 3478 49746
rect 3378 49696 3394 49730
rect 3462 49696 3478 49730
rect 3378 49658 3478 49696
rect 3536 49730 3636 49746
rect 3536 49696 3552 49730
rect 3620 49696 3636 49730
rect 3536 49658 3636 49696
rect 3694 49730 3794 49746
rect 3694 49696 3710 49730
rect 3778 49696 3794 49730
rect 3694 49658 3794 49696
rect 3852 49730 3952 49746
rect 3852 49696 3868 49730
rect 3936 49696 3952 49730
rect 3852 49658 3952 49696
rect 4010 49730 4110 49746
rect 4010 49696 4026 49730
rect 4094 49696 4110 49730
rect 4010 49658 4110 49696
rect -572 43620 -472 43658
rect -572 43586 -556 43620
rect -488 43586 -472 43620
rect -572 43570 -472 43586
rect -414 43620 -314 43658
rect -414 43586 -398 43620
rect -330 43586 -314 43620
rect -414 43570 -314 43586
rect -256 43620 -156 43658
rect -256 43586 -240 43620
rect -172 43586 -156 43620
rect -256 43570 -156 43586
rect -98 43620 2 43658
rect -98 43586 -82 43620
rect -14 43586 2 43620
rect -98 43570 2 43586
rect 60 43620 160 43658
rect 60 43586 76 43620
rect 144 43586 160 43620
rect 60 43570 160 43586
rect 218 43620 318 43658
rect 218 43586 234 43620
rect 302 43586 318 43620
rect 218 43570 318 43586
rect 376 43620 476 43658
rect 376 43586 392 43620
rect 460 43586 476 43620
rect 376 43570 476 43586
rect 534 43620 634 43658
rect 534 43586 550 43620
rect 618 43586 634 43620
rect 534 43570 634 43586
rect 692 43620 792 43658
rect 692 43586 708 43620
rect 776 43586 792 43620
rect 692 43570 792 43586
rect 850 43620 950 43658
rect 850 43586 866 43620
rect 934 43586 950 43620
rect 850 43570 950 43586
rect 1008 43620 1108 43658
rect 1008 43586 1024 43620
rect 1092 43586 1108 43620
rect 1008 43570 1108 43586
rect 1166 43620 1266 43658
rect 1166 43586 1182 43620
rect 1250 43586 1266 43620
rect 1166 43570 1266 43586
rect 1324 43620 1424 43658
rect 1324 43586 1340 43620
rect 1408 43586 1424 43620
rect 1324 43570 1424 43586
rect 1482 43620 1582 43658
rect 1482 43586 1498 43620
rect 1566 43586 1582 43620
rect 1482 43570 1582 43586
rect 1640 43620 1740 43658
rect 1640 43586 1656 43620
rect 1724 43586 1740 43620
rect 1640 43570 1740 43586
rect 1798 43620 1898 43658
rect 1798 43586 1814 43620
rect 1882 43586 1898 43620
rect 1798 43570 1898 43586
rect 1956 43620 2056 43658
rect 1956 43586 1972 43620
rect 2040 43586 2056 43620
rect 1956 43570 2056 43586
rect 2114 43620 2214 43658
rect 2114 43586 2130 43620
rect 2198 43586 2214 43620
rect 2114 43570 2214 43586
rect 2272 43620 2372 43658
rect 2272 43586 2288 43620
rect 2356 43586 2372 43620
rect 2272 43570 2372 43586
rect 2430 43620 2530 43658
rect 2430 43586 2446 43620
rect 2514 43586 2530 43620
rect 2430 43570 2530 43586
rect 2588 43620 2688 43658
rect 2588 43586 2604 43620
rect 2672 43586 2688 43620
rect 2588 43570 2688 43586
rect 2746 43620 2846 43658
rect 2746 43586 2762 43620
rect 2830 43586 2846 43620
rect 2746 43570 2846 43586
rect 2904 43620 3004 43658
rect 2904 43586 2920 43620
rect 2988 43586 3004 43620
rect 2904 43570 3004 43586
rect 3062 43620 3162 43658
rect 3062 43586 3078 43620
rect 3146 43586 3162 43620
rect 3062 43570 3162 43586
rect 3220 43620 3320 43658
rect 3220 43586 3236 43620
rect 3304 43586 3320 43620
rect 3220 43570 3320 43586
rect 3378 43620 3478 43658
rect 3378 43586 3394 43620
rect 3462 43586 3478 43620
rect 3378 43570 3478 43586
rect 3536 43620 3636 43658
rect 3536 43586 3552 43620
rect 3620 43586 3636 43620
rect 3536 43570 3636 43586
rect 3694 43620 3794 43658
rect 3694 43586 3710 43620
rect 3778 43586 3794 43620
rect 3694 43570 3794 43586
rect 3852 43620 3952 43658
rect 3852 43586 3868 43620
rect 3936 43586 3952 43620
rect 3852 43570 3952 43586
rect 4010 43620 4110 43658
rect 4010 43586 4026 43620
rect 4094 43586 4110 43620
rect 4010 43570 4110 43586
rect 5728 49730 5828 49746
rect 5728 49696 5744 49730
rect 5812 49696 5828 49730
rect 5728 49658 5828 49696
rect 5886 49730 5986 49746
rect 5886 49696 5902 49730
rect 5970 49696 5986 49730
rect 5886 49658 5986 49696
rect 6044 49730 6144 49746
rect 6044 49696 6060 49730
rect 6128 49696 6144 49730
rect 6044 49658 6144 49696
rect 6202 49730 6302 49746
rect 6202 49696 6218 49730
rect 6286 49696 6302 49730
rect 6202 49658 6302 49696
rect 6360 49730 6460 49746
rect 6360 49696 6376 49730
rect 6444 49696 6460 49730
rect 6360 49658 6460 49696
rect 6518 49730 6618 49746
rect 6518 49696 6534 49730
rect 6602 49696 6618 49730
rect 6518 49658 6618 49696
rect 6676 49730 6776 49746
rect 6676 49696 6692 49730
rect 6760 49696 6776 49730
rect 6676 49658 6776 49696
rect 6834 49730 6934 49746
rect 6834 49696 6850 49730
rect 6918 49696 6934 49730
rect 6834 49658 6934 49696
rect 6992 49730 7092 49746
rect 6992 49696 7008 49730
rect 7076 49696 7092 49730
rect 6992 49658 7092 49696
rect 7150 49730 7250 49746
rect 7150 49696 7166 49730
rect 7234 49696 7250 49730
rect 7150 49658 7250 49696
rect 7308 49730 7408 49746
rect 7308 49696 7324 49730
rect 7392 49696 7408 49730
rect 7308 49658 7408 49696
rect 7466 49730 7566 49746
rect 7466 49696 7482 49730
rect 7550 49696 7566 49730
rect 7466 49658 7566 49696
rect 7624 49730 7724 49746
rect 7624 49696 7640 49730
rect 7708 49696 7724 49730
rect 7624 49658 7724 49696
rect 7782 49730 7882 49746
rect 7782 49696 7798 49730
rect 7866 49696 7882 49730
rect 7782 49658 7882 49696
rect 7940 49730 8040 49746
rect 7940 49696 7956 49730
rect 8024 49696 8040 49730
rect 7940 49658 8040 49696
rect 8098 49730 8198 49746
rect 8098 49696 8114 49730
rect 8182 49696 8198 49730
rect 8098 49658 8198 49696
rect 8256 49730 8356 49746
rect 8256 49696 8272 49730
rect 8340 49696 8356 49730
rect 8256 49658 8356 49696
rect 8414 49730 8514 49746
rect 8414 49696 8430 49730
rect 8498 49696 8514 49730
rect 8414 49658 8514 49696
rect 8572 49730 8672 49746
rect 8572 49696 8588 49730
rect 8656 49696 8672 49730
rect 8572 49658 8672 49696
rect 8730 49730 8830 49746
rect 8730 49696 8746 49730
rect 8814 49696 8830 49730
rect 8730 49658 8830 49696
rect 8888 49730 8988 49746
rect 8888 49696 8904 49730
rect 8972 49696 8988 49730
rect 8888 49658 8988 49696
rect 9046 49730 9146 49746
rect 9046 49696 9062 49730
rect 9130 49696 9146 49730
rect 9046 49658 9146 49696
rect 9204 49730 9304 49746
rect 9204 49696 9220 49730
rect 9288 49696 9304 49730
rect 9204 49658 9304 49696
rect 9362 49730 9462 49746
rect 9362 49696 9378 49730
rect 9446 49696 9462 49730
rect 9362 49658 9462 49696
rect 9520 49730 9620 49746
rect 9520 49696 9536 49730
rect 9604 49696 9620 49730
rect 9520 49658 9620 49696
rect 9678 49730 9778 49746
rect 9678 49696 9694 49730
rect 9762 49696 9778 49730
rect 9678 49658 9778 49696
rect 9836 49730 9936 49746
rect 9836 49696 9852 49730
rect 9920 49696 9936 49730
rect 9836 49658 9936 49696
rect 9994 49730 10094 49746
rect 9994 49696 10010 49730
rect 10078 49696 10094 49730
rect 9994 49658 10094 49696
rect 10152 49730 10252 49746
rect 10152 49696 10168 49730
rect 10236 49696 10252 49730
rect 10152 49658 10252 49696
rect 10310 49730 10410 49746
rect 10310 49696 10326 49730
rect 10394 49696 10410 49730
rect 10310 49658 10410 49696
rect 5728 43620 5828 43658
rect 5728 43586 5744 43620
rect 5812 43586 5828 43620
rect 5728 43570 5828 43586
rect 5886 43620 5986 43658
rect 5886 43586 5902 43620
rect 5970 43586 5986 43620
rect 5886 43570 5986 43586
rect 6044 43620 6144 43658
rect 6044 43586 6060 43620
rect 6128 43586 6144 43620
rect 6044 43570 6144 43586
rect 6202 43620 6302 43658
rect 6202 43586 6218 43620
rect 6286 43586 6302 43620
rect 6202 43570 6302 43586
rect 6360 43620 6460 43658
rect 6360 43586 6376 43620
rect 6444 43586 6460 43620
rect 6360 43570 6460 43586
rect 6518 43620 6618 43658
rect 6518 43586 6534 43620
rect 6602 43586 6618 43620
rect 6518 43570 6618 43586
rect 6676 43620 6776 43658
rect 6676 43586 6692 43620
rect 6760 43586 6776 43620
rect 6676 43570 6776 43586
rect 6834 43620 6934 43658
rect 6834 43586 6850 43620
rect 6918 43586 6934 43620
rect 6834 43570 6934 43586
rect 6992 43620 7092 43658
rect 6992 43586 7008 43620
rect 7076 43586 7092 43620
rect 6992 43570 7092 43586
rect 7150 43620 7250 43658
rect 7150 43586 7166 43620
rect 7234 43586 7250 43620
rect 7150 43570 7250 43586
rect 7308 43620 7408 43658
rect 7308 43586 7324 43620
rect 7392 43586 7408 43620
rect 7308 43570 7408 43586
rect 7466 43620 7566 43658
rect 7466 43586 7482 43620
rect 7550 43586 7566 43620
rect 7466 43570 7566 43586
rect 7624 43620 7724 43658
rect 7624 43586 7640 43620
rect 7708 43586 7724 43620
rect 7624 43570 7724 43586
rect 7782 43620 7882 43658
rect 7782 43586 7798 43620
rect 7866 43586 7882 43620
rect 7782 43570 7882 43586
rect 7940 43620 8040 43658
rect 7940 43586 7956 43620
rect 8024 43586 8040 43620
rect 7940 43570 8040 43586
rect 8098 43620 8198 43658
rect 8098 43586 8114 43620
rect 8182 43586 8198 43620
rect 8098 43570 8198 43586
rect 8256 43620 8356 43658
rect 8256 43586 8272 43620
rect 8340 43586 8356 43620
rect 8256 43570 8356 43586
rect 8414 43620 8514 43658
rect 8414 43586 8430 43620
rect 8498 43586 8514 43620
rect 8414 43570 8514 43586
rect 8572 43620 8672 43658
rect 8572 43586 8588 43620
rect 8656 43586 8672 43620
rect 8572 43570 8672 43586
rect 8730 43620 8830 43658
rect 8730 43586 8746 43620
rect 8814 43586 8830 43620
rect 8730 43570 8830 43586
rect 8888 43620 8988 43658
rect 8888 43586 8904 43620
rect 8972 43586 8988 43620
rect 8888 43570 8988 43586
rect 9046 43620 9146 43658
rect 9046 43586 9062 43620
rect 9130 43586 9146 43620
rect 9046 43570 9146 43586
rect 9204 43620 9304 43658
rect 9204 43586 9220 43620
rect 9288 43586 9304 43620
rect 9204 43570 9304 43586
rect 9362 43620 9462 43658
rect 9362 43586 9378 43620
rect 9446 43586 9462 43620
rect 9362 43570 9462 43586
rect 9520 43620 9620 43658
rect 9520 43586 9536 43620
rect 9604 43586 9620 43620
rect 9520 43570 9620 43586
rect 9678 43620 9778 43658
rect 9678 43586 9694 43620
rect 9762 43586 9778 43620
rect 9678 43570 9778 43586
rect 9836 43620 9936 43658
rect 9836 43586 9852 43620
rect 9920 43586 9936 43620
rect 9836 43570 9936 43586
rect 9994 43620 10094 43658
rect 9994 43586 10010 43620
rect 10078 43586 10094 43620
rect 9994 43570 10094 43586
rect 10152 43620 10252 43658
rect 10152 43586 10168 43620
rect 10236 43586 10252 43620
rect 10152 43570 10252 43586
rect 10310 43620 10410 43658
rect 10310 43586 10326 43620
rect 10394 43586 10410 43620
rect 10310 43570 10410 43586
rect -13172 42730 -13072 42746
rect -13172 42696 -13156 42730
rect -13088 42696 -13072 42730
rect -13172 42658 -13072 42696
rect -13014 42730 -12914 42746
rect -13014 42696 -12998 42730
rect -12930 42696 -12914 42730
rect -13014 42658 -12914 42696
rect -12856 42730 -12756 42746
rect -12856 42696 -12840 42730
rect -12772 42696 -12756 42730
rect -12856 42658 -12756 42696
rect -12698 42730 -12598 42746
rect -12698 42696 -12682 42730
rect -12614 42696 -12598 42730
rect -12698 42658 -12598 42696
rect -12540 42730 -12440 42746
rect -12540 42696 -12524 42730
rect -12456 42696 -12440 42730
rect -12540 42658 -12440 42696
rect -12382 42730 -12282 42746
rect -12382 42696 -12366 42730
rect -12298 42696 -12282 42730
rect -12382 42658 -12282 42696
rect -12224 42730 -12124 42746
rect -12224 42696 -12208 42730
rect -12140 42696 -12124 42730
rect -12224 42658 -12124 42696
rect -12066 42730 -11966 42746
rect -12066 42696 -12050 42730
rect -11982 42696 -11966 42730
rect -12066 42658 -11966 42696
rect -11908 42730 -11808 42746
rect -11908 42696 -11892 42730
rect -11824 42696 -11808 42730
rect -11908 42658 -11808 42696
rect -11750 42730 -11650 42746
rect -11750 42696 -11734 42730
rect -11666 42696 -11650 42730
rect -11750 42658 -11650 42696
rect -11592 42730 -11492 42746
rect -11592 42696 -11576 42730
rect -11508 42696 -11492 42730
rect -11592 42658 -11492 42696
rect -11434 42730 -11334 42746
rect -11434 42696 -11418 42730
rect -11350 42696 -11334 42730
rect -11434 42658 -11334 42696
rect -11276 42730 -11176 42746
rect -11276 42696 -11260 42730
rect -11192 42696 -11176 42730
rect -11276 42658 -11176 42696
rect -11118 42730 -11018 42746
rect -11118 42696 -11102 42730
rect -11034 42696 -11018 42730
rect -11118 42658 -11018 42696
rect -10960 42730 -10860 42746
rect -10960 42696 -10944 42730
rect -10876 42696 -10860 42730
rect -10960 42658 -10860 42696
rect -10802 42730 -10702 42746
rect -10802 42696 -10786 42730
rect -10718 42696 -10702 42730
rect -10802 42658 -10702 42696
rect -10644 42730 -10544 42746
rect -10644 42696 -10628 42730
rect -10560 42696 -10544 42730
rect -10644 42658 -10544 42696
rect -10486 42730 -10386 42746
rect -10486 42696 -10470 42730
rect -10402 42696 -10386 42730
rect -10486 42658 -10386 42696
rect -10328 42730 -10228 42746
rect -10328 42696 -10312 42730
rect -10244 42696 -10228 42730
rect -10328 42658 -10228 42696
rect -10170 42730 -10070 42746
rect -10170 42696 -10154 42730
rect -10086 42696 -10070 42730
rect -10170 42658 -10070 42696
rect -10012 42730 -9912 42746
rect -10012 42696 -9996 42730
rect -9928 42696 -9912 42730
rect -10012 42658 -9912 42696
rect -9854 42730 -9754 42746
rect -9854 42696 -9838 42730
rect -9770 42696 -9754 42730
rect -9854 42658 -9754 42696
rect -9696 42730 -9596 42746
rect -9696 42696 -9680 42730
rect -9612 42696 -9596 42730
rect -9696 42658 -9596 42696
rect -9538 42730 -9438 42746
rect -9538 42696 -9522 42730
rect -9454 42696 -9438 42730
rect -9538 42658 -9438 42696
rect -9380 42730 -9280 42746
rect -9380 42696 -9364 42730
rect -9296 42696 -9280 42730
rect -9380 42658 -9280 42696
rect -9222 42730 -9122 42746
rect -9222 42696 -9206 42730
rect -9138 42696 -9122 42730
rect -9222 42658 -9122 42696
rect -9064 42730 -8964 42746
rect -9064 42696 -9048 42730
rect -8980 42696 -8964 42730
rect -9064 42658 -8964 42696
rect -8906 42730 -8806 42746
rect -8906 42696 -8890 42730
rect -8822 42696 -8806 42730
rect -8906 42658 -8806 42696
rect -8748 42730 -8648 42746
rect -8748 42696 -8732 42730
rect -8664 42696 -8648 42730
rect -8748 42658 -8648 42696
rect -8590 42730 -8490 42746
rect -8590 42696 -8574 42730
rect -8506 42696 -8490 42730
rect -8590 42658 -8490 42696
rect -13172 36620 -13072 36658
rect -13172 36586 -13156 36620
rect -13088 36586 -13072 36620
rect -13172 36570 -13072 36586
rect -13014 36620 -12914 36658
rect -13014 36586 -12998 36620
rect -12930 36586 -12914 36620
rect -13014 36570 -12914 36586
rect -12856 36620 -12756 36658
rect -12856 36586 -12840 36620
rect -12772 36586 -12756 36620
rect -12856 36570 -12756 36586
rect -12698 36620 -12598 36658
rect -12698 36586 -12682 36620
rect -12614 36586 -12598 36620
rect -12698 36570 -12598 36586
rect -12540 36620 -12440 36658
rect -12540 36586 -12524 36620
rect -12456 36586 -12440 36620
rect -12540 36570 -12440 36586
rect -12382 36620 -12282 36658
rect -12382 36586 -12366 36620
rect -12298 36586 -12282 36620
rect -12382 36570 -12282 36586
rect -12224 36620 -12124 36658
rect -12224 36586 -12208 36620
rect -12140 36586 -12124 36620
rect -12224 36570 -12124 36586
rect -12066 36620 -11966 36658
rect -12066 36586 -12050 36620
rect -11982 36586 -11966 36620
rect -12066 36570 -11966 36586
rect -11908 36620 -11808 36658
rect -11908 36586 -11892 36620
rect -11824 36586 -11808 36620
rect -11908 36570 -11808 36586
rect -11750 36620 -11650 36658
rect -11750 36586 -11734 36620
rect -11666 36586 -11650 36620
rect -11750 36570 -11650 36586
rect -11592 36620 -11492 36658
rect -11592 36586 -11576 36620
rect -11508 36586 -11492 36620
rect -11592 36570 -11492 36586
rect -11434 36620 -11334 36658
rect -11434 36586 -11418 36620
rect -11350 36586 -11334 36620
rect -11434 36570 -11334 36586
rect -11276 36620 -11176 36658
rect -11276 36586 -11260 36620
rect -11192 36586 -11176 36620
rect -11276 36570 -11176 36586
rect -11118 36620 -11018 36658
rect -11118 36586 -11102 36620
rect -11034 36586 -11018 36620
rect -11118 36570 -11018 36586
rect -10960 36620 -10860 36658
rect -10960 36586 -10944 36620
rect -10876 36586 -10860 36620
rect -10960 36570 -10860 36586
rect -10802 36620 -10702 36658
rect -10802 36586 -10786 36620
rect -10718 36586 -10702 36620
rect -10802 36570 -10702 36586
rect -10644 36620 -10544 36658
rect -10644 36586 -10628 36620
rect -10560 36586 -10544 36620
rect -10644 36570 -10544 36586
rect -10486 36620 -10386 36658
rect -10486 36586 -10470 36620
rect -10402 36586 -10386 36620
rect -10486 36570 -10386 36586
rect -10328 36620 -10228 36658
rect -10328 36586 -10312 36620
rect -10244 36586 -10228 36620
rect -10328 36570 -10228 36586
rect -10170 36620 -10070 36658
rect -10170 36586 -10154 36620
rect -10086 36586 -10070 36620
rect -10170 36570 -10070 36586
rect -10012 36620 -9912 36658
rect -10012 36586 -9996 36620
rect -9928 36586 -9912 36620
rect -10012 36570 -9912 36586
rect -9854 36620 -9754 36658
rect -9854 36586 -9838 36620
rect -9770 36586 -9754 36620
rect -9854 36570 -9754 36586
rect -9696 36620 -9596 36658
rect -9696 36586 -9680 36620
rect -9612 36586 -9596 36620
rect -9696 36570 -9596 36586
rect -9538 36620 -9438 36658
rect -9538 36586 -9522 36620
rect -9454 36586 -9438 36620
rect -9538 36570 -9438 36586
rect -9380 36620 -9280 36658
rect -9380 36586 -9364 36620
rect -9296 36586 -9280 36620
rect -9380 36570 -9280 36586
rect -9222 36620 -9122 36658
rect -9222 36586 -9206 36620
rect -9138 36586 -9122 36620
rect -9222 36570 -9122 36586
rect -9064 36620 -8964 36658
rect -9064 36586 -9048 36620
rect -8980 36586 -8964 36620
rect -9064 36570 -8964 36586
rect -8906 36620 -8806 36658
rect -8906 36586 -8890 36620
rect -8822 36586 -8806 36620
rect -8906 36570 -8806 36586
rect -8748 36620 -8648 36658
rect -8748 36586 -8732 36620
rect -8664 36586 -8648 36620
rect -8748 36570 -8648 36586
rect -8590 36620 -8490 36658
rect -8590 36586 -8574 36620
rect -8506 36586 -8490 36620
rect -8590 36570 -8490 36586
rect -6872 42730 -6772 42746
rect -6872 42696 -6856 42730
rect -6788 42696 -6772 42730
rect -6872 42658 -6772 42696
rect -6714 42730 -6614 42746
rect -6714 42696 -6698 42730
rect -6630 42696 -6614 42730
rect -6714 42658 -6614 42696
rect -6556 42730 -6456 42746
rect -6556 42696 -6540 42730
rect -6472 42696 -6456 42730
rect -6556 42658 -6456 42696
rect -6398 42730 -6298 42746
rect -6398 42696 -6382 42730
rect -6314 42696 -6298 42730
rect -6398 42658 -6298 42696
rect -6240 42730 -6140 42746
rect -6240 42696 -6224 42730
rect -6156 42696 -6140 42730
rect -6240 42658 -6140 42696
rect -6082 42730 -5982 42746
rect -6082 42696 -6066 42730
rect -5998 42696 -5982 42730
rect -6082 42658 -5982 42696
rect -5924 42730 -5824 42746
rect -5924 42696 -5908 42730
rect -5840 42696 -5824 42730
rect -5924 42658 -5824 42696
rect -5766 42730 -5666 42746
rect -5766 42696 -5750 42730
rect -5682 42696 -5666 42730
rect -5766 42658 -5666 42696
rect -5608 42730 -5508 42746
rect -5608 42696 -5592 42730
rect -5524 42696 -5508 42730
rect -5608 42658 -5508 42696
rect -5450 42730 -5350 42746
rect -5450 42696 -5434 42730
rect -5366 42696 -5350 42730
rect -5450 42658 -5350 42696
rect -5292 42730 -5192 42746
rect -5292 42696 -5276 42730
rect -5208 42696 -5192 42730
rect -5292 42658 -5192 42696
rect -5134 42730 -5034 42746
rect -5134 42696 -5118 42730
rect -5050 42696 -5034 42730
rect -5134 42658 -5034 42696
rect -4976 42730 -4876 42746
rect -4976 42696 -4960 42730
rect -4892 42696 -4876 42730
rect -4976 42658 -4876 42696
rect -4818 42730 -4718 42746
rect -4818 42696 -4802 42730
rect -4734 42696 -4718 42730
rect -4818 42658 -4718 42696
rect -4660 42730 -4560 42746
rect -4660 42696 -4644 42730
rect -4576 42696 -4560 42730
rect -4660 42658 -4560 42696
rect -4502 42730 -4402 42746
rect -4502 42696 -4486 42730
rect -4418 42696 -4402 42730
rect -4502 42658 -4402 42696
rect -4344 42730 -4244 42746
rect -4344 42696 -4328 42730
rect -4260 42696 -4244 42730
rect -4344 42658 -4244 42696
rect -4186 42730 -4086 42746
rect -4186 42696 -4170 42730
rect -4102 42696 -4086 42730
rect -4186 42658 -4086 42696
rect -4028 42730 -3928 42746
rect -4028 42696 -4012 42730
rect -3944 42696 -3928 42730
rect -4028 42658 -3928 42696
rect -3870 42730 -3770 42746
rect -3870 42696 -3854 42730
rect -3786 42696 -3770 42730
rect -3870 42658 -3770 42696
rect -3712 42730 -3612 42746
rect -3712 42696 -3696 42730
rect -3628 42696 -3612 42730
rect -3712 42658 -3612 42696
rect -3554 42730 -3454 42746
rect -3554 42696 -3538 42730
rect -3470 42696 -3454 42730
rect -3554 42658 -3454 42696
rect -3396 42730 -3296 42746
rect -3396 42696 -3380 42730
rect -3312 42696 -3296 42730
rect -3396 42658 -3296 42696
rect -3238 42730 -3138 42746
rect -3238 42696 -3222 42730
rect -3154 42696 -3138 42730
rect -3238 42658 -3138 42696
rect -3080 42730 -2980 42746
rect -3080 42696 -3064 42730
rect -2996 42696 -2980 42730
rect -3080 42658 -2980 42696
rect -2922 42730 -2822 42746
rect -2922 42696 -2906 42730
rect -2838 42696 -2822 42730
rect -2922 42658 -2822 42696
rect -2764 42730 -2664 42746
rect -2764 42696 -2748 42730
rect -2680 42696 -2664 42730
rect -2764 42658 -2664 42696
rect -2606 42730 -2506 42746
rect -2606 42696 -2590 42730
rect -2522 42696 -2506 42730
rect -2606 42658 -2506 42696
rect -2448 42730 -2348 42746
rect -2448 42696 -2432 42730
rect -2364 42696 -2348 42730
rect -2448 42658 -2348 42696
rect -2290 42730 -2190 42746
rect -2290 42696 -2274 42730
rect -2206 42696 -2190 42730
rect -2290 42658 -2190 42696
rect -6872 36620 -6772 36658
rect -6872 36586 -6856 36620
rect -6788 36586 -6772 36620
rect -6872 36570 -6772 36586
rect -6714 36620 -6614 36658
rect -6714 36586 -6698 36620
rect -6630 36586 -6614 36620
rect -6714 36570 -6614 36586
rect -6556 36620 -6456 36658
rect -6556 36586 -6540 36620
rect -6472 36586 -6456 36620
rect -6556 36570 -6456 36586
rect -6398 36620 -6298 36658
rect -6398 36586 -6382 36620
rect -6314 36586 -6298 36620
rect -6398 36570 -6298 36586
rect -6240 36620 -6140 36658
rect -6240 36586 -6224 36620
rect -6156 36586 -6140 36620
rect -6240 36570 -6140 36586
rect -6082 36620 -5982 36658
rect -6082 36586 -6066 36620
rect -5998 36586 -5982 36620
rect -6082 36570 -5982 36586
rect -5924 36620 -5824 36658
rect -5924 36586 -5908 36620
rect -5840 36586 -5824 36620
rect -5924 36570 -5824 36586
rect -5766 36620 -5666 36658
rect -5766 36586 -5750 36620
rect -5682 36586 -5666 36620
rect -5766 36570 -5666 36586
rect -5608 36620 -5508 36658
rect -5608 36586 -5592 36620
rect -5524 36586 -5508 36620
rect -5608 36570 -5508 36586
rect -5450 36620 -5350 36658
rect -5450 36586 -5434 36620
rect -5366 36586 -5350 36620
rect -5450 36570 -5350 36586
rect -5292 36620 -5192 36658
rect -5292 36586 -5276 36620
rect -5208 36586 -5192 36620
rect -5292 36570 -5192 36586
rect -5134 36620 -5034 36658
rect -5134 36586 -5118 36620
rect -5050 36586 -5034 36620
rect -5134 36570 -5034 36586
rect -4976 36620 -4876 36658
rect -4976 36586 -4960 36620
rect -4892 36586 -4876 36620
rect -4976 36570 -4876 36586
rect -4818 36620 -4718 36658
rect -4818 36586 -4802 36620
rect -4734 36586 -4718 36620
rect -4818 36570 -4718 36586
rect -4660 36620 -4560 36658
rect -4660 36586 -4644 36620
rect -4576 36586 -4560 36620
rect -4660 36570 -4560 36586
rect -4502 36620 -4402 36658
rect -4502 36586 -4486 36620
rect -4418 36586 -4402 36620
rect -4502 36570 -4402 36586
rect -4344 36620 -4244 36658
rect -4344 36586 -4328 36620
rect -4260 36586 -4244 36620
rect -4344 36570 -4244 36586
rect -4186 36620 -4086 36658
rect -4186 36586 -4170 36620
rect -4102 36586 -4086 36620
rect -4186 36570 -4086 36586
rect -4028 36620 -3928 36658
rect -4028 36586 -4012 36620
rect -3944 36586 -3928 36620
rect -4028 36570 -3928 36586
rect -3870 36620 -3770 36658
rect -3870 36586 -3854 36620
rect -3786 36586 -3770 36620
rect -3870 36570 -3770 36586
rect -3712 36620 -3612 36658
rect -3712 36586 -3696 36620
rect -3628 36586 -3612 36620
rect -3712 36570 -3612 36586
rect -3554 36620 -3454 36658
rect -3554 36586 -3538 36620
rect -3470 36586 -3454 36620
rect -3554 36570 -3454 36586
rect -3396 36620 -3296 36658
rect -3396 36586 -3380 36620
rect -3312 36586 -3296 36620
rect -3396 36570 -3296 36586
rect -3238 36620 -3138 36658
rect -3238 36586 -3222 36620
rect -3154 36586 -3138 36620
rect -3238 36570 -3138 36586
rect -3080 36620 -2980 36658
rect -3080 36586 -3064 36620
rect -2996 36586 -2980 36620
rect -3080 36570 -2980 36586
rect -2922 36620 -2822 36658
rect -2922 36586 -2906 36620
rect -2838 36586 -2822 36620
rect -2922 36570 -2822 36586
rect -2764 36620 -2664 36658
rect -2764 36586 -2748 36620
rect -2680 36586 -2664 36620
rect -2764 36570 -2664 36586
rect -2606 36620 -2506 36658
rect -2606 36586 -2590 36620
rect -2522 36586 -2506 36620
rect -2606 36570 -2506 36586
rect -2448 36620 -2348 36658
rect -2448 36586 -2432 36620
rect -2364 36586 -2348 36620
rect -2448 36570 -2348 36586
rect -2290 36620 -2190 36658
rect -2290 36586 -2274 36620
rect -2206 36586 -2190 36620
rect -2290 36570 -2190 36586
rect -572 42730 -472 42746
rect -572 42696 -556 42730
rect -488 42696 -472 42730
rect -572 42658 -472 42696
rect -414 42730 -314 42746
rect -414 42696 -398 42730
rect -330 42696 -314 42730
rect -414 42658 -314 42696
rect -256 42730 -156 42746
rect -256 42696 -240 42730
rect -172 42696 -156 42730
rect -256 42658 -156 42696
rect -98 42730 2 42746
rect -98 42696 -82 42730
rect -14 42696 2 42730
rect -98 42658 2 42696
rect 60 42730 160 42746
rect 60 42696 76 42730
rect 144 42696 160 42730
rect 60 42658 160 42696
rect 218 42730 318 42746
rect 218 42696 234 42730
rect 302 42696 318 42730
rect 218 42658 318 42696
rect 376 42730 476 42746
rect 376 42696 392 42730
rect 460 42696 476 42730
rect 376 42658 476 42696
rect 534 42730 634 42746
rect 534 42696 550 42730
rect 618 42696 634 42730
rect 534 42658 634 42696
rect 692 42730 792 42746
rect 692 42696 708 42730
rect 776 42696 792 42730
rect 692 42658 792 42696
rect 850 42730 950 42746
rect 850 42696 866 42730
rect 934 42696 950 42730
rect 850 42658 950 42696
rect 1008 42730 1108 42746
rect 1008 42696 1024 42730
rect 1092 42696 1108 42730
rect 1008 42658 1108 42696
rect 1166 42730 1266 42746
rect 1166 42696 1182 42730
rect 1250 42696 1266 42730
rect 1166 42658 1266 42696
rect 1324 42730 1424 42746
rect 1324 42696 1340 42730
rect 1408 42696 1424 42730
rect 1324 42658 1424 42696
rect 1482 42730 1582 42746
rect 1482 42696 1498 42730
rect 1566 42696 1582 42730
rect 1482 42658 1582 42696
rect 1640 42730 1740 42746
rect 1640 42696 1656 42730
rect 1724 42696 1740 42730
rect 1640 42658 1740 42696
rect 1798 42730 1898 42746
rect 1798 42696 1814 42730
rect 1882 42696 1898 42730
rect 1798 42658 1898 42696
rect 1956 42730 2056 42746
rect 1956 42696 1972 42730
rect 2040 42696 2056 42730
rect 1956 42658 2056 42696
rect 2114 42730 2214 42746
rect 2114 42696 2130 42730
rect 2198 42696 2214 42730
rect 2114 42658 2214 42696
rect 2272 42730 2372 42746
rect 2272 42696 2288 42730
rect 2356 42696 2372 42730
rect 2272 42658 2372 42696
rect 2430 42730 2530 42746
rect 2430 42696 2446 42730
rect 2514 42696 2530 42730
rect 2430 42658 2530 42696
rect 2588 42730 2688 42746
rect 2588 42696 2604 42730
rect 2672 42696 2688 42730
rect 2588 42658 2688 42696
rect 2746 42730 2846 42746
rect 2746 42696 2762 42730
rect 2830 42696 2846 42730
rect 2746 42658 2846 42696
rect 2904 42730 3004 42746
rect 2904 42696 2920 42730
rect 2988 42696 3004 42730
rect 2904 42658 3004 42696
rect 3062 42730 3162 42746
rect 3062 42696 3078 42730
rect 3146 42696 3162 42730
rect 3062 42658 3162 42696
rect 3220 42730 3320 42746
rect 3220 42696 3236 42730
rect 3304 42696 3320 42730
rect 3220 42658 3320 42696
rect 3378 42730 3478 42746
rect 3378 42696 3394 42730
rect 3462 42696 3478 42730
rect 3378 42658 3478 42696
rect 3536 42730 3636 42746
rect 3536 42696 3552 42730
rect 3620 42696 3636 42730
rect 3536 42658 3636 42696
rect 3694 42730 3794 42746
rect 3694 42696 3710 42730
rect 3778 42696 3794 42730
rect 3694 42658 3794 42696
rect 3852 42730 3952 42746
rect 3852 42696 3868 42730
rect 3936 42696 3952 42730
rect 3852 42658 3952 42696
rect 4010 42730 4110 42746
rect 4010 42696 4026 42730
rect 4094 42696 4110 42730
rect 4010 42658 4110 42696
rect -572 36620 -472 36658
rect -572 36586 -556 36620
rect -488 36586 -472 36620
rect -572 36570 -472 36586
rect -414 36620 -314 36658
rect -414 36586 -398 36620
rect -330 36586 -314 36620
rect -414 36570 -314 36586
rect -256 36620 -156 36658
rect -256 36586 -240 36620
rect -172 36586 -156 36620
rect -256 36570 -156 36586
rect -98 36620 2 36658
rect -98 36586 -82 36620
rect -14 36586 2 36620
rect -98 36570 2 36586
rect 60 36620 160 36658
rect 60 36586 76 36620
rect 144 36586 160 36620
rect 60 36570 160 36586
rect 218 36620 318 36658
rect 218 36586 234 36620
rect 302 36586 318 36620
rect 218 36570 318 36586
rect 376 36620 476 36658
rect 376 36586 392 36620
rect 460 36586 476 36620
rect 376 36570 476 36586
rect 534 36620 634 36658
rect 534 36586 550 36620
rect 618 36586 634 36620
rect 534 36570 634 36586
rect 692 36620 792 36658
rect 692 36586 708 36620
rect 776 36586 792 36620
rect 692 36570 792 36586
rect 850 36620 950 36658
rect 850 36586 866 36620
rect 934 36586 950 36620
rect 850 36570 950 36586
rect 1008 36620 1108 36658
rect 1008 36586 1024 36620
rect 1092 36586 1108 36620
rect 1008 36570 1108 36586
rect 1166 36620 1266 36658
rect 1166 36586 1182 36620
rect 1250 36586 1266 36620
rect 1166 36570 1266 36586
rect 1324 36620 1424 36658
rect 1324 36586 1340 36620
rect 1408 36586 1424 36620
rect 1324 36570 1424 36586
rect 1482 36620 1582 36658
rect 1482 36586 1498 36620
rect 1566 36586 1582 36620
rect 1482 36570 1582 36586
rect 1640 36620 1740 36658
rect 1640 36586 1656 36620
rect 1724 36586 1740 36620
rect 1640 36570 1740 36586
rect 1798 36620 1898 36658
rect 1798 36586 1814 36620
rect 1882 36586 1898 36620
rect 1798 36570 1898 36586
rect 1956 36620 2056 36658
rect 1956 36586 1972 36620
rect 2040 36586 2056 36620
rect 1956 36570 2056 36586
rect 2114 36620 2214 36658
rect 2114 36586 2130 36620
rect 2198 36586 2214 36620
rect 2114 36570 2214 36586
rect 2272 36620 2372 36658
rect 2272 36586 2288 36620
rect 2356 36586 2372 36620
rect 2272 36570 2372 36586
rect 2430 36620 2530 36658
rect 2430 36586 2446 36620
rect 2514 36586 2530 36620
rect 2430 36570 2530 36586
rect 2588 36620 2688 36658
rect 2588 36586 2604 36620
rect 2672 36586 2688 36620
rect 2588 36570 2688 36586
rect 2746 36620 2846 36658
rect 2746 36586 2762 36620
rect 2830 36586 2846 36620
rect 2746 36570 2846 36586
rect 2904 36620 3004 36658
rect 2904 36586 2920 36620
rect 2988 36586 3004 36620
rect 2904 36570 3004 36586
rect 3062 36620 3162 36658
rect 3062 36586 3078 36620
rect 3146 36586 3162 36620
rect 3062 36570 3162 36586
rect 3220 36620 3320 36658
rect 3220 36586 3236 36620
rect 3304 36586 3320 36620
rect 3220 36570 3320 36586
rect 3378 36620 3478 36658
rect 3378 36586 3394 36620
rect 3462 36586 3478 36620
rect 3378 36570 3478 36586
rect 3536 36620 3636 36658
rect 3536 36586 3552 36620
rect 3620 36586 3636 36620
rect 3536 36570 3636 36586
rect 3694 36620 3794 36658
rect 3694 36586 3710 36620
rect 3778 36586 3794 36620
rect 3694 36570 3794 36586
rect 3852 36620 3952 36658
rect 3852 36586 3868 36620
rect 3936 36586 3952 36620
rect 3852 36570 3952 36586
rect 4010 36620 4110 36658
rect 4010 36586 4026 36620
rect 4094 36586 4110 36620
rect 4010 36570 4110 36586
rect 5728 42730 5828 42746
rect 5728 42696 5744 42730
rect 5812 42696 5828 42730
rect 5728 42658 5828 42696
rect 5886 42730 5986 42746
rect 5886 42696 5902 42730
rect 5970 42696 5986 42730
rect 5886 42658 5986 42696
rect 6044 42730 6144 42746
rect 6044 42696 6060 42730
rect 6128 42696 6144 42730
rect 6044 42658 6144 42696
rect 6202 42730 6302 42746
rect 6202 42696 6218 42730
rect 6286 42696 6302 42730
rect 6202 42658 6302 42696
rect 6360 42730 6460 42746
rect 6360 42696 6376 42730
rect 6444 42696 6460 42730
rect 6360 42658 6460 42696
rect 6518 42730 6618 42746
rect 6518 42696 6534 42730
rect 6602 42696 6618 42730
rect 6518 42658 6618 42696
rect 6676 42730 6776 42746
rect 6676 42696 6692 42730
rect 6760 42696 6776 42730
rect 6676 42658 6776 42696
rect 6834 42730 6934 42746
rect 6834 42696 6850 42730
rect 6918 42696 6934 42730
rect 6834 42658 6934 42696
rect 6992 42730 7092 42746
rect 6992 42696 7008 42730
rect 7076 42696 7092 42730
rect 6992 42658 7092 42696
rect 7150 42730 7250 42746
rect 7150 42696 7166 42730
rect 7234 42696 7250 42730
rect 7150 42658 7250 42696
rect 7308 42730 7408 42746
rect 7308 42696 7324 42730
rect 7392 42696 7408 42730
rect 7308 42658 7408 42696
rect 7466 42730 7566 42746
rect 7466 42696 7482 42730
rect 7550 42696 7566 42730
rect 7466 42658 7566 42696
rect 7624 42730 7724 42746
rect 7624 42696 7640 42730
rect 7708 42696 7724 42730
rect 7624 42658 7724 42696
rect 7782 42730 7882 42746
rect 7782 42696 7798 42730
rect 7866 42696 7882 42730
rect 7782 42658 7882 42696
rect 7940 42730 8040 42746
rect 7940 42696 7956 42730
rect 8024 42696 8040 42730
rect 7940 42658 8040 42696
rect 8098 42730 8198 42746
rect 8098 42696 8114 42730
rect 8182 42696 8198 42730
rect 8098 42658 8198 42696
rect 8256 42730 8356 42746
rect 8256 42696 8272 42730
rect 8340 42696 8356 42730
rect 8256 42658 8356 42696
rect 8414 42730 8514 42746
rect 8414 42696 8430 42730
rect 8498 42696 8514 42730
rect 8414 42658 8514 42696
rect 8572 42730 8672 42746
rect 8572 42696 8588 42730
rect 8656 42696 8672 42730
rect 8572 42658 8672 42696
rect 8730 42730 8830 42746
rect 8730 42696 8746 42730
rect 8814 42696 8830 42730
rect 8730 42658 8830 42696
rect 8888 42730 8988 42746
rect 8888 42696 8904 42730
rect 8972 42696 8988 42730
rect 8888 42658 8988 42696
rect 9046 42730 9146 42746
rect 9046 42696 9062 42730
rect 9130 42696 9146 42730
rect 9046 42658 9146 42696
rect 9204 42730 9304 42746
rect 9204 42696 9220 42730
rect 9288 42696 9304 42730
rect 9204 42658 9304 42696
rect 9362 42730 9462 42746
rect 9362 42696 9378 42730
rect 9446 42696 9462 42730
rect 9362 42658 9462 42696
rect 9520 42730 9620 42746
rect 9520 42696 9536 42730
rect 9604 42696 9620 42730
rect 9520 42658 9620 42696
rect 9678 42730 9778 42746
rect 9678 42696 9694 42730
rect 9762 42696 9778 42730
rect 9678 42658 9778 42696
rect 9836 42730 9936 42746
rect 9836 42696 9852 42730
rect 9920 42696 9936 42730
rect 9836 42658 9936 42696
rect 9994 42730 10094 42746
rect 9994 42696 10010 42730
rect 10078 42696 10094 42730
rect 9994 42658 10094 42696
rect 10152 42730 10252 42746
rect 10152 42696 10168 42730
rect 10236 42696 10252 42730
rect 10152 42658 10252 42696
rect 10310 42730 10410 42746
rect 10310 42696 10326 42730
rect 10394 42696 10410 42730
rect 10310 42658 10410 42696
rect 5728 36620 5828 36658
rect 5728 36586 5744 36620
rect 5812 36586 5828 36620
rect 5728 36570 5828 36586
rect 5886 36620 5986 36658
rect 5886 36586 5902 36620
rect 5970 36586 5986 36620
rect 5886 36570 5986 36586
rect 6044 36620 6144 36658
rect 6044 36586 6060 36620
rect 6128 36586 6144 36620
rect 6044 36570 6144 36586
rect 6202 36620 6302 36658
rect 6202 36586 6218 36620
rect 6286 36586 6302 36620
rect 6202 36570 6302 36586
rect 6360 36620 6460 36658
rect 6360 36586 6376 36620
rect 6444 36586 6460 36620
rect 6360 36570 6460 36586
rect 6518 36620 6618 36658
rect 6518 36586 6534 36620
rect 6602 36586 6618 36620
rect 6518 36570 6618 36586
rect 6676 36620 6776 36658
rect 6676 36586 6692 36620
rect 6760 36586 6776 36620
rect 6676 36570 6776 36586
rect 6834 36620 6934 36658
rect 6834 36586 6850 36620
rect 6918 36586 6934 36620
rect 6834 36570 6934 36586
rect 6992 36620 7092 36658
rect 6992 36586 7008 36620
rect 7076 36586 7092 36620
rect 6992 36570 7092 36586
rect 7150 36620 7250 36658
rect 7150 36586 7166 36620
rect 7234 36586 7250 36620
rect 7150 36570 7250 36586
rect 7308 36620 7408 36658
rect 7308 36586 7324 36620
rect 7392 36586 7408 36620
rect 7308 36570 7408 36586
rect 7466 36620 7566 36658
rect 7466 36586 7482 36620
rect 7550 36586 7566 36620
rect 7466 36570 7566 36586
rect 7624 36620 7724 36658
rect 7624 36586 7640 36620
rect 7708 36586 7724 36620
rect 7624 36570 7724 36586
rect 7782 36620 7882 36658
rect 7782 36586 7798 36620
rect 7866 36586 7882 36620
rect 7782 36570 7882 36586
rect 7940 36620 8040 36658
rect 7940 36586 7956 36620
rect 8024 36586 8040 36620
rect 7940 36570 8040 36586
rect 8098 36620 8198 36658
rect 8098 36586 8114 36620
rect 8182 36586 8198 36620
rect 8098 36570 8198 36586
rect 8256 36620 8356 36658
rect 8256 36586 8272 36620
rect 8340 36586 8356 36620
rect 8256 36570 8356 36586
rect 8414 36620 8514 36658
rect 8414 36586 8430 36620
rect 8498 36586 8514 36620
rect 8414 36570 8514 36586
rect 8572 36620 8672 36658
rect 8572 36586 8588 36620
rect 8656 36586 8672 36620
rect 8572 36570 8672 36586
rect 8730 36620 8830 36658
rect 8730 36586 8746 36620
rect 8814 36586 8830 36620
rect 8730 36570 8830 36586
rect 8888 36620 8988 36658
rect 8888 36586 8904 36620
rect 8972 36586 8988 36620
rect 8888 36570 8988 36586
rect 9046 36620 9146 36658
rect 9046 36586 9062 36620
rect 9130 36586 9146 36620
rect 9046 36570 9146 36586
rect 9204 36620 9304 36658
rect 9204 36586 9220 36620
rect 9288 36586 9304 36620
rect 9204 36570 9304 36586
rect 9362 36620 9462 36658
rect 9362 36586 9378 36620
rect 9446 36586 9462 36620
rect 9362 36570 9462 36586
rect 9520 36620 9620 36658
rect 9520 36586 9536 36620
rect 9604 36586 9620 36620
rect 9520 36570 9620 36586
rect 9678 36620 9778 36658
rect 9678 36586 9694 36620
rect 9762 36586 9778 36620
rect 9678 36570 9778 36586
rect 9836 36620 9936 36658
rect 9836 36586 9852 36620
rect 9920 36586 9936 36620
rect 9836 36570 9936 36586
rect 9994 36620 10094 36658
rect 9994 36586 10010 36620
rect 10078 36586 10094 36620
rect 9994 36570 10094 36586
rect 10152 36620 10252 36658
rect 10152 36586 10168 36620
rect 10236 36586 10252 36620
rect 10152 36570 10252 36586
rect 10310 36620 10410 36658
rect 10310 36586 10326 36620
rect 10394 36586 10410 36620
rect 10310 36570 10410 36586
rect -13172 34430 -13072 34446
rect -13172 34396 -13156 34430
rect -13088 34396 -13072 34430
rect -13172 34358 -13072 34396
rect -13014 34430 -12914 34446
rect -13014 34396 -12998 34430
rect -12930 34396 -12914 34430
rect -13014 34358 -12914 34396
rect -12856 34430 -12756 34446
rect -12856 34396 -12840 34430
rect -12772 34396 -12756 34430
rect -12856 34358 -12756 34396
rect -12698 34430 -12598 34446
rect -12698 34396 -12682 34430
rect -12614 34396 -12598 34430
rect -12698 34358 -12598 34396
rect -12540 34430 -12440 34446
rect -12540 34396 -12524 34430
rect -12456 34396 -12440 34430
rect -12540 34358 -12440 34396
rect -12382 34430 -12282 34446
rect -12382 34396 -12366 34430
rect -12298 34396 -12282 34430
rect -12382 34358 -12282 34396
rect -12224 34430 -12124 34446
rect -12224 34396 -12208 34430
rect -12140 34396 -12124 34430
rect -12224 34358 -12124 34396
rect -12066 34430 -11966 34446
rect -12066 34396 -12050 34430
rect -11982 34396 -11966 34430
rect -12066 34358 -11966 34396
rect -11908 34430 -11808 34446
rect -11908 34396 -11892 34430
rect -11824 34396 -11808 34430
rect -11908 34358 -11808 34396
rect -11750 34430 -11650 34446
rect -11750 34396 -11734 34430
rect -11666 34396 -11650 34430
rect -11750 34358 -11650 34396
rect -11592 34430 -11492 34446
rect -11592 34396 -11576 34430
rect -11508 34396 -11492 34430
rect -11592 34358 -11492 34396
rect -11434 34430 -11334 34446
rect -11434 34396 -11418 34430
rect -11350 34396 -11334 34430
rect -11434 34358 -11334 34396
rect -11276 34430 -11176 34446
rect -11276 34396 -11260 34430
rect -11192 34396 -11176 34430
rect -11276 34358 -11176 34396
rect -11118 34430 -11018 34446
rect -11118 34396 -11102 34430
rect -11034 34396 -11018 34430
rect -11118 34358 -11018 34396
rect -10960 34430 -10860 34446
rect -10960 34396 -10944 34430
rect -10876 34396 -10860 34430
rect -10960 34358 -10860 34396
rect -10802 34430 -10702 34446
rect -10802 34396 -10786 34430
rect -10718 34396 -10702 34430
rect -10802 34358 -10702 34396
rect -10644 34430 -10544 34446
rect -10644 34396 -10628 34430
rect -10560 34396 -10544 34430
rect -10644 34358 -10544 34396
rect -10486 34430 -10386 34446
rect -10486 34396 -10470 34430
rect -10402 34396 -10386 34430
rect -10486 34358 -10386 34396
rect -10328 34430 -10228 34446
rect -10328 34396 -10312 34430
rect -10244 34396 -10228 34430
rect -10328 34358 -10228 34396
rect -10170 34430 -10070 34446
rect -10170 34396 -10154 34430
rect -10086 34396 -10070 34430
rect -10170 34358 -10070 34396
rect -10012 34430 -9912 34446
rect -10012 34396 -9996 34430
rect -9928 34396 -9912 34430
rect -10012 34358 -9912 34396
rect -9854 34430 -9754 34446
rect -9854 34396 -9838 34430
rect -9770 34396 -9754 34430
rect -9854 34358 -9754 34396
rect -9696 34430 -9596 34446
rect -9696 34396 -9680 34430
rect -9612 34396 -9596 34430
rect -9696 34358 -9596 34396
rect -9538 34430 -9438 34446
rect -9538 34396 -9522 34430
rect -9454 34396 -9438 34430
rect -9538 34358 -9438 34396
rect -9380 34430 -9280 34446
rect -9380 34396 -9364 34430
rect -9296 34396 -9280 34430
rect -9380 34358 -9280 34396
rect -9222 34430 -9122 34446
rect -9222 34396 -9206 34430
rect -9138 34396 -9122 34430
rect -9222 34358 -9122 34396
rect -9064 34430 -8964 34446
rect -9064 34396 -9048 34430
rect -8980 34396 -8964 34430
rect -9064 34358 -8964 34396
rect -8906 34430 -8806 34446
rect -8906 34396 -8890 34430
rect -8822 34396 -8806 34430
rect -8906 34358 -8806 34396
rect -8748 34430 -8648 34446
rect -8748 34396 -8732 34430
rect -8664 34396 -8648 34430
rect -8748 34358 -8648 34396
rect -8590 34430 -8490 34446
rect -8590 34396 -8574 34430
rect -8506 34396 -8490 34430
rect -8590 34358 -8490 34396
rect -13172 28320 -13072 28358
rect -13172 28286 -13156 28320
rect -13088 28286 -13072 28320
rect -13172 28270 -13072 28286
rect -13014 28320 -12914 28358
rect -13014 28286 -12998 28320
rect -12930 28286 -12914 28320
rect -13014 28270 -12914 28286
rect -12856 28320 -12756 28358
rect -12856 28286 -12840 28320
rect -12772 28286 -12756 28320
rect -12856 28270 -12756 28286
rect -12698 28320 -12598 28358
rect -12698 28286 -12682 28320
rect -12614 28286 -12598 28320
rect -12698 28270 -12598 28286
rect -12540 28320 -12440 28358
rect -12540 28286 -12524 28320
rect -12456 28286 -12440 28320
rect -12540 28270 -12440 28286
rect -12382 28320 -12282 28358
rect -12382 28286 -12366 28320
rect -12298 28286 -12282 28320
rect -12382 28270 -12282 28286
rect -12224 28320 -12124 28358
rect -12224 28286 -12208 28320
rect -12140 28286 -12124 28320
rect -12224 28270 -12124 28286
rect -12066 28320 -11966 28358
rect -12066 28286 -12050 28320
rect -11982 28286 -11966 28320
rect -12066 28270 -11966 28286
rect -11908 28320 -11808 28358
rect -11908 28286 -11892 28320
rect -11824 28286 -11808 28320
rect -11908 28270 -11808 28286
rect -11750 28320 -11650 28358
rect -11750 28286 -11734 28320
rect -11666 28286 -11650 28320
rect -11750 28270 -11650 28286
rect -11592 28320 -11492 28358
rect -11592 28286 -11576 28320
rect -11508 28286 -11492 28320
rect -11592 28270 -11492 28286
rect -11434 28320 -11334 28358
rect -11434 28286 -11418 28320
rect -11350 28286 -11334 28320
rect -11434 28270 -11334 28286
rect -11276 28320 -11176 28358
rect -11276 28286 -11260 28320
rect -11192 28286 -11176 28320
rect -11276 28270 -11176 28286
rect -11118 28320 -11018 28358
rect -11118 28286 -11102 28320
rect -11034 28286 -11018 28320
rect -11118 28270 -11018 28286
rect -10960 28320 -10860 28358
rect -10960 28286 -10944 28320
rect -10876 28286 -10860 28320
rect -10960 28270 -10860 28286
rect -10802 28320 -10702 28358
rect -10802 28286 -10786 28320
rect -10718 28286 -10702 28320
rect -10802 28270 -10702 28286
rect -10644 28320 -10544 28358
rect -10644 28286 -10628 28320
rect -10560 28286 -10544 28320
rect -10644 28270 -10544 28286
rect -10486 28320 -10386 28358
rect -10486 28286 -10470 28320
rect -10402 28286 -10386 28320
rect -10486 28270 -10386 28286
rect -10328 28320 -10228 28358
rect -10328 28286 -10312 28320
rect -10244 28286 -10228 28320
rect -10328 28270 -10228 28286
rect -10170 28320 -10070 28358
rect -10170 28286 -10154 28320
rect -10086 28286 -10070 28320
rect -10170 28270 -10070 28286
rect -10012 28320 -9912 28358
rect -10012 28286 -9996 28320
rect -9928 28286 -9912 28320
rect -10012 28270 -9912 28286
rect -9854 28320 -9754 28358
rect -9854 28286 -9838 28320
rect -9770 28286 -9754 28320
rect -9854 28270 -9754 28286
rect -9696 28320 -9596 28358
rect -9696 28286 -9680 28320
rect -9612 28286 -9596 28320
rect -9696 28270 -9596 28286
rect -9538 28320 -9438 28358
rect -9538 28286 -9522 28320
rect -9454 28286 -9438 28320
rect -9538 28270 -9438 28286
rect -9380 28320 -9280 28358
rect -9380 28286 -9364 28320
rect -9296 28286 -9280 28320
rect -9380 28270 -9280 28286
rect -9222 28320 -9122 28358
rect -9222 28286 -9206 28320
rect -9138 28286 -9122 28320
rect -9222 28270 -9122 28286
rect -9064 28320 -8964 28358
rect -9064 28286 -9048 28320
rect -8980 28286 -8964 28320
rect -9064 28270 -8964 28286
rect -8906 28320 -8806 28358
rect -8906 28286 -8890 28320
rect -8822 28286 -8806 28320
rect -8906 28270 -8806 28286
rect -8748 28320 -8648 28358
rect -8748 28286 -8732 28320
rect -8664 28286 -8648 28320
rect -8748 28270 -8648 28286
rect -8590 28320 -8490 28358
rect -8590 28286 -8574 28320
rect -8506 28286 -8490 28320
rect -8590 28270 -8490 28286
rect -6872 34430 -6772 34446
rect -6872 34396 -6856 34430
rect -6788 34396 -6772 34430
rect -6872 34358 -6772 34396
rect -6714 34430 -6614 34446
rect -6714 34396 -6698 34430
rect -6630 34396 -6614 34430
rect -6714 34358 -6614 34396
rect -6556 34430 -6456 34446
rect -6556 34396 -6540 34430
rect -6472 34396 -6456 34430
rect -6556 34358 -6456 34396
rect -6398 34430 -6298 34446
rect -6398 34396 -6382 34430
rect -6314 34396 -6298 34430
rect -6398 34358 -6298 34396
rect -6240 34430 -6140 34446
rect -6240 34396 -6224 34430
rect -6156 34396 -6140 34430
rect -6240 34358 -6140 34396
rect -6082 34430 -5982 34446
rect -6082 34396 -6066 34430
rect -5998 34396 -5982 34430
rect -6082 34358 -5982 34396
rect -5924 34430 -5824 34446
rect -5924 34396 -5908 34430
rect -5840 34396 -5824 34430
rect -5924 34358 -5824 34396
rect -5766 34430 -5666 34446
rect -5766 34396 -5750 34430
rect -5682 34396 -5666 34430
rect -5766 34358 -5666 34396
rect -5608 34430 -5508 34446
rect -5608 34396 -5592 34430
rect -5524 34396 -5508 34430
rect -5608 34358 -5508 34396
rect -5450 34430 -5350 34446
rect -5450 34396 -5434 34430
rect -5366 34396 -5350 34430
rect -5450 34358 -5350 34396
rect -5292 34430 -5192 34446
rect -5292 34396 -5276 34430
rect -5208 34396 -5192 34430
rect -5292 34358 -5192 34396
rect -5134 34430 -5034 34446
rect -5134 34396 -5118 34430
rect -5050 34396 -5034 34430
rect -5134 34358 -5034 34396
rect -4976 34430 -4876 34446
rect -4976 34396 -4960 34430
rect -4892 34396 -4876 34430
rect -4976 34358 -4876 34396
rect -4818 34430 -4718 34446
rect -4818 34396 -4802 34430
rect -4734 34396 -4718 34430
rect -4818 34358 -4718 34396
rect -4660 34430 -4560 34446
rect -4660 34396 -4644 34430
rect -4576 34396 -4560 34430
rect -4660 34358 -4560 34396
rect -4502 34430 -4402 34446
rect -4502 34396 -4486 34430
rect -4418 34396 -4402 34430
rect -4502 34358 -4402 34396
rect -4344 34430 -4244 34446
rect -4344 34396 -4328 34430
rect -4260 34396 -4244 34430
rect -4344 34358 -4244 34396
rect -4186 34430 -4086 34446
rect -4186 34396 -4170 34430
rect -4102 34396 -4086 34430
rect -4186 34358 -4086 34396
rect -4028 34430 -3928 34446
rect -4028 34396 -4012 34430
rect -3944 34396 -3928 34430
rect -4028 34358 -3928 34396
rect -3870 34430 -3770 34446
rect -3870 34396 -3854 34430
rect -3786 34396 -3770 34430
rect -3870 34358 -3770 34396
rect -3712 34430 -3612 34446
rect -3712 34396 -3696 34430
rect -3628 34396 -3612 34430
rect -3712 34358 -3612 34396
rect -3554 34430 -3454 34446
rect -3554 34396 -3538 34430
rect -3470 34396 -3454 34430
rect -3554 34358 -3454 34396
rect -3396 34430 -3296 34446
rect -3396 34396 -3380 34430
rect -3312 34396 -3296 34430
rect -3396 34358 -3296 34396
rect -3238 34430 -3138 34446
rect -3238 34396 -3222 34430
rect -3154 34396 -3138 34430
rect -3238 34358 -3138 34396
rect -3080 34430 -2980 34446
rect -3080 34396 -3064 34430
rect -2996 34396 -2980 34430
rect -3080 34358 -2980 34396
rect -2922 34430 -2822 34446
rect -2922 34396 -2906 34430
rect -2838 34396 -2822 34430
rect -2922 34358 -2822 34396
rect -2764 34430 -2664 34446
rect -2764 34396 -2748 34430
rect -2680 34396 -2664 34430
rect -2764 34358 -2664 34396
rect -2606 34430 -2506 34446
rect -2606 34396 -2590 34430
rect -2522 34396 -2506 34430
rect -2606 34358 -2506 34396
rect -2448 34430 -2348 34446
rect -2448 34396 -2432 34430
rect -2364 34396 -2348 34430
rect -2448 34358 -2348 34396
rect -2290 34430 -2190 34446
rect -2290 34396 -2274 34430
rect -2206 34396 -2190 34430
rect -2290 34358 -2190 34396
rect -6872 28320 -6772 28358
rect -6872 28286 -6856 28320
rect -6788 28286 -6772 28320
rect -6872 28270 -6772 28286
rect -6714 28320 -6614 28358
rect -6714 28286 -6698 28320
rect -6630 28286 -6614 28320
rect -6714 28270 -6614 28286
rect -6556 28320 -6456 28358
rect -6556 28286 -6540 28320
rect -6472 28286 -6456 28320
rect -6556 28270 -6456 28286
rect -6398 28320 -6298 28358
rect -6398 28286 -6382 28320
rect -6314 28286 -6298 28320
rect -6398 28270 -6298 28286
rect -6240 28320 -6140 28358
rect -6240 28286 -6224 28320
rect -6156 28286 -6140 28320
rect -6240 28270 -6140 28286
rect -6082 28320 -5982 28358
rect -6082 28286 -6066 28320
rect -5998 28286 -5982 28320
rect -6082 28270 -5982 28286
rect -5924 28320 -5824 28358
rect -5924 28286 -5908 28320
rect -5840 28286 -5824 28320
rect -5924 28270 -5824 28286
rect -5766 28320 -5666 28358
rect -5766 28286 -5750 28320
rect -5682 28286 -5666 28320
rect -5766 28270 -5666 28286
rect -5608 28320 -5508 28358
rect -5608 28286 -5592 28320
rect -5524 28286 -5508 28320
rect -5608 28270 -5508 28286
rect -5450 28320 -5350 28358
rect -5450 28286 -5434 28320
rect -5366 28286 -5350 28320
rect -5450 28270 -5350 28286
rect -5292 28320 -5192 28358
rect -5292 28286 -5276 28320
rect -5208 28286 -5192 28320
rect -5292 28270 -5192 28286
rect -5134 28320 -5034 28358
rect -5134 28286 -5118 28320
rect -5050 28286 -5034 28320
rect -5134 28270 -5034 28286
rect -4976 28320 -4876 28358
rect -4976 28286 -4960 28320
rect -4892 28286 -4876 28320
rect -4976 28270 -4876 28286
rect -4818 28320 -4718 28358
rect -4818 28286 -4802 28320
rect -4734 28286 -4718 28320
rect -4818 28270 -4718 28286
rect -4660 28320 -4560 28358
rect -4660 28286 -4644 28320
rect -4576 28286 -4560 28320
rect -4660 28270 -4560 28286
rect -4502 28320 -4402 28358
rect -4502 28286 -4486 28320
rect -4418 28286 -4402 28320
rect -4502 28270 -4402 28286
rect -4344 28320 -4244 28358
rect -4344 28286 -4328 28320
rect -4260 28286 -4244 28320
rect -4344 28270 -4244 28286
rect -4186 28320 -4086 28358
rect -4186 28286 -4170 28320
rect -4102 28286 -4086 28320
rect -4186 28270 -4086 28286
rect -4028 28320 -3928 28358
rect -4028 28286 -4012 28320
rect -3944 28286 -3928 28320
rect -4028 28270 -3928 28286
rect -3870 28320 -3770 28358
rect -3870 28286 -3854 28320
rect -3786 28286 -3770 28320
rect -3870 28270 -3770 28286
rect -3712 28320 -3612 28358
rect -3712 28286 -3696 28320
rect -3628 28286 -3612 28320
rect -3712 28270 -3612 28286
rect -3554 28320 -3454 28358
rect -3554 28286 -3538 28320
rect -3470 28286 -3454 28320
rect -3554 28270 -3454 28286
rect -3396 28320 -3296 28358
rect -3396 28286 -3380 28320
rect -3312 28286 -3296 28320
rect -3396 28270 -3296 28286
rect -3238 28320 -3138 28358
rect -3238 28286 -3222 28320
rect -3154 28286 -3138 28320
rect -3238 28270 -3138 28286
rect -3080 28320 -2980 28358
rect -3080 28286 -3064 28320
rect -2996 28286 -2980 28320
rect -3080 28270 -2980 28286
rect -2922 28320 -2822 28358
rect -2922 28286 -2906 28320
rect -2838 28286 -2822 28320
rect -2922 28270 -2822 28286
rect -2764 28320 -2664 28358
rect -2764 28286 -2748 28320
rect -2680 28286 -2664 28320
rect -2764 28270 -2664 28286
rect -2606 28320 -2506 28358
rect -2606 28286 -2590 28320
rect -2522 28286 -2506 28320
rect -2606 28270 -2506 28286
rect -2448 28320 -2348 28358
rect -2448 28286 -2432 28320
rect -2364 28286 -2348 28320
rect -2448 28270 -2348 28286
rect -2290 28320 -2190 28358
rect -2290 28286 -2274 28320
rect -2206 28286 -2190 28320
rect -2290 28270 -2190 28286
rect -572 34430 -472 34446
rect -572 34396 -556 34430
rect -488 34396 -472 34430
rect -572 34358 -472 34396
rect -414 34430 -314 34446
rect -414 34396 -398 34430
rect -330 34396 -314 34430
rect -414 34358 -314 34396
rect -256 34430 -156 34446
rect -256 34396 -240 34430
rect -172 34396 -156 34430
rect -256 34358 -156 34396
rect -98 34430 2 34446
rect -98 34396 -82 34430
rect -14 34396 2 34430
rect -98 34358 2 34396
rect 60 34430 160 34446
rect 60 34396 76 34430
rect 144 34396 160 34430
rect 60 34358 160 34396
rect 218 34430 318 34446
rect 218 34396 234 34430
rect 302 34396 318 34430
rect 218 34358 318 34396
rect 376 34430 476 34446
rect 376 34396 392 34430
rect 460 34396 476 34430
rect 376 34358 476 34396
rect 534 34430 634 34446
rect 534 34396 550 34430
rect 618 34396 634 34430
rect 534 34358 634 34396
rect 692 34430 792 34446
rect 692 34396 708 34430
rect 776 34396 792 34430
rect 692 34358 792 34396
rect 850 34430 950 34446
rect 850 34396 866 34430
rect 934 34396 950 34430
rect 850 34358 950 34396
rect 1008 34430 1108 34446
rect 1008 34396 1024 34430
rect 1092 34396 1108 34430
rect 1008 34358 1108 34396
rect 1166 34430 1266 34446
rect 1166 34396 1182 34430
rect 1250 34396 1266 34430
rect 1166 34358 1266 34396
rect 1324 34430 1424 34446
rect 1324 34396 1340 34430
rect 1408 34396 1424 34430
rect 1324 34358 1424 34396
rect 1482 34430 1582 34446
rect 1482 34396 1498 34430
rect 1566 34396 1582 34430
rect 1482 34358 1582 34396
rect 1640 34430 1740 34446
rect 1640 34396 1656 34430
rect 1724 34396 1740 34430
rect 1640 34358 1740 34396
rect 1798 34430 1898 34446
rect 1798 34396 1814 34430
rect 1882 34396 1898 34430
rect 1798 34358 1898 34396
rect 1956 34430 2056 34446
rect 1956 34396 1972 34430
rect 2040 34396 2056 34430
rect 1956 34358 2056 34396
rect 2114 34430 2214 34446
rect 2114 34396 2130 34430
rect 2198 34396 2214 34430
rect 2114 34358 2214 34396
rect 2272 34430 2372 34446
rect 2272 34396 2288 34430
rect 2356 34396 2372 34430
rect 2272 34358 2372 34396
rect 2430 34430 2530 34446
rect 2430 34396 2446 34430
rect 2514 34396 2530 34430
rect 2430 34358 2530 34396
rect 2588 34430 2688 34446
rect 2588 34396 2604 34430
rect 2672 34396 2688 34430
rect 2588 34358 2688 34396
rect 2746 34430 2846 34446
rect 2746 34396 2762 34430
rect 2830 34396 2846 34430
rect 2746 34358 2846 34396
rect 2904 34430 3004 34446
rect 2904 34396 2920 34430
rect 2988 34396 3004 34430
rect 2904 34358 3004 34396
rect 3062 34430 3162 34446
rect 3062 34396 3078 34430
rect 3146 34396 3162 34430
rect 3062 34358 3162 34396
rect 3220 34430 3320 34446
rect 3220 34396 3236 34430
rect 3304 34396 3320 34430
rect 3220 34358 3320 34396
rect 3378 34430 3478 34446
rect 3378 34396 3394 34430
rect 3462 34396 3478 34430
rect 3378 34358 3478 34396
rect 3536 34430 3636 34446
rect 3536 34396 3552 34430
rect 3620 34396 3636 34430
rect 3536 34358 3636 34396
rect 3694 34430 3794 34446
rect 3694 34396 3710 34430
rect 3778 34396 3794 34430
rect 3694 34358 3794 34396
rect 3852 34430 3952 34446
rect 3852 34396 3868 34430
rect 3936 34396 3952 34430
rect 3852 34358 3952 34396
rect 4010 34430 4110 34446
rect 4010 34396 4026 34430
rect 4094 34396 4110 34430
rect 4010 34358 4110 34396
rect -572 28320 -472 28358
rect -572 28286 -556 28320
rect -488 28286 -472 28320
rect -572 28270 -472 28286
rect -414 28320 -314 28358
rect -414 28286 -398 28320
rect -330 28286 -314 28320
rect -414 28270 -314 28286
rect -256 28320 -156 28358
rect -256 28286 -240 28320
rect -172 28286 -156 28320
rect -256 28270 -156 28286
rect -98 28320 2 28358
rect -98 28286 -82 28320
rect -14 28286 2 28320
rect -98 28270 2 28286
rect 60 28320 160 28358
rect 60 28286 76 28320
rect 144 28286 160 28320
rect 60 28270 160 28286
rect 218 28320 318 28358
rect 218 28286 234 28320
rect 302 28286 318 28320
rect 218 28270 318 28286
rect 376 28320 476 28358
rect 376 28286 392 28320
rect 460 28286 476 28320
rect 376 28270 476 28286
rect 534 28320 634 28358
rect 534 28286 550 28320
rect 618 28286 634 28320
rect 534 28270 634 28286
rect 692 28320 792 28358
rect 692 28286 708 28320
rect 776 28286 792 28320
rect 692 28270 792 28286
rect 850 28320 950 28358
rect 850 28286 866 28320
rect 934 28286 950 28320
rect 850 28270 950 28286
rect 1008 28320 1108 28358
rect 1008 28286 1024 28320
rect 1092 28286 1108 28320
rect 1008 28270 1108 28286
rect 1166 28320 1266 28358
rect 1166 28286 1182 28320
rect 1250 28286 1266 28320
rect 1166 28270 1266 28286
rect 1324 28320 1424 28358
rect 1324 28286 1340 28320
rect 1408 28286 1424 28320
rect 1324 28270 1424 28286
rect 1482 28320 1582 28358
rect 1482 28286 1498 28320
rect 1566 28286 1582 28320
rect 1482 28270 1582 28286
rect 1640 28320 1740 28358
rect 1640 28286 1656 28320
rect 1724 28286 1740 28320
rect 1640 28270 1740 28286
rect 1798 28320 1898 28358
rect 1798 28286 1814 28320
rect 1882 28286 1898 28320
rect 1798 28270 1898 28286
rect 1956 28320 2056 28358
rect 1956 28286 1972 28320
rect 2040 28286 2056 28320
rect 1956 28270 2056 28286
rect 2114 28320 2214 28358
rect 2114 28286 2130 28320
rect 2198 28286 2214 28320
rect 2114 28270 2214 28286
rect 2272 28320 2372 28358
rect 2272 28286 2288 28320
rect 2356 28286 2372 28320
rect 2272 28270 2372 28286
rect 2430 28320 2530 28358
rect 2430 28286 2446 28320
rect 2514 28286 2530 28320
rect 2430 28270 2530 28286
rect 2588 28320 2688 28358
rect 2588 28286 2604 28320
rect 2672 28286 2688 28320
rect 2588 28270 2688 28286
rect 2746 28320 2846 28358
rect 2746 28286 2762 28320
rect 2830 28286 2846 28320
rect 2746 28270 2846 28286
rect 2904 28320 3004 28358
rect 2904 28286 2920 28320
rect 2988 28286 3004 28320
rect 2904 28270 3004 28286
rect 3062 28320 3162 28358
rect 3062 28286 3078 28320
rect 3146 28286 3162 28320
rect 3062 28270 3162 28286
rect 3220 28320 3320 28358
rect 3220 28286 3236 28320
rect 3304 28286 3320 28320
rect 3220 28270 3320 28286
rect 3378 28320 3478 28358
rect 3378 28286 3394 28320
rect 3462 28286 3478 28320
rect 3378 28270 3478 28286
rect 3536 28320 3636 28358
rect 3536 28286 3552 28320
rect 3620 28286 3636 28320
rect 3536 28270 3636 28286
rect 3694 28320 3794 28358
rect 3694 28286 3710 28320
rect 3778 28286 3794 28320
rect 3694 28270 3794 28286
rect 3852 28320 3952 28358
rect 3852 28286 3868 28320
rect 3936 28286 3952 28320
rect 3852 28270 3952 28286
rect 4010 28320 4110 28358
rect 4010 28286 4026 28320
rect 4094 28286 4110 28320
rect 4010 28270 4110 28286
rect 5728 34430 5828 34446
rect 5728 34396 5744 34430
rect 5812 34396 5828 34430
rect 5728 34358 5828 34396
rect 5886 34430 5986 34446
rect 5886 34396 5902 34430
rect 5970 34396 5986 34430
rect 5886 34358 5986 34396
rect 6044 34430 6144 34446
rect 6044 34396 6060 34430
rect 6128 34396 6144 34430
rect 6044 34358 6144 34396
rect 6202 34430 6302 34446
rect 6202 34396 6218 34430
rect 6286 34396 6302 34430
rect 6202 34358 6302 34396
rect 6360 34430 6460 34446
rect 6360 34396 6376 34430
rect 6444 34396 6460 34430
rect 6360 34358 6460 34396
rect 6518 34430 6618 34446
rect 6518 34396 6534 34430
rect 6602 34396 6618 34430
rect 6518 34358 6618 34396
rect 6676 34430 6776 34446
rect 6676 34396 6692 34430
rect 6760 34396 6776 34430
rect 6676 34358 6776 34396
rect 6834 34430 6934 34446
rect 6834 34396 6850 34430
rect 6918 34396 6934 34430
rect 6834 34358 6934 34396
rect 6992 34430 7092 34446
rect 6992 34396 7008 34430
rect 7076 34396 7092 34430
rect 6992 34358 7092 34396
rect 7150 34430 7250 34446
rect 7150 34396 7166 34430
rect 7234 34396 7250 34430
rect 7150 34358 7250 34396
rect 7308 34430 7408 34446
rect 7308 34396 7324 34430
rect 7392 34396 7408 34430
rect 7308 34358 7408 34396
rect 7466 34430 7566 34446
rect 7466 34396 7482 34430
rect 7550 34396 7566 34430
rect 7466 34358 7566 34396
rect 7624 34430 7724 34446
rect 7624 34396 7640 34430
rect 7708 34396 7724 34430
rect 7624 34358 7724 34396
rect 7782 34430 7882 34446
rect 7782 34396 7798 34430
rect 7866 34396 7882 34430
rect 7782 34358 7882 34396
rect 7940 34430 8040 34446
rect 7940 34396 7956 34430
rect 8024 34396 8040 34430
rect 7940 34358 8040 34396
rect 8098 34430 8198 34446
rect 8098 34396 8114 34430
rect 8182 34396 8198 34430
rect 8098 34358 8198 34396
rect 8256 34430 8356 34446
rect 8256 34396 8272 34430
rect 8340 34396 8356 34430
rect 8256 34358 8356 34396
rect 8414 34430 8514 34446
rect 8414 34396 8430 34430
rect 8498 34396 8514 34430
rect 8414 34358 8514 34396
rect 8572 34430 8672 34446
rect 8572 34396 8588 34430
rect 8656 34396 8672 34430
rect 8572 34358 8672 34396
rect 8730 34430 8830 34446
rect 8730 34396 8746 34430
rect 8814 34396 8830 34430
rect 8730 34358 8830 34396
rect 8888 34430 8988 34446
rect 8888 34396 8904 34430
rect 8972 34396 8988 34430
rect 8888 34358 8988 34396
rect 9046 34430 9146 34446
rect 9046 34396 9062 34430
rect 9130 34396 9146 34430
rect 9046 34358 9146 34396
rect 9204 34430 9304 34446
rect 9204 34396 9220 34430
rect 9288 34396 9304 34430
rect 9204 34358 9304 34396
rect 9362 34430 9462 34446
rect 9362 34396 9378 34430
rect 9446 34396 9462 34430
rect 9362 34358 9462 34396
rect 9520 34430 9620 34446
rect 9520 34396 9536 34430
rect 9604 34396 9620 34430
rect 9520 34358 9620 34396
rect 9678 34430 9778 34446
rect 9678 34396 9694 34430
rect 9762 34396 9778 34430
rect 9678 34358 9778 34396
rect 9836 34430 9936 34446
rect 9836 34396 9852 34430
rect 9920 34396 9936 34430
rect 9836 34358 9936 34396
rect 9994 34430 10094 34446
rect 9994 34396 10010 34430
rect 10078 34396 10094 34430
rect 9994 34358 10094 34396
rect 10152 34430 10252 34446
rect 10152 34396 10168 34430
rect 10236 34396 10252 34430
rect 10152 34358 10252 34396
rect 10310 34430 10410 34446
rect 10310 34396 10326 34430
rect 10394 34396 10410 34430
rect 10310 34358 10410 34396
rect 5728 28320 5828 28358
rect 5728 28286 5744 28320
rect 5812 28286 5828 28320
rect 5728 28270 5828 28286
rect 5886 28320 5986 28358
rect 5886 28286 5902 28320
rect 5970 28286 5986 28320
rect 5886 28270 5986 28286
rect 6044 28320 6144 28358
rect 6044 28286 6060 28320
rect 6128 28286 6144 28320
rect 6044 28270 6144 28286
rect 6202 28320 6302 28358
rect 6202 28286 6218 28320
rect 6286 28286 6302 28320
rect 6202 28270 6302 28286
rect 6360 28320 6460 28358
rect 6360 28286 6376 28320
rect 6444 28286 6460 28320
rect 6360 28270 6460 28286
rect 6518 28320 6618 28358
rect 6518 28286 6534 28320
rect 6602 28286 6618 28320
rect 6518 28270 6618 28286
rect 6676 28320 6776 28358
rect 6676 28286 6692 28320
rect 6760 28286 6776 28320
rect 6676 28270 6776 28286
rect 6834 28320 6934 28358
rect 6834 28286 6850 28320
rect 6918 28286 6934 28320
rect 6834 28270 6934 28286
rect 6992 28320 7092 28358
rect 6992 28286 7008 28320
rect 7076 28286 7092 28320
rect 6992 28270 7092 28286
rect 7150 28320 7250 28358
rect 7150 28286 7166 28320
rect 7234 28286 7250 28320
rect 7150 28270 7250 28286
rect 7308 28320 7408 28358
rect 7308 28286 7324 28320
rect 7392 28286 7408 28320
rect 7308 28270 7408 28286
rect 7466 28320 7566 28358
rect 7466 28286 7482 28320
rect 7550 28286 7566 28320
rect 7466 28270 7566 28286
rect 7624 28320 7724 28358
rect 7624 28286 7640 28320
rect 7708 28286 7724 28320
rect 7624 28270 7724 28286
rect 7782 28320 7882 28358
rect 7782 28286 7798 28320
rect 7866 28286 7882 28320
rect 7782 28270 7882 28286
rect 7940 28320 8040 28358
rect 7940 28286 7956 28320
rect 8024 28286 8040 28320
rect 7940 28270 8040 28286
rect 8098 28320 8198 28358
rect 8098 28286 8114 28320
rect 8182 28286 8198 28320
rect 8098 28270 8198 28286
rect 8256 28320 8356 28358
rect 8256 28286 8272 28320
rect 8340 28286 8356 28320
rect 8256 28270 8356 28286
rect 8414 28320 8514 28358
rect 8414 28286 8430 28320
rect 8498 28286 8514 28320
rect 8414 28270 8514 28286
rect 8572 28320 8672 28358
rect 8572 28286 8588 28320
rect 8656 28286 8672 28320
rect 8572 28270 8672 28286
rect 8730 28320 8830 28358
rect 8730 28286 8746 28320
rect 8814 28286 8830 28320
rect 8730 28270 8830 28286
rect 8888 28320 8988 28358
rect 8888 28286 8904 28320
rect 8972 28286 8988 28320
rect 8888 28270 8988 28286
rect 9046 28320 9146 28358
rect 9046 28286 9062 28320
rect 9130 28286 9146 28320
rect 9046 28270 9146 28286
rect 9204 28320 9304 28358
rect 9204 28286 9220 28320
rect 9288 28286 9304 28320
rect 9204 28270 9304 28286
rect 9362 28320 9462 28358
rect 9362 28286 9378 28320
rect 9446 28286 9462 28320
rect 9362 28270 9462 28286
rect 9520 28320 9620 28358
rect 9520 28286 9536 28320
rect 9604 28286 9620 28320
rect 9520 28270 9620 28286
rect 9678 28320 9778 28358
rect 9678 28286 9694 28320
rect 9762 28286 9778 28320
rect 9678 28270 9778 28286
rect 9836 28320 9936 28358
rect 9836 28286 9852 28320
rect 9920 28286 9936 28320
rect 9836 28270 9936 28286
rect 9994 28320 10094 28358
rect 9994 28286 10010 28320
rect 10078 28286 10094 28320
rect 9994 28270 10094 28286
rect 10152 28320 10252 28358
rect 10152 28286 10168 28320
rect 10236 28286 10252 28320
rect 10152 28270 10252 28286
rect 10310 28320 10410 28358
rect 10310 28286 10326 28320
rect 10394 28286 10410 28320
rect 10310 28270 10410 28286
rect -13172 27430 -13072 27446
rect -13172 27396 -13156 27430
rect -13088 27396 -13072 27430
rect -13172 27358 -13072 27396
rect -13014 27430 -12914 27446
rect -13014 27396 -12998 27430
rect -12930 27396 -12914 27430
rect -13014 27358 -12914 27396
rect -12856 27430 -12756 27446
rect -12856 27396 -12840 27430
rect -12772 27396 -12756 27430
rect -12856 27358 -12756 27396
rect -12698 27430 -12598 27446
rect -12698 27396 -12682 27430
rect -12614 27396 -12598 27430
rect -12698 27358 -12598 27396
rect -12540 27430 -12440 27446
rect -12540 27396 -12524 27430
rect -12456 27396 -12440 27430
rect -12540 27358 -12440 27396
rect -12382 27430 -12282 27446
rect -12382 27396 -12366 27430
rect -12298 27396 -12282 27430
rect -12382 27358 -12282 27396
rect -12224 27430 -12124 27446
rect -12224 27396 -12208 27430
rect -12140 27396 -12124 27430
rect -12224 27358 -12124 27396
rect -12066 27430 -11966 27446
rect -12066 27396 -12050 27430
rect -11982 27396 -11966 27430
rect -12066 27358 -11966 27396
rect -11908 27430 -11808 27446
rect -11908 27396 -11892 27430
rect -11824 27396 -11808 27430
rect -11908 27358 -11808 27396
rect -11750 27430 -11650 27446
rect -11750 27396 -11734 27430
rect -11666 27396 -11650 27430
rect -11750 27358 -11650 27396
rect -11592 27430 -11492 27446
rect -11592 27396 -11576 27430
rect -11508 27396 -11492 27430
rect -11592 27358 -11492 27396
rect -11434 27430 -11334 27446
rect -11434 27396 -11418 27430
rect -11350 27396 -11334 27430
rect -11434 27358 -11334 27396
rect -11276 27430 -11176 27446
rect -11276 27396 -11260 27430
rect -11192 27396 -11176 27430
rect -11276 27358 -11176 27396
rect -11118 27430 -11018 27446
rect -11118 27396 -11102 27430
rect -11034 27396 -11018 27430
rect -11118 27358 -11018 27396
rect -10960 27430 -10860 27446
rect -10960 27396 -10944 27430
rect -10876 27396 -10860 27430
rect -10960 27358 -10860 27396
rect -10802 27430 -10702 27446
rect -10802 27396 -10786 27430
rect -10718 27396 -10702 27430
rect -10802 27358 -10702 27396
rect -10644 27430 -10544 27446
rect -10644 27396 -10628 27430
rect -10560 27396 -10544 27430
rect -10644 27358 -10544 27396
rect -10486 27430 -10386 27446
rect -10486 27396 -10470 27430
rect -10402 27396 -10386 27430
rect -10486 27358 -10386 27396
rect -10328 27430 -10228 27446
rect -10328 27396 -10312 27430
rect -10244 27396 -10228 27430
rect -10328 27358 -10228 27396
rect -10170 27430 -10070 27446
rect -10170 27396 -10154 27430
rect -10086 27396 -10070 27430
rect -10170 27358 -10070 27396
rect -10012 27430 -9912 27446
rect -10012 27396 -9996 27430
rect -9928 27396 -9912 27430
rect -10012 27358 -9912 27396
rect -9854 27430 -9754 27446
rect -9854 27396 -9838 27430
rect -9770 27396 -9754 27430
rect -9854 27358 -9754 27396
rect -9696 27430 -9596 27446
rect -9696 27396 -9680 27430
rect -9612 27396 -9596 27430
rect -9696 27358 -9596 27396
rect -9538 27430 -9438 27446
rect -9538 27396 -9522 27430
rect -9454 27396 -9438 27430
rect -9538 27358 -9438 27396
rect -9380 27430 -9280 27446
rect -9380 27396 -9364 27430
rect -9296 27396 -9280 27430
rect -9380 27358 -9280 27396
rect -9222 27430 -9122 27446
rect -9222 27396 -9206 27430
rect -9138 27396 -9122 27430
rect -9222 27358 -9122 27396
rect -9064 27430 -8964 27446
rect -9064 27396 -9048 27430
rect -8980 27396 -8964 27430
rect -9064 27358 -8964 27396
rect -8906 27430 -8806 27446
rect -8906 27396 -8890 27430
rect -8822 27396 -8806 27430
rect -8906 27358 -8806 27396
rect -8748 27430 -8648 27446
rect -8748 27396 -8732 27430
rect -8664 27396 -8648 27430
rect -8748 27358 -8648 27396
rect -8590 27430 -8490 27446
rect -8590 27396 -8574 27430
rect -8506 27396 -8490 27430
rect -8590 27358 -8490 27396
rect -13172 21320 -13072 21358
rect -13172 21286 -13156 21320
rect -13088 21286 -13072 21320
rect -13172 21270 -13072 21286
rect -13014 21320 -12914 21358
rect -13014 21286 -12998 21320
rect -12930 21286 -12914 21320
rect -13014 21270 -12914 21286
rect -12856 21320 -12756 21358
rect -12856 21286 -12840 21320
rect -12772 21286 -12756 21320
rect -12856 21270 -12756 21286
rect -12698 21320 -12598 21358
rect -12698 21286 -12682 21320
rect -12614 21286 -12598 21320
rect -12698 21270 -12598 21286
rect -12540 21320 -12440 21358
rect -12540 21286 -12524 21320
rect -12456 21286 -12440 21320
rect -12540 21270 -12440 21286
rect -12382 21320 -12282 21358
rect -12382 21286 -12366 21320
rect -12298 21286 -12282 21320
rect -12382 21270 -12282 21286
rect -12224 21320 -12124 21358
rect -12224 21286 -12208 21320
rect -12140 21286 -12124 21320
rect -12224 21270 -12124 21286
rect -12066 21320 -11966 21358
rect -12066 21286 -12050 21320
rect -11982 21286 -11966 21320
rect -12066 21270 -11966 21286
rect -11908 21320 -11808 21358
rect -11908 21286 -11892 21320
rect -11824 21286 -11808 21320
rect -11908 21270 -11808 21286
rect -11750 21320 -11650 21358
rect -11750 21286 -11734 21320
rect -11666 21286 -11650 21320
rect -11750 21270 -11650 21286
rect -11592 21320 -11492 21358
rect -11592 21286 -11576 21320
rect -11508 21286 -11492 21320
rect -11592 21270 -11492 21286
rect -11434 21320 -11334 21358
rect -11434 21286 -11418 21320
rect -11350 21286 -11334 21320
rect -11434 21270 -11334 21286
rect -11276 21320 -11176 21358
rect -11276 21286 -11260 21320
rect -11192 21286 -11176 21320
rect -11276 21270 -11176 21286
rect -11118 21320 -11018 21358
rect -11118 21286 -11102 21320
rect -11034 21286 -11018 21320
rect -11118 21270 -11018 21286
rect -10960 21320 -10860 21358
rect -10960 21286 -10944 21320
rect -10876 21286 -10860 21320
rect -10960 21270 -10860 21286
rect -10802 21320 -10702 21358
rect -10802 21286 -10786 21320
rect -10718 21286 -10702 21320
rect -10802 21270 -10702 21286
rect -10644 21320 -10544 21358
rect -10644 21286 -10628 21320
rect -10560 21286 -10544 21320
rect -10644 21270 -10544 21286
rect -10486 21320 -10386 21358
rect -10486 21286 -10470 21320
rect -10402 21286 -10386 21320
rect -10486 21270 -10386 21286
rect -10328 21320 -10228 21358
rect -10328 21286 -10312 21320
rect -10244 21286 -10228 21320
rect -10328 21270 -10228 21286
rect -10170 21320 -10070 21358
rect -10170 21286 -10154 21320
rect -10086 21286 -10070 21320
rect -10170 21270 -10070 21286
rect -10012 21320 -9912 21358
rect -10012 21286 -9996 21320
rect -9928 21286 -9912 21320
rect -10012 21270 -9912 21286
rect -9854 21320 -9754 21358
rect -9854 21286 -9838 21320
rect -9770 21286 -9754 21320
rect -9854 21270 -9754 21286
rect -9696 21320 -9596 21358
rect -9696 21286 -9680 21320
rect -9612 21286 -9596 21320
rect -9696 21270 -9596 21286
rect -9538 21320 -9438 21358
rect -9538 21286 -9522 21320
rect -9454 21286 -9438 21320
rect -9538 21270 -9438 21286
rect -9380 21320 -9280 21358
rect -9380 21286 -9364 21320
rect -9296 21286 -9280 21320
rect -9380 21270 -9280 21286
rect -9222 21320 -9122 21358
rect -9222 21286 -9206 21320
rect -9138 21286 -9122 21320
rect -9222 21270 -9122 21286
rect -9064 21320 -8964 21358
rect -9064 21286 -9048 21320
rect -8980 21286 -8964 21320
rect -9064 21270 -8964 21286
rect -8906 21320 -8806 21358
rect -8906 21286 -8890 21320
rect -8822 21286 -8806 21320
rect -8906 21270 -8806 21286
rect -8748 21320 -8648 21358
rect -8748 21286 -8732 21320
rect -8664 21286 -8648 21320
rect -8748 21270 -8648 21286
rect -8590 21320 -8490 21358
rect -8590 21286 -8574 21320
rect -8506 21286 -8490 21320
rect -8590 21270 -8490 21286
rect -6872 27430 -6772 27446
rect -6872 27396 -6856 27430
rect -6788 27396 -6772 27430
rect -6872 27358 -6772 27396
rect -6714 27430 -6614 27446
rect -6714 27396 -6698 27430
rect -6630 27396 -6614 27430
rect -6714 27358 -6614 27396
rect -6556 27430 -6456 27446
rect -6556 27396 -6540 27430
rect -6472 27396 -6456 27430
rect -6556 27358 -6456 27396
rect -6398 27430 -6298 27446
rect -6398 27396 -6382 27430
rect -6314 27396 -6298 27430
rect -6398 27358 -6298 27396
rect -6240 27430 -6140 27446
rect -6240 27396 -6224 27430
rect -6156 27396 -6140 27430
rect -6240 27358 -6140 27396
rect -6082 27430 -5982 27446
rect -6082 27396 -6066 27430
rect -5998 27396 -5982 27430
rect -6082 27358 -5982 27396
rect -5924 27430 -5824 27446
rect -5924 27396 -5908 27430
rect -5840 27396 -5824 27430
rect -5924 27358 -5824 27396
rect -5766 27430 -5666 27446
rect -5766 27396 -5750 27430
rect -5682 27396 -5666 27430
rect -5766 27358 -5666 27396
rect -5608 27430 -5508 27446
rect -5608 27396 -5592 27430
rect -5524 27396 -5508 27430
rect -5608 27358 -5508 27396
rect -5450 27430 -5350 27446
rect -5450 27396 -5434 27430
rect -5366 27396 -5350 27430
rect -5450 27358 -5350 27396
rect -5292 27430 -5192 27446
rect -5292 27396 -5276 27430
rect -5208 27396 -5192 27430
rect -5292 27358 -5192 27396
rect -5134 27430 -5034 27446
rect -5134 27396 -5118 27430
rect -5050 27396 -5034 27430
rect -5134 27358 -5034 27396
rect -4976 27430 -4876 27446
rect -4976 27396 -4960 27430
rect -4892 27396 -4876 27430
rect -4976 27358 -4876 27396
rect -4818 27430 -4718 27446
rect -4818 27396 -4802 27430
rect -4734 27396 -4718 27430
rect -4818 27358 -4718 27396
rect -4660 27430 -4560 27446
rect -4660 27396 -4644 27430
rect -4576 27396 -4560 27430
rect -4660 27358 -4560 27396
rect -4502 27430 -4402 27446
rect -4502 27396 -4486 27430
rect -4418 27396 -4402 27430
rect -4502 27358 -4402 27396
rect -4344 27430 -4244 27446
rect -4344 27396 -4328 27430
rect -4260 27396 -4244 27430
rect -4344 27358 -4244 27396
rect -4186 27430 -4086 27446
rect -4186 27396 -4170 27430
rect -4102 27396 -4086 27430
rect -4186 27358 -4086 27396
rect -4028 27430 -3928 27446
rect -4028 27396 -4012 27430
rect -3944 27396 -3928 27430
rect -4028 27358 -3928 27396
rect -3870 27430 -3770 27446
rect -3870 27396 -3854 27430
rect -3786 27396 -3770 27430
rect -3870 27358 -3770 27396
rect -3712 27430 -3612 27446
rect -3712 27396 -3696 27430
rect -3628 27396 -3612 27430
rect -3712 27358 -3612 27396
rect -3554 27430 -3454 27446
rect -3554 27396 -3538 27430
rect -3470 27396 -3454 27430
rect -3554 27358 -3454 27396
rect -3396 27430 -3296 27446
rect -3396 27396 -3380 27430
rect -3312 27396 -3296 27430
rect -3396 27358 -3296 27396
rect -3238 27430 -3138 27446
rect -3238 27396 -3222 27430
rect -3154 27396 -3138 27430
rect -3238 27358 -3138 27396
rect -3080 27430 -2980 27446
rect -3080 27396 -3064 27430
rect -2996 27396 -2980 27430
rect -3080 27358 -2980 27396
rect -2922 27430 -2822 27446
rect -2922 27396 -2906 27430
rect -2838 27396 -2822 27430
rect -2922 27358 -2822 27396
rect -2764 27430 -2664 27446
rect -2764 27396 -2748 27430
rect -2680 27396 -2664 27430
rect -2764 27358 -2664 27396
rect -2606 27430 -2506 27446
rect -2606 27396 -2590 27430
rect -2522 27396 -2506 27430
rect -2606 27358 -2506 27396
rect -2448 27430 -2348 27446
rect -2448 27396 -2432 27430
rect -2364 27396 -2348 27430
rect -2448 27358 -2348 27396
rect -2290 27430 -2190 27446
rect -2290 27396 -2274 27430
rect -2206 27396 -2190 27430
rect -2290 27358 -2190 27396
rect -6872 21320 -6772 21358
rect -6872 21286 -6856 21320
rect -6788 21286 -6772 21320
rect -6872 21270 -6772 21286
rect -6714 21320 -6614 21358
rect -6714 21286 -6698 21320
rect -6630 21286 -6614 21320
rect -6714 21270 -6614 21286
rect -6556 21320 -6456 21358
rect -6556 21286 -6540 21320
rect -6472 21286 -6456 21320
rect -6556 21270 -6456 21286
rect -6398 21320 -6298 21358
rect -6398 21286 -6382 21320
rect -6314 21286 -6298 21320
rect -6398 21270 -6298 21286
rect -6240 21320 -6140 21358
rect -6240 21286 -6224 21320
rect -6156 21286 -6140 21320
rect -6240 21270 -6140 21286
rect -6082 21320 -5982 21358
rect -6082 21286 -6066 21320
rect -5998 21286 -5982 21320
rect -6082 21270 -5982 21286
rect -5924 21320 -5824 21358
rect -5924 21286 -5908 21320
rect -5840 21286 -5824 21320
rect -5924 21270 -5824 21286
rect -5766 21320 -5666 21358
rect -5766 21286 -5750 21320
rect -5682 21286 -5666 21320
rect -5766 21270 -5666 21286
rect -5608 21320 -5508 21358
rect -5608 21286 -5592 21320
rect -5524 21286 -5508 21320
rect -5608 21270 -5508 21286
rect -5450 21320 -5350 21358
rect -5450 21286 -5434 21320
rect -5366 21286 -5350 21320
rect -5450 21270 -5350 21286
rect -5292 21320 -5192 21358
rect -5292 21286 -5276 21320
rect -5208 21286 -5192 21320
rect -5292 21270 -5192 21286
rect -5134 21320 -5034 21358
rect -5134 21286 -5118 21320
rect -5050 21286 -5034 21320
rect -5134 21270 -5034 21286
rect -4976 21320 -4876 21358
rect -4976 21286 -4960 21320
rect -4892 21286 -4876 21320
rect -4976 21270 -4876 21286
rect -4818 21320 -4718 21358
rect -4818 21286 -4802 21320
rect -4734 21286 -4718 21320
rect -4818 21270 -4718 21286
rect -4660 21320 -4560 21358
rect -4660 21286 -4644 21320
rect -4576 21286 -4560 21320
rect -4660 21270 -4560 21286
rect -4502 21320 -4402 21358
rect -4502 21286 -4486 21320
rect -4418 21286 -4402 21320
rect -4502 21270 -4402 21286
rect -4344 21320 -4244 21358
rect -4344 21286 -4328 21320
rect -4260 21286 -4244 21320
rect -4344 21270 -4244 21286
rect -4186 21320 -4086 21358
rect -4186 21286 -4170 21320
rect -4102 21286 -4086 21320
rect -4186 21270 -4086 21286
rect -4028 21320 -3928 21358
rect -4028 21286 -4012 21320
rect -3944 21286 -3928 21320
rect -4028 21270 -3928 21286
rect -3870 21320 -3770 21358
rect -3870 21286 -3854 21320
rect -3786 21286 -3770 21320
rect -3870 21270 -3770 21286
rect -3712 21320 -3612 21358
rect -3712 21286 -3696 21320
rect -3628 21286 -3612 21320
rect -3712 21270 -3612 21286
rect -3554 21320 -3454 21358
rect -3554 21286 -3538 21320
rect -3470 21286 -3454 21320
rect -3554 21270 -3454 21286
rect -3396 21320 -3296 21358
rect -3396 21286 -3380 21320
rect -3312 21286 -3296 21320
rect -3396 21270 -3296 21286
rect -3238 21320 -3138 21358
rect -3238 21286 -3222 21320
rect -3154 21286 -3138 21320
rect -3238 21270 -3138 21286
rect -3080 21320 -2980 21358
rect -3080 21286 -3064 21320
rect -2996 21286 -2980 21320
rect -3080 21270 -2980 21286
rect -2922 21320 -2822 21358
rect -2922 21286 -2906 21320
rect -2838 21286 -2822 21320
rect -2922 21270 -2822 21286
rect -2764 21320 -2664 21358
rect -2764 21286 -2748 21320
rect -2680 21286 -2664 21320
rect -2764 21270 -2664 21286
rect -2606 21320 -2506 21358
rect -2606 21286 -2590 21320
rect -2522 21286 -2506 21320
rect -2606 21270 -2506 21286
rect -2448 21320 -2348 21358
rect -2448 21286 -2432 21320
rect -2364 21286 -2348 21320
rect -2448 21270 -2348 21286
rect -2290 21320 -2190 21358
rect -2290 21286 -2274 21320
rect -2206 21286 -2190 21320
rect -2290 21270 -2190 21286
rect -572 27430 -472 27446
rect -572 27396 -556 27430
rect -488 27396 -472 27430
rect -572 27358 -472 27396
rect -414 27430 -314 27446
rect -414 27396 -398 27430
rect -330 27396 -314 27430
rect -414 27358 -314 27396
rect -256 27430 -156 27446
rect -256 27396 -240 27430
rect -172 27396 -156 27430
rect -256 27358 -156 27396
rect -98 27430 2 27446
rect -98 27396 -82 27430
rect -14 27396 2 27430
rect -98 27358 2 27396
rect 60 27430 160 27446
rect 60 27396 76 27430
rect 144 27396 160 27430
rect 60 27358 160 27396
rect 218 27430 318 27446
rect 218 27396 234 27430
rect 302 27396 318 27430
rect 218 27358 318 27396
rect 376 27430 476 27446
rect 376 27396 392 27430
rect 460 27396 476 27430
rect 376 27358 476 27396
rect 534 27430 634 27446
rect 534 27396 550 27430
rect 618 27396 634 27430
rect 534 27358 634 27396
rect 692 27430 792 27446
rect 692 27396 708 27430
rect 776 27396 792 27430
rect 692 27358 792 27396
rect 850 27430 950 27446
rect 850 27396 866 27430
rect 934 27396 950 27430
rect 850 27358 950 27396
rect 1008 27430 1108 27446
rect 1008 27396 1024 27430
rect 1092 27396 1108 27430
rect 1008 27358 1108 27396
rect 1166 27430 1266 27446
rect 1166 27396 1182 27430
rect 1250 27396 1266 27430
rect 1166 27358 1266 27396
rect 1324 27430 1424 27446
rect 1324 27396 1340 27430
rect 1408 27396 1424 27430
rect 1324 27358 1424 27396
rect 1482 27430 1582 27446
rect 1482 27396 1498 27430
rect 1566 27396 1582 27430
rect 1482 27358 1582 27396
rect 1640 27430 1740 27446
rect 1640 27396 1656 27430
rect 1724 27396 1740 27430
rect 1640 27358 1740 27396
rect 1798 27430 1898 27446
rect 1798 27396 1814 27430
rect 1882 27396 1898 27430
rect 1798 27358 1898 27396
rect 1956 27430 2056 27446
rect 1956 27396 1972 27430
rect 2040 27396 2056 27430
rect 1956 27358 2056 27396
rect 2114 27430 2214 27446
rect 2114 27396 2130 27430
rect 2198 27396 2214 27430
rect 2114 27358 2214 27396
rect 2272 27430 2372 27446
rect 2272 27396 2288 27430
rect 2356 27396 2372 27430
rect 2272 27358 2372 27396
rect 2430 27430 2530 27446
rect 2430 27396 2446 27430
rect 2514 27396 2530 27430
rect 2430 27358 2530 27396
rect 2588 27430 2688 27446
rect 2588 27396 2604 27430
rect 2672 27396 2688 27430
rect 2588 27358 2688 27396
rect 2746 27430 2846 27446
rect 2746 27396 2762 27430
rect 2830 27396 2846 27430
rect 2746 27358 2846 27396
rect 2904 27430 3004 27446
rect 2904 27396 2920 27430
rect 2988 27396 3004 27430
rect 2904 27358 3004 27396
rect 3062 27430 3162 27446
rect 3062 27396 3078 27430
rect 3146 27396 3162 27430
rect 3062 27358 3162 27396
rect 3220 27430 3320 27446
rect 3220 27396 3236 27430
rect 3304 27396 3320 27430
rect 3220 27358 3320 27396
rect 3378 27430 3478 27446
rect 3378 27396 3394 27430
rect 3462 27396 3478 27430
rect 3378 27358 3478 27396
rect 3536 27430 3636 27446
rect 3536 27396 3552 27430
rect 3620 27396 3636 27430
rect 3536 27358 3636 27396
rect 3694 27430 3794 27446
rect 3694 27396 3710 27430
rect 3778 27396 3794 27430
rect 3694 27358 3794 27396
rect 3852 27430 3952 27446
rect 3852 27396 3868 27430
rect 3936 27396 3952 27430
rect 3852 27358 3952 27396
rect 4010 27430 4110 27446
rect 4010 27396 4026 27430
rect 4094 27396 4110 27430
rect 4010 27358 4110 27396
rect -572 21320 -472 21358
rect -572 21286 -556 21320
rect -488 21286 -472 21320
rect -572 21270 -472 21286
rect -414 21320 -314 21358
rect -414 21286 -398 21320
rect -330 21286 -314 21320
rect -414 21270 -314 21286
rect -256 21320 -156 21358
rect -256 21286 -240 21320
rect -172 21286 -156 21320
rect -256 21270 -156 21286
rect -98 21320 2 21358
rect -98 21286 -82 21320
rect -14 21286 2 21320
rect -98 21270 2 21286
rect 60 21320 160 21358
rect 60 21286 76 21320
rect 144 21286 160 21320
rect 60 21270 160 21286
rect 218 21320 318 21358
rect 218 21286 234 21320
rect 302 21286 318 21320
rect 218 21270 318 21286
rect 376 21320 476 21358
rect 376 21286 392 21320
rect 460 21286 476 21320
rect 376 21270 476 21286
rect 534 21320 634 21358
rect 534 21286 550 21320
rect 618 21286 634 21320
rect 534 21270 634 21286
rect 692 21320 792 21358
rect 692 21286 708 21320
rect 776 21286 792 21320
rect 692 21270 792 21286
rect 850 21320 950 21358
rect 850 21286 866 21320
rect 934 21286 950 21320
rect 850 21270 950 21286
rect 1008 21320 1108 21358
rect 1008 21286 1024 21320
rect 1092 21286 1108 21320
rect 1008 21270 1108 21286
rect 1166 21320 1266 21358
rect 1166 21286 1182 21320
rect 1250 21286 1266 21320
rect 1166 21270 1266 21286
rect 1324 21320 1424 21358
rect 1324 21286 1340 21320
rect 1408 21286 1424 21320
rect 1324 21270 1424 21286
rect 1482 21320 1582 21358
rect 1482 21286 1498 21320
rect 1566 21286 1582 21320
rect 1482 21270 1582 21286
rect 1640 21320 1740 21358
rect 1640 21286 1656 21320
rect 1724 21286 1740 21320
rect 1640 21270 1740 21286
rect 1798 21320 1898 21358
rect 1798 21286 1814 21320
rect 1882 21286 1898 21320
rect 1798 21270 1898 21286
rect 1956 21320 2056 21358
rect 1956 21286 1972 21320
rect 2040 21286 2056 21320
rect 1956 21270 2056 21286
rect 2114 21320 2214 21358
rect 2114 21286 2130 21320
rect 2198 21286 2214 21320
rect 2114 21270 2214 21286
rect 2272 21320 2372 21358
rect 2272 21286 2288 21320
rect 2356 21286 2372 21320
rect 2272 21270 2372 21286
rect 2430 21320 2530 21358
rect 2430 21286 2446 21320
rect 2514 21286 2530 21320
rect 2430 21270 2530 21286
rect 2588 21320 2688 21358
rect 2588 21286 2604 21320
rect 2672 21286 2688 21320
rect 2588 21270 2688 21286
rect 2746 21320 2846 21358
rect 2746 21286 2762 21320
rect 2830 21286 2846 21320
rect 2746 21270 2846 21286
rect 2904 21320 3004 21358
rect 2904 21286 2920 21320
rect 2988 21286 3004 21320
rect 2904 21270 3004 21286
rect 3062 21320 3162 21358
rect 3062 21286 3078 21320
rect 3146 21286 3162 21320
rect 3062 21270 3162 21286
rect 3220 21320 3320 21358
rect 3220 21286 3236 21320
rect 3304 21286 3320 21320
rect 3220 21270 3320 21286
rect 3378 21320 3478 21358
rect 3378 21286 3394 21320
rect 3462 21286 3478 21320
rect 3378 21270 3478 21286
rect 3536 21320 3636 21358
rect 3536 21286 3552 21320
rect 3620 21286 3636 21320
rect 3536 21270 3636 21286
rect 3694 21320 3794 21358
rect 3694 21286 3710 21320
rect 3778 21286 3794 21320
rect 3694 21270 3794 21286
rect 3852 21320 3952 21358
rect 3852 21286 3868 21320
rect 3936 21286 3952 21320
rect 3852 21270 3952 21286
rect 4010 21320 4110 21358
rect 4010 21286 4026 21320
rect 4094 21286 4110 21320
rect 4010 21270 4110 21286
rect 5728 27430 5828 27446
rect 5728 27396 5744 27430
rect 5812 27396 5828 27430
rect 5728 27358 5828 27396
rect 5886 27430 5986 27446
rect 5886 27396 5902 27430
rect 5970 27396 5986 27430
rect 5886 27358 5986 27396
rect 6044 27430 6144 27446
rect 6044 27396 6060 27430
rect 6128 27396 6144 27430
rect 6044 27358 6144 27396
rect 6202 27430 6302 27446
rect 6202 27396 6218 27430
rect 6286 27396 6302 27430
rect 6202 27358 6302 27396
rect 6360 27430 6460 27446
rect 6360 27396 6376 27430
rect 6444 27396 6460 27430
rect 6360 27358 6460 27396
rect 6518 27430 6618 27446
rect 6518 27396 6534 27430
rect 6602 27396 6618 27430
rect 6518 27358 6618 27396
rect 6676 27430 6776 27446
rect 6676 27396 6692 27430
rect 6760 27396 6776 27430
rect 6676 27358 6776 27396
rect 6834 27430 6934 27446
rect 6834 27396 6850 27430
rect 6918 27396 6934 27430
rect 6834 27358 6934 27396
rect 6992 27430 7092 27446
rect 6992 27396 7008 27430
rect 7076 27396 7092 27430
rect 6992 27358 7092 27396
rect 7150 27430 7250 27446
rect 7150 27396 7166 27430
rect 7234 27396 7250 27430
rect 7150 27358 7250 27396
rect 7308 27430 7408 27446
rect 7308 27396 7324 27430
rect 7392 27396 7408 27430
rect 7308 27358 7408 27396
rect 7466 27430 7566 27446
rect 7466 27396 7482 27430
rect 7550 27396 7566 27430
rect 7466 27358 7566 27396
rect 7624 27430 7724 27446
rect 7624 27396 7640 27430
rect 7708 27396 7724 27430
rect 7624 27358 7724 27396
rect 7782 27430 7882 27446
rect 7782 27396 7798 27430
rect 7866 27396 7882 27430
rect 7782 27358 7882 27396
rect 7940 27430 8040 27446
rect 7940 27396 7956 27430
rect 8024 27396 8040 27430
rect 7940 27358 8040 27396
rect 8098 27430 8198 27446
rect 8098 27396 8114 27430
rect 8182 27396 8198 27430
rect 8098 27358 8198 27396
rect 8256 27430 8356 27446
rect 8256 27396 8272 27430
rect 8340 27396 8356 27430
rect 8256 27358 8356 27396
rect 8414 27430 8514 27446
rect 8414 27396 8430 27430
rect 8498 27396 8514 27430
rect 8414 27358 8514 27396
rect 8572 27430 8672 27446
rect 8572 27396 8588 27430
rect 8656 27396 8672 27430
rect 8572 27358 8672 27396
rect 8730 27430 8830 27446
rect 8730 27396 8746 27430
rect 8814 27396 8830 27430
rect 8730 27358 8830 27396
rect 8888 27430 8988 27446
rect 8888 27396 8904 27430
rect 8972 27396 8988 27430
rect 8888 27358 8988 27396
rect 9046 27430 9146 27446
rect 9046 27396 9062 27430
rect 9130 27396 9146 27430
rect 9046 27358 9146 27396
rect 9204 27430 9304 27446
rect 9204 27396 9220 27430
rect 9288 27396 9304 27430
rect 9204 27358 9304 27396
rect 9362 27430 9462 27446
rect 9362 27396 9378 27430
rect 9446 27396 9462 27430
rect 9362 27358 9462 27396
rect 9520 27430 9620 27446
rect 9520 27396 9536 27430
rect 9604 27396 9620 27430
rect 9520 27358 9620 27396
rect 9678 27430 9778 27446
rect 9678 27396 9694 27430
rect 9762 27396 9778 27430
rect 9678 27358 9778 27396
rect 9836 27430 9936 27446
rect 9836 27396 9852 27430
rect 9920 27396 9936 27430
rect 9836 27358 9936 27396
rect 9994 27430 10094 27446
rect 9994 27396 10010 27430
rect 10078 27396 10094 27430
rect 9994 27358 10094 27396
rect 10152 27430 10252 27446
rect 10152 27396 10168 27430
rect 10236 27396 10252 27430
rect 10152 27358 10252 27396
rect 10310 27430 10410 27446
rect 10310 27396 10326 27430
rect 10394 27396 10410 27430
rect 10310 27358 10410 27396
rect 5728 21320 5828 21358
rect 5728 21286 5744 21320
rect 5812 21286 5828 21320
rect 5728 21270 5828 21286
rect 5886 21320 5986 21358
rect 5886 21286 5902 21320
rect 5970 21286 5986 21320
rect 5886 21270 5986 21286
rect 6044 21320 6144 21358
rect 6044 21286 6060 21320
rect 6128 21286 6144 21320
rect 6044 21270 6144 21286
rect 6202 21320 6302 21358
rect 6202 21286 6218 21320
rect 6286 21286 6302 21320
rect 6202 21270 6302 21286
rect 6360 21320 6460 21358
rect 6360 21286 6376 21320
rect 6444 21286 6460 21320
rect 6360 21270 6460 21286
rect 6518 21320 6618 21358
rect 6518 21286 6534 21320
rect 6602 21286 6618 21320
rect 6518 21270 6618 21286
rect 6676 21320 6776 21358
rect 6676 21286 6692 21320
rect 6760 21286 6776 21320
rect 6676 21270 6776 21286
rect 6834 21320 6934 21358
rect 6834 21286 6850 21320
rect 6918 21286 6934 21320
rect 6834 21270 6934 21286
rect 6992 21320 7092 21358
rect 6992 21286 7008 21320
rect 7076 21286 7092 21320
rect 6992 21270 7092 21286
rect 7150 21320 7250 21358
rect 7150 21286 7166 21320
rect 7234 21286 7250 21320
rect 7150 21270 7250 21286
rect 7308 21320 7408 21358
rect 7308 21286 7324 21320
rect 7392 21286 7408 21320
rect 7308 21270 7408 21286
rect 7466 21320 7566 21358
rect 7466 21286 7482 21320
rect 7550 21286 7566 21320
rect 7466 21270 7566 21286
rect 7624 21320 7724 21358
rect 7624 21286 7640 21320
rect 7708 21286 7724 21320
rect 7624 21270 7724 21286
rect 7782 21320 7882 21358
rect 7782 21286 7798 21320
rect 7866 21286 7882 21320
rect 7782 21270 7882 21286
rect 7940 21320 8040 21358
rect 7940 21286 7956 21320
rect 8024 21286 8040 21320
rect 7940 21270 8040 21286
rect 8098 21320 8198 21358
rect 8098 21286 8114 21320
rect 8182 21286 8198 21320
rect 8098 21270 8198 21286
rect 8256 21320 8356 21358
rect 8256 21286 8272 21320
rect 8340 21286 8356 21320
rect 8256 21270 8356 21286
rect 8414 21320 8514 21358
rect 8414 21286 8430 21320
rect 8498 21286 8514 21320
rect 8414 21270 8514 21286
rect 8572 21320 8672 21358
rect 8572 21286 8588 21320
rect 8656 21286 8672 21320
rect 8572 21270 8672 21286
rect 8730 21320 8830 21358
rect 8730 21286 8746 21320
rect 8814 21286 8830 21320
rect 8730 21270 8830 21286
rect 8888 21320 8988 21358
rect 8888 21286 8904 21320
rect 8972 21286 8988 21320
rect 8888 21270 8988 21286
rect 9046 21320 9146 21358
rect 9046 21286 9062 21320
rect 9130 21286 9146 21320
rect 9046 21270 9146 21286
rect 9204 21320 9304 21358
rect 9204 21286 9220 21320
rect 9288 21286 9304 21320
rect 9204 21270 9304 21286
rect 9362 21320 9462 21358
rect 9362 21286 9378 21320
rect 9446 21286 9462 21320
rect 9362 21270 9462 21286
rect 9520 21320 9620 21358
rect 9520 21286 9536 21320
rect 9604 21286 9620 21320
rect 9520 21270 9620 21286
rect 9678 21320 9778 21358
rect 9678 21286 9694 21320
rect 9762 21286 9778 21320
rect 9678 21270 9778 21286
rect 9836 21320 9936 21358
rect 9836 21286 9852 21320
rect 9920 21286 9936 21320
rect 9836 21270 9936 21286
rect 9994 21320 10094 21358
rect 9994 21286 10010 21320
rect 10078 21286 10094 21320
rect 9994 21270 10094 21286
rect 10152 21320 10252 21358
rect 10152 21286 10168 21320
rect 10236 21286 10252 21320
rect 10152 21270 10252 21286
rect 10310 21320 10410 21358
rect 10310 21286 10326 21320
rect 10394 21286 10410 21320
rect 10310 21270 10410 21286
rect -13172 19130 -13072 19146
rect -13172 19096 -13156 19130
rect -13088 19096 -13072 19130
rect -13172 19058 -13072 19096
rect -13014 19130 -12914 19146
rect -13014 19096 -12998 19130
rect -12930 19096 -12914 19130
rect -13014 19058 -12914 19096
rect -12856 19130 -12756 19146
rect -12856 19096 -12840 19130
rect -12772 19096 -12756 19130
rect -12856 19058 -12756 19096
rect -12698 19130 -12598 19146
rect -12698 19096 -12682 19130
rect -12614 19096 -12598 19130
rect -12698 19058 -12598 19096
rect -12540 19130 -12440 19146
rect -12540 19096 -12524 19130
rect -12456 19096 -12440 19130
rect -12540 19058 -12440 19096
rect -12382 19130 -12282 19146
rect -12382 19096 -12366 19130
rect -12298 19096 -12282 19130
rect -12382 19058 -12282 19096
rect -12224 19130 -12124 19146
rect -12224 19096 -12208 19130
rect -12140 19096 -12124 19130
rect -12224 19058 -12124 19096
rect -12066 19130 -11966 19146
rect -12066 19096 -12050 19130
rect -11982 19096 -11966 19130
rect -12066 19058 -11966 19096
rect -11908 19130 -11808 19146
rect -11908 19096 -11892 19130
rect -11824 19096 -11808 19130
rect -11908 19058 -11808 19096
rect -11750 19130 -11650 19146
rect -11750 19096 -11734 19130
rect -11666 19096 -11650 19130
rect -11750 19058 -11650 19096
rect -11592 19130 -11492 19146
rect -11592 19096 -11576 19130
rect -11508 19096 -11492 19130
rect -11592 19058 -11492 19096
rect -11434 19130 -11334 19146
rect -11434 19096 -11418 19130
rect -11350 19096 -11334 19130
rect -11434 19058 -11334 19096
rect -11276 19130 -11176 19146
rect -11276 19096 -11260 19130
rect -11192 19096 -11176 19130
rect -11276 19058 -11176 19096
rect -11118 19130 -11018 19146
rect -11118 19096 -11102 19130
rect -11034 19096 -11018 19130
rect -11118 19058 -11018 19096
rect -10960 19130 -10860 19146
rect -10960 19096 -10944 19130
rect -10876 19096 -10860 19130
rect -10960 19058 -10860 19096
rect -10802 19130 -10702 19146
rect -10802 19096 -10786 19130
rect -10718 19096 -10702 19130
rect -10802 19058 -10702 19096
rect -10644 19130 -10544 19146
rect -10644 19096 -10628 19130
rect -10560 19096 -10544 19130
rect -10644 19058 -10544 19096
rect -10486 19130 -10386 19146
rect -10486 19096 -10470 19130
rect -10402 19096 -10386 19130
rect -10486 19058 -10386 19096
rect -10328 19130 -10228 19146
rect -10328 19096 -10312 19130
rect -10244 19096 -10228 19130
rect -10328 19058 -10228 19096
rect -10170 19130 -10070 19146
rect -10170 19096 -10154 19130
rect -10086 19096 -10070 19130
rect -10170 19058 -10070 19096
rect -10012 19130 -9912 19146
rect -10012 19096 -9996 19130
rect -9928 19096 -9912 19130
rect -10012 19058 -9912 19096
rect -9854 19130 -9754 19146
rect -9854 19096 -9838 19130
rect -9770 19096 -9754 19130
rect -9854 19058 -9754 19096
rect -9696 19130 -9596 19146
rect -9696 19096 -9680 19130
rect -9612 19096 -9596 19130
rect -9696 19058 -9596 19096
rect -9538 19130 -9438 19146
rect -9538 19096 -9522 19130
rect -9454 19096 -9438 19130
rect -9538 19058 -9438 19096
rect -9380 19130 -9280 19146
rect -9380 19096 -9364 19130
rect -9296 19096 -9280 19130
rect -9380 19058 -9280 19096
rect -9222 19130 -9122 19146
rect -9222 19096 -9206 19130
rect -9138 19096 -9122 19130
rect -9222 19058 -9122 19096
rect -9064 19130 -8964 19146
rect -9064 19096 -9048 19130
rect -8980 19096 -8964 19130
rect -9064 19058 -8964 19096
rect -8906 19130 -8806 19146
rect -8906 19096 -8890 19130
rect -8822 19096 -8806 19130
rect -8906 19058 -8806 19096
rect -8748 19130 -8648 19146
rect -8748 19096 -8732 19130
rect -8664 19096 -8648 19130
rect -8748 19058 -8648 19096
rect -8590 19130 -8490 19146
rect -8590 19096 -8574 19130
rect -8506 19096 -8490 19130
rect -8590 19058 -8490 19096
rect -13172 13020 -13072 13058
rect -13172 12986 -13156 13020
rect -13088 12986 -13072 13020
rect -13172 12970 -13072 12986
rect -13014 13020 -12914 13058
rect -13014 12986 -12998 13020
rect -12930 12986 -12914 13020
rect -13014 12970 -12914 12986
rect -12856 13020 -12756 13058
rect -12856 12986 -12840 13020
rect -12772 12986 -12756 13020
rect -12856 12970 -12756 12986
rect -12698 13020 -12598 13058
rect -12698 12986 -12682 13020
rect -12614 12986 -12598 13020
rect -12698 12970 -12598 12986
rect -12540 13020 -12440 13058
rect -12540 12986 -12524 13020
rect -12456 12986 -12440 13020
rect -12540 12970 -12440 12986
rect -12382 13020 -12282 13058
rect -12382 12986 -12366 13020
rect -12298 12986 -12282 13020
rect -12382 12970 -12282 12986
rect -12224 13020 -12124 13058
rect -12224 12986 -12208 13020
rect -12140 12986 -12124 13020
rect -12224 12970 -12124 12986
rect -12066 13020 -11966 13058
rect -12066 12986 -12050 13020
rect -11982 12986 -11966 13020
rect -12066 12970 -11966 12986
rect -11908 13020 -11808 13058
rect -11908 12986 -11892 13020
rect -11824 12986 -11808 13020
rect -11908 12970 -11808 12986
rect -11750 13020 -11650 13058
rect -11750 12986 -11734 13020
rect -11666 12986 -11650 13020
rect -11750 12970 -11650 12986
rect -11592 13020 -11492 13058
rect -11592 12986 -11576 13020
rect -11508 12986 -11492 13020
rect -11592 12970 -11492 12986
rect -11434 13020 -11334 13058
rect -11434 12986 -11418 13020
rect -11350 12986 -11334 13020
rect -11434 12970 -11334 12986
rect -11276 13020 -11176 13058
rect -11276 12986 -11260 13020
rect -11192 12986 -11176 13020
rect -11276 12970 -11176 12986
rect -11118 13020 -11018 13058
rect -11118 12986 -11102 13020
rect -11034 12986 -11018 13020
rect -11118 12970 -11018 12986
rect -10960 13020 -10860 13058
rect -10960 12986 -10944 13020
rect -10876 12986 -10860 13020
rect -10960 12970 -10860 12986
rect -10802 13020 -10702 13058
rect -10802 12986 -10786 13020
rect -10718 12986 -10702 13020
rect -10802 12970 -10702 12986
rect -10644 13020 -10544 13058
rect -10644 12986 -10628 13020
rect -10560 12986 -10544 13020
rect -10644 12970 -10544 12986
rect -10486 13020 -10386 13058
rect -10486 12986 -10470 13020
rect -10402 12986 -10386 13020
rect -10486 12970 -10386 12986
rect -10328 13020 -10228 13058
rect -10328 12986 -10312 13020
rect -10244 12986 -10228 13020
rect -10328 12970 -10228 12986
rect -10170 13020 -10070 13058
rect -10170 12986 -10154 13020
rect -10086 12986 -10070 13020
rect -10170 12970 -10070 12986
rect -10012 13020 -9912 13058
rect -10012 12986 -9996 13020
rect -9928 12986 -9912 13020
rect -10012 12970 -9912 12986
rect -9854 13020 -9754 13058
rect -9854 12986 -9838 13020
rect -9770 12986 -9754 13020
rect -9854 12970 -9754 12986
rect -9696 13020 -9596 13058
rect -9696 12986 -9680 13020
rect -9612 12986 -9596 13020
rect -9696 12970 -9596 12986
rect -9538 13020 -9438 13058
rect -9538 12986 -9522 13020
rect -9454 12986 -9438 13020
rect -9538 12970 -9438 12986
rect -9380 13020 -9280 13058
rect -9380 12986 -9364 13020
rect -9296 12986 -9280 13020
rect -9380 12970 -9280 12986
rect -9222 13020 -9122 13058
rect -9222 12986 -9206 13020
rect -9138 12986 -9122 13020
rect -9222 12970 -9122 12986
rect -9064 13020 -8964 13058
rect -9064 12986 -9048 13020
rect -8980 12986 -8964 13020
rect -9064 12970 -8964 12986
rect -8906 13020 -8806 13058
rect -8906 12986 -8890 13020
rect -8822 12986 -8806 13020
rect -8906 12970 -8806 12986
rect -8748 13020 -8648 13058
rect -8748 12986 -8732 13020
rect -8664 12986 -8648 13020
rect -8748 12970 -8648 12986
rect -8590 13020 -8490 13058
rect -8590 12986 -8574 13020
rect -8506 12986 -8490 13020
rect -8590 12970 -8490 12986
rect -6872 19130 -6772 19146
rect -6872 19096 -6856 19130
rect -6788 19096 -6772 19130
rect -6872 19058 -6772 19096
rect -6714 19130 -6614 19146
rect -6714 19096 -6698 19130
rect -6630 19096 -6614 19130
rect -6714 19058 -6614 19096
rect -6556 19130 -6456 19146
rect -6556 19096 -6540 19130
rect -6472 19096 -6456 19130
rect -6556 19058 -6456 19096
rect -6398 19130 -6298 19146
rect -6398 19096 -6382 19130
rect -6314 19096 -6298 19130
rect -6398 19058 -6298 19096
rect -6240 19130 -6140 19146
rect -6240 19096 -6224 19130
rect -6156 19096 -6140 19130
rect -6240 19058 -6140 19096
rect -6082 19130 -5982 19146
rect -6082 19096 -6066 19130
rect -5998 19096 -5982 19130
rect -6082 19058 -5982 19096
rect -5924 19130 -5824 19146
rect -5924 19096 -5908 19130
rect -5840 19096 -5824 19130
rect -5924 19058 -5824 19096
rect -5766 19130 -5666 19146
rect -5766 19096 -5750 19130
rect -5682 19096 -5666 19130
rect -5766 19058 -5666 19096
rect -5608 19130 -5508 19146
rect -5608 19096 -5592 19130
rect -5524 19096 -5508 19130
rect -5608 19058 -5508 19096
rect -5450 19130 -5350 19146
rect -5450 19096 -5434 19130
rect -5366 19096 -5350 19130
rect -5450 19058 -5350 19096
rect -5292 19130 -5192 19146
rect -5292 19096 -5276 19130
rect -5208 19096 -5192 19130
rect -5292 19058 -5192 19096
rect -5134 19130 -5034 19146
rect -5134 19096 -5118 19130
rect -5050 19096 -5034 19130
rect -5134 19058 -5034 19096
rect -4976 19130 -4876 19146
rect -4976 19096 -4960 19130
rect -4892 19096 -4876 19130
rect -4976 19058 -4876 19096
rect -4818 19130 -4718 19146
rect -4818 19096 -4802 19130
rect -4734 19096 -4718 19130
rect -4818 19058 -4718 19096
rect -4660 19130 -4560 19146
rect -4660 19096 -4644 19130
rect -4576 19096 -4560 19130
rect -4660 19058 -4560 19096
rect -4502 19130 -4402 19146
rect -4502 19096 -4486 19130
rect -4418 19096 -4402 19130
rect -4502 19058 -4402 19096
rect -4344 19130 -4244 19146
rect -4344 19096 -4328 19130
rect -4260 19096 -4244 19130
rect -4344 19058 -4244 19096
rect -4186 19130 -4086 19146
rect -4186 19096 -4170 19130
rect -4102 19096 -4086 19130
rect -4186 19058 -4086 19096
rect -4028 19130 -3928 19146
rect -4028 19096 -4012 19130
rect -3944 19096 -3928 19130
rect -4028 19058 -3928 19096
rect -3870 19130 -3770 19146
rect -3870 19096 -3854 19130
rect -3786 19096 -3770 19130
rect -3870 19058 -3770 19096
rect -3712 19130 -3612 19146
rect -3712 19096 -3696 19130
rect -3628 19096 -3612 19130
rect -3712 19058 -3612 19096
rect -3554 19130 -3454 19146
rect -3554 19096 -3538 19130
rect -3470 19096 -3454 19130
rect -3554 19058 -3454 19096
rect -3396 19130 -3296 19146
rect -3396 19096 -3380 19130
rect -3312 19096 -3296 19130
rect -3396 19058 -3296 19096
rect -3238 19130 -3138 19146
rect -3238 19096 -3222 19130
rect -3154 19096 -3138 19130
rect -3238 19058 -3138 19096
rect -3080 19130 -2980 19146
rect -3080 19096 -3064 19130
rect -2996 19096 -2980 19130
rect -3080 19058 -2980 19096
rect -2922 19130 -2822 19146
rect -2922 19096 -2906 19130
rect -2838 19096 -2822 19130
rect -2922 19058 -2822 19096
rect -2764 19130 -2664 19146
rect -2764 19096 -2748 19130
rect -2680 19096 -2664 19130
rect -2764 19058 -2664 19096
rect -2606 19130 -2506 19146
rect -2606 19096 -2590 19130
rect -2522 19096 -2506 19130
rect -2606 19058 -2506 19096
rect -2448 19130 -2348 19146
rect -2448 19096 -2432 19130
rect -2364 19096 -2348 19130
rect -2448 19058 -2348 19096
rect -2290 19130 -2190 19146
rect -2290 19096 -2274 19130
rect -2206 19096 -2190 19130
rect -2290 19058 -2190 19096
rect -6872 13020 -6772 13058
rect -6872 12986 -6856 13020
rect -6788 12986 -6772 13020
rect -6872 12970 -6772 12986
rect -6714 13020 -6614 13058
rect -6714 12986 -6698 13020
rect -6630 12986 -6614 13020
rect -6714 12970 -6614 12986
rect -6556 13020 -6456 13058
rect -6556 12986 -6540 13020
rect -6472 12986 -6456 13020
rect -6556 12970 -6456 12986
rect -6398 13020 -6298 13058
rect -6398 12986 -6382 13020
rect -6314 12986 -6298 13020
rect -6398 12970 -6298 12986
rect -6240 13020 -6140 13058
rect -6240 12986 -6224 13020
rect -6156 12986 -6140 13020
rect -6240 12970 -6140 12986
rect -6082 13020 -5982 13058
rect -6082 12986 -6066 13020
rect -5998 12986 -5982 13020
rect -6082 12970 -5982 12986
rect -5924 13020 -5824 13058
rect -5924 12986 -5908 13020
rect -5840 12986 -5824 13020
rect -5924 12970 -5824 12986
rect -5766 13020 -5666 13058
rect -5766 12986 -5750 13020
rect -5682 12986 -5666 13020
rect -5766 12970 -5666 12986
rect -5608 13020 -5508 13058
rect -5608 12986 -5592 13020
rect -5524 12986 -5508 13020
rect -5608 12970 -5508 12986
rect -5450 13020 -5350 13058
rect -5450 12986 -5434 13020
rect -5366 12986 -5350 13020
rect -5450 12970 -5350 12986
rect -5292 13020 -5192 13058
rect -5292 12986 -5276 13020
rect -5208 12986 -5192 13020
rect -5292 12970 -5192 12986
rect -5134 13020 -5034 13058
rect -5134 12986 -5118 13020
rect -5050 12986 -5034 13020
rect -5134 12970 -5034 12986
rect -4976 13020 -4876 13058
rect -4976 12986 -4960 13020
rect -4892 12986 -4876 13020
rect -4976 12970 -4876 12986
rect -4818 13020 -4718 13058
rect -4818 12986 -4802 13020
rect -4734 12986 -4718 13020
rect -4818 12970 -4718 12986
rect -4660 13020 -4560 13058
rect -4660 12986 -4644 13020
rect -4576 12986 -4560 13020
rect -4660 12970 -4560 12986
rect -4502 13020 -4402 13058
rect -4502 12986 -4486 13020
rect -4418 12986 -4402 13020
rect -4502 12970 -4402 12986
rect -4344 13020 -4244 13058
rect -4344 12986 -4328 13020
rect -4260 12986 -4244 13020
rect -4344 12970 -4244 12986
rect -4186 13020 -4086 13058
rect -4186 12986 -4170 13020
rect -4102 12986 -4086 13020
rect -4186 12970 -4086 12986
rect -4028 13020 -3928 13058
rect -4028 12986 -4012 13020
rect -3944 12986 -3928 13020
rect -4028 12970 -3928 12986
rect -3870 13020 -3770 13058
rect -3870 12986 -3854 13020
rect -3786 12986 -3770 13020
rect -3870 12970 -3770 12986
rect -3712 13020 -3612 13058
rect -3712 12986 -3696 13020
rect -3628 12986 -3612 13020
rect -3712 12970 -3612 12986
rect -3554 13020 -3454 13058
rect -3554 12986 -3538 13020
rect -3470 12986 -3454 13020
rect -3554 12970 -3454 12986
rect -3396 13020 -3296 13058
rect -3396 12986 -3380 13020
rect -3312 12986 -3296 13020
rect -3396 12970 -3296 12986
rect -3238 13020 -3138 13058
rect -3238 12986 -3222 13020
rect -3154 12986 -3138 13020
rect -3238 12970 -3138 12986
rect -3080 13020 -2980 13058
rect -3080 12986 -3064 13020
rect -2996 12986 -2980 13020
rect -3080 12970 -2980 12986
rect -2922 13020 -2822 13058
rect -2922 12986 -2906 13020
rect -2838 12986 -2822 13020
rect -2922 12970 -2822 12986
rect -2764 13020 -2664 13058
rect -2764 12986 -2748 13020
rect -2680 12986 -2664 13020
rect -2764 12970 -2664 12986
rect -2606 13020 -2506 13058
rect -2606 12986 -2590 13020
rect -2522 12986 -2506 13020
rect -2606 12970 -2506 12986
rect -2448 13020 -2348 13058
rect -2448 12986 -2432 13020
rect -2364 12986 -2348 13020
rect -2448 12970 -2348 12986
rect -2290 13020 -2190 13058
rect -2290 12986 -2274 13020
rect -2206 12986 -2190 13020
rect -2290 12970 -2190 12986
rect -572 19130 -472 19146
rect -572 19096 -556 19130
rect -488 19096 -472 19130
rect -572 19058 -472 19096
rect -414 19130 -314 19146
rect -414 19096 -398 19130
rect -330 19096 -314 19130
rect -414 19058 -314 19096
rect -256 19130 -156 19146
rect -256 19096 -240 19130
rect -172 19096 -156 19130
rect -256 19058 -156 19096
rect -98 19130 2 19146
rect -98 19096 -82 19130
rect -14 19096 2 19130
rect -98 19058 2 19096
rect 60 19130 160 19146
rect 60 19096 76 19130
rect 144 19096 160 19130
rect 60 19058 160 19096
rect 218 19130 318 19146
rect 218 19096 234 19130
rect 302 19096 318 19130
rect 218 19058 318 19096
rect 376 19130 476 19146
rect 376 19096 392 19130
rect 460 19096 476 19130
rect 376 19058 476 19096
rect 534 19130 634 19146
rect 534 19096 550 19130
rect 618 19096 634 19130
rect 534 19058 634 19096
rect 692 19130 792 19146
rect 692 19096 708 19130
rect 776 19096 792 19130
rect 692 19058 792 19096
rect 850 19130 950 19146
rect 850 19096 866 19130
rect 934 19096 950 19130
rect 850 19058 950 19096
rect 1008 19130 1108 19146
rect 1008 19096 1024 19130
rect 1092 19096 1108 19130
rect 1008 19058 1108 19096
rect 1166 19130 1266 19146
rect 1166 19096 1182 19130
rect 1250 19096 1266 19130
rect 1166 19058 1266 19096
rect 1324 19130 1424 19146
rect 1324 19096 1340 19130
rect 1408 19096 1424 19130
rect 1324 19058 1424 19096
rect 1482 19130 1582 19146
rect 1482 19096 1498 19130
rect 1566 19096 1582 19130
rect 1482 19058 1582 19096
rect 1640 19130 1740 19146
rect 1640 19096 1656 19130
rect 1724 19096 1740 19130
rect 1640 19058 1740 19096
rect 1798 19130 1898 19146
rect 1798 19096 1814 19130
rect 1882 19096 1898 19130
rect 1798 19058 1898 19096
rect 1956 19130 2056 19146
rect 1956 19096 1972 19130
rect 2040 19096 2056 19130
rect 1956 19058 2056 19096
rect 2114 19130 2214 19146
rect 2114 19096 2130 19130
rect 2198 19096 2214 19130
rect 2114 19058 2214 19096
rect 2272 19130 2372 19146
rect 2272 19096 2288 19130
rect 2356 19096 2372 19130
rect 2272 19058 2372 19096
rect 2430 19130 2530 19146
rect 2430 19096 2446 19130
rect 2514 19096 2530 19130
rect 2430 19058 2530 19096
rect 2588 19130 2688 19146
rect 2588 19096 2604 19130
rect 2672 19096 2688 19130
rect 2588 19058 2688 19096
rect 2746 19130 2846 19146
rect 2746 19096 2762 19130
rect 2830 19096 2846 19130
rect 2746 19058 2846 19096
rect 2904 19130 3004 19146
rect 2904 19096 2920 19130
rect 2988 19096 3004 19130
rect 2904 19058 3004 19096
rect 3062 19130 3162 19146
rect 3062 19096 3078 19130
rect 3146 19096 3162 19130
rect 3062 19058 3162 19096
rect 3220 19130 3320 19146
rect 3220 19096 3236 19130
rect 3304 19096 3320 19130
rect 3220 19058 3320 19096
rect 3378 19130 3478 19146
rect 3378 19096 3394 19130
rect 3462 19096 3478 19130
rect 3378 19058 3478 19096
rect 3536 19130 3636 19146
rect 3536 19096 3552 19130
rect 3620 19096 3636 19130
rect 3536 19058 3636 19096
rect 3694 19130 3794 19146
rect 3694 19096 3710 19130
rect 3778 19096 3794 19130
rect 3694 19058 3794 19096
rect 3852 19130 3952 19146
rect 3852 19096 3868 19130
rect 3936 19096 3952 19130
rect 3852 19058 3952 19096
rect 4010 19130 4110 19146
rect 4010 19096 4026 19130
rect 4094 19096 4110 19130
rect 4010 19058 4110 19096
rect -572 13020 -472 13058
rect -572 12986 -556 13020
rect -488 12986 -472 13020
rect -572 12970 -472 12986
rect -414 13020 -314 13058
rect -414 12986 -398 13020
rect -330 12986 -314 13020
rect -414 12970 -314 12986
rect -256 13020 -156 13058
rect -256 12986 -240 13020
rect -172 12986 -156 13020
rect -256 12970 -156 12986
rect -98 13020 2 13058
rect -98 12986 -82 13020
rect -14 12986 2 13020
rect -98 12970 2 12986
rect 60 13020 160 13058
rect 60 12986 76 13020
rect 144 12986 160 13020
rect 60 12970 160 12986
rect 218 13020 318 13058
rect 218 12986 234 13020
rect 302 12986 318 13020
rect 218 12970 318 12986
rect 376 13020 476 13058
rect 376 12986 392 13020
rect 460 12986 476 13020
rect 376 12970 476 12986
rect 534 13020 634 13058
rect 534 12986 550 13020
rect 618 12986 634 13020
rect 534 12970 634 12986
rect 692 13020 792 13058
rect 692 12986 708 13020
rect 776 12986 792 13020
rect 692 12970 792 12986
rect 850 13020 950 13058
rect 850 12986 866 13020
rect 934 12986 950 13020
rect 850 12970 950 12986
rect 1008 13020 1108 13058
rect 1008 12986 1024 13020
rect 1092 12986 1108 13020
rect 1008 12970 1108 12986
rect 1166 13020 1266 13058
rect 1166 12986 1182 13020
rect 1250 12986 1266 13020
rect 1166 12970 1266 12986
rect 1324 13020 1424 13058
rect 1324 12986 1340 13020
rect 1408 12986 1424 13020
rect 1324 12970 1424 12986
rect 1482 13020 1582 13058
rect 1482 12986 1498 13020
rect 1566 12986 1582 13020
rect 1482 12970 1582 12986
rect 1640 13020 1740 13058
rect 1640 12986 1656 13020
rect 1724 12986 1740 13020
rect 1640 12970 1740 12986
rect 1798 13020 1898 13058
rect 1798 12986 1814 13020
rect 1882 12986 1898 13020
rect 1798 12970 1898 12986
rect 1956 13020 2056 13058
rect 1956 12986 1972 13020
rect 2040 12986 2056 13020
rect 1956 12970 2056 12986
rect 2114 13020 2214 13058
rect 2114 12986 2130 13020
rect 2198 12986 2214 13020
rect 2114 12970 2214 12986
rect 2272 13020 2372 13058
rect 2272 12986 2288 13020
rect 2356 12986 2372 13020
rect 2272 12970 2372 12986
rect 2430 13020 2530 13058
rect 2430 12986 2446 13020
rect 2514 12986 2530 13020
rect 2430 12970 2530 12986
rect 2588 13020 2688 13058
rect 2588 12986 2604 13020
rect 2672 12986 2688 13020
rect 2588 12970 2688 12986
rect 2746 13020 2846 13058
rect 2746 12986 2762 13020
rect 2830 12986 2846 13020
rect 2746 12970 2846 12986
rect 2904 13020 3004 13058
rect 2904 12986 2920 13020
rect 2988 12986 3004 13020
rect 2904 12970 3004 12986
rect 3062 13020 3162 13058
rect 3062 12986 3078 13020
rect 3146 12986 3162 13020
rect 3062 12970 3162 12986
rect 3220 13020 3320 13058
rect 3220 12986 3236 13020
rect 3304 12986 3320 13020
rect 3220 12970 3320 12986
rect 3378 13020 3478 13058
rect 3378 12986 3394 13020
rect 3462 12986 3478 13020
rect 3378 12970 3478 12986
rect 3536 13020 3636 13058
rect 3536 12986 3552 13020
rect 3620 12986 3636 13020
rect 3536 12970 3636 12986
rect 3694 13020 3794 13058
rect 3694 12986 3710 13020
rect 3778 12986 3794 13020
rect 3694 12970 3794 12986
rect 3852 13020 3952 13058
rect 3852 12986 3868 13020
rect 3936 12986 3952 13020
rect 3852 12970 3952 12986
rect 4010 13020 4110 13058
rect 4010 12986 4026 13020
rect 4094 12986 4110 13020
rect 4010 12970 4110 12986
rect 5728 19130 5828 19146
rect 5728 19096 5744 19130
rect 5812 19096 5828 19130
rect 5728 19058 5828 19096
rect 5886 19130 5986 19146
rect 5886 19096 5902 19130
rect 5970 19096 5986 19130
rect 5886 19058 5986 19096
rect 6044 19130 6144 19146
rect 6044 19096 6060 19130
rect 6128 19096 6144 19130
rect 6044 19058 6144 19096
rect 6202 19130 6302 19146
rect 6202 19096 6218 19130
rect 6286 19096 6302 19130
rect 6202 19058 6302 19096
rect 6360 19130 6460 19146
rect 6360 19096 6376 19130
rect 6444 19096 6460 19130
rect 6360 19058 6460 19096
rect 6518 19130 6618 19146
rect 6518 19096 6534 19130
rect 6602 19096 6618 19130
rect 6518 19058 6618 19096
rect 6676 19130 6776 19146
rect 6676 19096 6692 19130
rect 6760 19096 6776 19130
rect 6676 19058 6776 19096
rect 6834 19130 6934 19146
rect 6834 19096 6850 19130
rect 6918 19096 6934 19130
rect 6834 19058 6934 19096
rect 6992 19130 7092 19146
rect 6992 19096 7008 19130
rect 7076 19096 7092 19130
rect 6992 19058 7092 19096
rect 7150 19130 7250 19146
rect 7150 19096 7166 19130
rect 7234 19096 7250 19130
rect 7150 19058 7250 19096
rect 7308 19130 7408 19146
rect 7308 19096 7324 19130
rect 7392 19096 7408 19130
rect 7308 19058 7408 19096
rect 7466 19130 7566 19146
rect 7466 19096 7482 19130
rect 7550 19096 7566 19130
rect 7466 19058 7566 19096
rect 7624 19130 7724 19146
rect 7624 19096 7640 19130
rect 7708 19096 7724 19130
rect 7624 19058 7724 19096
rect 7782 19130 7882 19146
rect 7782 19096 7798 19130
rect 7866 19096 7882 19130
rect 7782 19058 7882 19096
rect 7940 19130 8040 19146
rect 7940 19096 7956 19130
rect 8024 19096 8040 19130
rect 7940 19058 8040 19096
rect 8098 19130 8198 19146
rect 8098 19096 8114 19130
rect 8182 19096 8198 19130
rect 8098 19058 8198 19096
rect 8256 19130 8356 19146
rect 8256 19096 8272 19130
rect 8340 19096 8356 19130
rect 8256 19058 8356 19096
rect 8414 19130 8514 19146
rect 8414 19096 8430 19130
rect 8498 19096 8514 19130
rect 8414 19058 8514 19096
rect 8572 19130 8672 19146
rect 8572 19096 8588 19130
rect 8656 19096 8672 19130
rect 8572 19058 8672 19096
rect 8730 19130 8830 19146
rect 8730 19096 8746 19130
rect 8814 19096 8830 19130
rect 8730 19058 8830 19096
rect 8888 19130 8988 19146
rect 8888 19096 8904 19130
rect 8972 19096 8988 19130
rect 8888 19058 8988 19096
rect 9046 19130 9146 19146
rect 9046 19096 9062 19130
rect 9130 19096 9146 19130
rect 9046 19058 9146 19096
rect 9204 19130 9304 19146
rect 9204 19096 9220 19130
rect 9288 19096 9304 19130
rect 9204 19058 9304 19096
rect 9362 19130 9462 19146
rect 9362 19096 9378 19130
rect 9446 19096 9462 19130
rect 9362 19058 9462 19096
rect 9520 19130 9620 19146
rect 9520 19096 9536 19130
rect 9604 19096 9620 19130
rect 9520 19058 9620 19096
rect 9678 19130 9778 19146
rect 9678 19096 9694 19130
rect 9762 19096 9778 19130
rect 9678 19058 9778 19096
rect 9836 19130 9936 19146
rect 9836 19096 9852 19130
rect 9920 19096 9936 19130
rect 9836 19058 9936 19096
rect 9994 19130 10094 19146
rect 9994 19096 10010 19130
rect 10078 19096 10094 19130
rect 9994 19058 10094 19096
rect 10152 19130 10252 19146
rect 10152 19096 10168 19130
rect 10236 19096 10252 19130
rect 10152 19058 10252 19096
rect 10310 19130 10410 19146
rect 10310 19096 10326 19130
rect 10394 19096 10410 19130
rect 10310 19058 10410 19096
rect 5728 13020 5828 13058
rect 5728 12986 5744 13020
rect 5812 12986 5828 13020
rect 5728 12970 5828 12986
rect 5886 13020 5986 13058
rect 5886 12986 5902 13020
rect 5970 12986 5986 13020
rect 5886 12970 5986 12986
rect 6044 13020 6144 13058
rect 6044 12986 6060 13020
rect 6128 12986 6144 13020
rect 6044 12970 6144 12986
rect 6202 13020 6302 13058
rect 6202 12986 6218 13020
rect 6286 12986 6302 13020
rect 6202 12970 6302 12986
rect 6360 13020 6460 13058
rect 6360 12986 6376 13020
rect 6444 12986 6460 13020
rect 6360 12970 6460 12986
rect 6518 13020 6618 13058
rect 6518 12986 6534 13020
rect 6602 12986 6618 13020
rect 6518 12970 6618 12986
rect 6676 13020 6776 13058
rect 6676 12986 6692 13020
rect 6760 12986 6776 13020
rect 6676 12970 6776 12986
rect 6834 13020 6934 13058
rect 6834 12986 6850 13020
rect 6918 12986 6934 13020
rect 6834 12970 6934 12986
rect 6992 13020 7092 13058
rect 6992 12986 7008 13020
rect 7076 12986 7092 13020
rect 6992 12970 7092 12986
rect 7150 13020 7250 13058
rect 7150 12986 7166 13020
rect 7234 12986 7250 13020
rect 7150 12970 7250 12986
rect 7308 13020 7408 13058
rect 7308 12986 7324 13020
rect 7392 12986 7408 13020
rect 7308 12970 7408 12986
rect 7466 13020 7566 13058
rect 7466 12986 7482 13020
rect 7550 12986 7566 13020
rect 7466 12970 7566 12986
rect 7624 13020 7724 13058
rect 7624 12986 7640 13020
rect 7708 12986 7724 13020
rect 7624 12970 7724 12986
rect 7782 13020 7882 13058
rect 7782 12986 7798 13020
rect 7866 12986 7882 13020
rect 7782 12970 7882 12986
rect 7940 13020 8040 13058
rect 7940 12986 7956 13020
rect 8024 12986 8040 13020
rect 7940 12970 8040 12986
rect 8098 13020 8198 13058
rect 8098 12986 8114 13020
rect 8182 12986 8198 13020
rect 8098 12970 8198 12986
rect 8256 13020 8356 13058
rect 8256 12986 8272 13020
rect 8340 12986 8356 13020
rect 8256 12970 8356 12986
rect 8414 13020 8514 13058
rect 8414 12986 8430 13020
rect 8498 12986 8514 13020
rect 8414 12970 8514 12986
rect 8572 13020 8672 13058
rect 8572 12986 8588 13020
rect 8656 12986 8672 13020
rect 8572 12970 8672 12986
rect 8730 13020 8830 13058
rect 8730 12986 8746 13020
rect 8814 12986 8830 13020
rect 8730 12970 8830 12986
rect 8888 13020 8988 13058
rect 8888 12986 8904 13020
rect 8972 12986 8988 13020
rect 8888 12970 8988 12986
rect 9046 13020 9146 13058
rect 9046 12986 9062 13020
rect 9130 12986 9146 13020
rect 9046 12970 9146 12986
rect 9204 13020 9304 13058
rect 9204 12986 9220 13020
rect 9288 12986 9304 13020
rect 9204 12970 9304 12986
rect 9362 13020 9462 13058
rect 9362 12986 9378 13020
rect 9446 12986 9462 13020
rect 9362 12970 9462 12986
rect 9520 13020 9620 13058
rect 9520 12986 9536 13020
rect 9604 12986 9620 13020
rect 9520 12970 9620 12986
rect 9678 13020 9778 13058
rect 9678 12986 9694 13020
rect 9762 12986 9778 13020
rect 9678 12970 9778 12986
rect 9836 13020 9936 13058
rect 9836 12986 9852 13020
rect 9920 12986 9936 13020
rect 9836 12970 9936 12986
rect 9994 13020 10094 13058
rect 9994 12986 10010 13020
rect 10078 12986 10094 13020
rect 9994 12970 10094 12986
rect 10152 13020 10252 13058
rect 10152 12986 10168 13020
rect 10236 12986 10252 13020
rect 10152 12970 10252 12986
rect 10310 13020 10410 13058
rect 10310 12986 10326 13020
rect 10394 12986 10410 13020
rect 10310 12970 10410 12986
rect -13172 12130 -13072 12146
rect -13172 12096 -13156 12130
rect -13088 12096 -13072 12130
rect -13172 12058 -13072 12096
rect -13014 12130 -12914 12146
rect -13014 12096 -12998 12130
rect -12930 12096 -12914 12130
rect -13014 12058 -12914 12096
rect -12856 12130 -12756 12146
rect -12856 12096 -12840 12130
rect -12772 12096 -12756 12130
rect -12856 12058 -12756 12096
rect -12698 12130 -12598 12146
rect -12698 12096 -12682 12130
rect -12614 12096 -12598 12130
rect -12698 12058 -12598 12096
rect -12540 12130 -12440 12146
rect -12540 12096 -12524 12130
rect -12456 12096 -12440 12130
rect -12540 12058 -12440 12096
rect -12382 12130 -12282 12146
rect -12382 12096 -12366 12130
rect -12298 12096 -12282 12130
rect -12382 12058 -12282 12096
rect -12224 12130 -12124 12146
rect -12224 12096 -12208 12130
rect -12140 12096 -12124 12130
rect -12224 12058 -12124 12096
rect -12066 12130 -11966 12146
rect -12066 12096 -12050 12130
rect -11982 12096 -11966 12130
rect -12066 12058 -11966 12096
rect -11908 12130 -11808 12146
rect -11908 12096 -11892 12130
rect -11824 12096 -11808 12130
rect -11908 12058 -11808 12096
rect -11750 12130 -11650 12146
rect -11750 12096 -11734 12130
rect -11666 12096 -11650 12130
rect -11750 12058 -11650 12096
rect -11592 12130 -11492 12146
rect -11592 12096 -11576 12130
rect -11508 12096 -11492 12130
rect -11592 12058 -11492 12096
rect -11434 12130 -11334 12146
rect -11434 12096 -11418 12130
rect -11350 12096 -11334 12130
rect -11434 12058 -11334 12096
rect -11276 12130 -11176 12146
rect -11276 12096 -11260 12130
rect -11192 12096 -11176 12130
rect -11276 12058 -11176 12096
rect -11118 12130 -11018 12146
rect -11118 12096 -11102 12130
rect -11034 12096 -11018 12130
rect -11118 12058 -11018 12096
rect -10960 12130 -10860 12146
rect -10960 12096 -10944 12130
rect -10876 12096 -10860 12130
rect -10960 12058 -10860 12096
rect -10802 12130 -10702 12146
rect -10802 12096 -10786 12130
rect -10718 12096 -10702 12130
rect -10802 12058 -10702 12096
rect -10644 12130 -10544 12146
rect -10644 12096 -10628 12130
rect -10560 12096 -10544 12130
rect -10644 12058 -10544 12096
rect -10486 12130 -10386 12146
rect -10486 12096 -10470 12130
rect -10402 12096 -10386 12130
rect -10486 12058 -10386 12096
rect -10328 12130 -10228 12146
rect -10328 12096 -10312 12130
rect -10244 12096 -10228 12130
rect -10328 12058 -10228 12096
rect -10170 12130 -10070 12146
rect -10170 12096 -10154 12130
rect -10086 12096 -10070 12130
rect -10170 12058 -10070 12096
rect -10012 12130 -9912 12146
rect -10012 12096 -9996 12130
rect -9928 12096 -9912 12130
rect -10012 12058 -9912 12096
rect -9854 12130 -9754 12146
rect -9854 12096 -9838 12130
rect -9770 12096 -9754 12130
rect -9854 12058 -9754 12096
rect -9696 12130 -9596 12146
rect -9696 12096 -9680 12130
rect -9612 12096 -9596 12130
rect -9696 12058 -9596 12096
rect -9538 12130 -9438 12146
rect -9538 12096 -9522 12130
rect -9454 12096 -9438 12130
rect -9538 12058 -9438 12096
rect -9380 12130 -9280 12146
rect -9380 12096 -9364 12130
rect -9296 12096 -9280 12130
rect -9380 12058 -9280 12096
rect -9222 12130 -9122 12146
rect -9222 12096 -9206 12130
rect -9138 12096 -9122 12130
rect -9222 12058 -9122 12096
rect -9064 12130 -8964 12146
rect -9064 12096 -9048 12130
rect -8980 12096 -8964 12130
rect -9064 12058 -8964 12096
rect -8906 12130 -8806 12146
rect -8906 12096 -8890 12130
rect -8822 12096 -8806 12130
rect -8906 12058 -8806 12096
rect -8748 12130 -8648 12146
rect -8748 12096 -8732 12130
rect -8664 12096 -8648 12130
rect -8748 12058 -8648 12096
rect -8590 12130 -8490 12146
rect -8590 12096 -8574 12130
rect -8506 12096 -8490 12130
rect -8590 12058 -8490 12096
rect -13172 6020 -13072 6058
rect -13172 5986 -13156 6020
rect -13088 5986 -13072 6020
rect -13172 5970 -13072 5986
rect -13014 6020 -12914 6058
rect -13014 5986 -12998 6020
rect -12930 5986 -12914 6020
rect -13014 5970 -12914 5986
rect -12856 6020 -12756 6058
rect -12856 5986 -12840 6020
rect -12772 5986 -12756 6020
rect -12856 5970 -12756 5986
rect -12698 6020 -12598 6058
rect -12698 5986 -12682 6020
rect -12614 5986 -12598 6020
rect -12698 5970 -12598 5986
rect -12540 6020 -12440 6058
rect -12540 5986 -12524 6020
rect -12456 5986 -12440 6020
rect -12540 5970 -12440 5986
rect -12382 6020 -12282 6058
rect -12382 5986 -12366 6020
rect -12298 5986 -12282 6020
rect -12382 5970 -12282 5986
rect -12224 6020 -12124 6058
rect -12224 5986 -12208 6020
rect -12140 5986 -12124 6020
rect -12224 5970 -12124 5986
rect -12066 6020 -11966 6058
rect -12066 5986 -12050 6020
rect -11982 5986 -11966 6020
rect -12066 5970 -11966 5986
rect -11908 6020 -11808 6058
rect -11908 5986 -11892 6020
rect -11824 5986 -11808 6020
rect -11908 5970 -11808 5986
rect -11750 6020 -11650 6058
rect -11750 5986 -11734 6020
rect -11666 5986 -11650 6020
rect -11750 5970 -11650 5986
rect -11592 6020 -11492 6058
rect -11592 5986 -11576 6020
rect -11508 5986 -11492 6020
rect -11592 5970 -11492 5986
rect -11434 6020 -11334 6058
rect -11434 5986 -11418 6020
rect -11350 5986 -11334 6020
rect -11434 5970 -11334 5986
rect -11276 6020 -11176 6058
rect -11276 5986 -11260 6020
rect -11192 5986 -11176 6020
rect -11276 5970 -11176 5986
rect -11118 6020 -11018 6058
rect -11118 5986 -11102 6020
rect -11034 5986 -11018 6020
rect -11118 5970 -11018 5986
rect -10960 6020 -10860 6058
rect -10960 5986 -10944 6020
rect -10876 5986 -10860 6020
rect -10960 5970 -10860 5986
rect -10802 6020 -10702 6058
rect -10802 5986 -10786 6020
rect -10718 5986 -10702 6020
rect -10802 5970 -10702 5986
rect -10644 6020 -10544 6058
rect -10644 5986 -10628 6020
rect -10560 5986 -10544 6020
rect -10644 5970 -10544 5986
rect -10486 6020 -10386 6058
rect -10486 5986 -10470 6020
rect -10402 5986 -10386 6020
rect -10486 5970 -10386 5986
rect -10328 6020 -10228 6058
rect -10328 5986 -10312 6020
rect -10244 5986 -10228 6020
rect -10328 5970 -10228 5986
rect -10170 6020 -10070 6058
rect -10170 5986 -10154 6020
rect -10086 5986 -10070 6020
rect -10170 5970 -10070 5986
rect -10012 6020 -9912 6058
rect -10012 5986 -9996 6020
rect -9928 5986 -9912 6020
rect -10012 5970 -9912 5986
rect -9854 6020 -9754 6058
rect -9854 5986 -9838 6020
rect -9770 5986 -9754 6020
rect -9854 5970 -9754 5986
rect -9696 6020 -9596 6058
rect -9696 5986 -9680 6020
rect -9612 5986 -9596 6020
rect -9696 5970 -9596 5986
rect -9538 6020 -9438 6058
rect -9538 5986 -9522 6020
rect -9454 5986 -9438 6020
rect -9538 5970 -9438 5986
rect -9380 6020 -9280 6058
rect -9380 5986 -9364 6020
rect -9296 5986 -9280 6020
rect -9380 5970 -9280 5986
rect -9222 6020 -9122 6058
rect -9222 5986 -9206 6020
rect -9138 5986 -9122 6020
rect -9222 5970 -9122 5986
rect -9064 6020 -8964 6058
rect -9064 5986 -9048 6020
rect -8980 5986 -8964 6020
rect -9064 5970 -8964 5986
rect -8906 6020 -8806 6058
rect -8906 5986 -8890 6020
rect -8822 5986 -8806 6020
rect -8906 5970 -8806 5986
rect -8748 6020 -8648 6058
rect -8748 5986 -8732 6020
rect -8664 5986 -8648 6020
rect -8748 5970 -8648 5986
rect -8590 6020 -8490 6058
rect -8590 5986 -8574 6020
rect -8506 5986 -8490 6020
rect -8590 5970 -8490 5986
rect -6872 12130 -6772 12146
rect -6872 12096 -6856 12130
rect -6788 12096 -6772 12130
rect -6872 12058 -6772 12096
rect -6714 12130 -6614 12146
rect -6714 12096 -6698 12130
rect -6630 12096 -6614 12130
rect -6714 12058 -6614 12096
rect -6556 12130 -6456 12146
rect -6556 12096 -6540 12130
rect -6472 12096 -6456 12130
rect -6556 12058 -6456 12096
rect -6398 12130 -6298 12146
rect -6398 12096 -6382 12130
rect -6314 12096 -6298 12130
rect -6398 12058 -6298 12096
rect -6240 12130 -6140 12146
rect -6240 12096 -6224 12130
rect -6156 12096 -6140 12130
rect -6240 12058 -6140 12096
rect -6082 12130 -5982 12146
rect -6082 12096 -6066 12130
rect -5998 12096 -5982 12130
rect -6082 12058 -5982 12096
rect -5924 12130 -5824 12146
rect -5924 12096 -5908 12130
rect -5840 12096 -5824 12130
rect -5924 12058 -5824 12096
rect -5766 12130 -5666 12146
rect -5766 12096 -5750 12130
rect -5682 12096 -5666 12130
rect -5766 12058 -5666 12096
rect -5608 12130 -5508 12146
rect -5608 12096 -5592 12130
rect -5524 12096 -5508 12130
rect -5608 12058 -5508 12096
rect -5450 12130 -5350 12146
rect -5450 12096 -5434 12130
rect -5366 12096 -5350 12130
rect -5450 12058 -5350 12096
rect -5292 12130 -5192 12146
rect -5292 12096 -5276 12130
rect -5208 12096 -5192 12130
rect -5292 12058 -5192 12096
rect -5134 12130 -5034 12146
rect -5134 12096 -5118 12130
rect -5050 12096 -5034 12130
rect -5134 12058 -5034 12096
rect -4976 12130 -4876 12146
rect -4976 12096 -4960 12130
rect -4892 12096 -4876 12130
rect -4976 12058 -4876 12096
rect -4818 12130 -4718 12146
rect -4818 12096 -4802 12130
rect -4734 12096 -4718 12130
rect -4818 12058 -4718 12096
rect -4660 12130 -4560 12146
rect -4660 12096 -4644 12130
rect -4576 12096 -4560 12130
rect -4660 12058 -4560 12096
rect -4502 12130 -4402 12146
rect -4502 12096 -4486 12130
rect -4418 12096 -4402 12130
rect -4502 12058 -4402 12096
rect -4344 12130 -4244 12146
rect -4344 12096 -4328 12130
rect -4260 12096 -4244 12130
rect -4344 12058 -4244 12096
rect -4186 12130 -4086 12146
rect -4186 12096 -4170 12130
rect -4102 12096 -4086 12130
rect -4186 12058 -4086 12096
rect -4028 12130 -3928 12146
rect -4028 12096 -4012 12130
rect -3944 12096 -3928 12130
rect -4028 12058 -3928 12096
rect -3870 12130 -3770 12146
rect -3870 12096 -3854 12130
rect -3786 12096 -3770 12130
rect -3870 12058 -3770 12096
rect -3712 12130 -3612 12146
rect -3712 12096 -3696 12130
rect -3628 12096 -3612 12130
rect -3712 12058 -3612 12096
rect -3554 12130 -3454 12146
rect -3554 12096 -3538 12130
rect -3470 12096 -3454 12130
rect -3554 12058 -3454 12096
rect -3396 12130 -3296 12146
rect -3396 12096 -3380 12130
rect -3312 12096 -3296 12130
rect -3396 12058 -3296 12096
rect -3238 12130 -3138 12146
rect -3238 12096 -3222 12130
rect -3154 12096 -3138 12130
rect -3238 12058 -3138 12096
rect -3080 12130 -2980 12146
rect -3080 12096 -3064 12130
rect -2996 12096 -2980 12130
rect -3080 12058 -2980 12096
rect -2922 12130 -2822 12146
rect -2922 12096 -2906 12130
rect -2838 12096 -2822 12130
rect -2922 12058 -2822 12096
rect -2764 12130 -2664 12146
rect -2764 12096 -2748 12130
rect -2680 12096 -2664 12130
rect -2764 12058 -2664 12096
rect -2606 12130 -2506 12146
rect -2606 12096 -2590 12130
rect -2522 12096 -2506 12130
rect -2606 12058 -2506 12096
rect -2448 12130 -2348 12146
rect -2448 12096 -2432 12130
rect -2364 12096 -2348 12130
rect -2448 12058 -2348 12096
rect -2290 12130 -2190 12146
rect -2290 12096 -2274 12130
rect -2206 12096 -2190 12130
rect -2290 12058 -2190 12096
rect -6872 6020 -6772 6058
rect -6872 5986 -6856 6020
rect -6788 5986 -6772 6020
rect -6872 5970 -6772 5986
rect -6714 6020 -6614 6058
rect -6714 5986 -6698 6020
rect -6630 5986 -6614 6020
rect -6714 5970 -6614 5986
rect -6556 6020 -6456 6058
rect -6556 5986 -6540 6020
rect -6472 5986 -6456 6020
rect -6556 5970 -6456 5986
rect -6398 6020 -6298 6058
rect -6398 5986 -6382 6020
rect -6314 5986 -6298 6020
rect -6398 5970 -6298 5986
rect -6240 6020 -6140 6058
rect -6240 5986 -6224 6020
rect -6156 5986 -6140 6020
rect -6240 5970 -6140 5986
rect -6082 6020 -5982 6058
rect -6082 5986 -6066 6020
rect -5998 5986 -5982 6020
rect -6082 5970 -5982 5986
rect -5924 6020 -5824 6058
rect -5924 5986 -5908 6020
rect -5840 5986 -5824 6020
rect -5924 5970 -5824 5986
rect -5766 6020 -5666 6058
rect -5766 5986 -5750 6020
rect -5682 5986 -5666 6020
rect -5766 5970 -5666 5986
rect -5608 6020 -5508 6058
rect -5608 5986 -5592 6020
rect -5524 5986 -5508 6020
rect -5608 5970 -5508 5986
rect -5450 6020 -5350 6058
rect -5450 5986 -5434 6020
rect -5366 5986 -5350 6020
rect -5450 5970 -5350 5986
rect -5292 6020 -5192 6058
rect -5292 5986 -5276 6020
rect -5208 5986 -5192 6020
rect -5292 5970 -5192 5986
rect -5134 6020 -5034 6058
rect -5134 5986 -5118 6020
rect -5050 5986 -5034 6020
rect -5134 5970 -5034 5986
rect -4976 6020 -4876 6058
rect -4976 5986 -4960 6020
rect -4892 5986 -4876 6020
rect -4976 5970 -4876 5986
rect -4818 6020 -4718 6058
rect -4818 5986 -4802 6020
rect -4734 5986 -4718 6020
rect -4818 5970 -4718 5986
rect -4660 6020 -4560 6058
rect -4660 5986 -4644 6020
rect -4576 5986 -4560 6020
rect -4660 5970 -4560 5986
rect -4502 6020 -4402 6058
rect -4502 5986 -4486 6020
rect -4418 5986 -4402 6020
rect -4502 5970 -4402 5986
rect -4344 6020 -4244 6058
rect -4344 5986 -4328 6020
rect -4260 5986 -4244 6020
rect -4344 5970 -4244 5986
rect -4186 6020 -4086 6058
rect -4186 5986 -4170 6020
rect -4102 5986 -4086 6020
rect -4186 5970 -4086 5986
rect -4028 6020 -3928 6058
rect -4028 5986 -4012 6020
rect -3944 5986 -3928 6020
rect -4028 5970 -3928 5986
rect -3870 6020 -3770 6058
rect -3870 5986 -3854 6020
rect -3786 5986 -3770 6020
rect -3870 5970 -3770 5986
rect -3712 6020 -3612 6058
rect -3712 5986 -3696 6020
rect -3628 5986 -3612 6020
rect -3712 5970 -3612 5986
rect -3554 6020 -3454 6058
rect -3554 5986 -3538 6020
rect -3470 5986 -3454 6020
rect -3554 5970 -3454 5986
rect -3396 6020 -3296 6058
rect -3396 5986 -3380 6020
rect -3312 5986 -3296 6020
rect -3396 5970 -3296 5986
rect -3238 6020 -3138 6058
rect -3238 5986 -3222 6020
rect -3154 5986 -3138 6020
rect -3238 5970 -3138 5986
rect -3080 6020 -2980 6058
rect -3080 5986 -3064 6020
rect -2996 5986 -2980 6020
rect -3080 5970 -2980 5986
rect -2922 6020 -2822 6058
rect -2922 5986 -2906 6020
rect -2838 5986 -2822 6020
rect -2922 5970 -2822 5986
rect -2764 6020 -2664 6058
rect -2764 5986 -2748 6020
rect -2680 5986 -2664 6020
rect -2764 5970 -2664 5986
rect -2606 6020 -2506 6058
rect -2606 5986 -2590 6020
rect -2522 5986 -2506 6020
rect -2606 5970 -2506 5986
rect -2448 6020 -2348 6058
rect -2448 5986 -2432 6020
rect -2364 5986 -2348 6020
rect -2448 5970 -2348 5986
rect -2290 6020 -2190 6058
rect -2290 5986 -2274 6020
rect -2206 5986 -2190 6020
rect -2290 5970 -2190 5986
rect -572 12130 -472 12146
rect -572 12096 -556 12130
rect -488 12096 -472 12130
rect -572 12058 -472 12096
rect -414 12130 -314 12146
rect -414 12096 -398 12130
rect -330 12096 -314 12130
rect -414 12058 -314 12096
rect -256 12130 -156 12146
rect -256 12096 -240 12130
rect -172 12096 -156 12130
rect -256 12058 -156 12096
rect -98 12130 2 12146
rect -98 12096 -82 12130
rect -14 12096 2 12130
rect -98 12058 2 12096
rect 60 12130 160 12146
rect 60 12096 76 12130
rect 144 12096 160 12130
rect 60 12058 160 12096
rect 218 12130 318 12146
rect 218 12096 234 12130
rect 302 12096 318 12130
rect 218 12058 318 12096
rect 376 12130 476 12146
rect 376 12096 392 12130
rect 460 12096 476 12130
rect 376 12058 476 12096
rect 534 12130 634 12146
rect 534 12096 550 12130
rect 618 12096 634 12130
rect 534 12058 634 12096
rect 692 12130 792 12146
rect 692 12096 708 12130
rect 776 12096 792 12130
rect 692 12058 792 12096
rect 850 12130 950 12146
rect 850 12096 866 12130
rect 934 12096 950 12130
rect 850 12058 950 12096
rect 1008 12130 1108 12146
rect 1008 12096 1024 12130
rect 1092 12096 1108 12130
rect 1008 12058 1108 12096
rect 1166 12130 1266 12146
rect 1166 12096 1182 12130
rect 1250 12096 1266 12130
rect 1166 12058 1266 12096
rect 1324 12130 1424 12146
rect 1324 12096 1340 12130
rect 1408 12096 1424 12130
rect 1324 12058 1424 12096
rect 1482 12130 1582 12146
rect 1482 12096 1498 12130
rect 1566 12096 1582 12130
rect 1482 12058 1582 12096
rect 1640 12130 1740 12146
rect 1640 12096 1656 12130
rect 1724 12096 1740 12130
rect 1640 12058 1740 12096
rect 1798 12130 1898 12146
rect 1798 12096 1814 12130
rect 1882 12096 1898 12130
rect 1798 12058 1898 12096
rect 1956 12130 2056 12146
rect 1956 12096 1972 12130
rect 2040 12096 2056 12130
rect 1956 12058 2056 12096
rect 2114 12130 2214 12146
rect 2114 12096 2130 12130
rect 2198 12096 2214 12130
rect 2114 12058 2214 12096
rect 2272 12130 2372 12146
rect 2272 12096 2288 12130
rect 2356 12096 2372 12130
rect 2272 12058 2372 12096
rect 2430 12130 2530 12146
rect 2430 12096 2446 12130
rect 2514 12096 2530 12130
rect 2430 12058 2530 12096
rect 2588 12130 2688 12146
rect 2588 12096 2604 12130
rect 2672 12096 2688 12130
rect 2588 12058 2688 12096
rect 2746 12130 2846 12146
rect 2746 12096 2762 12130
rect 2830 12096 2846 12130
rect 2746 12058 2846 12096
rect 2904 12130 3004 12146
rect 2904 12096 2920 12130
rect 2988 12096 3004 12130
rect 2904 12058 3004 12096
rect 3062 12130 3162 12146
rect 3062 12096 3078 12130
rect 3146 12096 3162 12130
rect 3062 12058 3162 12096
rect 3220 12130 3320 12146
rect 3220 12096 3236 12130
rect 3304 12096 3320 12130
rect 3220 12058 3320 12096
rect 3378 12130 3478 12146
rect 3378 12096 3394 12130
rect 3462 12096 3478 12130
rect 3378 12058 3478 12096
rect 3536 12130 3636 12146
rect 3536 12096 3552 12130
rect 3620 12096 3636 12130
rect 3536 12058 3636 12096
rect 3694 12130 3794 12146
rect 3694 12096 3710 12130
rect 3778 12096 3794 12130
rect 3694 12058 3794 12096
rect 3852 12130 3952 12146
rect 3852 12096 3868 12130
rect 3936 12096 3952 12130
rect 3852 12058 3952 12096
rect 4010 12130 4110 12146
rect 4010 12096 4026 12130
rect 4094 12096 4110 12130
rect 4010 12058 4110 12096
rect -572 6020 -472 6058
rect -572 5986 -556 6020
rect -488 5986 -472 6020
rect -572 5970 -472 5986
rect -414 6020 -314 6058
rect -414 5986 -398 6020
rect -330 5986 -314 6020
rect -414 5970 -314 5986
rect -256 6020 -156 6058
rect -256 5986 -240 6020
rect -172 5986 -156 6020
rect -256 5970 -156 5986
rect -98 6020 2 6058
rect -98 5986 -82 6020
rect -14 5986 2 6020
rect -98 5970 2 5986
rect 60 6020 160 6058
rect 60 5986 76 6020
rect 144 5986 160 6020
rect 60 5970 160 5986
rect 218 6020 318 6058
rect 218 5986 234 6020
rect 302 5986 318 6020
rect 218 5970 318 5986
rect 376 6020 476 6058
rect 376 5986 392 6020
rect 460 5986 476 6020
rect 376 5970 476 5986
rect 534 6020 634 6058
rect 534 5986 550 6020
rect 618 5986 634 6020
rect 534 5970 634 5986
rect 692 6020 792 6058
rect 692 5986 708 6020
rect 776 5986 792 6020
rect 692 5970 792 5986
rect 850 6020 950 6058
rect 850 5986 866 6020
rect 934 5986 950 6020
rect 850 5970 950 5986
rect 1008 6020 1108 6058
rect 1008 5986 1024 6020
rect 1092 5986 1108 6020
rect 1008 5970 1108 5986
rect 1166 6020 1266 6058
rect 1166 5986 1182 6020
rect 1250 5986 1266 6020
rect 1166 5970 1266 5986
rect 1324 6020 1424 6058
rect 1324 5986 1340 6020
rect 1408 5986 1424 6020
rect 1324 5970 1424 5986
rect 1482 6020 1582 6058
rect 1482 5986 1498 6020
rect 1566 5986 1582 6020
rect 1482 5970 1582 5986
rect 1640 6020 1740 6058
rect 1640 5986 1656 6020
rect 1724 5986 1740 6020
rect 1640 5970 1740 5986
rect 1798 6020 1898 6058
rect 1798 5986 1814 6020
rect 1882 5986 1898 6020
rect 1798 5970 1898 5986
rect 1956 6020 2056 6058
rect 1956 5986 1972 6020
rect 2040 5986 2056 6020
rect 1956 5970 2056 5986
rect 2114 6020 2214 6058
rect 2114 5986 2130 6020
rect 2198 5986 2214 6020
rect 2114 5970 2214 5986
rect 2272 6020 2372 6058
rect 2272 5986 2288 6020
rect 2356 5986 2372 6020
rect 2272 5970 2372 5986
rect 2430 6020 2530 6058
rect 2430 5986 2446 6020
rect 2514 5986 2530 6020
rect 2430 5970 2530 5986
rect 2588 6020 2688 6058
rect 2588 5986 2604 6020
rect 2672 5986 2688 6020
rect 2588 5970 2688 5986
rect 2746 6020 2846 6058
rect 2746 5986 2762 6020
rect 2830 5986 2846 6020
rect 2746 5970 2846 5986
rect 2904 6020 3004 6058
rect 2904 5986 2920 6020
rect 2988 5986 3004 6020
rect 2904 5970 3004 5986
rect 3062 6020 3162 6058
rect 3062 5986 3078 6020
rect 3146 5986 3162 6020
rect 3062 5970 3162 5986
rect 3220 6020 3320 6058
rect 3220 5986 3236 6020
rect 3304 5986 3320 6020
rect 3220 5970 3320 5986
rect 3378 6020 3478 6058
rect 3378 5986 3394 6020
rect 3462 5986 3478 6020
rect 3378 5970 3478 5986
rect 3536 6020 3636 6058
rect 3536 5986 3552 6020
rect 3620 5986 3636 6020
rect 3536 5970 3636 5986
rect 3694 6020 3794 6058
rect 3694 5986 3710 6020
rect 3778 5986 3794 6020
rect 3694 5970 3794 5986
rect 3852 6020 3952 6058
rect 3852 5986 3868 6020
rect 3936 5986 3952 6020
rect 3852 5970 3952 5986
rect 4010 6020 4110 6058
rect 4010 5986 4026 6020
rect 4094 5986 4110 6020
rect 4010 5970 4110 5986
rect 5728 12130 5828 12146
rect 5728 12096 5744 12130
rect 5812 12096 5828 12130
rect 5728 12058 5828 12096
rect 5886 12130 5986 12146
rect 5886 12096 5902 12130
rect 5970 12096 5986 12130
rect 5886 12058 5986 12096
rect 6044 12130 6144 12146
rect 6044 12096 6060 12130
rect 6128 12096 6144 12130
rect 6044 12058 6144 12096
rect 6202 12130 6302 12146
rect 6202 12096 6218 12130
rect 6286 12096 6302 12130
rect 6202 12058 6302 12096
rect 6360 12130 6460 12146
rect 6360 12096 6376 12130
rect 6444 12096 6460 12130
rect 6360 12058 6460 12096
rect 6518 12130 6618 12146
rect 6518 12096 6534 12130
rect 6602 12096 6618 12130
rect 6518 12058 6618 12096
rect 6676 12130 6776 12146
rect 6676 12096 6692 12130
rect 6760 12096 6776 12130
rect 6676 12058 6776 12096
rect 6834 12130 6934 12146
rect 6834 12096 6850 12130
rect 6918 12096 6934 12130
rect 6834 12058 6934 12096
rect 6992 12130 7092 12146
rect 6992 12096 7008 12130
rect 7076 12096 7092 12130
rect 6992 12058 7092 12096
rect 7150 12130 7250 12146
rect 7150 12096 7166 12130
rect 7234 12096 7250 12130
rect 7150 12058 7250 12096
rect 7308 12130 7408 12146
rect 7308 12096 7324 12130
rect 7392 12096 7408 12130
rect 7308 12058 7408 12096
rect 7466 12130 7566 12146
rect 7466 12096 7482 12130
rect 7550 12096 7566 12130
rect 7466 12058 7566 12096
rect 7624 12130 7724 12146
rect 7624 12096 7640 12130
rect 7708 12096 7724 12130
rect 7624 12058 7724 12096
rect 7782 12130 7882 12146
rect 7782 12096 7798 12130
rect 7866 12096 7882 12130
rect 7782 12058 7882 12096
rect 7940 12130 8040 12146
rect 7940 12096 7956 12130
rect 8024 12096 8040 12130
rect 7940 12058 8040 12096
rect 8098 12130 8198 12146
rect 8098 12096 8114 12130
rect 8182 12096 8198 12130
rect 8098 12058 8198 12096
rect 8256 12130 8356 12146
rect 8256 12096 8272 12130
rect 8340 12096 8356 12130
rect 8256 12058 8356 12096
rect 8414 12130 8514 12146
rect 8414 12096 8430 12130
rect 8498 12096 8514 12130
rect 8414 12058 8514 12096
rect 8572 12130 8672 12146
rect 8572 12096 8588 12130
rect 8656 12096 8672 12130
rect 8572 12058 8672 12096
rect 8730 12130 8830 12146
rect 8730 12096 8746 12130
rect 8814 12096 8830 12130
rect 8730 12058 8830 12096
rect 8888 12130 8988 12146
rect 8888 12096 8904 12130
rect 8972 12096 8988 12130
rect 8888 12058 8988 12096
rect 9046 12130 9146 12146
rect 9046 12096 9062 12130
rect 9130 12096 9146 12130
rect 9046 12058 9146 12096
rect 9204 12130 9304 12146
rect 9204 12096 9220 12130
rect 9288 12096 9304 12130
rect 9204 12058 9304 12096
rect 9362 12130 9462 12146
rect 9362 12096 9378 12130
rect 9446 12096 9462 12130
rect 9362 12058 9462 12096
rect 9520 12130 9620 12146
rect 9520 12096 9536 12130
rect 9604 12096 9620 12130
rect 9520 12058 9620 12096
rect 9678 12130 9778 12146
rect 9678 12096 9694 12130
rect 9762 12096 9778 12130
rect 9678 12058 9778 12096
rect 9836 12130 9936 12146
rect 9836 12096 9852 12130
rect 9920 12096 9936 12130
rect 9836 12058 9936 12096
rect 9994 12130 10094 12146
rect 9994 12096 10010 12130
rect 10078 12096 10094 12130
rect 9994 12058 10094 12096
rect 10152 12130 10252 12146
rect 10152 12096 10168 12130
rect 10236 12096 10252 12130
rect 10152 12058 10252 12096
rect 10310 12130 10410 12146
rect 10310 12096 10326 12130
rect 10394 12096 10410 12130
rect 10310 12058 10410 12096
rect 5728 6020 5828 6058
rect 5728 5986 5744 6020
rect 5812 5986 5828 6020
rect 5728 5970 5828 5986
rect 5886 6020 5986 6058
rect 5886 5986 5902 6020
rect 5970 5986 5986 6020
rect 5886 5970 5986 5986
rect 6044 6020 6144 6058
rect 6044 5986 6060 6020
rect 6128 5986 6144 6020
rect 6044 5970 6144 5986
rect 6202 6020 6302 6058
rect 6202 5986 6218 6020
rect 6286 5986 6302 6020
rect 6202 5970 6302 5986
rect 6360 6020 6460 6058
rect 6360 5986 6376 6020
rect 6444 5986 6460 6020
rect 6360 5970 6460 5986
rect 6518 6020 6618 6058
rect 6518 5986 6534 6020
rect 6602 5986 6618 6020
rect 6518 5970 6618 5986
rect 6676 6020 6776 6058
rect 6676 5986 6692 6020
rect 6760 5986 6776 6020
rect 6676 5970 6776 5986
rect 6834 6020 6934 6058
rect 6834 5986 6850 6020
rect 6918 5986 6934 6020
rect 6834 5970 6934 5986
rect 6992 6020 7092 6058
rect 6992 5986 7008 6020
rect 7076 5986 7092 6020
rect 6992 5970 7092 5986
rect 7150 6020 7250 6058
rect 7150 5986 7166 6020
rect 7234 5986 7250 6020
rect 7150 5970 7250 5986
rect 7308 6020 7408 6058
rect 7308 5986 7324 6020
rect 7392 5986 7408 6020
rect 7308 5970 7408 5986
rect 7466 6020 7566 6058
rect 7466 5986 7482 6020
rect 7550 5986 7566 6020
rect 7466 5970 7566 5986
rect 7624 6020 7724 6058
rect 7624 5986 7640 6020
rect 7708 5986 7724 6020
rect 7624 5970 7724 5986
rect 7782 6020 7882 6058
rect 7782 5986 7798 6020
rect 7866 5986 7882 6020
rect 7782 5970 7882 5986
rect 7940 6020 8040 6058
rect 7940 5986 7956 6020
rect 8024 5986 8040 6020
rect 7940 5970 8040 5986
rect 8098 6020 8198 6058
rect 8098 5986 8114 6020
rect 8182 5986 8198 6020
rect 8098 5970 8198 5986
rect 8256 6020 8356 6058
rect 8256 5986 8272 6020
rect 8340 5986 8356 6020
rect 8256 5970 8356 5986
rect 8414 6020 8514 6058
rect 8414 5986 8430 6020
rect 8498 5986 8514 6020
rect 8414 5970 8514 5986
rect 8572 6020 8672 6058
rect 8572 5986 8588 6020
rect 8656 5986 8672 6020
rect 8572 5970 8672 5986
rect 8730 6020 8830 6058
rect 8730 5986 8746 6020
rect 8814 5986 8830 6020
rect 8730 5970 8830 5986
rect 8888 6020 8988 6058
rect 8888 5986 8904 6020
rect 8972 5986 8988 6020
rect 8888 5970 8988 5986
rect 9046 6020 9146 6058
rect 9046 5986 9062 6020
rect 9130 5986 9146 6020
rect 9046 5970 9146 5986
rect 9204 6020 9304 6058
rect 9204 5986 9220 6020
rect 9288 5986 9304 6020
rect 9204 5970 9304 5986
rect 9362 6020 9462 6058
rect 9362 5986 9378 6020
rect 9446 5986 9462 6020
rect 9362 5970 9462 5986
rect 9520 6020 9620 6058
rect 9520 5986 9536 6020
rect 9604 5986 9620 6020
rect 9520 5970 9620 5986
rect 9678 6020 9778 6058
rect 9678 5986 9694 6020
rect 9762 5986 9778 6020
rect 9678 5970 9778 5986
rect 9836 6020 9936 6058
rect 9836 5986 9852 6020
rect 9920 5986 9936 6020
rect 9836 5970 9936 5986
rect 9994 6020 10094 6058
rect 9994 5986 10010 6020
rect 10078 5986 10094 6020
rect 9994 5970 10094 5986
rect 10152 6020 10252 6058
rect 10152 5986 10168 6020
rect 10236 5986 10252 6020
rect 10152 5970 10252 5986
rect 10310 6020 10410 6058
rect 10310 5986 10326 6020
rect 10394 5986 10410 6020
rect 10310 5970 10410 5986
<< polycont >>
rect -13156 49696 -13088 49730
rect -12998 49696 -12930 49730
rect -12840 49696 -12772 49730
rect -12682 49696 -12614 49730
rect -12524 49696 -12456 49730
rect -12366 49696 -12298 49730
rect -12208 49696 -12140 49730
rect -12050 49696 -11982 49730
rect -11892 49696 -11824 49730
rect -11734 49696 -11666 49730
rect -11576 49696 -11508 49730
rect -11418 49696 -11350 49730
rect -11260 49696 -11192 49730
rect -11102 49696 -11034 49730
rect -10944 49696 -10876 49730
rect -10786 49696 -10718 49730
rect -10628 49696 -10560 49730
rect -10470 49696 -10402 49730
rect -10312 49696 -10244 49730
rect -10154 49696 -10086 49730
rect -9996 49696 -9928 49730
rect -9838 49696 -9770 49730
rect -9680 49696 -9612 49730
rect -9522 49696 -9454 49730
rect -9364 49696 -9296 49730
rect -9206 49696 -9138 49730
rect -9048 49696 -8980 49730
rect -8890 49696 -8822 49730
rect -8732 49696 -8664 49730
rect -8574 49696 -8506 49730
rect -13156 43586 -13088 43620
rect -12998 43586 -12930 43620
rect -12840 43586 -12772 43620
rect -12682 43586 -12614 43620
rect -12524 43586 -12456 43620
rect -12366 43586 -12298 43620
rect -12208 43586 -12140 43620
rect -12050 43586 -11982 43620
rect -11892 43586 -11824 43620
rect -11734 43586 -11666 43620
rect -11576 43586 -11508 43620
rect -11418 43586 -11350 43620
rect -11260 43586 -11192 43620
rect -11102 43586 -11034 43620
rect -10944 43586 -10876 43620
rect -10786 43586 -10718 43620
rect -10628 43586 -10560 43620
rect -10470 43586 -10402 43620
rect -10312 43586 -10244 43620
rect -10154 43586 -10086 43620
rect -9996 43586 -9928 43620
rect -9838 43586 -9770 43620
rect -9680 43586 -9612 43620
rect -9522 43586 -9454 43620
rect -9364 43586 -9296 43620
rect -9206 43586 -9138 43620
rect -9048 43586 -8980 43620
rect -8890 43586 -8822 43620
rect -8732 43586 -8664 43620
rect -8574 43586 -8506 43620
rect -6856 49696 -6788 49730
rect -6698 49696 -6630 49730
rect -6540 49696 -6472 49730
rect -6382 49696 -6314 49730
rect -6224 49696 -6156 49730
rect -6066 49696 -5998 49730
rect -5908 49696 -5840 49730
rect -5750 49696 -5682 49730
rect -5592 49696 -5524 49730
rect -5434 49696 -5366 49730
rect -5276 49696 -5208 49730
rect -5118 49696 -5050 49730
rect -4960 49696 -4892 49730
rect -4802 49696 -4734 49730
rect -4644 49696 -4576 49730
rect -4486 49696 -4418 49730
rect -4328 49696 -4260 49730
rect -4170 49696 -4102 49730
rect -4012 49696 -3944 49730
rect -3854 49696 -3786 49730
rect -3696 49696 -3628 49730
rect -3538 49696 -3470 49730
rect -3380 49696 -3312 49730
rect -3222 49696 -3154 49730
rect -3064 49696 -2996 49730
rect -2906 49696 -2838 49730
rect -2748 49696 -2680 49730
rect -2590 49696 -2522 49730
rect -2432 49696 -2364 49730
rect -2274 49696 -2206 49730
rect -6856 43586 -6788 43620
rect -6698 43586 -6630 43620
rect -6540 43586 -6472 43620
rect -6382 43586 -6314 43620
rect -6224 43586 -6156 43620
rect -6066 43586 -5998 43620
rect -5908 43586 -5840 43620
rect -5750 43586 -5682 43620
rect -5592 43586 -5524 43620
rect -5434 43586 -5366 43620
rect -5276 43586 -5208 43620
rect -5118 43586 -5050 43620
rect -4960 43586 -4892 43620
rect -4802 43586 -4734 43620
rect -4644 43586 -4576 43620
rect -4486 43586 -4418 43620
rect -4328 43586 -4260 43620
rect -4170 43586 -4102 43620
rect -4012 43586 -3944 43620
rect -3854 43586 -3786 43620
rect -3696 43586 -3628 43620
rect -3538 43586 -3470 43620
rect -3380 43586 -3312 43620
rect -3222 43586 -3154 43620
rect -3064 43586 -2996 43620
rect -2906 43586 -2838 43620
rect -2748 43586 -2680 43620
rect -2590 43586 -2522 43620
rect -2432 43586 -2364 43620
rect -2274 43586 -2206 43620
rect -556 49696 -488 49730
rect -398 49696 -330 49730
rect -240 49696 -172 49730
rect -82 49696 -14 49730
rect 76 49696 144 49730
rect 234 49696 302 49730
rect 392 49696 460 49730
rect 550 49696 618 49730
rect 708 49696 776 49730
rect 866 49696 934 49730
rect 1024 49696 1092 49730
rect 1182 49696 1250 49730
rect 1340 49696 1408 49730
rect 1498 49696 1566 49730
rect 1656 49696 1724 49730
rect 1814 49696 1882 49730
rect 1972 49696 2040 49730
rect 2130 49696 2198 49730
rect 2288 49696 2356 49730
rect 2446 49696 2514 49730
rect 2604 49696 2672 49730
rect 2762 49696 2830 49730
rect 2920 49696 2988 49730
rect 3078 49696 3146 49730
rect 3236 49696 3304 49730
rect 3394 49696 3462 49730
rect 3552 49696 3620 49730
rect 3710 49696 3778 49730
rect 3868 49696 3936 49730
rect 4026 49696 4094 49730
rect -556 43586 -488 43620
rect -398 43586 -330 43620
rect -240 43586 -172 43620
rect -82 43586 -14 43620
rect 76 43586 144 43620
rect 234 43586 302 43620
rect 392 43586 460 43620
rect 550 43586 618 43620
rect 708 43586 776 43620
rect 866 43586 934 43620
rect 1024 43586 1092 43620
rect 1182 43586 1250 43620
rect 1340 43586 1408 43620
rect 1498 43586 1566 43620
rect 1656 43586 1724 43620
rect 1814 43586 1882 43620
rect 1972 43586 2040 43620
rect 2130 43586 2198 43620
rect 2288 43586 2356 43620
rect 2446 43586 2514 43620
rect 2604 43586 2672 43620
rect 2762 43586 2830 43620
rect 2920 43586 2988 43620
rect 3078 43586 3146 43620
rect 3236 43586 3304 43620
rect 3394 43586 3462 43620
rect 3552 43586 3620 43620
rect 3710 43586 3778 43620
rect 3868 43586 3936 43620
rect 4026 43586 4094 43620
rect 5744 49696 5812 49730
rect 5902 49696 5970 49730
rect 6060 49696 6128 49730
rect 6218 49696 6286 49730
rect 6376 49696 6444 49730
rect 6534 49696 6602 49730
rect 6692 49696 6760 49730
rect 6850 49696 6918 49730
rect 7008 49696 7076 49730
rect 7166 49696 7234 49730
rect 7324 49696 7392 49730
rect 7482 49696 7550 49730
rect 7640 49696 7708 49730
rect 7798 49696 7866 49730
rect 7956 49696 8024 49730
rect 8114 49696 8182 49730
rect 8272 49696 8340 49730
rect 8430 49696 8498 49730
rect 8588 49696 8656 49730
rect 8746 49696 8814 49730
rect 8904 49696 8972 49730
rect 9062 49696 9130 49730
rect 9220 49696 9288 49730
rect 9378 49696 9446 49730
rect 9536 49696 9604 49730
rect 9694 49696 9762 49730
rect 9852 49696 9920 49730
rect 10010 49696 10078 49730
rect 10168 49696 10236 49730
rect 10326 49696 10394 49730
rect 5744 43586 5812 43620
rect 5902 43586 5970 43620
rect 6060 43586 6128 43620
rect 6218 43586 6286 43620
rect 6376 43586 6444 43620
rect 6534 43586 6602 43620
rect 6692 43586 6760 43620
rect 6850 43586 6918 43620
rect 7008 43586 7076 43620
rect 7166 43586 7234 43620
rect 7324 43586 7392 43620
rect 7482 43586 7550 43620
rect 7640 43586 7708 43620
rect 7798 43586 7866 43620
rect 7956 43586 8024 43620
rect 8114 43586 8182 43620
rect 8272 43586 8340 43620
rect 8430 43586 8498 43620
rect 8588 43586 8656 43620
rect 8746 43586 8814 43620
rect 8904 43586 8972 43620
rect 9062 43586 9130 43620
rect 9220 43586 9288 43620
rect 9378 43586 9446 43620
rect 9536 43586 9604 43620
rect 9694 43586 9762 43620
rect 9852 43586 9920 43620
rect 10010 43586 10078 43620
rect 10168 43586 10236 43620
rect 10326 43586 10394 43620
rect -13156 42696 -13088 42730
rect -12998 42696 -12930 42730
rect -12840 42696 -12772 42730
rect -12682 42696 -12614 42730
rect -12524 42696 -12456 42730
rect -12366 42696 -12298 42730
rect -12208 42696 -12140 42730
rect -12050 42696 -11982 42730
rect -11892 42696 -11824 42730
rect -11734 42696 -11666 42730
rect -11576 42696 -11508 42730
rect -11418 42696 -11350 42730
rect -11260 42696 -11192 42730
rect -11102 42696 -11034 42730
rect -10944 42696 -10876 42730
rect -10786 42696 -10718 42730
rect -10628 42696 -10560 42730
rect -10470 42696 -10402 42730
rect -10312 42696 -10244 42730
rect -10154 42696 -10086 42730
rect -9996 42696 -9928 42730
rect -9838 42696 -9770 42730
rect -9680 42696 -9612 42730
rect -9522 42696 -9454 42730
rect -9364 42696 -9296 42730
rect -9206 42696 -9138 42730
rect -9048 42696 -8980 42730
rect -8890 42696 -8822 42730
rect -8732 42696 -8664 42730
rect -8574 42696 -8506 42730
rect -13156 36586 -13088 36620
rect -12998 36586 -12930 36620
rect -12840 36586 -12772 36620
rect -12682 36586 -12614 36620
rect -12524 36586 -12456 36620
rect -12366 36586 -12298 36620
rect -12208 36586 -12140 36620
rect -12050 36586 -11982 36620
rect -11892 36586 -11824 36620
rect -11734 36586 -11666 36620
rect -11576 36586 -11508 36620
rect -11418 36586 -11350 36620
rect -11260 36586 -11192 36620
rect -11102 36586 -11034 36620
rect -10944 36586 -10876 36620
rect -10786 36586 -10718 36620
rect -10628 36586 -10560 36620
rect -10470 36586 -10402 36620
rect -10312 36586 -10244 36620
rect -10154 36586 -10086 36620
rect -9996 36586 -9928 36620
rect -9838 36586 -9770 36620
rect -9680 36586 -9612 36620
rect -9522 36586 -9454 36620
rect -9364 36586 -9296 36620
rect -9206 36586 -9138 36620
rect -9048 36586 -8980 36620
rect -8890 36586 -8822 36620
rect -8732 36586 -8664 36620
rect -8574 36586 -8506 36620
rect -6856 42696 -6788 42730
rect -6698 42696 -6630 42730
rect -6540 42696 -6472 42730
rect -6382 42696 -6314 42730
rect -6224 42696 -6156 42730
rect -6066 42696 -5998 42730
rect -5908 42696 -5840 42730
rect -5750 42696 -5682 42730
rect -5592 42696 -5524 42730
rect -5434 42696 -5366 42730
rect -5276 42696 -5208 42730
rect -5118 42696 -5050 42730
rect -4960 42696 -4892 42730
rect -4802 42696 -4734 42730
rect -4644 42696 -4576 42730
rect -4486 42696 -4418 42730
rect -4328 42696 -4260 42730
rect -4170 42696 -4102 42730
rect -4012 42696 -3944 42730
rect -3854 42696 -3786 42730
rect -3696 42696 -3628 42730
rect -3538 42696 -3470 42730
rect -3380 42696 -3312 42730
rect -3222 42696 -3154 42730
rect -3064 42696 -2996 42730
rect -2906 42696 -2838 42730
rect -2748 42696 -2680 42730
rect -2590 42696 -2522 42730
rect -2432 42696 -2364 42730
rect -2274 42696 -2206 42730
rect -6856 36586 -6788 36620
rect -6698 36586 -6630 36620
rect -6540 36586 -6472 36620
rect -6382 36586 -6314 36620
rect -6224 36586 -6156 36620
rect -6066 36586 -5998 36620
rect -5908 36586 -5840 36620
rect -5750 36586 -5682 36620
rect -5592 36586 -5524 36620
rect -5434 36586 -5366 36620
rect -5276 36586 -5208 36620
rect -5118 36586 -5050 36620
rect -4960 36586 -4892 36620
rect -4802 36586 -4734 36620
rect -4644 36586 -4576 36620
rect -4486 36586 -4418 36620
rect -4328 36586 -4260 36620
rect -4170 36586 -4102 36620
rect -4012 36586 -3944 36620
rect -3854 36586 -3786 36620
rect -3696 36586 -3628 36620
rect -3538 36586 -3470 36620
rect -3380 36586 -3312 36620
rect -3222 36586 -3154 36620
rect -3064 36586 -2996 36620
rect -2906 36586 -2838 36620
rect -2748 36586 -2680 36620
rect -2590 36586 -2522 36620
rect -2432 36586 -2364 36620
rect -2274 36586 -2206 36620
rect -556 42696 -488 42730
rect -398 42696 -330 42730
rect -240 42696 -172 42730
rect -82 42696 -14 42730
rect 76 42696 144 42730
rect 234 42696 302 42730
rect 392 42696 460 42730
rect 550 42696 618 42730
rect 708 42696 776 42730
rect 866 42696 934 42730
rect 1024 42696 1092 42730
rect 1182 42696 1250 42730
rect 1340 42696 1408 42730
rect 1498 42696 1566 42730
rect 1656 42696 1724 42730
rect 1814 42696 1882 42730
rect 1972 42696 2040 42730
rect 2130 42696 2198 42730
rect 2288 42696 2356 42730
rect 2446 42696 2514 42730
rect 2604 42696 2672 42730
rect 2762 42696 2830 42730
rect 2920 42696 2988 42730
rect 3078 42696 3146 42730
rect 3236 42696 3304 42730
rect 3394 42696 3462 42730
rect 3552 42696 3620 42730
rect 3710 42696 3778 42730
rect 3868 42696 3936 42730
rect 4026 42696 4094 42730
rect -556 36586 -488 36620
rect -398 36586 -330 36620
rect -240 36586 -172 36620
rect -82 36586 -14 36620
rect 76 36586 144 36620
rect 234 36586 302 36620
rect 392 36586 460 36620
rect 550 36586 618 36620
rect 708 36586 776 36620
rect 866 36586 934 36620
rect 1024 36586 1092 36620
rect 1182 36586 1250 36620
rect 1340 36586 1408 36620
rect 1498 36586 1566 36620
rect 1656 36586 1724 36620
rect 1814 36586 1882 36620
rect 1972 36586 2040 36620
rect 2130 36586 2198 36620
rect 2288 36586 2356 36620
rect 2446 36586 2514 36620
rect 2604 36586 2672 36620
rect 2762 36586 2830 36620
rect 2920 36586 2988 36620
rect 3078 36586 3146 36620
rect 3236 36586 3304 36620
rect 3394 36586 3462 36620
rect 3552 36586 3620 36620
rect 3710 36586 3778 36620
rect 3868 36586 3936 36620
rect 4026 36586 4094 36620
rect 5744 42696 5812 42730
rect 5902 42696 5970 42730
rect 6060 42696 6128 42730
rect 6218 42696 6286 42730
rect 6376 42696 6444 42730
rect 6534 42696 6602 42730
rect 6692 42696 6760 42730
rect 6850 42696 6918 42730
rect 7008 42696 7076 42730
rect 7166 42696 7234 42730
rect 7324 42696 7392 42730
rect 7482 42696 7550 42730
rect 7640 42696 7708 42730
rect 7798 42696 7866 42730
rect 7956 42696 8024 42730
rect 8114 42696 8182 42730
rect 8272 42696 8340 42730
rect 8430 42696 8498 42730
rect 8588 42696 8656 42730
rect 8746 42696 8814 42730
rect 8904 42696 8972 42730
rect 9062 42696 9130 42730
rect 9220 42696 9288 42730
rect 9378 42696 9446 42730
rect 9536 42696 9604 42730
rect 9694 42696 9762 42730
rect 9852 42696 9920 42730
rect 10010 42696 10078 42730
rect 10168 42696 10236 42730
rect 10326 42696 10394 42730
rect 5744 36586 5812 36620
rect 5902 36586 5970 36620
rect 6060 36586 6128 36620
rect 6218 36586 6286 36620
rect 6376 36586 6444 36620
rect 6534 36586 6602 36620
rect 6692 36586 6760 36620
rect 6850 36586 6918 36620
rect 7008 36586 7076 36620
rect 7166 36586 7234 36620
rect 7324 36586 7392 36620
rect 7482 36586 7550 36620
rect 7640 36586 7708 36620
rect 7798 36586 7866 36620
rect 7956 36586 8024 36620
rect 8114 36586 8182 36620
rect 8272 36586 8340 36620
rect 8430 36586 8498 36620
rect 8588 36586 8656 36620
rect 8746 36586 8814 36620
rect 8904 36586 8972 36620
rect 9062 36586 9130 36620
rect 9220 36586 9288 36620
rect 9378 36586 9446 36620
rect 9536 36586 9604 36620
rect 9694 36586 9762 36620
rect 9852 36586 9920 36620
rect 10010 36586 10078 36620
rect 10168 36586 10236 36620
rect 10326 36586 10394 36620
rect -13156 34396 -13088 34430
rect -12998 34396 -12930 34430
rect -12840 34396 -12772 34430
rect -12682 34396 -12614 34430
rect -12524 34396 -12456 34430
rect -12366 34396 -12298 34430
rect -12208 34396 -12140 34430
rect -12050 34396 -11982 34430
rect -11892 34396 -11824 34430
rect -11734 34396 -11666 34430
rect -11576 34396 -11508 34430
rect -11418 34396 -11350 34430
rect -11260 34396 -11192 34430
rect -11102 34396 -11034 34430
rect -10944 34396 -10876 34430
rect -10786 34396 -10718 34430
rect -10628 34396 -10560 34430
rect -10470 34396 -10402 34430
rect -10312 34396 -10244 34430
rect -10154 34396 -10086 34430
rect -9996 34396 -9928 34430
rect -9838 34396 -9770 34430
rect -9680 34396 -9612 34430
rect -9522 34396 -9454 34430
rect -9364 34396 -9296 34430
rect -9206 34396 -9138 34430
rect -9048 34396 -8980 34430
rect -8890 34396 -8822 34430
rect -8732 34396 -8664 34430
rect -8574 34396 -8506 34430
rect -13156 28286 -13088 28320
rect -12998 28286 -12930 28320
rect -12840 28286 -12772 28320
rect -12682 28286 -12614 28320
rect -12524 28286 -12456 28320
rect -12366 28286 -12298 28320
rect -12208 28286 -12140 28320
rect -12050 28286 -11982 28320
rect -11892 28286 -11824 28320
rect -11734 28286 -11666 28320
rect -11576 28286 -11508 28320
rect -11418 28286 -11350 28320
rect -11260 28286 -11192 28320
rect -11102 28286 -11034 28320
rect -10944 28286 -10876 28320
rect -10786 28286 -10718 28320
rect -10628 28286 -10560 28320
rect -10470 28286 -10402 28320
rect -10312 28286 -10244 28320
rect -10154 28286 -10086 28320
rect -9996 28286 -9928 28320
rect -9838 28286 -9770 28320
rect -9680 28286 -9612 28320
rect -9522 28286 -9454 28320
rect -9364 28286 -9296 28320
rect -9206 28286 -9138 28320
rect -9048 28286 -8980 28320
rect -8890 28286 -8822 28320
rect -8732 28286 -8664 28320
rect -8574 28286 -8506 28320
rect -6856 34396 -6788 34430
rect -6698 34396 -6630 34430
rect -6540 34396 -6472 34430
rect -6382 34396 -6314 34430
rect -6224 34396 -6156 34430
rect -6066 34396 -5998 34430
rect -5908 34396 -5840 34430
rect -5750 34396 -5682 34430
rect -5592 34396 -5524 34430
rect -5434 34396 -5366 34430
rect -5276 34396 -5208 34430
rect -5118 34396 -5050 34430
rect -4960 34396 -4892 34430
rect -4802 34396 -4734 34430
rect -4644 34396 -4576 34430
rect -4486 34396 -4418 34430
rect -4328 34396 -4260 34430
rect -4170 34396 -4102 34430
rect -4012 34396 -3944 34430
rect -3854 34396 -3786 34430
rect -3696 34396 -3628 34430
rect -3538 34396 -3470 34430
rect -3380 34396 -3312 34430
rect -3222 34396 -3154 34430
rect -3064 34396 -2996 34430
rect -2906 34396 -2838 34430
rect -2748 34396 -2680 34430
rect -2590 34396 -2522 34430
rect -2432 34396 -2364 34430
rect -2274 34396 -2206 34430
rect -6856 28286 -6788 28320
rect -6698 28286 -6630 28320
rect -6540 28286 -6472 28320
rect -6382 28286 -6314 28320
rect -6224 28286 -6156 28320
rect -6066 28286 -5998 28320
rect -5908 28286 -5840 28320
rect -5750 28286 -5682 28320
rect -5592 28286 -5524 28320
rect -5434 28286 -5366 28320
rect -5276 28286 -5208 28320
rect -5118 28286 -5050 28320
rect -4960 28286 -4892 28320
rect -4802 28286 -4734 28320
rect -4644 28286 -4576 28320
rect -4486 28286 -4418 28320
rect -4328 28286 -4260 28320
rect -4170 28286 -4102 28320
rect -4012 28286 -3944 28320
rect -3854 28286 -3786 28320
rect -3696 28286 -3628 28320
rect -3538 28286 -3470 28320
rect -3380 28286 -3312 28320
rect -3222 28286 -3154 28320
rect -3064 28286 -2996 28320
rect -2906 28286 -2838 28320
rect -2748 28286 -2680 28320
rect -2590 28286 -2522 28320
rect -2432 28286 -2364 28320
rect -2274 28286 -2206 28320
rect -556 34396 -488 34430
rect -398 34396 -330 34430
rect -240 34396 -172 34430
rect -82 34396 -14 34430
rect 76 34396 144 34430
rect 234 34396 302 34430
rect 392 34396 460 34430
rect 550 34396 618 34430
rect 708 34396 776 34430
rect 866 34396 934 34430
rect 1024 34396 1092 34430
rect 1182 34396 1250 34430
rect 1340 34396 1408 34430
rect 1498 34396 1566 34430
rect 1656 34396 1724 34430
rect 1814 34396 1882 34430
rect 1972 34396 2040 34430
rect 2130 34396 2198 34430
rect 2288 34396 2356 34430
rect 2446 34396 2514 34430
rect 2604 34396 2672 34430
rect 2762 34396 2830 34430
rect 2920 34396 2988 34430
rect 3078 34396 3146 34430
rect 3236 34396 3304 34430
rect 3394 34396 3462 34430
rect 3552 34396 3620 34430
rect 3710 34396 3778 34430
rect 3868 34396 3936 34430
rect 4026 34396 4094 34430
rect -556 28286 -488 28320
rect -398 28286 -330 28320
rect -240 28286 -172 28320
rect -82 28286 -14 28320
rect 76 28286 144 28320
rect 234 28286 302 28320
rect 392 28286 460 28320
rect 550 28286 618 28320
rect 708 28286 776 28320
rect 866 28286 934 28320
rect 1024 28286 1092 28320
rect 1182 28286 1250 28320
rect 1340 28286 1408 28320
rect 1498 28286 1566 28320
rect 1656 28286 1724 28320
rect 1814 28286 1882 28320
rect 1972 28286 2040 28320
rect 2130 28286 2198 28320
rect 2288 28286 2356 28320
rect 2446 28286 2514 28320
rect 2604 28286 2672 28320
rect 2762 28286 2830 28320
rect 2920 28286 2988 28320
rect 3078 28286 3146 28320
rect 3236 28286 3304 28320
rect 3394 28286 3462 28320
rect 3552 28286 3620 28320
rect 3710 28286 3778 28320
rect 3868 28286 3936 28320
rect 4026 28286 4094 28320
rect 5744 34396 5812 34430
rect 5902 34396 5970 34430
rect 6060 34396 6128 34430
rect 6218 34396 6286 34430
rect 6376 34396 6444 34430
rect 6534 34396 6602 34430
rect 6692 34396 6760 34430
rect 6850 34396 6918 34430
rect 7008 34396 7076 34430
rect 7166 34396 7234 34430
rect 7324 34396 7392 34430
rect 7482 34396 7550 34430
rect 7640 34396 7708 34430
rect 7798 34396 7866 34430
rect 7956 34396 8024 34430
rect 8114 34396 8182 34430
rect 8272 34396 8340 34430
rect 8430 34396 8498 34430
rect 8588 34396 8656 34430
rect 8746 34396 8814 34430
rect 8904 34396 8972 34430
rect 9062 34396 9130 34430
rect 9220 34396 9288 34430
rect 9378 34396 9446 34430
rect 9536 34396 9604 34430
rect 9694 34396 9762 34430
rect 9852 34396 9920 34430
rect 10010 34396 10078 34430
rect 10168 34396 10236 34430
rect 10326 34396 10394 34430
rect 5744 28286 5812 28320
rect 5902 28286 5970 28320
rect 6060 28286 6128 28320
rect 6218 28286 6286 28320
rect 6376 28286 6444 28320
rect 6534 28286 6602 28320
rect 6692 28286 6760 28320
rect 6850 28286 6918 28320
rect 7008 28286 7076 28320
rect 7166 28286 7234 28320
rect 7324 28286 7392 28320
rect 7482 28286 7550 28320
rect 7640 28286 7708 28320
rect 7798 28286 7866 28320
rect 7956 28286 8024 28320
rect 8114 28286 8182 28320
rect 8272 28286 8340 28320
rect 8430 28286 8498 28320
rect 8588 28286 8656 28320
rect 8746 28286 8814 28320
rect 8904 28286 8972 28320
rect 9062 28286 9130 28320
rect 9220 28286 9288 28320
rect 9378 28286 9446 28320
rect 9536 28286 9604 28320
rect 9694 28286 9762 28320
rect 9852 28286 9920 28320
rect 10010 28286 10078 28320
rect 10168 28286 10236 28320
rect 10326 28286 10394 28320
rect -13156 27396 -13088 27430
rect -12998 27396 -12930 27430
rect -12840 27396 -12772 27430
rect -12682 27396 -12614 27430
rect -12524 27396 -12456 27430
rect -12366 27396 -12298 27430
rect -12208 27396 -12140 27430
rect -12050 27396 -11982 27430
rect -11892 27396 -11824 27430
rect -11734 27396 -11666 27430
rect -11576 27396 -11508 27430
rect -11418 27396 -11350 27430
rect -11260 27396 -11192 27430
rect -11102 27396 -11034 27430
rect -10944 27396 -10876 27430
rect -10786 27396 -10718 27430
rect -10628 27396 -10560 27430
rect -10470 27396 -10402 27430
rect -10312 27396 -10244 27430
rect -10154 27396 -10086 27430
rect -9996 27396 -9928 27430
rect -9838 27396 -9770 27430
rect -9680 27396 -9612 27430
rect -9522 27396 -9454 27430
rect -9364 27396 -9296 27430
rect -9206 27396 -9138 27430
rect -9048 27396 -8980 27430
rect -8890 27396 -8822 27430
rect -8732 27396 -8664 27430
rect -8574 27396 -8506 27430
rect -13156 21286 -13088 21320
rect -12998 21286 -12930 21320
rect -12840 21286 -12772 21320
rect -12682 21286 -12614 21320
rect -12524 21286 -12456 21320
rect -12366 21286 -12298 21320
rect -12208 21286 -12140 21320
rect -12050 21286 -11982 21320
rect -11892 21286 -11824 21320
rect -11734 21286 -11666 21320
rect -11576 21286 -11508 21320
rect -11418 21286 -11350 21320
rect -11260 21286 -11192 21320
rect -11102 21286 -11034 21320
rect -10944 21286 -10876 21320
rect -10786 21286 -10718 21320
rect -10628 21286 -10560 21320
rect -10470 21286 -10402 21320
rect -10312 21286 -10244 21320
rect -10154 21286 -10086 21320
rect -9996 21286 -9928 21320
rect -9838 21286 -9770 21320
rect -9680 21286 -9612 21320
rect -9522 21286 -9454 21320
rect -9364 21286 -9296 21320
rect -9206 21286 -9138 21320
rect -9048 21286 -8980 21320
rect -8890 21286 -8822 21320
rect -8732 21286 -8664 21320
rect -8574 21286 -8506 21320
rect -6856 27396 -6788 27430
rect -6698 27396 -6630 27430
rect -6540 27396 -6472 27430
rect -6382 27396 -6314 27430
rect -6224 27396 -6156 27430
rect -6066 27396 -5998 27430
rect -5908 27396 -5840 27430
rect -5750 27396 -5682 27430
rect -5592 27396 -5524 27430
rect -5434 27396 -5366 27430
rect -5276 27396 -5208 27430
rect -5118 27396 -5050 27430
rect -4960 27396 -4892 27430
rect -4802 27396 -4734 27430
rect -4644 27396 -4576 27430
rect -4486 27396 -4418 27430
rect -4328 27396 -4260 27430
rect -4170 27396 -4102 27430
rect -4012 27396 -3944 27430
rect -3854 27396 -3786 27430
rect -3696 27396 -3628 27430
rect -3538 27396 -3470 27430
rect -3380 27396 -3312 27430
rect -3222 27396 -3154 27430
rect -3064 27396 -2996 27430
rect -2906 27396 -2838 27430
rect -2748 27396 -2680 27430
rect -2590 27396 -2522 27430
rect -2432 27396 -2364 27430
rect -2274 27396 -2206 27430
rect -6856 21286 -6788 21320
rect -6698 21286 -6630 21320
rect -6540 21286 -6472 21320
rect -6382 21286 -6314 21320
rect -6224 21286 -6156 21320
rect -6066 21286 -5998 21320
rect -5908 21286 -5840 21320
rect -5750 21286 -5682 21320
rect -5592 21286 -5524 21320
rect -5434 21286 -5366 21320
rect -5276 21286 -5208 21320
rect -5118 21286 -5050 21320
rect -4960 21286 -4892 21320
rect -4802 21286 -4734 21320
rect -4644 21286 -4576 21320
rect -4486 21286 -4418 21320
rect -4328 21286 -4260 21320
rect -4170 21286 -4102 21320
rect -4012 21286 -3944 21320
rect -3854 21286 -3786 21320
rect -3696 21286 -3628 21320
rect -3538 21286 -3470 21320
rect -3380 21286 -3312 21320
rect -3222 21286 -3154 21320
rect -3064 21286 -2996 21320
rect -2906 21286 -2838 21320
rect -2748 21286 -2680 21320
rect -2590 21286 -2522 21320
rect -2432 21286 -2364 21320
rect -2274 21286 -2206 21320
rect -556 27396 -488 27430
rect -398 27396 -330 27430
rect -240 27396 -172 27430
rect -82 27396 -14 27430
rect 76 27396 144 27430
rect 234 27396 302 27430
rect 392 27396 460 27430
rect 550 27396 618 27430
rect 708 27396 776 27430
rect 866 27396 934 27430
rect 1024 27396 1092 27430
rect 1182 27396 1250 27430
rect 1340 27396 1408 27430
rect 1498 27396 1566 27430
rect 1656 27396 1724 27430
rect 1814 27396 1882 27430
rect 1972 27396 2040 27430
rect 2130 27396 2198 27430
rect 2288 27396 2356 27430
rect 2446 27396 2514 27430
rect 2604 27396 2672 27430
rect 2762 27396 2830 27430
rect 2920 27396 2988 27430
rect 3078 27396 3146 27430
rect 3236 27396 3304 27430
rect 3394 27396 3462 27430
rect 3552 27396 3620 27430
rect 3710 27396 3778 27430
rect 3868 27396 3936 27430
rect 4026 27396 4094 27430
rect -556 21286 -488 21320
rect -398 21286 -330 21320
rect -240 21286 -172 21320
rect -82 21286 -14 21320
rect 76 21286 144 21320
rect 234 21286 302 21320
rect 392 21286 460 21320
rect 550 21286 618 21320
rect 708 21286 776 21320
rect 866 21286 934 21320
rect 1024 21286 1092 21320
rect 1182 21286 1250 21320
rect 1340 21286 1408 21320
rect 1498 21286 1566 21320
rect 1656 21286 1724 21320
rect 1814 21286 1882 21320
rect 1972 21286 2040 21320
rect 2130 21286 2198 21320
rect 2288 21286 2356 21320
rect 2446 21286 2514 21320
rect 2604 21286 2672 21320
rect 2762 21286 2830 21320
rect 2920 21286 2988 21320
rect 3078 21286 3146 21320
rect 3236 21286 3304 21320
rect 3394 21286 3462 21320
rect 3552 21286 3620 21320
rect 3710 21286 3778 21320
rect 3868 21286 3936 21320
rect 4026 21286 4094 21320
rect 5744 27396 5812 27430
rect 5902 27396 5970 27430
rect 6060 27396 6128 27430
rect 6218 27396 6286 27430
rect 6376 27396 6444 27430
rect 6534 27396 6602 27430
rect 6692 27396 6760 27430
rect 6850 27396 6918 27430
rect 7008 27396 7076 27430
rect 7166 27396 7234 27430
rect 7324 27396 7392 27430
rect 7482 27396 7550 27430
rect 7640 27396 7708 27430
rect 7798 27396 7866 27430
rect 7956 27396 8024 27430
rect 8114 27396 8182 27430
rect 8272 27396 8340 27430
rect 8430 27396 8498 27430
rect 8588 27396 8656 27430
rect 8746 27396 8814 27430
rect 8904 27396 8972 27430
rect 9062 27396 9130 27430
rect 9220 27396 9288 27430
rect 9378 27396 9446 27430
rect 9536 27396 9604 27430
rect 9694 27396 9762 27430
rect 9852 27396 9920 27430
rect 10010 27396 10078 27430
rect 10168 27396 10236 27430
rect 10326 27396 10394 27430
rect 5744 21286 5812 21320
rect 5902 21286 5970 21320
rect 6060 21286 6128 21320
rect 6218 21286 6286 21320
rect 6376 21286 6444 21320
rect 6534 21286 6602 21320
rect 6692 21286 6760 21320
rect 6850 21286 6918 21320
rect 7008 21286 7076 21320
rect 7166 21286 7234 21320
rect 7324 21286 7392 21320
rect 7482 21286 7550 21320
rect 7640 21286 7708 21320
rect 7798 21286 7866 21320
rect 7956 21286 8024 21320
rect 8114 21286 8182 21320
rect 8272 21286 8340 21320
rect 8430 21286 8498 21320
rect 8588 21286 8656 21320
rect 8746 21286 8814 21320
rect 8904 21286 8972 21320
rect 9062 21286 9130 21320
rect 9220 21286 9288 21320
rect 9378 21286 9446 21320
rect 9536 21286 9604 21320
rect 9694 21286 9762 21320
rect 9852 21286 9920 21320
rect 10010 21286 10078 21320
rect 10168 21286 10236 21320
rect 10326 21286 10394 21320
rect -13156 19096 -13088 19130
rect -12998 19096 -12930 19130
rect -12840 19096 -12772 19130
rect -12682 19096 -12614 19130
rect -12524 19096 -12456 19130
rect -12366 19096 -12298 19130
rect -12208 19096 -12140 19130
rect -12050 19096 -11982 19130
rect -11892 19096 -11824 19130
rect -11734 19096 -11666 19130
rect -11576 19096 -11508 19130
rect -11418 19096 -11350 19130
rect -11260 19096 -11192 19130
rect -11102 19096 -11034 19130
rect -10944 19096 -10876 19130
rect -10786 19096 -10718 19130
rect -10628 19096 -10560 19130
rect -10470 19096 -10402 19130
rect -10312 19096 -10244 19130
rect -10154 19096 -10086 19130
rect -9996 19096 -9928 19130
rect -9838 19096 -9770 19130
rect -9680 19096 -9612 19130
rect -9522 19096 -9454 19130
rect -9364 19096 -9296 19130
rect -9206 19096 -9138 19130
rect -9048 19096 -8980 19130
rect -8890 19096 -8822 19130
rect -8732 19096 -8664 19130
rect -8574 19096 -8506 19130
rect -13156 12986 -13088 13020
rect -12998 12986 -12930 13020
rect -12840 12986 -12772 13020
rect -12682 12986 -12614 13020
rect -12524 12986 -12456 13020
rect -12366 12986 -12298 13020
rect -12208 12986 -12140 13020
rect -12050 12986 -11982 13020
rect -11892 12986 -11824 13020
rect -11734 12986 -11666 13020
rect -11576 12986 -11508 13020
rect -11418 12986 -11350 13020
rect -11260 12986 -11192 13020
rect -11102 12986 -11034 13020
rect -10944 12986 -10876 13020
rect -10786 12986 -10718 13020
rect -10628 12986 -10560 13020
rect -10470 12986 -10402 13020
rect -10312 12986 -10244 13020
rect -10154 12986 -10086 13020
rect -9996 12986 -9928 13020
rect -9838 12986 -9770 13020
rect -9680 12986 -9612 13020
rect -9522 12986 -9454 13020
rect -9364 12986 -9296 13020
rect -9206 12986 -9138 13020
rect -9048 12986 -8980 13020
rect -8890 12986 -8822 13020
rect -8732 12986 -8664 13020
rect -8574 12986 -8506 13020
rect -6856 19096 -6788 19130
rect -6698 19096 -6630 19130
rect -6540 19096 -6472 19130
rect -6382 19096 -6314 19130
rect -6224 19096 -6156 19130
rect -6066 19096 -5998 19130
rect -5908 19096 -5840 19130
rect -5750 19096 -5682 19130
rect -5592 19096 -5524 19130
rect -5434 19096 -5366 19130
rect -5276 19096 -5208 19130
rect -5118 19096 -5050 19130
rect -4960 19096 -4892 19130
rect -4802 19096 -4734 19130
rect -4644 19096 -4576 19130
rect -4486 19096 -4418 19130
rect -4328 19096 -4260 19130
rect -4170 19096 -4102 19130
rect -4012 19096 -3944 19130
rect -3854 19096 -3786 19130
rect -3696 19096 -3628 19130
rect -3538 19096 -3470 19130
rect -3380 19096 -3312 19130
rect -3222 19096 -3154 19130
rect -3064 19096 -2996 19130
rect -2906 19096 -2838 19130
rect -2748 19096 -2680 19130
rect -2590 19096 -2522 19130
rect -2432 19096 -2364 19130
rect -2274 19096 -2206 19130
rect -6856 12986 -6788 13020
rect -6698 12986 -6630 13020
rect -6540 12986 -6472 13020
rect -6382 12986 -6314 13020
rect -6224 12986 -6156 13020
rect -6066 12986 -5998 13020
rect -5908 12986 -5840 13020
rect -5750 12986 -5682 13020
rect -5592 12986 -5524 13020
rect -5434 12986 -5366 13020
rect -5276 12986 -5208 13020
rect -5118 12986 -5050 13020
rect -4960 12986 -4892 13020
rect -4802 12986 -4734 13020
rect -4644 12986 -4576 13020
rect -4486 12986 -4418 13020
rect -4328 12986 -4260 13020
rect -4170 12986 -4102 13020
rect -4012 12986 -3944 13020
rect -3854 12986 -3786 13020
rect -3696 12986 -3628 13020
rect -3538 12986 -3470 13020
rect -3380 12986 -3312 13020
rect -3222 12986 -3154 13020
rect -3064 12986 -2996 13020
rect -2906 12986 -2838 13020
rect -2748 12986 -2680 13020
rect -2590 12986 -2522 13020
rect -2432 12986 -2364 13020
rect -2274 12986 -2206 13020
rect -556 19096 -488 19130
rect -398 19096 -330 19130
rect -240 19096 -172 19130
rect -82 19096 -14 19130
rect 76 19096 144 19130
rect 234 19096 302 19130
rect 392 19096 460 19130
rect 550 19096 618 19130
rect 708 19096 776 19130
rect 866 19096 934 19130
rect 1024 19096 1092 19130
rect 1182 19096 1250 19130
rect 1340 19096 1408 19130
rect 1498 19096 1566 19130
rect 1656 19096 1724 19130
rect 1814 19096 1882 19130
rect 1972 19096 2040 19130
rect 2130 19096 2198 19130
rect 2288 19096 2356 19130
rect 2446 19096 2514 19130
rect 2604 19096 2672 19130
rect 2762 19096 2830 19130
rect 2920 19096 2988 19130
rect 3078 19096 3146 19130
rect 3236 19096 3304 19130
rect 3394 19096 3462 19130
rect 3552 19096 3620 19130
rect 3710 19096 3778 19130
rect 3868 19096 3936 19130
rect 4026 19096 4094 19130
rect -556 12986 -488 13020
rect -398 12986 -330 13020
rect -240 12986 -172 13020
rect -82 12986 -14 13020
rect 76 12986 144 13020
rect 234 12986 302 13020
rect 392 12986 460 13020
rect 550 12986 618 13020
rect 708 12986 776 13020
rect 866 12986 934 13020
rect 1024 12986 1092 13020
rect 1182 12986 1250 13020
rect 1340 12986 1408 13020
rect 1498 12986 1566 13020
rect 1656 12986 1724 13020
rect 1814 12986 1882 13020
rect 1972 12986 2040 13020
rect 2130 12986 2198 13020
rect 2288 12986 2356 13020
rect 2446 12986 2514 13020
rect 2604 12986 2672 13020
rect 2762 12986 2830 13020
rect 2920 12986 2988 13020
rect 3078 12986 3146 13020
rect 3236 12986 3304 13020
rect 3394 12986 3462 13020
rect 3552 12986 3620 13020
rect 3710 12986 3778 13020
rect 3868 12986 3936 13020
rect 4026 12986 4094 13020
rect 5744 19096 5812 19130
rect 5902 19096 5970 19130
rect 6060 19096 6128 19130
rect 6218 19096 6286 19130
rect 6376 19096 6444 19130
rect 6534 19096 6602 19130
rect 6692 19096 6760 19130
rect 6850 19096 6918 19130
rect 7008 19096 7076 19130
rect 7166 19096 7234 19130
rect 7324 19096 7392 19130
rect 7482 19096 7550 19130
rect 7640 19096 7708 19130
rect 7798 19096 7866 19130
rect 7956 19096 8024 19130
rect 8114 19096 8182 19130
rect 8272 19096 8340 19130
rect 8430 19096 8498 19130
rect 8588 19096 8656 19130
rect 8746 19096 8814 19130
rect 8904 19096 8972 19130
rect 9062 19096 9130 19130
rect 9220 19096 9288 19130
rect 9378 19096 9446 19130
rect 9536 19096 9604 19130
rect 9694 19096 9762 19130
rect 9852 19096 9920 19130
rect 10010 19096 10078 19130
rect 10168 19096 10236 19130
rect 10326 19096 10394 19130
rect 5744 12986 5812 13020
rect 5902 12986 5970 13020
rect 6060 12986 6128 13020
rect 6218 12986 6286 13020
rect 6376 12986 6444 13020
rect 6534 12986 6602 13020
rect 6692 12986 6760 13020
rect 6850 12986 6918 13020
rect 7008 12986 7076 13020
rect 7166 12986 7234 13020
rect 7324 12986 7392 13020
rect 7482 12986 7550 13020
rect 7640 12986 7708 13020
rect 7798 12986 7866 13020
rect 7956 12986 8024 13020
rect 8114 12986 8182 13020
rect 8272 12986 8340 13020
rect 8430 12986 8498 13020
rect 8588 12986 8656 13020
rect 8746 12986 8814 13020
rect 8904 12986 8972 13020
rect 9062 12986 9130 13020
rect 9220 12986 9288 13020
rect 9378 12986 9446 13020
rect 9536 12986 9604 13020
rect 9694 12986 9762 13020
rect 9852 12986 9920 13020
rect 10010 12986 10078 13020
rect 10168 12986 10236 13020
rect 10326 12986 10394 13020
rect -13156 12096 -13088 12130
rect -12998 12096 -12930 12130
rect -12840 12096 -12772 12130
rect -12682 12096 -12614 12130
rect -12524 12096 -12456 12130
rect -12366 12096 -12298 12130
rect -12208 12096 -12140 12130
rect -12050 12096 -11982 12130
rect -11892 12096 -11824 12130
rect -11734 12096 -11666 12130
rect -11576 12096 -11508 12130
rect -11418 12096 -11350 12130
rect -11260 12096 -11192 12130
rect -11102 12096 -11034 12130
rect -10944 12096 -10876 12130
rect -10786 12096 -10718 12130
rect -10628 12096 -10560 12130
rect -10470 12096 -10402 12130
rect -10312 12096 -10244 12130
rect -10154 12096 -10086 12130
rect -9996 12096 -9928 12130
rect -9838 12096 -9770 12130
rect -9680 12096 -9612 12130
rect -9522 12096 -9454 12130
rect -9364 12096 -9296 12130
rect -9206 12096 -9138 12130
rect -9048 12096 -8980 12130
rect -8890 12096 -8822 12130
rect -8732 12096 -8664 12130
rect -8574 12096 -8506 12130
rect -13156 5986 -13088 6020
rect -12998 5986 -12930 6020
rect -12840 5986 -12772 6020
rect -12682 5986 -12614 6020
rect -12524 5986 -12456 6020
rect -12366 5986 -12298 6020
rect -12208 5986 -12140 6020
rect -12050 5986 -11982 6020
rect -11892 5986 -11824 6020
rect -11734 5986 -11666 6020
rect -11576 5986 -11508 6020
rect -11418 5986 -11350 6020
rect -11260 5986 -11192 6020
rect -11102 5986 -11034 6020
rect -10944 5986 -10876 6020
rect -10786 5986 -10718 6020
rect -10628 5986 -10560 6020
rect -10470 5986 -10402 6020
rect -10312 5986 -10244 6020
rect -10154 5986 -10086 6020
rect -9996 5986 -9928 6020
rect -9838 5986 -9770 6020
rect -9680 5986 -9612 6020
rect -9522 5986 -9454 6020
rect -9364 5986 -9296 6020
rect -9206 5986 -9138 6020
rect -9048 5986 -8980 6020
rect -8890 5986 -8822 6020
rect -8732 5986 -8664 6020
rect -8574 5986 -8506 6020
rect -6856 12096 -6788 12130
rect -6698 12096 -6630 12130
rect -6540 12096 -6472 12130
rect -6382 12096 -6314 12130
rect -6224 12096 -6156 12130
rect -6066 12096 -5998 12130
rect -5908 12096 -5840 12130
rect -5750 12096 -5682 12130
rect -5592 12096 -5524 12130
rect -5434 12096 -5366 12130
rect -5276 12096 -5208 12130
rect -5118 12096 -5050 12130
rect -4960 12096 -4892 12130
rect -4802 12096 -4734 12130
rect -4644 12096 -4576 12130
rect -4486 12096 -4418 12130
rect -4328 12096 -4260 12130
rect -4170 12096 -4102 12130
rect -4012 12096 -3944 12130
rect -3854 12096 -3786 12130
rect -3696 12096 -3628 12130
rect -3538 12096 -3470 12130
rect -3380 12096 -3312 12130
rect -3222 12096 -3154 12130
rect -3064 12096 -2996 12130
rect -2906 12096 -2838 12130
rect -2748 12096 -2680 12130
rect -2590 12096 -2522 12130
rect -2432 12096 -2364 12130
rect -2274 12096 -2206 12130
rect -6856 5986 -6788 6020
rect -6698 5986 -6630 6020
rect -6540 5986 -6472 6020
rect -6382 5986 -6314 6020
rect -6224 5986 -6156 6020
rect -6066 5986 -5998 6020
rect -5908 5986 -5840 6020
rect -5750 5986 -5682 6020
rect -5592 5986 -5524 6020
rect -5434 5986 -5366 6020
rect -5276 5986 -5208 6020
rect -5118 5986 -5050 6020
rect -4960 5986 -4892 6020
rect -4802 5986 -4734 6020
rect -4644 5986 -4576 6020
rect -4486 5986 -4418 6020
rect -4328 5986 -4260 6020
rect -4170 5986 -4102 6020
rect -4012 5986 -3944 6020
rect -3854 5986 -3786 6020
rect -3696 5986 -3628 6020
rect -3538 5986 -3470 6020
rect -3380 5986 -3312 6020
rect -3222 5986 -3154 6020
rect -3064 5986 -2996 6020
rect -2906 5986 -2838 6020
rect -2748 5986 -2680 6020
rect -2590 5986 -2522 6020
rect -2432 5986 -2364 6020
rect -2274 5986 -2206 6020
rect -556 12096 -488 12130
rect -398 12096 -330 12130
rect -240 12096 -172 12130
rect -82 12096 -14 12130
rect 76 12096 144 12130
rect 234 12096 302 12130
rect 392 12096 460 12130
rect 550 12096 618 12130
rect 708 12096 776 12130
rect 866 12096 934 12130
rect 1024 12096 1092 12130
rect 1182 12096 1250 12130
rect 1340 12096 1408 12130
rect 1498 12096 1566 12130
rect 1656 12096 1724 12130
rect 1814 12096 1882 12130
rect 1972 12096 2040 12130
rect 2130 12096 2198 12130
rect 2288 12096 2356 12130
rect 2446 12096 2514 12130
rect 2604 12096 2672 12130
rect 2762 12096 2830 12130
rect 2920 12096 2988 12130
rect 3078 12096 3146 12130
rect 3236 12096 3304 12130
rect 3394 12096 3462 12130
rect 3552 12096 3620 12130
rect 3710 12096 3778 12130
rect 3868 12096 3936 12130
rect 4026 12096 4094 12130
rect -556 5986 -488 6020
rect -398 5986 -330 6020
rect -240 5986 -172 6020
rect -82 5986 -14 6020
rect 76 5986 144 6020
rect 234 5986 302 6020
rect 392 5986 460 6020
rect 550 5986 618 6020
rect 708 5986 776 6020
rect 866 5986 934 6020
rect 1024 5986 1092 6020
rect 1182 5986 1250 6020
rect 1340 5986 1408 6020
rect 1498 5986 1566 6020
rect 1656 5986 1724 6020
rect 1814 5986 1882 6020
rect 1972 5986 2040 6020
rect 2130 5986 2198 6020
rect 2288 5986 2356 6020
rect 2446 5986 2514 6020
rect 2604 5986 2672 6020
rect 2762 5986 2830 6020
rect 2920 5986 2988 6020
rect 3078 5986 3146 6020
rect 3236 5986 3304 6020
rect 3394 5986 3462 6020
rect 3552 5986 3620 6020
rect 3710 5986 3778 6020
rect 3868 5986 3936 6020
rect 4026 5986 4094 6020
rect 5744 12096 5812 12130
rect 5902 12096 5970 12130
rect 6060 12096 6128 12130
rect 6218 12096 6286 12130
rect 6376 12096 6444 12130
rect 6534 12096 6602 12130
rect 6692 12096 6760 12130
rect 6850 12096 6918 12130
rect 7008 12096 7076 12130
rect 7166 12096 7234 12130
rect 7324 12096 7392 12130
rect 7482 12096 7550 12130
rect 7640 12096 7708 12130
rect 7798 12096 7866 12130
rect 7956 12096 8024 12130
rect 8114 12096 8182 12130
rect 8272 12096 8340 12130
rect 8430 12096 8498 12130
rect 8588 12096 8656 12130
rect 8746 12096 8814 12130
rect 8904 12096 8972 12130
rect 9062 12096 9130 12130
rect 9220 12096 9288 12130
rect 9378 12096 9446 12130
rect 9536 12096 9604 12130
rect 9694 12096 9762 12130
rect 9852 12096 9920 12130
rect 10010 12096 10078 12130
rect 10168 12096 10236 12130
rect 10326 12096 10394 12130
rect 5744 5986 5812 6020
rect 5902 5986 5970 6020
rect 6060 5986 6128 6020
rect 6218 5986 6286 6020
rect 6376 5986 6444 6020
rect 6534 5986 6602 6020
rect 6692 5986 6760 6020
rect 6850 5986 6918 6020
rect 7008 5986 7076 6020
rect 7166 5986 7234 6020
rect 7324 5986 7392 6020
rect 7482 5986 7550 6020
rect 7640 5986 7708 6020
rect 7798 5986 7866 6020
rect 7956 5986 8024 6020
rect 8114 5986 8182 6020
rect 8272 5986 8340 6020
rect 8430 5986 8498 6020
rect 8588 5986 8656 6020
rect 8746 5986 8814 6020
rect 8904 5986 8972 6020
rect 9062 5986 9130 6020
rect 9220 5986 9288 6020
rect 9378 5986 9446 6020
rect 9536 5986 9604 6020
rect 9694 5986 9762 6020
rect 9852 5986 9920 6020
rect 10010 5986 10078 6020
rect 10168 5986 10236 6020
rect 10326 5986 10394 6020
<< locali >>
rect -13352 49834 -13256 49868
rect -8406 49834 -8310 49868
rect -13352 49772 -13318 49834
rect -8344 49772 -8310 49834
rect -13172 49696 -13156 49730
rect -13088 49696 -13072 49730
rect -13014 49696 -12998 49730
rect -12930 49696 -12914 49730
rect -12856 49696 -12840 49730
rect -12772 49696 -12756 49730
rect -12698 49696 -12682 49730
rect -12614 49696 -12598 49730
rect -12540 49696 -12524 49730
rect -12456 49696 -12440 49730
rect -12382 49696 -12366 49730
rect -12298 49696 -12282 49730
rect -12224 49696 -12208 49730
rect -12140 49696 -12124 49730
rect -12066 49696 -12050 49730
rect -11982 49696 -11966 49730
rect -11908 49696 -11892 49730
rect -11824 49696 -11808 49730
rect -11750 49696 -11734 49730
rect -11666 49696 -11650 49730
rect -11592 49696 -11576 49730
rect -11508 49696 -11492 49730
rect -11434 49696 -11418 49730
rect -11350 49696 -11334 49730
rect -11276 49696 -11260 49730
rect -11192 49696 -11176 49730
rect -11118 49696 -11102 49730
rect -11034 49696 -11018 49730
rect -10960 49696 -10944 49730
rect -10876 49696 -10860 49730
rect -10802 49696 -10786 49730
rect -10718 49696 -10702 49730
rect -10644 49696 -10628 49730
rect -10560 49696 -10544 49730
rect -10486 49696 -10470 49730
rect -10402 49696 -10386 49730
rect -10328 49696 -10312 49730
rect -10244 49696 -10228 49730
rect -10170 49696 -10154 49730
rect -10086 49696 -10070 49730
rect -10012 49696 -9996 49730
rect -9928 49696 -9912 49730
rect -9854 49696 -9838 49730
rect -9770 49696 -9754 49730
rect -9696 49696 -9680 49730
rect -9612 49696 -9596 49730
rect -9538 49696 -9522 49730
rect -9454 49696 -9438 49730
rect -9380 49696 -9364 49730
rect -9296 49696 -9280 49730
rect -9222 49696 -9206 49730
rect -9138 49696 -9122 49730
rect -9064 49696 -9048 49730
rect -8980 49696 -8964 49730
rect -8906 49696 -8890 49730
rect -8822 49696 -8806 49730
rect -8748 49696 -8732 49730
rect -8664 49696 -8648 49730
rect -8590 49696 -8574 49730
rect -8506 49696 -8490 49730
rect -7052 49834 -6956 49868
rect -2106 49834 -2010 49868
rect -7052 49772 -7018 49834
rect -2044 49772 -2010 49834
rect -6872 49696 -6856 49730
rect -6788 49696 -6772 49730
rect -6714 49696 -6698 49730
rect -6630 49696 -6614 49730
rect -6556 49696 -6540 49730
rect -6472 49696 -6456 49730
rect -6398 49696 -6382 49730
rect -6314 49696 -6298 49730
rect -6240 49696 -6224 49730
rect -6156 49696 -6140 49730
rect -6082 49696 -6066 49730
rect -5998 49696 -5982 49730
rect -5924 49696 -5908 49730
rect -5840 49696 -5824 49730
rect -5766 49696 -5750 49730
rect -5682 49696 -5666 49730
rect -5608 49696 -5592 49730
rect -5524 49696 -5508 49730
rect -5450 49696 -5434 49730
rect -5366 49696 -5350 49730
rect -5292 49696 -5276 49730
rect -5208 49696 -5192 49730
rect -5134 49696 -5118 49730
rect -5050 49696 -5034 49730
rect -4976 49696 -4960 49730
rect -4892 49696 -4876 49730
rect -4818 49696 -4802 49730
rect -4734 49696 -4718 49730
rect -4660 49696 -4644 49730
rect -4576 49696 -4560 49730
rect -4502 49696 -4486 49730
rect -4418 49696 -4402 49730
rect -4344 49696 -4328 49730
rect -4260 49696 -4244 49730
rect -4186 49696 -4170 49730
rect -4102 49696 -4086 49730
rect -4028 49696 -4012 49730
rect -3944 49696 -3928 49730
rect -3870 49696 -3854 49730
rect -3786 49696 -3770 49730
rect -3712 49696 -3696 49730
rect -3628 49696 -3612 49730
rect -3554 49696 -3538 49730
rect -3470 49696 -3454 49730
rect -3396 49696 -3380 49730
rect -3312 49696 -3296 49730
rect -3238 49696 -3222 49730
rect -3154 49696 -3138 49730
rect -3080 49696 -3064 49730
rect -2996 49696 -2980 49730
rect -2922 49696 -2906 49730
rect -2838 49696 -2822 49730
rect -2764 49696 -2748 49730
rect -2680 49696 -2664 49730
rect -2606 49696 -2590 49730
rect -2522 49696 -2506 49730
rect -2448 49696 -2432 49730
rect -2364 49696 -2348 49730
rect -2290 49696 -2274 49730
rect -2206 49696 -2190 49730
rect -752 49834 -656 49868
rect 4194 49834 4290 49868
rect -752 49772 -718 49834
rect 4256 49772 4290 49834
rect -572 49696 -556 49730
rect -488 49696 -472 49730
rect -414 49696 -398 49730
rect -330 49696 -314 49730
rect -256 49696 -240 49730
rect -172 49696 -156 49730
rect -98 49696 -82 49730
rect -14 49696 2 49730
rect 60 49696 76 49730
rect 144 49696 160 49730
rect 218 49696 234 49730
rect 302 49696 318 49730
rect 376 49696 392 49730
rect 460 49696 476 49730
rect 534 49696 550 49730
rect 618 49696 634 49730
rect 692 49696 708 49730
rect 776 49696 792 49730
rect 850 49696 866 49730
rect 934 49696 950 49730
rect 1008 49696 1024 49730
rect 1092 49696 1108 49730
rect 1166 49696 1182 49730
rect 1250 49696 1266 49730
rect 1324 49696 1340 49730
rect 1408 49696 1424 49730
rect 1482 49696 1498 49730
rect 1566 49696 1582 49730
rect 1640 49696 1656 49730
rect 1724 49696 1740 49730
rect 1798 49696 1814 49730
rect 1882 49696 1898 49730
rect 1956 49696 1972 49730
rect 2040 49696 2056 49730
rect 2114 49696 2130 49730
rect 2198 49696 2214 49730
rect 2272 49696 2288 49730
rect 2356 49696 2372 49730
rect 2430 49696 2446 49730
rect 2514 49696 2530 49730
rect 2588 49696 2604 49730
rect 2672 49696 2688 49730
rect 2746 49696 2762 49730
rect 2830 49696 2846 49730
rect 2904 49696 2920 49730
rect 2988 49696 3004 49730
rect 3062 49696 3078 49730
rect 3146 49696 3162 49730
rect 3220 49696 3236 49730
rect 3304 49696 3320 49730
rect 3378 49696 3394 49730
rect 3462 49696 3478 49730
rect 3536 49696 3552 49730
rect 3620 49696 3636 49730
rect 3694 49696 3710 49730
rect 3778 49696 3794 49730
rect 3852 49696 3868 49730
rect 3936 49696 3952 49730
rect 4010 49696 4026 49730
rect 4094 49696 4110 49730
rect 5548 49834 5644 49868
rect 10494 49834 10590 49868
rect 5548 49772 5582 49834
rect 10556 49772 10590 49834
rect 5728 49696 5744 49730
rect 5812 49696 5828 49730
rect 5886 49696 5902 49730
rect 5970 49696 5986 49730
rect 6044 49696 6060 49730
rect 6128 49696 6144 49730
rect 6202 49696 6218 49730
rect 6286 49696 6302 49730
rect 6360 49696 6376 49730
rect 6444 49696 6460 49730
rect 6518 49696 6534 49730
rect 6602 49696 6618 49730
rect 6676 49696 6692 49730
rect 6760 49696 6776 49730
rect 6834 49696 6850 49730
rect 6918 49696 6934 49730
rect 6992 49696 7008 49730
rect 7076 49696 7092 49730
rect 7150 49696 7166 49730
rect 7234 49696 7250 49730
rect 7308 49696 7324 49730
rect 7392 49696 7408 49730
rect 7466 49696 7482 49730
rect 7550 49696 7566 49730
rect 7624 49696 7640 49730
rect 7708 49696 7724 49730
rect 7782 49696 7798 49730
rect 7866 49696 7882 49730
rect 7940 49696 7956 49730
rect 8024 49696 8040 49730
rect 8098 49696 8114 49730
rect 8182 49696 8198 49730
rect 8256 49696 8272 49730
rect 8340 49696 8356 49730
rect 8414 49696 8430 49730
rect 8498 49696 8514 49730
rect 8572 49696 8588 49730
rect 8656 49696 8672 49730
rect 8730 49696 8746 49730
rect 8814 49696 8830 49730
rect 8888 49696 8904 49730
rect 8972 49696 8988 49730
rect 9046 49696 9062 49730
rect 9130 49696 9146 49730
rect 9204 49696 9220 49730
rect 9288 49696 9304 49730
rect 9362 49696 9378 49730
rect 9446 49696 9462 49730
rect 9520 49696 9536 49730
rect 9604 49696 9620 49730
rect 9678 49696 9694 49730
rect 9762 49696 9778 49730
rect 9836 49696 9852 49730
rect 9920 49696 9936 49730
rect 9994 49696 10010 49730
rect 10078 49696 10094 49730
rect 10152 49696 10168 49730
rect 10236 49696 10252 49730
rect 10310 49696 10326 49730
rect 10394 49696 10410 49730
rect -13218 49646 -13184 49662
rect -13218 43654 -13184 43670
rect -13060 49646 -13026 49662
rect -13060 43654 -13026 43670
rect -12902 49646 -12868 49662
rect -12902 43654 -12868 43670
rect -12744 49646 -12710 49662
rect -12744 43654 -12710 43670
rect -12586 49646 -12552 49662
rect -12586 43654 -12552 43670
rect -12428 49646 -12394 49662
rect -12428 43654 -12394 43670
rect -12270 49646 -12236 49662
rect -12270 43654 -12236 43670
rect -12112 49646 -12078 49662
rect -12112 43654 -12078 43670
rect -11954 49646 -11920 49662
rect -11954 43654 -11920 43670
rect -11796 49646 -11762 49662
rect -11796 43654 -11762 43670
rect -11638 49646 -11604 49662
rect -11638 43654 -11604 43670
rect -11480 49646 -11446 49662
rect -11480 43654 -11446 43670
rect -11322 49646 -11288 49662
rect -11322 43654 -11288 43670
rect -11164 49646 -11130 49662
rect -11164 43654 -11130 43670
rect -11006 49646 -10972 49662
rect -11006 43654 -10972 43670
rect -10848 49646 -10814 49662
rect -10848 43654 -10814 43670
rect -10690 49646 -10656 49662
rect -10690 43654 -10656 43670
rect -10532 49646 -10498 49662
rect -10532 43654 -10498 43670
rect -10374 49646 -10340 49662
rect -10374 43654 -10340 43670
rect -10216 49646 -10182 49662
rect -10216 43654 -10182 43670
rect -10058 49646 -10024 49662
rect -10058 43654 -10024 43670
rect -9900 49646 -9866 49662
rect -9900 43654 -9866 43670
rect -9742 49646 -9708 49662
rect -9742 43654 -9708 43670
rect -9584 49646 -9550 49662
rect -9584 43654 -9550 43670
rect -9426 49646 -9392 49662
rect -9426 43654 -9392 43670
rect -9268 49646 -9234 49662
rect -9268 43654 -9234 43670
rect -9110 49646 -9076 49662
rect -9110 43654 -9076 43670
rect -8952 49646 -8918 49662
rect -8952 43654 -8918 43670
rect -8794 49646 -8760 49662
rect -8794 43654 -8760 43670
rect -8636 49646 -8602 49662
rect -8636 43654 -8602 43670
rect -8478 49646 -8444 49662
rect -8478 43654 -8444 43670
rect -6918 49646 -6884 49662
rect -6918 43654 -6884 43670
rect -6760 49646 -6726 49662
rect -6760 43654 -6726 43670
rect -6602 49646 -6568 49662
rect -6602 43654 -6568 43670
rect -6444 49646 -6410 49662
rect -6444 43654 -6410 43670
rect -6286 49646 -6252 49662
rect -6286 43654 -6252 43670
rect -6128 49646 -6094 49662
rect -6128 43654 -6094 43670
rect -5970 49646 -5936 49662
rect -5970 43654 -5936 43670
rect -5812 49646 -5778 49662
rect -5812 43654 -5778 43670
rect -5654 49646 -5620 49662
rect -5654 43654 -5620 43670
rect -5496 49646 -5462 49662
rect -5496 43654 -5462 43670
rect -5338 49646 -5304 49662
rect -5338 43654 -5304 43670
rect -5180 49646 -5146 49662
rect -5180 43654 -5146 43670
rect -5022 49646 -4988 49662
rect -5022 43654 -4988 43670
rect -4864 49646 -4830 49662
rect -4864 43654 -4830 43670
rect -4706 49646 -4672 49662
rect -4706 43654 -4672 43670
rect -4548 49646 -4514 49662
rect -4548 43654 -4514 43670
rect -4390 49646 -4356 49662
rect -4390 43654 -4356 43670
rect -4232 49646 -4198 49662
rect -4232 43654 -4198 43670
rect -4074 49646 -4040 49662
rect -4074 43654 -4040 43670
rect -3916 49646 -3882 49662
rect -3916 43654 -3882 43670
rect -3758 49646 -3724 49662
rect -3758 43654 -3724 43670
rect -3600 49646 -3566 49662
rect -3600 43654 -3566 43670
rect -3442 49646 -3408 49662
rect -3442 43654 -3408 43670
rect -3284 49646 -3250 49662
rect -3284 43654 -3250 43670
rect -3126 49646 -3092 49662
rect -3126 43654 -3092 43670
rect -2968 49646 -2934 49662
rect -2968 43654 -2934 43670
rect -2810 49646 -2776 49662
rect -2810 43654 -2776 43670
rect -2652 49646 -2618 49662
rect -2652 43654 -2618 43670
rect -2494 49646 -2460 49662
rect -2494 43654 -2460 43670
rect -2336 49646 -2302 49662
rect -2336 43654 -2302 43670
rect -2178 49646 -2144 49662
rect -2178 43654 -2144 43670
rect -618 49646 -584 49662
rect -618 43654 -584 43670
rect -460 49646 -426 49662
rect -460 43654 -426 43670
rect -302 49646 -268 49662
rect -302 43654 -268 43670
rect -144 49646 -110 49662
rect -144 43654 -110 43670
rect 14 49646 48 49662
rect 14 43654 48 43670
rect 172 49646 206 49662
rect 172 43654 206 43670
rect 330 49646 364 49662
rect 330 43654 364 43670
rect 488 49646 522 49662
rect 488 43654 522 43670
rect 646 49646 680 49662
rect 646 43654 680 43670
rect 804 49646 838 49662
rect 804 43654 838 43670
rect 962 49646 996 49662
rect 962 43654 996 43670
rect 1120 49646 1154 49662
rect 1120 43654 1154 43670
rect 1278 49646 1312 49662
rect 1278 43654 1312 43670
rect 1436 49646 1470 49662
rect 1436 43654 1470 43670
rect 1594 49646 1628 49662
rect 1594 43654 1628 43670
rect 1752 49646 1786 49662
rect 1752 43654 1786 43670
rect 1910 49646 1944 49662
rect 1910 43654 1944 43670
rect 2068 49646 2102 49662
rect 2068 43654 2102 43670
rect 2226 49646 2260 49662
rect 2226 43654 2260 43670
rect 2384 49646 2418 49662
rect 2384 43654 2418 43670
rect 2542 49646 2576 49662
rect 2542 43654 2576 43670
rect 2700 49646 2734 49662
rect 2700 43654 2734 43670
rect 2858 49646 2892 49662
rect 2858 43654 2892 43670
rect 3016 49646 3050 49662
rect 3016 43654 3050 43670
rect 3174 49646 3208 49662
rect 3174 43654 3208 43670
rect 3332 49646 3366 49662
rect 3332 43654 3366 43670
rect 3490 49646 3524 49662
rect 3490 43654 3524 43670
rect 3648 49646 3682 49662
rect 3648 43654 3682 43670
rect 3806 49646 3840 49662
rect 3806 43654 3840 43670
rect 3964 49646 3998 49662
rect 3964 43654 3998 43670
rect 4122 49646 4156 49662
rect 4122 43654 4156 43670
rect 5682 49646 5716 49662
rect 5682 43654 5716 43670
rect 5840 49646 5874 49662
rect 5840 43654 5874 43670
rect 5998 49646 6032 49662
rect 5998 43654 6032 43670
rect 6156 49646 6190 49662
rect 6156 43654 6190 43670
rect 6314 49646 6348 49662
rect 6314 43654 6348 43670
rect 6472 49646 6506 49662
rect 6472 43654 6506 43670
rect 6630 49646 6664 49662
rect 6630 43654 6664 43670
rect 6788 49646 6822 49662
rect 6788 43654 6822 43670
rect 6946 49646 6980 49662
rect 6946 43654 6980 43670
rect 7104 49646 7138 49662
rect 7104 43654 7138 43670
rect 7262 49646 7296 49662
rect 7262 43654 7296 43670
rect 7420 49646 7454 49662
rect 7420 43654 7454 43670
rect 7578 49646 7612 49662
rect 7578 43654 7612 43670
rect 7736 49646 7770 49662
rect 7736 43654 7770 43670
rect 7894 49646 7928 49662
rect 7894 43654 7928 43670
rect 8052 49646 8086 49662
rect 8052 43654 8086 43670
rect 8210 49646 8244 49662
rect 8210 43654 8244 43670
rect 8368 49646 8402 49662
rect 8368 43654 8402 43670
rect 8526 49646 8560 49662
rect 8526 43654 8560 43670
rect 8684 49646 8718 49662
rect 8684 43654 8718 43670
rect 8842 49646 8876 49662
rect 8842 43654 8876 43670
rect 9000 49646 9034 49662
rect 9000 43654 9034 43670
rect 9158 49646 9192 49662
rect 9158 43654 9192 43670
rect 9316 49646 9350 49662
rect 9316 43654 9350 43670
rect 9474 49646 9508 49662
rect 9474 43654 9508 43670
rect 9632 49646 9666 49662
rect 9632 43654 9666 43670
rect 9790 49646 9824 49662
rect 9790 43654 9824 43670
rect 9948 49646 9982 49662
rect 9948 43654 9982 43670
rect 10106 49646 10140 49662
rect 10106 43654 10140 43670
rect 10264 49646 10298 49662
rect 10264 43654 10298 43670
rect 10422 49646 10456 49662
rect 10422 43654 10456 43670
rect -13172 43586 -13156 43620
rect -13088 43586 -13072 43620
rect -13014 43586 -12998 43620
rect -12930 43586 -12914 43620
rect -12856 43586 -12840 43620
rect -12772 43586 -12756 43620
rect -12698 43586 -12682 43620
rect -12614 43586 -12598 43620
rect -12540 43586 -12524 43620
rect -12456 43586 -12440 43620
rect -12382 43586 -12366 43620
rect -12298 43586 -12282 43620
rect -12224 43586 -12208 43620
rect -12140 43586 -12124 43620
rect -12066 43586 -12050 43620
rect -11982 43586 -11966 43620
rect -11908 43586 -11892 43620
rect -11824 43586 -11808 43620
rect -11750 43586 -11734 43620
rect -11666 43586 -11650 43620
rect -11592 43586 -11576 43620
rect -11508 43586 -11492 43620
rect -11434 43586 -11418 43620
rect -11350 43586 -11334 43620
rect -11276 43586 -11260 43620
rect -11192 43586 -11176 43620
rect -11118 43586 -11102 43620
rect -11034 43586 -11018 43620
rect -10960 43586 -10944 43620
rect -10876 43586 -10860 43620
rect -10802 43586 -10786 43620
rect -10718 43586 -10702 43620
rect -10644 43586 -10628 43620
rect -10560 43586 -10544 43620
rect -10486 43586 -10470 43620
rect -10402 43586 -10386 43620
rect -10328 43586 -10312 43620
rect -10244 43586 -10228 43620
rect -10170 43586 -10154 43620
rect -10086 43586 -10070 43620
rect -10012 43586 -9996 43620
rect -9928 43586 -9912 43620
rect -9854 43586 -9838 43620
rect -9770 43586 -9754 43620
rect -9696 43586 -9680 43620
rect -9612 43586 -9596 43620
rect -9538 43586 -9522 43620
rect -9454 43586 -9438 43620
rect -9380 43586 -9364 43620
rect -9296 43586 -9280 43620
rect -9222 43586 -9206 43620
rect -9138 43586 -9122 43620
rect -9064 43586 -9048 43620
rect -8980 43586 -8964 43620
rect -8906 43586 -8890 43620
rect -8822 43586 -8806 43620
rect -8748 43586 -8732 43620
rect -8664 43586 -8648 43620
rect -8590 43586 -8574 43620
rect -8506 43586 -8490 43620
rect -13352 43482 -13318 43544
rect -8344 43482 -8310 43544
rect -13352 43448 -13256 43482
rect -8406 43448 -8310 43482
rect -6872 43586 -6856 43620
rect -6788 43586 -6772 43620
rect -6714 43586 -6698 43620
rect -6630 43586 -6614 43620
rect -6556 43586 -6540 43620
rect -6472 43586 -6456 43620
rect -6398 43586 -6382 43620
rect -6314 43586 -6298 43620
rect -6240 43586 -6224 43620
rect -6156 43586 -6140 43620
rect -6082 43586 -6066 43620
rect -5998 43586 -5982 43620
rect -5924 43586 -5908 43620
rect -5840 43586 -5824 43620
rect -5766 43586 -5750 43620
rect -5682 43586 -5666 43620
rect -5608 43586 -5592 43620
rect -5524 43586 -5508 43620
rect -5450 43586 -5434 43620
rect -5366 43586 -5350 43620
rect -5292 43586 -5276 43620
rect -5208 43586 -5192 43620
rect -5134 43586 -5118 43620
rect -5050 43586 -5034 43620
rect -4976 43586 -4960 43620
rect -4892 43586 -4876 43620
rect -4818 43586 -4802 43620
rect -4734 43586 -4718 43620
rect -4660 43586 -4644 43620
rect -4576 43586 -4560 43620
rect -4502 43586 -4486 43620
rect -4418 43586 -4402 43620
rect -4344 43586 -4328 43620
rect -4260 43586 -4244 43620
rect -4186 43586 -4170 43620
rect -4102 43586 -4086 43620
rect -4028 43586 -4012 43620
rect -3944 43586 -3928 43620
rect -3870 43586 -3854 43620
rect -3786 43586 -3770 43620
rect -3712 43586 -3696 43620
rect -3628 43586 -3612 43620
rect -3554 43586 -3538 43620
rect -3470 43586 -3454 43620
rect -3396 43586 -3380 43620
rect -3312 43586 -3296 43620
rect -3238 43586 -3222 43620
rect -3154 43586 -3138 43620
rect -3080 43586 -3064 43620
rect -2996 43586 -2980 43620
rect -2922 43586 -2906 43620
rect -2838 43586 -2822 43620
rect -2764 43586 -2748 43620
rect -2680 43586 -2664 43620
rect -2606 43586 -2590 43620
rect -2522 43586 -2506 43620
rect -2448 43586 -2432 43620
rect -2364 43586 -2348 43620
rect -2290 43586 -2274 43620
rect -2206 43586 -2190 43620
rect -7052 43482 -7018 43544
rect -2044 43482 -2010 43544
rect -7052 43448 -6956 43482
rect -2106 43448 -2010 43482
rect -572 43586 -556 43620
rect -488 43586 -472 43620
rect -414 43586 -398 43620
rect -330 43586 -314 43620
rect -256 43586 -240 43620
rect -172 43586 -156 43620
rect -98 43586 -82 43620
rect -14 43586 2 43620
rect 60 43586 76 43620
rect 144 43586 160 43620
rect 218 43586 234 43620
rect 302 43586 318 43620
rect 376 43586 392 43620
rect 460 43586 476 43620
rect 534 43586 550 43620
rect 618 43586 634 43620
rect 692 43586 708 43620
rect 776 43586 792 43620
rect 850 43586 866 43620
rect 934 43586 950 43620
rect 1008 43586 1024 43620
rect 1092 43586 1108 43620
rect 1166 43586 1182 43620
rect 1250 43586 1266 43620
rect 1324 43586 1340 43620
rect 1408 43586 1424 43620
rect 1482 43586 1498 43620
rect 1566 43586 1582 43620
rect 1640 43586 1656 43620
rect 1724 43586 1740 43620
rect 1798 43586 1814 43620
rect 1882 43586 1898 43620
rect 1956 43586 1972 43620
rect 2040 43586 2056 43620
rect 2114 43586 2130 43620
rect 2198 43586 2214 43620
rect 2272 43586 2288 43620
rect 2356 43586 2372 43620
rect 2430 43586 2446 43620
rect 2514 43586 2530 43620
rect 2588 43586 2604 43620
rect 2672 43586 2688 43620
rect 2746 43586 2762 43620
rect 2830 43586 2846 43620
rect 2904 43586 2920 43620
rect 2988 43586 3004 43620
rect 3062 43586 3078 43620
rect 3146 43586 3162 43620
rect 3220 43586 3236 43620
rect 3304 43586 3320 43620
rect 3378 43586 3394 43620
rect 3462 43586 3478 43620
rect 3536 43586 3552 43620
rect 3620 43586 3636 43620
rect 3694 43586 3710 43620
rect 3778 43586 3794 43620
rect 3852 43586 3868 43620
rect 3936 43586 3952 43620
rect 4010 43586 4026 43620
rect 4094 43586 4110 43620
rect -752 43482 -718 43544
rect 4256 43482 4290 43544
rect -752 43448 -656 43482
rect 4194 43448 4290 43482
rect 5728 43586 5744 43620
rect 5812 43586 5828 43620
rect 5886 43586 5902 43620
rect 5970 43586 5986 43620
rect 6044 43586 6060 43620
rect 6128 43586 6144 43620
rect 6202 43586 6218 43620
rect 6286 43586 6302 43620
rect 6360 43586 6376 43620
rect 6444 43586 6460 43620
rect 6518 43586 6534 43620
rect 6602 43586 6618 43620
rect 6676 43586 6692 43620
rect 6760 43586 6776 43620
rect 6834 43586 6850 43620
rect 6918 43586 6934 43620
rect 6992 43586 7008 43620
rect 7076 43586 7092 43620
rect 7150 43586 7166 43620
rect 7234 43586 7250 43620
rect 7308 43586 7324 43620
rect 7392 43586 7408 43620
rect 7466 43586 7482 43620
rect 7550 43586 7566 43620
rect 7624 43586 7640 43620
rect 7708 43586 7724 43620
rect 7782 43586 7798 43620
rect 7866 43586 7882 43620
rect 7940 43586 7956 43620
rect 8024 43586 8040 43620
rect 8098 43586 8114 43620
rect 8182 43586 8198 43620
rect 8256 43586 8272 43620
rect 8340 43586 8356 43620
rect 8414 43586 8430 43620
rect 8498 43586 8514 43620
rect 8572 43586 8588 43620
rect 8656 43586 8672 43620
rect 8730 43586 8746 43620
rect 8814 43586 8830 43620
rect 8888 43586 8904 43620
rect 8972 43586 8988 43620
rect 9046 43586 9062 43620
rect 9130 43586 9146 43620
rect 9204 43586 9220 43620
rect 9288 43586 9304 43620
rect 9362 43586 9378 43620
rect 9446 43586 9462 43620
rect 9520 43586 9536 43620
rect 9604 43586 9620 43620
rect 9678 43586 9694 43620
rect 9762 43586 9778 43620
rect 9836 43586 9852 43620
rect 9920 43586 9936 43620
rect 9994 43586 10010 43620
rect 10078 43586 10094 43620
rect 10152 43586 10168 43620
rect 10236 43586 10252 43620
rect 10310 43586 10326 43620
rect 10394 43586 10410 43620
rect 5548 43482 5582 43544
rect 10556 43482 10590 43544
rect 5548 43448 5644 43482
rect 10494 43448 10590 43482
rect -13352 42834 -13256 42868
rect -8406 42834 -8310 42868
rect -13352 42772 -13318 42834
rect -8344 42772 -8310 42834
rect -13172 42696 -13156 42730
rect -13088 42696 -13072 42730
rect -13014 42696 -12998 42730
rect -12930 42696 -12914 42730
rect -12856 42696 -12840 42730
rect -12772 42696 -12756 42730
rect -12698 42696 -12682 42730
rect -12614 42696 -12598 42730
rect -12540 42696 -12524 42730
rect -12456 42696 -12440 42730
rect -12382 42696 -12366 42730
rect -12298 42696 -12282 42730
rect -12224 42696 -12208 42730
rect -12140 42696 -12124 42730
rect -12066 42696 -12050 42730
rect -11982 42696 -11966 42730
rect -11908 42696 -11892 42730
rect -11824 42696 -11808 42730
rect -11750 42696 -11734 42730
rect -11666 42696 -11650 42730
rect -11592 42696 -11576 42730
rect -11508 42696 -11492 42730
rect -11434 42696 -11418 42730
rect -11350 42696 -11334 42730
rect -11276 42696 -11260 42730
rect -11192 42696 -11176 42730
rect -11118 42696 -11102 42730
rect -11034 42696 -11018 42730
rect -10960 42696 -10944 42730
rect -10876 42696 -10860 42730
rect -10802 42696 -10786 42730
rect -10718 42696 -10702 42730
rect -10644 42696 -10628 42730
rect -10560 42696 -10544 42730
rect -10486 42696 -10470 42730
rect -10402 42696 -10386 42730
rect -10328 42696 -10312 42730
rect -10244 42696 -10228 42730
rect -10170 42696 -10154 42730
rect -10086 42696 -10070 42730
rect -10012 42696 -9996 42730
rect -9928 42696 -9912 42730
rect -9854 42696 -9838 42730
rect -9770 42696 -9754 42730
rect -9696 42696 -9680 42730
rect -9612 42696 -9596 42730
rect -9538 42696 -9522 42730
rect -9454 42696 -9438 42730
rect -9380 42696 -9364 42730
rect -9296 42696 -9280 42730
rect -9222 42696 -9206 42730
rect -9138 42696 -9122 42730
rect -9064 42696 -9048 42730
rect -8980 42696 -8964 42730
rect -8906 42696 -8890 42730
rect -8822 42696 -8806 42730
rect -8748 42696 -8732 42730
rect -8664 42696 -8648 42730
rect -8590 42696 -8574 42730
rect -8506 42696 -8490 42730
rect -7052 42834 -6956 42868
rect -2106 42834 -2010 42868
rect -7052 42772 -7018 42834
rect -2044 42772 -2010 42834
rect -6872 42696 -6856 42730
rect -6788 42696 -6772 42730
rect -6714 42696 -6698 42730
rect -6630 42696 -6614 42730
rect -6556 42696 -6540 42730
rect -6472 42696 -6456 42730
rect -6398 42696 -6382 42730
rect -6314 42696 -6298 42730
rect -6240 42696 -6224 42730
rect -6156 42696 -6140 42730
rect -6082 42696 -6066 42730
rect -5998 42696 -5982 42730
rect -5924 42696 -5908 42730
rect -5840 42696 -5824 42730
rect -5766 42696 -5750 42730
rect -5682 42696 -5666 42730
rect -5608 42696 -5592 42730
rect -5524 42696 -5508 42730
rect -5450 42696 -5434 42730
rect -5366 42696 -5350 42730
rect -5292 42696 -5276 42730
rect -5208 42696 -5192 42730
rect -5134 42696 -5118 42730
rect -5050 42696 -5034 42730
rect -4976 42696 -4960 42730
rect -4892 42696 -4876 42730
rect -4818 42696 -4802 42730
rect -4734 42696 -4718 42730
rect -4660 42696 -4644 42730
rect -4576 42696 -4560 42730
rect -4502 42696 -4486 42730
rect -4418 42696 -4402 42730
rect -4344 42696 -4328 42730
rect -4260 42696 -4244 42730
rect -4186 42696 -4170 42730
rect -4102 42696 -4086 42730
rect -4028 42696 -4012 42730
rect -3944 42696 -3928 42730
rect -3870 42696 -3854 42730
rect -3786 42696 -3770 42730
rect -3712 42696 -3696 42730
rect -3628 42696 -3612 42730
rect -3554 42696 -3538 42730
rect -3470 42696 -3454 42730
rect -3396 42696 -3380 42730
rect -3312 42696 -3296 42730
rect -3238 42696 -3222 42730
rect -3154 42696 -3138 42730
rect -3080 42696 -3064 42730
rect -2996 42696 -2980 42730
rect -2922 42696 -2906 42730
rect -2838 42696 -2822 42730
rect -2764 42696 -2748 42730
rect -2680 42696 -2664 42730
rect -2606 42696 -2590 42730
rect -2522 42696 -2506 42730
rect -2448 42696 -2432 42730
rect -2364 42696 -2348 42730
rect -2290 42696 -2274 42730
rect -2206 42696 -2190 42730
rect -752 42834 -656 42868
rect 4194 42834 4290 42868
rect -752 42772 -718 42834
rect 4256 42772 4290 42834
rect -572 42696 -556 42730
rect -488 42696 -472 42730
rect -414 42696 -398 42730
rect -330 42696 -314 42730
rect -256 42696 -240 42730
rect -172 42696 -156 42730
rect -98 42696 -82 42730
rect -14 42696 2 42730
rect 60 42696 76 42730
rect 144 42696 160 42730
rect 218 42696 234 42730
rect 302 42696 318 42730
rect 376 42696 392 42730
rect 460 42696 476 42730
rect 534 42696 550 42730
rect 618 42696 634 42730
rect 692 42696 708 42730
rect 776 42696 792 42730
rect 850 42696 866 42730
rect 934 42696 950 42730
rect 1008 42696 1024 42730
rect 1092 42696 1108 42730
rect 1166 42696 1182 42730
rect 1250 42696 1266 42730
rect 1324 42696 1340 42730
rect 1408 42696 1424 42730
rect 1482 42696 1498 42730
rect 1566 42696 1582 42730
rect 1640 42696 1656 42730
rect 1724 42696 1740 42730
rect 1798 42696 1814 42730
rect 1882 42696 1898 42730
rect 1956 42696 1972 42730
rect 2040 42696 2056 42730
rect 2114 42696 2130 42730
rect 2198 42696 2214 42730
rect 2272 42696 2288 42730
rect 2356 42696 2372 42730
rect 2430 42696 2446 42730
rect 2514 42696 2530 42730
rect 2588 42696 2604 42730
rect 2672 42696 2688 42730
rect 2746 42696 2762 42730
rect 2830 42696 2846 42730
rect 2904 42696 2920 42730
rect 2988 42696 3004 42730
rect 3062 42696 3078 42730
rect 3146 42696 3162 42730
rect 3220 42696 3236 42730
rect 3304 42696 3320 42730
rect 3378 42696 3394 42730
rect 3462 42696 3478 42730
rect 3536 42696 3552 42730
rect 3620 42696 3636 42730
rect 3694 42696 3710 42730
rect 3778 42696 3794 42730
rect 3852 42696 3868 42730
rect 3936 42696 3952 42730
rect 4010 42696 4026 42730
rect 4094 42696 4110 42730
rect 5548 42834 5644 42868
rect 10494 42834 10590 42868
rect 5548 42772 5582 42834
rect 10556 42772 10590 42834
rect 5728 42696 5744 42730
rect 5812 42696 5828 42730
rect 5886 42696 5902 42730
rect 5970 42696 5986 42730
rect 6044 42696 6060 42730
rect 6128 42696 6144 42730
rect 6202 42696 6218 42730
rect 6286 42696 6302 42730
rect 6360 42696 6376 42730
rect 6444 42696 6460 42730
rect 6518 42696 6534 42730
rect 6602 42696 6618 42730
rect 6676 42696 6692 42730
rect 6760 42696 6776 42730
rect 6834 42696 6850 42730
rect 6918 42696 6934 42730
rect 6992 42696 7008 42730
rect 7076 42696 7092 42730
rect 7150 42696 7166 42730
rect 7234 42696 7250 42730
rect 7308 42696 7324 42730
rect 7392 42696 7408 42730
rect 7466 42696 7482 42730
rect 7550 42696 7566 42730
rect 7624 42696 7640 42730
rect 7708 42696 7724 42730
rect 7782 42696 7798 42730
rect 7866 42696 7882 42730
rect 7940 42696 7956 42730
rect 8024 42696 8040 42730
rect 8098 42696 8114 42730
rect 8182 42696 8198 42730
rect 8256 42696 8272 42730
rect 8340 42696 8356 42730
rect 8414 42696 8430 42730
rect 8498 42696 8514 42730
rect 8572 42696 8588 42730
rect 8656 42696 8672 42730
rect 8730 42696 8746 42730
rect 8814 42696 8830 42730
rect 8888 42696 8904 42730
rect 8972 42696 8988 42730
rect 9046 42696 9062 42730
rect 9130 42696 9146 42730
rect 9204 42696 9220 42730
rect 9288 42696 9304 42730
rect 9362 42696 9378 42730
rect 9446 42696 9462 42730
rect 9520 42696 9536 42730
rect 9604 42696 9620 42730
rect 9678 42696 9694 42730
rect 9762 42696 9778 42730
rect 9836 42696 9852 42730
rect 9920 42696 9936 42730
rect 9994 42696 10010 42730
rect 10078 42696 10094 42730
rect 10152 42696 10168 42730
rect 10236 42696 10252 42730
rect 10310 42696 10326 42730
rect 10394 42696 10410 42730
rect -13218 42646 -13184 42662
rect -13218 36654 -13184 36670
rect -13060 42646 -13026 42662
rect -13060 36654 -13026 36670
rect -12902 42646 -12868 42662
rect -12902 36654 -12868 36670
rect -12744 42646 -12710 42662
rect -12744 36654 -12710 36670
rect -12586 42646 -12552 42662
rect -12586 36654 -12552 36670
rect -12428 42646 -12394 42662
rect -12428 36654 -12394 36670
rect -12270 42646 -12236 42662
rect -12270 36654 -12236 36670
rect -12112 42646 -12078 42662
rect -12112 36654 -12078 36670
rect -11954 42646 -11920 42662
rect -11954 36654 -11920 36670
rect -11796 42646 -11762 42662
rect -11796 36654 -11762 36670
rect -11638 42646 -11604 42662
rect -11638 36654 -11604 36670
rect -11480 42646 -11446 42662
rect -11480 36654 -11446 36670
rect -11322 42646 -11288 42662
rect -11322 36654 -11288 36670
rect -11164 42646 -11130 42662
rect -11164 36654 -11130 36670
rect -11006 42646 -10972 42662
rect -11006 36654 -10972 36670
rect -10848 42646 -10814 42662
rect -10848 36654 -10814 36670
rect -10690 42646 -10656 42662
rect -10690 36654 -10656 36670
rect -10532 42646 -10498 42662
rect -10532 36654 -10498 36670
rect -10374 42646 -10340 42662
rect -10374 36654 -10340 36670
rect -10216 42646 -10182 42662
rect -10216 36654 -10182 36670
rect -10058 42646 -10024 42662
rect -10058 36654 -10024 36670
rect -9900 42646 -9866 42662
rect -9900 36654 -9866 36670
rect -9742 42646 -9708 42662
rect -9742 36654 -9708 36670
rect -9584 42646 -9550 42662
rect -9584 36654 -9550 36670
rect -9426 42646 -9392 42662
rect -9426 36654 -9392 36670
rect -9268 42646 -9234 42662
rect -9268 36654 -9234 36670
rect -9110 42646 -9076 42662
rect -9110 36654 -9076 36670
rect -8952 42646 -8918 42662
rect -8952 36654 -8918 36670
rect -8794 42646 -8760 42662
rect -8794 36654 -8760 36670
rect -8636 42646 -8602 42662
rect -8636 36654 -8602 36670
rect -8478 42646 -8444 42662
rect -8478 36654 -8444 36670
rect -6918 42646 -6884 42662
rect -6918 36654 -6884 36670
rect -6760 42646 -6726 42662
rect -6760 36654 -6726 36670
rect -6602 42646 -6568 42662
rect -6602 36654 -6568 36670
rect -6444 42646 -6410 42662
rect -6444 36654 -6410 36670
rect -6286 42646 -6252 42662
rect -6286 36654 -6252 36670
rect -6128 42646 -6094 42662
rect -6128 36654 -6094 36670
rect -5970 42646 -5936 42662
rect -5970 36654 -5936 36670
rect -5812 42646 -5778 42662
rect -5812 36654 -5778 36670
rect -5654 42646 -5620 42662
rect -5654 36654 -5620 36670
rect -5496 42646 -5462 42662
rect -5496 36654 -5462 36670
rect -5338 42646 -5304 42662
rect -5338 36654 -5304 36670
rect -5180 42646 -5146 42662
rect -5180 36654 -5146 36670
rect -5022 42646 -4988 42662
rect -5022 36654 -4988 36670
rect -4864 42646 -4830 42662
rect -4864 36654 -4830 36670
rect -4706 42646 -4672 42662
rect -4706 36654 -4672 36670
rect -4548 42646 -4514 42662
rect -4548 36654 -4514 36670
rect -4390 42646 -4356 42662
rect -4390 36654 -4356 36670
rect -4232 42646 -4198 42662
rect -4232 36654 -4198 36670
rect -4074 42646 -4040 42662
rect -4074 36654 -4040 36670
rect -3916 42646 -3882 42662
rect -3916 36654 -3882 36670
rect -3758 42646 -3724 42662
rect -3758 36654 -3724 36670
rect -3600 42646 -3566 42662
rect -3600 36654 -3566 36670
rect -3442 42646 -3408 42662
rect -3442 36654 -3408 36670
rect -3284 42646 -3250 42662
rect -3284 36654 -3250 36670
rect -3126 42646 -3092 42662
rect -3126 36654 -3092 36670
rect -2968 42646 -2934 42662
rect -2968 36654 -2934 36670
rect -2810 42646 -2776 42662
rect -2810 36654 -2776 36670
rect -2652 42646 -2618 42662
rect -2652 36654 -2618 36670
rect -2494 42646 -2460 42662
rect -2494 36654 -2460 36670
rect -2336 42646 -2302 42662
rect -2336 36654 -2302 36670
rect -2178 42646 -2144 42662
rect -2178 36654 -2144 36670
rect -618 42646 -584 42662
rect -618 36654 -584 36670
rect -460 42646 -426 42662
rect -460 36654 -426 36670
rect -302 42646 -268 42662
rect -302 36654 -268 36670
rect -144 42646 -110 42662
rect -144 36654 -110 36670
rect 14 42646 48 42662
rect 14 36654 48 36670
rect 172 42646 206 42662
rect 172 36654 206 36670
rect 330 42646 364 42662
rect 330 36654 364 36670
rect 488 42646 522 42662
rect 488 36654 522 36670
rect 646 42646 680 42662
rect 646 36654 680 36670
rect 804 42646 838 42662
rect 804 36654 838 36670
rect 962 42646 996 42662
rect 962 36654 996 36670
rect 1120 42646 1154 42662
rect 1120 36654 1154 36670
rect 1278 42646 1312 42662
rect 1278 36654 1312 36670
rect 1436 42646 1470 42662
rect 1436 36654 1470 36670
rect 1594 42646 1628 42662
rect 1594 36654 1628 36670
rect 1752 42646 1786 42662
rect 1752 36654 1786 36670
rect 1910 42646 1944 42662
rect 1910 36654 1944 36670
rect 2068 42646 2102 42662
rect 2068 36654 2102 36670
rect 2226 42646 2260 42662
rect 2226 36654 2260 36670
rect 2384 42646 2418 42662
rect 2384 36654 2418 36670
rect 2542 42646 2576 42662
rect 2542 36654 2576 36670
rect 2700 42646 2734 42662
rect 2700 36654 2734 36670
rect 2858 42646 2892 42662
rect 2858 36654 2892 36670
rect 3016 42646 3050 42662
rect 3016 36654 3050 36670
rect 3174 42646 3208 42662
rect 3174 36654 3208 36670
rect 3332 42646 3366 42662
rect 3332 36654 3366 36670
rect 3490 42646 3524 42662
rect 3490 36654 3524 36670
rect 3648 42646 3682 42662
rect 3648 36654 3682 36670
rect 3806 42646 3840 42662
rect 3806 36654 3840 36670
rect 3964 42646 3998 42662
rect 3964 36654 3998 36670
rect 4122 42646 4156 42662
rect 4122 36654 4156 36670
rect 5682 42646 5716 42662
rect 5682 36654 5716 36670
rect 5840 42646 5874 42662
rect 5840 36654 5874 36670
rect 5998 42646 6032 42662
rect 5998 36654 6032 36670
rect 6156 42646 6190 42662
rect 6156 36654 6190 36670
rect 6314 42646 6348 42662
rect 6314 36654 6348 36670
rect 6472 42646 6506 42662
rect 6472 36654 6506 36670
rect 6630 42646 6664 42662
rect 6630 36654 6664 36670
rect 6788 42646 6822 42662
rect 6788 36654 6822 36670
rect 6946 42646 6980 42662
rect 6946 36654 6980 36670
rect 7104 42646 7138 42662
rect 7104 36654 7138 36670
rect 7262 42646 7296 42662
rect 7262 36654 7296 36670
rect 7420 42646 7454 42662
rect 7420 36654 7454 36670
rect 7578 42646 7612 42662
rect 7578 36654 7612 36670
rect 7736 42646 7770 42662
rect 7736 36654 7770 36670
rect 7894 42646 7928 42662
rect 7894 36654 7928 36670
rect 8052 42646 8086 42662
rect 8052 36654 8086 36670
rect 8210 42646 8244 42662
rect 8210 36654 8244 36670
rect 8368 42646 8402 42662
rect 8368 36654 8402 36670
rect 8526 42646 8560 42662
rect 8526 36654 8560 36670
rect 8684 42646 8718 42662
rect 8684 36654 8718 36670
rect 8842 42646 8876 42662
rect 8842 36654 8876 36670
rect 9000 42646 9034 42662
rect 9000 36654 9034 36670
rect 9158 42646 9192 42662
rect 9158 36654 9192 36670
rect 9316 42646 9350 42662
rect 9316 36654 9350 36670
rect 9474 42646 9508 42662
rect 9474 36654 9508 36670
rect 9632 42646 9666 42662
rect 9632 36654 9666 36670
rect 9790 42646 9824 42662
rect 9790 36654 9824 36670
rect 9948 42646 9982 42662
rect 9948 36654 9982 36670
rect 10106 42646 10140 42662
rect 10106 36654 10140 36670
rect 10264 42646 10298 42662
rect 10264 36654 10298 36670
rect 10422 42646 10456 42662
rect 10422 36654 10456 36670
rect -13172 36586 -13156 36620
rect -13088 36586 -13072 36620
rect -13014 36586 -12998 36620
rect -12930 36586 -12914 36620
rect -12856 36586 -12840 36620
rect -12772 36586 -12756 36620
rect -12698 36586 -12682 36620
rect -12614 36586 -12598 36620
rect -12540 36586 -12524 36620
rect -12456 36586 -12440 36620
rect -12382 36586 -12366 36620
rect -12298 36586 -12282 36620
rect -12224 36586 -12208 36620
rect -12140 36586 -12124 36620
rect -12066 36586 -12050 36620
rect -11982 36586 -11966 36620
rect -11908 36586 -11892 36620
rect -11824 36586 -11808 36620
rect -11750 36586 -11734 36620
rect -11666 36586 -11650 36620
rect -11592 36586 -11576 36620
rect -11508 36586 -11492 36620
rect -11434 36586 -11418 36620
rect -11350 36586 -11334 36620
rect -11276 36586 -11260 36620
rect -11192 36586 -11176 36620
rect -11118 36586 -11102 36620
rect -11034 36586 -11018 36620
rect -10960 36586 -10944 36620
rect -10876 36586 -10860 36620
rect -10802 36586 -10786 36620
rect -10718 36586 -10702 36620
rect -10644 36586 -10628 36620
rect -10560 36586 -10544 36620
rect -10486 36586 -10470 36620
rect -10402 36586 -10386 36620
rect -10328 36586 -10312 36620
rect -10244 36586 -10228 36620
rect -10170 36586 -10154 36620
rect -10086 36586 -10070 36620
rect -10012 36586 -9996 36620
rect -9928 36586 -9912 36620
rect -9854 36586 -9838 36620
rect -9770 36586 -9754 36620
rect -9696 36586 -9680 36620
rect -9612 36586 -9596 36620
rect -9538 36586 -9522 36620
rect -9454 36586 -9438 36620
rect -9380 36586 -9364 36620
rect -9296 36586 -9280 36620
rect -9222 36586 -9206 36620
rect -9138 36586 -9122 36620
rect -9064 36586 -9048 36620
rect -8980 36586 -8964 36620
rect -8906 36586 -8890 36620
rect -8822 36586 -8806 36620
rect -8748 36586 -8732 36620
rect -8664 36586 -8648 36620
rect -8590 36586 -8574 36620
rect -8506 36586 -8490 36620
rect -13352 36482 -13318 36544
rect -8344 36482 -8310 36544
rect -13352 36448 -13256 36482
rect -8406 36448 -8310 36482
rect -6872 36586 -6856 36620
rect -6788 36586 -6772 36620
rect -6714 36586 -6698 36620
rect -6630 36586 -6614 36620
rect -6556 36586 -6540 36620
rect -6472 36586 -6456 36620
rect -6398 36586 -6382 36620
rect -6314 36586 -6298 36620
rect -6240 36586 -6224 36620
rect -6156 36586 -6140 36620
rect -6082 36586 -6066 36620
rect -5998 36586 -5982 36620
rect -5924 36586 -5908 36620
rect -5840 36586 -5824 36620
rect -5766 36586 -5750 36620
rect -5682 36586 -5666 36620
rect -5608 36586 -5592 36620
rect -5524 36586 -5508 36620
rect -5450 36586 -5434 36620
rect -5366 36586 -5350 36620
rect -5292 36586 -5276 36620
rect -5208 36586 -5192 36620
rect -5134 36586 -5118 36620
rect -5050 36586 -5034 36620
rect -4976 36586 -4960 36620
rect -4892 36586 -4876 36620
rect -4818 36586 -4802 36620
rect -4734 36586 -4718 36620
rect -4660 36586 -4644 36620
rect -4576 36586 -4560 36620
rect -4502 36586 -4486 36620
rect -4418 36586 -4402 36620
rect -4344 36586 -4328 36620
rect -4260 36586 -4244 36620
rect -4186 36586 -4170 36620
rect -4102 36586 -4086 36620
rect -4028 36586 -4012 36620
rect -3944 36586 -3928 36620
rect -3870 36586 -3854 36620
rect -3786 36586 -3770 36620
rect -3712 36586 -3696 36620
rect -3628 36586 -3612 36620
rect -3554 36586 -3538 36620
rect -3470 36586 -3454 36620
rect -3396 36586 -3380 36620
rect -3312 36586 -3296 36620
rect -3238 36586 -3222 36620
rect -3154 36586 -3138 36620
rect -3080 36586 -3064 36620
rect -2996 36586 -2980 36620
rect -2922 36586 -2906 36620
rect -2838 36586 -2822 36620
rect -2764 36586 -2748 36620
rect -2680 36586 -2664 36620
rect -2606 36586 -2590 36620
rect -2522 36586 -2506 36620
rect -2448 36586 -2432 36620
rect -2364 36586 -2348 36620
rect -2290 36586 -2274 36620
rect -2206 36586 -2190 36620
rect -7052 36482 -7018 36544
rect -2044 36482 -2010 36544
rect -7052 36448 -6956 36482
rect -2106 36448 -2010 36482
rect -572 36586 -556 36620
rect -488 36586 -472 36620
rect -414 36586 -398 36620
rect -330 36586 -314 36620
rect -256 36586 -240 36620
rect -172 36586 -156 36620
rect -98 36586 -82 36620
rect -14 36586 2 36620
rect 60 36586 76 36620
rect 144 36586 160 36620
rect 218 36586 234 36620
rect 302 36586 318 36620
rect 376 36586 392 36620
rect 460 36586 476 36620
rect 534 36586 550 36620
rect 618 36586 634 36620
rect 692 36586 708 36620
rect 776 36586 792 36620
rect 850 36586 866 36620
rect 934 36586 950 36620
rect 1008 36586 1024 36620
rect 1092 36586 1108 36620
rect 1166 36586 1182 36620
rect 1250 36586 1266 36620
rect 1324 36586 1340 36620
rect 1408 36586 1424 36620
rect 1482 36586 1498 36620
rect 1566 36586 1582 36620
rect 1640 36586 1656 36620
rect 1724 36586 1740 36620
rect 1798 36586 1814 36620
rect 1882 36586 1898 36620
rect 1956 36586 1972 36620
rect 2040 36586 2056 36620
rect 2114 36586 2130 36620
rect 2198 36586 2214 36620
rect 2272 36586 2288 36620
rect 2356 36586 2372 36620
rect 2430 36586 2446 36620
rect 2514 36586 2530 36620
rect 2588 36586 2604 36620
rect 2672 36586 2688 36620
rect 2746 36586 2762 36620
rect 2830 36586 2846 36620
rect 2904 36586 2920 36620
rect 2988 36586 3004 36620
rect 3062 36586 3078 36620
rect 3146 36586 3162 36620
rect 3220 36586 3236 36620
rect 3304 36586 3320 36620
rect 3378 36586 3394 36620
rect 3462 36586 3478 36620
rect 3536 36586 3552 36620
rect 3620 36586 3636 36620
rect 3694 36586 3710 36620
rect 3778 36586 3794 36620
rect 3852 36586 3868 36620
rect 3936 36586 3952 36620
rect 4010 36586 4026 36620
rect 4094 36586 4110 36620
rect -752 36482 -718 36544
rect 4256 36482 4290 36544
rect -752 36448 -656 36482
rect 4194 36448 4290 36482
rect 5728 36586 5744 36620
rect 5812 36586 5828 36620
rect 5886 36586 5902 36620
rect 5970 36586 5986 36620
rect 6044 36586 6060 36620
rect 6128 36586 6144 36620
rect 6202 36586 6218 36620
rect 6286 36586 6302 36620
rect 6360 36586 6376 36620
rect 6444 36586 6460 36620
rect 6518 36586 6534 36620
rect 6602 36586 6618 36620
rect 6676 36586 6692 36620
rect 6760 36586 6776 36620
rect 6834 36586 6850 36620
rect 6918 36586 6934 36620
rect 6992 36586 7008 36620
rect 7076 36586 7092 36620
rect 7150 36586 7166 36620
rect 7234 36586 7250 36620
rect 7308 36586 7324 36620
rect 7392 36586 7408 36620
rect 7466 36586 7482 36620
rect 7550 36586 7566 36620
rect 7624 36586 7640 36620
rect 7708 36586 7724 36620
rect 7782 36586 7798 36620
rect 7866 36586 7882 36620
rect 7940 36586 7956 36620
rect 8024 36586 8040 36620
rect 8098 36586 8114 36620
rect 8182 36586 8198 36620
rect 8256 36586 8272 36620
rect 8340 36586 8356 36620
rect 8414 36586 8430 36620
rect 8498 36586 8514 36620
rect 8572 36586 8588 36620
rect 8656 36586 8672 36620
rect 8730 36586 8746 36620
rect 8814 36586 8830 36620
rect 8888 36586 8904 36620
rect 8972 36586 8988 36620
rect 9046 36586 9062 36620
rect 9130 36586 9146 36620
rect 9204 36586 9220 36620
rect 9288 36586 9304 36620
rect 9362 36586 9378 36620
rect 9446 36586 9462 36620
rect 9520 36586 9536 36620
rect 9604 36586 9620 36620
rect 9678 36586 9694 36620
rect 9762 36586 9778 36620
rect 9836 36586 9852 36620
rect 9920 36586 9936 36620
rect 9994 36586 10010 36620
rect 10078 36586 10094 36620
rect 10152 36586 10168 36620
rect 10236 36586 10252 36620
rect 10310 36586 10326 36620
rect 10394 36586 10410 36620
rect 5548 36482 5582 36544
rect 10556 36482 10590 36544
rect 5548 36448 5644 36482
rect 10494 36448 10590 36482
rect -13352 34534 -13256 34568
rect -8406 34534 -8310 34568
rect -13352 34472 -13318 34534
rect -8344 34472 -8310 34534
rect -13172 34396 -13156 34430
rect -13088 34396 -13072 34430
rect -13014 34396 -12998 34430
rect -12930 34396 -12914 34430
rect -12856 34396 -12840 34430
rect -12772 34396 -12756 34430
rect -12698 34396 -12682 34430
rect -12614 34396 -12598 34430
rect -12540 34396 -12524 34430
rect -12456 34396 -12440 34430
rect -12382 34396 -12366 34430
rect -12298 34396 -12282 34430
rect -12224 34396 -12208 34430
rect -12140 34396 -12124 34430
rect -12066 34396 -12050 34430
rect -11982 34396 -11966 34430
rect -11908 34396 -11892 34430
rect -11824 34396 -11808 34430
rect -11750 34396 -11734 34430
rect -11666 34396 -11650 34430
rect -11592 34396 -11576 34430
rect -11508 34396 -11492 34430
rect -11434 34396 -11418 34430
rect -11350 34396 -11334 34430
rect -11276 34396 -11260 34430
rect -11192 34396 -11176 34430
rect -11118 34396 -11102 34430
rect -11034 34396 -11018 34430
rect -10960 34396 -10944 34430
rect -10876 34396 -10860 34430
rect -10802 34396 -10786 34430
rect -10718 34396 -10702 34430
rect -10644 34396 -10628 34430
rect -10560 34396 -10544 34430
rect -10486 34396 -10470 34430
rect -10402 34396 -10386 34430
rect -10328 34396 -10312 34430
rect -10244 34396 -10228 34430
rect -10170 34396 -10154 34430
rect -10086 34396 -10070 34430
rect -10012 34396 -9996 34430
rect -9928 34396 -9912 34430
rect -9854 34396 -9838 34430
rect -9770 34396 -9754 34430
rect -9696 34396 -9680 34430
rect -9612 34396 -9596 34430
rect -9538 34396 -9522 34430
rect -9454 34396 -9438 34430
rect -9380 34396 -9364 34430
rect -9296 34396 -9280 34430
rect -9222 34396 -9206 34430
rect -9138 34396 -9122 34430
rect -9064 34396 -9048 34430
rect -8980 34396 -8964 34430
rect -8906 34396 -8890 34430
rect -8822 34396 -8806 34430
rect -8748 34396 -8732 34430
rect -8664 34396 -8648 34430
rect -8590 34396 -8574 34430
rect -8506 34396 -8490 34430
rect -7052 34534 -6956 34568
rect -2106 34534 -2010 34568
rect -7052 34472 -7018 34534
rect -2044 34472 -2010 34534
rect -6872 34396 -6856 34430
rect -6788 34396 -6772 34430
rect -6714 34396 -6698 34430
rect -6630 34396 -6614 34430
rect -6556 34396 -6540 34430
rect -6472 34396 -6456 34430
rect -6398 34396 -6382 34430
rect -6314 34396 -6298 34430
rect -6240 34396 -6224 34430
rect -6156 34396 -6140 34430
rect -6082 34396 -6066 34430
rect -5998 34396 -5982 34430
rect -5924 34396 -5908 34430
rect -5840 34396 -5824 34430
rect -5766 34396 -5750 34430
rect -5682 34396 -5666 34430
rect -5608 34396 -5592 34430
rect -5524 34396 -5508 34430
rect -5450 34396 -5434 34430
rect -5366 34396 -5350 34430
rect -5292 34396 -5276 34430
rect -5208 34396 -5192 34430
rect -5134 34396 -5118 34430
rect -5050 34396 -5034 34430
rect -4976 34396 -4960 34430
rect -4892 34396 -4876 34430
rect -4818 34396 -4802 34430
rect -4734 34396 -4718 34430
rect -4660 34396 -4644 34430
rect -4576 34396 -4560 34430
rect -4502 34396 -4486 34430
rect -4418 34396 -4402 34430
rect -4344 34396 -4328 34430
rect -4260 34396 -4244 34430
rect -4186 34396 -4170 34430
rect -4102 34396 -4086 34430
rect -4028 34396 -4012 34430
rect -3944 34396 -3928 34430
rect -3870 34396 -3854 34430
rect -3786 34396 -3770 34430
rect -3712 34396 -3696 34430
rect -3628 34396 -3612 34430
rect -3554 34396 -3538 34430
rect -3470 34396 -3454 34430
rect -3396 34396 -3380 34430
rect -3312 34396 -3296 34430
rect -3238 34396 -3222 34430
rect -3154 34396 -3138 34430
rect -3080 34396 -3064 34430
rect -2996 34396 -2980 34430
rect -2922 34396 -2906 34430
rect -2838 34396 -2822 34430
rect -2764 34396 -2748 34430
rect -2680 34396 -2664 34430
rect -2606 34396 -2590 34430
rect -2522 34396 -2506 34430
rect -2448 34396 -2432 34430
rect -2364 34396 -2348 34430
rect -2290 34396 -2274 34430
rect -2206 34396 -2190 34430
rect -752 34534 -656 34568
rect 4194 34534 4290 34568
rect -752 34472 -718 34534
rect 4256 34472 4290 34534
rect -572 34396 -556 34430
rect -488 34396 -472 34430
rect -414 34396 -398 34430
rect -330 34396 -314 34430
rect -256 34396 -240 34430
rect -172 34396 -156 34430
rect -98 34396 -82 34430
rect -14 34396 2 34430
rect 60 34396 76 34430
rect 144 34396 160 34430
rect 218 34396 234 34430
rect 302 34396 318 34430
rect 376 34396 392 34430
rect 460 34396 476 34430
rect 534 34396 550 34430
rect 618 34396 634 34430
rect 692 34396 708 34430
rect 776 34396 792 34430
rect 850 34396 866 34430
rect 934 34396 950 34430
rect 1008 34396 1024 34430
rect 1092 34396 1108 34430
rect 1166 34396 1182 34430
rect 1250 34396 1266 34430
rect 1324 34396 1340 34430
rect 1408 34396 1424 34430
rect 1482 34396 1498 34430
rect 1566 34396 1582 34430
rect 1640 34396 1656 34430
rect 1724 34396 1740 34430
rect 1798 34396 1814 34430
rect 1882 34396 1898 34430
rect 1956 34396 1972 34430
rect 2040 34396 2056 34430
rect 2114 34396 2130 34430
rect 2198 34396 2214 34430
rect 2272 34396 2288 34430
rect 2356 34396 2372 34430
rect 2430 34396 2446 34430
rect 2514 34396 2530 34430
rect 2588 34396 2604 34430
rect 2672 34396 2688 34430
rect 2746 34396 2762 34430
rect 2830 34396 2846 34430
rect 2904 34396 2920 34430
rect 2988 34396 3004 34430
rect 3062 34396 3078 34430
rect 3146 34396 3162 34430
rect 3220 34396 3236 34430
rect 3304 34396 3320 34430
rect 3378 34396 3394 34430
rect 3462 34396 3478 34430
rect 3536 34396 3552 34430
rect 3620 34396 3636 34430
rect 3694 34396 3710 34430
rect 3778 34396 3794 34430
rect 3852 34396 3868 34430
rect 3936 34396 3952 34430
rect 4010 34396 4026 34430
rect 4094 34396 4110 34430
rect 5548 34534 5644 34568
rect 10494 34534 10590 34568
rect 5548 34472 5582 34534
rect 10556 34472 10590 34534
rect 5728 34396 5744 34430
rect 5812 34396 5828 34430
rect 5886 34396 5902 34430
rect 5970 34396 5986 34430
rect 6044 34396 6060 34430
rect 6128 34396 6144 34430
rect 6202 34396 6218 34430
rect 6286 34396 6302 34430
rect 6360 34396 6376 34430
rect 6444 34396 6460 34430
rect 6518 34396 6534 34430
rect 6602 34396 6618 34430
rect 6676 34396 6692 34430
rect 6760 34396 6776 34430
rect 6834 34396 6850 34430
rect 6918 34396 6934 34430
rect 6992 34396 7008 34430
rect 7076 34396 7092 34430
rect 7150 34396 7166 34430
rect 7234 34396 7250 34430
rect 7308 34396 7324 34430
rect 7392 34396 7408 34430
rect 7466 34396 7482 34430
rect 7550 34396 7566 34430
rect 7624 34396 7640 34430
rect 7708 34396 7724 34430
rect 7782 34396 7798 34430
rect 7866 34396 7882 34430
rect 7940 34396 7956 34430
rect 8024 34396 8040 34430
rect 8098 34396 8114 34430
rect 8182 34396 8198 34430
rect 8256 34396 8272 34430
rect 8340 34396 8356 34430
rect 8414 34396 8430 34430
rect 8498 34396 8514 34430
rect 8572 34396 8588 34430
rect 8656 34396 8672 34430
rect 8730 34396 8746 34430
rect 8814 34396 8830 34430
rect 8888 34396 8904 34430
rect 8972 34396 8988 34430
rect 9046 34396 9062 34430
rect 9130 34396 9146 34430
rect 9204 34396 9220 34430
rect 9288 34396 9304 34430
rect 9362 34396 9378 34430
rect 9446 34396 9462 34430
rect 9520 34396 9536 34430
rect 9604 34396 9620 34430
rect 9678 34396 9694 34430
rect 9762 34396 9778 34430
rect 9836 34396 9852 34430
rect 9920 34396 9936 34430
rect 9994 34396 10010 34430
rect 10078 34396 10094 34430
rect 10152 34396 10168 34430
rect 10236 34396 10252 34430
rect 10310 34396 10326 34430
rect 10394 34396 10410 34430
rect -13218 34346 -13184 34362
rect -13218 28354 -13184 28370
rect -13060 34346 -13026 34362
rect -13060 28354 -13026 28370
rect -12902 34346 -12868 34362
rect -12902 28354 -12868 28370
rect -12744 34346 -12710 34362
rect -12744 28354 -12710 28370
rect -12586 34346 -12552 34362
rect -12586 28354 -12552 28370
rect -12428 34346 -12394 34362
rect -12428 28354 -12394 28370
rect -12270 34346 -12236 34362
rect -12270 28354 -12236 28370
rect -12112 34346 -12078 34362
rect -12112 28354 -12078 28370
rect -11954 34346 -11920 34362
rect -11954 28354 -11920 28370
rect -11796 34346 -11762 34362
rect -11796 28354 -11762 28370
rect -11638 34346 -11604 34362
rect -11638 28354 -11604 28370
rect -11480 34346 -11446 34362
rect -11480 28354 -11446 28370
rect -11322 34346 -11288 34362
rect -11322 28354 -11288 28370
rect -11164 34346 -11130 34362
rect -11164 28354 -11130 28370
rect -11006 34346 -10972 34362
rect -11006 28354 -10972 28370
rect -10848 34346 -10814 34362
rect -10848 28354 -10814 28370
rect -10690 34346 -10656 34362
rect -10690 28354 -10656 28370
rect -10532 34346 -10498 34362
rect -10532 28354 -10498 28370
rect -10374 34346 -10340 34362
rect -10374 28354 -10340 28370
rect -10216 34346 -10182 34362
rect -10216 28354 -10182 28370
rect -10058 34346 -10024 34362
rect -10058 28354 -10024 28370
rect -9900 34346 -9866 34362
rect -9900 28354 -9866 28370
rect -9742 34346 -9708 34362
rect -9742 28354 -9708 28370
rect -9584 34346 -9550 34362
rect -9584 28354 -9550 28370
rect -9426 34346 -9392 34362
rect -9426 28354 -9392 28370
rect -9268 34346 -9234 34362
rect -9268 28354 -9234 28370
rect -9110 34346 -9076 34362
rect -9110 28354 -9076 28370
rect -8952 34346 -8918 34362
rect -8952 28354 -8918 28370
rect -8794 34346 -8760 34362
rect -8794 28354 -8760 28370
rect -8636 34346 -8602 34362
rect -8636 28354 -8602 28370
rect -8478 34346 -8444 34362
rect -8478 28354 -8444 28370
rect -6918 34346 -6884 34362
rect -6918 28354 -6884 28370
rect -6760 34346 -6726 34362
rect -6760 28354 -6726 28370
rect -6602 34346 -6568 34362
rect -6602 28354 -6568 28370
rect -6444 34346 -6410 34362
rect -6444 28354 -6410 28370
rect -6286 34346 -6252 34362
rect -6286 28354 -6252 28370
rect -6128 34346 -6094 34362
rect -6128 28354 -6094 28370
rect -5970 34346 -5936 34362
rect -5970 28354 -5936 28370
rect -5812 34346 -5778 34362
rect -5812 28354 -5778 28370
rect -5654 34346 -5620 34362
rect -5654 28354 -5620 28370
rect -5496 34346 -5462 34362
rect -5496 28354 -5462 28370
rect -5338 34346 -5304 34362
rect -5338 28354 -5304 28370
rect -5180 34346 -5146 34362
rect -5180 28354 -5146 28370
rect -5022 34346 -4988 34362
rect -5022 28354 -4988 28370
rect -4864 34346 -4830 34362
rect -4864 28354 -4830 28370
rect -4706 34346 -4672 34362
rect -4706 28354 -4672 28370
rect -4548 34346 -4514 34362
rect -4548 28354 -4514 28370
rect -4390 34346 -4356 34362
rect -4390 28354 -4356 28370
rect -4232 34346 -4198 34362
rect -4232 28354 -4198 28370
rect -4074 34346 -4040 34362
rect -4074 28354 -4040 28370
rect -3916 34346 -3882 34362
rect -3916 28354 -3882 28370
rect -3758 34346 -3724 34362
rect -3758 28354 -3724 28370
rect -3600 34346 -3566 34362
rect -3600 28354 -3566 28370
rect -3442 34346 -3408 34362
rect -3442 28354 -3408 28370
rect -3284 34346 -3250 34362
rect -3284 28354 -3250 28370
rect -3126 34346 -3092 34362
rect -3126 28354 -3092 28370
rect -2968 34346 -2934 34362
rect -2968 28354 -2934 28370
rect -2810 34346 -2776 34362
rect -2810 28354 -2776 28370
rect -2652 34346 -2618 34362
rect -2652 28354 -2618 28370
rect -2494 34346 -2460 34362
rect -2494 28354 -2460 28370
rect -2336 34346 -2302 34362
rect -2336 28354 -2302 28370
rect -2178 34346 -2144 34362
rect -2178 28354 -2144 28370
rect -618 34346 -584 34362
rect -618 28354 -584 28370
rect -460 34346 -426 34362
rect -460 28354 -426 28370
rect -302 34346 -268 34362
rect -302 28354 -268 28370
rect -144 34346 -110 34362
rect -144 28354 -110 28370
rect 14 34346 48 34362
rect 14 28354 48 28370
rect 172 34346 206 34362
rect 172 28354 206 28370
rect 330 34346 364 34362
rect 330 28354 364 28370
rect 488 34346 522 34362
rect 488 28354 522 28370
rect 646 34346 680 34362
rect 646 28354 680 28370
rect 804 34346 838 34362
rect 804 28354 838 28370
rect 962 34346 996 34362
rect 962 28354 996 28370
rect 1120 34346 1154 34362
rect 1120 28354 1154 28370
rect 1278 34346 1312 34362
rect 1278 28354 1312 28370
rect 1436 34346 1470 34362
rect 1436 28354 1470 28370
rect 1594 34346 1628 34362
rect 1594 28354 1628 28370
rect 1752 34346 1786 34362
rect 1752 28354 1786 28370
rect 1910 34346 1944 34362
rect 1910 28354 1944 28370
rect 2068 34346 2102 34362
rect 2068 28354 2102 28370
rect 2226 34346 2260 34362
rect 2226 28354 2260 28370
rect 2384 34346 2418 34362
rect 2384 28354 2418 28370
rect 2542 34346 2576 34362
rect 2542 28354 2576 28370
rect 2700 34346 2734 34362
rect 2700 28354 2734 28370
rect 2858 34346 2892 34362
rect 2858 28354 2892 28370
rect 3016 34346 3050 34362
rect 3016 28354 3050 28370
rect 3174 34346 3208 34362
rect 3174 28354 3208 28370
rect 3332 34346 3366 34362
rect 3332 28354 3366 28370
rect 3490 34346 3524 34362
rect 3490 28354 3524 28370
rect 3648 34346 3682 34362
rect 3648 28354 3682 28370
rect 3806 34346 3840 34362
rect 3806 28354 3840 28370
rect 3964 34346 3998 34362
rect 3964 28354 3998 28370
rect 4122 34346 4156 34362
rect 4122 28354 4156 28370
rect 5682 34346 5716 34362
rect 5682 28354 5716 28370
rect 5840 34346 5874 34362
rect 5840 28354 5874 28370
rect 5998 34346 6032 34362
rect 5998 28354 6032 28370
rect 6156 34346 6190 34362
rect 6156 28354 6190 28370
rect 6314 34346 6348 34362
rect 6314 28354 6348 28370
rect 6472 34346 6506 34362
rect 6472 28354 6506 28370
rect 6630 34346 6664 34362
rect 6630 28354 6664 28370
rect 6788 34346 6822 34362
rect 6788 28354 6822 28370
rect 6946 34346 6980 34362
rect 6946 28354 6980 28370
rect 7104 34346 7138 34362
rect 7104 28354 7138 28370
rect 7262 34346 7296 34362
rect 7262 28354 7296 28370
rect 7420 34346 7454 34362
rect 7420 28354 7454 28370
rect 7578 34346 7612 34362
rect 7578 28354 7612 28370
rect 7736 34346 7770 34362
rect 7736 28354 7770 28370
rect 7894 34346 7928 34362
rect 7894 28354 7928 28370
rect 8052 34346 8086 34362
rect 8052 28354 8086 28370
rect 8210 34346 8244 34362
rect 8210 28354 8244 28370
rect 8368 34346 8402 34362
rect 8368 28354 8402 28370
rect 8526 34346 8560 34362
rect 8526 28354 8560 28370
rect 8684 34346 8718 34362
rect 8684 28354 8718 28370
rect 8842 34346 8876 34362
rect 8842 28354 8876 28370
rect 9000 34346 9034 34362
rect 9000 28354 9034 28370
rect 9158 34346 9192 34362
rect 9158 28354 9192 28370
rect 9316 34346 9350 34362
rect 9316 28354 9350 28370
rect 9474 34346 9508 34362
rect 9474 28354 9508 28370
rect 9632 34346 9666 34362
rect 9632 28354 9666 28370
rect 9790 34346 9824 34362
rect 9790 28354 9824 28370
rect 9948 34346 9982 34362
rect 9948 28354 9982 28370
rect 10106 34346 10140 34362
rect 10106 28354 10140 28370
rect 10264 34346 10298 34362
rect 10264 28354 10298 28370
rect 10422 34346 10456 34362
rect 10422 28354 10456 28370
rect -13172 28286 -13156 28320
rect -13088 28286 -13072 28320
rect -13014 28286 -12998 28320
rect -12930 28286 -12914 28320
rect -12856 28286 -12840 28320
rect -12772 28286 -12756 28320
rect -12698 28286 -12682 28320
rect -12614 28286 -12598 28320
rect -12540 28286 -12524 28320
rect -12456 28286 -12440 28320
rect -12382 28286 -12366 28320
rect -12298 28286 -12282 28320
rect -12224 28286 -12208 28320
rect -12140 28286 -12124 28320
rect -12066 28286 -12050 28320
rect -11982 28286 -11966 28320
rect -11908 28286 -11892 28320
rect -11824 28286 -11808 28320
rect -11750 28286 -11734 28320
rect -11666 28286 -11650 28320
rect -11592 28286 -11576 28320
rect -11508 28286 -11492 28320
rect -11434 28286 -11418 28320
rect -11350 28286 -11334 28320
rect -11276 28286 -11260 28320
rect -11192 28286 -11176 28320
rect -11118 28286 -11102 28320
rect -11034 28286 -11018 28320
rect -10960 28286 -10944 28320
rect -10876 28286 -10860 28320
rect -10802 28286 -10786 28320
rect -10718 28286 -10702 28320
rect -10644 28286 -10628 28320
rect -10560 28286 -10544 28320
rect -10486 28286 -10470 28320
rect -10402 28286 -10386 28320
rect -10328 28286 -10312 28320
rect -10244 28286 -10228 28320
rect -10170 28286 -10154 28320
rect -10086 28286 -10070 28320
rect -10012 28286 -9996 28320
rect -9928 28286 -9912 28320
rect -9854 28286 -9838 28320
rect -9770 28286 -9754 28320
rect -9696 28286 -9680 28320
rect -9612 28286 -9596 28320
rect -9538 28286 -9522 28320
rect -9454 28286 -9438 28320
rect -9380 28286 -9364 28320
rect -9296 28286 -9280 28320
rect -9222 28286 -9206 28320
rect -9138 28286 -9122 28320
rect -9064 28286 -9048 28320
rect -8980 28286 -8964 28320
rect -8906 28286 -8890 28320
rect -8822 28286 -8806 28320
rect -8748 28286 -8732 28320
rect -8664 28286 -8648 28320
rect -8590 28286 -8574 28320
rect -8506 28286 -8490 28320
rect -13352 28182 -13318 28244
rect -8344 28182 -8310 28244
rect -13352 28148 -13256 28182
rect -8406 28148 -8310 28182
rect -6872 28286 -6856 28320
rect -6788 28286 -6772 28320
rect -6714 28286 -6698 28320
rect -6630 28286 -6614 28320
rect -6556 28286 -6540 28320
rect -6472 28286 -6456 28320
rect -6398 28286 -6382 28320
rect -6314 28286 -6298 28320
rect -6240 28286 -6224 28320
rect -6156 28286 -6140 28320
rect -6082 28286 -6066 28320
rect -5998 28286 -5982 28320
rect -5924 28286 -5908 28320
rect -5840 28286 -5824 28320
rect -5766 28286 -5750 28320
rect -5682 28286 -5666 28320
rect -5608 28286 -5592 28320
rect -5524 28286 -5508 28320
rect -5450 28286 -5434 28320
rect -5366 28286 -5350 28320
rect -5292 28286 -5276 28320
rect -5208 28286 -5192 28320
rect -5134 28286 -5118 28320
rect -5050 28286 -5034 28320
rect -4976 28286 -4960 28320
rect -4892 28286 -4876 28320
rect -4818 28286 -4802 28320
rect -4734 28286 -4718 28320
rect -4660 28286 -4644 28320
rect -4576 28286 -4560 28320
rect -4502 28286 -4486 28320
rect -4418 28286 -4402 28320
rect -4344 28286 -4328 28320
rect -4260 28286 -4244 28320
rect -4186 28286 -4170 28320
rect -4102 28286 -4086 28320
rect -4028 28286 -4012 28320
rect -3944 28286 -3928 28320
rect -3870 28286 -3854 28320
rect -3786 28286 -3770 28320
rect -3712 28286 -3696 28320
rect -3628 28286 -3612 28320
rect -3554 28286 -3538 28320
rect -3470 28286 -3454 28320
rect -3396 28286 -3380 28320
rect -3312 28286 -3296 28320
rect -3238 28286 -3222 28320
rect -3154 28286 -3138 28320
rect -3080 28286 -3064 28320
rect -2996 28286 -2980 28320
rect -2922 28286 -2906 28320
rect -2838 28286 -2822 28320
rect -2764 28286 -2748 28320
rect -2680 28286 -2664 28320
rect -2606 28286 -2590 28320
rect -2522 28286 -2506 28320
rect -2448 28286 -2432 28320
rect -2364 28286 -2348 28320
rect -2290 28286 -2274 28320
rect -2206 28286 -2190 28320
rect -7052 28182 -7018 28244
rect -2044 28182 -2010 28244
rect -7052 28148 -6956 28182
rect -2106 28148 -2010 28182
rect -572 28286 -556 28320
rect -488 28286 -472 28320
rect -414 28286 -398 28320
rect -330 28286 -314 28320
rect -256 28286 -240 28320
rect -172 28286 -156 28320
rect -98 28286 -82 28320
rect -14 28286 2 28320
rect 60 28286 76 28320
rect 144 28286 160 28320
rect 218 28286 234 28320
rect 302 28286 318 28320
rect 376 28286 392 28320
rect 460 28286 476 28320
rect 534 28286 550 28320
rect 618 28286 634 28320
rect 692 28286 708 28320
rect 776 28286 792 28320
rect 850 28286 866 28320
rect 934 28286 950 28320
rect 1008 28286 1024 28320
rect 1092 28286 1108 28320
rect 1166 28286 1182 28320
rect 1250 28286 1266 28320
rect 1324 28286 1340 28320
rect 1408 28286 1424 28320
rect 1482 28286 1498 28320
rect 1566 28286 1582 28320
rect 1640 28286 1656 28320
rect 1724 28286 1740 28320
rect 1798 28286 1814 28320
rect 1882 28286 1898 28320
rect 1956 28286 1972 28320
rect 2040 28286 2056 28320
rect 2114 28286 2130 28320
rect 2198 28286 2214 28320
rect 2272 28286 2288 28320
rect 2356 28286 2372 28320
rect 2430 28286 2446 28320
rect 2514 28286 2530 28320
rect 2588 28286 2604 28320
rect 2672 28286 2688 28320
rect 2746 28286 2762 28320
rect 2830 28286 2846 28320
rect 2904 28286 2920 28320
rect 2988 28286 3004 28320
rect 3062 28286 3078 28320
rect 3146 28286 3162 28320
rect 3220 28286 3236 28320
rect 3304 28286 3320 28320
rect 3378 28286 3394 28320
rect 3462 28286 3478 28320
rect 3536 28286 3552 28320
rect 3620 28286 3636 28320
rect 3694 28286 3710 28320
rect 3778 28286 3794 28320
rect 3852 28286 3868 28320
rect 3936 28286 3952 28320
rect 4010 28286 4026 28320
rect 4094 28286 4110 28320
rect -752 28182 -718 28244
rect 4256 28182 4290 28244
rect -752 28148 -656 28182
rect 4194 28148 4290 28182
rect 5728 28286 5744 28320
rect 5812 28286 5828 28320
rect 5886 28286 5902 28320
rect 5970 28286 5986 28320
rect 6044 28286 6060 28320
rect 6128 28286 6144 28320
rect 6202 28286 6218 28320
rect 6286 28286 6302 28320
rect 6360 28286 6376 28320
rect 6444 28286 6460 28320
rect 6518 28286 6534 28320
rect 6602 28286 6618 28320
rect 6676 28286 6692 28320
rect 6760 28286 6776 28320
rect 6834 28286 6850 28320
rect 6918 28286 6934 28320
rect 6992 28286 7008 28320
rect 7076 28286 7092 28320
rect 7150 28286 7166 28320
rect 7234 28286 7250 28320
rect 7308 28286 7324 28320
rect 7392 28286 7408 28320
rect 7466 28286 7482 28320
rect 7550 28286 7566 28320
rect 7624 28286 7640 28320
rect 7708 28286 7724 28320
rect 7782 28286 7798 28320
rect 7866 28286 7882 28320
rect 7940 28286 7956 28320
rect 8024 28286 8040 28320
rect 8098 28286 8114 28320
rect 8182 28286 8198 28320
rect 8256 28286 8272 28320
rect 8340 28286 8356 28320
rect 8414 28286 8430 28320
rect 8498 28286 8514 28320
rect 8572 28286 8588 28320
rect 8656 28286 8672 28320
rect 8730 28286 8746 28320
rect 8814 28286 8830 28320
rect 8888 28286 8904 28320
rect 8972 28286 8988 28320
rect 9046 28286 9062 28320
rect 9130 28286 9146 28320
rect 9204 28286 9220 28320
rect 9288 28286 9304 28320
rect 9362 28286 9378 28320
rect 9446 28286 9462 28320
rect 9520 28286 9536 28320
rect 9604 28286 9620 28320
rect 9678 28286 9694 28320
rect 9762 28286 9778 28320
rect 9836 28286 9852 28320
rect 9920 28286 9936 28320
rect 9994 28286 10010 28320
rect 10078 28286 10094 28320
rect 10152 28286 10168 28320
rect 10236 28286 10252 28320
rect 10310 28286 10326 28320
rect 10394 28286 10410 28320
rect 5548 28182 5582 28244
rect 10556 28182 10590 28244
rect 5548 28148 5644 28182
rect 10494 28148 10590 28182
rect -13352 27534 -13256 27568
rect -8406 27534 -8310 27568
rect -13352 27472 -13318 27534
rect -8344 27472 -8310 27534
rect -13172 27396 -13156 27430
rect -13088 27396 -13072 27430
rect -13014 27396 -12998 27430
rect -12930 27396 -12914 27430
rect -12856 27396 -12840 27430
rect -12772 27396 -12756 27430
rect -12698 27396 -12682 27430
rect -12614 27396 -12598 27430
rect -12540 27396 -12524 27430
rect -12456 27396 -12440 27430
rect -12382 27396 -12366 27430
rect -12298 27396 -12282 27430
rect -12224 27396 -12208 27430
rect -12140 27396 -12124 27430
rect -12066 27396 -12050 27430
rect -11982 27396 -11966 27430
rect -11908 27396 -11892 27430
rect -11824 27396 -11808 27430
rect -11750 27396 -11734 27430
rect -11666 27396 -11650 27430
rect -11592 27396 -11576 27430
rect -11508 27396 -11492 27430
rect -11434 27396 -11418 27430
rect -11350 27396 -11334 27430
rect -11276 27396 -11260 27430
rect -11192 27396 -11176 27430
rect -11118 27396 -11102 27430
rect -11034 27396 -11018 27430
rect -10960 27396 -10944 27430
rect -10876 27396 -10860 27430
rect -10802 27396 -10786 27430
rect -10718 27396 -10702 27430
rect -10644 27396 -10628 27430
rect -10560 27396 -10544 27430
rect -10486 27396 -10470 27430
rect -10402 27396 -10386 27430
rect -10328 27396 -10312 27430
rect -10244 27396 -10228 27430
rect -10170 27396 -10154 27430
rect -10086 27396 -10070 27430
rect -10012 27396 -9996 27430
rect -9928 27396 -9912 27430
rect -9854 27396 -9838 27430
rect -9770 27396 -9754 27430
rect -9696 27396 -9680 27430
rect -9612 27396 -9596 27430
rect -9538 27396 -9522 27430
rect -9454 27396 -9438 27430
rect -9380 27396 -9364 27430
rect -9296 27396 -9280 27430
rect -9222 27396 -9206 27430
rect -9138 27396 -9122 27430
rect -9064 27396 -9048 27430
rect -8980 27396 -8964 27430
rect -8906 27396 -8890 27430
rect -8822 27396 -8806 27430
rect -8748 27396 -8732 27430
rect -8664 27396 -8648 27430
rect -8590 27396 -8574 27430
rect -8506 27396 -8490 27430
rect -7052 27534 -6956 27568
rect -2106 27534 -2010 27568
rect -7052 27472 -7018 27534
rect -2044 27472 -2010 27534
rect -6872 27396 -6856 27430
rect -6788 27396 -6772 27430
rect -6714 27396 -6698 27430
rect -6630 27396 -6614 27430
rect -6556 27396 -6540 27430
rect -6472 27396 -6456 27430
rect -6398 27396 -6382 27430
rect -6314 27396 -6298 27430
rect -6240 27396 -6224 27430
rect -6156 27396 -6140 27430
rect -6082 27396 -6066 27430
rect -5998 27396 -5982 27430
rect -5924 27396 -5908 27430
rect -5840 27396 -5824 27430
rect -5766 27396 -5750 27430
rect -5682 27396 -5666 27430
rect -5608 27396 -5592 27430
rect -5524 27396 -5508 27430
rect -5450 27396 -5434 27430
rect -5366 27396 -5350 27430
rect -5292 27396 -5276 27430
rect -5208 27396 -5192 27430
rect -5134 27396 -5118 27430
rect -5050 27396 -5034 27430
rect -4976 27396 -4960 27430
rect -4892 27396 -4876 27430
rect -4818 27396 -4802 27430
rect -4734 27396 -4718 27430
rect -4660 27396 -4644 27430
rect -4576 27396 -4560 27430
rect -4502 27396 -4486 27430
rect -4418 27396 -4402 27430
rect -4344 27396 -4328 27430
rect -4260 27396 -4244 27430
rect -4186 27396 -4170 27430
rect -4102 27396 -4086 27430
rect -4028 27396 -4012 27430
rect -3944 27396 -3928 27430
rect -3870 27396 -3854 27430
rect -3786 27396 -3770 27430
rect -3712 27396 -3696 27430
rect -3628 27396 -3612 27430
rect -3554 27396 -3538 27430
rect -3470 27396 -3454 27430
rect -3396 27396 -3380 27430
rect -3312 27396 -3296 27430
rect -3238 27396 -3222 27430
rect -3154 27396 -3138 27430
rect -3080 27396 -3064 27430
rect -2996 27396 -2980 27430
rect -2922 27396 -2906 27430
rect -2838 27396 -2822 27430
rect -2764 27396 -2748 27430
rect -2680 27396 -2664 27430
rect -2606 27396 -2590 27430
rect -2522 27396 -2506 27430
rect -2448 27396 -2432 27430
rect -2364 27396 -2348 27430
rect -2290 27396 -2274 27430
rect -2206 27396 -2190 27430
rect -752 27534 -656 27568
rect 4194 27534 4290 27568
rect -752 27472 -718 27534
rect 4256 27472 4290 27534
rect -572 27396 -556 27430
rect -488 27396 -472 27430
rect -414 27396 -398 27430
rect -330 27396 -314 27430
rect -256 27396 -240 27430
rect -172 27396 -156 27430
rect -98 27396 -82 27430
rect -14 27396 2 27430
rect 60 27396 76 27430
rect 144 27396 160 27430
rect 218 27396 234 27430
rect 302 27396 318 27430
rect 376 27396 392 27430
rect 460 27396 476 27430
rect 534 27396 550 27430
rect 618 27396 634 27430
rect 692 27396 708 27430
rect 776 27396 792 27430
rect 850 27396 866 27430
rect 934 27396 950 27430
rect 1008 27396 1024 27430
rect 1092 27396 1108 27430
rect 1166 27396 1182 27430
rect 1250 27396 1266 27430
rect 1324 27396 1340 27430
rect 1408 27396 1424 27430
rect 1482 27396 1498 27430
rect 1566 27396 1582 27430
rect 1640 27396 1656 27430
rect 1724 27396 1740 27430
rect 1798 27396 1814 27430
rect 1882 27396 1898 27430
rect 1956 27396 1972 27430
rect 2040 27396 2056 27430
rect 2114 27396 2130 27430
rect 2198 27396 2214 27430
rect 2272 27396 2288 27430
rect 2356 27396 2372 27430
rect 2430 27396 2446 27430
rect 2514 27396 2530 27430
rect 2588 27396 2604 27430
rect 2672 27396 2688 27430
rect 2746 27396 2762 27430
rect 2830 27396 2846 27430
rect 2904 27396 2920 27430
rect 2988 27396 3004 27430
rect 3062 27396 3078 27430
rect 3146 27396 3162 27430
rect 3220 27396 3236 27430
rect 3304 27396 3320 27430
rect 3378 27396 3394 27430
rect 3462 27396 3478 27430
rect 3536 27396 3552 27430
rect 3620 27396 3636 27430
rect 3694 27396 3710 27430
rect 3778 27396 3794 27430
rect 3852 27396 3868 27430
rect 3936 27396 3952 27430
rect 4010 27396 4026 27430
rect 4094 27396 4110 27430
rect 5548 27534 5644 27568
rect 10494 27534 10590 27568
rect 5548 27472 5582 27534
rect 10556 27472 10590 27534
rect 5728 27396 5744 27430
rect 5812 27396 5828 27430
rect 5886 27396 5902 27430
rect 5970 27396 5986 27430
rect 6044 27396 6060 27430
rect 6128 27396 6144 27430
rect 6202 27396 6218 27430
rect 6286 27396 6302 27430
rect 6360 27396 6376 27430
rect 6444 27396 6460 27430
rect 6518 27396 6534 27430
rect 6602 27396 6618 27430
rect 6676 27396 6692 27430
rect 6760 27396 6776 27430
rect 6834 27396 6850 27430
rect 6918 27396 6934 27430
rect 6992 27396 7008 27430
rect 7076 27396 7092 27430
rect 7150 27396 7166 27430
rect 7234 27396 7250 27430
rect 7308 27396 7324 27430
rect 7392 27396 7408 27430
rect 7466 27396 7482 27430
rect 7550 27396 7566 27430
rect 7624 27396 7640 27430
rect 7708 27396 7724 27430
rect 7782 27396 7798 27430
rect 7866 27396 7882 27430
rect 7940 27396 7956 27430
rect 8024 27396 8040 27430
rect 8098 27396 8114 27430
rect 8182 27396 8198 27430
rect 8256 27396 8272 27430
rect 8340 27396 8356 27430
rect 8414 27396 8430 27430
rect 8498 27396 8514 27430
rect 8572 27396 8588 27430
rect 8656 27396 8672 27430
rect 8730 27396 8746 27430
rect 8814 27396 8830 27430
rect 8888 27396 8904 27430
rect 8972 27396 8988 27430
rect 9046 27396 9062 27430
rect 9130 27396 9146 27430
rect 9204 27396 9220 27430
rect 9288 27396 9304 27430
rect 9362 27396 9378 27430
rect 9446 27396 9462 27430
rect 9520 27396 9536 27430
rect 9604 27396 9620 27430
rect 9678 27396 9694 27430
rect 9762 27396 9778 27430
rect 9836 27396 9852 27430
rect 9920 27396 9936 27430
rect 9994 27396 10010 27430
rect 10078 27396 10094 27430
rect 10152 27396 10168 27430
rect 10236 27396 10252 27430
rect 10310 27396 10326 27430
rect 10394 27396 10410 27430
rect -13218 27346 -13184 27362
rect -13218 21354 -13184 21370
rect -13060 27346 -13026 27362
rect -13060 21354 -13026 21370
rect -12902 27346 -12868 27362
rect -12902 21354 -12868 21370
rect -12744 27346 -12710 27362
rect -12744 21354 -12710 21370
rect -12586 27346 -12552 27362
rect -12586 21354 -12552 21370
rect -12428 27346 -12394 27362
rect -12428 21354 -12394 21370
rect -12270 27346 -12236 27362
rect -12270 21354 -12236 21370
rect -12112 27346 -12078 27362
rect -12112 21354 -12078 21370
rect -11954 27346 -11920 27362
rect -11954 21354 -11920 21370
rect -11796 27346 -11762 27362
rect -11796 21354 -11762 21370
rect -11638 27346 -11604 27362
rect -11638 21354 -11604 21370
rect -11480 27346 -11446 27362
rect -11480 21354 -11446 21370
rect -11322 27346 -11288 27362
rect -11322 21354 -11288 21370
rect -11164 27346 -11130 27362
rect -11164 21354 -11130 21370
rect -11006 27346 -10972 27362
rect -11006 21354 -10972 21370
rect -10848 27346 -10814 27362
rect -10848 21354 -10814 21370
rect -10690 27346 -10656 27362
rect -10690 21354 -10656 21370
rect -10532 27346 -10498 27362
rect -10532 21354 -10498 21370
rect -10374 27346 -10340 27362
rect -10374 21354 -10340 21370
rect -10216 27346 -10182 27362
rect -10216 21354 -10182 21370
rect -10058 27346 -10024 27362
rect -10058 21354 -10024 21370
rect -9900 27346 -9866 27362
rect -9900 21354 -9866 21370
rect -9742 27346 -9708 27362
rect -9742 21354 -9708 21370
rect -9584 27346 -9550 27362
rect -9584 21354 -9550 21370
rect -9426 27346 -9392 27362
rect -9426 21354 -9392 21370
rect -9268 27346 -9234 27362
rect -9268 21354 -9234 21370
rect -9110 27346 -9076 27362
rect -9110 21354 -9076 21370
rect -8952 27346 -8918 27362
rect -8952 21354 -8918 21370
rect -8794 27346 -8760 27362
rect -8794 21354 -8760 21370
rect -8636 27346 -8602 27362
rect -8636 21354 -8602 21370
rect -8478 27346 -8444 27362
rect -8478 21354 -8444 21370
rect -6918 27346 -6884 27362
rect -6918 21354 -6884 21370
rect -6760 27346 -6726 27362
rect -6760 21354 -6726 21370
rect -6602 27346 -6568 27362
rect -6602 21354 -6568 21370
rect -6444 27346 -6410 27362
rect -6444 21354 -6410 21370
rect -6286 27346 -6252 27362
rect -6286 21354 -6252 21370
rect -6128 27346 -6094 27362
rect -6128 21354 -6094 21370
rect -5970 27346 -5936 27362
rect -5970 21354 -5936 21370
rect -5812 27346 -5778 27362
rect -5812 21354 -5778 21370
rect -5654 27346 -5620 27362
rect -5654 21354 -5620 21370
rect -5496 27346 -5462 27362
rect -5496 21354 -5462 21370
rect -5338 27346 -5304 27362
rect -5338 21354 -5304 21370
rect -5180 27346 -5146 27362
rect -5180 21354 -5146 21370
rect -5022 27346 -4988 27362
rect -5022 21354 -4988 21370
rect -4864 27346 -4830 27362
rect -4864 21354 -4830 21370
rect -4706 27346 -4672 27362
rect -4706 21354 -4672 21370
rect -4548 27346 -4514 27362
rect -4548 21354 -4514 21370
rect -4390 27346 -4356 27362
rect -4390 21354 -4356 21370
rect -4232 27346 -4198 27362
rect -4232 21354 -4198 21370
rect -4074 27346 -4040 27362
rect -4074 21354 -4040 21370
rect -3916 27346 -3882 27362
rect -3916 21354 -3882 21370
rect -3758 27346 -3724 27362
rect -3758 21354 -3724 21370
rect -3600 27346 -3566 27362
rect -3600 21354 -3566 21370
rect -3442 27346 -3408 27362
rect -3442 21354 -3408 21370
rect -3284 27346 -3250 27362
rect -3284 21354 -3250 21370
rect -3126 27346 -3092 27362
rect -3126 21354 -3092 21370
rect -2968 27346 -2934 27362
rect -2968 21354 -2934 21370
rect -2810 27346 -2776 27362
rect -2810 21354 -2776 21370
rect -2652 27346 -2618 27362
rect -2652 21354 -2618 21370
rect -2494 27346 -2460 27362
rect -2494 21354 -2460 21370
rect -2336 27346 -2302 27362
rect -2336 21354 -2302 21370
rect -2178 27346 -2144 27362
rect -2178 21354 -2144 21370
rect -618 27346 -584 27362
rect -618 21354 -584 21370
rect -460 27346 -426 27362
rect -460 21354 -426 21370
rect -302 27346 -268 27362
rect -302 21354 -268 21370
rect -144 27346 -110 27362
rect -144 21354 -110 21370
rect 14 27346 48 27362
rect 14 21354 48 21370
rect 172 27346 206 27362
rect 172 21354 206 21370
rect 330 27346 364 27362
rect 330 21354 364 21370
rect 488 27346 522 27362
rect 488 21354 522 21370
rect 646 27346 680 27362
rect 646 21354 680 21370
rect 804 27346 838 27362
rect 804 21354 838 21370
rect 962 27346 996 27362
rect 962 21354 996 21370
rect 1120 27346 1154 27362
rect 1120 21354 1154 21370
rect 1278 27346 1312 27362
rect 1278 21354 1312 21370
rect 1436 27346 1470 27362
rect 1436 21354 1470 21370
rect 1594 27346 1628 27362
rect 1594 21354 1628 21370
rect 1752 27346 1786 27362
rect 1752 21354 1786 21370
rect 1910 27346 1944 27362
rect 1910 21354 1944 21370
rect 2068 27346 2102 27362
rect 2068 21354 2102 21370
rect 2226 27346 2260 27362
rect 2226 21354 2260 21370
rect 2384 27346 2418 27362
rect 2384 21354 2418 21370
rect 2542 27346 2576 27362
rect 2542 21354 2576 21370
rect 2700 27346 2734 27362
rect 2700 21354 2734 21370
rect 2858 27346 2892 27362
rect 2858 21354 2892 21370
rect 3016 27346 3050 27362
rect 3016 21354 3050 21370
rect 3174 27346 3208 27362
rect 3174 21354 3208 21370
rect 3332 27346 3366 27362
rect 3332 21354 3366 21370
rect 3490 27346 3524 27362
rect 3490 21354 3524 21370
rect 3648 27346 3682 27362
rect 3648 21354 3682 21370
rect 3806 27346 3840 27362
rect 3806 21354 3840 21370
rect 3964 27346 3998 27362
rect 3964 21354 3998 21370
rect 4122 27346 4156 27362
rect 4122 21354 4156 21370
rect 5682 27346 5716 27362
rect 5682 21354 5716 21370
rect 5840 27346 5874 27362
rect 5840 21354 5874 21370
rect 5998 27346 6032 27362
rect 5998 21354 6032 21370
rect 6156 27346 6190 27362
rect 6156 21354 6190 21370
rect 6314 27346 6348 27362
rect 6314 21354 6348 21370
rect 6472 27346 6506 27362
rect 6472 21354 6506 21370
rect 6630 27346 6664 27362
rect 6630 21354 6664 21370
rect 6788 27346 6822 27362
rect 6788 21354 6822 21370
rect 6946 27346 6980 27362
rect 6946 21354 6980 21370
rect 7104 27346 7138 27362
rect 7104 21354 7138 21370
rect 7262 27346 7296 27362
rect 7262 21354 7296 21370
rect 7420 27346 7454 27362
rect 7420 21354 7454 21370
rect 7578 27346 7612 27362
rect 7578 21354 7612 21370
rect 7736 27346 7770 27362
rect 7736 21354 7770 21370
rect 7894 27346 7928 27362
rect 7894 21354 7928 21370
rect 8052 27346 8086 27362
rect 8052 21354 8086 21370
rect 8210 27346 8244 27362
rect 8210 21354 8244 21370
rect 8368 27346 8402 27362
rect 8368 21354 8402 21370
rect 8526 27346 8560 27362
rect 8526 21354 8560 21370
rect 8684 27346 8718 27362
rect 8684 21354 8718 21370
rect 8842 27346 8876 27362
rect 8842 21354 8876 21370
rect 9000 27346 9034 27362
rect 9000 21354 9034 21370
rect 9158 27346 9192 27362
rect 9158 21354 9192 21370
rect 9316 27346 9350 27362
rect 9316 21354 9350 21370
rect 9474 27346 9508 27362
rect 9474 21354 9508 21370
rect 9632 27346 9666 27362
rect 9632 21354 9666 21370
rect 9790 27346 9824 27362
rect 9790 21354 9824 21370
rect 9948 27346 9982 27362
rect 9948 21354 9982 21370
rect 10106 27346 10140 27362
rect 10106 21354 10140 21370
rect 10264 27346 10298 27362
rect 10264 21354 10298 21370
rect 10422 27346 10456 27362
rect 10422 21354 10456 21370
rect -13172 21286 -13156 21320
rect -13088 21286 -13072 21320
rect -13014 21286 -12998 21320
rect -12930 21286 -12914 21320
rect -12856 21286 -12840 21320
rect -12772 21286 -12756 21320
rect -12698 21286 -12682 21320
rect -12614 21286 -12598 21320
rect -12540 21286 -12524 21320
rect -12456 21286 -12440 21320
rect -12382 21286 -12366 21320
rect -12298 21286 -12282 21320
rect -12224 21286 -12208 21320
rect -12140 21286 -12124 21320
rect -12066 21286 -12050 21320
rect -11982 21286 -11966 21320
rect -11908 21286 -11892 21320
rect -11824 21286 -11808 21320
rect -11750 21286 -11734 21320
rect -11666 21286 -11650 21320
rect -11592 21286 -11576 21320
rect -11508 21286 -11492 21320
rect -11434 21286 -11418 21320
rect -11350 21286 -11334 21320
rect -11276 21286 -11260 21320
rect -11192 21286 -11176 21320
rect -11118 21286 -11102 21320
rect -11034 21286 -11018 21320
rect -10960 21286 -10944 21320
rect -10876 21286 -10860 21320
rect -10802 21286 -10786 21320
rect -10718 21286 -10702 21320
rect -10644 21286 -10628 21320
rect -10560 21286 -10544 21320
rect -10486 21286 -10470 21320
rect -10402 21286 -10386 21320
rect -10328 21286 -10312 21320
rect -10244 21286 -10228 21320
rect -10170 21286 -10154 21320
rect -10086 21286 -10070 21320
rect -10012 21286 -9996 21320
rect -9928 21286 -9912 21320
rect -9854 21286 -9838 21320
rect -9770 21286 -9754 21320
rect -9696 21286 -9680 21320
rect -9612 21286 -9596 21320
rect -9538 21286 -9522 21320
rect -9454 21286 -9438 21320
rect -9380 21286 -9364 21320
rect -9296 21286 -9280 21320
rect -9222 21286 -9206 21320
rect -9138 21286 -9122 21320
rect -9064 21286 -9048 21320
rect -8980 21286 -8964 21320
rect -8906 21286 -8890 21320
rect -8822 21286 -8806 21320
rect -8748 21286 -8732 21320
rect -8664 21286 -8648 21320
rect -8590 21286 -8574 21320
rect -8506 21286 -8490 21320
rect -13352 21182 -13318 21244
rect -8344 21182 -8310 21244
rect -13352 21148 -13256 21182
rect -8406 21148 -8310 21182
rect -6872 21286 -6856 21320
rect -6788 21286 -6772 21320
rect -6714 21286 -6698 21320
rect -6630 21286 -6614 21320
rect -6556 21286 -6540 21320
rect -6472 21286 -6456 21320
rect -6398 21286 -6382 21320
rect -6314 21286 -6298 21320
rect -6240 21286 -6224 21320
rect -6156 21286 -6140 21320
rect -6082 21286 -6066 21320
rect -5998 21286 -5982 21320
rect -5924 21286 -5908 21320
rect -5840 21286 -5824 21320
rect -5766 21286 -5750 21320
rect -5682 21286 -5666 21320
rect -5608 21286 -5592 21320
rect -5524 21286 -5508 21320
rect -5450 21286 -5434 21320
rect -5366 21286 -5350 21320
rect -5292 21286 -5276 21320
rect -5208 21286 -5192 21320
rect -5134 21286 -5118 21320
rect -5050 21286 -5034 21320
rect -4976 21286 -4960 21320
rect -4892 21286 -4876 21320
rect -4818 21286 -4802 21320
rect -4734 21286 -4718 21320
rect -4660 21286 -4644 21320
rect -4576 21286 -4560 21320
rect -4502 21286 -4486 21320
rect -4418 21286 -4402 21320
rect -4344 21286 -4328 21320
rect -4260 21286 -4244 21320
rect -4186 21286 -4170 21320
rect -4102 21286 -4086 21320
rect -4028 21286 -4012 21320
rect -3944 21286 -3928 21320
rect -3870 21286 -3854 21320
rect -3786 21286 -3770 21320
rect -3712 21286 -3696 21320
rect -3628 21286 -3612 21320
rect -3554 21286 -3538 21320
rect -3470 21286 -3454 21320
rect -3396 21286 -3380 21320
rect -3312 21286 -3296 21320
rect -3238 21286 -3222 21320
rect -3154 21286 -3138 21320
rect -3080 21286 -3064 21320
rect -2996 21286 -2980 21320
rect -2922 21286 -2906 21320
rect -2838 21286 -2822 21320
rect -2764 21286 -2748 21320
rect -2680 21286 -2664 21320
rect -2606 21286 -2590 21320
rect -2522 21286 -2506 21320
rect -2448 21286 -2432 21320
rect -2364 21286 -2348 21320
rect -2290 21286 -2274 21320
rect -2206 21286 -2190 21320
rect -7052 21182 -7018 21244
rect -2044 21182 -2010 21244
rect -7052 21148 -6956 21182
rect -2106 21148 -2010 21182
rect -572 21286 -556 21320
rect -488 21286 -472 21320
rect -414 21286 -398 21320
rect -330 21286 -314 21320
rect -256 21286 -240 21320
rect -172 21286 -156 21320
rect -98 21286 -82 21320
rect -14 21286 2 21320
rect 60 21286 76 21320
rect 144 21286 160 21320
rect 218 21286 234 21320
rect 302 21286 318 21320
rect 376 21286 392 21320
rect 460 21286 476 21320
rect 534 21286 550 21320
rect 618 21286 634 21320
rect 692 21286 708 21320
rect 776 21286 792 21320
rect 850 21286 866 21320
rect 934 21286 950 21320
rect 1008 21286 1024 21320
rect 1092 21286 1108 21320
rect 1166 21286 1182 21320
rect 1250 21286 1266 21320
rect 1324 21286 1340 21320
rect 1408 21286 1424 21320
rect 1482 21286 1498 21320
rect 1566 21286 1582 21320
rect 1640 21286 1656 21320
rect 1724 21286 1740 21320
rect 1798 21286 1814 21320
rect 1882 21286 1898 21320
rect 1956 21286 1972 21320
rect 2040 21286 2056 21320
rect 2114 21286 2130 21320
rect 2198 21286 2214 21320
rect 2272 21286 2288 21320
rect 2356 21286 2372 21320
rect 2430 21286 2446 21320
rect 2514 21286 2530 21320
rect 2588 21286 2604 21320
rect 2672 21286 2688 21320
rect 2746 21286 2762 21320
rect 2830 21286 2846 21320
rect 2904 21286 2920 21320
rect 2988 21286 3004 21320
rect 3062 21286 3078 21320
rect 3146 21286 3162 21320
rect 3220 21286 3236 21320
rect 3304 21286 3320 21320
rect 3378 21286 3394 21320
rect 3462 21286 3478 21320
rect 3536 21286 3552 21320
rect 3620 21286 3636 21320
rect 3694 21286 3710 21320
rect 3778 21286 3794 21320
rect 3852 21286 3868 21320
rect 3936 21286 3952 21320
rect 4010 21286 4026 21320
rect 4094 21286 4110 21320
rect -752 21182 -718 21244
rect 4256 21182 4290 21244
rect -752 21148 -656 21182
rect 4194 21148 4290 21182
rect 5728 21286 5744 21320
rect 5812 21286 5828 21320
rect 5886 21286 5902 21320
rect 5970 21286 5986 21320
rect 6044 21286 6060 21320
rect 6128 21286 6144 21320
rect 6202 21286 6218 21320
rect 6286 21286 6302 21320
rect 6360 21286 6376 21320
rect 6444 21286 6460 21320
rect 6518 21286 6534 21320
rect 6602 21286 6618 21320
rect 6676 21286 6692 21320
rect 6760 21286 6776 21320
rect 6834 21286 6850 21320
rect 6918 21286 6934 21320
rect 6992 21286 7008 21320
rect 7076 21286 7092 21320
rect 7150 21286 7166 21320
rect 7234 21286 7250 21320
rect 7308 21286 7324 21320
rect 7392 21286 7408 21320
rect 7466 21286 7482 21320
rect 7550 21286 7566 21320
rect 7624 21286 7640 21320
rect 7708 21286 7724 21320
rect 7782 21286 7798 21320
rect 7866 21286 7882 21320
rect 7940 21286 7956 21320
rect 8024 21286 8040 21320
rect 8098 21286 8114 21320
rect 8182 21286 8198 21320
rect 8256 21286 8272 21320
rect 8340 21286 8356 21320
rect 8414 21286 8430 21320
rect 8498 21286 8514 21320
rect 8572 21286 8588 21320
rect 8656 21286 8672 21320
rect 8730 21286 8746 21320
rect 8814 21286 8830 21320
rect 8888 21286 8904 21320
rect 8972 21286 8988 21320
rect 9046 21286 9062 21320
rect 9130 21286 9146 21320
rect 9204 21286 9220 21320
rect 9288 21286 9304 21320
rect 9362 21286 9378 21320
rect 9446 21286 9462 21320
rect 9520 21286 9536 21320
rect 9604 21286 9620 21320
rect 9678 21286 9694 21320
rect 9762 21286 9778 21320
rect 9836 21286 9852 21320
rect 9920 21286 9936 21320
rect 9994 21286 10010 21320
rect 10078 21286 10094 21320
rect 10152 21286 10168 21320
rect 10236 21286 10252 21320
rect 10310 21286 10326 21320
rect 10394 21286 10410 21320
rect 5548 21182 5582 21244
rect 10556 21182 10590 21244
rect 5548 21148 5644 21182
rect 10494 21148 10590 21182
rect -13352 19234 -13256 19268
rect -8406 19234 -8310 19268
rect -13352 19172 -13318 19234
rect -8344 19172 -8310 19234
rect -13172 19096 -13156 19130
rect -13088 19096 -13072 19130
rect -13014 19096 -12998 19130
rect -12930 19096 -12914 19130
rect -12856 19096 -12840 19130
rect -12772 19096 -12756 19130
rect -12698 19096 -12682 19130
rect -12614 19096 -12598 19130
rect -12540 19096 -12524 19130
rect -12456 19096 -12440 19130
rect -12382 19096 -12366 19130
rect -12298 19096 -12282 19130
rect -12224 19096 -12208 19130
rect -12140 19096 -12124 19130
rect -12066 19096 -12050 19130
rect -11982 19096 -11966 19130
rect -11908 19096 -11892 19130
rect -11824 19096 -11808 19130
rect -11750 19096 -11734 19130
rect -11666 19096 -11650 19130
rect -11592 19096 -11576 19130
rect -11508 19096 -11492 19130
rect -11434 19096 -11418 19130
rect -11350 19096 -11334 19130
rect -11276 19096 -11260 19130
rect -11192 19096 -11176 19130
rect -11118 19096 -11102 19130
rect -11034 19096 -11018 19130
rect -10960 19096 -10944 19130
rect -10876 19096 -10860 19130
rect -10802 19096 -10786 19130
rect -10718 19096 -10702 19130
rect -10644 19096 -10628 19130
rect -10560 19096 -10544 19130
rect -10486 19096 -10470 19130
rect -10402 19096 -10386 19130
rect -10328 19096 -10312 19130
rect -10244 19096 -10228 19130
rect -10170 19096 -10154 19130
rect -10086 19096 -10070 19130
rect -10012 19096 -9996 19130
rect -9928 19096 -9912 19130
rect -9854 19096 -9838 19130
rect -9770 19096 -9754 19130
rect -9696 19096 -9680 19130
rect -9612 19096 -9596 19130
rect -9538 19096 -9522 19130
rect -9454 19096 -9438 19130
rect -9380 19096 -9364 19130
rect -9296 19096 -9280 19130
rect -9222 19096 -9206 19130
rect -9138 19096 -9122 19130
rect -9064 19096 -9048 19130
rect -8980 19096 -8964 19130
rect -8906 19096 -8890 19130
rect -8822 19096 -8806 19130
rect -8748 19096 -8732 19130
rect -8664 19096 -8648 19130
rect -8590 19096 -8574 19130
rect -8506 19096 -8490 19130
rect -7052 19234 -6956 19268
rect -2106 19234 -2010 19268
rect -7052 19172 -7018 19234
rect -2044 19172 -2010 19234
rect -6872 19096 -6856 19130
rect -6788 19096 -6772 19130
rect -6714 19096 -6698 19130
rect -6630 19096 -6614 19130
rect -6556 19096 -6540 19130
rect -6472 19096 -6456 19130
rect -6398 19096 -6382 19130
rect -6314 19096 -6298 19130
rect -6240 19096 -6224 19130
rect -6156 19096 -6140 19130
rect -6082 19096 -6066 19130
rect -5998 19096 -5982 19130
rect -5924 19096 -5908 19130
rect -5840 19096 -5824 19130
rect -5766 19096 -5750 19130
rect -5682 19096 -5666 19130
rect -5608 19096 -5592 19130
rect -5524 19096 -5508 19130
rect -5450 19096 -5434 19130
rect -5366 19096 -5350 19130
rect -5292 19096 -5276 19130
rect -5208 19096 -5192 19130
rect -5134 19096 -5118 19130
rect -5050 19096 -5034 19130
rect -4976 19096 -4960 19130
rect -4892 19096 -4876 19130
rect -4818 19096 -4802 19130
rect -4734 19096 -4718 19130
rect -4660 19096 -4644 19130
rect -4576 19096 -4560 19130
rect -4502 19096 -4486 19130
rect -4418 19096 -4402 19130
rect -4344 19096 -4328 19130
rect -4260 19096 -4244 19130
rect -4186 19096 -4170 19130
rect -4102 19096 -4086 19130
rect -4028 19096 -4012 19130
rect -3944 19096 -3928 19130
rect -3870 19096 -3854 19130
rect -3786 19096 -3770 19130
rect -3712 19096 -3696 19130
rect -3628 19096 -3612 19130
rect -3554 19096 -3538 19130
rect -3470 19096 -3454 19130
rect -3396 19096 -3380 19130
rect -3312 19096 -3296 19130
rect -3238 19096 -3222 19130
rect -3154 19096 -3138 19130
rect -3080 19096 -3064 19130
rect -2996 19096 -2980 19130
rect -2922 19096 -2906 19130
rect -2838 19096 -2822 19130
rect -2764 19096 -2748 19130
rect -2680 19096 -2664 19130
rect -2606 19096 -2590 19130
rect -2522 19096 -2506 19130
rect -2448 19096 -2432 19130
rect -2364 19096 -2348 19130
rect -2290 19096 -2274 19130
rect -2206 19096 -2190 19130
rect -752 19234 -656 19268
rect 4194 19234 4290 19268
rect -752 19172 -718 19234
rect 4256 19172 4290 19234
rect -572 19096 -556 19130
rect -488 19096 -472 19130
rect -414 19096 -398 19130
rect -330 19096 -314 19130
rect -256 19096 -240 19130
rect -172 19096 -156 19130
rect -98 19096 -82 19130
rect -14 19096 2 19130
rect 60 19096 76 19130
rect 144 19096 160 19130
rect 218 19096 234 19130
rect 302 19096 318 19130
rect 376 19096 392 19130
rect 460 19096 476 19130
rect 534 19096 550 19130
rect 618 19096 634 19130
rect 692 19096 708 19130
rect 776 19096 792 19130
rect 850 19096 866 19130
rect 934 19096 950 19130
rect 1008 19096 1024 19130
rect 1092 19096 1108 19130
rect 1166 19096 1182 19130
rect 1250 19096 1266 19130
rect 1324 19096 1340 19130
rect 1408 19096 1424 19130
rect 1482 19096 1498 19130
rect 1566 19096 1582 19130
rect 1640 19096 1656 19130
rect 1724 19096 1740 19130
rect 1798 19096 1814 19130
rect 1882 19096 1898 19130
rect 1956 19096 1972 19130
rect 2040 19096 2056 19130
rect 2114 19096 2130 19130
rect 2198 19096 2214 19130
rect 2272 19096 2288 19130
rect 2356 19096 2372 19130
rect 2430 19096 2446 19130
rect 2514 19096 2530 19130
rect 2588 19096 2604 19130
rect 2672 19096 2688 19130
rect 2746 19096 2762 19130
rect 2830 19096 2846 19130
rect 2904 19096 2920 19130
rect 2988 19096 3004 19130
rect 3062 19096 3078 19130
rect 3146 19096 3162 19130
rect 3220 19096 3236 19130
rect 3304 19096 3320 19130
rect 3378 19096 3394 19130
rect 3462 19096 3478 19130
rect 3536 19096 3552 19130
rect 3620 19096 3636 19130
rect 3694 19096 3710 19130
rect 3778 19096 3794 19130
rect 3852 19096 3868 19130
rect 3936 19096 3952 19130
rect 4010 19096 4026 19130
rect 4094 19096 4110 19130
rect 5548 19234 5644 19268
rect 10494 19234 10590 19268
rect 5548 19172 5582 19234
rect 10556 19172 10590 19234
rect 5728 19096 5744 19130
rect 5812 19096 5828 19130
rect 5886 19096 5902 19130
rect 5970 19096 5986 19130
rect 6044 19096 6060 19130
rect 6128 19096 6144 19130
rect 6202 19096 6218 19130
rect 6286 19096 6302 19130
rect 6360 19096 6376 19130
rect 6444 19096 6460 19130
rect 6518 19096 6534 19130
rect 6602 19096 6618 19130
rect 6676 19096 6692 19130
rect 6760 19096 6776 19130
rect 6834 19096 6850 19130
rect 6918 19096 6934 19130
rect 6992 19096 7008 19130
rect 7076 19096 7092 19130
rect 7150 19096 7166 19130
rect 7234 19096 7250 19130
rect 7308 19096 7324 19130
rect 7392 19096 7408 19130
rect 7466 19096 7482 19130
rect 7550 19096 7566 19130
rect 7624 19096 7640 19130
rect 7708 19096 7724 19130
rect 7782 19096 7798 19130
rect 7866 19096 7882 19130
rect 7940 19096 7956 19130
rect 8024 19096 8040 19130
rect 8098 19096 8114 19130
rect 8182 19096 8198 19130
rect 8256 19096 8272 19130
rect 8340 19096 8356 19130
rect 8414 19096 8430 19130
rect 8498 19096 8514 19130
rect 8572 19096 8588 19130
rect 8656 19096 8672 19130
rect 8730 19096 8746 19130
rect 8814 19096 8830 19130
rect 8888 19096 8904 19130
rect 8972 19096 8988 19130
rect 9046 19096 9062 19130
rect 9130 19096 9146 19130
rect 9204 19096 9220 19130
rect 9288 19096 9304 19130
rect 9362 19096 9378 19130
rect 9446 19096 9462 19130
rect 9520 19096 9536 19130
rect 9604 19096 9620 19130
rect 9678 19096 9694 19130
rect 9762 19096 9778 19130
rect 9836 19096 9852 19130
rect 9920 19096 9936 19130
rect 9994 19096 10010 19130
rect 10078 19096 10094 19130
rect 10152 19096 10168 19130
rect 10236 19096 10252 19130
rect 10310 19096 10326 19130
rect 10394 19096 10410 19130
rect -13218 19046 -13184 19062
rect -13218 13054 -13184 13070
rect -13060 19046 -13026 19062
rect -13060 13054 -13026 13070
rect -12902 19046 -12868 19062
rect -12902 13054 -12868 13070
rect -12744 19046 -12710 19062
rect -12744 13054 -12710 13070
rect -12586 19046 -12552 19062
rect -12586 13054 -12552 13070
rect -12428 19046 -12394 19062
rect -12428 13054 -12394 13070
rect -12270 19046 -12236 19062
rect -12270 13054 -12236 13070
rect -12112 19046 -12078 19062
rect -12112 13054 -12078 13070
rect -11954 19046 -11920 19062
rect -11954 13054 -11920 13070
rect -11796 19046 -11762 19062
rect -11796 13054 -11762 13070
rect -11638 19046 -11604 19062
rect -11638 13054 -11604 13070
rect -11480 19046 -11446 19062
rect -11480 13054 -11446 13070
rect -11322 19046 -11288 19062
rect -11322 13054 -11288 13070
rect -11164 19046 -11130 19062
rect -11164 13054 -11130 13070
rect -11006 19046 -10972 19062
rect -11006 13054 -10972 13070
rect -10848 19046 -10814 19062
rect -10848 13054 -10814 13070
rect -10690 19046 -10656 19062
rect -10690 13054 -10656 13070
rect -10532 19046 -10498 19062
rect -10532 13054 -10498 13070
rect -10374 19046 -10340 19062
rect -10374 13054 -10340 13070
rect -10216 19046 -10182 19062
rect -10216 13054 -10182 13070
rect -10058 19046 -10024 19062
rect -10058 13054 -10024 13070
rect -9900 19046 -9866 19062
rect -9900 13054 -9866 13070
rect -9742 19046 -9708 19062
rect -9742 13054 -9708 13070
rect -9584 19046 -9550 19062
rect -9584 13054 -9550 13070
rect -9426 19046 -9392 19062
rect -9426 13054 -9392 13070
rect -9268 19046 -9234 19062
rect -9268 13054 -9234 13070
rect -9110 19046 -9076 19062
rect -9110 13054 -9076 13070
rect -8952 19046 -8918 19062
rect -8952 13054 -8918 13070
rect -8794 19046 -8760 19062
rect -8794 13054 -8760 13070
rect -8636 19046 -8602 19062
rect -8636 13054 -8602 13070
rect -8478 19046 -8444 19062
rect -8478 13054 -8444 13070
rect -6918 19046 -6884 19062
rect -6918 13054 -6884 13070
rect -6760 19046 -6726 19062
rect -6760 13054 -6726 13070
rect -6602 19046 -6568 19062
rect -6602 13054 -6568 13070
rect -6444 19046 -6410 19062
rect -6444 13054 -6410 13070
rect -6286 19046 -6252 19062
rect -6286 13054 -6252 13070
rect -6128 19046 -6094 19062
rect -6128 13054 -6094 13070
rect -5970 19046 -5936 19062
rect -5970 13054 -5936 13070
rect -5812 19046 -5778 19062
rect -5812 13054 -5778 13070
rect -5654 19046 -5620 19062
rect -5654 13054 -5620 13070
rect -5496 19046 -5462 19062
rect -5496 13054 -5462 13070
rect -5338 19046 -5304 19062
rect -5338 13054 -5304 13070
rect -5180 19046 -5146 19062
rect -5180 13054 -5146 13070
rect -5022 19046 -4988 19062
rect -5022 13054 -4988 13070
rect -4864 19046 -4830 19062
rect -4864 13054 -4830 13070
rect -4706 19046 -4672 19062
rect -4706 13054 -4672 13070
rect -4548 19046 -4514 19062
rect -4548 13054 -4514 13070
rect -4390 19046 -4356 19062
rect -4390 13054 -4356 13070
rect -4232 19046 -4198 19062
rect -4232 13054 -4198 13070
rect -4074 19046 -4040 19062
rect -4074 13054 -4040 13070
rect -3916 19046 -3882 19062
rect -3916 13054 -3882 13070
rect -3758 19046 -3724 19062
rect -3758 13054 -3724 13070
rect -3600 19046 -3566 19062
rect -3600 13054 -3566 13070
rect -3442 19046 -3408 19062
rect -3442 13054 -3408 13070
rect -3284 19046 -3250 19062
rect -3284 13054 -3250 13070
rect -3126 19046 -3092 19062
rect -3126 13054 -3092 13070
rect -2968 19046 -2934 19062
rect -2968 13054 -2934 13070
rect -2810 19046 -2776 19062
rect -2810 13054 -2776 13070
rect -2652 19046 -2618 19062
rect -2652 13054 -2618 13070
rect -2494 19046 -2460 19062
rect -2494 13054 -2460 13070
rect -2336 19046 -2302 19062
rect -2336 13054 -2302 13070
rect -2178 19046 -2144 19062
rect -2178 13054 -2144 13070
rect -618 19046 -584 19062
rect -618 13054 -584 13070
rect -460 19046 -426 19062
rect -460 13054 -426 13070
rect -302 19046 -268 19062
rect -302 13054 -268 13070
rect -144 19046 -110 19062
rect -144 13054 -110 13070
rect 14 19046 48 19062
rect 14 13054 48 13070
rect 172 19046 206 19062
rect 172 13054 206 13070
rect 330 19046 364 19062
rect 330 13054 364 13070
rect 488 19046 522 19062
rect 488 13054 522 13070
rect 646 19046 680 19062
rect 646 13054 680 13070
rect 804 19046 838 19062
rect 804 13054 838 13070
rect 962 19046 996 19062
rect 962 13054 996 13070
rect 1120 19046 1154 19062
rect 1120 13054 1154 13070
rect 1278 19046 1312 19062
rect 1278 13054 1312 13070
rect 1436 19046 1470 19062
rect 1436 13054 1470 13070
rect 1594 19046 1628 19062
rect 1594 13054 1628 13070
rect 1752 19046 1786 19062
rect 1752 13054 1786 13070
rect 1910 19046 1944 19062
rect 1910 13054 1944 13070
rect 2068 19046 2102 19062
rect 2068 13054 2102 13070
rect 2226 19046 2260 19062
rect 2226 13054 2260 13070
rect 2384 19046 2418 19062
rect 2384 13054 2418 13070
rect 2542 19046 2576 19062
rect 2542 13054 2576 13070
rect 2700 19046 2734 19062
rect 2700 13054 2734 13070
rect 2858 19046 2892 19062
rect 2858 13054 2892 13070
rect 3016 19046 3050 19062
rect 3016 13054 3050 13070
rect 3174 19046 3208 19062
rect 3174 13054 3208 13070
rect 3332 19046 3366 19062
rect 3332 13054 3366 13070
rect 3490 19046 3524 19062
rect 3490 13054 3524 13070
rect 3648 19046 3682 19062
rect 3648 13054 3682 13070
rect 3806 19046 3840 19062
rect 3806 13054 3840 13070
rect 3964 19046 3998 19062
rect 3964 13054 3998 13070
rect 4122 19046 4156 19062
rect 4122 13054 4156 13070
rect 5682 19046 5716 19062
rect 5682 13054 5716 13070
rect 5840 19046 5874 19062
rect 5840 13054 5874 13070
rect 5998 19046 6032 19062
rect 5998 13054 6032 13070
rect 6156 19046 6190 19062
rect 6156 13054 6190 13070
rect 6314 19046 6348 19062
rect 6314 13054 6348 13070
rect 6472 19046 6506 19062
rect 6472 13054 6506 13070
rect 6630 19046 6664 19062
rect 6630 13054 6664 13070
rect 6788 19046 6822 19062
rect 6788 13054 6822 13070
rect 6946 19046 6980 19062
rect 6946 13054 6980 13070
rect 7104 19046 7138 19062
rect 7104 13054 7138 13070
rect 7262 19046 7296 19062
rect 7262 13054 7296 13070
rect 7420 19046 7454 19062
rect 7420 13054 7454 13070
rect 7578 19046 7612 19062
rect 7578 13054 7612 13070
rect 7736 19046 7770 19062
rect 7736 13054 7770 13070
rect 7894 19046 7928 19062
rect 7894 13054 7928 13070
rect 8052 19046 8086 19062
rect 8052 13054 8086 13070
rect 8210 19046 8244 19062
rect 8210 13054 8244 13070
rect 8368 19046 8402 19062
rect 8368 13054 8402 13070
rect 8526 19046 8560 19062
rect 8526 13054 8560 13070
rect 8684 19046 8718 19062
rect 8684 13054 8718 13070
rect 8842 19046 8876 19062
rect 8842 13054 8876 13070
rect 9000 19046 9034 19062
rect 9000 13054 9034 13070
rect 9158 19046 9192 19062
rect 9158 13054 9192 13070
rect 9316 19046 9350 19062
rect 9316 13054 9350 13070
rect 9474 19046 9508 19062
rect 9474 13054 9508 13070
rect 9632 19046 9666 19062
rect 9632 13054 9666 13070
rect 9790 19046 9824 19062
rect 9790 13054 9824 13070
rect 9948 19046 9982 19062
rect 9948 13054 9982 13070
rect 10106 19046 10140 19062
rect 10106 13054 10140 13070
rect 10264 19046 10298 19062
rect 10264 13054 10298 13070
rect 10422 19046 10456 19062
rect 10422 13054 10456 13070
rect -13172 12986 -13156 13020
rect -13088 12986 -13072 13020
rect -13014 12986 -12998 13020
rect -12930 12986 -12914 13020
rect -12856 12986 -12840 13020
rect -12772 12986 -12756 13020
rect -12698 12986 -12682 13020
rect -12614 12986 -12598 13020
rect -12540 12986 -12524 13020
rect -12456 12986 -12440 13020
rect -12382 12986 -12366 13020
rect -12298 12986 -12282 13020
rect -12224 12986 -12208 13020
rect -12140 12986 -12124 13020
rect -12066 12986 -12050 13020
rect -11982 12986 -11966 13020
rect -11908 12986 -11892 13020
rect -11824 12986 -11808 13020
rect -11750 12986 -11734 13020
rect -11666 12986 -11650 13020
rect -11592 12986 -11576 13020
rect -11508 12986 -11492 13020
rect -11434 12986 -11418 13020
rect -11350 12986 -11334 13020
rect -11276 12986 -11260 13020
rect -11192 12986 -11176 13020
rect -11118 12986 -11102 13020
rect -11034 12986 -11018 13020
rect -10960 12986 -10944 13020
rect -10876 12986 -10860 13020
rect -10802 12986 -10786 13020
rect -10718 12986 -10702 13020
rect -10644 12986 -10628 13020
rect -10560 12986 -10544 13020
rect -10486 12986 -10470 13020
rect -10402 12986 -10386 13020
rect -10328 12986 -10312 13020
rect -10244 12986 -10228 13020
rect -10170 12986 -10154 13020
rect -10086 12986 -10070 13020
rect -10012 12986 -9996 13020
rect -9928 12986 -9912 13020
rect -9854 12986 -9838 13020
rect -9770 12986 -9754 13020
rect -9696 12986 -9680 13020
rect -9612 12986 -9596 13020
rect -9538 12986 -9522 13020
rect -9454 12986 -9438 13020
rect -9380 12986 -9364 13020
rect -9296 12986 -9280 13020
rect -9222 12986 -9206 13020
rect -9138 12986 -9122 13020
rect -9064 12986 -9048 13020
rect -8980 12986 -8964 13020
rect -8906 12986 -8890 13020
rect -8822 12986 -8806 13020
rect -8748 12986 -8732 13020
rect -8664 12986 -8648 13020
rect -8590 12986 -8574 13020
rect -8506 12986 -8490 13020
rect -13352 12882 -13318 12944
rect -8344 12882 -8310 12944
rect -13352 12848 -13256 12882
rect -8406 12848 -8310 12882
rect -6872 12986 -6856 13020
rect -6788 12986 -6772 13020
rect -6714 12986 -6698 13020
rect -6630 12986 -6614 13020
rect -6556 12986 -6540 13020
rect -6472 12986 -6456 13020
rect -6398 12986 -6382 13020
rect -6314 12986 -6298 13020
rect -6240 12986 -6224 13020
rect -6156 12986 -6140 13020
rect -6082 12986 -6066 13020
rect -5998 12986 -5982 13020
rect -5924 12986 -5908 13020
rect -5840 12986 -5824 13020
rect -5766 12986 -5750 13020
rect -5682 12986 -5666 13020
rect -5608 12986 -5592 13020
rect -5524 12986 -5508 13020
rect -5450 12986 -5434 13020
rect -5366 12986 -5350 13020
rect -5292 12986 -5276 13020
rect -5208 12986 -5192 13020
rect -5134 12986 -5118 13020
rect -5050 12986 -5034 13020
rect -4976 12986 -4960 13020
rect -4892 12986 -4876 13020
rect -4818 12986 -4802 13020
rect -4734 12986 -4718 13020
rect -4660 12986 -4644 13020
rect -4576 12986 -4560 13020
rect -4502 12986 -4486 13020
rect -4418 12986 -4402 13020
rect -4344 12986 -4328 13020
rect -4260 12986 -4244 13020
rect -4186 12986 -4170 13020
rect -4102 12986 -4086 13020
rect -4028 12986 -4012 13020
rect -3944 12986 -3928 13020
rect -3870 12986 -3854 13020
rect -3786 12986 -3770 13020
rect -3712 12986 -3696 13020
rect -3628 12986 -3612 13020
rect -3554 12986 -3538 13020
rect -3470 12986 -3454 13020
rect -3396 12986 -3380 13020
rect -3312 12986 -3296 13020
rect -3238 12986 -3222 13020
rect -3154 12986 -3138 13020
rect -3080 12986 -3064 13020
rect -2996 12986 -2980 13020
rect -2922 12986 -2906 13020
rect -2838 12986 -2822 13020
rect -2764 12986 -2748 13020
rect -2680 12986 -2664 13020
rect -2606 12986 -2590 13020
rect -2522 12986 -2506 13020
rect -2448 12986 -2432 13020
rect -2364 12986 -2348 13020
rect -2290 12986 -2274 13020
rect -2206 12986 -2190 13020
rect -7052 12882 -7018 12944
rect -2044 12882 -2010 12944
rect -7052 12848 -6956 12882
rect -2106 12848 -2010 12882
rect -572 12986 -556 13020
rect -488 12986 -472 13020
rect -414 12986 -398 13020
rect -330 12986 -314 13020
rect -256 12986 -240 13020
rect -172 12986 -156 13020
rect -98 12986 -82 13020
rect -14 12986 2 13020
rect 60 12986 76 13020
rect 144 12986 160 13020
rect 218 12986 234 13020
rect 302 12986 318 13020
rect 376 12986 392 13020
rect 460 12986 476 13020
rect 534 12986 550 13020
rect 618 12986 634 13020
rect 692 12986 708 13020
rect 776 12986 792 13020
rect 850 12986 866 13020
rect 934 12986 950 13020
rect 1008 12986 1024 13020
rect 1092 12986 1108 13020
rect 1166 12986 1182 13020
rect 1250 12986 1266 13020
rect 1324 12986 1340 13020
rect 1408 12986 1424 13020
rect 1482 12986 1498 13020
rect 1566 12986 1582 13020
rect 1640 12986 1656 13020
rect 1724 12986 1740 13020
rect 1798 12986 1814 13020
rect 1882 12986 1898 13020
rect 1956 12986 1972 13020
rect 2040 12986 2056 13020
rect 2114 12986 2130 13020
rect 2198 12986 2214 13020
rect 2272 12986 2288 13020
rect 2356 12986 2372 13020
rect 2430 12986 2446 13020
rect 2514 12986 2530 13020
rect 2588 12986 2604 13020
rect 2672 12986 2688 13020
rect 2746 12986 2762 13020
rect 2830 12986 2846 13020
rect 2904 12986 2920 13020
rect 2988 12986 3004 13020
rect 3062 12986 3078 13020
rect 3146 12986 3162 13020
rect 3220 12986 3236 13020
rect 3304 12986 3320 13020
rect 3378 12986 3394 13020
rect 3462 12986 3478 13020
rect 3536 12986 3552 13020
rect 3620 12986 3636 13020
rect 3694 12986 3710 13020
rect 3778 12986 3794 13020
rect 3852 12986 3868 13020
rect 3936 12986 3952 13020
rect 4010 12986 4026 13020
rect 4094 12986 4110 13020
rect -752 12882 -718 12944
rect 4256 12882 4290 12944
rect -752 12848 -656 12882
rect 4194 12848 4290 12882
rect 5728 12986 5744 13020
rect 5812 12986 5828 13020
rect 5886 12986 5902 13020
rect 5970 12986 5986 13020
rect 6044 12986 6060 13020
rect 6128 12986 6144 13020
rect 6202 12986 6218 13020
rect 6286 12986 6302 13020
rect 6360 12986 6376 13020
rect 6444 12986 6460 13020
rect 6518 12986 6534 13020
rect 6602 12986 6618 13020
rect 6676 12986 6692 13020
rect 6760 12986 6776 13020
rect 6834 12986 6850 13020
rect 6918 12986 6934 13020
rect 6992 12986 7008 13020
rect 7076 12986 7092 13020
rect 7150 12986 7166 13020
rect 7234 12986 7250 13020
rect 7308 12986 7324 13020
rect 7392 12986 7408 13020
rect 7466 12986 7482 13020
rect 7550 12986 7566 13020
rect 7624 12986 7640 13020
rect 7708 12986 7724 13020
rect 7782 12986 7798 13020
rect 7866 12986 7882 13020
rect 7940 12986 7956 13020
rect 8024 12986 8040 13020
rect 8098 12986 8114 13020
rect 8182 12986 8198 13020
rect 8256 12986 8272 13020
rect 8340 12986 8356 13020
rect 8414 12986 8430 13020
rect 8498 12986 8514 13020
rect 8572 12986 8588 13020
rect 8656 12986 8672 13020
rect 8730 12986 8746 13020
rect 8814 12986 8830 13020
rect 8888 12986 8904 13020
rect 8972 12986 8988 13020
rect 9046 12986 9062 13020
rect 9130 12986 9146 13020
rect 9204 12986 9220 13020
rect 9288 12986 9304 13020
rect 9362 12986 9378 13020
rect 9446 12986 9462 13020
rect 9520 12986 9536 13020
rect 9604 12986 9620 13020
rect 9678 12986 9694 13020
rect 9762 12986 9778 13020
rect 9836 12986 9852 13020
rect 9920 12986 9936 13020
rect 9994 12986 10010 13020
rect 10078 12986 10094 13020
rect 10152 12986 10168 13020
rect 10236 12986 10252 13020
rect 10310 12986 10326 13020
rect 10394 12986 10410 13020
rect 5548 12882 5582 12944
rect 10556 12882 10590 12944
rect 5548 12848 5644 12882
rect 10494 12848 10590 12882
rect -13352 12234 -13256 12268
rect -8406 12234 -8310 12268
rect -13352 12172 -13318 12234
rect -8344 12172 -8310 12234
rect -13172 12096 -13156 12130
rect -13088 12096 -13072 12130
rect -13014 12096 -12998 12130
rect -12930 12096 -12914 12130
rect -12856 12096 -12840 12130
rect -12772 12096 -12756 12130
rect -12698 12096 -12682 12130
rect -12614 12096 -12598 12130
rect -12540 12096 -12524 12130
rect -12456 12096 -12440 12130
rect -12382 12096 -12366 12130
rect -12298 12096 -12282 12130
rect -12224 12096 -12208 12130
rect -12140 12096 -12124 12130
rect -12066 12096 -12050 12130
rect -11982 12096 -11966 12130
rect -11908 12096 -11892 12130
rect -11824 12096 -11808 12130
rect -11750 12096 -11734 12130
rect -11666 12096 -11650 12130
rect -11592 12096 -11576 12130
rect -11508 12096 -11492 12130
rect -11434 12096 -11418 12130
rect -11350 12096 -11334 12130
rect -11276 12096 -11260 12130
rect -11192 12096 -11176 12130
rect -11118 12096 -11102 12130
rect -11034 12096 -11018 12130
rect -10960 12096 -10944 12130
rect -10876 12096 -10860 12130
rect -10802 12096 -10786 12130
rect -10718 12096 -10702 12130
rect -10644 12096 -10628 12130
rect -10560 12096 -10544 12130
rect -10486 12096 -10470 12130
rect -10402 12096 -10386 12130
rect -10328 12096 -10312 12130
rect -10244 12096 -10228 12130
rect -10170 12096 -10154 12130
rect -10086 12096 -10070 12130
rect -10012 12096 -9996 12130
rect -9928 12096 -9912 12130
rect -9854 12096 -9838 12130
rect -9770 12096 -9754 12130
rect -9696 12096 -9680 12130
rect -9612 12096 -9596 12130
rect -9538 12096 -9522 12130
rect -9454 12096 -9438 12130
rect -9380 12096 -9364 12130
rect -9296 12096 -9280 12130
rect -9222 12096 -9206 12130
rect -9138 12096 -9122 12130
rect -9064 12096 -9048 12130
rect -8980 12096 -8964 12130
rect -8906 12096 -8890 12130
rect -8822 12096 -8806 12130
rect -8748 12096 -8732 12130
rect -8664 12096 -8648 12130
rect -8590 12096 -8574 12130
rect -8506 12096 -8490 12130
rect -7052 12234 -6956 12268
rect -2106 12234 -2010 12268
rect -7052 12172 -7018 12234
rect -2044 12172 -2010 12234
rect -6872 12096 -6856 12130
rect -6788 12096 -6772 12130
rect -6714 12096 -6698 12130
rect -6630 12096 -6614 12130
rect -6556 12096 -6540 12130
rect -6472 12096 -6456 12130
rect -6398 12096 -6382 12130
rect -6314 12096 -6298 12130
rect -6240 12096 -6224 12130
rect -6156 12096 -6140 12130
rect -6082 12096 -6066 12130
rect -5998 12096 -5982 12130
rect -5924 12096 -5908 12130
rect -5840 12096 -5824 12130
rect -5766 12096 -5750 12130
rect -5682 12096 -5666 12130
rect -5608 12096 -5592 12130
rect -5524 12096 -5508 12130
rect -5450 12096 -5434 12130
rect -5366 12096 -5350 12130
rect -5292 12096 -5276 12130
rect -5208 12096 -5192 12130
rect -5134 12096 -5118 12130
rect -5050 12096 -5034 12130
rect -4976 12096 -4960 12130
rect -4892 12096 -4876 12130
rect -4818 12096 -4802 12130
rect -4734 12096 -4718 12130
rect -4660 12096 -4644 12130
rect -4576 12096 -4560 12130
rect -4502 12096 -4486 12130
rect -4418 12096 -4402 12130
rect -4344 12096 -4328 12130
rect -4260 12096 -4244 12130
rect -4186 12096 -4170 12130
rect -4102 12096 -4086 12130
rect -4028 12096 -4012 12130
rect -3944 12096 -3928 12130
rect -3870 12096 -3854 12130
rect -3786 12096 -3770 12130
rect -3712 12096 -3696 12130
rect -3628 12096 -3612 12130
rect -3554 12096 -3538 12130
rect -3470 12096 -3454 12130
rect -3396 12096 -3380 12130
rect -3312 12096 -3296 12130
rect -3238 12096 -3222 12130
rect -3154 12096 -3138 12130
rect -3080 12096 -3064 12130
rect -2996 12096 -2980 12130
rect -2922 12096 -2906 12130
rect -2838 12096 -2822 12130
rect -2764 12096 -2748 12130
rect -2680 12096 -2664 12130
rect -2606 12096 -2590 12130
rect -2522 12096 -2506 12130
rect -2448 12096 -2432 12130
rect -2364 12096 -2348 12130
rect -2290 12096 -2274 12130
rect -2206 12096 -2190 12130
rect -752 12234 -656 12268
rect 4194 12234 4290 12268
rect -752 12172 -718 12234
rect 4256 12172 4290 12234
rect -572 12096 -556 12130
rect -488 12096 -472 12130
rect -414 12096 -398 12130
rect -330 12096 -314 12130
rect -256 12096 -240 12130
rect -172 12096 -156 12130
rect -98 12096 -82 12130
rect -14 12096 2 12130
rect 60 12096 76 12130
rect 144 12096 160 12130
rect 218 12096 234 12130
rect 302 12096 318 12130
rect 376 12096 392 12130
rect 460 12096 476 12130
rect 534 12096 550 12130
rect 618 12096 634 12130
rect 692 12096 708 12130
rect 776 12096 792 12130
rect 850 12096 866 12130
rect 934 12096 950 12130
rect 1008 12096 1024 12130
rect 1092 12096 1108 12130
rect 1166 12096 1182 12130
rect 1250 12096 1266 12130
rect 1324 12096 1340 12130
rect 1408 12096 1424 12130
rect 1482 12096 1498 12130
rect 1566 12096 1582 12130
rect 1640 12096 1656 12130
rect 1724 12096 1740 12130
rect 1798 12096 1814 12130
rect 1882 12096 1898 12130
rect 1956 12096 1972 12130
rect 2040 12096 2056 12130
rect 2114 12096 2130 12130
rect 2198 12096 2214 12130
rect 2272 12096 2288 12130
rect 2356 12096 2372 12130
rect 2430 12096 2446 12130
rect 2514 12096 2530 12130
rect 2588 12096 2604 12130
rect 2672 12096 2688 12130
rect 2746 12096 2762 12130
rect 2830 12096 2846 12130
rect 2904 12096 2920 12130
rect 2988 12096 3004 12130
rect 3062 12096 3078 12130
rect 3146 12096 3162 12130
rect 3220 12096 3236 12130
rect 3304 12096 3320 12130
rect 3378 12096 3394 12130
rect 3462 12096 3478 12130
rect 3536 12096 3552 12130
rect 3620 12096 3636 12130
rect 3694 12096 3710 12130
rect 3778 12096 3794 12130
rect 3852 12096 3868 12130
rect 3936 12096 3952 12130
rect 4010 12096 4026 12130
rect 4094 12096 4110 12130
rect 5548 12234 5644 12268
rect 10494 12234 10590 12268
rect 5548 12172 5582 12234
rect 10556 12172 10590 12234
rect 5728 12096 5744 12130
rect 5812 12096 5828 12130
rect 5886 12096 5902 12130
rect 5970 12096 5986 12130
rect 6044 12096 6060 12130
rect 6128 12096 6144 12130
rect 6202 12096 6218 12130
rect 6286 12096 6302 12130
rect 6360 12096 6376 12130
rect 6444 12096 6460 12130
rect 6518 12096 6534 12130
rect 6602 12096 6618 12130
rect 6676 12096 6692 12130
rect 6760 12096 6776 12130
rect 6834 12096 6850 12130
rect 6918 12096 6934 12130
rect 6992 12096 7008 12130
rect 7076 12096 7092 12130
rect 7150 12096 7166 12130
rect 7234 12096 7250 12130
rect 7308 12096 7324 12130
rect 7392 12096 7408 12130
rect 7466 12096 7482 12130
rect 7550 12096 7566 12130
rect 7624 12096 7640 12130
rect 7708 12096 7724 12130
rect 7782 12096 7798 12130
rect 7866 12096 7882 12130
rect 7940 12096 7956 12130
rect 8024 12096 8040 12130
rect 8098 12096 8114 12130
rect 8182 12096 8198 12130
rect 8256 12096 8272 12130
rect 8340 12096 8356 12130
rect 8414 12096 8430 12130
rect 8498 12096 8514 12130
rect 8572 12096 8588 12130
rect 8656 12096 8672 12130
rect 8730 12096 8746 12130
rect 8814 12096 8830 12130
rect 8888 12096 8904 12130
rect 8972 12096 8988 12130
rect 9046 12096 9062 12130
rect 9130 12096 9146 12130
rect 9204 12096 9220 12130
rect 9288 12096 9304 12130
rect 9362 12096 9378 12130
rect 9446 12096 9462 12130
rect 9520 12096 9536 12130
rect 9604 12096 9620 12130
rect 9678 12096 9694 12130
rect 9762 12096 9778 12130
rect 9836 12096 9852 12130
rect 9920 12096 9936 12130
rect 9994 12096 10010 12130
rect 10078 12096 10094 12130
rect 10152 12096 10168 12130
rect 10236 12096 10252 12130
rect 10310 12096 10326 12130
rect 10394 12096 10410 12130
rect -13218 12046 -13184 12062
rect -13218 6054 -13184 6070
rect -13060 12046 -13026 12062
rect -13060 6054 -13026 6070
rect -12902 12046 -12868 12062
rect -12902 6054 -12868 6070
rect -12744 12046 -12710 12062
rect -12744 6054 -12710 6070
rect -12586 12046 -12552 12062
rect -12586 6054 -12552 6070
rect -12428 12046 -12394 12062
rect -12428 6054 -12394 6070
rect -12270 12046 -12236 12062
rect -12270 6054 -12236 6070
rect -12112 12046 -12078 12062
rect -12112 6054 -12078 6070
rect -11954 12046 -11920 12062
rect -11954 6054 -11920 6070
rect -11796 12046 -11762 12062
rect -11796 6054 -11762 6070
rect -11638 12046 -11604 12062
rect -11638 6054 -11604 6070
rect -11480 12046 -11446 12062
rect -11480 6054 -11446 6070
rect -11322 12046 -11288 12062
rect -11322 6054 -11288 6070
rect -11164 12046 -11130 12062
rect -11164 6054 -11130 6070
rect -11006 12046 -10972 12062
rect -11006 6054 -10972 6070
rect -10848 12046 -10814 12062
rect -10848 6054 -10814 6070
rect -10690 12046 -10656 12062
rect -10690 6054 -10656 6070
rect -10532 12046 -10498 12062
rect -10532 6054 -10498 6070
rect -10374 12046 -10340 12062
rect -10374 6054 -10340 6070
rect -10216 12046 -10182 12062
rect -10216 6054 -10182 6070
rect -10058 12046 -10024 12062
rect -10058 6054 -10024 6070
rect -9900 12046 -9866 12062
rect -9900 6054 -9866 6070
rect -9742 12046 -9708 12062
rect -9742 6054 -9708 6070
rect -9584 12046 -9550 12062
rect -9584 6054 -9550 6070
rect -9426 12046 -9392 12062
rect -9426 6054 -9392 6070
rect -9268 12046 -9234 12062
rect -9268 6054 -9234 6070
rect -9110 12046 -9076 12062
rect -9110 6054 -9076 6070
rect -8952 12046 -8918 12062
rect -8952 6054 -8918 6070
rect -8794 12046 -8760 12062
rect -8794 6054 -8760 6070
rect -8636 12046 -8602 12062
rect -8636 6054 -8602 6070
rect -8478 12046 -8444 12062
rect -8478 6054 -8444 6070
rect -6918 12046 -6884 12062
rect -6918 6054 -6884 6070
rect -6760 12046 -6726 12062
rect -6760 6054 -6726 6070
rect -6602 12046 -6568 12062
rect -6602 6054 -6568 6070
rect -6444 12046 -6410 12062
rect -6444 6054 -6410 6070
rect -6286 12046 -6252 12062
rect -6286 6054 -6252 6070
rect -6128 12046 -6094 12062
rect -6128 6054 -6094 6070
rect -5970 12046 -5936 12062
rect -5970 6054 -5936 6070
rect -5812 12046 -5778 12062
rect -5812 6054 -5778 6070
rect -5654 12046 -5620 12062
rect -5654 6054 -5620 6070
rect -5496 12046 -5462 12062
rect -5496 6054 -5462 6070
rect -5338 12046 -5304 12062
rect -5338 6054 -5304 6070
rect -5180 12046 -5146 12062
rect -5180 6054 -5146 6070
rect -5022 12046 -4988 12062
rect -5022 6054 -4988 6070
rect -4864 12046 -4830 12062
rect -4864 6054 -4830 6070
rect -4706 12046 -4672 12062
rect -4706 6054 -4672 6070
rect -4548 12046 -4514 12062
rect -4548 6054 -4514 6070
rect -4390 12046 -4356 12062
rect -4390 6054 -4356 6070
rect -4232 12046 -4198 12062
rect -4232 6054 -4198 6070
rect -4074 12046 -4040 12062
rect -4074 6054 -4040 6070
rect -3916 12046 -3882 12062
rect -3916 6054 -3882 6070
rect -3758 12046 -3724 12062
rect -3758 6054 -3724 6070
rect -3600 12046 -3566 12062
rect -3600 6054 -3566 6070
rect -3442 12046 -3408 12062
rect -3442 6054 -3408 6070
rect -3284 12046 -3250 12062
rect -3284 6054 -3250 6070
rect -3126 12046 -3092 12062
rect -3126 6054 -3092 6070
rect -2968 12046 -2934 12062
rect -2968 6054 -2934 6070
rect -2810 12046 -2776 12062
rect -2810 6054 -2776 6070
rect -2652 12046 -2618 12062
rect -2652 6054 -2618 6070
rect -2494 12046 -2460 12062
rect -2494 6054 -2460 6070
rect -2336 12046 -2302 12062
rect -2336 6054 -2302 6070
rect -2178 12046 -2144 12062
rect -2178 6054 -2144 6070
rect -618 12046 -584 12062
rect -618 6054 -584 6070
rect -460 12046 -426 12062
rect -460 6054 -426 6070
rect -302 12046 -268 12062
rect -302 6054 -268 6070
rect -144 12046 -110 12062
rect -144 6054 -110 6070
rect 14 12046 48 12062
rect 14 6054 48 6070
rect 172 12046 206 12062
rect 172 6054 206 6070
rect 330 12046 364 12062
rect 330 6054 364 6070
rect 488 12046 522 12062
rect 488 6054 522 6070
rect 646 12046 680 12062
rect 646 6054 680 6070
rect 804 12046 838 12062
rect 804 6054 838 6070
rect 962 12046 996 12062
rect 962 6054 996 6070
rect 1120 12046 1154 12062
rect 1120 6054 1154 6070
rect 1278 12046 1312 12062
rect 1278 6054 1312 6070
rect 1436 12046 1470 12062
rect 1436 6054 1470 6070
rect 1594 12046 1628 12062
rect 1594 6054 1628 6070
rect 1752 12046 1786 12062
rect 1752 6054 1786 6070
rect 1910 12046 1944 12062
rect 1910 6054 1944 6070
rect 2068 12046 2102 12062
rect 2068 6054 2102 6070
rect 2226 12046 2260 12062
rect 2226 6054 2260 6070
rect 2384 12046 2418 12062
rect 2384 6054 2418 6070
rect 2542 12046 2576 12062
rect 2542 6054 2576 6070
rect 2700 12046 2734 12062
rect 2700 6054 2734 6070
rect 2858 12046 2892 12062
rect 2858 6054 2892 6070
rect 3016 12046 3050 12062
rect 3016 6054 3050 6070
rect 3174 12046 3208 12062
rect 3174 6054 3208 6070
rect 3332 12046 3366 12062
rect 3332 6054 3366 6070
rect 3490 12046 3524 12062
rect 3490 6054 3524 6070
rect 3648 12046 3682 12062
rect 3648 6054 3682 6070
rect 3806 12046 3840 12062
rect 3806 6054 3840 6070
rect 3964 12046 3998 12062
rect 3964 6054 3998 6070
rect 4122 12046 4156 12062
rect 4122 6054 4156 6070
rect 5682 12046 5716 12062
rect 5682 6054 5716 6070
rect 5840 12046 5874 12062
rect 5840 6054 5874 6070
rect 5998 12046 6032 12062
rect 5998 6054 6032 6070
rect 6156 12046 6190 12062
rect 6156 6054 6190 6070
rect 6314 12046 6348 12062
rect 6314 6054 6348 6070
rect 6472 12046 6506 12062
rect 6472 6054 6506 6070
rect 6630 12046 6664 12062
rect 6630 6054 6664 6070
rect 6788 12046 6822 12062
rect 6788 6054 6822 6070
rect 6946 12046 6980 12062
rect 6946 6054 6980 6070
rect 7104 12046 7138 12062
rect 7104 6054 7138 6070
rect 7262 12046 7296 12062
rect 7262 6054 7296 6070
rect 7420 12046 7454 12062
rect 7420 6054 7454 6070
rect 7578 12046 7612 12062
rect 7578 6054 7612 6070
rect 7736 12046 7770 12062
rect 7736 6054 7770 6070
rect 7894 12046 7928 12062
rect 7894 6054 7928 6070
rect 8052 12046 8086 12062
rect 8052 6054 8086 6070
rect 8210 12046 8244 12062
rect 8210 6054 8244 6070
rect 8368 12046 8402 12062
rect 8368 6054 8402 6070
rect 8526 12046 8560 12062
rect 8526 6054 8560 6070
rect 8684 12046 8718 12062
rect 8684 6054 8718 6070
rect 8842 12046 8876 12062
rect 8842 6054 8876 6070
rect 9000 12046 9034 12062
rect 9000 6054 9034 6070
rect 9158 12046 9192 12062
rect 9158 6054 9192 6070
rect 9316 12046 9350 12062
rect 9316 6054 9350 6070
rect 9474 12046 9508 12062
rect 9474 6054 9508 6070
rect 9632 12046 9666 12062
rect 9632 6054 9666 6070
rect 9790 12046 9824 12062
rect 9790 6054 9824 6070
rect 9948 12046 9982 12062
rect 9948 6054 9982 6070
rect 10106 12046 10140 12062
rect 10106 6054 10140 6070
rect 10264 12046 10298 12062
rect 10264 6054 10298 6070
rect 10422 12046 10456 12062
rect 10422 6054 10456 6070
rect -13172 5986 -13156 6020
rect -13088 5986 -13072 6020
rect -13014 5986 -12998 6020
rect -12930 5986 -12914 6020
rect -12856 5986 -12840 6020
rect -12772 5986 -12756 6020
rect -12698 5986 -12682 6020
rect -12614 5986 -12598 6020
rect -12540 5986 -12524 6020
rect -12456 5986 -12440 6020
rect -12382 5986 -12366 6020
rect -12298 5986 -12282 6020
rect -12224 5986 -12208 6020
rect -12140 5986 -12124 6020
rect -12066 5986 -12050 6020
rect -11982 5986 -11966 6020
rect -11908 5986 -11892 6020
rect -11824 5986 -11808 6020
rect -11750 5986 -11734 6020
rect -11666 5986 -11650 6020
rect -11592 5986 -11576 6020
rect -11508 5986 -11492 6020
rect -11434 5986 -11418 6020
rect -11350 5986 -11334 6020
rect -11276 5986 -11260 6020
rect -11192 5986 -11176 6020
rect -11118 5986 -11102 6020
rect -11034 5986 -11018 6020
rect -10960 5986 -10944 6020
rect -10876 5986 -10860 6020
rect -10802 5986 -10786 6020
rect -10718 5986 -10702 6020
rect -10644 5986 -10628 6020
rect -10560 5986 -10544 6020
rect -10486 5986 -10470 6020
rect -10402 5986 -10386 6020
rect -10328 5986 -10312 6020
rect -10244 5986 -10228 6020
rect -10170 5986 -10154 6020
rect -10086 5986 -10070 6020
rect -10012 5986 -9996 6020
rect -9928 5986 -9912 6020
rect -9854 5986 -9838 6020
rect -9770 5986 -9754 6020
rect -9696 5986 -9680 6020
rect -9612 5986 -9596 6020
rect -9538 5986 -9522 6020
rect -9454 5986 -9438 6020
rect -9380 5986 -9364 6020
rect -9296 5986 -9280 6020
rect -9222 5986 -9206 6020
rect -9138 5986 -9122 6020
rect -9064 5986 -9048 6020
rect -8980 5986 -8964 6020
rect -8906 5986 -8890 6020
rect -8822 5986 -8806 6020
rect -8748 5986 -8732 6020
rect -8664 5986 -8648 6020
rect -8590 5986 -8574 6020
rect -8506 5986 -8490 6020
rect -13352 5882 -13318 5944
rect -8344 5882 -8310 5944
rect -13352 5848 -13256 5882
rect -8406 5848 -8310 5882
rect -6872 5986 -6856 6020
rect -6788 5986 -6772 6020
rect -6714 5986 -6698 6020
rect -6630 5986 -6614 6020
rect -6556 5986 -6540 6020
rect -6472 5986 -6456 6020
rect -6398 5986 -6382 6020
rect -6314 5986 -6298 6020
rect -6240 5986 -6224 6020
rect -6156 5986 -6140 6020
rect -6082 5986 -6066 6020
rect -5998 5986 -5982 6020
rect -5924 5986 -5908 6020
rect -5840 5986 -5824 6020
rect -5766 5986 -5750 6020
rect -5682 5986 -5666 6020
rect -5608 5986 -5592 6020
rect -5524 5986 -5508 6020
rect -5450 5986 -5434 6020
rect -5366 5986 -5350 6020
rect -5292 5986 -5276 6020
rect -5208 5986 -5192 6020
rect -5134 5986 -5118 6020
rect -5050 5986 -5034 6020
rect -4976 5986 -4960 6020
rect -4892 5986 -4876 6020
rect -4818 5986 -4802 6020
rect -4734 5986 -4718 6020
rect -4660 5986 -4644 6020
rect -4576 5986 -4560 6020
rect -4502 5986 -4486 6020
rect -4418 5986 -4402 6020
rect -4344 5986 -4328 6020
rect -4260 5986 -4244 6020
rect -4186 5986 -4170 6020
rect -4102 5986 -4086 6020
rect -4028 5986 -4012 6020
rect -3944 5986 -3928 6020
rect -3870 5986 -3854 6020
rect -3786 5986 -3770 6020
rect -3712 5986 -3696 6020
rect -3628 5986 -3612 6020
rect -3554 5986 -3538 6020
rect -3470 5986 -3454 6020
rect -3396 5986 -3380 6020
rect -3312 5986 -3296 6020
rect -3238 5986 -3222 6020
rect -3154 5986 -3138 6020
rect -3080 5986 -3064 6020
rect -2996 5986 -2980 6020
rect -2922 5986 -2906 6020
rect -2838 5986 -2822 6020
rect -2764 5986 -2748 6020
rect -2680 5986 -2664 6020
rect -2606 5986 -2590 6020
rect -2522 5986 -2506 6020
rect -2448 5986 -2432 6020
rect -2364 5986 -2348 6020
rect -2290 5986 -2274 6020
rect -2206 5986 -2190 6020
rect -7052 5882 -7018 5944
rect -2044 5882 -2010 5944
rect -7052 5848 -6956 5882
rect -2106 5848 -2010 5882
rect -572 5986 -556 6020
rect -488 5986 -472 6020
rect -414 5986 -398 6020
rect -330 5986 -314 6020
rect -256 5986 -240 6020
rect -172 5986 -156 6020
rect -98 5986 -82 6020
rect -14 5986 2 6020
rect 60 5986 76 6020
rect 144 5986 160 6020
rect 218 5986 234 6020
rect 302 5986 318 6020
rect 376 5986 392 6020
rect 460 5986 476 6020
rect 534 5986 550 6020
rect 618 5986 634 6020
rect 692 5986 708 6020
rect 776 5986 792 6020
rect 850 5986 866 6020
rect 934 5986 950 6020
rect 1008 5986 1024 6020
rect 1092 5986 1108 6020
rect 1166 5986 1182 6020
rect 1250 5986 1266 6020
rect 1324 5986 1340 6020
rect 1408 5986 1424 6020
rect 1482 5986 1498 6020
rect 1566 5986 1582 6020
rect 1640 5986 1656 6020
rect 1724 5986 1740 6020
rect 1798 5986 1814 6020
rect 1882 5986 1898 6020
rect 1956 5986 1972 6020
rect 2040 5986 2056 6020
rect 2114 5986 2130 6020
rect 2198 5986 2214 6020
rect 2272 5986 2288 6020
rect 2356 5986 2372 6020
rect 2430 5986 2446 6020
rect 2514 5986 2530 6020
rect 2588 5986 2604 6020
rect 2672 5986 2688 6020
rect 2746 5986 2762 6020
rect 2830 5986 2846 6020
rect 2904 5986 2920 6020
rect 2988 5986 3004 6020
rect 3062 5986 3078 6020
rect 3146 5986 3162 6020
rect 3220 5986 3236 6020
rect 3304 5986 3320 6020
rect 3378 5986 3394 6020
rect 3462 5986 3478 6020
rect 3536 5986 3552 6020
rect 3620 5986 3636 6020
rect 3694 5986 3710 6020
rect 3778 5986 3794 6020
rect 3852 5986 3868 6020
rect 3936 5986 3952 6020
rect 4010 5986 4026 6020
rect 4094 5986 4110 6020
rect -752 5882 -718 5944
rect 4256 5882 4290 5944
rect -752 5848 -656 5882
rect 4194 5848 4290 5882
rect 5728 5986 5744 6020
rect 5812 5986 5828 6020
rect 5886 5986 5902 6020
rect 5970 5986 5986 6020
rect 6044 5986 6060 6020
rect 6128 5986 6144 6020
rect 6202 5986 6218 6020
rect 6286 5986 6302 6020
rect 6360 5986 6376 6020
rect 6444 5986 6460 6020
rect 6518 5986 6534 6020
rect 6602 5986 6618 6020
rect 6676 5986 6692 6020
rect 6760 5986 6776 6020
rect 6834 5986 6850 6020
rect 6918 5986 6934 6020
rect 6992 5986 7008 6020
rect 7076 5986 7092 6020
rect 7150 5986 7166 6020
rect 7234 5986 7250 6020
rect 7308 5986 7324 6020
rect 7392 5986 7408 6020
rect 7466 5986 7482 6020
rect 7550 5986 7566 6020
rect 7624 5986 7640 6020
rect 7708 5986 7724 6020
rect 7782 5986 7798 6020
rect 7866 5986 7882 6020
rect 7940 5986 7956 6020
rect 8024 5986 8040 6020
rect 8098 5986 8114 6020
rect 8182 5986 8198 6020
rect 8256 5986 8272 6020
rect 8340 5986 8356 6020
rect 8414 5986 8430 6020
rect 8498 5986 8514 6020
rect 8572 5986 8588 6020
rect 8656 5986 8672 6020
rect 8730 5986 8746 6020
rect 8814 5986 8830 6020
rect 8888 5986 8904 6020
rect 8972 5986 8988 6020
rect 9046 5986 9062 6020
rect 9130 5986 9146 6020
rect 9204 5986 9220 6020
rect 9288 5986 9304 6020
rect 9362 5986 9378 6020
rect 9446 5986 9462 6020
rect 9520 5986 9536 6020
rect 9604 5986 9620 6020
rect 9678 5986 9694 6020
rect 9762 5986 9778 6020
rect 9836 5986 9852 6020
rect 9920 5986 9936 6020
rect 9994 5986 10010 6020
rect 10078 5986 10094 6020
rect 10152 5986 10168 6020
rect 10236 5986 10252 6020
rect 10310 5986 10326 6020
rect 10394 5986 10410 6020
rect 5548 5882 5582 5944
rect 10556 5882 10590 5944
rect 5548 5848 5644 5882
rect 10494 5848 10590 5882
<< viali >>
rect -13164 49868 -8441 49870
rect -6864 49868 -2141 49870
rect -564 49868 4159 49870
rect 5736 49868 10459 49870
rect -13164 49834 -8441 49868
rect -13164 49832 -8441 49834
rect -13156 49696 -13088 49730
rect -12998 49696 -12930 49730
rect -12840 49696 -12772 49730
rect -12682 49696 -12614 49730
rect -12524 49696 -12456 49730
rect -12366 49696 -12298 49730
rect -12208 49696 -12140 49730
rect -12050 49696 -11982 49730
rect -11892 49696 -11824 49730
rect -11734 49696 -11666 49730
rect -11576 49696 -11508 49730
rect -11418 49696 -11350 49730
rect -11260 49696 -11192 49730
rect -11102 49696 -11034 49730
rect -10944 49696 -10876 49730
rect -10786 49696 -10718 49730
rect -10628 49696 -10560 49730
rect -10470 49696 -10402 49730
rect -10312 49696 -10244 49730
rect -10154 49696 -10086 49730
rect -9996 49696 -9928 49730
rect -9838 49696 -9770 49730
rect -9680 49696 -9612 49730
rect -9522 49696 -9454 49730
rect -9364 49696 -9296 49730
rect -9206 49696 -9138 49730
rect -9048 49696 -8980 49730
rect -8890 49696 -8822 49730
rect -8732 49696 -8664 49730
rect -8574 49696 -8506 49730
rect -6864 49834 -2141 49868
rect -6864 49832 -2141 49834
rect -6856 49696 -6788 49730
rect -6698 49696 -6630 49730
rect -6540 49696 -6472 49730
rect -6382 49696 -6314 49730
rect -6224 49696 -6156 49730
rect -6066 49696 -5998 49730
rect -5908 49696 -5840 49730
rect -5750 49696 -5682 49730
rect -5592 49696 -5524 49730
rect -5434 49696 -5366 49730
rect -5276 49696 -5208 49730
rect -5118 49696 -5050 49730
rect -4960 49696 -4892 49730
rect -4802 49696 -4734 49730
rect -4644 49696 -4576 49730
rect -4486 49696 -4418 49730
rect -4328 49696 -4260 49730
rect -4170 49696 -4102 49730
rect -4012 49696 -3944 49730
rect -3854 49696 -3786 49730
rect -3696 49696 -3628 49730
rect -3538 49696 -3470 49730
rect -3380 49696 -3312 49730
rect -3222 49696 -3154 49730
rect -3064 49696 -2996 49730
rect -2906 49696 -2838 49730
rect -2748 49696 -2680 49730
rect -2590 49696 -2522 49730
rect -2432 49696 -2364 49730
rect -2274 49696 -2206 49730
rect -564 49834 4159 49868
rect -564 49832 4159 49834
rect -556 49696 -488 49730
rect -398 49696 -330 49730
rect -240 49696 -172 49730
rect -82 49696 -14 49730
rect 76 49696 144 49730
rect 234 49696 302 49730
rect 392 49696 460 49730
rect 550 49696 618 49730
rect 708 49696 776 49730
rect 866 49696 934 49730
rect 1024 49696 1092 49730
rect 1182 49696 1250 49730
rect 1340 49696 1408 49730
rect 1498 49696 1566 49730
rect 1656 49696 1724 49730
rect 1814 49696 1882 49730
rect 1972 49696 2040 49730
rect 2130 49696 2198 49730
rect 2288 49696 2356 49730
rect 2446 49696 2514 49730
rect 2604 49696 2672 49730
rect 2762 49696 2830 49730
rect 2920 49696 2988 49730
rect 3078 49696 3146 49730
rect 3236 49696 3304 49730
rect 3394 49696 3462 49730
rect 3552 49696 3620 49730
rect 3710 49696 3778 49730
rect 3868 49696 3936 49730
rect 4026 49696 4094 49730
rect 5736 49834 10459 49868
rect 5736 49832 10459 49834
rect 5744 49696 5812 49730
rect 5902 49696 5970 49730
rect 6060 49696 6128 49730
rect 6218 49696 6286 49730
rect 6376 49696 6444 49730
rect 6534 49696 6602 49730
rect 6692 49696 6760 49730
rect 6850 49696 6918 49730
rect 7008 49696 7076 49730
rect 7166 49696 7234 49730
rect 7324 49696 7392 49730
rect 7482 49696 7550 49730
rect 7640 49696 7708 49730
rect 7798 49696 7866 49730
rect 7956 49696 8024 49730
rect 8114 49696 8182 49730
rect 8272 49696 8340 49730
rect 8430 49696 8498 49730
rect 8588 49696 8656 49730
rect 8746 49696 8814 49730
rect 8904 49696 8972 49730
rect 9062 49696 9130 49730
rect 9220 49696 9288 49730
rect 9378 49696 9446 49730
rect 9536 49696 9604 49730
rect 9694 49696 9762 49730
rect 9852 49696 9920 49730
rect 10010 49696 10078 49730
rect 10168 49696 10236 49730
rect 10326 49696 10394 49730
rect -13354 43636 -13352 49680
rect -13352 43636 -13318 49680
rect -13318 43636 -13316 49680
rect -13218 43670 -13184 49646
rect -13060 43670 -13026 49646
rect -12902 43670 -12868 49646
rect -12744 43670 -12710 49646
rect -12586 43670 -12552 49646
rect -12428 43670 -12394 49646
rect -12270 43670 -12236 49646
rect -12112 43670 -12078 49646
rect -11954 43670 -11920 49646
rect -11796 43670 -11762 49646
rect -11638 43670 -11604 49646
rect -11480 43670 -11446 49646
rect -11322 43670 -11288 49646
rect -11164 43670 -11130 49646
rect -11006 43670 -10972 49646
rect -10848 43670 -10814 49646
rect -10690 43670 -10656 49646
rect -10532 43670 -10498 49646
rect -10374 43670 -10340 49646
rect -10216 43670 -10182 49646
rect -10058 43670 -10024 49646
rect -9900 43670 -9866 49646
rect -9742 43670 -9708 49646
rect -9584 43670 -9550 49646
rect -9426 43670 -9392 49646
rect -9268 43670 -9234 49646
rect -9110 43670 -9076 49646
rect -8952 43670 -8918 49646
rect -8794 43670 -8760 49646
rect -8636 43670 -8602 49646
rect -8478 43670 -8444 49646
rect -8346 43636 -8344 49680
rect -8344 43636 -8310 49680
rect -8310 43636 -8308 49680
rect -7054 43636 -7052 49680
rect -7052 43636 -7018 49680
rect -7018 43636 -7016 49680
rect -6918 43670 -6884 49646
rect -6760 43670 -6726 49646
rect -6602 43670 -6568 49646
rect -6444 43670 -6410 49646
rect -6286 43670 -6252 49646
rect -6128 43670 -6094 49646
rect -5970 43670 -5936 49646
rect -5812 43670 -5778 49646
rect -5654 43670 -5620 49646
rect -5496 43670 -5462 49646
rect -5338 43670 -5304 49646
rect -5180 43670 -5146 49646
rect -5022 43670 -4988 49646
rect -4864 43670 -4830 49646
rect -4706 43670 -4672 49646
rect -4548 43670 -4514 49646
rect -4390 43670 -4356 49646
rect -4232 43670 -4198 49646
rect -4074 43670 -4040 49646
rect -3916 43670 -3882 49646
rect -3758 43670 -3724 49646
rect -3600 43670 -3566 49646
rect -3442 43670 -3408 49646
rect -3284 43670 -3250 49646
rect -3126 43670 -3092 49646
rect -2968 43670 -2934 49646
rect -2810 43670 -2776 49646
rect -2652 43670 -2618 49646
rect -2494 43670 -2460 49646
rect -2336 43670 -2302 49646
rect -2178 43670 -2144 49646
rect -2046 43636 -2044 49680
rect -2044 43636 -2010 49680
rect -2010 43636 -2008 49680
rect -754 43636 -752 49680
rect -752 43636 -718 49680
rect -718 43636 -716 49680
rect -618 43670 -584 49646
rect -460 43670 -426 49646
rect -302 43670 -268 49646
rect -144 43670 -110 49646
rect 14 43670 48 49646
rect 172 43670 206 49646
rect 330 43670 364 49646
rect 488 43670 522 49646
rect 646 43670 680 49646
rect 804 43670 838 49646
rect 962 43670 996 49646
rect 1120 43670 1154 49646
rect 1278 43670 1312 49646
rect 1436 43670 1470 49646
rect 1594 43670 1628 49646
rect 1752 43670 1786 49646
rect 1910 43670 1944 49646
rect 2068 43670 2102 49646
rect 2226 43670 2260 49646
rect 2384 43670 2418 49646
rect 2542 43670 2576 49646
rect 2700 43670 2734 49646
rect 2858 43670 2892 49646
rect 3016 43670 3050 49646
rect 3174 43670 3208 49646
rect 3332 43670 3366 49646
rect 3490 43670 3524 49646
rect 3648 43670 3682 49646
rect 3806 43670 3840 49646
rect 3964 43670 3998 49646
rect 4122 43670 4156 49646
rect 4254 43636 4256 49680
rect 4256 43636 4290 49680
rect 4290 43636 4292 49680
rect 5546 43636 5548 49680
rect 5548 43636 5582 49680
rect 5582 43636 5584 49680
rect 5682 43670 5716 49646
rect 5840 43670 5874 49646
rect 5998 43670 6032 49646
rect 6156 43670 6190 49646
rect 6314 43670 6348 49646
rect 6472 43670 6506 49646
rect 6630 43670 6664 49646
rect 6788 43670 6822 49646
rect 6946 43670 6980 49646
rect 7104 43670 7138 49646
rect 7262 43670 7296 49646
rect 7420 43670 7454 49646
rect 7578 43670 7612 49646
rect 7736 43670 7770 49646
rect 7894 43670 7928 49646
rect 8052 43670 8086 49646
rect 8210 43670 8244 49646
rect 8368 43670 8402 49646
rect 8526 43670 8560 49646
rect 8684 43670 8718 49646
rect 8842 43670 8876 49646
rect 9000 43670 9034 49646
rect 9158 43670 9192 49646
rect 9316 43670 9350 49646
rect 9474 43670 9508 49646
rect 9632 43670 9666 49646
rect 9790 43670 9824 49646
rect 9948 43670 9982 49646
rect 10106 43670 10140 49646
rect 10264 43670 10298 49646
rect 10422 43670 10456 49646
rect 10554 43636 10556 49680
rect 10556 43636 10590 49680
rect 10590 43636 10592 49680
rect -13156 43586 -13088 43620
rect -12998 43586 -12930 43620
rect -12840 43586 -12772 43620
rect -12682 43586 -12614 43620
rect -12524 43586 -12456 43620
rect -12366 43586 -12298 43620
rect -12208 43586 -12140 43620
rect -12050 43586 -11982 43620
rect -11892 43586 -11824 43620
rect -11734 43586 -11666 43620
rect -11576 43586 -11508 43620
rect -11418 43586 -11350 43620
rect -11260 43586 -11192 43620
rect -11102 43586 -11034 43620
rect -10944 43586 -10876 43620
rect -10786 43586 -10718 43620
rect -10628 43586 -10560 43620
rect -10470 43586 -10402 43620
rect -10312 43586 -10244 43620
rect -10154 43586 -10086 43620
rect -9996 43586 -9928 43620
rect -9838 43586 -9770 43620
rect -9680 43586 -9612 43620
rect -9522 43586 -9454 43620
rect -9364 43586 -9296 43620
rect -9206 43586 -9138 43620
rect -9048 43586 -8980 43620
rect -8890 43586 -8822 43620
rect -8732 43586 -8664 43620
rect -8574 43586 -8506 43620
rect -13164 43482 -8498 43484
rect -13164 43448 -8498 43482
rect -6856 43586 -6788 43620
rect -6698 43586 -6630 43620
rect -6540 43586 -6472 43620
rect -6382 43586 -6314 43620
rect -6224 43586 -6156 43620
rect -6066 43586 -5998 43620
rect -5908 43586 -5840 43620
rect -5750 43586 -5682 43620
rect -5592 43586 -5524 43620
rect -5434 43586 -5366 43620
rect -5276 43586 -5208 43620
rect -5118 43586 -5050 43620
rect -4960 43586 -4892 43620
rect -4802 43586 -4734 43620
rect -4644 43586 -4576 43620
rect -4486 43586 -4418 43620
rect -4328 43586 -4260 43620
rect -4170 43586 -4102 43620
rect -4012 43586 -3944 43620
rect -3854 43586 -3786 43620
rect -3696 43586 -3628 43620
rect -3538 43586 -3470 43620
rect -3380 43586 -3312 43620
rect -3222 43586 -3154 43620
rect -3064 43586 -2996 43620
rect -2906 43586 -2838 43620
rect -2748 43586 -2680 43620
rect -2590 43586 -2522 43620
rect -2432 43586 -2364 43620
rect -2274 43586 -2206 43620
rect -6864 43482 -2198 43484
rect -6864 43448 -2198 43482
rect -556 43586 -488 43620
rect -398 43586 -330 43620
rect -240 43586 -172 43620
rect -82 43586 -14 43620
rect 76 43586 144 43620
rect 234 43586 302 43620
rect 392 43586 460 43620
rect 550 43586 618 43620
rect 708 43586 776 43620
rect 866 43586 934 43620
rect 1024 43586 1092 43620
rect 1182 43586 1250 43620
rect 1340 43586 1408 43620
rect 1498 43586 1566 43620
rect 1656 43586 1724 43620
rect 1814 43586 1882 43620
rect 1972 43586 2040 43620
rect 2130 43586 2198 43620
rect 2288 43586 2356 43620
rect 2446 43586 2514 43620
rect 2604 43586 2672 43620
rect 2762 43586 2830 43620
rect 2920 43586 2988 43620
rect 3078 43586 3146 43620
rect 3236 43586 3304 43620
rect 3394 43586 3462 43620
rect 3552 43586 3620 43620
rect 3710 43586 3778 43620
rect 3868 43586 3936 43620
rect 4026 43586 4094 43620
rect -564 43482 4102 43484
rect -564 43448 4102 43482
rect 5744 43586 5812 43620
rect 5902 43586 5970 43620
rect 6060 43586 6128 43620
rect 6218 43586 6286 43620
rect 6376 43586 6444 43620
rect 6534 43586 6602 43620
rect 6692 43586 6760 43620
rect 6850 43586 6918 43620
rect 7008 43586 7076 43620
rect 7166 43586 7234 43620
rect 7324 43586 7392 43620
rect 7482 43586 7550 43620
rect 7640 43586 7708 43620
rect 7798 43586 7866 43620
rect 7956 43586 8024 43620
rect 8114 43586 8182 43620
rect 8272 43586 8340 43620
rect 8430 43586 8498 43620
rect 8588 43586 8656 43620
rect 8746 43586 8814 43620
rect 8904 43586 8972 43620
rect 9062 43586 9130 43620
rect 9220 43586 9288 43620
rect 9378 43586 9446 43620
rect 9536 43586 9604 43620
rect 9694 43586 9762 43620
rect 9852 43586 9920 43620
rect 10010 43586 10078 43620
rect 10168 43586 10236 43620
rect 10326 43586 10394 43620
rect 5736 43482 10402 43484
rect 5736 43448 10402 43482
rect -13164 43446 -8498 43448
rect -6864 43446 -2198 43448
rect -564 43446 4102 43448
rect 5736 43446 10402 43448
rect -13164 42868 -8441 42870
rect -6864 42868 -2141 42870
rect -564 42868 4159 42870
rect 5736 42868 10459 42870
rect -13164 42834 -8441 42868
rect -13164 42832 -8441 42834
rect -13156 42696 -13088 42730
rect -12998 42696 -12930 42730
rect -12840 42696 -12772 42730
rect -12682 42696 -12614 42730
rect -12524 42696 -12456 42730
rect -12366 42696 -12298 42730
rect -12208 42696 -12140 42730
rect -12050 42696 -11982 42730
rect -11892 42696 -11824 42730
rect -11734 42696 -11666 42730
rect -11576 42696 -11508 42730
rect -11418 42696 -11350 42730
rect -11260 42696 -11192 42730
rect -11102 42696 -11034 42730
rect -10944 42696 -10876 42730
rect -10786 42696 -10718 42730
rect -10628 42696 -10560 42730
rect -10470 42696 -10402 42730
rect -10312 42696 -10244 42730
rect -10154 42696 -10086 42730
rect -9996 42696 -9928 42730
rect -9838 42696 -9770 42730
rect -9680 42696 -9612 42730
rect -9522 42696 -9454 42730
rect -9364 42696 -9296 42730
rect -9206 42696 -9138 42730
rect -9048 42696 -8980 42730
rect -8890 42696 -8822 42730
rect -8732 42696 -8664 42730
rect -8574 42696 -8506 42730
rect -6864 42834 -2141 42868
rect -6864 42832 -2141 42834
rect -6856 42696 -6788 42730
rect -6698 42696 -6630 42730
rect -6540 42696 -6472 42730
rect -6382 42696 -6314 42730
rect -6224 42696 -6156 42730
rect -6066 42696 -5998 42730
rect -5908 42696 -5840 42730
rect -5750 42696 -5682 42730
rect -5592 42696 -5524 42730
rect -5434 42696 -5366 42730
rect -5276 42696 -5208 42730
rect -5118 42696 -5050 42730
rect -4960 42696 -4892 42730
rect -4802 42696 -4734 42730
rect -4644 42696 -4576 42730
rect -4486 42696 -4418 42730
rect -4328 42696 -4260 42730
rect -4170 42696 -4102 42730
rect -4012 42696 -3944 42730
rect -3854 42696 -3786 42730
rect -3696 42696 -3628 42730
rect -3538 42696 -3470 42730
rect -3380 42696 -3312 42730
rect -3222 42696 -3154 42730
rect -3064 42696 -2996 42730
rect -2906 42696 -2838 42730
rect -2748 42696 -2680 42730
rect -2590 42696 -2522 42730
rect -2432 42696 -2364 42730
rect -2274 42696 -2206 42730
rect -564 42834 4159 42868
rect -564 42832 4159 42834
rect -556 42696 -488 42730
rect -398 42696 -330 42730
rect -240 42696 -172 42730
rect -82 42696 -14 42730
rect 76 42696 144 42730
rect 234 42696 302 42730
rect 392 42696 460 42730
rect 550 42696 618 42730
rect 708 42696 776 42730
rect 866 42696 934 42730
rect 1024 42696 1092 42730
rect 1182 42696 1250 42730
rect 1340 42696 1408 42730
rect 1498 42696 1566 42730
rect 1656 42696 1724 42730
rect 1814 42696 1882 42730
rect 1972 42696 2040 42730
rect 2130 42696 2198 42730
rect 2288 42696 2356 42730
rect 2446 42696 2514 42730
rect 2604 42696 2672 42730
rect 2762 42696 2830 42730
rect 2920 42696 2988 42730
rect 3078 42696 3146 42730
rect 3236 42696 3304 42730
rect 3394 42696 3462 42730
rect 3552 42696 3620 42730
rect 3710 42696 3778 42730
rect 3868 42696 3936 42730
rect 4026 42696 4094 42730
rect 5736 42834 10459 42868
rect 5736 42832 10459 42834
rect 5744 42696 5812 42730
rect 5902 42696 5970 42730
rect 6060 42696 6128 42730
rect 6218 42696 6286 42730
rect 6376 42696 6444 42730
rect 6534 42696 6602 42730
rect 6692 42696 6760 42730
rect 6850 42696 6918 42730
rect 7008 42696 7076 42730
rect 7166 42696 7234 42730
rect 7324 42696 7392 42730
rect 7482 42696 7550 42730
rect 7640 42696 7708 42730
rect 7798 42696 7866 42730
rect 7956 42696 8024 42730
rect 8114 42696 8182 42730
rect 8272 42696 8340 42730
rect 8430 42696 8498 42730
rect 8588 42696 8656 42730
rect 8746 42696 8814 42730
rect 8904 42696 8972 42730
rect 9062 42696 9130 42730
rect 9220 42696 9288 42730
rect 9378 42696 9446 42730
rect 9536 42696 9604 42730
rect 9694 42696 9762 42730
rect 9852 42696 9920 42730
rect 10010 42696 10078 42730
rect 10168 42696 10236 42730
rect 10326 42696 10394 42730
rect -13354 36636 -13352 42680
rect -13352 36636 -13318 42680
rect -13318 36636 -13316 42680
rect -13218 36670 -13184 42646
rect -13060 36670 -13026 42646
rect -12902 36670 -12868 42646
rect -12744 36670 -12710 42646
rect -12586 36670 -12552 42646
rect -12428 36670 -12394 42646
rect -12270 36670 -12236 42646
rect -12112 36670 -12078 42646
rect -11954 36670 -11920 42646
rect -11796 36670 -11762 42646
rect -11638 36670 -11604 42646
rect -11480 36670 -11446 42646
rect -11322 36670 -11288 42646
rect -11164 36670 -11130 42646
rect -11006 36670 -10972 42646
rect -10848 36670 -10814 42646
rect -10690 36670 -10656 42646
rect -10532 36670 -10498 42646
rect -10374 36670 -10340 42646
rect -10216 36670 -10182 42646
rect -10058 36670 -10024 42646
rect -9900 36670 -9866 42646
rect -9742 36670 -9708 42646
rect -9584 36670 -9550 42646
rect -9426 36670 -9392 42646
rect -9268 36670 -9234 42646
rect -9110 36670 -9076 42646
rect -8952 36670 -8918 42646
rect -8794 36670 -8760 42646
rect -8636 36670 -8602 42646
rect -8478 36670 -8444 42646
rect -8346 36636 -8344 42680
rect -8344 36636 -8310 42680
rect -8310 36636 -8308 42680
rect -7054 36636 -7052 42680
rect -7052 36636 -7018 42680
rect -7018 36636 -7016 42680
rect -6918 36670 -6884 42646
rect -6760 36670 -6726 42646
rect -6602 36670 -6568 42646
rect -6444 36670 -6410 42646
rect -6286 36670 -6252 42646
rect -6128 36670 -6094 42646
rect -5970 36670 -5936 42646
rect -5812 36670 -5778 42646
rect -5654 36670 -5620 42646
rect -5496 36670 -5462 42646
rect -5338 36670 -5304 42646
rect -5180 36670 -5146 42646
rect -5022 36670 -4988 42646
rect -4864 36670 -4830 42646
rect -4706 36670 -4672 42646
rect -4548 36670 -4514 42646
rect -4390 36670 -4356 42646
rect -4232 36670 -4198 42646
rect -4074 36670 -4040 42646
rect -3916 36670 -3882 42646
rect -3758 36670 -3724 42646
rect -3600 36670 -3566 42646
rect -3442 36670 -3408 42646
rect -3284 36670 -3250 42646
rect -3126 36670 -3092 42646
rect -2968 36670 -2934 42646
rect -2810 36670 -2776 42646
rect -2652 36670 -2618 42646
rect -2494 36670 -2460 42646
rect -2336 36670 -2302 42646
rect -2178 36670 -2144 42646
rect -2046 36636 -2044 42680
rect -2044 36636 -2010 42680
rect -2010 36636 -2008 42680
rect -754 36636 -752 42680
rect -752 36636 -718 42680
rect -718 36636 -716 42680
rect -618 36670 -584 42646
rect -460 36670 -426 42646
rect -302 36670 -268 42646
rect -144 36670 -110 42646
rect 14 36670 48 42646
rect 172 36670 206 42646
rect 330 36670 364 42646
rect 488 36670 522 42646
rect 646 36670 680 42646
rect 804 36670 838 42646
rect 962 36670 996 42646
rect 1120 36670 1154 42646
rect 1278 36670 1312 42646
rect 1436 36670 1470 42646
rect 1594 36670 1628 42646
rect 1752 36670 1786 42646
rect 1910 36670 1944 42646
rect 2068 36670 2102 42646
rect 2226 36670 2260 42646
rect 2384 36670 2418 42646
rect 2542 36670 2576 42646
rect 2700 36670 2734 42646
rect 2858 36670 2892 42646
rect 3016 36670 3050 42646
rect 3174 36670 3208 42646
rect 3332 36670 3366 42646
rect 3490 36670 3524 42646
rect 3648 36670 3682 42646
rect 3806 36670 3840 42646
rect 3964 36670 3998 42646
rect 4122 36670 4156 42646
rect 4254 36636 4256 42680
rect 4256 36636 4290 42680
rect 4290 36636 4292 42680
rect 5546 36636 5548 42680
rect 5548 36636 5582 42680
rect 5582 36636 5584 42680
rect 5682 36670 5716 42646
rect 5840 36670 5874 42646
rect 5998 36670 6032 42646
rect 6156 36670 6190 42646
rect 6314 36670 6348 42646
rect 6472 36670 6506 42646
rect 6630 36670 6664 42646
rect 6788 36670 6822 42646
rect 6946 36670 6980 42646
rect 7104 36670 7138 42646
rect 7262 36670 7296 42646
rect 7420 36670 7454 42646
rect 7578 36670 7612 42646
rect 7736 36670 7770 42646
rect 7894 36670 7928 42646
rect 8052 36670 8086 42646
rect 8210 36670 8244 42646
rect 8368 36670 8402 42646
rect 8526 36670 8560 42646
rect 8684 36670 8718 42646
rect 8842 36670 8876 42646
rect 9000 36670 9034 42646
rect 9158 36670 9192 42646
rect 9316 36670 9350 42646
rect 9474 36670 9508 42646
rect 9632 36670 9666 42646
rect 9790 36670 9824 42646
rect 9948 36670 9982 42646
rect 10106 36670 10140 42646
rect 10264 36670 10298 42646
rect 10422 36670 10456 42646
rect 10554 36636 10556 42680
rect 10556 36636 10590 42680
rect 10590 36636 10592 42680
rect -13156 36586 -13088 36620
rect -12998 36586 -12930 36620
rect -12840 36586 -12772 36620
rect -12682 36586 -12614 36620
rect -12524 36586 -12456 36620
rect -12366 36586 -12298 36620
rect -12208 36586 -12140 36620
rect -12050 36586 -11982 36620
rect -11892 36586 -11824 36620
rect -11734 36586 -11666 36620
rect -11576 36586 -11508 36620
rect -11418 36586 -11350 36620
rect -11260 36586 -11192 36620
rect -11102 36586 -11034 36620
rect -10944 36586 -10876 36620
rect -10786 36586 -10718 36620
rect -10628 36586 -10560 36620
rect -10470 36586 -10402 36620
rect -10312 36586 -10244 36620
rect -10154 36586 -10086 36620
rect -9996 36586 -9928 36620
rect -9838 36586 -9770 36620
rect -9680 36586 -9612 36620
rect -9522 36586 -9454 36620
rect -9364 36586 -9296 36620
rect -9206 36586 -9138 36620
rect -9048 36586 -8980 36620
rect -8890 36586 -8822 36620
rect -8732 36586 -8664 36620
rect -8574 36586 -8506 36620
rect -13164 36482 -8498 36484
rect -13164 36448 -8498 36482
rect -6856 36586 -6788 36620
rect -6698 36586 -6630 36620
rect -6540 36586 -6472 36620
rect -6382 36586 -6314 36620
rect -6224 36586 -6156 36620
rect -6066 36586 -5998 36620
rect -5908 36586 -5840 36620
rect -5750 36586 -5682 36620
rect -5592 36586 -5524 36620
rect -5434 36586 -5366 36620
rect -5276 36586 -5208 36620
rect -5118 36586 -5050 36620
rect -4960 36586 -4892 36620
rect -4802 36586 -4734 36620
rect -4644 36586 -4576 36620
rect -4486 36586 -4418 36620
rect -4328 36586 -4260 36620
rect -4170 36586 -4102 36620
rect -4012 36586 -3944 36620
rect -3854 36586 -3786 36620
rect -3696 36586 -3628 36620
rect -3538 36586 -3470 36620
rect -3380 36586 -3312 36620
rect -3222 36586 -3154 36620
rect -3064 36586 -2996 36620
rect -2906 36586 -2838 36620
rect -2748 36586 -2680 36620
rect -2590 36586 -2522 36620
rect -2432 36586 -2364 36620
rect -2274 36586 -2206 36620
rect -6864 36482 -2198 36484
rect -6864 36448 -2198 36482
rect -556 36586 -488 36620
rect -398 36586 -330 36620
rect -240 36586 -172 36620
rect -82 36586 -14 36620
rect 76 36586 144 36620
rect 234 36586 302 36620
rect 392 36586 460 36620
rect 550 36586 618 36620
rect 708 36586 776 36620
rect 866 36586 934 36620
rect 1024 36586 1092 36620
rect 1182 36586 1250 36620
rect 1340 36586 1408 36620
rect 1498 36586 1566 36620
rect 1656 36586 1724 36620
rect 1814 36586 1882 36620
rect 1972 36586 2040 36620
rect 2130 36586 2198 36620
rect 2288 36586 2356 36620
rect 2446 36586 2514 36620
rect 2604 36586 2672 36620
rect 2762 36586 2830 36620
rect 2920 36586 2988 36620
rect 3078 36586 3146 36620
rect 3236 36586 3304 36620
rect 3394 36586 3462 36620
rect 3552 36586 3620 36620
rect 3710 36586 3778 36620
rect 3868 36586 3936 36620
rect 4026 36586 4094 36620
rect -564 36482 4102 36484
rect -564 36448 4102 36482
rect 5744 36586 5812 36620
rect 5902 36586 5970 36620
rect 6060 36586 6128 36620
rect 6218 36586 6286 36620
rect 6376 36586 6444 36620
rect 6534 36586 6602 36620
rect 6692 36586 6760 36620
rect 6850 36586 6918 36620
rect 7008 36586 7076 36620
rect 7166 36586 7234 36620
rect 7324 36586 7392 36620
rect 7482 36586 7550 36620
rect 7640 36586 7708 36620
rect 7798 36586 7866 36620
rect 7956 36586 8024 36620
rect 8114 36586 8182 36620
rect 8272 36586 8340 36620
rect 8430 36586 8498 36620
rect 8588 36586 8656 36620
rect 8746 36586 8814 36620
rect 8904 36586 8972 36620
rect 9062 36586 9130 36620
rect 9220 36586 9288 36620
rect 9378 36586 9446 36620
rect 9536 36586 9604 36620
rect 9694 36586 9762 36620
rect 9852 36586 9920 36620
rect 10010 36586 10078 36620
rect 10168 36586 10236 36620
rect 10326 36586 10394 36620
rect 5736 36482 10402 36484
rect 5736 36448 10402 36482
rect -13164 36446 -8498 36448
rect -6864 36446 -2198 36448
rect -564 36446 4102 36448
rect 5736 36446 10402 36448
rect -13164 34568 -8441 34570
rect -6864 34568 -2141 34570
rect -564 34568 4159 34570
rect 5736 34568 10459 34570
rect -13164 34534 -8441 34568
rect -13164 34532 -8441 34534
rect -13156 34396 -13088 34430
rect -12998 34396 -12930 34430
rect -12840 34396 -12772 34430
rect -12682 34396 -12614 34430
rect -12524 34396 -12456 34430
rect -12366 34396 -12298 34430
rect -12208 34396 -12140 34430
rect -12050 34396 -11982 34430
rect -11892 34396 -11824 34430
rect -11734 34396 -11666 34430
rect -11576 34396 -11508 34430
rect -11418 34396 -11350 34430
rect -11260 34396 -11192 34430
rect -11102 34396 -11034 34430
rect -10944 34396 -10876 34430
rect -10786 34396 -10718 34430
rect -10628 34396 -10560 34430
rect -10470 34396 -10402 34430
rect -10312 34396 -10244 34430
rect -10154 34396 -10086 34430
rect -9996 34396 -9928 34430
rect -9838 34396 -9770 34430
rect -9680 34396 -9612 34430
rect -9522 34396 -9454 34430
rect -9364 34396 -9296 34430
rect -9206 34396 -9138 34430
rect -9048 34396 -8980 34430
rect -8890 34396 -8822 34430
rect -8732 34396 -8664 34430
rect -8574 34396 -8506 34430
rect -6864 34534 -2141 34568
rect -6864 34532 -2141 34534
rect -6856 34396 -6788 34430
rect -6698 34396 -6630 34430
rect -6540 34396 -6472 34430
rect -6382 34396 -6314 34430
rect -6224 34396 -6156 34430
rect -6066 34396 -5998 34430
rect -5908 34396 -5840 34430
rect -5750 34396 -5682 34430
rect -5592 34396 -5524 34430
rect -5434 34396 -5366 34430
rect -5276 34396 -5208 34430
rect -5118 34396 -5050 34430
rect -4960 34396 -4892 34430
rect -4802 34396 -4734 34430
rect -4644 34396 -4576 34430
rect -4486 34396 -4418 34430
rect -4328 34396 -4260 34430
rect -4170 34396 -4102 34430
rect -4012 34396 -3944 34430
rect -3854 34396 -3786 34430
rect -3696 34396 -3628 34430
rect -3538 34396 -3470 34430
rect -3380 34396 -3312 34430
rect -3222 34396 -3154 34430
rect -3064 34396 -2996 34430
rect -2906 34396 -2838 34430
rect -2748 34396 -2680 34430
rect -2590 34396 -2522 34430
rect -2432 34396 -2364 34430
rect -2274 34396 -2206 34430
rect -564 34534 4159 34568
rect -564 34532 4159 34534
rect -556 34396 -488 34430
rect -398 34396 -330 34430
rect -240 34396 -172 34430
rect -82 34396 -14 34430
rect 76 34396 144 34430
rect 234 34396 302 34430
rect 392 34396 460 34430
rect 550 34396 618 34430
rect 708 34396 776 34430
rect 866 34396 934 34430
rect 1024 34396 1092 34430
rect 1182 34396 1250 34430
rect 1340 34396 1408 34430
rect 1498 34396 1566 34430
rect 1656 34396 1724 34430
rect 1814 34396 1882 34430
rect 1972 34396 2040 34430
rect 2130 34396 2198 34430
rect 2288 34396 2356 34430
rect 2446 34396 2514 34430
rect 2604 34396 2672 34430
rect 2762 34396 2830 34430
rect 2920 34396 2988 34430
rect 3078 34396 3146 34430
rect 3236 34396 3304 34430
rect 3394 34396 3462 34430
rect 3552 34396 3620 34430
rect 3710 34396 3778 34430
rect 3868 34396 3936 34430
rect 4026 34396 4094 34430
rect 5736 34534 10459 34568
rect 5736 34532 10459 34534
rect 5744 34396 5812 34430
rect 5902 34396 5970 34430
rect 6060 34396 6128 34430
rect 6218 34396 6286 34430
rect 6376 34396 6444 34430
rect 6534 34396 6602 34430
rect 6692 34396 6760 34430
rect 6850 34396 6918 34430
rect 7008 34396 7076 34430
rect 7166 34396 7234 34430
rect 7324 34396 7392 34430
rect 7482 34396 7550 34430
rect 7640 34396 7708 34430
rect 7798 34396 7866 34430
rect 7956 34396 8024 34430
rect 8114 34396 8182 34430
rect 8272 34396 8340 34430
rect 8430 34396 8498 34430
rect 8588 34396 8656 34430
rect 8746 34396 8814 34430
rect 8904 34396 8972 34430
rect 9062 34396 9130 34430
rect 9220 34396 9288 34430
rect 9378 34396 9446 34430
rect 9536 34396 9604 34430
rect 9694 34396 9762 34430
rect 9852 34396 9920 34430
rect 10010 34396 10078 34430
rect 10168 34396 10236 34430
rect 10326 34396 10394 34430
rect -13354 28336 -13352 34380
rect -13352 28336 -13318 34380
rect -13318 28336 -13316 34380
rect -13218 28370 -13184 34346
rect -13060 28370 -13026 34346
rect -12902 28370 -12868 34346
rect -12744 28370 -12710 34346
rect -12586 28370 -12552 34346
rect -12428 28370 -12394 34346
rect -12270 28370 -12236 34346
rect -12112 28370 -12078 34346
rect -11954 28370 -11920 34346
rect -11796 28370 -11762 34346
rect -11638 28370 -11604 34346
rect -11480 28370 -11446 34346
rect -11322 28370 -11288 34346
rect -11164 28370 -11130 34346
rect -11006 28370 -10972 34346
rect -10848 28370 -10814 34346
rect -10690 28370 -10656 34346
rect -10532 28370 -10498 34346
rect -10374 28370 -10340 34346
rect -10216 28370 -10182 34346
rect -10058 28370 -10024 34346
rect -9900 28370 -9866 34346
rect -9742 28370 -9708 34346
rect -9584 28370 -9550 34346
rect -9426 28370 -9392 34346
rect -9268 28370 -9234 34346
rect -9110 28370 -9076 34346
rect -8952 28370 -8918 34346
rect -8794 28370 -8760 34346
rect -8636 28370 -8602 34346
rect -8478 28370 -8444 34346
rect -8346 28336 -8344 34380
rect -8344 28336 -8310 34380
rect -8310 28336 -8308 34380
rect -7054 28336 -7052 34380
rect -7052 28336 -7018 34380
rect -7018 28336 -7016 34380
rect -6918 28370 -6884 34346
rect -6760 28370 -6726 34346
rect -6602 28370 -6568 34346
rect -6444 28370 -6410 34346
rect -6286 28370 -6252 34346
rect -6128 28370 -6094 34346
rect -5970 28370 -5936 34346
rect -5812 28370 -5778 34346
rect -5654 28370 -5620 34346
rect -5496 28370 -5462 34346
rect -5338 28370 -5304 34346
rect -5180 28370 -5146 34346
rect -5022 28370 -4988 34346
rect -4864 28370 -4830 34346
rect -4706 28370 -4672 34346
rect -4548 28370 -4514 34346
rect -4390 28370 -4356 34346
rect -4232 28370 -4198 34346
rect -4074 28370 -4040 34346
rect -3916 28370 -3882 34346
rect -3758 28370 -3724 34346
rect -3600 28370 -3566 34346
rect -3442 28370 -3408 34346
rect -3284 28370 -3250 34346
rect -3126 28370 -3092 34346
rect -2968 28370 -2934 34346
rect -2810 28370 -2776 34346
rect -2652 28370 -2618 34346
rect -2494 28370 -2460 34346
rect -2336 28370 -2302 34346
rect -2178 28370 -2144 34346
rect -2046 28336 -2044 34380
rect -2044 28336 -2010 34380
rect -2010 28336 -2008 34380
rect -754 28336 -752 34380
rect -752 28336 -718 34380
rect -718 28336 -716 34380
rect -618 28370 -584 34346
rect -460 28370 -426 34346
rect -302 28370 -268 34346
rect -144 28370 -110 34346
rect 14 28370 48 34346
rect 172 28370 206 34346
rect 330 28370 364 34346
rect 488 28370 522 34346
rect 646 28370 680 34346
rect 804 28370 838 34346
rect 962 28370 996 34346
rect 1120 28370 1154 34346
rect 1278 28370 1312 34346
rect 1436 28370 1470 34346
rect 1594 28370 1628 34346
rect 1752 28370 1786 34346
rect 1910 28370 1944 34346
rect 2068 28370 2102 34346
rect 2226 28370 2260 34346
rect 2384 28370 2418 34346
rect 2542 28370 2576 34346
rect 2700 28370 2734 34346
rect 2858 28370 2892 34346
rect 3016 28370 3050 34346
rect 3174 28370 3208 34346
rect 3332 28370 3366 34346
rect 3490 28370 3524 34346
rect 3648 28370 3682 34346
rect 3806 28370 3840 34346
rect 3964 28370 3998 34346
rect 4122 28370 4156 34346
rect 4254 28336 4256 34380
rect 4256 28336 4290 34380
rect 4290 28336 4292 34380
rect 5546 28336 5548 34380
rect 5548 28336 5582 34380
rect 5582 28336 5584 34380
rect 5682 28370 5716 34346
rect 5840 28370 5874 34346
rect 5998 28370 6032 34346
rect 6156 28370 6190 34346
rect 6314 28370 6348 34346
rect 6472 28370 6506 34346
rect 6630 28370 6664 34346
rect 6788 28370 6822 34346
rect 6946 28370 6980 34346
rect 7104 28370 7138 34346
rect 7262 28370 7296 34346
rect 7420 28370 7454 34346
rect 7578 28370 7612 34346
rect 7736 28370 7770 34346
rect 7894 28370 7928 34346
rect 8052 28370 8086 34346
rect 8210 28370 8244 34346
rect 8368 28370 8402 34346
rect 8526 28370 8560 34346
rect 8684 28370 8718 34346
rect 8842 28370 8876 34346
rect 9000 28370 9034 34346
rect 9158 28370 9192 34346
rect 9316 28370 9350 34346
rect 9474 28370 9508 34346
rect 9632 28370 9666 34346
rect 9790 28370 9824 34346
rect 9948 28370 9982 34346
rect 10106 28370 10140 34346
rect 10264 28370 10298 34346
rect 10422 28370 10456 34346
rect 10554 28336 10556 34380
rect 10556 28336 10590 34380
rect 10590 28336 10592 34380
rect -13156 28286 -13088 28320
rect -12998 28286 -12930 28320
rect -12840 28286 -12772 28320
rect -12682 28286 -12614 28320
rect -12524 28286 -12456 28320
rect -12366 28286 -12298 28320
rect -12208 28286 -12140 28320
rect -12050 28286 -11982 28320
rect -11892 28286 -11824 28320
rect -11734 28286 -11666 28320
rect -11576 28286 -11508 28320
rect -11418 28286 -11350 28320
rect -11260 28286 -11192 28320
rect -11102 28286 -11034 28320
rect -10944 28286 -10876 28320
rect -10786 28286 -10718 28320
rect -10628 28286 -10560 28320
rect -10470 28286 -10402 28320
rect -10312 28286 -10244 28320
rect -10154 28286 -10086 28320
rect -9996 28286 -9928 28320
rect -9838 28286 -9770 28320
rect -9680 28286 -9612 28320
rect -9522 28286 -9454 28320
rect -9364 28286 -9296 28320
rect -9206 28286 -9138 28320
rect -9048 28286 -8980 28320
rect -8890 28286 -8822 28320
rect -8732 28286 -8664 28320
rect -8574 28286 -8506 28320
rect -13164 28182 -8498 28184
rect -13164 28148 -8498 28182
rect -6856 28286 -6788 28320
rect -6698 28286 -6630 28320
rect -6540 28286 -6472 28320
rect -6382 28286 -6314 28320
rect -6224 28286 -6156 28320
rect -6066 28286 -5998 28320
rect -5908 28286 -5840 28320
rect -5750 28286 -5682 28320
rect -5592 28286 -5524 28320
rect -5434 28286 -5366 28320
rect -5276 28286 -5208 28320
rect -5118 28286 -5050 28320
rect -4960 28286 -4892 28320
rect -4802 28286 -4734 28320
rect -4644 28286 -4576 28320
rect -4486 28286 -4418 28320
rect -4328 28286 -4260 28320
rect -4170 28286 -4102 28320
rect -4012 28286 -3944 28320
rect -3854 28286 -3786 28320
rect -3696 28286 -3628 28320
rect -3538 28286 -3470 28320
rect -3380 28286 -3312 28320
rect -3222 28286 -3154 28320
rect -3064 28286 -2996 28320
rect -2906 28286 -2838 28320
rect -2748 28286 -2680 28320
rect -2590 28286 -2522 28320
rect -2432 28286 -2364 28320
rect -2274 28286 -2206 28320
rect -6864 28182 -2198 28184
rect -6864 28148 -2198 28182
rect -556 28286 -488 28320
rect -398 28286 -330 28320
rect -240 28286 -172 28320
rect -82 28286 -14 28320
rect 76 28286 144 28320
rect 234 28286 302 28320
rect 392 28286 460 28320
rect 550 28286 618 28320
rect 708 28286 776 28320
rect 866 28286 934 28320
rect 1024 28286 1092 28320
rect 1182 28286 1250 28320
rect 1340 28286 1408 28320
rect 1498 28286 1566 28320
rect 1656 28286 1724 28320
rect 1814 28286 1882 28320
rect 1972 28286 2040 28320
rect 2130 28286 2198 28320
rect 2288 28286 2356 28320
rect 2446 28286 2514 28320
rect 2604 28286 2672 28320
rect 2762 28286 2830 28320
rect 2920 28286 2988 28320
rect 3078 28286 3146 28320
rect 3236 28286 3304 28320
rect 3394 28286 3462 28320
rect 3552 28286 3620 28320
rect 3710 28286 3778 28320
rect 3868 28286 3936 28320
rect 4026 28286 4094 28320
rect -564 28182 4102 28184
rect -564 28148 4102 28182
rect 5744 28286 5812 28320
rect 5902 28286 5970 28320
rect 6060 28286 6128 28320
rect 6218 28286 6286 28320
rect 6376 28286 6444 28320
rect 6534 28286 6602 28320
rect 6692 28286 6760 28320
rect 6850 28286 6918 28320
rect 7008 28286 7076 28320
rect 7166 28286 7234 28320
rect 7324 28286 7392 28320
rect 7482 28286 7550 28320
rect 7640 28286 7708 28320
rect 7798 28286 7866 28320
rect 7956 28286 8024 28320
rect 8114 28286 8182 28320
rect 8272 28286 8340 28320
rect 8430 28286 8498 28320
rect 8588 28286 8656 28320
rect 8746 28286 8814 28320
rect 8904 28286 8972 28320
rect 9062 28286 9130 28320
rect 9220 28286 9288 28320
rect 9378 28286 9446 28320
rect 9536 28286 9604 28320
rect 9694 28286 9762 28320
rect 9852 28286 9920 28320
rect 10010 28286 10078 28320
rect 10168 28286 10236 28320
rect 10326 28286 10394 28320
rect 5736 28182 10402 28184
rect 5736 28148 10402 28182
rect -13164 28146 -8498 28148
rect -6864 28146 -2198 28148
rect -564 28146 4102 28148
rect 5736 28146 10402 28148
rect -13164 27568 -8441 27570
rect -6864 27568 -2141 27570
rect -564 27568 4159 27570
rect 5736 27568 10459 27570
rect -13164 27534 -8441 27568
rect -13164 27532 -8441 27534
rect -13156 27396 -13088 27430
rect -12998 27396 -12930 27430
rect -12840 27396 -12772 27430
rect -12682 27396 -12614 27430
rect -12524 27396 -12456 27430
rect -12366 27396 -12298 27430
rect -12208 27396 -12140 27430
rect -12050 27396 -11982 27430
rect -11892 27396 -11824 27430
rect -11734 27396 -11666 27430
rect -11576 27396 -11508 27430
rect -11418 27396 -11350 27430
rect -11260 27396 -11192 27430
rect -11102 27396 -11034 27430
rect -10944 27396 -10876 27430
rect -10786 27396 -10718 27430
rect -10628 27396 -10560 27430
rect -10470 27396 -10402 27430
rect -10312 27396 -10244 27430
rect -10154 27396 -10086 27430
rect -9996 27396 -9928 27430
rect -9838 27396 -9770 27430
rect -9680 27396 -9612 27430
rect -9522 27396 -9454 27430
rect -9364 27396 -9296 27430
rect -9206 27396 -9138 27430
rect -9048 27396 -8980 27430
rect -8890 27396 -8822 27430
rect -8732 27396 -8664 27430
rect -8574 27396 -8506 27430
rect -6864 27534 -2141 27568
rect -6864 27532 -2141 27534
rect -6856 27396 -6788 27430
rect -6698 27396 -6630 27430
rect -6540 27396 -6472 27430
rect -6382 27396 -6314 27430
rect -6224 27396 -6156 27430
rect -6066 27396 -5998 27430
rect -5908 27396 -5840 27430
rect -5750 27396 -5682 27430
rect -5592 27396 -5524 27430
rect -5434 27396 -5366 27430
rect -5276 27396 -5208 27430
rect -5118 27396 -5050 27430
rect -4960 27396 -4892 27430
rect -4802 27396 -4734 27430
rect -4644 27396 -4576 27430
rect -4486 27396 -4418 27430
rect -4328 27396 -4260 27430
rect -4170 27396 -4102 27430
rect -4012 27396 -3944 27430
rect -3854 27396 -3786 27430
rect -3696 27396 -3628 27430
rect -3538 27396 -3470 27430
rect -3380 27396 -3312 27430
rect -3222 27396 -3154 27430
rect -3064 27396 -2996 27430
rect -2906 27396 -2838 27430
rect -2748 27396 -2680 27430
rect -2590 27396 -2522 27430
rect -2432 27396 -2364 27430
rect -2274 27396 -2206 27430
rect -564 27534 4159 27568
rect -564 27532 4159 27534
rect -556 27396 -488 27430
rect -398 27396 -330 27430
rect -240 27396 -172 27430
rect -82 27396 -14 27430
rect 76 27396 144 27430
rect 234 27396 302 27430
rect 392 27396 460 27430
rect 550 27396 618 27430
rect 708 27396 776 27430
rect 866 27396 934 27430
rect 1024 27396 1092 27430
rect 1182 27396 1250 27430
rect 1340 27396 1408 27430
rect 1498 27396 1566 27430
rect 1656 27396 1724 27430
rect 1814 27396 1882 27430
rect 1972 27396 2040 27430
rect 2130 27396 2198 27430
rect 2288 27396 2356 27430
rect 2446 27396 2514 27430
rect 2604 27396 2672 27430
rect 2762 27396 2830 27430
rect 2920 27396 2988 27430
rect 3078 27396 3146 27430
rect 3236 27396 3304 27430
rect 3394 27396 3462 27430
rect 3552 27396 3620 27430
rect 3710 27396 3778 27430
rect 3868 27396 3936 27430
rect 4026 27396 4094 27430
rect 5736 27534 10459 27568
rect 5736 27532 10459 27534
rect 5744 27396 5812 27430
rect 5902 27396 5970 27430
rect 6060 27396 6128 27430
rect 6218 27396 6286 27430
rect 6376 27396 6444 27430
rect 6534 27396 6602 27430
rect 6692 27396 6760 27430
rect 6850 27396 6918 27430
rect 7008 27396 7076 27430
rect 7166 27396 7234 27430
rect 7324 27396 7392 27430
rect 7482 27396 7550 27430
rect 7640 27396 7708 27430
rect 7798 27396 7866 27430
rect 7956 27396 8024 27430
rect 8114 27396 8182 27430
rect 8272 27396 8340 27430
rect 8430 27396 8498 27430
rect 8588 27396 8656 27430
rect 8746 27396 8814 27430
rect 8904 27396 8972 27430
rect 9062 27396 9130 27430
rect 9220 27396 9288 27430
rect 9378 27396 9446 27430
rect 9536 27396 9604 27430
rect 9694 27396 9762 27430
rect 9852 27396 9920 27430
rect 10010 27396 10078 27430
rect 10168 27396 10236 27430
rect 10326 27396 10394 27430
rect -13354 21336 -13352 27380
rect -13352 21336 -13318 27380
rect -13318 21336 -13316 27380
rect -13218 21370 -13184 27346
rect -13060 21370 -13026 27346
rect -12902 21370 -12868 27346
rect -12744 21370 -12710 27346
rect -12586 21370 -12552 27346
rect -12428 21370 -12394 27346
rect -12270 21370 -12236 27346
rect -12112 21370 -12078 27346
rect -11954 21370 -11920 27346
rect -11796 21370 -11762 27346
rect -11638 21370 -11604 27346
rect -11480 21370 -11446 27346
rect -11322 21370 -11288 27346
rect -11164 21370 -11130 27346
rect -11006 21370 -10972 27346
rect -10848 21370 -10814 27346
rect -10690 21370 -10656 27346
rect -10532 21370 -10498 27346
rect -10374 21370 -10340 27346
rect -10216 21370 -10182 27346
rect -10058 21370 -10024 27346
rect -9900 21370 -9866 27346
rect -9742 21370 -9708 27346
rect -9584 21370 -9550 27346
rect -9426 21370 -9392 27346
rect -9268 21370 -9234 27346
rect -9110 21370 -9076 27346
rect -8952 21370 -8918 27346
rect -8794 21370 -8760 27346
rect -8636 21370 -8602 27346
rect -8478 21370 -8444 27346
rect -8346 21336 -8344 27380
rect -8344 21336 -8310 27380
rect -8310 21336 -8308 27380
rect -7054 21336 -7052 27380
rect -7052 21336 -7018 27380
rect -7018 21336 -7016 27380
rect -6918 21370 -6884 27346
rect -6760 21370 -6726 27346
rect -6602 21370 -6568 27346
rect -6444 21370 -6410 27346
rect -6286 21370 -6252 27346
rect -6128 21370 -6094 27346
rect -5970 21370 -5936 27346
rect -5812 21370 -5778 27346
rect -5654 21370 -5620 27346
rect -5496 21370 -5462 27346
rect -5338 21370 -5304 27346
rect -5180 21370 -5146 27346
rect -5022 21370 -4988 27346
rect -4864 21370 -4830 27346
rect -4706 21370 -4672 27346
rect -4548 21370 -4514 27346
rect -4390 21370 -4356 27346
rect -4232 21370 -4198 27346
rect -4074 21370 -4040 27346
rect -3916 21370 -3882 27346
rect -3758 21370 -3724 27346
rect -3600 21370 -3566 27346
rect -3442 21370 -3408 27346
rect -3284 21370 -3250 27346
rect -3126 21370 -3092 27346
rect -2968 21370 -2934 27346
rect -2810 21370 -2776 27346
rect -2652 21370 -2618 27346
rect -2494 21370 -2460 27346
rect -2336 21370 -2302 27346
rect -2178 21370 -2144 27346
rect -2046 21336 -2044 27380
rect -2044 21336 -2010 27380
rect -2010 21336 -2008 27380
rect -754 21336 -752 27380
rect -752 21336 -718 27380
rect -718 21336 -716 27380
rect -618 21370 -584 27346
rect -460 21370 -426 27346
rect -302 21370 -268 27346
rect -144 21370 -110 27346
rect 14 21370 48 27346
rect 172 21370 206 27346
rect 330 21370 364 27346
rect 488 21370 522 27346
rect 646 21370 680 27346
rect 804 21370 838 27346
rect 962 21370 996 27346
rect 1120 21370 1154 27346
rect 1278 21370 1312 27346
rect 1436 21370 1470 27346
rect 1594 21370 1628 27346
rect 1752 21370 1786 27346
rect 1910 21370 1944 27346
rect 2068 21370 2102 27346
rect 2226 21370 2260 27346
rect 2384 21370 2418 27346
rect 2542 21370 2576 27346
rect 2700 21370 2734 27346
rect 2858 21370 2892 27346
rect 3016 21370 3050 27346
rect 3174 21370 3208 27346
rect 3332 21370 3366 27346
rect 3490 21370 3524 27346
rect 3648 21370 3682 27346
rect 3806 21370 3840 27346
rect 3964 21370 3998 27346
rect 4122 21370 4156 27346
rect 4254 21336 4256 27380
rect 4256 21336 4290 27380
rect 4290 21336 4292 27380
rect 5546 21336 5548 27380
rect 5548 21336 5582 27380
rect 5582 21336 5584 27380
rect 5682 21370 5716 27346
rect 5840 21370 5874 27346
rect 5998 21370 6032 27346
rect 6156 21370 6190 27346
rect 6314 21370 6348 27346
rect 6472 21370 6506 27346
rect 6630 21370 6664 27346
rect 6788 21370 6822 27346
rect 6946 21370 6980 27346
rect 7104 21370 7138 27346
rect 7262 21370 7296 27346
rect 7420 21370 7454 27346
rect 7578 21370 7612 27346
rect 7736 21370 7770 27346
rect 7894 21370 7928 27346
rect 8052 21370 8086 27346
rect 8210 21370 8244 27346
rect 8368 21370 8402 27346
rect 8526 21370 8560 27346
rect 8684 21370 8718 27346
rect 8842 21370 8876 27346
rect 9000 21370 9034 27346
rect 9158 21370 9192 27346
rect 9316 21370 9350 27346
rect 9474 21370 9508 27346
rect 9632 21370 9666 27346
rect 9790 21370 9824 27346
rect 9948 21370 9982 27346
rect 10106 21370 10140 27346
rect 10264 21370 10298 27346
rect 10422 21370 10456 27346
rect 10554 21336 10556 27380
rect 10556 21336 10590 27380
rect 10590 21336 10592 27380
rect -13156 21286 -13088 21320
rect -12998 21286 -12930 21320
rect -12840 21286 -12772 21320
rect -12682 21286 -12614 21320
rect -12524 21286 -12456 21320
rect -12366 21286 -12298 21320
rect -12208 21286 -12140 21320
rect -12050 21286 -11982 21320
rect -11892 21286 -11824 21320
rect -11734 21286 -11666 21320
rect -11576 21286 -11508 21320
rect -11418 21286 -11350 21320
rect -11260 21286 -11192 21320
rect -11102 21286 -11034 21320
rect -10944 21286 -10876 21320
rect -10786 21286 -10718 21320
rect -10628 21286 -10560 21320
rect -10470 21286 -10402 21320
rect -10312 21286 -10244 21320
rect -10154 21286 -10086 21320
rect -9996 21286 -9928 21320
rect -9838 21286 -9770 21320
rect -9680 21286 -9612 21320
rect -9522 21286 -9454 21320
rect -9364 21286 -9296 21320
rect -9206 21286 -9138 21320
rect -9048 21286 -8980 21320
rect -8890 21286 -8822 21320
rect -8732 21286 -8664 21320
rect -8574 21286 -8506 21320
rect -13164 21182 -8498 21184
rect -13164 21148 -8498 21182
rect -6856 21286 -6788 21320
rect -6698 21286 -6630 21320
rect -6540 21286 -6472 21320
rect -6382 21286 -6314 21320
rect -6224 21286 -6156 21320
rect -6066 21286 -5998 21320
rect -5908 21286 -5840 21320
rect -5750 21286 -5682 21320
rect -5592 21286 -5524 21320
rect -5434 21286 -5366 21320
rect -5276 21286 -5208 21320
rect -5118 21286 -5050 21320
rect -4960 21286 -4892 21320
rect -4802 21286 -4734 21320
rect -4644 21286 -4576 21320
rect -4486 21286 -4418 21320
rect -4328 21286 -4260 21320
rect -4170 21286 -4102 21320
rect -4012 21286 -3944 21320
rect -3854 21286 -3786 21320
rect -3696 21286 -3628 21320
rect -3538 21286 -3470 21320
rect -3380 21286 -3312 21320
rect -3222 21286 -3154 21320
rect -3064 21286 -2996 21320
rect -2906 21286 -2838 21320
rect -2748 21286 -2680 21320
rect -2590 21286 -2522 21320
rect -2432 21286 -2364 21320
rect -2274 21286 -2206 21320
rect -6864 21182 -2198 21184
rect -6864 21148 -2198 21182
rect -556 21286 -488 21320
rect -398 21286 -330 21320
rect -240 21286 -172 21320
rect -82 21286 -14 21320
rect 76 21286 144 21320
rect 234 21286 302 21320
rect 392 21286 460 21320
rect 550 21286 618 21320
rect 708 21286 776 21320
rect 866 21286 934 21320
rect 1024 21286 1092 21320
rect 1182 21286 1250 21320
rect 1340 21286 1408 21320
rect 1498 21286 1566 21320
rect 1656 21286 1724 21320
rect 1814 21286 1882 21320
rect 1972 21286 2040 21320
rect 2130 21286 2198 21320
rect 2288 21286 2356 21320
rect 2446 21286 2514 21320
rect 2604 21286 2672 21320
rect 2762 21286 2830 21320
rect 2920 21286 2988 21320
rect 3078 21286 3146 21320
rect 3236 21286 3304 21320
rect 3394 21286 3462 21320
rect 3552 21286 3620 21320
rect 3710 21286 3778 21320
rect 3868 21286 3936 21320
rect 4026 21286 4094 21320
rect -564 21182 4102 21184
rect -564 21148 4102 21182
rect 5744 21286 5812 21320
rect 5902 21286 5970 21320
rect 6060 21286 6128 21320
rect 6218 21286 6286 21320
rect 6376 21286 6444 21320
rect 6534 21286 6602 21320
rect 6692 21286 6760 21320
rect 6850 21286 6918 21320
rect 7008 21286 7076 21320
rect 7166 21286 7234 21320
rect 7324 21286 7392 21320
rect 7482 21286 7550 21320
rect 7640 21286 7708 21320
rect 7798 21286 7866 21320
rect 7956 21286 8024 21320
rect 8114 21286 8182 21320
rect 8272 21286 8340 21320
rect 8430 21286 8498 21320
rect 8588 21286 8656 21320
rect 8746 21286 8814 21320
rect 8904 21286 8972 21320
rect 9062 21286 9130 21320
rect 9220 21286 9288 21320
rect 9378 21286 9446 21320
rect 9536 21286 9604 21320
rect 9694 21286 9762 21320
rect 9852 21286 9920 21320
rect 10010 21286 10078 21320
rect 10168 21286 10236 21320
rect 10326 21286 10394 21320
rect 5736 21182 10402 21184
rect 5736 21148 10402 21182
rect -13164 21146 -8498 21148
rect -6864 21146 -2198 21148
rect -564 21146 4102 21148
rect 5736 21146 10402 21148
rect -13164 19268 -8441 19270
rect -6864 19268 -2141 19270
rect -564 19268 4159 19270
rect 5736 19268 10459 19270
rect -13164 19234 -8441 19268
rect -13164 19232 -8441 19234
rect -13156 19096 -13088 19130
rect -12998 19096 -12930 19130
rect -12840 19096 -12772 19130
rect -12682 19096 -12614 19130
rect -12524 19096 -12456 19130
rect -12366 19096 -12298 19130
rect -12208 19096 -12140 19130
rect -12050 19096 -11982 19130
rect -11892 19096 -11824 19130
rect -11734 19096 -11666 19130
rect -11576 19096 -11508 19130
rect -11418 19096 -11350 19130
rect -11260 19096 -11192 19130
rect -11102 19096 -11034 19130
rect -10944 19096 -10876 19130
rect -10786 19096 -10718 19130
rect -10628 19096 -10560 19130
rect -10470 19096 -10402 19130
rect -10312 19096 -10244 19130
rect -10154 19096 -10086 19130
rect -9996 19096 -9928 19130
rect -9838 19096 -9770 19130
rect -9680 19096 -9612 19130
rect -9522 19096 -9454 19130
rect -9364 19096 -9296 19130
rect -9206 19096 -9138 19130
rect -9048 19096 -8980 19130
rect -8890 19096 -8822 19130
rect -8732 19096 -8664 19130
rect -8574 19096 -8506 19130
rect -6864 19234 -2141 19268
rect -6864 19232 -2141 19234
rect -6856 19096 -6788 19130
rect -6698 19096 -6630 19130
rect -6540 19096 -6472 19130
rect -6382 19096 -6314 19130
rect -6224 19096 -6156 19130
rect -6066 19096 -5998 19130
rect -5908 19096 -5840 19130
rect -5750 19096 -5682 19130
rect -5592 19096 -5524 19130
rect -5434 19096 -5366 19130
rect -5276 19096 -5208 19130
rect -5118 19096 -5050 19130
rect -4960 19096 -4892 19130
rect -4802 19096 -4734 19130
rect -4644 19096 -4576 19130
rect -4486 19096 -4418 19130
rect -4328 19096 -4260 19130
rect -4170 19096 -4102 19130
rect -4012 19096 -3944 19130
rect -3854 19096 -3786 19130
rect -3696 19096 -3628 19130
rect -3538 19096 -3470 19130
rect -3380 19096 -3312 19130
rect -3222 19096 -3154 19130
rect -3064 19096 -2996 19130
rect -2906 19096 -2838 19130
rect -2748 19096 -2680 19130
rect -2590 19096 -2522 19130
rect -2432 19096 -2364 19130
rect -2274 19096 -2206 19130
rect -564 19234 4159 19268
rect -564 19232 4159 19234
rect -556 19096 -488 19130
rect -398 19096 -330 19130
rect -240 19096 -172 19130
rect -82 19096 -14 19130
rect 76 19096 144 19130
rect 234 19096 302 19130
rect 392 19096 460 19130
rect 550 19096 618 19130
rect 708 19096 776 19130
rect 866 19096 934 19130
rect 1024 19096 1092 19130
rect 1182 19096 1250 19130
rect 1340 19096 1408 19130
rect 1498 19096 1566 19130
rect 1656 19096 1724 19130
rect 1814 19096 1882 19130
rect 1972 19096 2040 19130
rect 2130 19096 2198 19130
rect 2288 19096 2356 19130
rect 2446 19096 2514 19130
rect 2604 19096 2672 19130
rect 2762 19096 2830 19130
rect 2920 19096 2988 19130
rect 3078 19096 3146 19130
rect 3236 19096 3304 19130
rect 3394 19096 3462 19130
rect 3552 19096 3620 19130
rect 3710 19096 3778 19130
rect 3868 19096 3936 19130
rect 4026 19096 4094 19130
rect 5736 19234 10459 19268
rect 5736 19232 10459 19234
rect 5744 19096 5812 19130
rect 5902 19096 5970 19130
rect 6060 19096 6128 19130
rect 6218 19096 6286 19130
rect 6376 19096 6444 19130
rect 6534 19096 6602 19130
rect 6692 19096 6760 19130
rect 6850 19096 6918 19130
rect 7008 19096 7076 19130
rect 7166 19096 7234 19130
rect 7324 19096 7392 19130
rect 7482 19096 7550 19130
rect 7640 19096 7708 19130
rect 7798 19096 7866 19130
rect 7956 19096 8024 19130
rect 8114 19096 8182 19130
rect 8272 19096 8340 19130
rect 8430 19096 8498 19130
rect 8588 19096 8656 19130
rect 8746 19096 8814 19130
rect 8904 19096 8972 19130
rect 9062 19096 9130 19130
rect 9220 19096 9288 19130
rect 9378 19096 9446 19130
rect 9536 19096 9604 19130
rect 9694 19096 9762 19130
rect 9852 19096 9920 19130
rect 10010 19096 10078 19130
rect 10168 19096 10236 19130
rect 10326 19096 10394 19130
rect -13354 13036 -13352 19080
rect -13352 13036 -13318 19080
rect -13318 13036 -13316 19080
rect -13218 13070 -13184 19046
rect -13060 13070 -13026 19046
rect -12902 13070 -12868 19046
rect -12744 13070 -12710 19046
rect -12586 13070 -12552 19046
rect -12428 13070 -12394 19046
rect -12270 13070 -12236 19046
rect -12112 13070 -12078 19046
rect -11954 13070 -11920 19046
rect -11796 13070 -11762 19046
rect -11638 13070 -11604 19046
rect -11480 13070 -11446 19046
rect -11322 13070 -11288 19046
rect -11164 13070 -11130 19046
rect -11006 13070 -10972 19046
rect -10848 13070 -10814 19046
rect -10690 13070 -10656 19046
rect -10532 13070 -10498 19046
rect -10374 13070 -10340 19046
rect -10216 13070 -10182 19046
rect -10058 13070 -10024 19046
rect -9900 13070 -9866 19046
rect -9742 13070 -9708 19046
rect -9584 13070 -9550 19046
rect -9426 13070 -9392 19046
rect -9268 13070 -9234 19046
rect -9110 13070 -9076 19046
rect -8952 13070 -8918 19046
rect -8794 13070 -8760 19046
rect -8636 13070 -8602 19046
rect -8478 13070 -8444 19046
rect -8346 13036 -8344 19080
rect -8344 13036 -8310 19080
rect -8310 13036 -8308 19080
rect -7054 13036 -7052 19080
rect -7052 13036 -7018 19080
rect -7018 13036 -7016 19080
rect -6918 13070 -6884 19046
rect -6760 13070 -6726 19046
rect -6602 13070 -6568 19046
rect -6444 13070 -6410 19046
rect -6286 13070 -6252 19046
rect -6128 13070 -6094 19046
rect -5970 13070 -5936 19046
rect -5812 13070 -5778 19046
rect -5654 13070 -5620 19046
rect -5496 13070 -5462 19046
rect -5338 13070 -5304 19046
rect -5180 13070 -5146 19046
rect -5022 13070 -4988 19046
rect -4864 13070 -4830 19046
rect -4706 13070 -4672 19046
rect -4548 13070 -4514 19046
rect -4390 13070 -4356 19046
rect -4232 13070 -4198 19046
rect -4074 13070 -4040 19046
rect -3916 13070 -3882 19046
rect -3758 13070 -3724 19046
rect -3600 13070 -3566 19046
rect -3442 13070 -3408 19046
rect -3284 13070 -3250 19046
rect -3126 13070 -3092 19046
rect -2968 13070 -2934 19046
rect -2810 13070 -2776 19046
rect -2652 13070 -2618 19046
rect -2494 13070 -2460 19046
rect -2336 13070 -2302 19046
rect -2178 13070 -2144 19046
rect -2046 13036 -2044 19080
rect -2044 13036 -2010 19080
rect -2010 13036 -2008 19080
rect -754 13036 -752 19080
rect -752 13036 -718 19080
rect -718 13036 -716 19080
rect -618 13070 -584 19046
rect -460 13070 -426 19046
rect -302 13070 -268 19046
rect -144 13070 -110 19046
rect 14 13070 48 19046
rect 172 13070 206 19046
rect 330 13070 364 19046
rect 488 13070 522 19046
rect 646 13070 680 19046
rect 804 13070 838 19046
rect 962 13070 996 19046
rect 1120 13070 1154 19046
rect 1278 13070 1312 19046
rect 1436 13070 1470 19046
rect 1594 13070 1628 19046
rect 1752 13070 1786 19046
rect 1910 13070 1944 19046
rect 2068 13070 2102 19046
rect 2226 13070 2260 19046
rect 2384 13070 2418 19046
rect 2542 13070 2576 19046
rect 2700 13070 2734 19046
rect 2858 13070 2892 19046
rect 3016 13070 3050 19046
rect 3174 13070 3208 19046
rect 3332 13070 3366 19046
rect 3490 13070 3524 19046
rect 3648 13070 3682 19046
rect 3806 13070 3840 19046
rect 3964 13070 3998 19046
rect 4122 13070 4156 19046
rect 4254 13036 4256 19080
rect 4256 13036 4290 19080
rect 4290 13036 4292 19080
rect 5546 13036 5548 19080
rect 5548 13036 5582 19080
rect 5582 13036 5584 19080
rect 5682 13070 5716 19046
rect 5840 13070 5874 19046
rect 5998 13070 6032 19046
rect 6156 13070 6190 19046
rect 6314 13070 6348 19046
rect 6472 13070 6506 19046
rect 6630 13070 6664 19046
rect 6788 13070 6822 19046
rect 6946 13070 6980 19046
rect 7104 13070 7138 19046
rect 7262 13070 7296 19046
rect 7420 13070 7454 19046
rect 7578 13070 7612 19046
rect 7736 13070 7770 19046
rect 7894 13070 7928 19046
rect 8052 13070 8086 19046
rect 8210 13070 8244 19046
rect 8368 13070 8402 19046
rect 8526 13070 8560 19046
rect 8684 13070 8718 19046
rect 8842 13070 8876 19046
rect 9000 13070 9034 19046
rect 9158 13070 9192 19046
rect 9316 13070 9350 19046
rect 9474 13070 9508 19046
rect 9632 13070 9666 19046
rect 9790 13070 9824 19046
rect 9948 13070 9982 19046
rect 10106 13070 10140 19046
rect 10264 13070 10298 19046
rect 10422 13070 10456 19046
rect 10554 13036 10556 19080
rect 10556 13036 10590 19080
rect 10590 13036 10592 19080
rect -13156 12986 -13088 13020
rect -12998 12986 -12930 13020
rect -12840 12986 -12772 13020
rect -12682 12986 -12614 13020
rect -12524 12986 -12456 13020
rect -12366 12986 -12298 13020
rect -12208 12986 -12140 13020
rect -12050 12986 -11982 13020
rect -11892 12986 -11824 13020
rect -11734 12986 -11666 13020
rect -11576 12986 -11508 13020
rect -11418 12986 -11350 13020
rect -11260 12986 -11192 13020
rect -11102 12986 -11034 13020
rect -10944 12986 -10876 13020
rect -10786 12986 -10718 13020
rect -10628 12986 -10560 13020
rect -10470 12986 -10402 13020
rect -10312 12986 -10244 13020
rect -10154 12986 -10086 13020
rect -9996 12986 -9928 13020
rect -9838 12986 -9770 13020
rect -9680 12986 -9612 13020
rect -9522 12986 -9454 13020
rect -9364 12986 -9296 13020
rect -9206 12986 -9138 13020
rect -9048 12986 -8980 13020
rect -8890 12986 -8822 13020
rect -8732 12986 -8664 13020
rect -8574 12986 -8506 13020
rect -13164 12882 -8498 12884
rect -13164 12848 -8498 12882
rect -6856 12986 -6788 13020
rect -6698 12986 -6630 13020
rect -6540 12986 -6472 13020
rect -6382 12986 -6314 13020
rect -6224 12986 -6156 13020
rect -6066 12986 -5998 13020
rect -5908 12986 -5840 13020
rect -5750 12986 -5682 13020
rect -5592 12986 -5524 13020
rect -5434 12986 -5366 13020
rect -5276 12986 -5208 13020
rect -5118 12986 -5050 13020
rect -4960 12986 -4892 13020
rect -4802 12986 -4734 13020
rect -4644 12986 -4576 13020
rect -4486 12986 -4418 13020
rect -4328 12986 -4260 13020
rect -4170 12986 -4102 13020
rect -4012 12986 -3944 13020
rect -3854 12986 -3786 13020
rect -3696 12986 -3628 13020
rect -3538 12986 -3470 13020
rect -3380 12986 -3312 13020
rect -3222 12986 -3154 13020
rect -3064 12986 -2996 13020
rect -2906 12986 -2838 13020
rect -2748 12986 -2680 13020
rect -2590 12986 -2522 13020
rect -2432 12986 -2364 13020
rect -2274 12986 -2206 13020
rect -6864 12882 -2198 12884
rect -6864 12848 -2198 12882
rect -556 12986 -488 13020
rect -398 12986 -330 13020
rect -240 12986 -172 13020
rect -82 12986 -14 13020
rect 76 12986 144 13020
rect 234 12986 302 13020
rect 392 12986 460 13020
rect 550 12986 618 13020
rect 708 12986 776 13020
rect 866 12986 934 13020
rect 1024 12986 1092 13020
rect 1182 12986 1250 13020
rect 1340 12986 1408 13020
rect 1498 12986 1566 13020
rect 1656 12986 1724 13020
rect 1814 12986 1882 13020
rect 1972 12986 2040 13020
rect 2130 12986 2198 13020
rect 2288 12986 2356 13020
rect 2446 12986 2514 13020
rect 2604 12986 2672 13020
rect 2762 12986 2830 13020
rect 2920 12986 2988 13020
rect 3078 12986 3146 13020
rect 3236 12986 3304 13020
rect 3394 12986 3462 13020
rect 3552 12986 3620 13020
rect 3710 12986 3778 13020
rect 3868 12986 3936 13020
rect 4026 12986 4094 13020
rect -564 12882 4102 12884
rect -564 12848 4102 12882
rect 5744 12986 5812 13020
rect 5902 12986 5970 13020
rect 6060 12986 6128 13020
rect 6218 12986 6286 13020
rect 6376 12986 6444 13020
rect 6534 12986 6602 13020
rect 6692 12986 6760 13020
rect 6850 12986 6918 13020
rect 7008 12986 7076 13020
rect 7166 12986 7234 13020
rect 7324 12986 7392 13020
rect 7482 12986 7550 13020
rect 7640 12986 7708 13020
rect 7798 12986 7866 13020
rect 7956 12986 8024 13020
rect 8114 12986 8182 13020
rect 8272 12986 8340 13020
rect 8430 12986 8498 13020
rect 8588 12986 8656 13020
rect 8746 12986 8814 13020
rect 8904 12986 8972 13020
rect 9062 12986 9130 13020
rect 9220 12986 9288 13020
rect 9378 12986 9446 13020
rect 9536 12986 9604 13020
rect 9694 12986 9762 13020
rect 9852 12986 9920 13020
rect 10010 12986 10078 13020
rect 10168 12986 10236 13020
rect 10326 12986 10394 13020
rect 5736 12882 10402 12884
rect 5736 12848 10402 12882
rect -13164 12846 -8498 12848
rect -6864 12846 -2198 12848
rect -564 12846 4102 12848
rect 5736 12846 10402 12848
rect -13164 12268 -8441 12270
rect -6864 12268 -2141 12270
rect -564 12268 4159 12270
rect 5736 12268 10459 12270
rect -13164 12234 -8441 12268
rect -13164 12232 -8441 12234
rect -13156 12096 -13088 12130
rect -12998 12096 -12930 12130
rect -12840 12096 -12772 12130
rect -12682 12096 -12614 12130
rect -12524 12096 -12456 12130
rect -12366 12096 -12298 12130
rect -12208 12096 -12140 12130
rect -12050 12096 -11982 12130
rect -11892 12096 -11824 12130
rect -11734 12096 -11666 12130
rect -11576 12096 -11508 12130
rect -11418 12096 -11350 12130
rect -11260 12096 -11192 12130
rect -11102 12096 -11034 12130
rect -10944 12096 -10876 12130
rect -10786 12096 -10718 12130
rect -10628 12096 -10560 12130
rect -10470 12096 -10402 12130
rect -10312 12096 -10244 12130
rect -10154 12096 -10086 12130
rect -9996 12096 -9928 12130
rect -9838 12096 -9770 12130
rect -9680 12096 -9612 12130
rect -9522 12096 -9454 12130
rect -9364 12096 -9296 12130
rect -9206 12096 -9138 12130
rect -9048 12096 -8980 12130
rect -8890 12096 -8822 12130
rect -8732 12096 -8664 12130
rect -8574 12096 -8506 12130
rect -6864 12234 -2141 12268
rect -6864 12232 -2141 12234
rect -6856 12096 -6788 12130
rect -6698 12096 -6630 12130
rect -6540 12096 -6472 12130
rect -6382 12096 -6314 12130
rect -6224 12096 -6156 12130
rect -6066 12096 -5998 12130
rect -5908 12096 -5840 12130
rect -5750 12096 -5682 12130
rect -5592 12096 -5524 12130
rect -5434 12096 -5366 12130
rect -5276 12096 -5208 12130
rect -5118 12096 -5050 12130
rect -4960 12096 -4892 12130
rect -4802 12096 -4734 12130
rect -4644 12096 -4576 12130
rect -4486 12096 -4418 12130
rect -4328 12096 -4260 12130
rect -4170 12096 -4102 12130
rect -4012 12096 -3944 12130
rect -3854 12096 -3786 12130
rect -3696 12096 -3628 12130
rect -3538 12096 -3470 12130
rect -3380 12096 -3312 12130
rect -3222 12096 -3154 12130
rect -3064 12096 -2996 12130
rect -2906 12096 -2838 12130
rect -2748 12096 -2680 12130
rect -2590 12096 -2522 12130
rect -2432 12096 -2364 12130
rect -2274 12096 -2206 12130
rect -564 12234 4159 12268
rect -564 12232 4159 12234
rect -556 12096 -488 12130
rect -398 12096 -330 12130
rect -240 12096 -172 12130
rect -82 12096 -14 12130
rect 76 12096 144 12130
rect 234 12096 302 12130
rect 392 12096 460 12130
rect 550 12096 618 12130
rect 708 12096 776 12130
rect 866 12096 934 12130
rect 1024 12096 1092 12130
rect 1182 12096 1250 12130
rect 1340 12096 1408 12130
rect 1498 12096 1566 12130
rect 1656 12096 1724 12130
rect 1814 12096 1882 12130
rect 1972 12096 2040 12130
rect 2130 12096 2198 12130
rect 2288 12096 2356 12130
rect 2446 12096 2514 12130
rect 2604 12096 2672 12130
rect 2762 12096 2830 12130
rect 2920 12096 2988 12130
rect 3078 12096 3146 12130
rect 3236 12096 3304 12130
rect 3394 12096 3462 12130
rect 3552 12096 3620 12130
rect 3710 12096 3778 12130
rect 3868 12096 3936 12130
rect 4026 12096 4094 12130
rect 5736 12234 10459 12268
rect 5736 12232 10459 12234
rect 5744 12096 5812 12130
rect 5902 12096 5970 12130
rect 6060 12096 6128 12130
rect 6218 12096 6286 12130
rect 6376 12096 6444 12130
rect 6534 12096 6602 12130
rect 6692 12096 6760 12130
rect 6850 12096 6918 12130
rect 7008 12096 7076 12130
rect 7166 12096 7234 12130
rect 7324 12096 7392 12130
rect 7482 12096 7550 12130
rect 7640 12096 7708 12130
rect 7798 12096 7866 12130
rect 7956 12096 8024 12130
rect 8114 12096 8182 12130
rect 8272 12096 8340 12130
rect 8430 12096 8498 12130
rect 8588 12096 8656 12130
rect 8746 12096 8814 12130
rect 8904 12096 8972 12130
rect 9062 12096 9130 12130
rect 9220 12096 9288 12130
rect 9378 12096 9446 12130
rect 9536 12096 9604 12130
rect 9694 12096 9762 12130
rect 9852 12096 9920 12130
rect 10010 12096 10078 12130
rect 10168 12096 10236 12130
rect 10326 12096 10394 12130
rect -13354 6036 -13352 12080
rect -13352 6036 -13318 12080
rect -13318 6036 -13316 12080
rect -13218 6070 -13184 12046
rect -13060 6070 -13026 12046
rect -12902 6070 -12868 12046
rect -12744 6070 -12710 12046
rect -12586 6070 -12552 12046
rect -12428 6070 -12394 12046
rect -12270 6070 -12236 12046
rect -12112 6070 -12078 12046
rect -11954 6070 -11920 12046
rect -11796 6070 -11762 12046
rect -11638 6070 -11604 12046
rect -11480 6070 -11446 12046
rect -11322 6070 -11288 12046
rect -11164 6070 -11130 12046
rect -11006 6070 -10972 12046
rect -10848 6070 -10814 12046
rect -10690 6070 -10656 12046
rect -10532 6070 -10498 12046
rect -10374 6070 -10340 12046
rect -10216 6070 -10182 12046
rect -10058 6070 -10024 12046
rect -9900 6070 -9866 12046
rect -9742 6070 -9708 12046
rect -9584 6070 -9550 12046
rect -9426 6070 -9392 12046
rect -9268 6070 -9234 12046
rect -9110 6070 -9076 12046
rect -8952 6070 -8918 12046
rect -8794 6070 -8760 12046
rect -8636 6070 -8602 12046
rect -8478 6070 -8444 12046
rect -8346 6036 -8344 12080
rect -8344 6036 -8310 12080
rect -8310 6036 -8308 12080
rect -7054 6036 -7052 12080
rect -7052 6036 -7018 12080
rect -7018 6036 -7016 12080
rect -6918 6070 -6884 12046
rect -6760 6070 -6726 12046
rect -6602 6070 -6568 12046
rect -6444 6070 -6410 12046
rect -6286 6070 -6252 12046
rect -6128 6070 -6094 12046
rect -5970 6070 -5936 12046
rect -5812 6070 -5778 12046
rect -5654 6070 -5620 12046
rect -5496 6070 -5462 12046
rect -5338 6070 -5304 12046
rect -5180 6070 -5146 12046
rect -5022 6070 -4988 12046
rect -4864 6070 -4830 12046
rect -4706 6070 -4672 12046
rect -4548 6070 -4514 12046
rect -4390 6070 -4356 12046
rect -4232 6070 -4198 12046
rect -4074 6070 -4040 12046
rect -3916 6070 -3882 12046
rect -3758 6070 -3724 12046
rect -3600 6070 -3566 12046
rect -3442 6070 -3408 12046
rect -3284 6070 -3250 12046
rect -3126 6070 -3092 12046
rect -2968 6070 -2934 12046
rect -2810 6070 -2776 12046
rect -2652 6070 -2618 12046
rect -2494 6070 -2460 12046
rect -2336 6070 -2302 12046
rect -2178 6070 -2144 12046
rect -2046 6036 -2044 12080
rect -2044 6036 -2010 12080
rect -2010 6036 -2008 12080
rect -754 6036 -752 12080
rect -752 6036 -718 12080
rect -718 6036 -716 12080
rect -618 6070 -584 12046
rect -460 6070 -426 12046
rect -302 6070 -268 12046
rect -144 6070 -110 12046
rect 14 6070 48 12046
rect 172 6070 206 12046
rect 330 6070 364 12046
rect 488 6070 522 12046
rect 646 6070 680 12046
rect 804 6070 838 12046
rect 962 6070 996 12046
rect 1120 6070 1154 12046
rect 1278 6070 1312 12046
rect 1436 6070 1470 12046
rect 1594 6070 1628 12046
rect 1752 6070 1786 12046
rect 1910 6070 1944 12046
rect 2068 6070 2102 12046
rect 2226 6070 2260 12046
rect 2384 6070 2418 12046
rect 2542 6070 2576 12046
rect 2700 6070 2734 12046
rect 2858 6070 2892 12046
rect 3016 6070 3050 12046
rect 3174 6070 3208 12046
rect 3332 6070 3366 12046
rect 3490 6070 3524 12046
rect 3648 6070 3682 12046
rect 3806 6070 3840 12046
rect 3964 6070 3998 12046
rect 4122 6070 4156 12046
rect 4254 6036 4256 12080
rect 4256 6036 4290 12080
rect 4290 6036 4292 12080
rect 5546 6036 5548 12080
rect 5548 6036 5582 12080
rect 5582 6036 5584 12080
rect 5682 6070 5716 12046
rect 5840 6070 5874 12046
rect 5998 6070 6032 12046
rect 6156 6070 6190 12046
rect 6314 6070 6348 12046
rect 6472 6070 6506 12046
rect 6630 6070 6664 12046
rect 6788 6070 6822 12046
rect 6946 6070 6980 12046
rect 7104 6070 7138 12046
rect 7262 6070 7296 12046
rect 7420 6070 7454 12046
rect 7578 6070 7612 12046
rect 7736 6070 7770 12046
rect 7894 6070 7928 12046
rect 8052 6070 8086 12046
rect 8210 6070 8244 12046
rect 8368 6070 8402 12046
rect 8526 6070 8560 12046
rect 8684 6070 8718 12046
rect 8842 6070 8876 12046
rect 9000 6070 9034 12046
rect 9158 6070 9192 12046
rect 9316 6070 9350 12046
rect 9474 6070 9508 12046
rect 9632 6070 9666 12046
rect 9790 6070 9824 12046
rect 9948 6070 9982 12046
rect 10106 6070 10140 12046
rect 10264 6070 10298 12046
rect 10422 6070 10456 12046
rect 10554 6036 10556 12080
rect 10556 6036 10590 12080
rect 10590 6036 10592 12080
rect -13156 5986 -13088 6020
rect -12998 5986 -12930 6020
rect -12840 5986 -12772 6020
rect -12682 5986 -12614 6020
rect -12524 5986 -12456 6020
rect -12366 5986 -12298 6020
rect -12208 5986 -12140 6020
rect -12050 5986 -11982 6020
rect -11892 5986 -11824 6020
rect -11734 5986 -11666 6020
rect -11576 5986 -11508 6020
rect -11418 5986 -11350 6020
rect -11260 5986 -11192 6020
rect -11102 5986 -11034 6020
rect -10944 5986 -10876 6020
rect -10786 5986 -10718 6020
rect -10628 5986 -10560 6020
rect -10470 5986 -10402 6020
rect -10312 5986 -10244 6020
rect -10154 5986 -10086 6020
rect -9996 5986 -9928 6020
rect -9838 5986 -9770 6020
rect -9680 5986 -9612 6020
rect -9522 5986 -9454 6020
rect -9364 5986 -9296 6020
rect -9206 5986 -9138 6020
rect -9048 5986 -8980 6020
rect -8890 5986 -8822 6020
rect -8732 5986 -8664 6020
rect -8574 5986 -8506 6020
rect -13164 5882 -8498 5884
rect -13164 5848 -8498 5882
rect -6856 5986 -6788 6020
rect -6698 5986 -6630 6020
rect -6540 5986 -6472 6020
rect -6382 5986 -6314 6020
rect -6224 5986 -6156 6020
rect -6066 5986 -5998 6020
rect -5908 5986 -5840 6020
rect -5750 5986 -5682 6020
rect -5592 5986 -5524 6020
rect -5434 5986 -5366 6020
rect -5276 5986 -5208 6020
rect -5118 5986 -5050 6020
rect -4960 5986 -4892 6020
rect -4802 5986 -4734 6020
rect -4644 5986 -4576 6020
rect -4486 5986 -4418 6020
rect -4328 5986 -4260 6020
rect -4170 5986 -4102 6020
rect -4012 5986 -3944 6020
rect -3854 5986 -3786 6020
rect -3696 5986 -3628 6020
rect -3538 5986 -3470 6020
rect -3380 5986 -3312 6020
rect -3222 5986 -3154 6020
rect -3064 5986 -2996 6020
rect -2906 5986 -2838 6020
rect -2748 5986 -2680 6020
rect -2590 5986 -2522 6020
rect -2432 5986 -2364 6020
rect -2274 5986 -2206 6020
rect -6864 5882 -2198 5884
rect -6864 5848 -2198 5882
rect -556 5986 -488 6020
rect -398 5986 -330 6020
rect -240 5986 -172 6020
rect -82 5986 -14 6020
rect 76 5986 144 6020
rect 234 5986 302 6020
rect 392 5986 460 6020
rect 550 5986 618 6020
rect 708 5986 776 6020
rect 866 5986 934 6020
rect 1024 5986 1092 6020
rect 1182 5986 1250 6020
rect 1340 5986 1408 6020
rect 1498 5986 1566 6020
rect 1656 5986 1724 6020
rect 1814 5986 1882 6020
rect 1972 5986 2040 6020
rect 2130 5986 2198 6020
rect 2288 5986 2356 6020
rect 2446 5986 2514 6020
rect 2604 5986 2672 6020
rect 2762 5986 2830 6020
rect 2920 5986 2988 6020
rect 3078 5986 3146 6020
rect 3236 5986 3304 6020
rect 3394 5986 3462 6020
rect 3552 5986 3620 6020
rect 3710 5986 3778 6020
rect 3868 5986 3936 6020
rect 4026 5986 4094 6020
rect -564 5882 4102 5884
rect -564 5848 4102 5882
rect 5744 5986 5812 6020
rect 5902 5986 5970 6020
rect 6060 5986 6128 6020
rect 6218 5986 6286 6020
rect 6376 5986 6444 6020
rect 6534 5986 6602 6020
rect 6692 5986 6760 6020
rect 6850 5986 6918 6020
rect 7008 5986 7076 6020
rect 7166 5986 7234 6020
rect 7324 5986 7392 6020
rect 7482 5986 7550 6020
rect 7640 5986 7708 6020
rect 7798 5986 7866 6020
rect 7956 5986 8024 6020
rect 8114 5986 8182 6020
rect 8272 5986 8340 6020
rect 8430 5986 8498 6020
rect 8588 5986 8656 6020
rect 8746 5986 8814 6020
rect 8904 5986 8972 6020
rect 9062 5986 9130 6020
rect 9220 5986 9288 6020
rect 9378 5986 9446 6020
rect 9536 5986 9604 6020
rect 9694 5986 9762 6020
rect 9852 5986 9920 6020
rect 10010 5986 10078 6020
rect 10168 5986 10236 6020
rect 10326 5986 10394 6020
rect 5736 5882 10402 5884
rect 5736 5848 10402 5882
rect -13164 5846 -8498 5848
rect -6864 5846 -2198 5848
rect -564 5846 4102 5848
rect 5736 5846 10402 5848
<< metal1 >>
rect -13370 49870 -8290 49880
rect -13370 49832 -13164 49870
rect -8441 49832 -8290 49870
rect -13370 49822 -8290 49832
rect -13370 49820 -13300 49822
rect -8360 49820 -8290 49822
rect -13168 49730 -13148 49790
rect -8514 49730 -8494 49790
rect -13168 49696 -13156 49730
rect -8506 49696 -8494 49730
rect -13168 49690 -13148 49696
rect -8514 49690 -8494 49696
rect -13235 49646 -13169 49658
rect -13235 49638 -13218 49646
rect -13184 49638 -13169 49646
rect -13235 43670 -13218 43678
rect -13184 43670 -13169 43678
rect -13235 43658 -13169 43670
rect -13077 49646 -13011 49658
rect -13077 49638 -13060 49646
rect -13026 49638 -13011 49646
rect -13077 43670 -13060 43678
rect -13026 43670 -13011 43678
rect -13077 43658 -13011 43670
rect -12919 49646 -12853 49658
rect -12919 49638 -12902 49646
rect -12868 49638 -12853 49646
rect -12919 43670 -12902 43678
rect -12868 43670 -12853 43678
rect -12919 43658 -12853 43670
rect -12761 49646 -12695 49658
rect -12761 49638 -12744 49646
rect -12710 49638 -12695 49646
rect -12761 43670 -12744 43678
rect -12710 43670 -12695 43678
rect -12761 43658 -12695 43670
rect -12603 49646 -12537 49658
rect -12603 49638 -12586 49646
rect -12552 49638 -12537 49646
rect -12603 43670 -12586 43678
rect -12552 43670 -12537 43678
rect -12603 43658 -12537 43670
rect -12445 49646 -12379 49658
rect -12445 49638 -12428 49646
rect -12394 49638 -12379 49646
rect -12445 43670 -12428 43678
rect -12394 43670 -12379 43678
rect -12445 43658 -12379 43670
rect -12287 49646 -12221 49658
rect -12287 49638 -12270 49646
rect -12236 49638 -12221 49646
rect -12287 43670 -12270 43678
rect -12236 43670 -12221 43678
rect -12287 43658 -12221 43670
rect -12129 49646 -12063 49658
rect -12129 49638 -12112 49646
rect -12078 49638 -12063 49646
rect -12129 43670 -12112 43678
rect -12078 43670 -12063 43678
rect -12129 43658 -12063 43670
rect -11971 49646 -11905 49658
rect -11971 49638 -11954 49646
rect -11920 49638 -11905 49646
rect -11971 43670 -11954 43678
rect -11920 43670 -11905 43678
rect -11971 43658 -11905 43670
rect -11813 49646 -11747 49658
rect -11813 49638 -11796 49646
rect -11762 49638 -11747 49646
rect -11813 43670 -11796 43678
rect -11762 43670 -11747 43678
rect -11813 43658 -11747 43670
rect -11655 49646 -11589 49658
rect -11655 49638 -11638 49646
rect -11604 49638 -11589 49646
rect -11655 43670 -11638 43678
rect -11604 43670 -11589 43678
rect -11655 43658 -11589 43670
rect -11497 49646 -11431 49658
rect -11497 49638 -11480 49646
rect -11446 49638 -11431 49646
rect -11497 43670 -11480 43678
rect -11446 43670 -11431 43678
rect -11497 43658 -11431 43670
rect -11339 49646 -11273 49658
rect -11339 49638 -11322 49646
rect -11288 49638 -11273 49646
rect -11339 43670 -11322 43678
rect -11288 43670 -11273 43678
rect -11339 43658 -11273 43670
rect -11181 49646 -11115 49658
rect -11181 49638 -11164 49646
rect -11130 49638 -11115 49646
rect -11181 43670 -11164 43678
rect -11130 43670 -11115 43678
rect -11181 43658 -11115 43670
rect -11023 49646 -10957 49658
rect -11023 49638 -11006 49646
rect -10972 49638 -10957 49646
rect -11023 43670 -11006 43678
rect -10972 43670 -10957 43678
rect -11023 43658 -10957 43670
rect -10865 49646 -10799 49658
rect -10865 49638 -10848 49646
rect -10814 49638 -10799 49646
rect -10865 43670 -10848 43678
rect -10814 43670 -10799 43678
rect -10865 43658 -10799 43670
rect -10707 49646 -10641 49658
rect -10707 49638 -10690 49646
rect -10656 49638 -10641 49646
rect -10707 43670 -10690 43678
rect -10656 43670 -10641 43678
rect -10707 43658 -10641 43670
rect -10549 49646 -10483 49658
rect -10549 49638 -10532 49646
rect -10498 49638 -10483 49646
rect -10549 43670 -10532 43678
rect -10498 43670 -10483 43678
rect -10549 43658 -10483 43670
rect -10391 49646 -10325 49658
rect -10391 49638 -10374 49646
rect -10340 49638 -10325 49646
rect -10391 43670 -10374 43678
rect -10340 43670 -10325 43678
rect -10391 43658 -10325 43670
rect -10233 49646 -10167 49658
rect -10233 49638 -10216 49646
rect -10182 49638 -10167 49646
rect -10233 43670 -10216 43678
rect -10182 43670 -10167 43678
rect -10233 43658 -10167 43670
rect -10075 49646 -10009 49658
rect -10075 49638 -10058 49646
rect -10024 49638 -10009 49646
rect -10075 43670 -10058 43678
rect -10024 43670 -10009 43678
rect -10075 43658 -10009 43670
rect -9917 49646 -9851 49658
rect -9917 49638 -9900 49646
rect -9866 49638 -9851 49646
rect -9917 43670 -9900 43678
rect -9866 43670 -9851 43678
rect -9917 43658 -9851 43670
rect -9759 49646 -9693 49658
rect -9759 49638 -9742 49646
rect -9708 49638 -9693 49646
rect -9759 43670 -9742 43678
rect -9708 43670 -9693 43678
rect -9759 43658 -9693 43670
rect -9601 49646 -9535 49658
rect -9601 49638 -9584 49646
rect -9550 49638 -9535 49646
rect -9601 43670 -9584 43678
rect -9550 43670 -9535 43678
rect -9601 43658 -9535 43670
rect -9443 49646 -9377 49658
rect -9443 49638 -9426 49646
rect -9392 49638 -9377 49646
rect -9443 43670 -9426 43678
rect -9392 43670 -9377 43678
rect -9443 43658 -9377 43670
rect -9285 49646 -9219 49658
rect -9285 49638 -9268 49646
rect -9234 49638 -9219 49646
rect -9285 43670 -9268 43678
rect -9234 43670 -9219 43678
rect -9285 43658 -9219 43670
rect -9127 49646 -9061 49658
rect -9127 49638 -9110 49646
rect -9076 49638 -9061 49646
rect -9127 43670 -9110 43678
rect -9076 43670 -9061 43678
rect -9127 43658 -9061 43670
rect -8969 49646 -8903 49658
rect -8969 49638 -8952 49646
rect -8918 49638 -8903 49646
rect -8969 43670 -8952 43678
rect -8918 43670 -8903 43678
rect -8969 43658 -8903 43670
rect -8811 49646 -8745 49658
rect -8811 49638 -8794 49646
rect -8760 49638 -8745 49646
rect -8811 43670 -8794 43678
rect -8760 43670 -8745 43678
rect -8811 43658 -8745 43670
rect -8653 49646 -8587 49658
rect -8653 49638 -8636 49646
rect -8602 49638 -8587 49646
rect -8653 43670 -8636 43678
rect -8602 43670 -8587 43678
rect -8653 43658 -8587 43670
rect -8495 49646 -8429 49658
rect -8495 49638 -8478 49646
rect -8444 49638 -8429 49646
rect -8495 43670 -8478 43678
rect -8444 43670 -8429 43678
rect -8495 43658 -8429 43670
rect -13168 43620 -13148 43626
rect -8514 43620 -8494 43626
rect -13168 43586 -13156 43620
rect -8506 43586 -8494 43620
rect -13168 43526 -13148 43586
rect -8514 43526 -8494 43586
rect -13370 43494 -13300 43500
rect -8360 43494 -8290 43500
rect -13370 43484 -8290 43494
rect -13370 43446 -13164 43484
rect -8498 43446 -8290 43484
rect -13370 43430 -8290 43446
rect -7070 49870 -1990 49880
rect -7070 49832 -6864 49870
rect -2141 49832 -1990 49870
rect -7070 49822 -1990 49832
rect -7070 49820 -7000 49822
rect -2060 49820 -1990 49822
rect -6868 49730 -6848 49790
rect -2214 49730 -2194 49790
rect -6868 49696 -6856 49730
rect -2206 49696 -2194 49730
rect -6868 49690 -6848 49696
rect -2214 49690 -2194 49696
rect -6935 49646 -6869 49658
rect -6935 49638 -6918 49646
rect -6884 49638 -6869 49646
rect -6935 43670 -6918 43678
rect -6884 43670 -6869 43678
rect -6935 43658 -6869 43670
rect -6777 49646 -6711 49658
rect -6777 49638 -6760 49646
rect -6726 49638 -6711 49646
rect -6777 43670 -6760 43678
rect -6726 43670 -6711 43678
rect -6777 43658 -6711 43670
rect -6619 49646 -6553 49658
rect -6619 49638 -6602 49646
rect -6568 49638 -6553 49646
rect -6619 43670 -6602 43678
rect -6568 43670 -6553 43678
rect -6619 43658 -6553 43670
rect -6461 49646 -6395 49658
rect -6461 49638 -6444 49646
rect -6410 49638 -6395 49646
rect -6461 43670 -6444 43678
rect -6410 43670 -6395 43678
rect -6461 43658 -6395 43670
rect -6303 49646 -6237 49658
rect -6303 49638 -6286 49646
rect -6252 49638 -6237 49646
rect -6303 43670 -6286 43678
rect -6252 43670 -6237 43678
rect -6303 43658 -6237 43670
rect -6145 49646 -6079 49658
rect -6145 49638 -6128 49646
rect -6094 49638 -6079 49646
rect -6145 43670 -6128 43678
rect -6094 43670 -6079 43678
rect -6145 43658 -6079 43670
rect -5987 49646 -5921 49658
rect -5987 49638 -5970 49646
rect -5936 49638 -5921 49646
rect -5987 43670 -5970 43678
rect -5936 43670 -5921 43678
rect -5987 43658 -5921 43670
rect -5829 49646 -5763 49658
rect -5829 49638 -5812 49646
rect -5778 49638 -5763 49646
rect -5829 43670 -5812 43678
rect -5778 43670 -5763 43678
rect -5829 43658 -5763 43670
rect -5671 49646 -5605 49658
rect -5671 49638 -5654 49646
rect -5620 49638 -5605 49646
rect -5671 43670 -5654 43678
rect -5620 43670 -5605 43678
rect -5671 43658 -5605 43670
rect -5513 49646 -5447 49658
rect -5513 49638 -5496 49646
rect -5462 49638 -5447 49646
rect -5513 43670 -5496 43678
rect -5462 43670 -5447 43678
rect -5513 43658 -5447 43670
rect -5355 49646 -5289 49658
rect -5355 49638 -5338 49646
rect -5304 49638 -5289 49646
rect -5355 43670 -5338 43678
rect -5304 43670 -5289 43678
rect -5355 43658 -5289 43670
rect -5197 49646 -5131 49658
rect -5197 49638 -5180 49646
rect -5146 49638 -5131 49646
rect -5197 43670 -5180 43678
rect -5146 43670 -5131 43678
rect -5197 43658 -5131 43670
rect -5039 49646 -4973 49658
rect -5039 49638 -5022 49646
rect -4988 49638 -4973 49646
rect -5039 43670 -5022 43678
rect -4988 43670 -4973 43678
rect -5039 43658 -4973 43670
rect -4881 49646 -4815 49658
rect -4881 49638 -4864 49646
rect -4830 49638 -4815 49646
rect -4881 43670 -4864 43678
rect -4830 43670 -4815 43678
rect -4881 43658 -4815 43670
rect -4723 49646 -4657 49658
rect -4723 49638 -4706 49646
rect -4672 49638 -4657 49646
rect -4723 43670 -4706 43678
rect -4672 43670 -4657 43678
rect -4723 43658 -4657 43670
rect -4565 49646 -4499 49658
rect -4565 49638 -4548 49646
rect -4514 49638 -4499 49646
rect -4565 43670 -4548 43678
rect -4514 43670 -4499 43678
rect -4565 43658 -4499 43670
rect -4407 49646 -4341 49658
rect -4407 49638 -4390 49646
rect -4356 49638 -4341 49646
rect -4407 43670 -4390 43678
rect -4356 43670 -4341 43678
rect -4407 43658 -4341 43670
rect -4249 49646 -4183 49658
rect -4249 49638 -4232 49646
rect -4198 49638 -4183 49646
rect -4249 43670 -4232 43678
rect -4198 43670 -4183 43678
rect -4249 43658 -4183 43670
rect -4091 49646 -4025 49658
rect -4091 49638 -4074 49646
rect -4040 49638 -4025 49646
rect -4091 43670 -4074 43678
rect -4040 43670 -4025 43678
rect -4091 43658 -4025 43670
rect -3933 49646 -3867 49658
rect -3933 49638 -3916 49646
rect -3882 49638 -3867 49646
rect -3933 43670 -3916 43678
rect -3882 43670 -3867 43678
rect -3933 43658 -3867 43670
rect -3775 49646 -3709 49658
rect -3775 49638 -3758 49646
rect -3724 49638 -3709 49646
rect -3775 43670 -3758 43678
rect -3724 43670 -3709 43678
rect -3775 43658 -3709 43670
rect -3617 49646 -3551 49658
rect -3617 49638 -3600 49646
rect -3566 49638 -3551 49646
rect -3617 43670 -3600 43678
rect -3566 43670 -3551 43678
rect -3617 43658 -3551 43670
rect -3459 49646 -3393 49658
rect -3459 49638 -3442 49646
rect -3408 49638 -3393 49646
rect -3459 43670 -3442 43678
rect -3408 43670 -3393 43678
rect -3459 43658 -3393 43670
rect -3301 49646 -3235 49658
rect -3301 49638 -3284 49646
rect -3250 49638 -3235 49646
rect -3301 43670 -3284 43678
rect -3250 43670 -3235 43678
rect -3301 43658 -3235 43670
rect -3143 49646 -3077 49658
rect -3143 49638 -3126 49646
rect -3092 49638 -3077 49646
rect -3143 43670 -3126 43678
rect -3092 43670 -3077 43678
rect -3143 43658 -3077 43670
rect -2985 49646 -2919 49658
rect -2985 49638 -2968 49646
rect -2934 49638 -2919 49646
rect -2985 43670 -2968 43678
rect -2934 43670 -2919 43678
rect -2985 43658 -2919 43670
rect -2827 49646 -2761 49658
rect -2827 49638 -2810 49646
rect -2776 49638 -2761 49646
rect -2827 43670 -2810 43678
rect -2776 43670 -2761 43678
rect -2827 43658 -2761 43670
rect -2669 49646 -2603 49658
rect -2669 49638 -2652 49646
rect -2618 49638 -2603 49646
rect -2669 43670 -2652 43678
rect -2618 43670 -2603 43678
rect -2669 43658 -2603 43670
rect -2511 49646 -2445 49658
rect -2511 49638 -2494 49646
rect -2460 49638 -2445 49646
rect -2511 43670 -2494 43678
rect -2460 43670 -2445 43678
rect -2511 43658 -2445 43670
rect -2353 49646 -2287 49658
rect -2353 49638 -2336 49646
rect -2302 49638 -2287 49646
rect -2353 43670 -2336 43678
rect -2302 43670 -2287 43678
rect -2353 43658 -2287 43670
rect -2195 49646 -2129 49658
rect -2195 49638 -2178 49646
rect -2144 49638 -2129 49646
rect -2195 43670 -2178 43678
rect -2144 43670 -2129 43678
rect -2195 43658 -2129 43670
rect -6868 43620 -6848 43626
rect -2214 43620 -2194 43626
rect -6868 43586 -6856 43620
rect -2206 43586 -2194 43620
rect -6868 43526 -6848 43586
rect -2214 43526 -2194 43586
rect -7070 43494 -7000 43500
rect -2060 43494 -1990 43500
rect -7070 43484 -1990 43494
rect -7070 43446 -6864 43484
rect -2198 43446 -1990 43484
rect -7070 43430 -1990 43446
rect -770 49870 4310 49880
rect -770 49832 -564 49870
rect 4159 49832 4310 49870
rect -770 49822 4310 49832
rect -770 49820 -700 49822
rect 4240 49820 4310 49822
rect -568 49730 -548 49790
rect 4086 49730 4106 49790
rect -568 49696 -556 49730
rect 4094 49696 4106 49730
rect -568 49690 -548 49696
rect 4086 49690 4106 49696
rect -635 49646 -569 49658
rect -635 49638 -618 49646
rect -584 49638 -569 49646
rect -635 43670 -618 43678
rect -584 43670 -569 43678
rect -635 43658 -569 43670
rect -477 49646 -411 49658
rect -477 49638 -460 49646
rect -426 49638 -411 49646
rect -477 43670 -460 43678
rect -426 43670 -411 43678
rect -477 43658 -411 43670
rect -319 49646 -253 49658
rect -319 49638 -302 49646
rect -268 49638 -253 49646
rect -319 43670 -302 43678
rect -268 43670 -253 43678
rect -319 43658 -253 43670
rect -161 49646 -95 49658
rect -161 49638 -144 49646
rect -110 49638 -95 49646
rect -161 43670 -144 43678
rect -110 43670 -95 43678
rect -161 43658 -95 43670
rect -3 49646 63 49658
rect -3 49638 14 49646
rect 48 49638 63 49646
rect -3 43670 14 43678
rect 48 43670 63 43678
rect -3 43658 63 43670
rect 155 49646 221 49658
rect 155 49638 172 49646
rect 206 49638 221 49646
rect 155 43670 172 43678
rect 206 43670 221 43678
rect 155 43658 221 43670
rect 313 49646 379 49658
rect 313 49638 330 49646
rect 364 49638 379 49646
rect 313 43670 330 43678
rect 364 43670 379 43678
rect 313 43658 379 43670
rect 471 49646 537 49658
rect 471 49638 488 49646
rect 522 49638 537 49646
rect 471 43670 488 43678
rect 522 43670 537 43678
rect 471 43658 537 43670
rect 629 49646 695 49658
rect 629 49638 646 49646
rect 680 49638 695 49646
rect 629 43670 646 43678
rect 680 43670 695 43678
rect 629 43658 695 43670
rect 787 49646 853 49658
rect 787 49638 804 49646
rect 838 49638 853 49646
rect 787 43670 804 43678
rect 838 43670 853 43678
rect 787 43658 853 43670
rect 945 49646 1011 49658
rect 945 49638 962 49646
rect 996 49638 1011 49646
rect 945 43670 962 43678
rect 996 43670 1011 43678
rect 945 43658 1011 43670
rect 1103 49646 1169 49658
rect 1103 49638 1120 49646
rect 1154 49638 1169 49646
rect 1103 43670 1120 43678
rect 1154 43670 1169 43678
rect 1103 43658 1169 43670
rect 1261 49646 1327 49658
rect 1261 49638 1278 49646
rect 1312 49638 1327 49646
rect 1261 43670 1278 43678
rect 1312 43670 1327 43678
rect 1261 43658 1327 43670
rect 1419 49646 1485 49658
rect 1419 49638 1436 49646
rect 1470 49638 1485 49646
rect 1419 43670 1436 43678
rect 1470 43670 1485 43678
rect 1419 43658 1485 43670
rect 1577 49646 1643 49658
rect 1577 49638 1594 49646
rect 1628 49638 1643 49646
rect 1577 43670 1594 43678
rect 1628 43670 1643 43678
rect 1577 43658 1643 43670
rect 1735 49646 1801 49658
rect 1735 49638 1752 49646
rect 1786 49638 1801 49646
rect 1735 43670 1752 43678
rect 1786 43670 1801 43678
rect 1735 43658 1801 43670
rect 1893 49646 1959 49658
rect 1893 49638 1910 49646
rect 1944 49638 1959 49646
rect 1893 43670 1910 43678
rect 1944 43670 1959 43678
rect 1893 43658 1959 43670
rect 2051 49646 2117 49658
rect 2051 49638 2068 49646
rect 2102 49638 2117 49646
rect 2051 43670 2068 43678
rect 2102 43670 2117 43678
rect 2051 43658 2117 43670
rect 2209 49646 2275 49658
rect 2209 49638 2226 49646
rect 2260 49638 2275 49646
rect 2209 43670 2226 43678
rect 2260 43670 2275 43678
rect 2209 43658 2275 43670
rect 2367 49646 2433 49658
rect 2367 49638 2384 49646
rect 2418 49638 2433 49646
rect 2367 43670 2384 43678
rect 2418 43670 2433 43678
rect 2367 43658 2433 43670
rect 2525 49646 2591 49658
rect 2525 49638 2542 49646
rect 2576 49638 2591 49646
rect 2525 43670 2542 43678
rect 2576 43670 2591 43678
rect 2525 43658 2591 43670
rect 2683 49646 2749 49658
rect 2683 49638 2700 49646
rect 2734 49638 2749 49646
rect 2683 43670 2700 43678
rect 2734 43670 2749 43678
rect 2683 43658 2749 43670
rect 2841 49646 2907 49658
rect 2841 49638 2858 49646
rect 2892 49638 2907 49646
rect 2841 43670 2858 43678
rect 2892 43670 2907 43678
rect 2841 43658 2907 43670
rect 2999 49646 3065 49658
rect 2999 49638 3016 49646
rect 3050 49638 3065 49646
rect 2999 43670 3016 43678
rect 3050 43670 3065 43678
rect 2999 43658 3065 43670
rect 3157 49646 3223 49658
rect 3157 49638 3174 49646
rect 3208 49638 3223 49646
rect 3157 43670 3174 43678
rect 3208 43670 3223 43678
rect 3157 43658 3223 43670
rect 3315 49646 3381 49658
rect 3315 49638 3332 49646
rect 3366 49638 3381 49646
rect 3315 43670 3332 43678
rect 3366 43670 3381 43678
rect 3315 43658 3381 43670
rect 3473 49646 3539 49658
rect 3473 49638 3490 49646
rect 3524 49638 3539 49646
rect 3473 43670 3490 43678
rect 3524 43670 3539 43678
rect 3473 43658 3539 43670
rect 3631 49646 3697 49658
rect 3631 49638 3648 49646
rect 3682 49638 3697 49646
rect 3631 43670 3648 43678
rect 3682 43670 3697 43678
rect 3631 43658 3697 43670
rect 3789 49646 3855 49658
rect 3789 49638 3806 49646
rect 3840 49638 3855 49646
rect 3789 43670 3806 43678
rect 3840 43670 3855 43678
rect 3789 43658 3855 43670
rect 3947 49646 4013 49658
rect 3947 49638 3964 49646
rect 3998 49638 4013 49646
rect 3947 43670 3964 43678
rect 3998 43670 4013 43678
rect 3947 43658 4013 43670
rect 4105 49646 4171 49658
rect 4105 49638 4122 49646
rect 4156 49638 4171 49646
rect 4105 43670 4122 43678
rect 4156 43670 4171 43678
rect 4105 43658 4171 43670
rect -568 43620 -548 43626
rect 4086 43620 4106 43626
rect -568 43586 -556 43620
rect 4094 43586 4106 43620
rect -568 43526 -548 43586
rect 4086 43526 4106 43586
rect -770 43494 -700 43500
rect 4240 43494 4310 43500
rect -770 43484 4310 43494
rect -770 43446 -564 43484
rect 4102 43446 4310 43484
rect -770 43430 4310 43446
rect 5530 49870 10610 49880
rect 5530 49832 5736 49870
rect 10459 49832 10610 49870
rect 5530 49822 10610 49832
rect 5530 49820 5600 49822
rect 10540 49820 10610 49822
rect 5732 49730 5752 49790
rect 10386 49730 10406 49790
rect 5732 49696 5744 49730
rect 10394 49696 10406 49730
rect 5732 49690 5752 49696
rect 10386 49690 10406 49696
rect 5665 49646 5731 49658
rect 5665 49638 5682 49646
rect 5716 49638 5731 49646
rect 5665 43670 5682 43678
rect 5716 43670 5731 43678
rect 5665 43658 5731 43670
rect 5823 49646 5889 49658
rect 5823 49638 5840 49646
rect 5874 49638 5889 49646
rect 5823 43670 5840 43678
rect 5874 43670 5889 43678
rect 5823 43658 5889 43670
rect 5981 49646 6047 49658
rect 5981 49638 5998 49646
rect 6032 49638 6047 49646
rect 5981 43670 5998 43678
rect 6032 43670 6047 43678
rect 5981 43658 6047 43670
rect 6139 49646 6205 49658
rect 6139 49638 6156 49646
rect 6190 49638 6205 49646
rect 6139 43670 6156 43678
rect 6190 43670 6205 43678
rect 6139 43658 6205 43670
rect 6297 49646 6363 49658
rect 6297 49638 6314 49646
rect 6348 49638 6363 49646
rect 6297 43670 6314 43678
rect 6348 43670 6363 43678
rect 6297 43658 6363 43670
rect 6455 49646 6521 49658
rect 6455 49638 6472 49646
rect 6506 49638 6521 49646
rect 6455 43670 6472 43678
rect 6506 43670 6521 43678
rect 6455 43658 6521 43670
rect 6613 49646 6679 49658
rect 6613 49638 6630 49646
rect 6664 49638 6679 49646
rect 6613 43670 6630 43678
rect 6664 43670 6679 43678
rect 6613 43658 6679 43670
rect 6771 49646 6837 49658
rect 6771 49638 6788 49646
rect 6822 49638 6837 49646
rect 6771 43670 6788 43678
rect 6822 43670 6837 43678
rect 6771 43658 6837 43670
rect 6929 49646 6995 49658
rect 6929 49638 6946 49646
rect 6980 49638 6995 49646
rect 6929 43670 6946 43678
rect 6980 43670 6995 43678
rect 6929 43658 6995 43670
rect 7087 49646 7153 49658
rect 7087 49638 7104 49646
rect 7138 49638 7153 49646
rect 7087 43670 7104 43678
rect 7138 43670 7153 43678
rect 7087 43658 7153 43670
rect 7245 49646 7311 49658
rect 7245 49638 7262 49646
rect 7296 49638 7311 49646
rect 7245 43670 7262 43678
rect 7296 43670 7311 43678
rect 7245 43658 7311 43670
rect 7403 49646 7469 49658
rect 7403 49638 7420 49646
rect 7454 49638 7469 49646
rect 7403 43670 7420 43678
rect 7454 43670 7469 43678
rect 7403 43658 7469 43670
rect 7561 49646 7627 49658
rect 7561 49638 7578 49646
rect 7612 49638 7627 49646
rect 7561 43670 7578 43678
rect 7612 43670 7627 43678
rect 7561 43658 7627 43670
rect 7719 49646 7785 49658
rect 7719 49638 7736 49646
rect 7770 49638 7785 49646
rect 7719 43670 7736 43678
rect 7770 43670 7785 43678
rect 7719 43658 7785 43670
rect 7877 49646 7943 49658
rect 7877 49638 7894 49646
rect 7928 49638 7943 49646
rect 7877 43670 7894 43678
rect 7928 43670 7943 43678
rect 7877 43658 7943 43670
rect 8035 49646 8101 49658
rect 8035 49638 8052 49646
rect 8086 49638 8101 49646
rect 8035 43670 8052 43678
rect 8086 43670 8101 43678
rect 8035 43658 8101 43670
rect 8193 49646 8259 49658
rect 8193 49638 8210 49646
rect 8244 49638 8259 49646
rect 8193 43670 8210 43678
rect 8244 43670 8259 43678
rect 8193 43658 8259 43670
rect 8351 49646 8417 49658
rect 8351 49638 8368 49646
rect 8402 49638 8417 49646
rect 8351 43670 8368 43678
rect 8402 43670 8417 43678
rect 8351 43658 8417 43670
rect 8509 49646 8575 49658
rect 8509 49638 8526 49646
rect 8560 49638 8575 49646
rect 8509 43670 8526 43678
rect 8560 43670 8575 43678
rect 8509 43658 8575 43670
rect 8667 49646 8733 49658
rect 8667 49638 8684 49646
rect 8718 49638 8733 49646
rect 8667 43670 8684 43678
rect 8718 43670 8733 43678
rect 8667 43658 8733 43670
rect 8825 49646 8891 49658
rect 8825 49638 8842 49646
rect 8876 49638 8891 49646
rect 8825 43670 8842 43678
rect 8876 43670 8891 43678
rect 8825 43658 8891 43670
rect 8983 49646 9049 49658
rect 8983 49638 9000 49646
rect 9034 49638 9049 49646
rect 8983 43670 9000 43678
rect 9034 43670 9049 43678
rect 8983 43658 9049 43670
rect 9141 49646 9207 49658
rect 9141 49638 9158 49646
rect 9192 49638 9207 49646
rect 9141 43670 9158 43678
rect 9192 43670 9207 43678
rect 9141 43658 9207 43670
rect 9299 49646 9365 49658
rect 9299 49638 9316 49646
rect 9350 49638 9365 49646
rect 9299 43670 9316 43678
rect 9350 43670 9365 43678
rect 9299 43658 9365 43670
rect 9457 49646 9523 49658
rect 9457 49638 9474 49646
rect 9508 49638 9523 49646
rect 9457 43670 9474 43678
rect 9508 43670 9523 43678
rect 9457 43658 9523 43670
rect 9615 49646 9681 49658
rect 9615 49638 9632 49646
rect 9666 49638 9681 49646
rect 9615 43670 9632 43678
rect 9666 43670 9681 43678
rect 9615 43658 9681 43670
rect 9773 49646 9839 49658
rect 9773 49638 9790 49646
rect 9824 49638 9839 49646
rect 9773 43670 9790 43678
rect 9824 43670 9839 43678
rect 9773 43658 9839 43670
rect 9931 49646 9997 49658
rect 9931 49638 9948 49646
rect 9982 49638 9997 49646
rect 9931 43670 9948 43678
rect 9982 43670 9997 43678
rect 9931 43658 9997 43670
rect 10089 49646 10155 49658
rect 10089 49638 10106 49646
rect 10140 49638 10155 49646
rect 10089 43670 10106 43678
rect 10140 43670 10155 43678
rect 10089 43658 10155 43670
rect 10247 49646 10313 49658
rect 10247 49638 10264 49646
rect 10298 49638 10313 49646
rect 10247 43670 10264 43678
rect 10298 43670 10313 43678
rect 10247 43658 10313 43670
rect 10405 49646 10471 49658
rect 10405 49638 10422 49646
rect 10456 49638 10471 49646
rect 10405 43670 10422 43678
rect 10456 43670 10471 43678
rect 10405 43658 10471 43670
rect 5732 43620 5752 43626
rect 10386 43620 10406 43626
rect 5732 43586 5744 43620
rect 10394 43586 10406 43620
rect 5732 43526 5752 43586
rect 10386 43526 10406 43586
rect 5530 43494 5600 43500
rect 10540 43494 10610 43500
rect 5530 43484 10610 43494
rect 5530 43446 5736 43484
rect 10402 43446 10610 43484
rect 5530 43430 10610 43446
rect -13370 42870 -8290 42880
rect -13370 42832 -13164 42870
rect -8441 42832 -8290 42870
rect -13370 42822 -8290 42832
rect -13370 42820 -13300 42822
rect -8360 42820 -8290 42822
rect -13168 42730 -13148 42790
rect -8514 42730 -8494 42790
rect -13168 42696 -13156 42730
rect -8506 42696 -8494 42730
rect -13168 42690 -13148 42696
rect -8514 42690 -8494 42696
rect -13235 42646 -13169 42658
rect -13235 42638 -13218 42646
rect -13184 42638 -13169 42646
rect -13235 36670 -13218 36678
rect -13184 36670 -13169 36678
rect -13235 36658 -13169 36670
rect -13077 42646 -13011 42658
rect -13077 42638 -13060 42646
rect -13026 42638 -13011 42646
rect -13077 36670 -13060 36678
rect -13026 36670 -13011 36678
rect -13077 36658 -13011 36670
rect -12919 42646 -12853 42658
rect -12919 42638 -12902 42646
rect -12868 42638 -12853 42646
rect -12919 36670 -12902 36678
rect -12868 36670 -12853 36678
rect -12919 36658 -12853 36670
rect -12761 42646 -12695 42658
rect -12761 42638 -12744 42646
rect -12710 42638 -12695 42646
rect -12761 36670 -12744 36678
rect -12710 36670 -12695 36678
rect -12761 36658 -12695 36670
rect -12603 42646 -12537 42658
rect -12603 42638 -12586 42646
rect -12552 42638 -12537 42646
rect -12603 36670 -12586 36678
rect -12552 36670 -12537 36678
rect -12603 36658 -12537 36670
rect -12445 42646 -12379 42658
rect -12445 42638 -12428 42646
rect -12394 42638 -12379 42646
rect -12445 36670 -12428 36678
rect -12394 36670 -12379 36678
rect -12445 36658 -12379 36670
rect -12287 42646 -12221 42658
rect -12287 42638 -12270 42646
rect -12236 42638 -12221 42646
rect -12287 36670 -12270 36678
rect -12236 36670 -12221 36678
rect -12287 36658 -12221 36670
rect -12129 42646 -12063 42658
rect -12129 42638 -12112 42646
rect -12078 42638 -12063 42646
rect -12129 36670 -12112 36678
rect -12078 36670 -12063 36678
rect -12129 36658 -12063 36670
rect -11971 42646 -11905 42658
rect -11971 42638 -11954 42646
rect -11920 42638 -11905 42646
rect -11971 36670 -11954 36678
rect -11920 36670 -11905 36678
rect -11971 36658 -11905 36670
rect -11813 42646 -11747 42658
rect -11813 42638 -11796 42646
rect -11762 42638 -11747 42646
rect -11813 36670 -11796 36678
rect -11762 36670 -11747 36678
rect -11813 36658 -11747 36670
rect -11655 42646 -11589 42658
rect -11655 42638 -11638 42646
rect -11604 42638 -11589 42646
rect -11655 36670 -11638 36678
rect -11604 36670 -11589 36678
rect -11655 36658 -11589 36670
rect -11497 42646 -11431 42658
rect -11497 42638 -11480 42646
rect -11446 42638 -11431 42646
rect -11497 36670 -11480 36678
rect -11446 36670 -11431 36678
rect -11497 36658 -11431 36670
rect -11339 42646 -11273 42658
rect -11339 42638 -11322 42646
rect -11288 42638 -11273 42646
rect -11339 36670 -11322 36678
rect -11288 36670 -11273 36678
rect -11339 36658 -11273 36670
rect -11181 42646 -11115 42658
rect -11181 42638 -11164 42646
rect -11130 42638 -11115 42646
rect -11181 36670 -11164 36678
rect -11130 36670 -11115 36678
rect -11181 36658 -11115 36670
rect -11023 42646 -10957 42658
rect -11023 42638 -11006 42646
rect -10972 42638 -10957 42646
rect -11023 36670 -11006 36678
rect -10972 36670 -10957 36678
rect -11023 36658 -10957 36670
rect -10865 42646 -10799 42658
rect -10865 42638 -10848 42646
rect -10814 42638 -10799 42646
rect -10865 36670 -10848 36678
rect -10814 36670 -10799 36678
rect -10865 36658 -10799 36670
rect -10707 42646 -10641 42658
rect -10707 42638 -10690 42646
rect -10656 42638 -10641 42646
rect -10707 36670 -10690 36678
rect -10656 36670 -10641 36678
rect -10707 36658 -10641 36670
rect -10549 42646 -10483 42658
rect -10549 42638 -10532 42646
rect -10498 42638 -10483 42646
rect -10549 36670 -10532 36678
rect -10498 36670 -10483 36678
rect -10549 36658 -10483 36670
rect -10391 42646 -10325 42658
rect -10391 42638 -10374 42646
rect -10340 42638 -10325 42646
rect -10391 36670 -10374 36678
rect -10340 36670 -10325 36678
rect -10391 36658 -10325 36670
rect -10233 42646 -10167 42658
rect -10233 42638 -10216 42646
rect -10182 42638 -10167 42646
rect -10233 36670 -10216 36678
rect -10182 36670 -10167 36678
rect -10233 36658 -10167 36670
rect -10075 42646 -10009 42658
rect -10075 42638 -10058 42646
rect -10024 42638 -10009 42646
rect -10075 36670 -10058 36678
rect -10024 36670 -10009 36678
rect -10075 36658 -10009 36670
rect -9917 42646 -9851 42658
rect -9917 42638 -9900 42646
rect -9866 42638 -9851 42646
rect -9917 36670 -9900 36678
rect -9866 36670 -9851 36678
rect -9917 36658 -9851 36670
rect -9759 42646 -9693 42658
rect -9759 42638 -9742 42646
rect -9708 42638 -9693 42646
rect -9759 36670 -9742 36678
rect -9708 36670 -9693 36678
rect -9759 36658 -9693 36670
rect -9601 42646 -9535 42658
rect -9601 42638 -9584 42646
rect -9550 42638 -9535 42646
rect -9601 36670 -9584 36678
rect -9550 36670 -9535 36678
rect -9601 36658 -9535 36670
rect -9443 42646 -9377 42658
rect -9443 42638 -9426 42646
rect -9392 42638 -9377 42646
rect -9443 36670 -9426 36678
rect -9392 36670 -9377 36678
rect -9443 36658 -9377 36670
rect -9285 42646 -9219 42658
rect -9285 42638 -9268 42646
rect -9234 42638 -9219 42646
rect -9285 36670 -9268 36678
rect -9234 36670 -9219 36678
rect -9285 36658 -9219 36670
rect -9127 42646 -9061 42658
rect -9127 42638 -9110 42646
rect -9076 42638 -9061 42646
rect -9127 36670 -9110 36678
rect -9076 36670 -9061 36678
rect -9127 36658 -9061 36670
rect -8969 42646 -8903 42658
rect -8969 42638 -8952 42646
rect -8918 42638 -8903 42646
rect -8969 36670 -8952 36678
rect -8918 36670 -8903 36678
rect -8969 36658 -8903 36670
rect -8811 42646 -8745 42658
rect -8811 42638 -8794 42646
rect -8760 42638 -8745 42646
rect -8811 36670 -8794 36678
rect -8760 36670 -8745 36678
rect -8811 36658 -8745 36670
rect -8653 42646 -8587 42658
rect -8653 42638 -8636 42646
rect -8602 42638 -8587 42646
rect -8653 36670 -8636 36678
rect -8602 36670 -8587 36678
rect -8653 36658 -8587 36670
rect -8495 42646 -8429 42658
rect -8495 42638 -8478 42646
rect -8444 42638 -8429 42646
rect -8495 36670 -8478 36678
rect -8444 36670 -8429 36678
rect -8495 36658 -8429 36670
rect -13168 36620 -13148 36626
rect -8514 36620 -8494 36626
rect -13168 36586 -13156 36620
rect -8506 36586 -8494 36620
rect -13168 36526 -13148 36586
rect -8514 36526 -8494 36586
rect -13370 36494 -13300 36500
rect -8360 36494 -8290 36500
rect -13370 36484 -8290 36494
rect -13370 36446 -13164 36484
rect -8498 36446 -8290 36484
rect -13370 36430 -8290 36446
rect -7070 42870 -1990 42880
rect -7070 42832 -6864 42870
rect -2141 42832 -1990 42870
rect -7070 42822 -1990 42832
rect -7070 42820 -7000 42822
rect -2060 42820 -1990 42822
rect -6868 42730 -6848 42790
rect -2214 42730 -2194 42790
rect -6868 42696 -6856 42730
rect -2206 42696 -2194 42730
rect -6868 42690 -6848 42696
rect -2214 42690 -2194 42696
rect -6935 42646 -6869 42658
rect -6935 42638 -6918 42646
rect -6884 42638 -6869 42646
rect -6935 36670 -6918 36678
rect -6884 36670 -6869 36678
rect -6935 36658 -6869 36670
rect -6777 42646 -6711 42658
rect -6777 42638 -6760 42646
rect -6726 42638 -6711 42646
rect -6777 36670 -6760 36678
rect -6726 36670 -6711 36678
rect -6777 36658 -6711 36670
rect -6619 42646 -6553 42658
rect -6619 42638 -6602 42646
rect -6568 42638 -6553 42646
rect -6619 36670 -6602 36678
rect -6568 36670 -6553 36678
rect -6619 36658 -6553 36670
rect -6461 42646 -6395 42658
rect -6461 42638 -6444 42646
rect -6410 42638 -6395 42646
rect -6461 36670 -6444 36678
rect -6410 36670 -6395 36678
rect -6461 36658 -6395 36670
rect -6303 42646 -6237 42658
rect -6303 42638 -6286 42646
rect -6252 42638 -6237 42646
rect -6303 36670 -6286 36678
rect -6252 36670 -6237 36678
rect -6303 36658 -6237 36670
rect -6145 42646 -6079 42658
rect -6145 42638 -6128 42646
rect -6094 42638 -6079 42646
rect -6145 36670 -6128 36678
rect -6094 36670 -6079 36678
rect -6145 36658 -6079 36670
rect -5987 42646 -5921 42658
rect -5987 42638 -5970 42646
rect -5936 42638 -5921 42646
rect -5987 36670 -5970 36678
rect -5936 36670 -5921 36678
rect -5987 36658 -5921 36670
rect -5829 42646 -5763 42658
rect -5829 42638 -5812 42646
rect -5778 42638 -5763 42646
rect -5829 36670 -5812 36678
rect -5778 36670 -5763 36678
rect -5829 36658 -5763 36670
rect -5671 42646 -5605 42658
rect -5671 42638 -5654 42646
rect -5620 42638 -5605 42646
rect -5671 36670 -5654 36678
rect -5620 36670 -5605 36678
rect -5671 36658 -5605 36670
rect -5513 42646 -5447 42658
rect -5513 42638 -5496 42646
rect -5462 42638 -5447 42646
rect -5513 36670 -5496 36678
rect -5462 36670 -5447 36678
rect -5513 36658 -5447 36670
rect -5355 42646 -5289 42658
rect -5355 42638 -5338 42646
rect -5304 42638 -5289 42646
rect -5355 36670 -5338 36678
rect -5304 36670 -5289 36678
rect -5355 36658 -5289 36670
rect -5197 42646 -5131 42658
rect -5197 42638 -5180 42646
rect -5146 42638 -5131 42646
rect -5197 36670 -5180 36678
rect -5146 36670 -5131 36678
rect -5197 36658 -5131 36670
rect -5039 42646 -4973 42658
rect -5039 42638 -5022 42646
rect -4988 42638 -4973 42646
rect -5039 36670 -5022 36678
rect -4988 36670 -4973 36678
rect -5039 36658 -4973 36670
rect -4881 42646 -4815 42658
rect -4881 42638 -4864 42646
rect -4830 42638 -4815 42646
rect -4881 36670 -4864 36678
rect -4830 36670 -4815 36678
rect -4881 36658 -4815 36670
rect -4723 42646 -4657 42658
rect -4723 42638 -4706 42646
rect -4672 42638 -4657 42646
rect -4723 36670 -4706 36678
rect -4672 36670 -4657 36678
rect -4723 36658 -4657 36670
rect -4565 42646 -4499 42658
rect -4565 42638 -4548 42646
rect -4514 42638 -4499 42646
rect -4565 36670 -4548 36678
rect -4514 36670 -4499 36678
rect -4565 36658 -4499 36670
rect -4407 42646 -4341 42658
rect -4407 42638 -4390 42646
rect -4356 42638 -4341 42646
rect -4407 36670 -4390 36678
rect -4356 36670 -4341 36678
rect -4407 36658 -4341 36670
rect -4249 42646 -4183 42658
rect -4249 42638 -4232 42646
rect -4198 42638 -4183 42646
rect -4249 36670 -4232 36678
rect -4198 36670 -4183 36678
rect -4249 36658 -4183 36670
rect -4091 42646 -4025 42658
rect -4091 42638 -4074 42646
rect -4040 42638 -4025 42646
rect -4091 36670 -4074 36678
rect -4040 36670 -4025 36678
rect -4091 36658 -4025 36670
rect -3933 42646 -3867 42658
rect -3933 42638 -3916 42646
rect -3882 42638 -3867 42646
rect -3933 36670 -3916 36678
rect -3882 36670 -3867 36678
rect -3933 36658 -3867 36670
rect -3775 42646 -3709 42658
rect -3775 42638 -3758 42646
rect -3724 42638 -3709 42646
rect -3775 36670 -3758 36678
rect -3724 36670 -3709 36678
rect -3775 36658 -3709 36670
rect -3617 42646 -3551 42658
rect -3617 42638 -3600 42646
rect -3566 42638 -3551 42646
rect -3617 36670 -3600 36678
rect -3566 36670 -3551 36678
rect -3617 36658 -3551 36670
rect -3459 42646 -3393 42658
rect -3459 42638 -3442 42646
rect -3408 42638 -3393 42646
rect -3459 36670 -3442 36678
rect -3408 36670 -3393 36678
rect -3459 36658 -3393 36670
rect -3301 42646 -3235 42658
rect -3301 42638 -3284 42646
rect -3250 42638 -3235 42646
rect -3301 36670 -3284 36678
rect -3250 36670 -3235 36678
rect -3301 36658 -3235 36670
rect -3143 42646 -3077 42658
rect -3143 42638 -3126 42646
rect -3092 42638 -3077 42646
rect -3143 36670 -3126 36678
rect -3092 36670 -3077 36678
rect -3143 36658 -3077 36670
rect -2985 42646 -2919 42658
rect -2985 42638 -2968 42646
rect -2934 42638 -2919 42646
rect -2985 36670 -2968 36678
rect -2934 36670 -2919 36678
rect -2985 36658 -2919 36670
rect -2827 42646 -2761 42658
rect -2827 42638 -2810 42646
rect -2776 42638 -2761 42646
rect -2827 36670 -2810 36678
rect -2776 36670 -2761 36678
rect -2827 36658 -2761 36670
rect -2669 42646 -2603 42658
rect -2669 42638 -2652 42646
rect -2618 42638 -2603 42646
rect -2669 36670 -2652 36678
rect -2618 36670 -2603 36678
rect -2669 36658 -2603 36670
rect -2511 42646 -2445 42658
rect -2511 42638 -2494 42646
rect -2460 42638 -2445 42646
rect -2511 36670 -2494 36678
rect -2460 36670 -2445 36678
rect -2511 36658 -2445 36670
rect -2353 42646 -2287 42658
rect -2353 42638 -2336 42646
rect -2302 42638 -2287 42646
rect -2353 36670 -2336 36678
rect -2302 36670 -2287 36678
rect -2353 36658 -2287 36670
rect -2195 42646 -2129 42658
rect -2195 42638 -2178 42646
rect -2144 42638 -2129 42646
rect -2195 36670 -2178 36678
rect -2144 36670 -2129 36678
rect -2195 36658 -2129 36670
rect -6868 36620 -6848 36626
rect -2214 36620 -2194 36626
rect -6868 36586 -6856 36620
rect -2206 36586 -2194 36620
rect -6868 36526 -6848 36586
rect -2214 36526 -2194 36586
rect -7070 36494 -7000 36500
rect -2060 36494 -1990 36500
rect -7070 36484 -1990 36494
rect -7070 36446 -6864 36484
rect -2198 36446 -1990 36484
rect -7070 36430 -1990 36446
rect -770 42870 4310 42880
rect -770 42832 -564 42870
rect 4159 42832 4310 42870
rect -770 42822 4310 42832
rect -770 42820 -700 42822
rect 4240 42820 4310 42822
rect -568 42730 -548 42790
rect 4086 42730 4106 42790
rect -568 42696 -556 42730
rect 4094 42696 4106 42730
rect -568 42690 -548 42696
rect 4086 42690 4106 42696
rect -635 42646 -569 42658
rect -635 42638 -618 42646
rect -584 42638 -569 42646
rect -635 36670 -618 36678
rect -584 36670 -569 36678
rect -635 36658 -569 36670
rect -477 42646 -411 42658
rect -477 42638 -460 42646
rect -426 42638 -411 42646
rect -477 36670 -460 36678
rect -426 36670 -411 36678
rect -477 36658 -411 36670
rect -319 42646 -253 42658
rect -319 42638 -302 42646
rect -268 42638 -253 42646
rect -319 36670 -302 36678
rect -268 36670 -253 36678
rect -319 36658 -253 36670
rect -161 42646 -95 42658
rect -161 42638 -144 42646
rect -110 42638 -95 42646
rect -161 36670 -144 36678
rect -110 36670 -95 36678
rect -161 36658 -95 36670
rect -3 42646 63 42658
rect -3 42638 14 42646
rect 48 42638 63 42646
rect -3 36670 14 36678
rect 48 36670 63 36678
rect -3 36658 63 36670
rect 155 42646 221 42658
rect 155 42638 172 42646
rect 206 42638 221 42646
rect 155 36670 172 36678
rect 206 36670 221 36678
rect 155 36658 221 36670
rect 313 42646 379 42658
rect 313 42638 330 42646
rect 364 42638 379 42646
rect 313 36670 330 36678
rect 364 36670 379 36678
rect 313 36658 379 36670
rect 471 42646 537 42658
rect 471 42638 488 42646
rect 522 42638 537 42646
rect 471 36670 488 36678
rect 522 36670 537 36678
rect 471 36658 537 36670
rect 629 42646 695 42658
rect 629 42638 646 42646
rect 680 42638 695 42646
rect 629 36670 646 36678
rect 680 36670 695 36678
rect 629 36658 695 36670
rect 787 42646 853 42658
rect 787 42638 804 42646
rect 838 42638 853 42646
rect 787 36670 804 36678
rect 838 36670 853 36678
rect 787 36658 853 36670
rect 945 42646 1011 42658
rect 945 42638 962 42646
rect 996 42638 1011 42646
rect 945 36670 962 36678
rect 996 36670 1011 36678
rect 945 36658 1011 36670
rect 1103 42646 1169 42658
rect 1103 42638 1120 42646
rect 1154 42638 1169 42646
rect 1103 36670 1120 36678
rect 1154 36670 1169 36678
rect 1103 36658 1169 36670
rect 1261 42646 1327 42658
rect 1261 42638 1278 42646
rect 1312 42638 1327 42646
rect 1261 36670 1278 36678
rect 1312 36670 1327 36678
rect 1261 36658 1327 36670
rect 1419 42646 1485 42658
rect 1419 42638 1436 42646
rect 1470 42638 1485 42646
rect 1419 36670 1436 36678
rect 1470 36670 1485 36678
rect 1419 36658 1485 36670
rect 1577 42646 1643 42658
rect 1577 42638 1594 42646
rect 1628 42638 1643 42646
rect 1577 36670 1594 36678
rect 1628 36670 1643 36678
rect 1577 36658 1643 36670
rect 1735 42646 1801 42658
rect 1735 42638 1752 42646
rect 1786 42638 1801 42646
rect 1735 36670 1752 36678
rect 1786 36670 1801 36678
rect 1735 36658 1801 36670
rect 1893 42646 1959 42658
rect 1893 42638 1910 42646
rect 1944 42638 1959 42646
rect 1893 36670 1910 36678
rect 1944 36670 1959 36678
rect 1893 36658 1959 36670
rect 2051 42646 2117 42658
rect 2051 42638 2068 42646
rect 2102 42638 2117 42646
rect 2051 36670 2068 36678
rect 2102 36670 2117 36678
rect 2051 36658 2117 36670
rect 2209 42646 2275 42658
rect 2209 42638 2226 42646
rect 2260 42638 2275 42646
rect 2209 36670 2226 36678
rect 2260 36670 2275 36678
rect 2209 36658 2275 36670
rect 2367 42646 2433 42658
rect 2367 42638 2384 42646
rect 2418 42638 2433 42646
rect 2367 36670 2384 36678
rect 2418 36670 2433 36678
rect 2367 36658 2433 36670
rect 2525 42646 2591 42658
rect 2525 42638 2542 42646
rect 2576 42638 2591 42646
rect 2525 36670 2542 36678
rect 2576 36670 2591 36678
rect 2525 36658 2591 36670
rect 2683 42646 2749 42658
rect 2683 42638 2700 42646
rect 2734 42638 2749 42646
rect 2683 36670 2700 36678
rect 2734 36670 2749 36678
rect 2683 36658 2749 36670
rect 2841 42646 2907 42658
rect 2841 42638 2858 42646
rect 2892 42638 2907 42646
rect 2841 36670 2858 36678
rect 2892 36670 2907 36678
rect 2841 36658 2907 36670
rect 2999 42646 3065 42658
rect 2999 42638 3016 42646
rect 3050 42638 3065 42646
rect 2999 36670 3016 36678
rect 3050 36670 3065 36678
rect 2999 36658 3065 36670
rect 3157 42646 3223 42658
rect 3157 42638 3174 42646
rect 3208 42638 3223 42646
rect 3157 36670 3174 36678
rect 3208 36670 3223 36678
rect 3157 36658 3223 36670
rect 3315 42646 3381 42658
rect 3315 42638 3332 42646
rect 3366 42638 3381 42646
rect 3315 36670 3332 36678
rect 3366 36670 3381 36678
rect 3315 36658 3381 36670
rect 3473 42646 3539 42658
rect 3473 42638 3490 42646
rect 3524 42638 3539 42646
rect 3473 36670 3490 36678
rect 3524 36670 3539 36678
rect 3473 36658 3539 36670
rect 3631 42646 3697 42658
rect 3631 42638 3648 42646
rect 3682 42638 3697 42646
rect 3631 36670 3648 36678
rect 3682 36670 3697 36678
rect 3631 36658 3697 36670
rect 3789 42646 3855 42658
rect 3789 42638 3806 42646
rect 3840 42638 3855 42646
rect 3789 36670 3806 36678
rect 3840 36670 3855 36678
rect 3789 36658 3855 36670
rect 3947 42646 4013 42658
rect 3947 42638 3964 42646
rect 3998 42638 4013 42646
rect 3947 36670 3964 36678
rect 3998 36670 4013 36678
rect 3947 36658 4013 36670
rect 4105 42646 4171 42658
rect 4105 42638 4122 42646
rect 4156 42638 4171 42646
rect 4105 36670 4122 36678
rect 4156 36670 4171 36678
rect 4105 36658 4171 36670
rect -568 36620 -548 36626
rect 4086 36620 4106 36626
rect -568 36586 -556 36620
rect 4094 36586 4106 36620
rect -568 36526 -548 36586
rect 4086 36526 4106 36586
rect -770 36494 -700 36500
rect 4240 36494 4310 36500
rect -770 36484 4310 36494
rect -770 36446 -564 36484
rect 4102 36446 4310 36484
rect -770 36430 4310 36446
rect 5530 42870 10610 42880
rect 5530 42832 5736 42870
rect 10459 42832 10610 42870
rect 5530 42822 10610 42832
rect 5530 42820 5600 42822
rect 10540 42820 10610 42822
rect 5732 42730 5752 42790
rect 10386 42730 10406 42790
rect 5732 42696 5744 42730
rect 10394 42696 10406 42730
rect 5732 42690 5752 42696
rect 10386 42690 10406 42696
rect 5665 42646 5731 42658
rect 5665 42638 5682 42646
rect 5716 42638 5731 42646
rect 5665 36670 5682 36678
rect 5716 36670 5731 36678
rect 5665 36658 5731 36670
rect 5823 42646 5889 42658
rect 5823 42638 5840 42646
rect 5874 42638 5889 42646
rect 5823 36670 5840 36678
rect 5874 36670 5889 36678
rect 5823 36658 5889 36670
rect 5981 42646 6047 42658
rect 5981 42638 5998 42646
rect 6032 42638 6047 42646
rect 5981 36670 5998 36678
rect 6032 36670 6047 36678
rect 5981 36658 6047 36670
rect 6139 42646 6205 42658
rect 6139 42638 6156 42646
rect 6190 42638 6205 42646
rect 6139 36670 6156 36678
rect 6190 36670 6205 36678
rect 6139 36658 6205 36670
rect 6297 42646 6363 42658
rect 6297 42638 6314 42646
rect 6348 42638 6363 42646
rect 6297 36670 6314 36678
rect 6348 36670 6363 36678
rect 6297 36658 6363 36670
rect 6455 42646 6521 42658
rect 6455 42638 6472 42646
rect 6506 42638 6521 42646
rect 6455 36670 6472 36678
rect 6506 36670 6521 36678
rect 6455 36658 6521 36670
rect 6613 42646 6679 42658
rect 6613 42638 6630 42646
rect 6664 42638 6679 42646
rect 6613 36670 6630 36678
rect 6664 36670 6679 36678
rect 6613 36658 6679 36670
rect 6771 42646 6837 42658
rect 6771 42638 6788 42646
rect 6822 42638 6837 42646
rect 6771 36670 6788 36678
rect 6822 36670 6837 36678
rect 6771 36658 6837 36670
rect 6929 42646 6995 42658
rect 6929 42638 6946 42646
rect 6980 42638 6995 42646
rect 6929 36670 6946 36678
rect 6980 36670 6995 36678
rect 6929 36658 6995 36670
rect 7087 42646 7153 42658
rect 7087 42638 7104 42646
rect 7138 42638 7153 42646
rect 7087 36670 7104 36678
rect 7138 36670 7153 36678
rect 7087 36658 7153 36670
rect 7245 42646 7311 42658
rect 7245 42638 7262 42646
rect 7296 42638 7311 42646
rect 7245 36670 7262 36678
rect 7296 36670 7311 36678
rect 7245 36658 7311 36670
rect 7403 42646 7469 42658
rect 7403 42638 7420 42646
rect 7454 42638 7469 42646
rect 7403 36670 7420 36678
rect 7454 36670 7469 36678
rect 7403 36658 7469 36670
rect 7561 42646 7627 42658
rect 7561 42638 7578 42646
rect 7612 42638 7627 42646
rect 7561 36670 7578 36678
rect 7612 36670 7627 36678
rect 7561 36658 7627 36670
rect 7719 42646 7785 42658
rect 7719 42638 7736 42646
rect 7770 42638 7785 42646
rect 7719 36670 7736 36678
rect 7770 36670 7785 36678
rect 7719 36658 7785 36670
rect 7877 42646 7943 42658
rect 7877 42638 7894 42646
rect 7928 42638 7943 42646
rect 7877 36670 7894 36678
rect 7928 36670 7943 36678
rect 7877 36658 7943 36670
rect 8035 42646 8101 42658
rect 8035 42638 8052 42646
rect 8086 42638 8101 42646
rect 8035 36670 8052 36678
rect 8086 36670 8101 36678
rect 8035 36658 8101 36670
rect 8193 42646 8259 42658
rect 8193 42638 8210 42646
rect 8244 42638 8259 42646
rect 8193 36670 8210 36678
rect 8244 36670 8259 36678
rect 8193 36658 8259 36670
rect 8351 42646 8417 42658
rect 8351 42638 8368 42646
rect 8402 42638 8417 42646
rect 8351 36670 8368 36678
rect 8402 36670 8417 36678
rect 8351 36658 8417 36670
rect 8509 42646 8575 42658
rect 8509 42638 8526 42646
rect 8560 42638 8575 42646
rect 8509 36670 8526 36678
rect 8560 36670 8575 36678
rect 8509 36658 8575 36670
rect 8667 42646 8733 42658
rect 8667 42638 8684 42646
rect 8718 42638 8733 42646
rect 8667 36670 8684 36678
rect 8718 36670 8733 36678
rect 8667 36658 8733 36670
rect 8825 42646 8891 42658
rect 8825 42638 8842 42646
rect 8876 42638 8891 42646
rect 8825 36670 8842 36678
rect 8876 36670 8891 36678
rect 8825 36658 8891 36670
rect 8983 42646 9049 42658
rect 8983 42638 9000 42646
rect 9034 42638 9049 42646
rect 8983 36670 9000 36678
rect 9034 36670 9049 36678
rect 8983 36658 9049 36670
rect 9141 42646 9207 42658
rect 9141 42638 9158 42646
rect 9192 42638 9207 42646
rect 9141 36670 9158 36678
rect 9192 36670 9207 36678
rect 9141 36658 9207 36670
rect 9299 42646 9365 42658
rect 9299 42638 9316 42646
rect 9350 42638 9365 42646
rect 9299 36670 9316 36678
rect 9350 36670 9365 36678
rect 9299 36658 9365 36670
rect 9457 42646 9523 42658
rect 9457 42638 9474 42646
rect 9508 42638 9523 42646
rect 9457 36670 9474 36678
rect 9508 36670 9523 36678
rect 9457 36658 9523 36670
rect 9615 42646 9681 42658
rect 9615 42638 9632 42646
rect 9666 42638 9681 42646
rect 9615 36670 9632 36678
rect 9666 36670 9681 36678
rect 9615 36658 9681 36670
rect 9773 42646 9839 42658
rect 9773 42638 9790 42646
rect 9824 42638 9839 42646
rect 9773 36670 9790 36678
rect 9824 36670 9839 36678
rect 9773 36658 9839 36670
rect 9931 42646 9997 42658
rect 9931 42638 9948 42646
rect 9982 42638 9997 42646
rect 9931 36670 9948 36678
rect 9982 36670 9997 36678
rect 9931 36658 9997 36670
rect 10089 42646 10155 42658
rect 10089 42638 10106 42646
rect 10140 42638 10155 42646
rect 10089 36670 10106 36678
rect 10140 36670 10155 36678
rect 10089 36658 10155 36670
rect 10247 42646 10313 42658
rect 10247 42638 10264 42646
rect 10298 42638 10313 42646
rect 10247 36670 10264 36678
rect 10298 36670 10313 36678
rect 10247 36658 10313 36670
rect 10405 42646 10471 42658
rect 10405 42638 10422 42646
rect 10456 42638 10471 42646
rect 10405 36670 10422 36678
rect 10456 36670 10471 36678
rect 10405 36658 10471 36670
rect 5732 36620 5752 36626
rect 10386 36620 10406 36626
rect 5732 36586 5744 36620
rect 10394 36586 10406 36620
rect 5732 36526 5752 36586
rect 10386 36526 10406 36586
rect 5530 36494 5600 36500
rect 10540 36494 10610 36500
rect 5530 36484 10610 36494
rect 5530 36446 5736 36484
rect 10402 36446 10610 36484
rect 5530 36430 10610 36446
rect -13370 34570 -8290 34580
rect -13370 34532 -13164 34570
rect -8441 34532 -8290 34570
rect -13370 34522 -8290 34532
rect -13370 34520 -13300 34522
rect -8360 34520 -8290 34522
rect -13168 34430 -13148 34490
rect -8514 34430 -8494 34490
rect -13168 34396 -13156 34430
rect -8506 34396 -8494 34430
rect -13168 34390 -13148 34396
rect -8514 34390 -8494 34396
rect -13235 34346 -13169 34358
rect -13235 34338 -13218 34346
rect -13184 34338 -13169 34346
rect -13235 28370 -13218 28378
rect -13184 28370 -13169 28378
rect -13235 28358 -13169 28370
rect -13077 34346 -13011 34358
rect -13077 34338 -13060 34346
rect -13026 34338 -13011 34346
rect -13077 28370 -13060 28378
rect -13026 28370 -13011 28378
rect -13077 28358 -13011 28370
rect -12919 34346 -12853 34358
rect -12919 34338 -12902 34346
rect -12868 34338 -12853 34346
rect -12919 28370 -12902 28378
rect -12868 28370 -12853 28378
rect -12919 28358 -12853 28370
rect -12761 34346 -12695 34358
rect -12761 34338 -12744 34346
rect -12710 34338 -12695 34346
rect -12761 28370 -12744 28378
rect -12710 28370 -12695 28378
rect -12761 28358 -12695 28370
rect -12603 34346 -12537 34358
rect -12603 34338 -12586 34346
rect -12552 34338 -12537 34346
rect -12603 28370 -12586 28378
rect -12552 28370 -12537 28378
rect -12603 28358 -12537 28370
rect -12445 34346 -12379 34358
rect -12445 34338 -12428 34346
rect -12394 34338 -12379 34346
rect -12445 28370 -12428 28378
rect -12394 28370 -12379 28378
rect -12445 28358 -12379 28370
rect -12287 34346 -12221 34358
rect -12287 34338 -12270 34346
rect -12236 34338 -12221 34346
rect -12287 28370 -12270 28378
rect -12236 28370 -12221 28378
rect -12287 28358 -12221 28370
rect -12129 34346 -12063 34358
rect -12129 34338 -12112 34346
rect -12078 34338 -12063 34346
rect -12129 28370 -12112 28378
rect -12078 28370 -12063 28378
rect -12129 28358 -12063 28370
rect -11971 34346 -11905 34358
rect -11971 34338 -11954 34346
rect -11920 34338 -11905 34346
rect -11971 28370 -11954 28378
rect -11920 28370 -11905 28378
rect -11971 28358 -11905 28370
rect -11813 34346 -11747 34358
rect -11813 34338 -11796 34346
rect -11762 34338 -11747 34346
rect -11813 28370 -11796 28378
rect -11762 28370 -11747 28378
rect -11813 28358 -11747 28370
rect -11655 34346 -11589 34358
rect -11655 34338 -11638 34346
rect -11604 34338 -11589 34346
rect -11655 28370 -11638 28378
rect -11604 28370 -11589 28378
rect -11655 28358 -11589 28370
rect -11497 34346 -11431 34358
rect -11497 34338 -11480 34346
rect -11446 34338 -11431 34346
rect -11497 28370 -11480 28378
rect -11446 28370 -11431 28378
rect -11497 28358 -11431 28370
rect -11339 34346 -11273 34358
rect -11339 34338 -11322 34346
rect -11288 34338 -11273 34346
rect -11339 28370 -11322 28378
rect -11288 28370 -11273 28378
rect -11339 28358 -11273 28370
rect -11181 34346 -11115 34358
rect -11181 34338 -11164 34346
rect -11130 34338 -11115 34346
rect -11181 28370 -11164 28378
rect -11130 28370 -11115 28378
rect -11181 28358 -11115 28370
rect -11023 34346 -10957 34358
rect -11023 34338 -11006 34346
rect -10972 34338 -10957 34346
rect -11023 28370 -11006 28378
rect -10972 28370 -10957 28378
rect -11023 28358 -10957 28370
rect -10865 34346 -10799 34358
rect -10865 34338 -10848 34346
rect -10814 34338 -10799 34346
rect -10865 28370 -10848 28378
rect -10814 28370 -10799 28378
rect -10865 28358 -10799 28370
rect -10707 34346 -10641 34358
rect -10707 34338 -10690 34346
rect -10656 34338 -10641 34346
rect -10707 28370 -10690 28378
rect -10656 28370 -10641 28378
rect -10707 28358 -10641 28370
rect -10549 34346 -10483 34358
rect -10549 34338 -10532 34346
rect -10498 34338 -10483 34346
rect -10549 28370 -10532 28378
rect -10498 28370 -10483 28378
rect -10549 28358 -10483 28370
rect -10391 34346 -10325 34358
rect -10391 34338 -10374 34346
rect -10340 34338 -10325 34346
rect -10391 28370 -10374 28378
rect -10340 28370 -10325 28378
rect -10391 28358 -10325 28370
rect -10233 34346 -10167 34358
rect -10233 34338 -10216 34346
rect -10182 34338 -10167 34346
rect -10233 28370 -10216 28378
rect -10182 28370 -10167 28378
rect -10233 28358 -10167 28370
rect -10075 34346 -10009 34358
rect -10075 34338 -10058 34346
rect -10024 34338 -10009 34346
rect -10075 28370 -10058 28378
rect -10024 28370 -10009 28378
rect -10075 28358 -10009 28370
rect -9917 34346 -9851 34358
rect -9917 34338 -9900 34346
rect -9866 34338 -9851 34346
rect -9917 28370 -9900 28378
rect -9866 28370 -9851 28378
rect -9917 28358 -9851 28370
rect -9759 34346 -9693 34358
rect -9759 34338 -9742 34346
rect -9708 34338 -9693 34346
rect -9759 28370 -9742 28378
rect -9708 28370 -9693 28378
rect -9759 28358 -9693 28370
rect -9601 34346 -9535 34358
rect -9601 34338 -9584 34346
rect -9550 34338 -9535 34346
rect -9601 28370 -9584 28378
rect -9550 28370 -9535 28378
rect -9601 28358 -9535 28370
rect -9443 34346 -9377 34358
rect -9443 34338 -9426 34346
rect -9392 34338 -9377 34346
rect -9443 28370 -9426 28378
rect -9392 28370 -9377 28378
rect -9443 28358 -9377 28370
rect -9285 34346 -9219 34358
rect -9285 34338 -9268 34346
rect -9234 34338 -9219 34346
rect -9285 28370 -9268 28378
rect -9234 28370 -9219 28378
rect -9285 28358 -9219 28370
rect -9127 34346 -9061 34358
rect -9127 34338 -9110 34346
rect -9076 34338 -9061 34346
rect -9127 28370 -9110 28378
rect -9076 28370 -9061 28378
rect -9127 28358 -9061 28370
rect -8969 34346 -8903 34358
rect -8969 34338 -8952 34346
rect -8918 34338 -8903 34346
rect -8969 28370 -8952 28378
rect -8918 28370 -8903 28378
rect -8969 28358 -8903 28370
rect -8811 34346 -8745 34358
rect -8811 34338 -8794 34346
rect -8760 34338 -8745 34346
rect -8811 28370 -8794 28378
rect -8760 28370 -8745 28378
rect -8811 28358 -8745 28370
rect -8653 34346 -8587 34358
rect -8653 34338 -8636 34346
rect -8602 34338 -8587 34346
rect -8653 28370 -8636 28378
rect -8602 28370 -8587 28378
rect -8653 28358 -8587 28370
rect -8495 34346 -8429 34358
rect -8495 34338 -8478 34346
rect -8444 34338 -8429 34346
rect -8495 28370 -8478 28378
rect -8444 28370 -8429 28378
rect -8495 28358 -8429 28370
rect -13168 28320 -13148 28326
rect -8514 28320 -8494 28326
rect -13168 28286 -13156 28320
rect -8506 28286 -8494 28320
rect -13168 28226 -13148 28286
rect -8514 28226 -8494 28286
rect -13370 28194 -13300 28200
rect -8360 28194 -8290 28200
rect -13370 28184 -8290 28194
rect -13370 28146 -13164 28184
rect -8498 28146 -8290 28184
rect -13370 28130 -8290 28146
rect -7070 34570 -1990 34580
rect -7070 34532 -6864 34570
rect -2141 34532 -1990 34570
rect -7070 34522 -1990 34532
rect -7070 34520 -7000 34522
rect -2060 34520 -1990 34522
rect -6868 34430 -6848 34490
rect -2214 34430 -2194 34490
rect -6868 34396 -6856 34430
rect -2206 34396 -2194 34430
rect -6868 34390 -6848 34396
rect -2214 34390 -2194 34396
rect -6935 34346 -6869 34358
rect -6935 34338 -6918 34346
rect -6884 34338 -6869 34346
rect -6935 28370 -6918 28378
rect -6884 28370 -6869 28378
rect -6935 28358 -6869 28370
rect -6777 34346 -6711 34358
rect -6777 34338 -6760 34346
rect -6726 34338 -6711 34346
rect -6777 28370 -6760 28378
rect -6726 28370 -6711 28378
rect -6777 28358 -6711 28370
rect -6619 34346 -6553 34358
rect -6619 34338 -6602 34346
rect -6568 34338 -6553 34346
rect -6619 28370 -6602 28378
rect -6568 28370 -6553 28378
rect -6619 28358 -6553 28370
rect -6461 34346 -6395 34358
rect -6461 34338 -6444 34346
rect -6410 34338 -6395 34346
rect -6461 28370 -6444 28378
rect -6410 28370 -6395 28378
rect -6461 28358 -6395 28370
rect -6303 34346 -6237 34358
rect -6303 34338 -6286 34346
rect -6252 34338 -6237 34346
rect -6303 28370 -6286 28378
rect -6252 28370 -6237 28378
rect -6303 28358 -6237 28370
rect -6145 34346 -6079 34358
rect -6145 34338 -6128 34346
rect -6094 34338 -6079 34346
rect -6145 28370 -6128 28378
rect -6094 28370 -6079 28378
rect -6145 28358 -6079 28370
rect -5987 34346 -5921 34358
rect -5987 34338 -5970 34346
rect -5936 34338 -5921 34346
rect -5987 28370 -5970 28378
rect -5936 28370 -5921 28378
rect -5987 28358 -5921 28370
rect -5829 34346 -5763 34358
rect -5829 34338 -5812 34346
rect -5778 34338 -5763 34346
rect -5829 28370 -5812 28378
rect -5778 28370 -5763 28378
rect -5829 28358 -5763 28370
rect -5671 34346 -5605 34358
rect -5671 34338 -5654 34346
rect -5620 34338 -5605 34346
rect -5671 28370 -5654 28378
rect -5620 28370 -5605 28378
rect -5671 28358 -5605 28370
rect -5513 34346 -5447 34358
rect -5513 34338 -5496 34346
rect -5462 34338 -5447 34346
rect -5513 28370 -5496 28378
rect -5462 28370 -5447 28378
rect -5513 28358 -5447 28370
rect -5355 34346 -5289 34358
rect -5355 34338 -5338 34346
rect -5304 34338 -5289 34346
rect -5355 28370 -5338 28378
rect -5304 28370 -5289 28378
rect -5355 28358 -5289 28370
rect -5197 34346 -5131 34358
rect -5197 34338 -5180 34346
rect -5146 34338 -5131 34346
rect -5197 28370 -5180 28378
rect -5146 28370 -5131 28378
rect -5197 28358 -5131 28370
rect -5039 34346 -4973 34358
rect -5039 34338 -5022 34346
rect -4988 34338 -4973 34346
rect -5039 28370 -5022 28378
rect -4988 28370 -4973 28378
rect -5039 28358 -4973 28370
rect -4881 34346 -4815 34358
rect -4881 34338 -4864 34346
rect -4830 34338 -4815 34346
rect -4881 28370 -4864 28378
rect -4830 28370 -4815 28378
rect -4881 28358 -4815 28370
rect -4723 34346 -4657 34358
rect -4723 34338 -4706 34346
rect -4672 34338 -4657 34346
rect -4723 28370 -4706 28378
rect -4672 28370 -4657 28378
rect -4723 28358 -4657 28370
rect -4565 34346 -4499 34358
rect -4565 34338 -4548 34346
rect -4514 34338 -4499 34346
rect -4565 28370 -4548 28378
rect -4514 28370 -4499 28378
rect -4565 28358 -4499 28370
rect -4407 34346 -4341 34358
rect -4407 34338 -4390 34346
rect -4356 34338 -4341 34346
rect -4407 28370 -4390 28378
rect -4356 28370 -4341 28378
rect -4407 28358 -4341 28370
rect -4249 34346 -4183 34358
rect -4249 34338 -4232 34346
rect -4198 34338 -4183 34346
rect -4249 28370 -4232 28378
rect -4198 28370 -4183 28378
rect -4249 28358 -4183 28370
rect -4091 34346 -4025 34358
rect -4091 34338 -4074 34346
rect -4040 34338 -4025 34346
rect -4091 28370 -4074 28378
rect -4040 28370 -4025 28378
rect -4091 28358 -4025 28370
rect -3933 34346 -3867 34358
rect -3933 34338 -3916 34346
rect -3882 34338 -3867 34346
rect -3933 28370 -3916 28378
rect -3882 28370 -3867 28378
rect -3933 28358 -3867 28370
rect -3775 34346 -3709 34358
rect -3775 34338 -3758 34346
rect -3724 34338 -3709 34346
rect -3775 28370 -3758 28378
rect -3724 28370 -3709 28378
rect -3775 28358 -3709 28370
rect -3617 34346 -3551 34358
rect -3617 34338 -3600 34346
rect -3566 34338 -3551 34346
rect -3617 28370 -3600 28378
rect -3566 28370 -3551 28378
rect -3617 28358 -3551 28370
rect -3459 34346 -3393 34358
rect -3459 34338 -3442 34346
rect -3408 34338 -3393 34346
rect -3459 28370 -3442 28378
rect -3408 28370 -3393 28378
rect -3459 28358 -3393 28370
rect -3301 34346 -3235 34358
rect -3301 34338 -3284 34346
rect -3250 34338 -3235 34346
rect -3301 28370 -3284 28378
rect -3250 28370 -3235 28378
rect -3301 28358 -3235 28370
rect -3143 34346 -3077 34358
rect -3143 34338 -3126 34346
rect -3092 34338 -3077 34346
rect -3143 28370 -3126 28378
rect -3092 28370 -3077 28378
rect -3143 28358 -3077 28370
rect -2985 34346 -2919 34358
rect -2985 34338 -2968 34346
rect -2934 34338 -2919 34346
rect -2985 28370 -2968 28378
rect -2934 28370 -2919 28378
rect -2985 28358 -2919 28370
rect -2827 34346 -2761 34358
rect -2827 34338 -2810 34346
rect -2776 34338 -2761 34346
rect -2827 28370 -2810 28378
rect -2776 28370 -2761 28378
rect -2827 28358 -2761 28370
rect -2669 34346 -2603 34358
rect -2669 34338 -2652 34346
rect -2618 34338 -2603 34346
rect -2669 28370 -2652 28378
rect -2618 28370 -2603 28378
rect -2669 28358 -2603 28370
rect -2511 34346 -2445 34358
rect -2511 34338 -2494 34346
rect -2460 34338 -2445 34346
rect -2511 28370 -2494 28378
rect -2460 28370 -2445 28378
rect -2511 28358 -2445 28370
rect -2353 34346 -2287 34358
rect -2353 34338 -2336 34346
rect -2302 34338 -2287 34346
rect -2353 28370 -2336 28378
rect -2302 28370 -2287 28378
rect -2353 28358 -2287 28370
rect -2195 34346 -2129 34358
rect -2195 34338 -2178 34346
rect -2144 34338 -2129 34346
rect -2195 28370 -2178 28378
rect -2144 28370 -2129 28378
rect -2195 28358 -2129 28370
rect -6868 28320 -6848 28326
rect -2214 28320 -2194 28326
rect -6868 28286 -6856 28320
rect -2206 28286 -2194 28320
rect -6868 28226 -6848 28286
rect -2214 28226 -2194 28286
rect -7070 28194 -7000 28200
rect -2060 28194 -1990 28200
rect -7070 28184 -1990 28194
rect -7070 28146 -6864 28184
rect -2198 28146 -1990 28184
rect -7070 28130 -1990 28146
rect -770 34570 4310 34580
rect -770 34532 -564 34570
rect 4159 34532 4310 34570
rect -770 34522 4310 34532
rect -770 34520 -700 34522
rect 4240 34520 4310 34522
rect -568 34430 -548 34490
rect 4086 34430 4106 34490
rect -568 34396 -556 34430
rect 4094 34396 4106 34430
rect -568 34390 -548 34396
rect 4086 34390 4106 34396
rect -635 34346 -569 34358
rect -635 34338 -618 34346
rect -584 34338 -569 34346
rect -635 28370 -618 28378
rect -584 28370 -569 28378
rect -635 28358 -569 28370
rect -477 34346 -411 34358
rect -477 34338 -460 34346
rect -426 34338 -411 34346
rect -477 28370 -460 28378
rect -426 28370 -411 28378
rect -477 28358 -411 28370
rect -319 34346 -253 34358
rect -319 34338 -302 34346
rect -268 34338 -253 34346
rect -319 28370 -302 28378
rect -268 28370 -253 28378
rect -319 28358 -253 28370
rect -161 34346 -95 34358
rect -161 34338 -144 34346
rect -110 34338 -95 34346
rect -161 28370 -144 28378
rect -110 28370 -95 28378
rect -161 28358 -95 28370
rect -3 34346 63 34358
rect -3 34338 14 34346
rect 48 34338 63 34346
rect -3 28370 14 28378
rect 48 28370 63 28378
rect -3 28358 63 28370
rect 155 34346 221 34358
rect 155 34338 172 34346
rect 206 34338 221 34346
rect 155 28370 172 28378
rect 206 28370 221 28378
rect 155 28358 221 28370
rect 313 34346 379 34358
rect 313 34338 330 34346
rect 364 34338 379 34346
rect 313 28370 330 28378
rect 364 28370 379 28378
rect 313 28358 379 28370
rect 471 34346 537 34358
rect 471 34338 488 34346
rect 522 34338 537 34346
rect 471 28370 488 28378
rect 522 28370 537 28378
rect 471 28358 537 28370
rect 629 34346 695 34358
rect 629 34338 646 34346
rect 680 34338 695 34346
rect 629 28370 646 28378
rect 680 28370 695 28378
rect 629 28358 695 28370
rect 787 34346 853 34358
rect 787 34338 804 34346
rect 838 34338 853 34346
rect 787 28370 804 28378
rect 838 28370 853 28378
rect 787 28358 853 28370
rect 945 34346 1011 34358
rect 945 34338 962 34346
rect 996 34338 1011 34346
rect 945 28370 962 28378
rect 996 28370 1011 28378
rect 945 28358 1011 28370
rect 1103 34346 1169 34358
rect 1103 34338 1120 34346
rect 1154 34338 1169 34346
rect 1103 28370 1120 28378
rect 1154 28370 1169 28378
rect 1103 28358 1169 28370
rect 1261 34346 1327 34358
rect 1261 34338 1278 34346
rect 1312 34338 1327 34346
rect 1261 28370 1278 28378
rect 1312 28370 1327 28378
rect 1261 28358 1327 28370
rect 1419 34346 1485 34358
rect 1419 34338 1436 34346
rect 1470 34338 1485 34346
rect 1419 28370 1436 28378
rect 1470 28370 1485 28378
rect 1419 28358 1485 28370
rect 1577 34346 1643 34358
rect 1577 34338 1594 34346
rect 1628 34338 1643 34346
rect 1577 28370 1594 28378
rect 1628 28370 1643 28378
rect 1577 28358 1643 28370
rect 1735 34346 1801 34358
rect 1735 34338 1752 34346
rect 1786 34338 1801 34346
rect 1735 28370 1752 28378
rect 1786 28370 1801 28378
rect 1735 28358 1801 28370
rect 1893 34346 1959 34358
rect 1893 34338 1910 34346
rect 1944 34338 1959 34346
rect 1893 28370 1910 28378
rect 1944 28370 1959 28378
rect 1893 28358 1959 28370
rect 2051 34346 2117 34358
rect 2051 34338 2068 34346
rect 2102 34338 2117 34346
rect 2051 28370 2068 28378
rect 2102 28370 2117 28378
rect 2051 28358 2117 28370
rect 2209 34346 2275 34358
rect 2209 34338 2226 34346
rect 2260 34338 2275 34346
rect 2209 28370 2226 28378
rect 2260 28370 2275 28378
rect 2209 28358 2275 28370
rect 2367 34346 2433 34358
rect 2367 34338 2384 34346
rect 2418 34338 2433 34346
rect 2367 28370 2384 28378
rect 2418 28370 2433 28378
rect 2367 28358 2433 28370
rect 2525 34346 2591 34358
rect 2525 34338 2542 34346
rect 2576 34338 2591 34346
rect 2525 28370 2542 28378
rect 2576 28370 2591 28378
rect 2525 28358 2591 28370
rect 2683 34346 2749 34358
rect 2683 34338 2700 34346
rect 2734 34338 2749 34346
rect 2683 28370 2700 28378
rect 2734 28370 2749 28378
rect 2683 28358 2749 28370
rect 2841 34346 2907 34358
rect 2841 34338 2858 34346
rect 2892 34338 2907 34346
rect 2841 28370 2858 28378
rect 2892 28370 2907 28378
rect 2841 28358 2907 28370
rect 2999 34346 3065 34358
rect 2999 34338 3016 34346
rect 3050 34338 3065 34346
rect 2999 28370 3016 28378
rect 3050 28370 3065 28378
rect 2999 28358 3065 28370
rect 3157 34346 3223 34358
rect 3157 34338 3174 34346
rect 3208 34338 3223 34346
rect 3157 28370 3174 28378
rect 3208 28370 3223 28378
rect 3157 28358 3223 28370
rect 3315 34346 3381 34358
rect 3315 34338 3332 34346
rect 3366 34338 3381 34346
rect 3315 28370 3332 28378
rect 3366 28370 3381 28378
rect 3315 28358 3381 28370
rect 3473 34346 3539 34358
rect 3473 34338 3490 34346
rect 3524 34338 3539 34346
rect 3473 28370 3490 28378
rect 3524 28370 3539 28378
rect 3473 28358 3539 28370
rect 3631 34346 3697 34358
rect 3631 34338 3648 34346
rect 3682 34338 3697 34346
rect 3631 28370 3648 28378
rect 3682 28370 3697 28378
rect 3631 28358 3697 28370
rect 3789 34346 3855 34358
rect 3789 34338 3806 34346
rect 3840 34338 3855 34346
rect 3789 28370 3806 28378
rect 3840 28370 3855 28378
rect 3789 28358 3855 28370
rect 3947 34346 4013 34358
rect 3947 34338 3964 34346
rect 3998 34338 4013 34346
rect 3947 28370 3964 28378
rect 3998 28370 4013 28378
rect 3947 28358 4013 28370
rect 4105 34346 4171 34358
rect 4105 34338 4122 34346
rect 4156 34338 4171 34346
rect 4105 28370 4122 28378
rect 4156 28370 4171 28378
rect 4105 28358 4171 28370
rect -568 28320 -548 28326
rect 4086 28320 4106 28326
rect -568 28286 -556 28320
rect 4094 28286 4106 28320
rect -568 28226 -548 28286
rect 4086 28226 4106 28286
rect -770 28194 -700 28200
rect 4240 28194 4310 28200
rect -770 28184 4310 28194
rect -770 28146 -564 28184
rect 4102 28146 4310 28184
rect -770 28130 4310 28146
rect 5530 34570 10610 34580
rect 5530 34532 5736 34570
rect 10459 34532 10610 34570
rect 5530 34522 10610 34532
rect 5530 34520 5600 34522
rect 10540 34520 10610 34522
rect 5732 34430 5752 34490
rect 10386 34430 10406 34490
rect 5732 34396 5744 34430
rect 10394 34396 10406 34430
rect 5732 34390 5752 34396
rect 10386 34390 10406 34396
rect 5665 34346 5731 34358
rect 5665 34338 5682 34346
rect 5716 34338 5731 34346
rect 5665 28370 5682 28378
rect 5716 28370 5731 28378
rect 5665 28358 5731 28370
rect 5823 34346 5889 34358
rect 5823 34338 5840 34346
rect 5874 34338 5889 34346
rect 5823 28370 5840 28378
rect 5874 28370 5889 28378
rect 5823 28358 5889 28370
rect 5981 34346 6047 34358
rect 5981 34338 5998 34346
rect 6032 34338 6047 34346
rect 5981 28370 5998 28378
rect 6032 28370 6047 28378
rect 5981 28358 6047 28370
rect 6139 34346 6205 34358
rect 6139 34338 6156 34346
rect 6190 34338 6205 34346
rect 6139 28370 6156 28378
rect 6190 28370 6205 28378
rect 6139 28358 6205 28370
rect 6297 34346 6363 34358
rect 6297 34338 6314 34346
rect 6348 34338 6363 34346
rect 6297 28370 6314 28378
rect 6348 28370 6363 28378
rect 6297 28358 6363 28370
rect 6455 34346 6521 34358
rect 6455 34338 6472 34346
rect 6506 34338 6521 34346
rect 6455 28370 6472 28378
rect 6506 28370 6521 28378
rect 6455 28358 6521 28370
rect 6613 34346 6679 34358
rect 6613 34338 6630 34346
rect 6664 34338 6679 34346
rect 6613 28370 6630 28378
rect 6664 28370 6679 28378
rect 6613 28358 6679 28370
rect 6771 34346 6837 34358
rect 6771 34338 6788 34346
rect 6822 34338 6837 34346
rect 6771 28370 6788 28378
rect 6822 28370 6837 28378
rect 6771 28358 6837 28370
rect 6929 34346 6995 34358
rect 6929 34338 6946 34346
rect 6980 34338 6995 34346
rect 6929 28370 6946 28378
rect 6980 28370 6995 28378
rect 6929 28358 6995 28370
rect 7087 34346 7153 34358
rect 7087 34338 7104 34346
rect 7138 34338 7153 34346
rect 7087 28370 7104 28378
rect 7138 28370 7153 28378
rect 7087 28358 7153 28370
rect 7245 34346 7311 34358
rect 7245 34338 7262 34346
rect 7296 34338 7311 34346
rect 7245 28370 7262 28378
rect 7296 28370 7311 28378
rect 7245 28358 7311 28370
rect 7403 34346 7469 34358
rect 7403 34338 7420 34346
rect 7454 34338 7469 34346
rect 7403 28370 7420 28378
rect 7454 28370 7469 28378
rect 7403 28358 7469 28370
rect 7561 34346 7627 34358
rect 7561 34338 7578 34346
rect 7612 34338 7627 34346
rect 7561 28370 7578 28378
rect 7612 28370 7627 28378
rect 7561 28358 7627 28370
rect 7719 34346 7785 34358
rect 7719 34338 7736 34346
rect 7770 34338 7785 34346
rect 7719 28370 7736 28378
rect 7770 28370 7785 28378
rect 7719 28358 7785 28370
rect 7877 34346 7943 34358
rect 7877 34338 7894 34346
rect 7928 34338 7943 34346
rect 7877 28370 7894 28378
rect 7928 28370 7943 28378
rect 7877 28358 7943 28370
rect 8035 34346 8101 34358
rect 8035 34338 8052 34346
rect 8086 34338 8101 34346
rect 8035 28370 8052 28378
rect 8086 28370 8101 28378
rect 8035 28358 8101 28370
rect 8193 34346 8259 34358
rect 8193 34338 8210 34346
rect 8244 34338 8259 34346
rect 8193 28370 8210 28378
rect 8244 28370 8259 28378
rect 8193 28358 8259 28370
rect 8351 34346 8417 34358
rect 8351 34338 8368 34346
rect 8402 34338 8417 34346
rect 8351 28370 8368 28378
rect 8402 28370 8417 28378
rect 8351 28358 8417 28370
rect 8509 34346 8575 34358
rect 8509 34338 8526 34346
rect 8560 34338 8575 34346
rect 8509 28370 8526 28378
rect 8560 28370 8575 28378
rect 8509 28358 8575 28370
rect 8667 34346 8733 34358
rect 8667 34338 8684 34346
rect 8718 34338 8733 34346
rect 8667 28370 8684 28378
rect 8718 28370 8733 28378
rect 8667 28358 8733 28370
rect 8825 34346 8891 34358
rect 8825 34338 8842 34346
rect 8876 34338 8891 34346
rect 8825 28370 8842 28378
rect 8876 28370 8891 28378
rect 8825 28358 8891 28370
rect 8983 34346 9049 34358
rect 8983 34338 9000 34346
rect 9034 34338 9049 34346
rect 8983 28370 9000 28378
rect 9034 28370 9049 28378
rect 8983 28358 9049 28370
rect 9141 34346 9207 34358
rect 9141 34338 9158 34346
rect 9192 34338 9207 34346
rect 9141 28370 9158 28378
rect 9192 28370 9207 28378
rect 9141 28358 9207 28370
rect 9299 34346 9365 34358
rect 9299 34338 9316 34346
rect 9350 34338 9365 34346
rect 9299 28370 9316 28378
rect 9350 28370 9365 28378
rect 9299 28358 9365 28370
rect 9457 34346 9523 34358
rect 9457 34338 9474 34346
rect 9508 34338 9523 34346
rect 9457 28370 9474 28378
rect 9508 28370 9523 28378
rect 9457 28358 9523 28370
rect 9615 34346 9681 34358
rect 9615 34338 9632 34346
rect 9666 34338 9681 34346
rect 9615 28370 9632 28378
rect 9666 28370 9681 28378
rect 9615 28358 9681 28370
rect 9773 34346 9839 34358
rect 9773 34338 9790 34346
rect 9824 34338 9839 34346
rect 9773 28370 9790 28378
rect 9824 28370 9839 28378
rect 9773 28358 9839 28370
rect 9931 34346 9997 34358
rect 9931 34338 9948 34346
rect 9982 34338 9997 34346
rect 9931 28370 9948 28378
rect 9982 28370 9997 28378
rect 9931 28358 9997 28370
rect 10089 34346 10155 34358
rect 10089 34338 10106 34346
rect 10140 34338 10155 34346
rect 10089 28370 10106 28378
rect 10140 28370 10155 28378
rect 10089 28358 10155 28370
rect 10247 34346 10313 34358
rect 10247 34338 10264 34346
rect 10298 34338 10313 34346
rect 10247 28370 10264 28378
rect 10298 28370 10313 28378
rect 10247 28358 10313 28370
rect 10405 34346 10471 34358
rect 10405 34338 10422 34346
rect 10456 34338 10471 34346
rect 10405 28370 10422 28378
rect 10456 28370 10471 28378
rect 10405 28358 10471 28370
rect 5732 28320 5752 28326
rect 10386 28320 10406 28326
rect 5732 28286 5744 28320
rect 10394 28286 10406 28320
rect 5732 28226 5752 28286
rect 10386 28226 10406 28286
rect 5530 28194 5600 28200
rect 10540 28194 10610 28200
rect 5530 28184 10610 28194
rect 5530 28146 5736 28184
rect 10402 28146 10610 28184
rect 5530 28130 10610 28146
rect -13370 27570 -8290 27580
rect -13370 27532 -13164 27570
rect -8441 27532 -8290 27570
rect -13370 27522 -8290 27532
rect -13370 27520 -13300 27522
rect -8360 27520 -8290 27522
rect -13168 27430 -13148 27490
rect -8514 27430 -8494 27490
rect -13168 27396 -13156 27430
rect -8506 27396 -8494 27430
rect -13168 27390 -13148 27396
rect -8514 27390 -8494 27396
rect -13235 27346 -13169 27358
rect -13235 27338 -13218 27346
rect -13184 27338 -13169 27346
rect -13235 21370 -13218 21378
rect -13184 21370 -13169 21378
rect -13235 21358 -13169 21370
rect -13077 27346 -13011 27358
rect -13077 27338 -13060 27346
rect -13026 27338 -13011 27346
rect -13077 21370 -13060 21378
rect -13026 21370 -13011 21378
rect -13077 21358 -13011 21370
rect -12919 27346 -12853 27358
rect -12919 27338 -12902 27346
rect -12868 27338 -12853 27346
rect -12919 21370 -12902 21378
rect -12868 21370 -12853 21378
rect -12919 21358 -12853 21370
rect -12761 27346 -12695 27358
rect -12761 27338 -12744 27346
rect -12710 27338 -12695 27346
rect -12761 21370 -12744 21378
rect -12710 21370 -12695 21378
rect -12761 21358 -12695 21370
rect -12603 27346 -12537 27358
rect -12603 27338 -12586 27346
rect -12552 27338 -12537 27346
rect -12603 21370 -12586 21378
rect -12552 21370 -12537 21378
rect -12603 21358 -12537 21370
rect -12445 27346 -12379 27358
rect -12445 27338 -12428 27346
rect -12394 27338 -12379 27346
rect -12445 21370 -12428 21378
rect -12394 21370 -12379 21378
rect -12445 21358 -12379 21370
rect -12287 27346 -12221 27358
rect -12287 27338 -12270 27346
rect -12236 27338 -12221 27346
rect -12287 21370 -12270 21378
rect -12236 21370 -12221 21378
rect -12287 21358 -12221 21370
rect -12129 27346 -12063 27358
rect -12129 27338 -12112 27346
rect -12078 27338 -12063 27346
rect -12129 21370 -12112 21378
rect -12078 21370 -12063 21378
rect -12129 21358 -12063 21370
rect -11971 27346 -11905 27358
rect -11971 27338 -11954 27346
rect -11920 27338 -11905 27346
rect -11971 21370 -11954 21378
rect -11920 21370 -11905 21378
rect -11971 21358 -11905 21370
rect -11813 27346 -11747 27358
rect -11813 27338 -11796 27346
rect -11762 27338 -11747 27346
rect -11813 21370 -11796 21378
rect -11762 21370 -11747 21378
rect -11813 21358 -11747 21370
rect -11655 27346 -11589 27358
rect -11655 27338 -11638 27346
rect -11604 27338 -11589 27346
rect -11655 21370 -11638 21378
rect -11604 21370 -11589 21378
rect -11655 21358 -11589 21370
rect -11497 27346 -11431 27358
rect -11497 27338 -11480 27346
rect -11446 27338 -11431 27346
rect -11497 21370 -11480 21378
rect -11446 21370 -11431 21378
rect -11497 21358 -11431 21370
rect -11339 27346 -11273 27358
rect -11339 27338 -11322 27346
rect -11288 27338 -11273 27346
rect -11339 21370 -11322 21378
rect -11288 21370 -11273 21378
rect -11339 21358 -11273 21370
rect -11181 27346 -11115 27358
rect -11181 27338 -11164 27346
rect -11130 27338 -11115 27346
rect -11181 21370 -11164 21378
rect -11130 21370 -11115 21378
rect -11181 21358 -11115 21370
rect -11023 27346 -10957 27358
rect -11023 27338 -11006 27346
rect -10972 27338 -10957 27346
rect -11023 21370 -11006 21378
rect -10972 21370 -10957 21378
rect -11023 21358 -10957 21370
rect -10865 27346 -10799 27358
rect -10865 27338 -10848 27346
rect -10814 27338 -10799 27346
rect -10865 21370 -10848 21378
rect -10814 21370 -10799 21378
rect -10865 21358 -10799 21370
rect -10707 27346 -10641 27358
rect -10707 27338 -10690 27346
rect -10656 27338 -10641 27346
rect -10707 21370 -10690 21378
rect -10656 21370 -10641 21378
rect -10707 21358 -10641 21370
rect -10549 27346 -10483 27358
rect -10549 27338 -10532 27346
rect -10498 27338 -10483 27346
rect -10549 21370 -10532 21378
rect -10498 21370 -10483 21378
rect -10549 21358 -10483 21370
rect -10391 27346 -10325 27358
rect -10391 27338 -10374 27346
rect -10340 27338 -10325 27346
rect -10391 21370 -10374 21378
rect -10340 21370 -10325 21378
rect -10391 21358 -10325 21370
rect -10233 27346 -10167 27358
rect -10233 27338 -10216 27346
rect -10182 27338 -10167 27346
rect -10233 21370 -10216 21378
rect -10182 21370 -10167 21378
rect -10233 21358 -10167 21370
rect -10075 27346 -10009 27358
rect -10075 27338 -10058 27346
rect -10024 27338 -10009 27346
rect -10075 21370 -10058 21378
rect -10024 21370 -10009 21378
rect -10075 21358 -10009 21370
rect -9917 27346 -9851 27358
rect -9917 27338 -9900 27346
rect -9866 27338 -9851 27346
rect -9917 21370 -9900 21378
rect -9866 21370 -9851 21378
rect -9917 21358 -9851 21370
rect -9759 27346 -9693 27358
rect -9759 27338 -9742 27346
rect -9708 27338 -9693 27346
rect -9759 21370 -9742 21378
rect -9708 21370 -9693 21378
rect -9759 21358 -9693 21370
rect -9601 27346 -9535 27358
rect -9601 27338 -9584 27346
rect -9550 27338 -9535 27346
rect -9601 21370 -9584 21378
rect -9550 21370 -9535 21378
rect -9601 21358 -9535 21370
rect -9443 27346 -9377 27358
rect -9443 27338 -9426 27346
rect -9392 27338 -9377 27346
rect -9443 21370 -9426 21378
rect -9392 21370 -9377 21378
rect -9443 21358 -9377 21370
rect -9285 27346 -9219 27358
rect -9285 27338 -9268 27346
rect -9234 27338 -9219 27346
rect -9285 21370 -9268 21378
rect -9234 21370 -9219 21378
rect -9285 21358 -9219 21370
rect -9127 27346 -9061 27358
rect -9127 27338 -9110 27346
rect -9076 27338 -9061 27346
rect -9127 21370 -9110 21378
rect -9076 21370 -9061 21378
rect -9127 21358 -9061 21370
rect -8969 27346 -8903 27358
rect -8969 27338 -8952 27346
rect -8918 27338 -8903 27346
rect -8969 21370 -8952 21378
rect -8918 21370 -8903 21378
rect -8969 21358 -8903 21370
rect -8811 27346 -8745 27358
rect -8811 27338 -8794 27346
rect -8760 27338 -8745 27346
rect -8811 21370 -8794 21378
rect -8760 21370 -8745 21378
rect -8811 21358 -8745 21370
rect -8653 27346 -8587 27358
rect -8653 27338 -8636 27346
rect -8602 27338 -8587 27346
rect -8653 21370 -8636 21378
rect -8602 21370 -8587 21378
rect -8653 21358 -8587 21370
rect -8495 27346 -8429 27358
rect -8495 27338 -8478 27346
rect -8444 27338 -8429 27346
rect -8495 21370 -8478 21378
rect -8444 21370 -8429 21378
rect -8495 21358 -8429 21370
rect -13168 21320 -13148 21326
rect -8514 21320 -8494 21326
rect -13168 21286 -13156 21320
rect -8506 21286 -8494 21320
rect -13168 21226 -13148 21286
rect -8514 21226 -8494 21286
rect -13370 21194 -13300 21200
rect -8360 21194 -8290 21200
rect -13370 21184 -8290 21194
rect -13370 21146 -13164 21184
rect -8498 21146 -8290 21184
rect -13370 21130 -8290 21146
rect -7070 27570 -1990 27580
rect -7070 27532 -6864 27570
rect -2141 27532 -1990 27570
rect -7070 27522 -1990 27532
rect -7070 27520 -7000 27522
rect -2060 27520 -1990 27522
rect -6868 27430 -6848 27490
rect -2214 27430 -2194 27490
rect -6868 27396 -6856 27430
rect -2206 27396 -2194 27430
rect -6868 27390 -6848 27396
rect -2214 27390 -2194 27396
rect -6935 27346 -6869 27358
rect -6935 27338 -6918 27346
rect -6884 27338 -6869 27346
rect -6935 21370 -6918 21378
rect -6884 21370 -6869 21378
rect -6935 21358 -6869 21370
rect -6777 27346 -6711 27358
rect -6777 27338 -6760 27346
rect -6726 27338 -6711 27346
rect -6777 21370 -6760 21378
rect -6726 21370 -6711 21378
rect -6777 21358 -6711 21370
rect -6619 27346 -6553 27358
rect -6619 27338 -6602 27346
rect -6568 27338 -6553 27346
rect -6619 21370 -6602 21378
rect -6568 21370 -6553 21378
rect -6619 21358 -6553 21370
rect -6461 27346 -6395 27358
rect -6461 27338 -6444 27346
rect -6410 27338 -6395 27346
rect -6461 21370 -6444 21378
rect -6410 21370 -6395 21378
rect -6461 21358 -6395 21370
rect -6303 27346 -6237 27358
rect -6303 27338 -6286 27346
rect -6252 27338 -6237 27346
rect -6303 21370 -6286 21378
rect -6252 21370 -6237 21378
rect -6303 21358 -6237 21370
rect -6145 27346 -6079 27358
rect -6145 27338 -6128 27346
rect -6094 27338 -6079 27346
rect -6145 21370 -6128 21378
rect -6094 21370 -6079 21378
rect -6145 21358 -6079 21370
rect -5987 27346 -5921 27358
rect -5987 27338 -5970 27346
rect -5936 27338 -5921 27346
rect -5987 21370 -5970 21378
rect -5936 21370 -5921 21378
rect -5987 21358 -5921 21370
rect -5829 27346 -5763 27358
rect -5829 27338 -5812 27346
rect -5778 27338 -5763 27346
rect -5829 21370 -5812 21378
rect -5778 21370 -5763 21378
rect -5829 21358 -5763 21370
rect -5671 27346 -5605 27358
rect -5671 27338 -5654 27346
rect -5620 27338 -5605 27346
rect -5671 21370 -5654 21378
rect -5620 21370 -5605 21378
rect -5671 21358 -5605 21370
rect -5513 27346 -5447 27358
rect -5513 27338 -5496 27346
rect -5462 27338 -5447 27346
rect -5513 21370 -5496 21378
rect -5462 21370 -5447 21378
rect -5513 21358 -5447 21370
rect -5355 27346 -5289 27358
rect -5355 27338 -5338 27346
rect -5304 27338 -5289 27346
rect -5355 21370 -5338 21378
rect -5304 21370 -5289 21378
rect -5355 21358 -5289 21370
rect -5197 27346 -5131 27358
rect -5197 27338 -5180 27346
rect -5146 27338 -5131 27346
rect -5197 21370 -5180 21378
rect -5146 21370 -5131 21378
rect -5197 21358 -5131 21370
rect -5039 27346 -4973 27358
rect -5039 27338 -5022 27346
rect -4988 27338 -4973 27346
rect -5039 21370 -5022 21378
rect -4988 21370 -4973 21378
rect -5039 21358 -4973 21370
rect -4881 27346 -4815 27358
rect -4881 27338 -4864 27346
rect -4830 27338 -4815 27346
rect -4881 21370 -4864 21378
rect -4830 21370 -4815 21378
rect -4881 21358 -4815 21370
rect -4723 27346 -4657 27358
rect -4723 27338 -4706 27346
rect -4672 27338 -4657 27346
rect -4723 21370 -4706 21378
rect -4672 21370 -4657 21378
rect -4723 21358 -4657 21370
rect -4565 27346 -4499 27358
rect -4565 27338 -4548 27346
rect -4514 27338 -4499 27346
rect -4565 21370 -4548 21378
rect -4514 21370 -4499 21378
rect -4565 21358 -4499 21370
rect -4407 27346 -4341 27358
rect -4407 27338 -4390 27346
rect -4356 27338 -4341 27346
rect -4407 21370 -4390 21378
rect -4356 21370 -4341 21378
rect -4407 21358 -4341 21370
rect -4249 27346 -4183 27358
rect -4249 27338 -4232 27346
rect -4198 27338 -4183 27346
rect -4249 21370 -4232 21378
rect -4198 21370 -4183 21378
rect -4249 21358 -4183 21370
rect -4091 27346 -4025 27358
rect -4091 27338 -4074 27346
rect -4040 27338 -4025 27346
rect -4091 21370 -4074 21378
rect -4040 21370 -4025 21378
rect -4091 21358 -4025 21370
rect -3933 27346 -3867 27358
rect -3933 27338 -3916 27346
rect -3882 27338 -3867 27346
rect -3933 21370 -3916 21378
rect -3882 21370 -3867 21378
rect -3933 21358 -3867 21370
rect -3775 27346 -3709 27358
rect -3775 27338 -3758 27346
rect -3724 27338 -3709 27346
rect -3775 21370 -3758 21378
rect -3724 21370 -3709 21378
rect -3775 21358 -3709 21370
rect -3617 27346 -3551 27358
rect -3617 27338 -3600 27346
rect -3566 27338 -3551 27346
rect -3617 21370 -3600 21378
rect -3566 21370 -3551 21378
rect -3617 21358 -3551 21370
rect -3459 27346 -3393 27358
rect -3459 27338 -3442 27346
rect -3408 27338 -3393 27346
rect -3459 21370 -3442 21378
rect -3408 21370 -3393 21378
rect -3459 21358 -3393 21370
rect -3301 27346 -3235 27358
rect -3301 27338 -3284 27346
rect -3250 27338 -3235 27346
rect -3301 21370 -3284 21378
rect -3250 21370 -3235 21378
rect -3301 21358 -3235 21370
rect -3143 27346 -3077 27358
rect -3143 27338 -3126 27346
rect -3092 27338 -3077 27346
rect -3143 21370 -3126 21378
rect -3092 21370 -3077 21378
rect -3143 21358 -3077 21370
rect -2985 27346 -2919 27358
rect -2985 27338 -2968 27346
rect -2934 27338 -2919 27346
rect -2985 21370 -2968 21378
rect -2934 21370 -2919 21378
rect -2985 21358 -2919 21370
rect -2827 27346 -2761 27358
rect -2827 27338 -2810 27346
rect -2776 27338 -2761 27346
rect -2827 21370 -2810 21378
rect -2776 21370 -2761 21378
rect -2827 21358 -2761 21370
rect -2669 27346 -2603 27358
rect -2669 27338 -2652 27346
rect -2618 27338 -2603 27346
rect -2669 21370 -2652 21378
rect -2618 21370 -2603 21378
rect -2669 21358 -2603 21370
rect -2511 27346 -2445 27358
rect -2511 27338 -2494 27346
rect -2460 27338 -2445 27346
rect -2511 21370 -2494 21378
rect -2460 21370 -2445 21378
rect -2511 21358 -2445 21370
rect -2353 27346 -2287 27358
rect -2353 27338 -2336 27346
rect -2302 27338 -2287 27346
rect -2353 21370 -2336 21378
rect -2302 21370 -2287 21378
rect -2353 21358 -2287 21370
rect -2195 27346 -2129 27358
rect -2195 27338 -2178 27346
rect -2144 27338 -2129 27346
rect -2195 21370 -2178 21378
rect -2144 21370 -2129 21378
rect -2195 21358 -2129 21370
rect -6868 21320 -6848 21326
rect -2214 21320 -2194 21326
rect -6868 21286 -6856 21320
rect -2206 21286 -2194 21320
rect -6868 21226 -6848 21286
rect -2214 21226 -2194 21286
rect -7070 21194 -7000 21200
rect -2060 21194 -1990 21200
rect -7070 21184 -1990 21194
rect -7070 21146 -6864 21184
rect -2198 21146 -1990 21184
rect -7070 21130 -1990 21146
rect -770 27570 4310 27580
rect -770 27532 -564 27570
rect 4159 27532 4310 27570
rect -770 27522 4310 27532
rect -770 27520 -700 27522
rect 4240 27520 4310 27522
rect -568 27430 -548 27490
rect 4086 27430 4106 27490
rect -568 27396 -556 27430
rect 4094 27396 4106 27430
rect -568 27390 -548 27396
rect 4086 27390 4106 27396
rect -635 27346 -569 27358
rect -635 27338 -618 27346
rect -584 27338 -569 27346
rect -635 21370 -618 21378
rect -584 21370 -569 21378
rect -635 21358 -569 21370
rect -477 27346 -411 27358
rect -477 27338 -460 27346
rect -426 27338 -411 27346
rect -477 21370 -460 21378
rect -426 21370 -411 21378
rect -477 21358 -411 21370
rect -319 27346 -253 27358
rect -319 27338 -302 27346
rect -268 27338 -253 27346
rect -319 21370 -302 21378
rect -268 21370 -253 21378
rect -319 21358 -253 21370
rect -161 27346 -95 27358
rect -161 27338 -144 27346
rect -110 27338 -95 27346
rect -161 21370 -144 21378
rect -110 21370 -95 21378
rect -161 21358 -95 21370
rect -3 27346 63 27358
rect -3 27338 14 27346
rect 48 27338 63 27346
rect -3 21370 14 21378
rect 48 21370 63 21378
rect -3 21358 63 21370
rect 155 27346 221 27358
rect 155 27338 172 27346
rect 206 27338 221 27346
rect 155 21370 172 21378
rect 206 21370 221 21378
rect 155 21358 221 21370
rect 313 27346 379 27358
rect 313 27338 330 27346
rect 364 27338 379 27346
rect 313 21370 330 21378
rect 364 21370 379 21378
rect 313 21358 379 21370
rect 471 27346 537 27358
rect 471 27338 488 27346
rect 522 27338 537 27346
rect 471 21370 488 21378
rect 522 21370 537 21378
rect 471 21358 537 21370
rect 629 27346 695 27358
rect 629 27338 646 27346
rect 680 27338 695 27346
rect 629 21370 646 21378
rect 680 21370 695 21378
rect 629 21358 695 21370
rect 787 27346 853 27358
rect 787 27338 804 27346
rect 838 27338 853 27346
rect 787 21370 804 21378
rect 838 21370 853 21378
rect 787 21358 853 21370
rect 945 27346 1011 27358
rect 945 27338 962 27346
rect 996 27338 1011 27346
rect 945 21370 962 21378
rect 996 21370 1011 21378
rect 945 21358 1011 21370
rect 1103 27346 1169 27358
rect 1103 27338 1120 27346
rect 1154 27338 1169 27346
rect 1103 21370 1120 21378
rect 1154 21370 1169 21378
rect 1103 21358 1169 21370
rect 1261 27346 1327 27358
rect 1261 27338 1278 27346
rect 1312 27338 1327 27346
rect 1261 21370 1278 21378
rect 1312 21370 1327 21378
rect 1261 21358 1327 21370
rect 1419 27346 1485 27358
rect 1419 27338 1436 27346
rect 1470 27338 1485 27346
rect 1419 21370 1436 21378
rect 1470 21370 1485 21378
rect 1419 21358 1485 21370
rect 1577 27346 1643 27358
rect 1577 27338 1594 27346
rect 1628 27338 1643 27346
rect 1577 21370 1594 21378
rect 1628 21370 1643 21378
rect 1577 21358 1643 21370
rect 1735 27346 1801 27358
rect 1735 27338 1752 27346
rect 1786 27338 1801 27346
rect 1735 21370 1752 21378
rect 1786 21370 1801 21378
rect 1735 21358 1801 21370
rect 1893 27346 1959 27358
rect 1893 27338 1910 27346
rect 1944 27338 1959 27346
rect 1893 21370 1910 21378
rect 1944 21370 1959 21378
rect 1893 21358 1959 21370
rect 2051 27346 2117 27358
rect 2051 27338 2068 27346
rect 2102 27338 2117 27346
rect 2051 21370 2068 21378
rect 2102 21370 2117 21378
rect 2051 21358 2117 21370
rect 2209 27346 2275 27358
rect 2209 27338 2226 27346
rect 2260 27338 2275 27346
rect 2209 21370 2226 21378
rect 2260 21370 2275 21378
rect 2209 21358 2275 21370
rect 2367 27346 2433 27358
rect 2367 27338 2384 27346
rect 2418 27338 2433 27346
rect 2367 21370 2384 21378
rect 2418 21370 2433 21378
rect 2367 21358 2433 21370
rect 2525 27346 2591 27358
rect 2525 27338 2542 27346
rect 2576 27338 2591 27346
rect 2525 21370 2542 21378
rect 2576 21370 2591 21378
rect 2525 21358 2591 21370
rect 2683 27346 2749 27358
rect 2683 27338 2700 27346
rect 2734 27338 2749 27346
rect 2683 21370 2700 21378
rect 2734 21370 2749 21378
rect 2683 21358 2749 21370
rect 2841 27346 2907 27358
rect 2841 27338 2858 27346
rect 2892 27338 2907 27346
rect 2841 21370 2858 21378
rect 2892 21370 2907 21378
rect 2841 21358 2907 21370
rect 2999 27346 3065 27358
rect 2999 27338 3016 27346
rect 3050 27338 3065 27346
rect 2999 21370 3016 21378
rect 3050 21370 3065 21378
rect 2999 21358 3065 21370
rect 3157 27346 3223 27358
rect 3157 27338 3174 27346
rect 3208 27338 3223 27346
rect 3157 21370 3174 21378
rect 3208 21370 3223 21378
rect 3157 21358 3223 21370
rect 3315 27346 3381 27358
rect 3315 27338 3332 27346
rect 3366 27338 3381 27346
rect 3315 21370 3332 21378
rect 3366 21370 3381 21378
rect 3315 21358 3381 21370
rect 3473 27346 3539 27358
rect 3473 27338 3490 27346
rect 3524 27338 3539 27346
rect 3473 21370 3490 21378
rect 3524 21370 3539 21378
rect 3473 21358 3539 21370
rect 3631 27346 3697 27358
rect 3631 27338 3648 27346
rect 3682 27338 3697 27346
rect 3631 21370 3648 21378
rect 3682 21370 3697 21378
rect 3631 21358 3697 21370
rect 3789 27346 3855 27358
rect 3789 27338 3806 27346
rect 3840 27338 3855 27346
rect 3789 21370 3806 21378
rect 3840 21370 3855 21378
rect 3789 21358 3855 21370
rect 3947 27346 4013 27358
rect 3947 27338 3964 27346
rect 3998 27338 4013 27346
rect 3947 21370 3964 21378
rect 3998 21370 4013 21378
rect 3947 21358 4013 21370
rect 4105 27346 4171 27358
rect 4105 27338 4122 27346
rect 4156 27338 4171 27346
rect 4105 21370 4122 21378
rect 4156 21370 4171 21378
rect 4105 21358 4171 21370
rect -568 21320 -548 21326
rect 4086 21320 4106 21326
rect -568 21286 -556 21320
rect 4094 21286 4106 21320
rect -568 21226 -548 21286
rect 4086 21226 4106 21286
rect -770 21194 -700 21200
rect 4240 21194 4310 21200
rect -770 21184 4310 21194
rect -770 21146 -564 21184
rect 4102 21146 4310 21184
rect -770 21130 4310 21146
rect 5530 27570 10610 27580
rect 5530 27532 5736 27570
rect 10459 27532 10610 27570
rect 5530 27522 10610 27532
rect 5530 27520 5600 27522
rect 10540 27520 10610 27522
rect 5732 27430 5752 27490
rect 10386 27430 10406 27490
rect 5732 27396 5744 27430
rect 10394 27396 10406 27430
rect 5732 27390 5752 27396
rect 10386 27390 10406 27396
rect 5665 27346 5731 27358
rect 5665 27338 5682 27346
rect 5716 27338 5731 27346
rect 5665 21370 5682 21378
rect 5716 21370 5731 21378
rect 5665 21358 5731 21370
rect 5823 27346 5889 27358
rect 5823 27338 5840 27346
rect 5874 27338 5889 27346
rect 5823 21370 5840 21378
rect 5874 21370 5889 21378
rect 5823 21358 5889 21370
rect 5981 27346 6047 27358
rect 5981 27338 5998 27346
rect 6032 27338 6047 27346
rect 5981 21370 5998 21378
rect 6032 21370 6047 21378
rect 5981 21358 6047 21370
rect 6139 27346 6205 27358
rect 6139 27338 6156 27346
rect 6190 27338 6205 27346
rect 6139 21370 6156 21378
rect 6190 21370 6205 21378
rect 6139 21358 6205 21370
rect 6297 27346 6363 27358
rect 6297 27338 6314 27346
rect 6348 27338 6363 27346
rect 6297 21370 6314 21378
rect 6348 21370 6363 21378
rect 6297 21358 6363 21370
rect 6455 27346 6521 27358
rect 6455 27338 6472 27346
rect 6506 27338 6521 27346
rect 6455 21370 6472 21378
rect 6506 21370 6521 21378
rect 6455 21358 6521 21370
rect 6613 27346 6679 27358
rect 6613 27338 6630 27346
rect 6664 27338 6679 27346
rect 6613 21370 6630 21378
rect 6664 21370 6679 21378
rect 6613 21358 6679 21370
rect 6771 27346 6837 27358
rect 6771 27338 6788 27346
rect 6822 27338 6837 27346
rect 6771 21370 6788 21378
rect 6822 21370 6837 21378
rect 6771 21358 6837 21370
rect 6929 27346 6995 27358
rect 6929 27338 6946 27346
rect 6980 27338 6995 27346
rect 6929 21370 6946 21378
rect 6980 21370 6995 21378
rect 6929 21358 6995 21370
rect 7087 27346 7153 27358
rect 7087 27338 7104 27346
rect 7138 27338 7153 27346
rect 7087 21370 7104 21378
rect 7138 21370 7153 21378
rect 7087 21358 7153 21370
rect 7245 27346 7311 27358
rect 7245 27338 7262 27346
rect 7296 27338 7311 27346
rect 7245 21370 7262 21378
rect 7296 21370 7311 21378
rect 7245 21358 7311 21370
rect 7403 27346 7469 27358
rect 7403 27338 7420 27346
rect 7454 27338 7469 27346
rect 7403 21370 7420 21378
rect 7454 21370 7469 21378
rect 7403 21358 7469 21370
rect 7561 27346 7627 27358
rect 7561 27338 7578 27346
rect 7612 27338 7627 27346
rect 7561 21370 7578 21378
rect 7612 21370 7627 21378
rect 7561 21358 7627 21370
rect 7719 27346 7785 27358
rect 7719 27338 7736 27346
rect 7770 27338 7785 27346
rect 7719 21370 7736 21378
rect 7770 21370 7785 21378
rect 7719 21358 7785 21370
rect 7877 27346 7943 27358
rect 7877 27338 7894 27346
rect 7928 27338 7943 27346
rect 7877 21370 7894 21378
rect 7928 21370 7943 21378
rect 7877 21358 7943 21370
rect 8035 27346 8101 27358
rect 8035 27338 8052 27346
rect 8086 27338 8101 27346
rect 8035 21370 8052 21378
rect 8086 21370 8101 21378
rect 8035 21358 8101 21370
rect 8193 27346 8259 27358
rect 8193 27338 8210 27346
rect 8244 27338 8259 27346
rect 8193 21370 8210 21378
rect 8244 21370 8259 21378
rect 8193 21358 8259 21370
rect 8351 27346 8417 27358
rect 8351 27338 8368 27346
rect 8402 27338 8417 27346
rect 8351 21370 8368 21378
rect 8402 21370 8417 21378
rect 8351 21358 8417 21370
rect 8509 27346 8575 27358
rect 8509 27338 8526 27346
rect 8560 27338 8575 27346
rect 8509 21370 8526 21378
rect 8560 21370 8575 21378
rect 8509 21358 8575 21370
rect 8667 27346 8733 27358
rect 8667 27338 8684 27346
rect 8718 27338 8733 27346
rect 8667 21370 8684 21378
rect 8718 21370 8733 21378
rect 8667 21358 8733 21370
rect 8825 27346 8891 27358
rect 8825 27338 8842 27346
rect 8876 27338 8891 27346
rect 8825 21370 8842 21378
rect 8876 21370 8891 21378
rect 8825 21358 8891 21370
rect 8983 27346 9049 27358
rect 8983 27338 9000 27346
rect 9034 27338 9049 27346
rect 8983 21370 9000 21378
rect 9034 21370 9049 21378
rect 8983 21358 9049 21370
rect 9141 27346 9207 27358
rect 9141 27338 9158 27346
rect 9192 27338 9207 27346
rect 9141 21370 9158 21378
rect 9192 21370 9207 21378
rect 9141 21358 9207 21370
rect 9299 27346 9365 27358
rect 9299 27338 9316 27346
rect 9350 27338 9365 27346
rect 9299 21370 9316 21378
rect 9350 21370 9365 21378
rect 9299 21358 9365 21370
rect 9457 27346 9523 27358
rect 9457 27338 9474 27346
rect 9508 27338 9523 27346
rect 9457 21370 9474 21378
rect 9508 21370 9523 21378
rect 9457 21358 9523 21370
rect 9615 27346 9681 27358
rect 9615 27338 9632 27346
rect 9666 27338 9681 27346
rect 9615 21370 9632 21378
rect 9666 21370 9681 21378
rect 9615 21358 9681 21370
rect 9773 27346 9839 27358
rect 9773 27338 9790 27346
rect 9824 27338 9839 27346
rect 9773 21370 9790 21378
rect 9824 21370 9839 21378
rect 9773 21358 9839 21370
rect 9931 27346 9997 27358
rect 9931 27338 9948 27346
rect 9982 27338 9997 27346
rect 9931 21370 9948 21378
rect 9982 21370 9997 21378
rect 9931 21358 9997 21370
rect 10089 27346 10155 27358
rect 10089 27338 10106 27346
rect 10140 27338 10155 27346
rect 10089 21370 10106 21378
rect 10140 21370 10155 21378
rect 10089 21358 10155 21370
rect 10247 27346 10313 27358
rect 10247 27338 10264 27346
rect 10298 27338 10313 27346
rect 10247 21370 10264 21378
rect 10298 21370 10313 21378
rect 10247 21358 10313 21370
rect 10405 27346 10471 27358
rect 10405 27338 10422 27346
rect 10456 27338 10471 27346
rect 10405 21370 10422 21378
rect 10456 21370 10471 21378
rect 10405 21358 10471 21370
rect 5732 21320 5752 21326
rect 10386 21320 10406 21326
rect 5732 21286 5744 21320
rect 10394 21286 10406 21320
rect 5732 21226 5752 21286
rect 10386 21226 10406 21286
rect 5530 21194 5600 21200
rect 10540 21194 10610 21200
rect 5530 21184 10610 21194
rect 5530 21146 5736 21184
rect 10402 21146 10610 21184
rect 5530 21130 10610 21146
rect -13370 19270 -8290 19280
rect -13370 19232 -13164 19270
rect -8441 19232 -8290 19270
rect -13370 19222 -8290 19232
rect -13370 19220 -13300 19222
rect -8360 19220 -8290 19222
rect -13168 19130 -13148 19190
rect -8514 19130 -8494 19190
rect -13168 19096 -13156 19130
rect -8506 19096 -8494 19130
rect -13168 19090 -13148 19096
rect -8514 19090 -8494 19096
rect -13235 19046 -13169 19058
rect -13235 19038 -13218 19046
rect -13184 19038 -13169 19046
rect -13235 13070 -13218 13078
rect -13184 13070 -13169 13078
rect -13235 13058 -13169 13070
rect -13077 19046 -13011 19058
rect -13077 19038 -13060 19046
rect -13026 19038 -13011 19046
rect -13077 13070 -13060 13078
rect -13026 13070 -13011 13078
rect -13077 13058 -13011 13070
rect -12919 19046 -12853 19058
rect -12919 19038 -12902 19046
rect -12868 19038 -12853 19046
rect -12919 13070 -12902 13078
rect -12868 13070 -12853 13078
rect -12919 13058 -12853 13070
rect -12761 19046 -12695 19058
rect -12761 19038 -12744 19046
rect -12710 19038 -12695 19046
rect -12761 13070 -12744 13078
rect -12710 13070 -12695 13078
rect -12761 13058 -12695 13070
rect -12603 19046 -12537 19058
rect -12603 19038 -12586 19046
rect -12552 19038 -12537 19046
rect -12603 13070 -12586 13078
rect -12552 13070 -12537 13078
rect -12603 13058 -12537 13070
rect -12445 19046 -12379 19058
rect -12445 19038 -12428 19046
rect -12394 19038 -12379 19046
rect -12445 13070 -12428 13078
rect -12394 13070 -12379 13078
rect -12445 13058 -12379 13070
rect -12287 19046 -12221 19058
rect -12287 19038 -12270 19046
rect -12236 19038 -12221 19046
rect -12287 13070 -12270 13078
rect -12236 13070 -12221 13078
rect -12287 13058 -12221 13070
rect -12129 19046 -12063 19058
rect -12129 19038 -12112 19046
rect -12078 19038 -12063 19046
rect -12129 13070 -12112 13078
rect -12078 13070 -12063 13078
rect -12129 13058 -12063 13070
rect -11971 19046 -11905 19058
rect -11971 19038 -11954 19046
rect -11920 19038 -11905 19046
rect -11971 13070 -11954 13078
rect -11920 13070 -11905 13078
rect -11971 13058 -11905 13070
rect -11813 19046 -11747 19058
rect -11813 19038 -11796 19046
rect -11762 19038 -11747 19046
rect -11813 13070 -11796 13078
rect -11762 13070 -11747 13078
rect -11813 13058 -11747 13070
rect -11655 19046 -11589 19058
rect -11655 19038 -11638 19046
rect -11604 19038 -11589 19046
rect -11655 13070 -11638 13078
rect -11604 13070 -11589 13078
rect -11655 13058 -11589 13070
rect -11497 19046 -11431 19058
rect -11497 19038 -11480 19046
rect -11446 19038 -11431 19046
rect -11497 13070 -11480 13078
rect -11446 13070 -11431 13078
rect -11497 13058 -11431 13070
rect -11339 19046 -11273 19058
rect -11339 19038 -11322 19046
rect -11288 19038 -11273 19046
rect -11339 13070 -11322 13078
rect -11288 13070 -11273 13078
rect -11339 13058 -11273 13070
rect -11181 19046 -11115 19058
rect -11181 19038 -11164 19046
rect -11130 19038 -11115 19046
rect -11181 13070 -11164 13078
rect -11130 13070 -11115 13078
rect -11181 13058 -11115 13070
rect -11023 19046 -10957 19058
rect -11023 19038 -11006 19046
rect -10972 19038 -10957 19046
rect -11023 13070 -11006 13078
rect -10972 13070 -10957 13078
rect -11023 13058 -10957 13070
rect -10865 19046 -10799 19058
rect -10865 19038 -10848 19046
rect -10814 19038 -10799 19046
rect -10865 13070 -10848 13078
rect -10814 13070 -10799 13078
rect -10865 13058 -10799 13070
rect -10707 19046 -10641 19058
rect -10707 19038 -10690 19046
rect -10656 19038 -10641 19046
rect -10707 13070 -10690 13078
rect -10656 13070 -10641 13078
rect -10707 13058 -10641 13070
rect -10549 19046 -10483 19058
rect -10549 19038 -10532 19046
rect -10498 19038 -10483 19046
rect -10549 13070 -10532 13078
rect -10498 13070 -10483 13078
rect -10549 13058 -10483 13070
rect -10391 19046 -10325 19058
rect -10391 19038 -10374 19046
rect -10340 19038 -10325 19046
rect -10391 13070 -10374 13078
rect -10340 13070 -10325 13078
rect -10391 13058 -10325 13070
rect -10233 19046 -10167 19058
rect -10233 19038 -10216 19046
rect -10182 19038 -10167 19046
rect -10233 13070 -10216 13078
rect -10182 13070 -10167 13078
rect -10233 13058 -10167 13070
rect -10075 19046 -10009 19058
rect -10075 19038 -10058 19046
rect -10024 19038 -10009 19046
rect -10075 13070 -10058 13078
rect -10024 13070 -10009 13078
rect -10075 13058 -10009 13070
rect -9917 19046 -9851 19058
rect -9917 19038 -9900 19046
rect -9866 19038 -9851 19046
rect -9917 13070 -9900 13078
rect -9866 13070 -9851 13078
rect -9917 13058 -9851 13070
rect -9759 19046 -9693 19058
rect -9759 19038 -9742 19046
rect -9708 19038 -9693 19046
rect -9759 13070 -9742 13078
rect -9708 13070 -9693 13078
rect -9759 13058 -9693 13070
rect -9601 19046 -9535 19058
rect -9601 19038 -9584 19046
rect -9550 19038 -9535 19046
rect -9601 13070 -9584 13078
rect -9550 13070 -9535 13078
rect -9601 13058 -9535 13070
rect -9443 19046 -9377 19058
rect -9443 19038 -9426 19046
rect -9392 19038 -9377 19046
rect -9443 13070 -9426 13078
rect -9392 13070 -9377 13078
rect -9443 13058 -9377 13070
rect -9285 19046 -9219 19058
rect -9285 19038 -9268 19046
rect -9234 19038 -9219 19046
rect -9285 13070 -9268 13078
rect -9234 13070 -9219 13078
rect -9285 13058 -9219 13070
rect -9127 19046 -9061 19058
rect -9127 19038 -9110 19046
rect -9076 19038 -9061 19046
rect -9127 13070 -9110 13078
rect -9076 13070 -9061 13078
rect -9127 13058 -9061 13070
rect -8969 19046 -8903 19058
rect -8969 19038 -8952 19046
rect -8918 19038 -8903 19046
rect -8969 13070 -8952 13078
rect -8918 13070 -8903 13078
rect -8969 13058 -8903 13070
rect -8811 19046 -8745 19058
rect -8811 19038 -8794 19046
rect -8760 19038 -8745 19046
rect -8811 13070 -8794 13078
rect -8760 13070 -8745 13078
rect -8811 13058 -8745 13070
rect -8653 19046 -8587 19058
rect -8653 19038 -8636 19046
rect -8602 19038 -8587 19046
rect -8653 13070 -8636 13078
rect -8602 13070 -8587 13078
rect -8653 13058 -8587 13070
rect -8495 19046 -8429 19058
rect -8495 19038 -8478 19046
rect -8444 19038 -8429 19046
rect -8495 13070 -8478 13078
rect -8444 13070 -8429 13078
rect -8495 13058 -8429 13070
rect -13168 13020 -13148 13026
rect -8514 13020 -8494 13026
rect -13168 12986 -13156 13020
rect -8506 12986 -8494 13020
rect -13168 12926 -13148 12986
rect -8514 12926 -8494 12986
rect -13370 12894 -13300 12900
rect -8360 12894 -8290 12900
rect -13370 12884 -8290 12894
rect -13370 12846 -13164 12884
rect -8498 12846 -8290 12884
rect -13370 12830 -8290 12846
rect -7070 19270 -1990 19280
rect -7070 19232 -6864 19270
rect -2141 19232 -1990 19270
rect -7070 19222 -1990 19232
rect -7070 19220 -7000 19222
rect -2060 19220 -1990 19222
rect -6868 19130 -6848 19190
rect -2214 19130 -2194 19190
rect -6868 19096 -6856 19130
rect -2206 19096 -2194 19130
rect -6868 19090 -6848 19096
rect -2214 19090 -2194 19096
rect -6935 19046 -6869 19058
rect -6935 19038 -6918 19046
rect -6884 19038 -6869 19046
rect -6935 13070 -6918 13078
rect -6884 13070 -6869 13078
rect -6935 13058 -6869 13070
rect -6777 19046 -6711 19058
rect -6777 19038 -6760 19046
rect -6726 19038 -6711 19046
rect -6777 13070 -6760 13078
rect -6726 13070 -6711 13078
rect -6777 13058 -6711 13070
rect -6619 19046 -6553 19058
rect -6619 19038 -6602 19046
rect -6568 19038 -6553 19046
rect -6619 13070 -6602 13078
rect -6568 13070 -6553 13078
rect -6619 13058 -6553 13070
rect -6461 19046 -6395 19058
rect -6461 19038 -6444 19046
rect -6410 19038 -6395 19046
rect -6461 13070 -6444 13078
rect -6410 13070 -6395 13078
rect -6461 13058 -6395 13070
rect -6303 19046 -6237 19058
rect -6303 19038 -6286 19046
rect -6252 19038 -6237 19046
rect -6303 13070 -6286 13078
rect -6252 13070 -6237 13078
rect -6303 13058 -6237 13070
rect -6145 19046 -6079 19058
rect -6145 19038 -6128 19046
rect -6094 19038 -6079 19046
rect -6145 13070 -6128 13078
rect -6094 13070 -6079 13078
rect -6145 13058 -6079 13070
rect -5987 19046 -5921 19058
rect -5987 19038 -5970 19046
rect -5936 19038 -5921 19046
rect -5987 13070 -5970 13078
rect -5936 13070 -5921 13078
rect -5987 13058 -5921 13070
rect -5829 19046 -5763 19058
rect -5829 19038 -5812 19046
rect -5778 19038 -5763 19046
rect -5829 13070 -5812 13078
rect -5778 13070 -5763 13078
rect -5829 13058 -5763 13070
rect -5671 19046 -5605 19058
rect -5671 19038 -5654 19046
rect -5620 19038 -5605 19046
rect -5671 13070 -5654 13078
rect -5620 13070 -5605 13078
rect -5671 13058 -5605 13070
rect -5513 19046 -5447 19058
rect -5513 19038 -5496 19046
rect -5462 19038 -5447 19046
rect -5513 13070 -5496 13078
rect -5462 13070 -5447 13078
rect -5513 13058 -5447 13070
rect -5355 19046 -5289 19058
rect -5355 19038 -5338 19046
rect -5304 19038 -5289 19046
rect -5355 13070 -5338 13078
rect -5304 13070 -5289 13078
rect -5355 13058 -5289 13070
rect -5197 19046 -5131 19058
rect -5197 19038 -5180 19046
rect -5146 19038 -5131 19046
rect -5197 13070 -5180 13078
rect -5146 13070 -5131 13078
rect -5197 13058 -5131 13070
rect -5039 19046 -4973 19058
rect -5039 19038 -5022 19046
rect -4988 19038 -4973 19046
rect -5039 13070 -5022 13078
rect -4988 13070 -4973 13078
rect -5039 13058 -4973 13070
rect -4881 19046 -4815 19058
rect -4881 19038 -4864 19046
rect -4830 19038 -4815 19046
rect -4881 13070 -4864 13078
rect -4830 13070 -4815 13078
rect -4881 13058 -4815 13070
rect -4723 19046 -4657 19058
rect -4723 19038 -4706 19046
rect -4672 19038 -4657 19046
rect -4723 13070 -4706 13078
rect -4672 13070 -4657 13078
rect -4723 13058 -4657 13070
rect -4565 19046 -4499 19058
rect -4565 19038 -4548 19046
rect -4514 19038 -4499 19046
rect -4565 13070 -4548 13078
rect -4514 13070 -4499 13078
rect -4565 13058 -4499 13070
rect -4407 19046 -4341 19058
rect -4407 19038 -4390 19046
rect -4356 19038 -4341 19046
rect -4407 13070 -4390 13078
rect -4356 13070 -4341 13078
rect -4407 13058 -4341 13070
rect -4249 19046 -4183 19058
rect -4249 19038 -4232 19046
rect -4198 19038 -4183 19046
rect -4249 13070 -4232 13078
rect -4198 13070 -4183 13078
rect -4249 13058 -4183 13070
rect -4091 19046 -4025 19058
rect -4091 19038 -4074 19046
rect -4040 19038 -4025 19046
rect -4091 13070 -4074 13078
rect -4040 13070 -4025 13078
rect -4091 13058 -4025 13070
rect -3933 19046 -3867 19058
rect -3933 19038 -3916 19046
rect -3882 19038 -3867 19046
rect -3933 13070 -3916 13078
rect -3882 13070 -3867 13078
rect -3933 13058 -3867 13070
rect -3775 19046 -3709 19058
rect -3775 19038 -3758 19046
rect -3724 19038 -3709 19046
rect -3775 13070 -3758 13078
rect -3724 13070 -3709 13078
rect -3775 13058 -3709 13070
rect -3617 19046 -3551 19058
rect -3617 19038 -3600 19046
rect -3566 19038 -3551 19046
rect -3617 13070 -3600 13078
rect -3566 13070 -3551 13078
rect -3617 13058 -3551 13070
rect -3459 19046 -3393 19058
rect -3459 19038 -3442 19046
rect -3408 19038 -3393 19046
rect -3459 13070 -3442 13078
rect -3408 13070 -3393 13078
rect -3459 13058 -3393 13070
rect -3301 19046 -3235 19058
rect -3301 19038 -3284 19046
rect -3250 19038 -3235 19046
rect -3301 13070 -3284 13078
rect -3250 13070 -3235 13078
rect -3301 13058 -3235 13070
rect -3143 19046 -3077 19058
rect -3143 19038 -3126 19046
rect -3092 19038 -3077 19046
rect -3143 13070 -3126 13078
rect -3092 13070 -3077 13078
rect -3143 13058 -3077 13070
rect -2985 19046 -2919 19058
rect -2985 19038 -2968 19046
rect -2934 19038 -2919 19046
rect -2985 13070 -2968 13078
rect -2934 13070 -2919 13078
rect -2985 13058 -2919 13070
rect -2827 19046 -2761 19058
rect -2827 19038 -2810 19046
rect -2776 19038 -2761 19046
rect -2827 13070 -2810 13078
rect -2776 13070 -2761 13078
rect -2827 13058 -2761 13070
rect -2669 19046 -2603 19058
rect -2669 19038 -2652 19046
rect -2618 19038 -2603 19046
rect -2669 13070 -2652 13078
rect -2618 13070 -2603 13078
rect -2669 13058 -2603 13070
rect -2511 19046 -2445 19058
rect -2511 19038 -2494 19046
rect -2460 19038 -2445 19046
rect -2511 13070 -2494 13078
rect -2460 13070 -2445 13078
rect -2511 13058 -2445 13070
rect -2353 19046 -2287 19058
rect -2353 19038 -2336 19046
rect -2302 19038 -2287 19046
rect -2353 13070 -2336 13078
rect -2302 13070 -2287 13078
rect -2353 13058 -2287 13070
rect -2195 19046 -2129 19058
rect -2195 19038 -2178 19046
rect -2144 19038 -2129 19046
rect -2195 13070 -2178 13078
rect -2144 13070 -2129 13078
rect -2195 13058 -2129 13070
rect -6868 13020 -6848 13026
rect -2214 13020 -2194 13026
rect -6868 12986 -6856 13020
rect -2206 12986 -2194 13020
rect -6868 12926 -6848 12986
rect -2214 12926 -2194 12986
rect -7070 12894 -7000 12900
rect -2060 12894 -1990 12900
rect -7070 12884 -1990 12894
rect -7070 12846 -6864 12884
rect -2198 12846 -1990 12884
rect -7070 12830 -1990 12846
rect -770 19270 4310 19280
rect -770 19232 -564 19270
rect 4159 19232 4310 19270
rect -770 19222 4310 19232
rect -770 19220 -700 19222
rect 4240 19220 4310 19222
rect -568 19130 -548 19190
rect 4086 19130 4106 19190
rect -568 19096 -556 19130
rect 4094 19096 4106 19130
rect -568 19090 -548 19096
rect 4086 19090 4106 19096
rect -635 19046 -569 19058
rect -635 19038 -618 19046
rect -584 19038 -569 19046
rect -635 13070 -618 13078
rect -584 13070 -569 13078
rect -635 13058 -569 13070
rect -477 19046 -411 19058
rect -477 19038 -460 19046
rect -426 19038 -411 19046
rect -477 13070 -460 13078
rect -426 13070 -411 13078
rect -477 13058 -411 13070
rect -319 19046 -253 19058
rect -319 19038 -302 19046
rect -268 19038 -253 19046
rect -319 13070 -302 13078
rect -268 13070 -253 13078
rect -319 13058 -253 13070
rect -161 19046 -95 19058
rect -161 19038 -144 19046
rect -110 19038 -95 19046
rect -161 13070 -144 13078
rect -110 13070 -95 13078
rect -161 13058 -95 13070
rect -3 19046 63 19058
rect -3 19038 14 19046
rect 48 19038 63 19046
rect -3 13070 14 13078
rect 48 13070 63 13078
rect -3 13058 63 13070
rect 155 19046 221 19058
rect 155 19038 172 19046
rect 206 19038 221 19046
rect 155 13070 172 13078
rect 206 13070 221 13078
rect 155 13058 221 13070
rect 313 19046 379 19058
rect 313 19038 330 19046
rect 364 19038 379 19046
rect 313 13070 330 13078
rect 364 13070 379 13078
rect 313 13058 379 13070
rect 471 19046 537 19058
rect 471 19038 488 19046
rect 522 19038 537 19046
rect 471 13070 488 13078
rect 522 13070 537 13078
rect 471 13058 537 13070
rect 629 19046 695 19058
rect 629 19038 646 19046
rect 680 19038 695 19046
rect 629 13070 646 13078
rect 680 13070 695 13078
rect 629 13058 695 13070
rect 787 19046 853 19058
rect 787 19038 804 19046
rect 838 19038 853 19046
rect 787 13070 804 13078
rect 838 13070 853 13078
rect 787 13058 853 13070
rect 945 19046 1011 19058
rect 945 19038 962 19046
rect 996 19038 1011 19046
rect 945 13070 962 13078
rect 996 13070 1011 13078
rect 945 13058 1011 13070
rect 1103 19046 1169 19058
rect 1103 19038 1120 19046
rect 1154 19038 1169 19046
rect 1103 13070 1120 13078
rect 1154 13070 1169 13078
rect 1103 13058 1169 13070
rect 1261 19046 1327 19058
rect 1261 19038 1278 19046
rect 1312 19038 1327 19046
rect 1261 13070 1278 13078
rect 1312 13070 1327 13078
rect 1261 13058 1327 13070
rect 1419 19046 1485 19058
rect 1419 19038 1436 19046
rect 1470 19038 1485 19046
rect 1419 13070 1436 13078
rect 1470 13070 1485 13078
rect 1419 13058 1485 13070
rect 1577 19046 1643 19058
rect 1577 19038 1594 19046
rect 1628 19038 1643 19046
rect 1577 13070 1594 13078
rect 1628 13070 1643 13078
rect 1577 13058 1643 13070
rect 1735 19046 1801 19058
rect 1735 19038 1752 19046
rect 1786 19038 1801 19046
rect 1735 13070 1752 13078
rect 1786 13070 1801 13078
rect 1735 13058 1801 13070
rect 1893 19046 1959 19058
rect 1893 19038 1910 19046
rect 1944 19038 1959 19046
rect 1893 13070 1910 13078
rect 1944 13070 1959 13078
rect 1893 13058 1959 13070
rect 2051 19046 2117 19058
rect 2051 19038 2068 19046
rect 2102 19038 2117 19046
rect 2051 13070 2068 13078
rect 2102 13070 2117 13078
rect 2051 13058 2117 13070
rect 2209 19046 2275 19058
rect 2209 19038 2226 19046
rect 2260 19038 2275 19046
rect 2209 13070 2226 13078
rect 2260 13070 2275 13078
rect 2209 13058 2275 13070
rect 2367 19046 2433 19058
rect 2367 19038 2384 19046
rect 2418 19038 2433 19046
rect 2367 13070 2384 13078
rect 2418 13070 2433 13078
rect 2367 13058 2433 13070
rect 2525 19046 2591 19058
rect 2525 19038 2542 19046
rect 2576 19038 2591 19046
rect 2525 13070 2542 13078
rect 2576 13070 2591 13078
rect 2525 13058 2591 13070
rect 2683 19046 2749 19058
rect 2683 19038 2700 19046
rect 2734 19038 2749 19046
rect 2683 13070 2700 13078
rect 2734 13070 2749 13078
rect 2683 13058 2749 13070
rect 2841 19046 2907 19058
rect 2841 19038 2858 19046
rect 2892 19038 2907 19046
rect 2841 13070 2858 13078
rect 2892 13070 2907 13078
rect 2841 13058 2907 13070
rect 2999 19046 3065 19058
rect 2999 19038 3016 19046
rect 3050 19038 3065 19046
rect 2999 13070 3016 13078
rect 3050 13070 3065 13078
rect 2999 13058 3065 13070
rect 3157 19046 3223 19058
rect 3157 19038 3174 19046
rect 3208 19038 3223 19046
rect 3157 13070 3174 13078
rect 3208 13070 3223 13078
rect 3157 13058 3223 13070
rect 3315 19046 3381 19058
rect 3315 19038 3332 19046
rect 3366 19038 3381 19046
rect 3315 13070 3332 13078
rect 3366 13070 3381 13078
rect 3315 13058 3381 13070
rect 3473 19046 3539 19058
rect 3473 19038 3490 19046
rect 3524 19038 3539 19046
rect 3473 13070 3490 13078
rect 3524 13070 3539 13078
rect 3473 13058 3539 13070
rect 3631 19046 3697 19058
rect 3631 19038 3648 19046
rect 3682 19038 3697 19046
rect 3631 13070 3648 13078
rect 3682 13070 3697 13078
rect 3631 13058 3697 13070
rect 3789 19046 3855 19058
rect 3789 19038 3806 19046
rect 3840 19038 3855 19046
rect 3789 13070 3806 13078
rect 3840 13070 3855 13078
rect 3789 13058 3855 13070
rect 3947 19046 4013 19058
rect 3947 19038 3964 19046
rect 3998 19038 4013 19046
rect 3947 13070 3964 13078
rect 3998 13070 4013 13078
rect 3947 13058 4013 13070
rect 4105 19046 4171 19058
rect 4105 19038 4122 19046
rect 4156 19038 4171 19046
rect 4105 13070 4122 13078
rect 4156 13070 4171 13078
rect 4105 13058 4171 13070
rect -568 13020 -548 13026
rect 4086 13020 4106 13026
rect -568 12986 -556 13020
rect 4094 12986 4106 13020
rect -568 12926 -548 12986
rect 4086 12926 4106 12986
rect -770 12894 -700 12900
rect 4240 12894 4310 12900
rect -770 12884 4310 12894
rect -770 12846 -564 12884
rect 4102 12846 4310 12884
rect -770 12830 4310 12846
rect 5530 19270 10610 19280
rect 5530 19232 5736 19270
rect 10459 19232 10610 19270
rect 5530 19222 10610 19232
rect 5530 19220 5600 19222
rect 10540 19220 10610 19222
rect 5732 19130 5752 19190
rect 10386 19130 10406 19190
rect 5732 19096 5744 19130
rect 10394 19096 10406 19130
rect 5732 19090 5752 19096
rect 10386 19090 10406 19096
rect 5665 19046 5731 19058
rect 5665 19038 5682 19046
rect 5716 19038 5731 19046
rect 5665 13070 5682 13078
rect 5716 13070 5731 13078
rect 5665 13058 5731 13070
rect 5823 19046 5889 19058
rect 5823 19038 5840 19046
rect 5874 19038 5889 19046
rect 5823 13070 5840 13078
rect 5874 13070 5889 13078
rect 5823 13058 5889 13070
rect 5981 19046 6047 19058
rect 5981 19038 5998 19046
rect 6032 19038 6047 19046
rect 5981 13070 5998 13078
rect 6032 13070 6047 13078
rect 5981 13058 6047 13070
rect 6139 19046 6205 19058
rect 6139 19038 6156 19046
rect 6190 19038 6205 19046
rect 6139 13070 6156 13078
rect 6190 13070 6205 13078
rect 6139 13058 6205 13070
rect 6297 19046 6363 19058
rect 6297 19038 6314 19046
rect 6348 19038 6363 19046
rect 6297 13070 6314 13078
rect 6348 13070 6363 13078
rect 6297 13058 6363 13070
rect 6455 19046 6521 19058
rect 6455 19038 6472 19046
rect 6506 19038 6521 19046
rect 6455 13070 6472 13078
rect 6506 13070 6521 13078
rect 6455 13058 6521 13070
rect 6613 19046 6679 19058
rect 6613 19038 6630 19046
rect 6664 19038 6679 19046
rect 6613 13070 6630 13078
rect 6664 13070 6679 13078
rect 6613 13058 6679 13070
rect 6771 19046 6837 19058
rect 6771 19038 6788 19046
rect 6822 19038 6837 19046
rect 6771 13070 6788 13078
rect 6822 13070 6837 13078
rect 6771 13058 6837 13070
rect 6929 19046 6995 19058
rect 6929 19038 6946 19046
rect 6980 19038 6995 19046
rect 6929 13070 6946 13078
rect 6980 13070 6995 13078
rect 6929 13058 6995 13070
rect 7087 19046 7153 19058
rect 7087 19038 7104 19046
rect 7138 19038 7153 19046
rect 7087 13070 7104 13078
rect 7138 13070 7153 13078
rect 7087 13058 7153 13070
rect 7245 19046 7311 19058
rect 7245 19038 7262 19046
rect 7296 19038 7311 19046
rect 7245 13070 7262 13078
rect 7296 13070 7311 13078
rect 7245 13058 7311 13070
rect 7403 19046 7469 19058
rect 7403 19038 7420 19046
rect 7454 19038 7469 19046
rect 7403 13070 7420 13078
rect 7454 13070 7469 13078
rect 7403 13058 7469 13070
rect 7561 19046 7627 19058
rect 7561 19038 7578 19046
rect 7612 19038 7627 19046
rect 7561 13070 7578 13078
rect 7612 13070 7627 13078
rect 7561 13058 7627 13070
rect 7719 19046 7785 19058
rect 7719 19038 7736 19046
rect 7770 19038 7785 19046
rect 7719 13070 7736 13078
rect 7770 13070 7785 13078
rect 7719 13058 7785 13070
rect 7877 19046 7943 19058
rect 7877 19038 7894 19046
rect 7928 19038 7943 19046
rect 7877 13070 7894 13078
rect 7928 13070 7943 13078
rect 7877 13058 7943 13070
rect 8035 19046 8101 19058
rect 8035 19038 8052 19046
rect 8086 19038 8101 19046
rect 8035 13070 8052 13078
rect 8086 13070 8101 13078
rect 8035 13058 8101 13070
rect 8193 19046 8259 19058
rect 8193 19038 8210 19046
rect 8244 19038 8259 19046
rect 8193 13070 8210 13078
rect 8244 13070 8259 13078
rect 8193 13058 8259 13070
rect 8351 19046 8417 19058
rect 8351 19038 8368 19046
rect 8402 19038 8417 19046
rect 8351 13070 8368 13078
rect 8402 13070 8417 13078
rect 8351 13058 8417 13070
rect 8509 19046 8575 19058
rect 8509 19038 8526 19046
rect 8560 19038 8575 19046
rect 8509 13070 8526 13078
rect 8560 13070 8575 13078
rect 8509 13058 8575 13070
rect 8667 19046 8733 19058
rect 8667 19038 8684 19046
rect 8718 19038 8733 19046
rect 8667 13070 8684 13078
rect 8718 13070 8733 13078
rect 8667 13058 8733 13070
rect 8825 19046 8891 19058
rect 8825 19038 8842 19046
rect 8876 19038 8891 19046
rect 8825 13070 8842 13078
rect 8876 13070 8891 13078
rect 8825 13058 8891 13070
rect 8983 19046 9049 19058
rect 8983 19038 9000 19046
rect 9034 19038 9049 19046
rect 8983 13070 9000 13078
rect 9034 13070 9049 13078
rect 8983 13058 9049 13070
rect 9141 19046 9207 19058
rect 9141 19038 9158 19046
rect 9192 19038 9207 19046
rect 9141 13070 9158 13078
rect 9192 13070 9207 13078
rect 9141 13058 9207 13070
rect 9299 19046 9365 19058
rect 9299 19038 9316 19046
rect 9350 19038 9365 19046
rect 9299 13070 9316 13078
rect 9350 13070 9365 13078
rect 9299 13058 9365 13070
rect 9457 19046 9523 19058
rect 9457 19038 9474 19046
rect 9508 19038 9523 19046
rect 9457 13070 9474 13078
rect 9508 13070 9523 13078
rect 9457 13058 9523 13070
rect 9615 19046 9681 19058
rect 9615 19038 9632 19046
rect 9666 19038 9681 19046
rect 9615 13070 9632 13078
rect 9666 13070 9681 13078
rect 9615 13058 9681 13070
rect 9773 19046 9839 19058
rect 9773 19038 9790 19046
rect 9824 19038 9839 19046
rect 9773 13070 9790 13078
rect 9824 13070 9839 13078
rect 9773 13058 9839 13070
rect 9931 19046 9997 19058
rect 9931 19038 9948 19046
rect 9982 19038 9997 19046
rect 9931 13070 9948 13078
rect 9982 13070 9997 13078
rect 9931 13058 9997 13070
rect 10089 19046 10155 19058
rect 10089 19038 10106 19046
rect 10140 19038 10155 19046
rect 10089 13070 10106 13078
rect 10140 13070 10155 13078
rect 10089 13058 10155 13070
rect 10247 19046 10313 19058
rect 10247 19038 10264 19046
rect 10298 19038 10313 19046
rect 10247 13070 10264 13078
rect 10298 13070 10313 13078
rect 10247 13058 10313 13070
rect 10405 19046 10471 19058
rect 10405 19038 10422 19046
rect 10456 19038 10471 19046
rect 10405 13070 10422 13078
rect 10456 13070 10471 13078
rect 10405 13058 10471 13070
rect 5732 13020 5752 13026
rect 10386 13020 10406 13026
rect 5732 12986 5744 13020
rect 10394 12986 10406 13020
rect 5732 12926 5752 12986
rect 10386 12926 10406 12986
rect 5530 12894 5600 12900
rect 10540 12894 10610 12900
rect 5530 12884 10610 12894
rect 5530 12846 5736 12884
rect 10402 12846 10610 12884
rect 5530 12830 10610 12846
rect -13370 12270 -8290 12280
rect -13370 12232 -13164 12270
rect -8441 12232 -8290 12270
rect -13370 12222 -8290 12232
rect -13370 12220 -13300 12222
rect -8360 12220 -8290 12222
rect -13168 12130 -13148 12190
rect -8514 12130 -8494 12190
rect -13168 12096 -13156 12130
rect -8506 12096 -8494 12130
rect -13168 12090 -13148 12096
rect -8514 12090 -8494 12096
rect -13235 12046 -13169 12058
rect -13235 12038 -13218 12046
rect -13184 12038 -13169 12046
rect -13235 6070 -13218 6078
rect -13184 6070 -13169 6078
rect -13235 6058 -13169 6070
rect -13077 12046 -13011 12058
rect -13077 12038 -13060 12046
rect -13026 12038 -13011 12046
rect -13077 6070 -13060 6078
rect -13026 6070 -13011 6078
rect -13077 6058 -13011 6070
rect -12919 12046 -12853 12058
rect -12919 12038 -12902 12046
rect -12868 12038 -12853 12046
rect -12919 6070 -12902 6078
rect -12868 6070 -12853 6078
rect -12919 6058 -12853 6070
rect -12761 12046 -12695 12058
rect -12761 12038 -12744 12046
rect -12710 12038 -12695 12046
rect -12761 6070 -12744 6078
rect -12710 6070 -12695 6078
rect -12761 6058 -12695 6070
rect -12603 12046 -12537 12058
rect -12603 12038 -12586 12046
rect -12552 12038 -12537 12046
rect -12603 6070 -12586 6078
rect -12552 6070 -12537 6078
rect -12603 6058 -12537 6070
rect -12445 12046 -12379 12058
rect -12445 12038 -12428 12046
rect -12394 12038 -12379 12046
rect -12445 6070 -12428 6078
rect -12394 6070 -12379 6078
rect -12445 6058 -12379 6070
rect -12287 12046 -12221 12058
rect -12287 12038 -12270 12046
rect -12236 12038 -12221 12046
rect -12287 6070 -12270 6078
rect -12236 6070 -12221 6078
rect -12287 6058 -12221 6070
rect -12129 12046 -12063 12058
rect -12129 12038 -12112 12046
rect -12078 12038 -12063 12046
rect -12129 6070 -12112 6078
rect -12078 6070 -12063 6078
rect -12129 6058 -12063 6070
rect -11971 12046 -11905 12058
rect -11971 12038 -11954 12046
rect -11920 12038 -11905 12046
rect -11971 6070 -11954 6078
rect -11920 6070 -11905 6078
rect -11971 6058 -11905 6070
rect -11813 12046 -11747 12058
rect -11813 12038 -11796 12046
rect -11762 12038 -11747 12046
rect -11813 6070 -11796 6078
rect -11762 6070 -11747 6078
rect -11813 6058 -11747 6070
rect -11655 12046 -11589 12058
rect -11655 12038 -11638 12046
rect -11604 12038 -11589 12046
rect -11655 6070 -11638 6078
rect -11604 6070 -11589 6078
rect -11655 6058 -11589 6070
rect -11497 12046 -11431 12058
rect -11497 12038 -11480 12046
rect -11446 12038 -11431 12046
rect -11497 6070 -11480 6078
rect -11446 6070 -11431 6078
rect -11497 6058 -11431 6070
rect -11339 12046 -11273 12058
rect -11339 12038 -11322 12046
rect -11288 12038 -11273 12046
rect -11339 6070 -11322 6078
rect -11288 6070 -11273 6078
rect -11339 6058 -11273 6070
rect -11181 12046 -11115 12058
rect -11181 12038 -11164 12046
rect -11130 12038 -11115 12046
rect -11181 6070 -11164 6078
rect -11130 6070 -11115 6078
rect -11181 6058 -11115 6070
rect -11023 12046 -10957 12058
rect -11023 12038 -11006 12046
rect -10972 12038 -10957 12046
rect -11023 6070 -11006 6078
rect -10972 6070 -10957 6078
rect -11023 6058 -10957 6070
rect -10865 12046 -10799 12058
rect -10865 12038 -10848 12046
rect -10814 12038 -10799 12046
rect -10865 6070 -10848 6078
rect -10814 6070 -10799 6078
rect -10865 6058 -10799 6070
rect -10707 12046 -10641 12058
rect -10707 12038 -10690 12046
rect -10656 12038 -10641 12046
rect -10707 6070 -10690 6078
rect -10656 6070 -10641 6078
rect -10707 6058 -10641 6070
rect -10549 12046 -10483 12058
rect -10549 12038 -10532 12046
rect -10498 12038 -10483 12046
rect -10549 6070 -10532 6078
rect -10498 6070 -10483 6078
rect -10549 6058 -10483 6070
rect -10391 12046 -10325 12058
rect -10391 12038 -10374 12046
rect -10340 12038 -10325 12046
rect -10391 6070 -10374 6078
rect -10340 6070 -10325 6078
rect -10391 6058 -10325 6070
rect -10233 12046 -10167 12058
rect -10233 12038 -10216 12046
rect -10182 12038 -10167 12046
rect -10233 6070 -10216 6078
rect -10182 6070 -10167 6078
rect -10233 6058 -10167 6070
rect -10075 12046 -10009 12058
rect -10075 12038 -10058 12046
rect -10024 12038 -10009 12046
rect -10075 6070 -10058 6078
rect -10024 6070 -10009 6078
rect -10075 6058 -10009 6070
rect -9917 12046 -9851 12058
rect -9917 12038 -9900 12046
rect -9866 12038 -9851 12046
rect -9917 6070 -9900 6078
rect -9866 6070 -9851 6078
rect -9917 6058 -9851 6070
rect -9759 12046 -9693 12058
rect -9759 12038 -9742 12046
rect -9708 12038 -9693 12046
rect -9759 6070 -9742 6078
rect -9708 6070 -9693 6078
rect -9759 6058 -9693 6070
rect -9601 12046 -9535 12058
rect -9601 12038 -9584 12046
rect -9550 12038 -9535 12046
rect -9601 6070 -9584 6078
rect -9550 6070 -9535 6078
rect -9601 6058 -9535 6070
rect -9443 12046 -9377 12058
rect -9443 12038 -9426 12046
rect -9392 12038 -9377 12046
rect -9443 6070 -9426 6078
rect -9392 6070 -9377 6078
rect -9443 6058 -9377 6070
rect -9285 12046 -9219 12058
rect -9285 12038 -9268 12046
rect -9234 12038 -9219 12046
rect -9285 6070 -9268 6078
rect -9234 6070 -9219 6078
rect -9285 6058 -9219 6070
rect -9127 12046 -9061 12058
rect -9127 12038 -9110 12046
rect -9076 12038 -9061 12046
rect -9127 6070 -9110 6078
rect -9076 6070 -9061 6078
rect -9127 6058 -9061 6070
rect -8969 12046 -8903 12058
rect -8969 12038 -8952 12046
rect -8918 12038 -8903 12046
rect -8969 6070 -8952 6078
rect -8918 6070 -8903 6078
rect -8969 6058 -8903 6070
rect -8811 12046 -8745 12058
rect -8811 12038 -8794 12046
rect -8760 12038 -8745 12046
rect -8811 6070 -8794 6078
rect -8760 6070 -8745 6078
rect -8811 6058 -8745 6070
rect -8653 12046 -8587 12058
rect -8653 12038 -8636 12046
rect -8602 12038 -8587 12046
rect -8653 6070 -8636 6078
rect -8602 6070 -8587 6078
rect -8653 6058 -8587 6070
rect -8495 12046 -8429 12058
rect -8495 12038 -8478 12046
rect -8444 12038 -8429 12046
rect -8495 6070 -8478 6078
rect -8444 6070 -8429 6078
rect -8495 6058 -8429 6070
rect -13168 6020 -13148 6026
rect -8514 6020 -8494 6026
rect -13168 5986 -13156 6020
rect -8506 5986 -8494 6020
rect -13168 5926 -13148 5986
rect -8514 5926 -8494 5986
rect -13370 5894 -13300 5900
rect -8360 5894 -8290 5900
rect -13370 5884 -8290 5894
rect -13370 5846 -13164 5884
rect -8498 5846 -8290 5884
rect -13370 5830 -8290 5846
rect -7070 12270 -1990 12280
rect -7070 12232 -6864 12270
rect -2141 12232 -1990 12270
rect -7070 12222 -1990 12232
rect -7070 12220 -7000 12222
rect -2060 12220 -1990 12222
rect -6868 12130 -6848 12190
rect -2214 12130 -2194 12190
rect -6868 12096 -6856 12130
rect -2206 12096 -2194 12130
rect -6868 12090 -6848 12096
rect -2214 12090 -2194 12096
rect -6935 12046 -6869 12058
rect -6935 12038 -6918 12046
rect -6884 12038 -6869 12046
rect -6935 6070 -6918 6078
rect -6884 6070 -6869 6078
rect -6935 6058 -6869 6070
rect -6777 12046 -6711 12058
rect -6777 12038 -6760 12046
rect -6726 12038 -6711 12046
rect -6777 6070 -6760 6078
rect -6726 6070 -6711 6078
rect -6777 6058 -6711 6070
rect -6619 12046 -6553 12058
rect -6619 12038 -6602 12046
rect -6568 12038 -6553 12046
rect -6619 6070 -6602 6078
rect -6568 6070 -6553 6078
rect -6619 6058 -6553 6070
rect -6461 12046 -6395 12058
rect -6461 12038 -6444 12046
rect -6410 12038 -6395 12046
rect -6461 6070 -6444 6078
rect -6410 6070 -6395 6078
rect -6461 6058 -6395 6070
rect -6303 12046 -6237 12058
rect -6303 12038 -6286 12046
rect -6252 12038 -6237 12046
rect -6303 6070 -6286 6078
rect -6252 6070 -6237 6078
rect -6303 6058 -6237 6070
rect -6145 12046 -6079 12058
rect -6145 12038 -6128 12046
rect -6094 12038 -6079 12046
rect -6145 6070 -6128 6078
rect -6094 6070 -6079 6078
rect -6145 6058 -6079 6070
rect -5987 12046 -5921 12058
rect -5987 12038 -5970 12046
rect -5936 12038 -5921 12046
rect -5987 6070 -5970 6078
rect -5936 6070 -5921 6078
rect -5987 6058 -5921 6070
rect -5829 12046 -5763 12058
rect -5829 12038 -5812 12046
rect -5778 12038 -5763 12046
rect -5829 6070 -5812 6078
rect -5778 6070 -5763 6078
rect -5829 6058 -5763 6070
rect -5671 12046 -5605 12058
rect -5671 12038 -5654 12046
rect -5620 12038 -5605 12046
rect -5671 6070 -5654 6078
rect -5620 6070 -5605 6078
rect -5671 6058 -5605 6070
rect -5513 12046 -5447 12058
rect -5513 12038 -5496 12046
rect -5462 12038 -5447 12046
rect -5513 6070 -5496 6078
rect -5462 6070 -5447 6078
rect -5513 6058 -5447 6070
rect -5355 12046 -5289 12058
rect -5355 12038 -5338 12046
rect -5304 12038 -5289 12046
rect -5355 6070 -5338 6078
rect -5304 6070 -5289 6078
rect -5355 6058 -5289 6070
rect -5197 12046 -5131 12058
rect -5197 12038 -5180 12046
rect -5146 12038 -5131 12046
rect -5197 6070 -5180 6078
rect -5146 6070 -5131 6078
rect -5197 6058 -5131 6070
rect -5039 12046 -4973 12058
rect -5039 12038 -5022 12046
rect -4988 12038 -4973 12046
rect -5039 6070 -5022 6078
rect -4988 6070 -4973 6078
rect -5039 6058 -4973 6070
rect -4881 12046 -4815 12058
rect -4881 12038 -4864 12046
rect -4830 12038 -4815 12046
rect -4881 6070 -4864 6078
rect -4830 6070 -4815 6078
rect -4881 6058 -4815 6070
rect -4723 12046 -4657 12058
rect -4723 12038 -4706 12046
rect -4672 12038 -4657 12046
rect -4723 6070 -4706 6078
rect -4672 6070 -4657 6078
rect -4723 6058 -4657 6070
rect -4565 12046 -4499 12058
rect -4565 12038 -4548 12046
rect -4514 12038 -4499 12046
rect -4565 6070 -4548 6078
rect -4514 6070 -4499 6078
rect -4565 6058 -4499 6070
rect -4407 12046 -4341 12058
rect -4407 12038 -4390 12046
rect -4356 12038 -4341 12046
rect -4407 6070 -4390 6078
rect -4356 6070 -4341 6078
rect -4407 6058 -4341 6070
rect -4249 12046 -4183 12058
rect -4249 12038 -4232 12046
rect -4198 12038 -4183 12046
rect -4249 6070 -4232 6078
rect -4198 6070 -4183 6078
rect -4249 6058 -4183 6070
rect -4091 12046 -4025 12058
rect -4091 12038 -4074 12046
rect -4040 12038 -4025 12046
rect -4091 6070 -4074 6078
rect -4040 6070 -4025 6078
rect -4091 6058 -4025 6070
rect -3933 12046 -3867 12058
rect -3933 12038 -3916 12046
rect -3882 12038 -3867 12046
rect -3933 6070 -3916 6078
rect -3882 6070 -3867 6078
rect -3933 6058 -3867 6070
rect -3775 12046 -3709 12058
rect -3775 12038 -3758 12046
rect -3724 12038 -3709 12046
rect -3775 6070 -3758 6078
rect -3724 6070 -3709 6078
rect -3775 6058 -3709 6070
rect -3617 12046 -3551 12058
rect -3617 12038 -3600 12046
rect -3566 12038 -3551 12046
rect -3617 6070 -3600 6078
rect -3566 6070 -3551 6078
rect -3617 6058 -3551 6070
rect -3459 12046 -3393 12058
rect -3459 12038 -3442 12046
rect -3408 12038 -3393 12046
rect -3459 6070 -3442 6078
rect -3408 6070 -3393 6078
rect -3459 6058 -3393 6070
rect -3301 12046 -3235 12058
rect -3301 12038 -3284 12046
rect -3250 12038 -3235 12046
rect -3301 6070 -3284 6078
rect -3250 6070 -3235 6078
rect -3301 6058 -3235 6070
rect -3143 12046 -3077 12058
rect -3143 12038 -3126 12046
rect -3092 12038 -3077 12046
rect -3143 6070 -3126 6078
rect -3092 6070 -3077 6078
rect -3143 6058 -3077 6070
rect -2985 12046 -2919 12058
rect -2985 12038 -2968 12046
rect -2934 12038 -2919 12046
rect -2985 6070 -2968 6078
rect -2934 6070 -2919 6078
rect -2985 6058 -2919 6070
rect -2827 12046 -2761 12058
rect -2827 12038 -2810 12046
rect -2776 12038 -2761 12046
rect -2827 6070 -2810 6078
rect -2776 6070 -2761 6078
rect -2827 6058 -2761 6070
rect -2669 12046 -2603 12058
rect -2669 12038 -2652 12046
rect -2618 12038 -2603 12046
rect -2669 6070 -2652 6078
rect -2618 6070 -2603 6078
rect -2669 6058 -2603 6070
rect -2511 12046 -2445 12058
rect -2511 12038 -2494 12046
rect -2460 12038 -2445 12046
rect -2511 6070 -2494 6078
rect -2460 6070 -2445 6078
rect -2511 6058 -2445 6070
rect -2353 12046 -2287 12058
rect -2353 12038 -2336 12046
rect -2302 12038 -2287 12046
rect -2353 6070 -2336 6078
rect -2302 6070 -2287 6078
rect -2353 6058 -2287 6070
rect -2195 12046 -2129 12058
rect -2195 12038 -2178 12046
rect -2144 12038 -2129 12046
rect -2195 6070 -2178 6078
rect -2144 6070 -2129 6078
rect -2195 6058 -2129 6070
rect -6868 6020 -6848 6026
rect -2214 6020 -2194 6026
rect -6868 5986 -6856 6020
rect -2206 5986 -2194 6020
rect -6868 5926 -6848 5986
rect -2214 5926 -2194 5986
rect -7070 5894 -7000 5900
rect -2060 5894 -1990 5900
rect -7070 5884 -1990 5894
rect -7070 5846 -6864 5884
rect -2198 5846 -1990 5884
rect -7070 5830 -1990 5846
rect -770 12270 4310 12280
rect -770 12232 -564 12270
rect 4159 12232 4310 12270
rect -770 12222 4310 12232
rect -770 12220 -700 12222
rect 4240 12220 4310 12222
rect -568 12130 -548 12190
rect 4086 12130 4106 12190
rect -568 12096 -556 12130
rect 4094 12096 4106 12130
rect -568 12090 -548 12096
rect 4086 12090 4106 12096
rect -635 12046 -569 12058
rect -635 12038 -618 12046
rect -584 12038 -569 12046
rect -635 6070 -618 6078
rect -584 6070 -569 6078
rect -635 6058 -569 6070
rect -477 12046 -411 12058
rect -477 12038 -460 12046
rect -426 12038 -411 12046
rect -477 6070 -460 6078
rect -426 6070 -411 6078
rect -477 6058 -411 6070
rect -319 12046 -253 12058
rect -319 12038 -302 12046
rect -268 12038 -253 12046
rect -319 6070 -302 6078
rect -268 6070 -253 6078
rect -319 6058 -253 6070
rect -161 12046 -95 12058
rect -161 12038 -144 12046
rect -110 12038 -95 12046
rect -161 6070 -144 6078
rect -110 6070 -95 6078
rect -161 6058 -95 6070
rect -3 12046 63 12058
rect -3 12038 14 12046
rect 48 12038 63 12046
rect -3 6070 14 6078
rect 48 6070 63 6078
rect -3 6058 63 6070
rect 155 12046 221 12058
rect 155 12038 172 12046
rect 206 12038 221 12046
rect 155 6070 172 6078
rect 206 6070 221 6078
rect 155 6058 221 6070
rect 313 12046 379 12058
rect 313 12038 330 12046
rect 364 12038 379 12046
rect 313 6070 330 6078
rect 364 6070 379 6078
rect 313 6058 379 6070
rect 471 12046 537 12058
rect 471 12038 488 12046
rect 522 12038 537 12046
rect 471 6070 488 6078
rect 522 6070 537 6078
rect 471 6058 537 6070
rect 629 12046 695 12058
rect 629 12038 646 12046
rect 680 12038 695 12046
rect 629 6070 646 6078
rect 680 6070 695 6078
rect 629 6058 695 6070
rect 787 12046 853 12058
rect 787 12038 804 12046
rect 838 12038 853 12046
rect 787 6070 804 6078
rect 838 6070 853 6078
rect 787 6058 853 6070
rect 945 12046 1011 12058
rect 945 12038 962 12046
rect 996 12038 1011 12046
rect 945 6070 962 6078
rect 996 6070 1011 6078
rect 945 6058 1011 6070
rect 1103 12046 1169 12058
rect 1103 12038 1120 12046
rect 1154 12038 1169 12046
rect 1103 6070 1120 6078
rect 1154 6070 1169 6078
rect 1103 6058 1169 6070
rect 1261 12046 1327 12058
rect 1261 12038 1278 12046
rect 1312 12038 1327 12046
rect 1261 6070 1278 6078
rect 1312 6070 1327 6078
rect 1261 6058 1327 6070
rect 1419 12046 1485 12058
rect 1419 12038 1436 12046
rect 1470 12038 1485 12046
rect 1419 6070 1436 6078
rect 1470 6070 1485 6078
rect 1419 6058 1485 6070
rect 1577 12046 1643 12058
rect 1577 12038 1594 12046
rect 1628 12038 1643 12046
rect 1577 6070 1594 6078
rect 1628 6070 1643 6078
rect 1577 6058 1643 6070
rect 1735 12046 1801 12058
rect 1735 12038 1752 12046
rect 1786 12038 1801 12046
rect 1735 6070 1752 6078
rect 1786 6070 1801 6078
rect 1735 6058 1801 6070
rect 1893 12046 1959 12058
rect 1893 12038 1910 12046
rect 1944 12038 1959 12046
rect 1893 6070 1910 6078
rect 1944 6070 1959 6078
rect 1893 6058 1959 6070
rect 2051 12046 2117 12058
rect 2051 12038 2068 12046
rect 2102 12038 2117 12046
rect 2051 6070 2068 6078
rect 2102 6070 2117 6078
rect 2051 6058 2117 6070
rect 2209 12046 2275 12058
rect 2209 12038 2226 12046
rect 2260 12038 2275 12046
rect 2209 6070 2226 6078
rect 2260 6070 2275 6078
rect 2209 6058 2275 6070
rect 2367 12046 2433 12058
rect 2367 12038 2384 12046
rect 2418 12038 2433 12046
rect 2367 6070 2384 6078
rect 2418 6070 2433 6078
rect 2367 6058 2433 6070
rect 2525 12046 2591 12058
rect 2525 12038 2542 12046
rect 2576 12038 2591 12046
rect 2525 6070 2542 6078
rect 2576 6070 2591 6078
rect 2525 6058 2591 6070
rect 2683 12046 2749 12058
rect 2683 12038 2700 12046
rect 2734 12038 2749 12046
rect 2683 6070 2700 6078
rect 2734 6070 2749 6078
rect 2683 6058 2749 6070
rect 2841 12046 2907 12058
rect 2841 12038 2858 12046
rect 2892 12038 2907 12046
rect 2841 6070 2858 6078
rect 2892 6070 2907 6078
rect 2841 6058 2907 6070
rect 2999 12046 3065 12058
rect 2999 12038 3016 12046
rect 3050 12038 3065 12046
rect 2999 6070 3016 6078
rect 3050 6070 3065 6078
rect 2999 6058 3065 6070
rect 3157 12046 3223 12058
rect 3157 12038 3174 12046
rect 3208 12038 3223 12046
rect 3157 6070 3174 6078
rect 3208 6070 3223 6078
rect 3157 6058 3223 6070
rect 3315 12046 3381 12058
rect 3315 12038 3332 12046
rect 3366 12038 3381 12046
rect 3315 6070 3332 6078
rect 3366 6070 3381 6078
rect 3315 6058 3381 6070
rect 3473 12046 3539 12058
rect 3473 12038 3490 12046
rect 3524 12038 3539 12046
rect 3473 6070 3490 6078
rect 3524 6070 3539 6078
rect 3473 6058 3539 6070
rect 3631 12046 3697 12058
rect 3631 12038 3648 12046
rect 3682 12038 3697 12046
rect 3631 6070 3648 6078
rect 3682 6070 3697 6078
rect 3631 6058 3697 6070
rect 3789 12046 3855 12058
rect 3789 12038 3806 12046
rect 3840 12038 3855 12046
rect 3789 6070 3806 6078
rect 3840 6070 3855 6078
rect 3789 6058 3855 6070
rect 3947 12046 4013 12058
rect 3947 12038 3964 12046
rect 3998 12038 4013 12046
rect 3947 6070 3964 6078
rect 3998 6070 4013 6078
rect 3947 6058 4013 6070
rect 4105 12046 4171 12058
rect 4105 12038 4122 12046
rect 4156 12038 4171 12046
rect 4105 6070 4122 6078
rect 4156 6070 4171 6078
rect 4105 6058 4171 6070
rect -568 6020 -548 6026
rect 4086 6020 4106 6026
rect -568 5986 -556 6020
rect 4094 5986 4106 6020
rect -568 5926 -548 5986
rect 4086 5926 4106 5986
rect -770 5894 -700 5900
rect 4240 5894 4310 5900
rect -770 5884 4310 5894
rect -770 5846 -564 5884
rect 4102 5846 4310 5884
rect -770 5830 4310 5846
rect 5530 12270 10610 12280
rect 5530 12232 5736 12270
rect 10459 12232 10610 12270
rect 5530 12222 10610 12232
rect 5530 12220 5600 12222
rect 10540 12220 10610 12222
rect 5732 12130 5752 12190
rect 10386 12130 10406 12190
rect 5732 12096 5744 12130
rect 10394 12096 10406 12130
rect 5732 12090 5752 12096
rect 10386 12090 10406 12096
rect 5665 12046 5731 12058
rect 5665 12038 5682 12046
rect 5716 12038 5731 12046
rect 5665 6070 5682 6078
rect 5716 6070 5731 6078
rect 5665 6058 5731 6070
rect 5823 12046 5889 12058
rect 5823 12038 5840 12046
rect 5874 12038 5889 12046
rect 5823 6070 5840 6078
rect 5874 6070 5889 6078
rect 5823 6058 5889 6070
rect 5981 12046 6047 12058
rect 5981 12038 5998 12046
rect 6032 12038 6047 12046
rect 5981 6070 5998 6078
rect 6032 6070 6047 6078
rect 5981 6058 6047 6070
rect 6139 12046 6205 12058
rect 6139 12038 6156 12046
rect 6190 12038 6205 12046
rect 6139 6070 6156 6078
rect 6190 6070 6205 6078
rect 6139 6058 6205 6070
rect 6297 12046 6363 12058
rect 6297 12038 6314 12046
rect 6348 12038 6363 12046
rect 6297 6070 6314 6078
rect 6348 6070 6363 6078
rect 6297 6058 6363 6070
rect 6455 12046 6521 12058
rect 6455 12038 6472 12046
rect 6506 12038 6521 12046
rect 6455 6070 6472 6078
rect 6506 6070 6521 6078
rect 6455 6058 6521 6070
rect 6613 12046 6679 12058
rect 6613 12038 6630 12046
rect 6664 12038 6679 12046
rect 6613 6070 6630 6078
rect 6664 6070 6679 6078
rect 6613 6058 6679 6070
rect 6771 12046 6837 12058
rect 6771 12038 6788 12046
rect 6822 12038 6837 12046
rect 6771 6070 6788 6078
rect 6822 6070 6837 6078
rect 6771 6058 6837 6070
rect 6929 12046 6995 12058
rect 6929 12038 6946 12046
rect 6980 12038 6995 12046
rect 6929 6070 6946 6078
rect 6980 6070 6995 6078
rect 6929 6058 6995 6070
rect 7087 12046 7153 12058
rect 7087 12038 7104 12046
rect 7138 12038 7153 12046
rect 7087 6070 7104 6078
rect 7138 6070 7153 6078
rect 7087 6058 7153 6070
rect 7245 12046 7311 12058
rect 7245 12038 7262 12046
rect 7296 12038 7311 12046
rect 7245 6070 7262 6078
rect 7296 6070 7311 6078
rect 7245 6058 7311 6070
rect 7403 12046 7469 12058
rect 7403 12038 7420 12046
rect 7454 12038 7469 12046
rect 7403 6070 7420 6078
rect 7454 6070 7469 6078
rect 7403 6058 7469 6070
rect 7561 12046 7627 12058
rect 7561 12038 7578 12046
rect 7612 12038 7627 12046
rect 7561 6070 7578 6078
rect 7612 6070 7627 6078
rect 7561 6058 7627 6070
rect 7719 12046 7785 12058
rect 7719 12038 7736 12046
rect 7770 12038 7785 12046
rect 7719 6070 7736 6078
rect 7770 6070 7785 6078
rect 7719 6058 7785 6070
rect 7877 12046 7943 12058
rect 7877 12038 7894 12046
rect 7928 12038 7943 12046
rect 7877 6070 7894 6078
rect 7928 6070 7943 6078
rect 7877 6058 7943 6070
rect 8035 12046 8101 12058
rect 8035 12038 8052 12046
rect 8086 12038 8101 12046
rect 8035 6070 8052 6078
rect 8086 6070 8101 6078
rect 8035 6058 8101 6070
rect 8193 12046 8259 12058
rect 8193 12038 8210 12046
rect 8244 12038 8259 12046
rect 8193 6070 8210 6078
rect 8244 6070 8259 6078
rect 8193 6058 8259 6070
rect 8351 12046 8417 12058
rect 8351 12038 8368 12046
rect 8402 12038 8417 12046
rect 8351 6070 8368 6078
rect 8402 6070 8417 6078
rect 8351 6058 8417 6070
rect 8509 12046 8575 12058
rect 8509 12038 8526 12046
rect 8560 12038 8575 12046
rect 8509 6070 8526 6078
rect 8560 6070 8575 6078
rect 8509 6058 8575 6070
rect 8667 12046 8733 12058
rect 8667 12038 8684 12046
rect 8718 12038 8733 12046
rect 8667 6070 8684 6078
rect 8718 6070 8733 6078
rect 8667 6058 8733 6070
rect 8825 12046 8891 12058
rect 8825 12038 8842 12046
rect 8876 12038 8891 12046
rect 8825 6070 8842 6078
rect 8876 6070 8891 6078
rect 8825 6058 8891 6070
rect 8983 12046 9049 12058
rect 8983 12038 9000 12046
rect 9034 12038 9049 12046
rect 8983 6070 9000 6078
rect 9034 6070 9049 6078
rect 8983 6058 9049 6070
rect 9141 12046 9207 12058
rect 9141 12038 9158 12046
rect 9192 12038 9207 12046
rect 9141 6070 9158 6078
rect 9192 6070 9207 6078
rect 9141 6058 9207 6070
rect 9299 12046 9365 12058
rect 9299 12038 9316 12046
rect 9350 12038 9365 12046
rect 9299 6070 9316 6078
rect 9350 6070 9365 6078
rect 9299 6058 9365 6070
rect 9457 12046 9523 12058
rect 9457 12038 9474 12046
rect 9508 12038 9523 12046
rect 9457 6070 9474 6078
rect 9508 6070 9523 6078
rect 9457 6058 9523 6070
rect 9615 12046 9681 12058
rect 9615 12038 9632 12046
rect 9666 12038 9681 12046
rect 9615 6070 9632 6078
rect 9666 6070 9681 6078
rect 9615 6058 9681 6070
rect 9773 12046 9839 12058
rect 9773 12038 9790 12046
rect 9824 12038 9839 12046
rect 9773 6070 9790 6078
rect 9824 6070 9839 6078
rect 9773 6058 9839 6070
rect 9931 12046 9997 12058
rect 9931 12038 9948 12046
rect 9982 12038 9997 12046
rect 9931 6070 9948 6078
rect 9982 6070 9997 6078
rect 9931 6058 9997 6070
rect 10089 12046 10155 12058
rect 10089 12038 10106 12046
rect 10140 12038 10155 12046
rect 10089 6070 10106 6078
rect 10140 6070 10155 6078
rect 10089 6058 10155 6070
rect 10247 12046 10313 12058
rect 10247 12038 10264 12046
rect 10298 12038 10313 12046
rect 10247 6070 10264 6078
rect 10298 6070 10313 6078
rect 10247 6058 10313 6070
rect 10405 12046 10471 12058
rect 10405 12038 10422 12046
rect 10456 12038 10471 12046
rect 10405 6070 10422 6078
rect 10456 6070 10471 6078
rect 10405 6058 10471 6070
rect 5732 6020 5752 6026
rect 10386 6020 10406 6026
rect 5732 5986 5744 6020
rect 10394 5986 10406 6020
rect 5732 5926 5752 5986
rect 10386 5926 10406 5986
rect 5530 5894 5600 5900
rect 10540 5894 10610 5900
rect 5530 5884 10610 5894
rect 5530 5846 5736 5884
rect 10402 5846 10610 5884
rect 5530 5830 10610 5846
<< via1 >>
rect -13370 49680 -13300 49820
rect -13148 49730 -8514 49790
rect -13148 49696 -13088 49730
rect -13088 49696 -12998 49730
rect -12998 49696 -12930 49730
rect -12930 49696 -12840 49730
rect -12840 49696 -12772 49730
rect -12772 49696 -12682 49730
rect -12682 49696 -12614 49730
rect -12614 49696 -12524 49730
rect -12524 49696 -12456 49730
rect -12456 49696 -12366 49730
rect -12366 49696 -12298 49730
rect -12298 49696 -12208 49730
rect -12208 49696 -12140 49730
rect -12140 49696 -12050 49730
rect -12050 49696 -11982 49730
rect -11982 49696 -11892 49730
rect -11892 49696 -11824 49730
rect -11824 49696 -11734 49730
rect -11734 49696 -11666 49730
rect -11666 49696 -11576 49730
rect -11576 49696 -11508 49730
rect -11508 49696 -11418 49730
rect -11418 49696 -11350 49730
rect -11350 49696 -11260 49730
rect -11260 49696 -11192 49730
rect -11192 49696 -11102 49730
rect -11102 49696 -11034 49730
rect -11034 49696 -10944 49730
rect -10944 49696 -10876 49730
rect -10876 49696 -10786 49730
rect -10786 49696 -10718 49730
rect -10718 49696 -10628 49730
rect -10628 49696 -10560 49730
rect -10560 49696 -10470 49730
rect -10470 49696 -10402 49730
rect -10402 49696 -10312 49730
rect -10312 49696 -10244 49730
rect -10244 49696 -10154 49730
rect -10154 49696 -10086 49730
rect -10086 49696 -9996 49730
rect -9996 49696 -9928 49730
rect -9928 49696 -9838 49730
rect -9838 49696 -9770 49730
rect -9770 49696 -9680 49730
rect -9680 49696 -9612 49730
rect -9612 49696 -9522 49730
rect -9522 49696 -9454 49730
rect -9454 49696 -9364 49730
rect -9364 49696 -9296 49730
rect -9296 49696 -9206 49730
rect -9206 49696 -9138 49730
rect -9138 49696 -9048 49730
rect -9048 49696 -8980 49730
rect -8980 49696 -8890 49730
rect -8890 49696 -8822 49730
rect -8822 49696 -8732 49730
rect -8732 49696 -8664 49730
rect -8664 49696 -8574 49730
rect -8574 49696 -8514 49730
rect -13148 49690 -8514 49696
rect -13370 43636 -13354 49680
rect -13354 43636 -13316 49680
rect -13316 43636 -13300 49680
rect -8360 49680 -8290 49820
rect -13235 43678 -13218 49638
rect -13218 43678 -13184 49638
rect -13184 43678 -13169 49638
rect -13077 43678 -13060 49638
rect -13060 43678 -13026 49638
rect -13026 43678 -13011 49638
rect -12919 43678 -12902 49638
rect -12902 43678 -12868 49638
rect -12868 43678 -12853 49638
rect -12761 43678 -12744 49638
rect -12744 43678 -12710 49638
rect -12710 43678 -12695 49638
rect -12603 43678 -12586 49638
rect -12586 43678 -12552 49638
rect -12552 43678 -12537 49638
rect -12445 43678 -12428 49638
rect -12428 43678 -12394 49638
rect -12394 43678 -12379 49638
rect -12287 43678 -12270 49638
rect -12270 43678 -12236 49638
rect -12236 43678 -12221 49638
rect -12129 43678 -12112 49638
rect -12112 43678 -12078 49638
rect -12078 43678 -12063 49638
rect -11971 43678 -11954 49638
rect -11954 43678 -11920 49638
rect -11920 43678 -11905 49638
rect -11813 43678 -11796 49638
rect -11796 43678 -11762 49638
rect -11762 43678 -11747 49638
rect -11655 43678 -11638 49638
rect -11638 43678 -11604 49638
rect -11604 43678 -11589 49638
rect -11497 43678 -11480 49638
rect -11480 43678 -11446 49638
rect -11446 43678 -11431 49638
rect -11339 43678 -11322 49638
rect -11322 43678 -11288 49638
rect -11288 43678 -11273 49638
rect -11181 43678 -11164 49638
rect -11164 43678 -11130 49638
rect -11130 43678 -11115 49638
rect -11023 43678 -11006 49638
rect -11006 43678 -10972 49638
rect -10972 43678 -10957 49638
rect -10865 43678 -10848 49638
rect -10848 43678 -10814 49638
rect -10814 43678 -10799 49638
rect -10707 43678 -10690 49638
rect -10690 43678 -10656 49638
rect -10656 43678 -10641 49638
rect -10549 43678 -10532 49638
rect -10532 43678 -10498 49638
rect -10498 43678 -10483 49638
rect -10391 43678 -10374 49638
rect -10374 43678 -10340 49638
rect -10340 43678 -10325 49638
rect -10233 43678 -10216 49638
rect -10216 43678 -10182 49638
rect -10182 43678 -10167 49638
rect -10075 43678 -10058 49638
rect -10058 43678 -10024 49638
rect -10024 43678 -10009 49638
rect -9917 43678 -9900 49638
rect -9900 43678 -9866 49638
rect -9866 43678 -9851 49638
rect -9759 43678 -9742 49638
rect -9742 43678 -9708 49638
rect -9708 43678 -9693 49638
rect -9601 43678 -9584 49638
rect -9584 43678 -9550 49638
rect -9550 43678 -9535 49638
rect -9443 43678 -9426 49638
rect -9426 43678 -9392 49638
rect -9392 43678 -9377 49638
rect -9285 43678 -9268 49638
rect -9268 43678 -9234 49638
rect -9234 43678 -9219 49638
rect -9127 43678 -9110 49638
rect -9110 43678 -9076 49638
rect -9076 43678 -9061 49638
rect -8969 43678 -8952 49638
rect -8952 43678 -8918 49638
rect -8918 43678 -8903 49638
rect -8811 43678 -8794 49638
rect -8794 43678 -8760 49638
rect -8760 43678 -8745 49638
rect -8653 43678 -8636 49638
rect -8636 43678 -8602 49638
rect -8602 43678 -8587 49638
rect -8495 43678 -8478 49638
rect -8478 43678 -8444 49638
rect -8444 43678 -8429 49638
rect -13370 43500 -13300 43636
rect -8360 43636 -8346 49680
rect -8346 43636 -8308 49680
rect -8308 43636 -8290 49680
rect -13148 43620 -8514 43626
rect -13148 43586 -13088 43620
rect -13088 43586 -12998 43620
rect -12998 43586 -12930 43620
rect -12930 43586 -12840 43620
rect -12840 43586 -12772 43620
rect -12772 43586 -12682 43620
rect -12682 43586 -12614 43620
rect -12614 43586 -12524 43620
rect -12524 43586 -12456 43620
rect -12456 43586 -12366 43620
rect -12366 43586 -12298 43620
rect -12298 43586 -12208 43620
rect -12208 43586 -12140 43620
rect -12140 43586 -12050 43620
rect -12050 43586 -11982 43620
rect -11982 43586 -11892 43620
rect -11892 43586 -11824 43620
rect -11824 43586 -11734 43620
rect -11734 43586 -11666 43620
rect -11666 43586 -11576 43620
rect -11576 43586 -11508 43620
rect -11508 43586 -11418 43620
rect -11418 43586 -11350 43620
rect -11350 43586 -11260 43620
rect -11260 43586 -11192 43620
rect -11192 43586 -11102 43620
rect -11102 43586 -11034 43620
rect -11034 43586 -10944 43620
rect -10944 43586 -10876 43620
rect -10876 43586 -10786 43620
rect -10786 43586 -10718 43620
rect -10718 43586 -10628 43620
rect -10628 43586 -10560 43620
rect -10560 43586 -10470 43620
rect -10470 43586 -10402 43620
rect -10402 43586 -10312 43620
rect -10312 43586 -10244 43620
rect -10244 43586 -10154 43620
rect -10154 43586 -10086 43620
rect -10086 43586 -9996 43620
rect -9996 43586 -9928 43620
rect -9928 43586 -9838 43620
rect -9838 43586 -9770 43620
rect -9770 43586 -9680 43620
rect -9680 43586 -9612 43620
rect -9612 43586 -9522 43620
rect -9522 43586 -9454 43620
rect -9454 43586 -9364 43620
rect -9364 43586 -9296 43620
rect -9296 43586 -9206 43620
rect -9206 43586 -9138 43620
rect -9138 43586 -9048 43620
rect -9048 43586 -8980 43620
rect -8980 43586 -8890 43620
rect -8890 43586 -8822 43620
rect -8822 43586 -8732 43620
rect -8732 43586 -8664 43620
rect -8664 43586 -8574 43620
rect -8574 43586 -8514 43620
rect -13148 43526 -8514 43586
rect -8360 43500 -8290 43636
rect -7070 49680 -7000 49820
rect -6848 49730 -2214 49790
rect -6848 49696 -6788 49730
rect -6788 49696 -6698 49730
rect -6698 49696 -6630 49730
rect -6630 49696 -6540 49730
rect -6540 49696 -6472 49730
rect -6472 49696 -6382 49730
rect -6382 49696 -6314 49730
rect -6314 49696 -6224 49730
rect -6224 49696 -6156 49730
rect -6156 49696 -6066 49730
rect -6066 49696 -5998 49730
rect -5998 49696 -5908 49730
rect -5908 49696 -5840 49730
rect -5840 49696 -5750 49730
rect -5750 49696 -5682 49730
rect -5682 49696 -5592 49730
rect -5592 49696 -5524 49730
rect -5524 49696 -5434 49730
rect -5434 49696 -5366 49730
rect -5366 49696 -5276 49730
rect -5276 49696 -5208 49730
rect -5208 49696 -5118 49730
rect -5118 49696 -5050 49730
rect -5050 49696 -4960 49730
rect -4960 49696 -4892 49730
rect -4892 49696 -4802 49730
rect -4802 49696 -4734 49730
rect -4734 49696 -4644 49730
rect -4644 49696 -4576 49730
rect -4576 49696 -4486 49730
rect -4486 49696 -4418 49730
rect -4418 49696 -4328 49730
rect -4328 49696 -4260 49730
rect -4260 49696 -4170 49730
rect -4170 49696 -4102 49730
rect -4102 49696 -4012 49730
rect -4012 49696 -3944 49730
rect -3944 49696 -3854 49730
rect -3854 49696 -3786 49730
rect -3786 49696 -3696 49730
rect -3696 49696 -3628 49730
rect -3628 49696 -3538 49730
rect -3538 49696 -3470 49730
rect -3470 49696 -3380 49730
rect -3380 49696 -3312 49730
rect -3312 49696 -3222 49730
rect -3222 49696 -3154 49730
rect -3154 49696 -3064 49730
rect -3064 49696 -2996 49730
rect -2996 49696 -2906 49730
rect -2906 49696 -2838 49730
rect -2838 49696 -2748 49730
rect -2748 49696 -2680 49730
rect -2680 49696 -2590 49730
rect -2590 49696 -2522 49730
rect -2522 49696 -2432 49730
rect -2432 49696 -2364 49730
rect -2364 49696 -2274 49730
rect -2274 49696 -2214 49730
rect -6848 49690 -2214 49696
rect -7070 43636 -7054 49680
rect -7054 43636 -7016 49680
rect -7016 43636 -7000 49680
rect -2060 49680 -1990 49820
rect -6935 43678 -6918 49638
rect -6918 43678 -6884 49638
rect -6884 43678 -6869 49638
rect -6777 43678 -6760 49638
rect -6760 43678 -6726 49638
rect -6726 43678 -6711 49638
rect -6619 43678 -6602 49638
rect -6602 43678 -6568 49638
rect -6568 43678 -6553 49638
rect -6461 43678 -6444 49638
rect -6444 43678 -6410 49638
rect -6410 43678 -6395 49638
rect -6303 43678 -6286 49638
rect -6286 43678 -6252 49638
rect -6252 43678 -6237 49638
rect -6145 43678 -6128 49638
rect -6128 43678 -6094 49638
rect -6094 43678 -6079 49638
rect -5987 43678 -5970 49638
rect -5970 43678 -5936 49638
rect -5936 43678 -5921 49638
rect -5829 43678 -5812 49638
rect -5812 43678 -5778 49638
rect -5778 43678 -5763 49638
rect -5671 43678 -5654 49638
rect -5654 43678 -5620 49638
rect -5620 43678 -5605 49638
rect -5513 43678 -5496 49638
rect -5496 43678 -5462 49638
rect -5462 43678 -5447 49638
rect -5355 43678 -5338 49638
rect -5338 43678 -5304 49638
rect -5304 43678 -5289 49638
rect -5197 43678 -5180 49638
rect -5180 43678 -5146 49638
rect -5146 43678 -5131 49638
rect -5039 43678 -5022 49638
rect -5022 43678 -4988 49638
rect -4988 43678 -4973 49638
rect -4881 43678 -4864 49638
rect -4864 43678 -4830 49638
rect -4830 43678 -4815 49638
rect -4723 43678 -4706 49638
rect -4706 43678 -4672 49638
rect -4672 43678 -4657 49638
rect -4565 43678 -4548 49638
rect -4548 43678 -4514 49638
rect -4514 43678 -4499 49638
rect -4407 43678 -4390 49638
rect -4390 43678 -4356 49638
rect -4356 43678 -4341 49638
rect -4249 43678 -4232 49638
rect -4232 43678 -4198 49638
rect -4198 43678 -4183 49638
rect -4091 43678 -4074 49638
rect -4074 43678 -4040 49638
rect -4040 43678 -4025 49638
rect -3933 43678 -3916 49638
rect -3916 43678 -3882 49638
rect -3882 43678 -3867 49638
rect -3775 43678 -3758 49638
rect -3758 43678 -3724 49638
rect -3724 43678 -3709 49638
rect -3617 43678 -3600 49638
rect -3600 43678 -3566 49638
rect -3566 43678 -3551 49638
rect -3459 43678 -3442 49638
rect -3442 43678 -3408 49638
rect -3408 43678 -3393 49638
rect -3301 43678 -3284 49638
rect -3284 43678 -3250 49638
rect -3250 43678 -3235 49638
rect -3143 43678 -3126 49638
rect -3126 43678 -3092 49638
rect -3092 43678 -3077 49638
rect -2985 43678 -2968 49638
rect -2968 43678 -2934 49638
rect -2934 43678 -2919 49638
rect -2827 43678 -2810 49638
rect -2810 43678 -2776 49638
rect -2776 43678 -2761 49638
rect -2669 43678 -2652 49638
rect -2652 43678 -2618 49638
rect -2618 43678 -2603 49638
rect -2511 43678 -2494 49638
rect -2494 43678 -2460 49638
rect -2460 43678 -2445 49638
rect -2353 43678 -2336 49638
rect -2336 43678 -2302 49638
rect -2302 43678 -2287 49638
rect -2195 43678 -2178 49638
rect -2178 43678 -2144 49638
rect -2144 43678 -2129 49638
rect -7070 43500 -7000 43636
rect -2060 43636 -2046 49680
rect -2046 43636 -2008 49680
rect -2008 43636 -1990 49680
rect -6848 43620 -2214 43626
rect -6848 43586 -6788 43620
rect -6788 43586 -6698 43620
rect -6698 43586 -6630 43620
rect -6630 43586 -6540 43620
rect -6540 43586 -6472 43620
rect -6472 43586 -6382 43620
rect -6382 43586 -6314 43620
rect -6314 43586 -6224 43620
rect -6224 43586 -6156 43620
rect -6156 43586 -6066 43620
rect -6066 43586 -5998 43620
rect -5998 43586 -5908 43620
rect -5908 43586 -5840 43620
rect -5840 43586 -5750 43620
rect -5750 43586 -5682 43620
rect -5682 43586 -5592 43620
rect -5592 43586 -5524 43620
rect -5524 43586 -5434 43620
rect -5434 43586 -5366 43620
rect -5366 43586 -5276 43620
rect -5276 43586 -5208 43620
rect -5208 43586 -5118 43620
rect -5118 43586 -5050 43620
rect -5050 43586 -4960 43620
rect -4960 43586 -4892 43620
rect -4892 43586 -4802 43620
rect -4802 43586 -4734 43620
rect -4734 43586 -4644 43620
rect -4644 43586 -4576 43620
rect -4576 43586 -4486 43620
rect -4486 43586 -4418 43620
rect -4418 43586 -4328 43620
rect -4328 43586 -4260 43620
rect -4260 43586 -4170 43620
rect -4170 43586 -4102 43620
rect -4102 43586 -4012 43620
rect -4012 43586 -3944 43620
rect -3944 43586 -3854 43620
rect -3854 43586 -3786 43620
rect -3786 43586 -3696 43620
rect -3696 43586 -3628 43620
rect -3628 43586 -3538 43620
rect -3538 43586 -3470 43620
rect -3470 43586 -3380 43620
rect -3380 43586 -3312 43620
rect -3312 43586 -3222 43620
rect -3222 43586 -3154 43620
rect -3154 43586 -3064 43620
rect -3064 43586 -2996 43620
rect -2996 43586 -2906 43620
rect -2906 43586 -2838 43620
rect -2838 43586 -2748 43620
rect -2748 43586 -2680 43620
rect -2680 43586 -2590 43620
rect -2590 43586 -2522 43620
rect -2522 43586 -2432 43620
rect -2432 43586 -2364 43620
rect -2364 43586 -2274 43620
rect -2274 43586 -2214 43620
rect -6848 43526 -2214 43586
rect -2060 43500 -1990 43636
rect -770 49680 -700 49820
rect -548 49730 4086 49790
rect -548 49696 -488 49730
rect -488 49696 -398 49730
rect -398 49696 -330 49730
rect -330 49696 -240 49730
rect -240 49696 -172 49730
rect -172 49696 -82 49730
rect -82 49696 -14 49730
rect -14 49696 76 49730
rect 76 49696 144 49730
rect 144 49696 234 49730
rect 234 49696 302 49730
rect 302 49696 392 49730
rect 392 49696 460 49730
rect 460 49696 550 49730
rect 550 49696 618 49730
rect 618 49696 708 49730
rect 708 49696 776 49730
rect 776 49696 866 49730
rect 866 49696 934 49730
rect 934 49696 1024 49730
rect 1024 49696 1092 49730
rect 1092 49696 1182 49730
rect 1182 49696 1250 49730
rect 1250 49696 1340 49730
rect 1340 49696 1408 49730
rect 1408 49696 1498 49730
rect 1498 49696 1566 49730
rect 1566 49696 1656 49730
rect 1656 49696 1724 49730
rect 1724 49696 1814 49730
rect 1814 49696 1882 49730
rect 1882 49696 1972 49730
rect 1972 49696 2040 49730
rect 2040 49696 2130 49730
rect 2130 49696 2198 49730
rect 2198 49696 2288 49730
rect 2288 49696 2356 49730
rect 2356 49696 2446 49730
rect 2446 49696 2514 49730
rect 2514 49696 2604 49730
rect 2604 49696 2672 49730
rect 2672 49696 2762 49730
rect 2762 49696 2830 49730
rect 2830 49696 2920 49730
rect 2920 49696 2988 49730
rect 2988 49696 3078 49730
rect 3078 49696 3146 49730
rect 3146 49696 3236 49730
rect 3236 49696 3304 49730
rect 3304 49696 3394 49730
rect 3394 49696 3462 49730
rect 3462 49696 3552 49730
rect 3552 49696 3620 49730
rect 3620 49696 3710 49730
rect 3710 49696 3778 49730
rect 3778 49696 3868 49730
rect 3868 49696 3936 49730
rect 3936 49696 4026 49730
rect 4026 49696 4086 49730
rect -548 49690 4086 49696
rect -770 43636 -754 49680
rect -754 43636 -716 49680
rect -716 43636 -700 49680
rect 4240 49680 4310 49820
rect -635 43678 -618 49638
rect -618 43678 -584 49638
rect -584 43678 -569 49638
rect -477 43678 -460 49638
rect -460 43678 -426 49638
rect -426 43678 -411 49638
rect -319 43678 -302 49638
rect -302 43678 -268 49638
rect -268 43678 -253 49638
rect -161 43678 -144 49638
rect -144 43678 -110 49638
rect -110 43678 -95 49638
rect -3 43678 14 49638
rect 14 43678 48 49638
rect 48 43678 63 49638
rect 155 43678 172 49638
rect 172 43678 206 49638
rect 206 43678 221 49638
rect 313 43678 330 49638
rect 330 43678 364 49638
rect 364 43678 379 49638
rect 471 43678 488 49638
rect 488 43678 522 49638
rect 522 43678 537 49638
rect 629 43678 646 49638
rect 646 43678 680 49638
rect 680 43678 695 49638
rect 787 43678 804 49638
rect 804 43678 838 49638
rect 838 43678 853 49638
rect 945 43678 962 49638
rect 962 43678 996 49638
rect 996 43678 1011 49638
rect 1103 43678 1120 49638
rect 1120 43678 1154 49638
rect 1154 43678 1169 49638
rect 1261 43678 1278 49638
rect 1278 43678 1312 49638
rect 1312 43678 1327 49638
rect 1419 43678 1436 49638
rect 1436 43678 1470 49638
rect 1470 43678 1485 49638
rect 1577 43678 1594 49638
rect 1594 43678 1628 49638
rect 1628 43678 1643 49638
rect 1735 43678 1752 49638
rect 1752 43678 1786 49638
rect 1786 43678 1801 49638
rect 1893 43678 1910 49638
rect 1910 43678 1944 49638
rect 1944 43678 1959 49638
rect 2051 43678 2068 49638
rect 2068 43678 2102 49638
rect 2102 43678 2117 49638
rect 2209 43678 2226 49638
rect 2226 43678 2260 49638
rect 2260 43678 2275 49638
rect 2367 43678 2384 49638
rect 2384 43678 2418 49638
rect 2418 43678 2433 49638
rect 2525 43678 2542 49638
rect 2542 43678 2576 49638
rect 2576 43678 2591 49638
rect 2683 43678 2700 49638
rect 2700 43678 2734 49638
rect 2734 43678 2749 49638
rect 2841 43678 2858 49638
rect 2858 43678 2892 49638
rect 2892 43678 2907 49638
rect 2999 43678 3016 49638
rect 3016 43678 3050 49638
rect 3050 43678 3065 49638
rect 3157 43678 3174 49638
rect 3174 43678 3208 49638
rect 3208 43678 3223 49638
rect 3315 43678 3332 49638
rect 3332 43678 3366 49638
rect 3366 43678 3381 49638
rect 3473 43678 3490 49638
rect 3490 43678 3524 49638
rect 3524 43678 3539 49638
rect 3631 43678 3648 49638
rect 3648 43678 3682 49638
rect 3682 43678 3697 49638
rect 3789 43678 3806 49638
rect 3806 43678 3840 49638
rect 3840 43678 3855 49638
rect 3947 43678 3964 49638
rect 3964 43678 3998 49638
rect 3998 43678 4013 49638
rect 4105 43678 4122 49638
rect 4122 43678 4156 49638
rect 4156 43678 4171 49638
rect -770 43500 -700 43636
rect 4240 43636 4254 49680
rect 4254 43636 4292 49680
rect 4292 43636 4310 49680
rect -548 43620 4086 43626
rect -548 43586 -488 43620
rect -488 43586 -398 43620
rect -398 43586 -330 43620
rect -330 43586 -240 43620
rect -240 43586 -172 43620
rect -172 43586 -82 43620
rect -82 43586 -14 43620
rect -14 43586 76 43620
rect 76 43586 144 43620
rect 144 43586 234 43620
rect 234 43586 302 43620
rect 302 43586 392 43620
rect 392 43586 460 43620
rect 460 43586 550 43620
rect 550 43586 618 43620
rect 618 43586 708 43620
rect 708 43586 776 43620
rect 776 43586 866 43620
rect 866 43586 934 43620
rect 934 43586 1024 43620
rect 1024 43586 1092 43620
rect 1092 43586 1182 43620
rect 1182 43586 1250 43620
rect 1250 43586 1340 43620
rect 1340 43586 1408 43620
rect 1408 43586 1498 43620
rect 1498 43586 1566 43620
rect 1566 43586 1656 43620
rect 1656 43586 1724 43620
rect 1724 43586 1814 43620
rect 1814 43586 1882 43620
rect 1882 43586 1972 43620
rect 1972 43586 2040 43620
rect 2040 43586 2130 43620
rect 2130 43586 2198 43620
rect 2198 43586 2288 43620
rect 2288 43586 2356 43620
rect 2356 43586 2446 43620
rect 2446 43586 2514 43620
rect 2514 43586 2604 43620
rect 2604 43586 2672 43620
rect 2672 43586 2762 43620
rect 2762 43586 2830 43620
rect 2830 43586 2920 43620
rect 2920 43586 2988 43620
rect 2988 43586 3078 43620
rect 3078 43586 3146 43620
rect 3146 43586 3236 43620
rect 3236 43586 3304 43620
rect 3304 43586 3394 43620
rect 3394 43586 3462 43620
rect 3462 43586 3552 43620
rect 3552 43586 3620 43620
rect 3620 43586 3710 43620
rect 3710 43586 3778 43620
rect 3778 43586 3868 43620
rect 3868 43586 3936 43620
rect 3936 43586 4026 43620
rect 4026 43586 4086 43620
rect -548 43526 4086 43586
rect 4240 43500 4310 43636
rect 5530 49680 5600 49820
rect 5752 49730 10386 49790
rect 5752 49696 5812 49730
rect 5812 49696 5902 49730
rect 5902 49696 5970 49730
rect 5970 49696 6060 49730
rect 6060 49696 6128 49730
rect 6128 49696 6218 49730
rect 6218 49696 6286 49730
rect 6286 49696 6376 49730
rect 6376 49696 6444 49730
rect 6444 49696 6534 49730
rect 6534 49696 6602 49730
rect 6602 49696 6692 49730
rect 6692 49696 6760 49730
rect 6760 49696 6850 49730
rect 6850 49696 6918 49730
rect 6918 49696 7008 49730
rect 7008 49696 7076 49730
rect 7076 49696 7166 49730
rect 7166 49696 7234 49730
rect 7234 49696 7324 49730
rect 7324 49696 7392 49730
rect 7392 49696 7482 49730
rect 7482 49696 7550 49730
rect 7550 49696 7640 49730
rect 7640 49696 7708 49730
rect 7708 49696 7798 49730
rect 7798 49696 7866 49730
rect 7866 49696 7956 49730
rect 7956 49696 8024 49730
rect 8024 49696 8114 49730
rect 8114 49696 8182 49730
rect 8182 49696 8272 49730
rect 8272 49696 8340 49730
rect 8340 49696 8430 49730
rect 8430 49696 8498 49730
rect 8498 49696 8588 49730
rect 8588 49696 8656 49730
rect 8656 49696 8746 49730
rect 8746 49696 8814 49730
rect 8814 49696 8904 49730
rect 8904 49696 8972 49730
rect 8972 49696 9062 49730
rect 9062 49696 9130 49730
rect 9130 49696 9220 49730
rect 9220 49696 9288 49730
rect 9288 49696 9378 49730
rect 9378 49696 9446 49730
rect 9446 49696 9536 49730
rect 9536 49696 9604 49730
rect 9604 49696 9694 49730
rect 9694 49696 9762 49730
rect 9762 49696 9852 49730
rect 9852 49696 9920 49730
rect 9920 49696 10010 49730
rect 10010 49696 10078 49730
rect 10078 49696 10168 49730
rect 10168 49696 10236 49730
rect 10236 49696 10326 49730
rect 10326 49696 10386 49730
rect 5752 49690 10386 49696
rect 5530 43636 5546 49680
rect 5546 43636 5584 49680
rect 5584 43636 5600 49680
rect 10540 49680 10610 49820
rect 5665 43678 5682 49638
rect 5682 43678 5716 49638
rect 5716 43678 5731 49638
rect 5823 43678 5840 49638
rect 5840 43678 5874 49638
rect 5874 43678 5889 49638
rect 5981 43678 5998 49638
rect 5998 43678 6032 49638
rect 6032 43678 6047 49638
rect 6139 43678 6156 49638
rect 6156 43678 6190 49638
rect 6190 43678 6205 49638
rect 6297 43678 6314 49638
rect 6314 43678 6348 49638
rect 6348 43678 6363 49638
rect 6455 43678 6472 49638
rect 6472 43678 6506 49638
rect 6506 43678 6521 49638
rect 6613 43678 6630 49638
rect 6630 43678 6664 49638
rect 6664 43678 6679 49638
rect 6771 43678 6788 49638
rect 6788 43678 6822 49638
rect 6822 43678 6837 49638
rect 6929 43678 6946 49638
rect 6946 43678 6980 49638
rect 6980 43678 6995 49638
rect 7087 43678 7104 49638
rect 7104 43678 7138 49638
rect 7138 43678 7153 49638
rect 7245 43678 7262 49638
rect 7262 43678 7296 49638
rect 7296 43678 7311 49638
rect 7403 43678 7420 49638
rect 7420 43678 7454 49638
rect 7454 43678 7469 49638
rect 7561 43678 7578 49638
rect 7578 43678 7612 49638
rect 7612 43678 7627 49638
rect 7719 43678 7736 49638
rect 7736 43678 7770 49638
rect 7770 43678 7785 49638
rect 7877 43678 7894 49638
rect 7894 43678 7928 49638
rect 7928 43678 7943 49638
rect 8035 43678 8052 49638
rect 8052 43678 8086 49638
rect 8086 43678 8101 49638
rect 8193 43678 8210 49638
rect 8210 43678 8244 49638
rect 8244 43678 8259 49638
rect 8351 43678 8368 49638
rect 8368 43678 8402 49638
rect 8402 43678 8417 49638
rect 8509 43678 8526 49638
rect 8526 43678 8560 49638
rect 8560 43678 8575 49638
rect 8667 43678 8684 49638
rect 8684 43678 8718 49638
rect 8718 43678 8733 49638
rect 8825 43678 8842 49638
rect 8842 43678 8876 49638
rect 8876 43678 8891 49638
rect 8983 43678 9000 49638
rect 9000 43678 9034 49638
rect 9034 43678 9049 49638
rect 9141 43678 9158 49638
rect 9158 43678 9192 49638
rect 9192 43678 9207 49638
rect 9299 43678 9316 49638
rect 9316 43678 9350 49638
rect 9350 43678 9365 49638
rect 9457 43678 9474 49638
rect 9474 43678 9508 49638
rect 9508 43678 9523 49638
rect 9615 43678 9632 49638
rect 9632 43678 9666 49638
rect 9666 43678 9681 49638
rect 9773 43678 9790 49638
rect 9790 43678 9824 49638
rect 9824 43678 9839 49638
rect 9931 43678 9948 49638
rect 9948 43678 9982 49638
rect 9982 43678 9997 49638
rect 10089 43678 10106 49638
rect 10106 43678 10140 49638
rect 10140 43678 10155 49638
rect 10247 43678 10264 49638
rect 10264 43678 10298 49638
rect 10298 43678 10313 49638
rect 10405 43678 10422 49638
rect 10422 43678 10456 49638
rect 10456 43678 10471 49638
rect 5530 43500 5600 43636
rect 10540 43636 10554 49680
rect 10554 43636 10592 49680
rect 10592 43636 10610 49680
rect 5752 43620 10386 43626
rect 5752 43586 5812 43620
rect 5812 43586 5902 43620
rect 5902 43586 5970 43620
rect 5970 43586 6060 43620
rect 6060 43586 6128 43620
rect 6128 43586 6218 43620
rect 6218 43586 6286 43620
rect 6286 43586 6376 43620
rect 6376 43586 6444 43620
rect 6444 43586 6534 43620
rect 6534 43586 6602 43620
rect 6602 43586 6692 43620
rect 6692 43586 6760 43620
rect 6760 43586 6850 43620
rect 6850 43586 6918 43620
rect 6918 43586 7008 43620
rect 7008 43586 7076 43620
rect 7076 43586 7166 43620
rect 7166 43586 7234 43620
rect 7234 43586 7324 43620
rect 7324 43586 7392 43620
rect 7392 43586 7482 43620
rect 7482 43586 7550 43620
rect 7550 43586 7640 43620
rect 7640 43586 7708 43620
rect 7708 43586 7798 43620
rect 7798 43586 7866 43620
rect 7866 43586 7956 43620
rect 7956 43586 8024 43620
rect 8024 43586 8114 43620
rect 8114 43586 8182 43620
rect 8182 43586 8272 43620
rect 8272 43586 8340 43620
rect 8340 43586 8430 43620
rect 8430 43586 8498 43620
rect 8498 43586 8588 43620
rect 8588 43586 8656 43620
rect 8656 43586 8746 43620
rect 8746 43586 8814 43620
rect 8814 43586 8904 43620
rect 8904 43586 8972 43620
rect 8972 43586 9062 43620
rect 9062 43586 9130 43620
rect 9130 43586 9220 43620
rect 9220 43586 9288 43620
rect 9288 43586 9378 43620
rect 9378 43586 9446 43620
rect 9446 43586 9536 43620
rect 9536 43586 9604 43620
rect 9604 43586 9694 43620
rect 9694 43586 9762 43620
rect 9762 43586 9852 43620
rect 9852 43586 9920 43620
rect 9920 43586 10010 43620
rect 10010 43586 10078 43620
rect 10078 43586 10168 43620
rect 10168 43586 10236 43620
rect 10236 43586 10326 43620
rect 10326 43586 10386 43620
rect 5752 43526 10386 43586
rect 10540 43500 10610 43636
rect -13370 42680 -13300 42820
rect -13148 42730 -8514 42790
rect -13148 42696 -13088 42730
rect -13088 42696 -12998 42730
rect -12998 42696 -12930 42730
rect -12930 42696 -12840 42730
rect -12840 42696 -12772 42730
rect -12772 42696 -12682 42730
rect -12682 42696 -12614 42730
rect -12614 42696 -12524 42730
rect -12524 42696 -12456 42730
rect -12456 42696 -12366 42730
rect -12366 42696 -12298 42730
rect -12298 42696 -12208 42730
rect -12208 42696 -12140 42730
rect -12140 42696 -12050 42730
rect -12050 42696 -11982 42730
rect -11982 42696 -11892 42730
rect -11892 42696 -11824 42730
rect -11824 42696 -11734 42730
rect -11734 42696 -11666 42730
rect -11666 42696 -11576 42730
rect -11576 42696 -11508 42730
rect -11508 42696 -11418 42730
rect -11418 42696 -11350 42730
rect -11350 42696 -11260 42730
rect -11260 42696 -11192 42730
rect -11192 42696 -11102 42730
rect -11102 42696 -11034 42730
rect -11034 42696 -10944 42730
rect -10944 42696 -10876 42730
rect -10876 42696 -10786 42730
rect -10786 42696 -10718 42730
rect -10718 42696 -10628 42730
rect -10628 42696 -10560 42730
rect -10560 42696 -10470 42730
rect -10470 42696 -10402 42730
rect -10402 42696 -10312 42730
rect -10312 42696 -10244 42730
rect -10244 42696 -10154 42730
rect -10154 42696 -10086 42730
rect -10086 42696 -9996 42730
rect -9996 42696 -9928 42730
rect -9928 42696 -9838 42730
rect -9838 42696 -9770 42730
rect -9770 42696 -9680 42730
rect -9680 42696 -9612 42730
rect -9612 42696 -9522 42730
rect -9522 42696 -9454 42730
rect -9454 42696 -9364 42730
rect -9364 42696 -9296 42730
rect -9296 42696 -9206 42730
rect -9206 42696 -9138 42730
rect -9138 42696 -9048 42730
rect -9048 42696 -8980 42730
rect -8980 42696 -8890 42730
rect -8890 42696 -8822 42730
rect -8822 42696 -8732 42730
rect -8732 42696 -8664 42730
rect -8664 42696 -8574 42730
rect -8574 42696 -8514 42730
rect -13148 42690 -8514 42696
rect -13370 36636 -13354 42680
rect -13354 36636 -13316 42680
rect -13316 36636 -13300 42680
rect -8360 42680 -8290 42820
rect -13235 36678 -13218 42638
rect -13218 36678 -13184 42638
rect -13184 36678 -13169 42638
rect -13077 36678 -13060 42638
rect -13060 36678 -13026 42638
rect -13026 36678 -13011 42638
rect -12919 36678 -12902 42638
rect -12902 36678 -12868 42638
rect -12868 36678 -12853 42638
rect -12761 36678 -12744 42638
rect -12744 36678 -12710 42638
rect -12710 36678 -12695 42638
rect -12603 36678 -12586 42638
rect -12586 36678 -12552 42638
rect -12552 36678 -12537 42638
rect -12445 36678 -12428 42638
rect -12428 36678 -12394 42638
rect -12394 36678 -12379 42638
rect -12287 36678 -12270 42638
rect -12270 36678 -12236 42638
rect -12236 36678 -12221 42638
rect -12129 36678 -12112 42638
rect -12112 36678 -12078 42638
rect -12078 36678 -12063 42638
rect -11971 36678 -11954 42638
rect -11954 36678 -11920 42638
rect -11920 36678 -11905 42638
rect -11813 36678 -11796 42638
rect -11796 36678 -11762 42638
rect -11762 36678 -11747 42638
rect -11655 36678 -11638 42638
rect -11638 36678 -11604 42638
rect -11604 36678 -11589 42638
rect -11497 36678 -11480 42638
rect -11480 36678 -11446 42638
rect -11446 36678 -11431 42638
rect -11339 36678 -11322 42638
rect -11322 36678 -11288 42638
rect -11288 36678 -11273 42638
rect -11181 36678 -11164 42638
rect -11164 36678 -11130 42638
rect -11130 36678 -11115 42638
rect -11023 36678 -11006 42638
rect -11006 36678 -10972 42638
rect -10972 36678 -10957 42638
rect -10865 36678 -10848 42638
rect -10848 36678 -10814 42638
rect -10814 36678 -10799 42638
rect -10707 36678 -10690 42638
rect -10690 36678 -10656 42638
rect -10656 36678 -10641 42638
rect -10549 36678 -10532 42638
rect -10532 36678 -10498 42638
rect -10498 36678 -10483 42638
rect -10391 36678 -10374 42638
rect -10374 36678 -10340 42638
rect -10340 36678 -10325 42638
rect -10233 36678 -10216 42638
rect -10216 36678 -10182 42638
rect -10182 36678 -10167 42638
rect -10075 36678 -10058 42638
rect -10058 36678 -10024 42638
rect -10024 36678 -10009 42638
rect -9917 36678 -9900 42638
rect -9900 36678 -9866 42638
rect -9866 36678 -9851 42638
rect -9759 36678 -9742 42638
rect -9742 36678 -9708 42638
rect -9708 36678 -9693 42638
rect -9601 36678 -9584 42638
rect -9584 36678 -9550 42638
rect -9550 36678 -9535 42638
rect -9443 36678 -9426 42638
rect -9426 36678 -9392 42638
rect -9392 36678 -9377 42638
rect -9285 36678 -9268 42638
rect -9268 36678 -9234 42638
rect -9234 36678 -9219 42638
rect -9127 36678 -9110 42638
rect -9110 36678 -9076 42638
rect -9076 36678 -9061 42638
rect -8969 36678 -8952 42638
rect -8952 36678 -8918 42638
rect -8918 36678 -8903 42638
rect -8811 36678 -8794 42638
rect -8794 36678 -8760 42638
rect -8760 36678 -8745 42638
rect -8653 36678 -8636 42638
rect -8636 36678 -8602 42638
rect -8602 36678 -8587 42638
rect -8495 36678 -8478 42638
rect -8478 36678 -8444 42638
rect -8444 36678 -8429 42638
rect -13370 36500 -13300 36636
rect -8360 36636 -8346 42680
rect -8346 36636 -8308 42680
rect -8308 36636 -8290 42680
rect -13148 36620 -8514 36626
rect -13148 36586 -13088 36620
rect -13088 36586 -12998 36620
rect -12998 36586 -12930 36620
rect -12930 36586 -12840 36620
rect -12840 36586 -12772 36620
rect -12772 36586 -12682 36620
rect -12682 36586 -12614 36620
rect -12614 36586 -12524 36620
rect -12524 36586 -12456 36620
rect -12456 36586 -12366 36620
rect -12366 36586 -12298 36620
rect -12298 36586 -12208 36620
rect -12208 36586 -12140 36620
rect -12140 36586 -12050 36620
rect -12050 36586 -11982 36620
rect -11982 36586 -11892 36620
rect -11892 36586 -11824 36620
rect -11824 36586 -11734 36620
rect -11734 36586 -11666 36620
rect -11666 36586 -11576 36620
rect -11576 36586 -11508 36620
rect -11508 36586 -11418 36620
rect -11418 36586 -11350 36620
rect -11350 36586 -11260 36620
rect -11260 36586 -11192 36620
rect -11192 36586 -11102 36620
rect -11102 36586 -11034 36620
rect -11034 36586 -10944 36620
rect -10944 36586 -10876 36620
rect -10876 36586 -10786 36620
rect -10786 36586 -10718 36620
rect -10718 36586 -10628 36620
rect -10628 36586 -10560 36620
rect -10560 36586 -10470 36620
rect -10470 36586 -10402 36620
rect -10402 36586 -10312 36620
rect -10312 36586 -10244 36620
rect -10244 36586 -10154 36620
rect -10154 36586 -10086 36620
rect -10086 36586 -9996 36620
rect -9996 36586 -9928 36620
rect -9928 36586 -9838 36620
rect -9838 36586 -9770 36620
rect -9770 36586 -9680 36620
rect -9680 36586 -9612 36620
rect -9612 36586 -9522 36620
rect -9522 36586 -9454 36620
rect -9454 36586 -9364 36620
rect -9364 36586 -9296 36620
rect -9296 36586 -9206 36620
rect -9206 36586 -9138 36620
rect -9138 36586 -9048 36620
rect -9048 36586 -8980 36620
rect -8980 36586 -8890 36620
rect -8890 36586 -8822 36620
rect -8822 36586 -8732 36620
rect -8732 36586 -8664 36620
rect -8664 36586 -8574 36620
rect -8574 36586 -8514 36620
rect -13148 36526 -8514 36586
rect -8360 36500 -8290 36636
rect -7070 42680 -7000 42820
rect -6848 42730 -2214 42790
rect -6848 42696 -6788 42730
rect -6788 42696 -6698 42730
rect -6698 42696 -6630 42730
rect -6630 42696 -6540 42730
rect -6540 42696 -6472 42730
rect -6472 42696 -6382 42730
rect -6382 42696 -6314 42730
rect -6314 42696 -6224 42730
rect -6224 42696 -6156 42730
rect -6156 42696 -6066 42730
rect -6066 42696 -5998 42730
rect -5998 42696 -5908 42730
rect -5908 42696 -5840 42730
rect -5840 42696 -5750 42730
rect -5750 42696 -5682 42730
rect -5682 42696 -5592 42730
rect -5592 42696 -5524 42730
rect -5524 42696 -5434 42730
rect -5434 42696 -5366 42730
rect -5366 42696 -5276 42730
rect -5276 42696 -5208 42730
rect -5208 42696 -5118 42730
rect -5118 42696 -5050 42730
rect -5050 42696 -4960 42730
rect -4960 42696 -4892 42730
rect -4892 42696 -4802 42730
rect -4802 42696 -4734 42730
rect -4734 42696 -4644 42730
rect -4644 42696 -4576 42730
rect -4576 42696 -4486 42730
rect -4486 42696 -4418 42730
rect -4418 42696 -4328 42730
rect -4328 42696 -4260 42730
rect -4260 42696 -4170 42730
rect -4170 42696 -4102 42730
rect -4102 42696 -4012 42730
rect -4012 42696 -3944 42730
rect -3944 42696 -3854 42730
rect -3854 42696 -3786 42730
rect -3786 42696 -3696 42730
rect -3696 42696 -3628 42730
rect -3628 42696 -3538 42730
rect -3538 42696 -3470 42730
rect -3470 42696 -3380 42730
rect -3380 42696 -3312 42730
rect -3312 42696 -3222 42730
rect -3222 42696 -3154 42730
rect -3154 42696 -3064 42730
rect -3064 42696 -2996 42730
rect -2996 42696 -2906 42730
rect -2906 42696 -2838 42730
rect -2838 42696 -2748 42730
rect -2748 42696 -2680 42730
rect -2680 42696 -2590 42730
rect -2590 42696 -2522 42730
rect -2522 42696 -2432 42730
rect -2432 42696 -2364 42730
rect -2364 42696 -2274 42730
rect -2274 42696 -2214 42730
rect -6848 42690 -2214 42696
rect -7070 36636 -7054 42680
rect -7054 36636 -7016 42680
rect -7016 36636 -7000 42680
rect -2060 42680 -1990 42820
rect -6935 36678 -6918 42638
rect -6918 36678 -6884 42638
rect -6884 36678 -6869 42638
rect -6777 36678 -6760 42638
rect -6760 36678 -6726 42638
rect -6726 36678 -6711 42638
rect -6619 36678 -6602 42638
rect -6602 36678 -6568 42638
rect -6568 36678 -6553 42638
rect -6461 36678 -6444 42638
rect -6444 36678 -6410 42638
rect -6410 36678 -6395 42638
rect -6303 36678 -6286 42638
rect -6286 36678 -6252 42638
rect -6252 36678 -6237 42638
rect -6145 36678 -6128 42638
rect -6128 36678 -6094 42638
rect -6094 36678 -6079 42638
rect -5987 36678 -5970 42638
rect -5970 36678 -5936 42638
rect -5936 36678 -5921 42638
rect -5829 36678 -5812 42638
rect -5812 36678 -5778 42638
rect -5778 36678 -5763 42638
rect -5671 36678 -5654 42638
rect -5654 36678 -5620 42638
rect -5620 36678 -5605 42638
rect -5513 36678 -5496 42638
rect -5496 36678 -5462 42638
rect -5462 36678 -5447 42638
rect -5355 36678 -5338 42638
rect -5338 36678 -5304 42638
rect -5304 36678 -5289 42638
rect -5197 36678 -5180 42638
rect -5180 36678 -5146 42638
rect -5146 36678 -5131 42638
rect -5039 36678 -5022 42638
rect -5022 36678 -4988 42638
rect -4988 36678 -4973 42638
rect -4881 36678 -4864 42638
rect -4864 36678 -4830 42638
rect -4830 36678 -4815 42638
rect -4723 36678 -4706 42638
rect -4706 36678 -4672 42638
rect -4672 36678 -4657 42638
rect -4565 36678 -4548 42638
rect -4548 36678 -4514 42638
rect -4514 36678 -4499 42638
rect -4407 36678 -4390 42638
rect -4390 36678 -4356 42638
rect -4356 36678 -4341 42638
rect -4249 36678 -4232 42638
rect -4232 36678 -4198 42638
rect -4198 36678 -4183 42638
rect -4091 36678 -4074 42638
rect -4074 36678 -4040 42638
rect -4040 36678 -4025 42638
rect -3933 36678 -3916 42638
rect -3916 36678 -3882 42638
rect -3882 36678 -3867 42638
rect -3775 36678 -3758 42638
rect -3758 36678 -3724 42638
rect -3724 36678 -3709 42638
rect -3617 36678 -3600 42638
rect -3600 36678 -3566 42638
rect -3566 36678 -3551 42638
rect -3459 36678 -3442 42638
rect -3442 36678 -3408 42638
rect -3408 36678 -3393 42638
rect -3301 36678 -3284 42638
rect -3284 36678 -3250 42638
rect -3250 36678 -3235 42638
rect -3143 36678 -3126 42638
rect -3126 36678 -3092 42638
rect -3092 36678 -3077 42638
rect -2985 36678 -2968 42638
rect -2968 36678 -2934 42638
rect -2934 36678 -2919 42638
rect -2827 36678 -2810 42638
rect -2810 36678 -2776 42638
rect -2776 36678 -2761 42638
rect -2669 36678 -2652 42638
rect -2652 36678 -2618 42638
rect -2618 36678 -2603 42638
rect -2511 36678 -2494 42638
rect -2494 36678 -2460 42638
rect -2460 36678 -2445 42638
rect -2353 36678 -2336 42638
rect -2336 36678 -2302 42638
rect -2302 36678 -2287 42638
rect -2195 36678 -2178 42638
rect -2178 36678 -2144 42638
rect -2144 36678 -2129 42638
rect -7070 36500 -7000 36636
rect -2060 36636 -2046 42680
rect -2046 36636 -2008 42680
rect -2008 36636 -1990 42680
rect -6848 36620 -2214 36626
rect -6848 36586 -6788 36620
rect -6788 36586 -6698 36620
rect -6698 36586 -6630 36620
rect -6630 36586 -6540 36620
rect -6540 36586 -6472 36620
rect -6472 36586 -6382 36620
rect -6382 36586 -6314 36620
rect -6314 36586 -6224 36620
rect -6224 36586 -6156 36620
rect -6156 36586 -6066 36620
rect -6066 36586 -5998 36620
rect -5998 36586 -5908 36620
rect -5908 36586 -5840 36620
rect -5840 36586 -5750 36620
rect -5750 36586 -5682 36620
rect -5682 36586 -5592 36620
rect -5592 36586 -5524 36620
rect -5524 36586 -5434 36620
rect -5434 36586 -5366 36620
rect -5366 36586 -5276 36620
rect -5276 36586 -5208 36620
rect -5208 36586 -5118 36620
rect -5118 36586 -5050 36620
rect -5050 36586 -4960 36620
rect -4960 36586 -4892 36620
rect -4892 36586 -4802 36620
rect -4802 36586 -4734 36620
rect -4734 36586 -4644 36620
rect -4644 36586 -4576 36620
rect -4576 36586 -4486 36620
rect -4486 36586 -4418 36620
rect -4418 36586 -4328 36620
rect -4328 36586 -4260 36620
rect -4260 36586 -4170 36620
rect -4170 36586 -4102 36620
rect -4102 36586 -4012 36620
rect -4012 36586 -3944 36620
rect -3944 36586 -3854 36620
rect -3854 36586 -3786 36620
rect -3786 36586 -3696 36620
rect -3696 36586 -3628 36620
rect -3628 36586 -3538 36620
rect -3538 36586 -3470 36620
rect -3470 36586 -3380 36620
rect -3380 36586 -3312 36620
rect -3312 36586 -3222 36620
rect -3222 36586 -3154 36620
rect -3154 36586 -3064 36620
rect -3064 36586 -2996 36620
rect -2996 36586 -2906 36620
rect -2906 36586 -2838 36620
rect -2838 36586 -2748 36620
rect -2748 36586 -2680 36620
rect -2680 36586 -2590 36620
rect -2590 36586 -2522 36620
rect -2522 36586 -2432 36620
rect -2432 36586 -2364 36620
rect -2364 36586 -2274 36620
rect -2274 36586 -2214 36620
rect -6848 36526 -2214 36586
rect -2060 36500 -1990 36636
rect -770 42680 -700 42820
rect -548 42730 4086 42790
rect -548 42696 -488 42730
rect -488 42696 -398 42730
rect -398 42696 -330 42730
rect -330 42696 -240 42730
rect -240 42696 -172 42730
rect -172 42696 -82 42730
rect -82 42696 -14 42730
rect -14 42696 76 42730
rect 76 42696 144 42730
rect 144 42696 234 42730
rect 234 42696 302 42730
rect 302 42696 392 42730
rect 392 42696 460 42730
rect 460 42696 550 42730
rect 550 42696 618 42730
rect 618 42696 708 42730
rect 708 42696 776 42730
rect 776 42696 866 42730
rect 866 42696 934 42730
rect 934 42696 1024 42730
rect 1024 42696 1092 42730
rect 1092 42696 1182 42730
rect 1182 42696 1250 42730
rect 1250 42696 1340 42730
rect 1340 42696 1408 42730
rect 1408 42696 1498 42730
rect 1498 42696 1566 42730
rect 1566 42696 1656 42730
rect 1656 42696 1724 42730
rect 1724 42696 1814 42730
rect 1814 42696 1882 42730
rect 1882 42696 1972 42730
rect 1972 42696 2040 42730
rect 2040 42696 2130 42730
rect 2130 42696 2198 42730
rect 2198 42696 2288 42730
rect 2288 42696 2356 42730
rect 2356 42696 2446 42730
rect 2446 42696 2514 42730
rect 2514 42696 2604 42730
rect 2604 42696 2672 42730
rect 2672 42696 2762 42730
rect 2762 42696 2830 42730
rect 2830 42696 2920 42730
rect 2920 42696 2988 42730
rect 2988 42696 3078 42730
rect 3078 42696 3146 42730
rect 3146 42696 3236 42730
rect 3236 42696 3304 42730
rect 3304 42696 3394 42730
rect 3394 42696 3462 42730
rect 3462 42696 3552 42730
rect 3552 42696 3620 42730
rect 3620 42696 3710 42730
rect 3710 42696 3778 42730
rect 3778 42696 3868 42730
rect 3868 42696 3936 42730
rect 3936 42696 4026 42730
rect 4026 42696 4086 42730
rect -548 42690 4086 42696
rect -770 36636 -754 42680
rect -754 36636 -716 42680
rect -716 36636 -700 42680
rect 4240 42680 4310 42820
rect -635 36678 -618 42638
rect -618 36678 -584 42638
rect -584 36678 -569 42638
rect -477 36678 -460 42638
rect -460 36678 -426 42638
rect -426 36678 -411 42638
rect -319 36678 -302 42638
rect -302 36678 -268 42638
rect -268 36678 -253 42638
rect -161 36678 -144 42638
rect -144 36678 -110 42638
rect -110 36678 -95 42638
rect -3 36678 14 42638
rect 14 36678 48 42638
rect 48 36678 63 42638
rect 155 36678 172 42638
rect 172 36678 206 42638
rect 206 36678 221 42638
rect 313 36678 330 42638
rect 330 36678 364 42638
rect 364 36678 379 42638
rect 471 36678 488 42638
rect 488 36678 522 42638
rect 522 36678 537 42638
rect 629 36678 646 42638
rect 646 36678 680 42638
rect 680 36678 695 42638
rect 787 36678 804 42638
rect 804 36678 838 42638
rect 838 36678 853 42638
rect 945 36678 962 42638
rect 962 36678 996 42638
rect 996 36678 1011 42638
rect 1103 36678 1120 42638
rect 1120 36678 1154 42638
rect 1154 36678 1169 42638
rect 1261 36678 1278 42638
rect 1278 36678 1312 42638
rect 1312 36678 1327 42638
rect 1419 36678 1436 42638
rect 1436 36678 1470 42638
rect 1470 36678 1485 42638
rect 1577 36678 1594 42638
rect 1594 36678 1628 42638
rect 1628 36678 1643 42638
rect 1735 36678 1752 42638
rect 1752 36678 1786 42638
rect 1786 36678 1801 42638
rect 1893 36678 1910 42638
rect 1910 36678 1944 42638
rect 1944 36678 1959 42638
rect 2051 36678 2068 42638
rect 2068 36678 2102 42638
rect 2102 36678 2117 42638
rect 2209 36678 2226 42638
rect 2226 36678 2260 42638
rect 2260 36678 2275 42638
rect 2367 36678 2384 42638
rect 2384 36678 2418 42638
rect 2418 36678 2433 42638
rect 2525 36678 2542 42638
rect 2542 36678 2576 42638
rect 2576 36678 2591 42638
rect 2683 36678 2700 42638
rect 2700 36678 2734 42638
rect 2734 36678 2749 42638
rect 2841 36678 2858 42638
rect 2858 36678 2892 42638
rect 2892 36678 2907 42638
rect 2999 36678 3016 42638
rect 3016 36678 3050 42638
rect 3050 36678 3065 42638
rect 3157 36678 3174 42638
rect 3174 36678 3208 42638
rect 3208 36678 3223 42638
rect 3315 36678 3332 42638
rect 3332 36678 3366 42638
rect 3366 36678 3381 42638
rect 3473 36678 3490 42638
rect 3490 36678 3524 42638
rect 3524 36678 3539 42638
rect 3631 36678 3648 42638
rect 3648 36678 3682 42638
rect 3682 36678 3697 42638
rect 3789 36678 3806 42638
rect 3806 36678 3840 42638
rect 3840 36678 3855 42638
rect 3947 36678 3964 42638
rect 3964 36678 3998 42638
rect 3998 36678 4013 42638
rect 4105 36678 4122 42638
rect 4122 36678 4156 42638
rect 4156 36678 4171 42638
rect -770 36500 -700 36636
rect 4240 36636 4254 42680
rect 4254 36636 4292 42680
rect 4292 36636 4310 42680
rect -548 36620 4086 36626
rect -548 36586 -488 36620
rect -488 36586 -398 36620
rect -398 36586 -330 36620
rect -330 36586 -240 36620
rect -240 36586 -172 36620
rect -172 36586 -82 36620
rect -82 36586 -14 36620
rect -14 36586 76 36620
rect 76 36586 144 36620
rect 144 36586 234 36620
rect 234 36586 302 36620
rect 302 36586 392 36620
rect 392 36586 460 36620
rect 460 36586 550 36620
rect 550 36586 618 36620
rect 618 36586 708 36620
rect 708 36586 776 36620
rect 776 36586 866 36620
rect 866 36586 934 36620
rect 934 36586 1024 36620
rect 1024 36586 1092 36620
rect 1092 36586 1182 36620
rect 1182 36586 1250 36620
rect 1250 36586 1340 36620
rect 1340 36586 1408 36620
rect 1408 36586 1498 36620
rect 1498 36586 1566 36620
rect 1566 36586 1656 36620
rect 1656 36586 1724 36620
rect 1724 36586 1814 36620
rect 1814 36586 1882 36620
rect 1882 36586 1972 36620
rect 1972 36586 2040 36620
rect 2040 36586 2130 36620
rect 2130 36586 2198 36620
rect 2198 36586 2288 36620
rect 2288 36586 2356 36620
rect 2356 36586 2446 36620
rect 2446 36586 2514 36620
rect 2514 36586 2604 36620
rect 2604 36586 2672 36620
rect 2672 36586 2762 36620
rect 2762 36586 2830 36620
rect 2830 36586 2920 36620
rect 2920 36586 2988 36620
rect 2988 36586 3078 36620
rect 3078 36586 3146 36620
rect 3146 36586 3236 36620
rect 3236 36586 3304 36620
rect 3304 36586 3394 36620
rect 3394 36586 3462 36620
rect 3462 36586 3552 36620
rect 3552 36586 3620 36620
rect 3620 36586 3710 36620
rect 3710 36586 3778 36620
rect 3778 36586 3868 36620
rect 3868 36586 3936 36620
rect 3936 36586 4026 36620
rect 4026 36586 4086 36620
rect -548 36526 4086 36586
rect 4240 36500 4310 36636
rect 5530 42680 5600 42820
rect 5752 42730 10386 42790
rect 5752 42696 5812 42730
rect 5812 42696 5902 42730
rect 5902 42696 5970 42730
rect 5970 42696 6060 42730
rect 6060 42696 6128 42730
rect 6128 42696 6218 42730
rect 6218 42696 6286 42730
rect 6286 42696 6376 42730
rect 6376 42696 6444 42730
rect 6444 42696 6534 42730
rect 6534 42696 6602 42730
rect 6602 42696 6692 42730
rect 6692 42696 6760 42730
rect 6760 42696 6850 42730
rect 6850 42696 6918 42730
rect 6918 42696 7008 42730
rect 7008 42696 7076 42730
rect 7076 42696 7166 42730
rect 7166 42696 7234 42730
rect 7234 42696 7324 42730
rect 7324 42696 7392 42730
rect 7392 42696 7482 42730
rect 7482 42696 7550 42730
rect 7550 42696 7640 42730
rect 7640 42696 7708 42730
rect 7708 42696 7798 42730
rect 7798 42696 7866 42730
rect 7866 42696 7956 42730
rect 7956 42696 8024 42730
rect 8024 42696 8114 42730
rect 8114 42696 8182 42730
rect 8182 42696 8272 42730
rect 8272 42696 8340 42730
rect 8340 42696 8430 42730
rect 8430 42696 8498 42730
rect 8498 42696 8588 42730
rect 8588 42696 8656 42730
rect 8656 42696 8746 42730
rect 8746 42696 8814 42730
rect 8814 42696 8904 42730
rect 8904 42696 8972 42730
rect 8972 42696 9062 42730
rect 9062 42696 9130 42730
rect 9130 42696 9220 42730
rect 9220 42696 9288 42730
rect 9288 42696 9378 42730
rect 9378 42696 9446 42730
rect 9446 42696 9536 42730
rect 9536 42696 9604 42730
rect 9604 42696 9694 42730
rect 9694 42696 9762 42730
rect 9762 42696 9852 42730
rect 9852 42696 9920 42730
rect 9920 42696 10010 42730
rect 10010 42696 10078 42730
rect 10078 42696 10168 42730
rect 10168 42696 10236 42730
rect 10236 42696 10326 42730
rect 10326 42696 10386 42730
rect 5752 42690 10386 42696
rect 5530 36636 5546 42680
rect 5546 36636 5584 42680
rect 5584 36636 5600 42680
rect 10540 42680 10610 42820
rect 5665 36678 5682 42638
rect 5682 36678 5716 42638
rect 5716 36678 5731 42638
rect 5823 36678 5840 42638
rect 5840 36678 5874 42638
rect 5874 36678 5889 42638
rect 5981 36678 5998 42638
rect 5998 36678 6032 42638
rect 6032 36678 6047 42638
rect 6139 36678 6156 42638
rect 6156 36678 6190 42638
rect 6190 36678 6205 42638
rect 6297 36678 6314 42638
rect 6314 36678 6348 42638
rect 6348 36678 6363 42638
rect 6455 36678 6472 42638
rect 6472 36678 6506 42638
rect 6506 36678 6521 42638
rect 6613 36678 6630 42638
rect 6630 36678 6664 42638
rect 6664 36678 6679 42638
rect 6771 36678 6788 42638
rect 6788 36678 6822 42638
rect 6822 36678 6837 42638
rect 6929 36678 6946 42638
rect 6946 36678 6980 42638
rect 6980 36678 6995 42638
rect 7087 36678 7104 42638
rect 7104 36678 7138 42638
rect 7138 36678 7153 42638
rect 7245 36678 7262 42638
rect 7262 36678 7296 42638
rect 7296 36678 7311 42638
rect 7403 36678 7420 42638
rect 7420 36678 7454 42638
rect 7454 36678 7469 42638
rect 7561 36678 7578 42638
rect 7578 36678 7612 42638
rect 7612 36678 7627 42638
rect 7719 36678 7736 42638
rect 7736 36678 7770 42638
rect 7770 36678 7785 42638
rect 7877 36678 7894 42638
rect 7894 36678 7928 42638
rect 7928 36678 7943 42638
rect 8035 36678 8052 42638
rect 8052 36678 8086 42638
rect 8086 36678 8101 42638
rect 8193 36678 8210 42638
rect 8210 36678 8244 42638
rect 8244 36678 8259 42638
rect 8351 36678 8368 42638
rect 8368 36678 8402 42638
rect 8402 36678 8417 42638
rect 8509 36678 8526 42638
rect 8526 36678 8560 42638
rect 8560 36678 8575 42638
rect 8667 36678 8684 42638
rect 8684 36678 8718 42638
rect 8718 36678 8733 42638
rect 8825 36678 8842 42638
rect 8842 36678 8876 42638
rect 8876 36678 8891 42638
rect 8983 36678 9000 42638
rect 9000 36678 9034 42638
rect 9034 36678 9049 42638
rect 9141 36678 9158 42638
rect 9158 36678 9192 42638
rect 9192 36678 9207 42638
rect 9299 36678 9316 42638
rect 9316 36678 9350 42638
rect 9350 36678 9365 42638
rect 9457 36678 9474 42638
rect 9474 36678 9508 42638
rect 9508 36678 9523 42638
rect 9615 36678 9632 42638
rect 9632 36678 9666 42638
rect 9666 36678 9681 42638
rect 9773 36678 9790 42638
rect 9790 36678 9824 42638
rect 9824 36678 9839 42638
rect 9931 36678 9948 42638
rect 9948 36678 9982 42638
rect 9982 36678 9997 42638
rect 10089 36678 10106 42638
rect 10106 36678 10140 42638
rect 10140 36678 10155 42638
rect 10247 36678 10264 42638
rect 10264 36678 10298 42638
rect 10298 36678 10313 42638
rect 10405 36678 10422 42638
rect 10422 36678 10456 42638
rect 10456 36678 10471 42638
rect 5530 36500 5600 36636
rect 10540 36636 10554 42680
rect 10554 36636 10592 42680
rect 10592 36636 10610 42680
rect 5752 36620 10386 36626
rect 5752 36586 5812 36620
rect 5812 36586 5902 36620
rect 5902 36586 5970 36620
rect 5970 36586 6060 36620
rect 6060 36586 6128 36620
rect 6128 36586 6218 36620
rect 6218 36586 6286 36620
rect 6286 36586 6376 36620
rect 6376 36586 6444 36620
rect 6444 36586 6534 36620
rect 6534 36586 6602 36620
rect 6602 36586 6692 36620
rect 6692 36586 6760 36620
rect 6760 36586 6850 36620
rect 6850 36586 6918 36620
rect 6918 36586 7008 36620
rect 7008 36586 7076 36620
rect 7076 36586 7166 36620
rect 7166 36586 7234 36620
rect 7234 36586 7324 36620
rect 7324 36586 7392 36620
rect 7392 36586 7482 36620
rect 7482 36586 7550 36620
rect 7550 36586 7640 36620
rect 7640 36586 7708 36620
rect 7708 36586 7798 36620
rect 7798 36586 7866 36620
rect 7866 36586 7956 36620
rect 7956 36586 8024 36620
rect 8024 36586 8114 36620
rect 8114 36586 8182 36620
rect 8182 36586 8272 36620
rect 8272 36586 8340 36620
rect 8340 36586 8430 36620
rect 8430 36586 8498 36620
rect 8498 36586 8588 36620
rect 8588 36586 8656 36620
rect 8656 36586 8746 36620
rect 8746 36586 8814 36620
rect 8814 36586 8904 36620
rect 8904 36586 8972 36620
rect 8972 36586 9062 36620
rect 9062 36586 9130 36620
rect 9130 36586 9220 36620
rect 9220 36586 9288 36620
rect 9288 36586 9378 36620
rect 9378 36586 9446 36620
rect 9446 36586 9536 36620
rect 9536 36586 9604 36620
rect 9604 36586 9694 36620
rect 9694 36586 9762 36620
rect 9762 36586 9852 36620
rect 9852 36586 9920 36620
rect 9920 36586 10010 36620
rect 10010 36586 10078 36620
rect 10078 36586 10168 36620
rect 10168 36586 10236 36620
rect 10236 36586 10326 36620
rect 10326 36586 10386 36620
rect 5752 36526 10386 36586
rect 10540 36500 10610 36636
rect -13370 34380 -13300 34520
rect -13148 34430 -8514 34490
rect -13148 34396 -13088 34430
rect -13088 34396 -12998 34430
rect -12998 34396 -12930 34430
rect -12930 34396 -12840 34430
rect -12840 34396 -12772 34430
rect -12772 34396 -12682 34430
rect -12682 34396 -12614 34430
rect -12614 34396 -12524 34430
rect -12524 34396 -12456 34430
rect -12456 34396 -12366 34430
rect -12366 34396 -12298 34430
rect -12298 34396 -12208 34430
rect -12208 34396 -12140 34430
rect -12140 34396 -12050 34430
rect -12050 34396 -11982 34430
rect -11982 34396 -11892 34430
rect -11892 34396 -11824 34430
rect -11824 34396 -11734 34430
rect -11734 34396 -11666 34430
rect -11666 34396 -11576 34430
rect -11576 34396 -11508 34430
rect -11508 34396 -11418 34430
rect -11418 34396 -11350 34430
rect -11350 34396 -11260 34430
rect -11260 34396 -11192 34430
rect -11192 34396 -11102 34430
rect -11102 34396 -11034 34430
rect -11034 34396 -10944 34430
rect -10944 34396 -10876 34430
rect -10876 34396 -10786 34430
rect -10786 34396 -10718 34430
rect -10718 34396 -10628 34430
rect -10628 34396 -10560 34430
rect -10560 34396 -10470 34430
rect -10470 34396 -10402 34430
rect -10402 34396 -10312 34430
rect -10312 34396 -10244 34430
rect -10244 34396 -10154 34430
rect -10154 34396 -10086 34430
rect -10086 34396 -9996 34430
rect -9996 34396 -9928 34430
rect -9928 34396 -9838 34430
rect -9838 34396 -9770 34430
rect -9770 34396 -9680 34430
rect -9680 34396 -9612 34430
rect -9612 34396 -9522 34430
rect -9522 34396 -9454 34430
rect -9454 34396 -9364 34430
rect -9364 34396 -9296 34430
rect -9296 34396 -9206 34430
rect -9206 34396 -9138 34430
rect -9138 34396 -9048 34430
rect -9048 34396 -8980 34430
rect -8980 34396 -8890 34430
rect -8890 34396 -8822 34430
rect -8822 34396 -8732 34430
rect -8732 34396 -8664 34430
rect -8664 34396 -8574 34430
rect -8574 34396 -8514 34430
rect -13148 34390 -8514 34396
rect -13370 28336 -13354 34380
rect -13354 28336 -13316 34380
rect -13316 28336 -13300 34380
rect -8360 34380 -8290 34520
rect -13235 28378 -13218 34338
rect -13218 28378 -13184 34338
rect -13184 28378 -13169 34338
rect -13077 28378 -13060 34338
rect -13060 28378 -13026 34338
rect -13026 28378 -13011 34338
rect -12919 28378 -12902 34338
rect -12902 28378 -12868 34338
rect -12868 28378 -12853 34338
rect -12761 28378 -12744 34338
rect -12744 28378 -12710 34338
rect -12710 28378 -12695 34338
rect -12603 28378 -12586 34338
rect -12586 28378 -12552 34338
rect -12552 28378 -12537 34338
rect -12445 28378 -12428 34338
rect -12428 28378 -12394 34338
rect -12394 28378 -12379 34338
rect -12287 28378 -12270 34338
rect -12270 28378 -12236 34338
rect -12236 28378 -12221 34338
rect -12129 28378 -12112 34338
rect -12112 28378 -12078 34338
rect -12078 28378 -12063 34338
rect -11971 28378 -11954 34338
rect -11954 28378 -11920 34338
rect -11920 28378 -11905 34338
rect -11813 28378 -11796 34338
rect -11796 28378 -11762 34338
rect -11762 28378 -11747 34338
rect -11655 28378 -11638 34338
rect -11638 28378 -11604 34338
rect -11604 28378 -11589 34338
rect -11497 28378 -11480 34338
rect -11480 28378 -11446 34338
rect -11446 28378 -11431 34338
rect -11339 28378 -11322 34338
rect -11322 28378 -11288 34338
rect -11288 28378 -11273 34338
rect -11181 28378 -11164 34338
rect -11164 28378 -11130 34338
rect -11130 28378 -11115 34338
rect -11023 28378 -11006 34338
rect -11006 28378 -10972 34338
rect -10972 28378 -10957 34338
rect -10865 28378 -10848 34338
rect -10848 28378 -10814 34338
rect -10814 28378 -10799 34338
rect -10707 28378 -10690 34338
rect -10690 28378 -10656 34338
rect -10656 28378 -10641 34338
rect -10549 28378 -10532 34338
rect -10532 28378 -10498 34338
rect -10498 28378 -10483 34338
rect -10391 28378 -10374 34338
rect -10374 28378 -10340 34338
rect -10340 28378 -10325 34338
rect -10233 28378 -10216 34338
rect -10216 28378 -10182 34338
rect -10182 28378 -10167 34338
rect -10075 28378 -10058 34338
rect -10058 28378 -10024 34338
rect -10024 28378 -10009 34338
rect -9917 28378 -9900 34338
rect -9900 28378 -9866 34338
rect -9866 28378 -9851 34338
rect -9759 28378 -9742 34338
rect -9742 28378 -9708 34338
rect -9708 28378 -9693 34338
rect -9601 28378 -9584 34338
rect -9584 28378 -9550 34338
rect -9550 28378 -9535 34338
rect -9443 28378 -9426 34338
rect -9426 28378 -9392 34338
rect -9392 28378 -9377 34338
rect -9285 28378 -9268 34338
rect -9268 28378 -9234 34338
rect -9234 28378 -9219 34338
rect -9127 28378 -9110 34338
rect -9110 28378 -9076 34338
rect -9076 28378 -9061 34338
rect -8969 28378 -8952 34338
rect -8952 28378 -8918 34338
rect -8918 28378 -8903 34338
rect -8811 28378 -8794 34338
rect -8794 28378 -8760 34338
rect -8760 28378 -8745 34338
rect -8653 28378 -8636 34338
rect -8636 28378 -8602 34338
rect -8602 28378 -8587 34338
rect -8495 28378 -8478 34338
rect -8478 28378 -8444 34338
rect -8444 28378 -8429 34338
rect -13370 28200 -13300 28336
rect -8360 28336 -8346 34380
rect -8346 28336 -8308 34380
rect -8308 28336 -8290 34380
rect -13148 28320 -8514 28326
rect -13148 28286 -13088 28320
rect -13088 28286 -12998 28320
rect -12998 28286 -12930 28320
rect -12930 28286 -12840 28320
rect -12840 28286 -12772 28320
rect -12772 28286 -12682 28320
rect -12682 28286 -12614 28320
rect -12614 28286 -12524 28320
rect -12524 28286 -12456 28320
rect -12456 28286 -12366 28320
rect -12366 28286 -12298 28320
rect -12298 28286 -12208 28320
rect -12208 28286 -12140 28320
rect -12140 28286 -12050 28320
rect -12050 28286 -11982 28320
rect -11982 28286 -11892 28320
rect -11892 28286 -11824 28320
rect -11824 28286 -11734 28320
rect -11734 28286 -11666 28320
rect -11666 28286 -11576 28320
rect -11576 28286 -11508 28320
rect -11508 28286 -11418 28320
rect -11418 28286 -11350 28320
rect -11350 28286 -11260 28320
rect -11260 28286 -11192 28320
rect -11192 28286 -11102 28320
rect -11102 28286 -11034 28320
rect -11034 28286 -10944 28320
rect -10944 28286 -10876 28320
rect -10876 28286 -10786 28320
rect -10786 28286 -10718 28320
rect -10718 28286 -10628 28320
rect -10628 28286 -10560 28320
rect -10560 28286 -10470 28320
rect -10470 28286 -10402 28320
rect -10402 28286 -10312 28320
rect -10312 28286 -10244 28320
rect -10244 28286 -10154 28320
rect -10154 28286 -10086 28320
rect -10086 28286 -9996 28320
rect -9996 28286 -9928 28320
rect -9928 28286 -9838 28320
rect -9838 28286 -9770 28320
rect -9770 28286 -9680 28320
rect -9680 28286 -9612 28320
rect -9612 28286 -9522 28320
rect -9522 28286 -9454 28320
rect -9454 28286 -9364 28320
rect -9364 28286 -9296 28320
rect -9296 28286 -9206 28320
rect -9206 28286 -9138 28320
rect -9138 28286 -9048 28320
rect -9048 28286 -8980 28320
rect -8980 28286 -8890 28320
rect -8890 28286 -8822 28320
rect -8822 28286 -8732 28320
rect -8732 28286 -8664 28320
rect -8664 28286 -8574 28320
rect -8574 28286 -8514 28320
rect -13148 28226 -8514 28286
rect -8360 28200 -8290 28336
rect -7070 34380 -7000 34520
rect -6848 34430 -2214 34490
rect -6848 34396 -6788 34430
rect -6788 34396 -6698 34430
rect -6698 34396 -6630 34430
rect -6630 34396 -6540 34430
rect -6540 34396 -6472 34430
rect -6472 34396 -6382 34430
rect -6382 34396 -6314 34430
rect -6314 34396 -6224 34430
rect -6224 34396 -6156 34430
rect -6156 34396 -6066 34430
rect -6066 34396 -5998 34430
rect -5998 34396 -5908 34430
rect -5908 34396 -5840 34430
rect -5840 34396 -5750 34430
rect -5750 34396 -5682 34430
rect -5682 34396 -5592 34430
rect -5592 34396 -5524 34430
rect -5524 34396 -5434 34430
rect -5434 34396 -5366 34430
rect -5366 34396 -5276 34430
rect -5276 34396 -5208 34430
rect -5208 34396 -5118 34430
rect -5118 34396 -5050 34430
rect -5050 34396 -4960 34430
rect -4960 34396 -4892 34430
rect -4892 34396 -4802 34430
rect -4802 34396 -4734 34430
rect -4734 34396 -4644 34430
rect -4644 34396 -4576 34430
rect -4576 34396 -4486 34430
rect -4486 34396 -4418 34430
rect -4418 34396 -4328 34430
rect -4328 34396 -4260 34430
rect -4260 34396 -4170 34430
rect -4170 34396 -4102 34430
rect -4102 34396 -4012 34430
rect -4012 34396 -3944 34430
rect -3944 34396 -3854 34430
rect -3854 34396 -3786 34430
rect -3786 34396 -3696 34430
rect -3696 34396 -3628 34430
rect -3628 34396 -3538 34430
rect -3538 34396 -3470 34430
rect -3470 34396 -3380 34430
rect -3380 34396 -3312 34430
rect -3312 34396 -3222 34430
rect -3222 34396 -3154 34430
rect -3154 34396 -3064 34430
rect -3064 34396 -2996 34430
rect -2996 34396 -2906 34430
rect -2906 34396 -2838 34430
rect -2838 34396 -2748 34430
rect -2748 34396 -2680 34430
rect -2680 34396 -2590 34430
rect -2590 34396 -2522 34430
rect -2522 34396 -2432 34430
rect -2432 34396 -2364 34430
rect -2364 34396 -2274 34430
rect -2274 34396 -2214 34430
rect -6848 34390 -2214 34396
rect -7070 28336 -7054 34380
rect -7054 28336 -7016 34380
rect -7016 28336 -7000 34380
rect -2060 34380 -1990 34520
rect -6935 28378 -6918 34338
rect -6918 28378 -6884 34338
rect -6884 28378 -6869 34338
rect -6777 28378 -6760 34338
rect -6760 28378 -6726 34338
rect -6726 28378 -6711 34338
rect -6619 28378 -6602 34338
rect -6602 28378 -6568 34338
rect -6568 28378 -6553 34338
rect -6461 28378 -6444 34338
rect -6444 28378 -6410 34338
rect -6410 28378 -6395 34338
rect -6303 28378 -6286 34338
rect -6286 28378 -6252 34338
rect -6252 28378 -6237 34338
rect -6145 28378 -6128 34338
rect -6128 28378 -6094 34338
rect -6094 28378 -6079 34338
rect -5987 28378 -5970 34338
rect -5970 28378 -5936 34338
rect -5936 28378 -5921 34338
rect -5829 28378 -5812 34338
rect -5812 28378 -5778 34338
rect -5778 28378 -5763 34338
rect -5671 28378 -5654 34338
rect -5654 28378 -5620 34338
rect -5620 28378 -5605 34338
rect -5513 28378 -5496 34338
rect -5496 28378 -5462 34338
rect -5462 28378 -5447 34338
rect -5355 28378 -5338 34338
rect -5338 28378 -5304 34338
rect -5304 28378 -5289 34338
rect -5197 28378 -5180 34338
rect -5180 28378 -5146 34338
rect -5146 28378 -5131 34338
rect -5039 28378 -5022 34338
rect -5022 28378 -4988 34338
rect -4988 28378 -4973 34338
rect -4881 28378 -4864 34338
rect -4864 28378 -4830 34338
rect -4830 28378 -4815 34338
rect -4723 28378 -4706 34338
rect -4706 28378 -4672 34338
rect -4672 28378 -4657 34338
rect -4565 28378 -4548 34338
rect -4548 28378 -4514 34338
rect -4514 28378 -4499 34338
rect -4407 28378 -4390 34338
rect -4390 28378 -4356 34338
rect -4356 28378 -4341 34338
rect -4249 28378 -4232 34338
rect -4232 28378 -4198 34338
rect -4198 28378 -4183 34338
rect -4091 28378 -4074 34338
rect -4074 28378 -4040 34338
rect -4040 28378 -4025 34338
rect -3933 28378 -3916 34338
rect -3916 28378 -3882 34338
rect -3882 28378 -3867 34338
rect -3775 28378 -3758 34338
rect -3758 28378 -3724 34338
rect -3724 28378 -3709 34338
rect -3617 28378 -3600 34338
rect -3600 28378 -3566 34338
rect -3566 28378 -3551 34338
rect -3459 28378 -3442 34338
rect -3442 28378 -3408 34338
rect -3408 28378 -3393 34338
rect -3301 28378 -3284 34338
rect -3284 28378 -3250 34338
rect -3250 28378 -3235 34338
rect -3143 28378 -3126 34338
rect -3126 28378 -3092 34338
rect -3092 28378 -3077 34338
rect -2985 28378 -2968 34338
rect -2968 28378 -2934 34338
rect -2934 28378 -2919 34338
rect -2827 28378 -2810 34338
rect -2810 28378 -2776 34338
rect -2776 28378 -2761 34338
rect -2669 28378 -2652 34338
rect -2652 28378 -2618 34338
rect -2618 28378 -2603 34338
rect -2511 28378 -2494 34338
rect -2494 28378 -2460 34338
rect -2460 28378 -2445 34338
rect -2353 28378 -2336 34338
rect -2336 28378 -2302 34338
rect -2302 28378 -2287 34338
rect -2195 28378 -2178 34338
rect -2178 28378 -2144 34338
rect -2144 28378 -2129 34338
rect -7070 28200 -7000 28336
rect -2060 28336 -2046 34380
rect -2046 28336 -2008 34380
rect -2008 28336 -1990 34380
rect -6848 28320 -2214 28326
rect -6848 28286 -6788 28320
rect -6788 28286 -6698 28320
rect -6698 28286 -6630 28320
rect -6630 28286 -6540 28320
rect -6540 28286 -6472 28320
rect -6472 28286 -6382 28320
rect -6382 28286 -6314 28320
rect -6314 28286 -6224 28320
rect -6224 28286 -6156 28320
rect -6156 28286 -6066 28320
rect -6066 28286 -5998 28320
rect -5998 28286 -5908 28320
rect -5908 28286 -5840 28320
rect -5840 28286 -5750 28320
rect -5750 28286 -5682 28320
rect -5682 28286 -5592 28320
rect -5592 28286 -5524 28320
rect -5524 28286 -5434 28320
rect -5434 28286 -5366 28320
rect -5366 28286 -5276 28320
rect -5276 28286 -5208 28320
rect -5208 28286 -5118 28320
rect -5118 28286 -5050 28320
rect -5050 28286 -4960 28320
rect -4960 28286 -4892 28320
rect -4892 28286 -4802 28320
rect -4802 28286 -4734 28320
rect -4734 28286 -4644 28320
rect -4644 28286 -4576 28320
rect -4576 28286 -4486 28320
rect -4486 28286 -4418 28320
rect -4418 28286 -4328 28320
rect -4328 28286 -4260 28320
rect -4260 28286 -4170 28320
rect -4170 28286 -4102 28320
rect -4102 28286 -4012 28320
rect -4012 28286 -3944 28320
rect -3944 28286 -3854 28320
rect -3854 28286 -3786 28320
rect -3786 28286 -3696 28320
rect -3696 28286 -3628 28320
rect -3628 28286 -3538 28320
rect -3538 28286 -3470 28320
rect -3470 28286 -3380 28320
rect -3380 28286 -3312 28320
rect -3312 28286 -3222 28320
rect -3222 28286 -3154 28320
rect -3154 28286 -3064 28320
rect -3064 28286 -2996 28320
rect -2996 28286 -2906 28320
rect -2906 28286 -2838 28320
rect -2838 28286 -2748 28320
rect -2748 28286 -2680 28320
rect -2680 28286 -2590 28320
rect -2590 28286 -2522 28320
rect -2522 28286 -2432 28320
rect -2432 28286 -2364 28320
rect -2364 28286 -2274 28320
rect -2274 28286 -2214 28320
rect -6848 28226 -2214 28286
rect -2060 28200 -1990 28336
rect -770 34380 -700 34520
rect -548 34430 4086 34490
rect -548 34396 -488 34430
rect -488 34396 -398 34430
rect -398 34396 -330 34430
rect -330 34396 -240 34430
rect -240 34396 -172 34430
rect -172 34396 -82 34430
rect -82 34396 -14 34430
rect -14 34396 76 34430
rect 76 34396 144 34430
rect 144 34396 234 34430
rect 234 34396 302 34430
rect 302 34396 392 34430
rect 392 34396 460 34430
rect 460 34396 550 34430
rect 550 34396 618 34430
rect 618 34396 708 34430
rect 708 34396 776 34430
rect 776 34396 866 34430
rect 866 34396 934 34430
rect 934 34396 1024 34430
rect 1024 34396 1092 34430
rect 1092 34396 1182 34430
rect 1182 34396 1250 34430
rect 1250 34396 1340 34430
rect 1340 34396 1408 34430
rect 1408 34396 1498 34430
rect 1498 34396 1566 34430
rect 1566 34396 1656 34430
rect 1656 34396 1724 34430
rect 1724 34396 1814 34430
rect 1814 34396 1882 34430
rect 1882 34396 1972 34430
rect 1972 34396 2040 34430
rect 2040 34396 2130 34430
rect 2130 34396 2198 34430
rect 2198 34396 2288 34430
rect 2288 34396 2356 34430
rect 2356 34396 2446 34430
rect 2446 34396 2514 34430
rect 2514 34396 2604 34430
rect 2604 34396 2672 34430
rect 2672 34396 2762 34430
rect 2762 34396 2830 34430
rect 2830 34396 2920 34430
rect 2920 34396 2988 34430
rect 2988 34396 3078 34430
rect 3078 34396 3146 34430
rect 3146 34396 3236 34430
rect 3236 34396 3304 34430
rect 3304 34396 3394 34430
rect 3394 34396 3462 34430
rect 3462 34396 3552 34430
rect 3552 34396 3620 34430
rect 3620 34396 3710 34430
rect 3710 34396 3778 34430
rect 3778 34396 3868 34430
rect 3868 34396 3936 34430
rect 3936 34396 4026 34430
rect 4026 34396 4086 34430
rect -548 34390 4086 34396
rect -770 28336 -754 34380
rect -754 28336 -716 34380
rect -716 28336 -700 34380
rect 4240 34380 4310 34520
rect -635 28378 -618 34338
rect -618 28378 -584 34338
rect -584 28378 -569 34338
rect -477 28378 -460 34338
rect -460 28378 -426 34338
rect -426 28378 -411 34338
rect -319 28378 -302 34338
rect -302 28378 -268 34338
rect -268 28378 -253 34338
rect -161 28378 -144 34338
rect -144 28378 -110 34338
rect -110 28378 -95 34338
rect -3 28378 14 34338
rect 14 28378 48 34338
rect 48 28378 63 34338
rect 155 28378 172 34338
rect 172 28378 206 34338
rect 206 28378 221 34338
rect 313 28378 330 34338
rect 330 28378 364 34338
rect 364 28378 379 34338
rect 471 28378 488 34338
rect 488 28378 522 34338
rect 522 28378 537 34338
rect 629 28378 646 34338
rect 646 28378 680 34338
rect 680 28378 695 34338
rect 787 28378 804 34338
rect 804 28378 838 34338
rect 838 28378 853 34338
rect 945 28378 962 34338
rect 962 28378 996 34338
rect 996 28378 1011 34338
rect 1103 28378 1120 34338
rect 1120 28378 1154 34338
rect 1154 28378 1169 34338
rect 1261 28378 1278 34338
rect 1278 28378 1312 34338
rect 1312 28378 1327 34338
rect 1419 28378 1436 34338
rect 1436 28378 1470 34338
rect 1470 28378 1485 34338
rect 1577 28378 1594 34338
rect 1594 28378 1628 34338
rect 1628 28378 1643 34338
rect 1735 28378 1752 34338
rect 1752 28378 1786 34338
rect 1786 28378 1801 34338
rect 1893 28378 1910 34338
rect 1910 28378 1944 34338
rect 1944 28378 1959 34338
rect 2051 28378 2068 34338
rect 2068 28378 2102 34338
rect 2102 28378 2117 34338
rect 2209 28378 2226 34338
rect 2226 28378 2260 34338
rect 2260 28378 2275 34338
rect 2367 28378 2384 34338
rect 2384 28378 2418 34338
rect 2418 28378 2433 34338
rect 2525 28378 2542 34338
rect 2542 28378 2576 34338
rect 2576 28378 2591 34338
rect 2683 28378 2700 34338
rect 2700 28378 2734 34338
rect 2734 28378 2749 34338
rect 2841 28378 2858 34338
rect 2858 28378 2892 34338
rect 2892 28378 2907 34338
rect 2999 28378 3016 34338
rect 3016 28378 3050 34338
rect 3050 28378 3065 34338
rect 3157 28378 3174 34338
rect 3174 28378 3208 34338
rect 3208 28378 3223 34338
rect 3315 28378 3332 34338
rect 3332 28378 3366 34338
rect 3366 28378 3381 34338
rect 3473 28378 3490 34338
rect 3490 28378 3524 34338
rect 3524 28378 3539 34338
rect 3631 28378 3648 34338
rect 3648 28378 3682 34338
rect 3682 28378 3697 34338
rect 3789 28378 3806 34338
rect 3806 28378 3840 34338
rect 3840 28378 3855 34338
rect 3947 28378 3964 34338
rect 3964 28378 3998 34338
rect 3998 28378 4013 34338
rect 4105 28378 4122 34338
rect 4122 28378 4156 34338
rect 4156 28378 4171 34338
rect -770 28200 -700 28336
rect 4240 28336 4254 34380
rect 4254 28336 4292 34380
rect 4292 28336 4310 34380
rect -548 28320 4086 28326
rect -548 28286 -488 28320
rect -488 28286 -398 28320
rect -398 28286 -330 28320
rect -330 28286 -240 28320
rect -240 28286 -172 28320
rect -172 28286 -82 28320
rect -82 28286 -14 28320
rect -14 28286 76 28320
rect 76 28286 144 28320
rect 144 28286 234 28320
rect 234 28286 302 28320
rect 302 28286 392 28320
rect 392 28286 460 28320
rect 460 28286 550 28320
rect 550 28286 618 28320
rect 618 28286 708 28320
rect 708 28286 776 28320
rect 776 28286 866 28320
rect 866 28286 934 28320
rect 934 28286 1024 28320
rect 1024 28286 1092 28320
rect 1092 28286 1182 28320
rect 1182 28286 1250 28320
rect 1250 28286 1340 28320
rect 1340 28286 1408 28320
rect 1408 28286 1498 28320
rect 1498 28286 1566 28320
rect 1566 28286 1656 28320
rect 1656 28286 1724 28320
rect 1724 28286 1814 28320
rect 1814 28286 1882 28320
rect 1882 28286 1972 28320
rect 1972 28286 2040 28320
rect 2040 28286 2130 28320
rect 2130 28286 2198 28320
rect 2198 28286 2288 28320
rect 2288 28286 2356 28320
rect 2356 28286 2446 28320
rect 2446 28286 2514 28320
rect 2514 28286 2604 28320
rect 2604 28286 2672 28320
rect 2672 28286 2762 28320
rect 2762 28286 2830 28320
rect 2830 28286 2920 28320
rect 2920 28286 2988 28320
rect 2988 28286 3078 28320
rect 3078 28286 3146 28320
rect 3146 28286 3236 28320
rect 3236 28286 3304 28320
rect 3304 28286 3394 28320
rect 3394 28286 3462 28320
rect 3462 28286 3552 28320
rect 3552 28286 3620 28320
rect 3620 28286 3710 28320
rect 3710 28286 3778 28320
rect 3778 28286 3868 28320
rect 3868 28286 3936 28320
rect 3936 28286 4026 28320
rect 4026 28286 4086 28320
rect -548 28226 4086 28286
rect 4240 28200 4310 28336
rect 5530 34380 5600 34520
rect 5752 34430 10386 34490
rect 5752 34396 5812 34430
rect 5812 34396 5902 34430
rect 5902 34396 5970 34430
rect 5970 34396 6060 34430
rect 6060 34396 6128 34430
rect 6128 34396 6218 34430
rect 6218 34396 6286 34430
rect 6286 34396 6376 34430
rect 6376 34396 6444 34430
rect 6444 34396 6534 34430
rect 6534 34396 6602 34430
rect 6602 34396 6692 34430
rect 6692 34396 6760 34430
rect 6760 34396 6850 34430
rect 6850 34396 6918 34430
rect 6918 34396 7008 34430
rect 7008 34396 7076 34430
rect 7076 34396 7166 34430
rect 7166 34396 7234 34430
rect 7234 34396 7324 34430
rect 7324 34396 7392 34430
rect 7392 34396 7482 34430
rect 7482 34396 7550 34430
rect 7550 34396 7640 34430
rect 7640 34396 7708 34430
rect 7708 34396 7798 34430
rect 7798 34396 7866 34430
rect 7866 34396 7956 34430
rect 7956 34396 8024 34430
rect 8024 34396 8114 34430
rect 8114 34396 8182 34430
rect 8182 34396 8272 34430
rect 8272 34396 8340 34430
rect 8340 34396 8430 34430
rect 8430 34396 8498 34430
rect 8498 34396 8588 34430
rect 8588 34396 8656 34430
rect 8656 34396 8746 34430
rect 8746 34396 8814 34430
rect 8814 34396 8904 34430
rect 8904 34396 8972 34430
rect 8972 34396 9062 34430
rect 9062 34396 9130 34430
rect 9130 34396 9220 34430
rect 9220 34396 9288 34430
rect 9288 34396 9378 34430
rect 9378 34396 9446 34430
rect 9446 34396 9536 34430
rect 9536 34396 9604 34430
rect 9604 34396 9694 34430
rect 9694 34396 9762 34430
rect 9762 34396 9852 34430
rect 9852 34396 9920 34430
rect 9920 34396 10010 34430
rect 10010 34396 10078 34430
rect 10078 34396 10168 34430
rect 10168 34396 10236 34430
rect 10236 34396 10326 34430
rect 10326 34396 10386 34430
rect 5752 34390 10386 34396
rect 5530 28336 5546 34380
rect 5546 28336 5584 34380
rect 5584 28336 5600 34380
rect 10540 34380 10610 34520
rect 5665 28378 5682 34338
rect 5682 28378 5716 34338
rect 5716 28378 5731 34338
rect 5823 28378 5840 34338
rect 5840 28378 5874 34338
rect 5874 28378 5889 34338
rect 5981 28378 5998 34338
rect 5998 28378 6032 34338
rect 6032 28378 6047 34338
rect 6139 28378 6156 34338
rect 6156 28378 6190 34338
rect 6190 28378 6205 34338
rect 6297 28378 6314 34338
rect 6314 28378 6348 34338
rect 6348 28378 6363 34338
rect 6455 28378 6472 34338
rect 6472 28378 6506 34338
rect 6506 28378 6521 34338
rect 6613 28378 6630 34338
rect 6630 28378 6664 34338
rect 6664 28378 6679 34338
rect 6771 28378 6788 34338
rect 6788 28378 6822 34338
rect 6822 28378 6837 34338
rect 6929 28378 6946 34338
rect 6946 28378 6980 34338
rect 6980 28378 6995 34338
rect 7087 28378 7104 34338
rect 7104 28378 7138 34338
rect 7138 28378 7153 34338
rect 7245 28378 7262 34338
rect 7262 28378 7296 34338
rect 7296 28378 7311 34338
rect 7403 28378 7420 34338
rect 7420 28378 7454 34338
rect 7454 28378 7469 34338
rect 7561 28378 7578 34338
rect 7578 28378 7612 34338
rect 7612 28378 7627 34338
rect 7719 28378 7736 34338
rect 7736 28378 7770 34338
rect 7770 28378 7785 34338
rect 7877 28378 7894 34338
rect 7894 28378 7928 34338
rect 7928 28378 7943 34338
rect 8035 28378 8052 34338
rect 8052 28378 8086 34338
rect 8086 28378 8101 34338
rect 8193 28378 8210 34338
rect 8210 28378 8244 34338
rect 8244 28378 8259 34338
rect 8351 28378 8368 34338
rect 8368 28378 8402 34338
rect 8402 28378 8417 34338
rect 8509 28378 8526 34338
rect 8526 28378 8560 34338
rect 8560 28378 8575 34338
rect 8667 28378 8684 34338
rect 8684 28378 8718 34338
rect 8718 28378 8733 34338
rect 8825 28378 8842 34338
rect 8842 28378 8876 34338
rect 8876 28378 8891 34338
rect 8983 28378 9000 34338
rect 9000 28378 9034 34338
rect 9034 28378 9049 34338
rect 9141 28378 9158 34338
rect 9158 28378 9192 34338
rect 9192 28378 9207 34338
rect 9299 28378 9316 34338
rect 9316 28378 9350 34338
rect 9350 28378 9365 34338
rect 9457 28378 9474 34338
rect 9474 28378 9508 34338
rect 9508 28378 9523 34338
rect 9615 28378 9632 34338
rect 9632 28378 9666 34338
rect 9666 28378 9681 34338
rect 9773 28378 9790 34338
rect 9790 28378 9824 34338
rect 9824 28378 9839 34338
rect 9931 28378 9948 34338
rect 9948 28378 9982 34338
rect 9982 28378 9997 34338
rect 10089 28378 10106 34338
rect 10106 28378 10140 34338
rect 10140 28378 10155 34338
rect 10247 28378 10264 34338
rect 10264 28378 10298 34338
rect 10298 28378 10313 34338
rect 10405 28378 10422 34338
rect 10422 28378 10456 34338
rect 10456 28378 10471 34338
rect 5530 28200 5600 28336
rect 10540 28336 10554 34380
rect 10554 28336 10592 34380
rect 10592 28336 10610 34380
rect 5752 28320 10386 28326
rect 5752 28286 5812 28320
rect 5812 28286 5902 28320
rect 5902 28286 5970 28320
rect 5970 28286 6060 28320
rect 6060 28286 6128 28320
rect 6128 28286 6218 28320
rect 6218 28286 6286 28320
rect 6286 28286 6376 28320
rect 6376 28286 6444 28320
rect 6444 28286 6534 28320
rect 6534 28286 6602 28320
rect 6602 28286 6692 28320
rect 6692 28286 6760 28320
rect 6760 28286 6850 28320
rect 6850 28286 6918 28320
rect 6918 28286 7008 28320
rect 7008 28286 7076 28320
rect 7076 28286 7166 28320
rect 7166 28286 7234 28320
rect 7234 28286 7324 28320
rect 7324 28286 7392 28320
rect 7392 28286 7482 28320
rect 7482 28286 7550 28320
rect 7550 28286 7640 28320
rect 7640 28286 7708 28320
rect 7708 28286 7798 28320
rect 7798 28286 7866 28320
rect 7866 28286 7956 28320
rect 7956 28286 8024 28320
rect 8024 28286 8114 28320
rect 8114 28286 8182 28320
rect 8182 28286 8272 28320
rect 8272 28286 8340 28320
rect 8340 28286 8430 28320
rect 8430 28286 8498 28320
rect 8498 28286 8588 28320
rect 8588 28286 8656 28320
rect 8656 28286 8746 28320
rect 8746 28286 8814 28320
rect 8814 28286 8904 28320
rect 8904 28286 8972 28320
rect 8972 28286 9062 28320
rect 9062 28286 9130 28320
rect 9130 28286 9220 28320
rect 9220 28286 9288 28320
rect 9288 28286 9378 28320
rect 9378 28286 9446 28320
rect 9446 28286 9536 28320
rect 9536 28286 9604 28320
rect 9604 28286 9694 28320
rect 9694 28286 9762 28320
rect 9762 28286 9852 28320
rect 9852 28286 9920 28320
rect 9920 28286 10010 28320
rect 10010 28286 10078 28320
rect 10078 28286 10168 28320
rect 10168 28286 10236 28320
rect 10236 28286 10326 28320
rect 10326 28286 10386 28320
rect 5752 28226 10386 28286
rect 10540 28200 10610 28336
rect -13370 27380 -13300 27520
rect -13148 27430 -8514 27490
rect -13148 27396 -13088 27430
rect -13088 27396 -12998 27430
rect -12998 27396 -12930 27430
rect -12930 27396 -12840 27430
rect -12840 27396 -12772 27430
rect -12772 27396 -12682 27430
rect -12682 27396 -12614 27430
rect -12614 27396 -12524 27430
rect -12524 27396 -12456 27430
rect -12456 27396 -12366 27430
rect -12366 27396 -12298 27430
rect -12298 27396 -12208 27430
rect -12208 27396 -12140 27430
rect -12140 27396 -12050 27430
rect -12050 27396 -11982 27430
rect -11982 27396 -11892 27430
rect -11892 27396 -11824 27430
rect -11824 27396 -11734 27430
rect -11734 27396 -11666 27430
rect -11666 27396 -11576 27430
rect -11576 27396 -11508 27430
rect -11508 27396 -11418 27430
rect -11418 27396 -11350 27430
rect -11350 27396 -11260 27430
rect -11260 27396 -11192 27430
rect -11192 27396 -11102 27430
rect -11102 27396 -11034 27430
rect -11034 27396 -10944 27430
rect -10944 27396 -10876 27430
rect -10876 27396 -10786 27430
rect -10786 27396 -10718 27430
rect -10718 27396 -10628 27430
rect -10628 27396 -10560 27430
rect -10560 27396 -10470 27430
rect -10470 27396 -10402 27430
rect -10402 27396 -10312 27430
rect -10312 27396 -10244 27430
rect -10244 27396 -10154 27430
rect -10154 27396 -10086 27430
rect -10086 27396 -9996 27430
rect -9996 27396 -9928 27430
rect -9928 27396 -9838 27430
rect -9838 27396 -9770 27430
rect -9770 27396 -9680 27430
rect -9680 27396 -9612 27430
rect -9612 27396 -9522 27430
rect -9522 27396 -9454 27430
rect -9454 27396 -9364 27430
rect -9364 27396 -9296 27430
rect -9296 27396 -9206 27430
rect -9206 27396 -9138 27430
rect -9138 27396 -9048 27430
rect -9048 27396 -8980 27430
rect -8980 27396 -8890 27430
rect -8890 27396 -8822 27430
rect -8822 27396 -8732 27430
rect -8732 27396 -8664 27430
rect -8664 27396 -8574 27430
rect -8574 27396 -8514 27430
rect -13148 27390 -8514 27396
rect -13370 21336 -13354 27380
rect -13354 21336 -13316 27380
rect -13316 21336 -13300 27380
rect -8360 27380 -8290 27520
rect -13235 21378 -13218 27338
rect -13218 21378 -13184 27338
rect -13184 21378 -13169 27338
rect -13077 21378 -13060 27338
rect -13060 21378 -13026 27338
rect -13026 21378 -13011 27338
rect -12919 21378 -12902 27338
rect -12902 21378 -12868 27338
rect -12868 21378 -12853 27338
rect -12761 21378 -12744 27338
rect -12744 21378 -12710 27338
rect -12710 21378 -12695 27338
rect -12603 21378 -12586 27338
rect -12586 21378 -12552 27338
rect -12552 21378 -12537 27338
rect -12445 21378 -12428 27338
rect -12428 21378 -12394 27338
rect -12394 21378 -12379 27338
rect -12287 21378 -12270 27338
rect -12270 21378 -12236 27338
rect -12236 21378 -12221 27338
rect -12129 21378 -12112 27338
rect -12112 21378 -12078 27338
rect -12078 21378 -12063 27338
rect -11971 21378 -11954 27338
rect -11954 21378 -11920 27338
rect -11920 21378 -11905 27338
rect -11813 21378 -11796 27338
rect -11796 21378 -11762 27338
rect -11762 21378 -11747 27338
rect -11655 21378 -11638 27338
rect -11638 21378 -11604 27338
rect -11604 21378 -11589 27338
rect -11497 21378 -11480 27338
rect -11480 21378 -11446 27338
rect -11446 21378 -11431 27338
rect -11339 21378 -11322 27338
rect -11322 21378 -11288 27338
rect -11288 21378 -11273 27338
rect -11181 21378 -11164 27338
rect -11164 21378 -11130 27338
rect -11130 21378 -11115 27338
rect -11023 21378 -11006 27338
rect -11006 21378 -10972 27338
rect -10972 21378 -10957 27338
rect -10865 21378 -10848 27338
rect -10848 21378 -10814 27338
rect -10814 21378 -10799 27338
rect -10707 21378 -10690 27338
rect -10690 21378 -10656 27338
rect -10656 21378 -10641 27338
rect -10549 21378 -10532 27338
rect -10532 21378 -10498 27338
rect -10498 21378 -10483 27338
rect -10391 21378 -10374 27338
rect -10374 21378 -10340 27338
rect -10340 21378 -10325 27338
rect -10233 21378 -10216 27338
rect -10216 21378 -10182 27338
rect -10182 21378 -10167 27338
rect -10075 21378 -10058 27338
rect -10058 21378 -10024 27338
rect -10024 21378 -10009 27338
rect -9917 21378 -9900 27338
rect -9900 21378 -9866 27338
rect -9866 21378 -9851 27338
rect -9759 21378 -9742 27338
rect -9742 21378 -9708 27338
rect -9708 21378 -9693 27338
rect -9601 21378 -9584 27338
rect -9584 21378 -9550 27338
rect -9550 21378 -9535 27338
rect -9443 21378 -9426 27338
rect -9426 21378 -9392 27338
rect -9392 21378 -9377 27338
rect -9285 21378 -9268 27338
rect -9268 21378 -9234 27338
rect -9234 21378 -9219 27338
rect -9127 21378 -9110 27338
rect -9110 21378 -9076 27338
rect -9076 21378 -9061 27338
rect -8969 21378 -8952 27338
rect -8952 21378 -8918 27338
rect -8918 21378 -8903 27338
rect -8811 21378 -8794 27338
rect -8794 21378 -8760 27338
rect -8760 21378 -8745 27338
rect -8653 21378 -8636 27338
rect -8636 21378 -8602 27338
rect -8602 21378 -8587 27338
rect -8495 21378 -8478 27338
rect -8478 21378 -8444 27338
rect -8444 21378 -8429 27338
rect -13370 21200 -13300 21336
rect -8360 21336 -8346 27380
rect -8346 21336 -8308 27380
rect -8308 21336 -8290 27380
rect -13148 21320 -8514 21326
rect -13148 21286 -13088 21320
rect -13088 21286 -12998 21320
rect -12998 21286 -12930 21320
rect -12930 21286 -12840 21320
rect -12840 21286 -12772 21320
rect -12772 21286 -12682 21320
rect -12682 21286 -12614 21320
rect -12614 21286 -12524 21320
rect -12524 21286 -12456 21320
rect -12456 21286 -12366 21320
rect -12366 21286 -12298 21320
rect -12298 21286 -12208 21320
rect -12208 21286 -12140 21320
rect -12140 21286 -12050 21320
rect -12050 21286 -11982 21320
rect -11982 21286 -11892 21320
rect -11892 21286 -11824 21320
rect -11824 21286 -11734 21320
rect -11734 21286 -11666 21320
rect -11666 21286 -11576 21320
rect -11576 21286 -11508 21320
rect -11508 21286 -11418 21320
rect -11418 21286 -11350 21320
rect -11350 21286 -11260 21320
rect -11260 21286 -11192 21320
rect -11192 21286 -11102 21320
rect -11102 21286 -11034 21320
rect -11034 21286 -10944 21320
rect -10944 21286 -10876 21320
rect -10876 21286 -10786 21320
rect -10786 21286 -10718 21320
rect -10718 21286 -10628 21320
rect -10628 21286 -10560 21320
rect -10560 21286 -10470 21320
rect -10470 21286 -10402 21320
rect -10402 21286 -10312 21320
rect -10312 21286 -10244 21320
rect -10244 21286 -10154 21320
rect -10154 21286 -10086 21320
rect -10086 21286 -9996 21320
rect -9996 21286 -9928 21320
rect -9928 21286 -9838 21320
rect -9838 21286 -9770 21320
rect -9770 21286 -9680 21320
rect -9680 21286 -9612 21320
rect -9612 21286 -9522 21320
rect -9522 21286 -9454 21320
rect -9454 21286 -9364 21320
rect -9364 21286 -9296 21320
rect -9296 21286 -9206 21320
rect -9206 21286 -9138 21320
rect -9138 21286 -9048 21320
rect -9048 21286 -8980 21320
rect -8980 21286 -8890 21320
rect -8890 21286 -8822 21320
rect -8822 21286 -8732 21320
rect -8732 21286 -8664 21320
rect -8664 21286 -8574 21320
rect -8574 21286 -8514 21320
rect -13148 21226 -8514 21286
rect -8360 21200 -8290 21336
rect -7070 27380 -7000 27520
rect -6848 27430 -2214 27490
rect -6848 27396 -6788 27430
rect -6788 27396 -6698 27430
rect -6698 27396 -6630 27430
rect -6630 27396 -6540 27430
rect -6540 27396 -6472 27430
rect -6472 27396 -6382 27430
rect -6382 27396 -6314 27430
rect -6314 27396 -6224 27430
rect -6224 27396 -6156 27430
rect -6156 27396 -6066 27430
rect -6066 27396 -5998 27430
rect -5998 27396 -5908 27430
rect -5908 27396 -5840 27430
rect -5840 27396 -5750 27430
rect -5750 27396 -5682 27430
rect -5682 27396 -5592 27430
rect -5592 27396 -5524 27430
rect -5524 27396 -5434 27430
rect -5434 27396 -5366 27430
rect -5366 27396 -5276 27430
rect -5276 27396 -5208 27430
rect -5208 27396 -5118 27430
rect -5118 27396 -5050 27430
rect -5050 27396 -4960 27430
rect -4960 27396 -4892 27430
rect -4892 27396 -4802 27430
rect -4802 27396 -4734 27430
rect -4734 27396 -4644 27430
rect -4644 27396 -4576 27430
rect -4576 27396 -4486 27430
rect -4486 27396 -4418 27430
rect -4418 27396 -4328 27430
rect -4328 27396 -4260 27430
rect -4260 27396 -4170 27430
rect -4170 27396 -4102 27430
rect -4102 27396 -4012 27430
rect -4012 27396 -3944 27430
rect -3944 27396 -3854 27430
rect -3854 27396 -3786 27430
rect -3786 27396 -3696 27430
rect -3696 27396 -3628 27430
rect -3628 27396 -3538 27430
rect -3538 27396 -3470 27430
rect -3470 27396 -3380 27430
rect -3380 27396 -3312 27430
rect -3312 27396 -3222 27430
rect -3222 27396 -3154 27430
rect -3154 27396 -3064 27430
rect -3064 27396 -2996 27430
rect -2996 27396 -2906 27430
rect -2906 27396 -2838 27430
rect -2838 27396 -2748 27430
rect -2748 27396 -2680 27430
rect -2680 27396 -2590 27430
rect -2590 27396 -2522 27430
rect -2522 27396 -2432 27430
rect -2432 27396 -2364 27430
rect -2364 27396 -2274 27430
rect -2274 27396 -2214 27430
rect -6848 27390 -2214 27396
rect -7070 21336 -7054 27380
rect -7054 21336 -7016 27380
rect -7016 21336 -7000 27380
rect -2060 27380 -1990 27520
rect -6935 21378 -6918 27338
rect -6918 21378 -6884 27338
rect -6884 21378 -6869 27338
rect -6777 21378 -6760 27338
rect -6760 21378 -6726 27338
rect -6726 21378 -6711 27338
rect -6619 21378 -6602 27338
rect -6602 21378 -6568 27338
rect -6568 21378 -6553 27338
rect -6461 21378 -6444 27338
rect -6444 21378 -6410 27338
rect -6410 21378 -6395 27338
rect -6303 21378 -6286 27338
rect -6286 21378 -6252 27338
rect -6252 21378 -6237 27338
rect -6145 21378 -6128 27338
rect -6128 21378 -6094 27338
rect -6094 21378 -6079 27338
rect -5987 21378 -5970 27338
rect -5970 21378 -5936 27338
rect -5936 21378 -5921 27338
rect -5829 21378 -5812 27338
rect -5812 21378 -5778 27338
rect -5778 21378 -5763 27338
rect -5671 21378 -5654 27338
rect -5654 21378 -5620 27338
rect -5620 21378 -5605 27338
rect -5513 21378 -5496 27338
rect -5496 21378 -5462 27338
rect -5462 21378 -5447 27338
rect -5355 21378 -5338 27338
rect -5338 21378 -5304 27338
rect -5304 21378 -5289 27338
rect -5197 21378 -5180 27338
rect -5180 21378 -5146 27338
rect -5146 21378 -5131 27338
rect -5039 21378 -5022 27338
rect -5022 21378 -4988 27338
rect -4988 21378 -4973 27338
rect -4881 21378 -4864 27338
rect -4864 21378 -4830 27338
rect -4830 21378 -4815 27338
rect -4723 21378 -4706 27338
rect -4706 21378 -4672 27338
rect -4672 21378 -4657 27338
rect -4565 21378 -4548 27338
rect -4548 21378 -4514 27338
rect -4514 21378 -4499 27338
rect -4407 21378 -4390 27338
rect -4390 21378 -4356 27338
rect -4356 21378 -4341 27338
rect -4249 21378 -4232 27338
rect -4232 21378 -4198 27338
rect -4198 21378 -4183 27338
rect -4091 21378 -4074 27338
rect -4074 21378 -4040 27338
rect -4040 21378 -4025 27338
rect -3933 21378 -3916 27338
rect -3916 21378 -3882 27338
rect -3882 21378 -3867 27338
rect -3775 21378 -3758 27338
rect -3758 21378 -3724 27338
rect -3724 21378 -3709 27338
rect -3617 21378 -3600 27338
rect -3600 21378 -3566 27338
rect -3566 21378 -3551 27338
rect -3459 21378 -3442 27338
rect -3442 21378 -3408 27338
rect -3408 21378 -3393 27338
rect -3301 21378 -3284 27338
rect -3284 21378 -3250 27338
rect -3250 21378 -3235 27338
rect -3143 21378 -3126 27338
rect -3126 21378 -3092 27338
rect -3092 21378 -3077 27338
rect -2985 21378 -2968 27338
rect -2968 21378 -2934 27338
rect -2934 21378 -2919 27338
rect -2827 21378 -2810 27338
rect -2810 21378 -2776 27338
rect -2776 21378 -2761 27338
rect -2669 21378 -2652 27338
rect -2652 21378 -2618 27338
rect -2618 21378 -2603 27338
rect -2511 21378 -2494 27338
rect -2494 21378 -2460 27338
rect -2460 21378 -2445 27338
rect -2353 21378 -2336 27338
rect -2336 21378 -2302 27338
rect -2302 21378 -2287 27338
rect -2195 21378 -2178 27338
rect -2178 21378 -2144 27338
rect -2144 21378 -2129 27338
rect -7070 21200 -7000 21336
rect -2060 21336 -2046 27380
rect -2046 21336 -2008 27380
rect -2008 21336 -1990 27380
rect -6848 21320 -2214 21326
rect -6848 21286 -6788 21320
rect -6788 21286 -6698 21320
rect -6698 21286 -6630 21320
rect -6630 21286 -6540 21320
rect -6540 21286 -6472 21320
rect -6472 21286 -6382 21320
rect -6382 21286 -6314 21320
rect -6314 21286 -6224 21320
rect -6224 21286 -6156 21320
rect -6156 21286 -6066 21320
rect -6066 21286 -5998 21320
rect -5998 21286 -5908 21320
rect -5908 21286 -5840 21320
rect -5840 21286 -5750 21320
rect -5750 21286 -5682 21320
rect -5682 21286 -5592 21320
rect -5592 21286 -5524 21320
rect -5524 21286 -5434 21320
rect -5434 21286 -5366 21320
rect -5366 21286 -5276 21320
rect -5276 21286 -5208 21320
rect -5208 21286 -5118 21320
rect -5118 21286 -5050 21320
rect -5050 21286 -4960 21320
rect -4960 21286 -4892 21320
rect -4892 21286 -4802 21320
rect -4802 21286 -4734 21320
rect -4734 21286 -4644 21320
rect -4644 21286 -4576 21320
rect -4576 21286 -4486 21320
rect -4486 21286 -4418 21320
rect -4418 21286 -4328 21320
rect -4328 21286 -4260 21320
rect -4260 21286 -4170 21320
rect -4170 21286 -4102 21320
rect -4102 21286 -4012 21320
rect -4012 21286 -3944 21320
rect -3944 21286 -3854 21320
rect -3854 21286 -3786 21320
rect -3786 21286 -3696 21320
rect -3696 21286 -3628 21320
rect -3628 21286 -3538 21320
rect -3538 21286 -3470 21320
rect -3470 21286 -3380 21320
rect -3380 21286 -3312 21320
rect -3312 21286 -3222 21320
rect -3222 21286 -3154 21320
rect -3154 21286 -3064 21320
rect -3064 21286 -2996 21320
rect -2996 21286 -2906 21320
rect -2906 21286 -2838 21320
rect -2838 21286 -2748 21320
rect -2748 21286 -2680 21320
rect -2680 21286 -2590 21320
rect -2590 21286 -2522 21320
rect -2522 21286 -2432 21320
rect -2432 21286 -2364 21320
rect -2364 21286 -2274 21320
rect -2274 21286 -2214 21320
rect -6848 21226 -2214 21286
rect -2060 21200 -1990 21336
rect -770 27380 -700 27520
rect -548 27430 4086 27490
rect -548 27396 -488 27430
rect -488 27396 -398 27430
rect -398 27396 -330 27430
rect -330 27396 -240 27430
rect -240 27396 -172 27430
rect -172 27396 -82 27430
rect -82 27396 -14 27430
rect -14 27396 76 27430
rect 76 27396 144 27430
rect 144 27396 234 27430
rect 234 27396 302 27430
rect 302 27396 392 27430
rect 392 27396 460 27430
rect 460 27396 550 27430
rect 550 27396 618 27430
rect 618 27396 708 27430
rect 708 27396 776 27430
rect 776 27396 866 27430
rect 866 27396 934 27430
rect 934 27396 1024 27430
rect 1024 27396 1092 27430
rect 1092 27396 1182 27430
rect 1182 27396 1250 27430
rect 1250 27396 1340 27430
rect 1340 27396 1408 27430
rect 1408 27396 1498 27430
rect 1498 27396 1566 27430
rect 1566 27396 1656 27430
rect 1656 27396 1724 27430
rect 1724 27396 1814 27430
rect 1814 27396 1882 27430
rect 1882 27396 1972 27430
rect 1972 27396 2040 27430
rect 2040 27396 2130 27430
rect 2130 27396 2198 27430
rect 2198 27396 2288 27430
rect 2288 27396 2356 27430
rect 2356 27396 2446 27430
rect 2446 27396 2514 27430
rect 2514 27396 2604 27430
rect 2604 27396 2672 27430
rect 2672 27396 2762 27430
rect 2762 27396 2830 27430
rect 2830 27396 2920 27430
rect 2920 27396 2988 27430
rect 2988 27396 3078 27430
rect 3078 27396 3146 27430
rect 3146 27396 3236 27430
rect 3236 27396 3304 27430
rect 3304 27396 3394 27430
rect 3394 27396 3462 27430
rect 3462 27396 3552 27430
rect 3552 27396 3620 27430
rect 3620 27396 3710 27430
rect 3710 27396 3778 27430
rect 3778 27396 3868 27430
rect 3868 27396 3936 27430
rect 3936 27396 4026 27430
rect 4026 27396 4086 27430
rect -548 27390 4086 27396
rect -770 21336 -754 27380
rect -754 21336 -716 27380
rect -716 21336 -700 27380
rect 4240 27380 4310 27520
rect -635 21378 -618 27338
rect -618 21378 -584 27338
rect -584 21378 -569 27338
rect -477 21378 -460 27338
rect -460 21378 -426 27338
rect -426 21378 -411 27338
rect -319 21378 -302 27338
rect -302 21378 -268 27338
rect -268 21378 -253 27338
rect -161 21378 -144 27338
rect -144 21378 -110 27338
rect -110 21378 -95 27338
rect -3 21378 14 27338
rect 14 21378 48 27338
rect 48 21378 63 27338
rect 155 21378 172 27338
rect 172 21378 206 27338
rect 206 21378 221 27338
rect 313 21378 330 27338
rect 330 21378 364 27338
rect 364 21378 379 27338
rect 471 21378 488 27338
rect 488 21378 522 27338
rect 522 21378 537 27338
rect 629 21378 646 27338
rect 646 21378 680 27338
rect 680 21378 695 27338
rect 787 21378 804 27338
rect 804 21378 838 27338
rect 838 21378 853 27338
rect 945 21378 962 27338
rect 962 21378 996 27338
rect 996 21378 1011 27338
rect 1103 21378 1120 27338
rect 1120 21378 1154 27338
rect 1154 21378 1169 27338
rect 1261 21378 1278 27338
rect 1278 21378 1312 27338
rect 1312 21378 1327 27338
rect 1419 21378 1436 27338
rect 1436 21378 1470 27338
rect 1470 21378 1485 27338
rect 1577 21378 1594 27338
rect 1594 21378 1628 27338
rect 1628 21378 1643 27338
rect 1735 21378 1752 27338
rect 1752 21378 1786 27338
rect 1786 21378 1801 27338
rect 1893 21378 1910 27338
rect 1910 21378 1944 27338
rect 1944 21378 1959 27338
rect 2051 21378 2068 27338
rect 2068 21378 2102 27338
rect 2102 21378 2117 27338
rect 2209 21378 2226 27338
rect 2226 21378 2260 27338
rect 2260 21378 2275 27338
rect 2367 21378 2384 27338
rect 2384 21378 2418 27338
rect 2418 21378 2433 27338
rect 2525 21378 2542 27338
rect 2542 21378 2576 27338
rect 2576 21378 2591 27338
rect 2683 21378 2700 27338
rect 2700 21378 2734 27338
rect 2734 21378 2749 27338
rect 2841 21378 2858 27338
rect 2858 21378 2892 27338
rect 2892 21378 2907 27338
rect 2999 21378 3016 27338
rect 3016 21378 3050 27338
rect 3050 21378 3065 27338
rect 3157 21378 3174 27338
rect 3174 21378 3208 27338
rect 3208 21378 3223 27338
rect 3315 21378 3332 27338
rect 3332 21378 3366 27338
rect 3366 21378 3381 27338
rect 3473 21378 3490 27338
rect 3490 21378 3524 27338
rect 3524 21378 3539 27338
rect 3631 21378 3648 27338
rect 3648 21378 3682 27338
rect 3682 21378 3697 27338
rect 3789 21378 3806 27338
rect 3806 21378 3840 27338
rect 3840 21378 3855 27338
rect 3947 21378 3964 27338
rect 3964 21378 3998 27338
rect 3998 21378 4013 27338
rect 4105 21378 4122 27338
rect 4122 21378 4156 27338
rect 4156 21378 4171 27338
rect -770 21200 -700 21336
rect 4240 21336 4254 27380
rect 4254 21336 4292 27380
rect 4292 21336 4310 27380
rect -548 21320 4086 21326
rect -548 21286 -488 21320
rect -488 21286 -398 21320
rect -398 21286 -330 21320
rect -330 21286 -240 21320
rect -240 21286 -172 21320
rect -172 21286 -82 21320
rect -82 21286 -14 21320
rect -14 21286 76 21320
rect 76 21286 144 21320
rect 144 21286 234 21320
rect 234 21286 302 21320
rect 302 21286 392 21320
rect 392 21286 460 21320
rect 460 21286 550 21320
rect 550 21286 618 21320
rect 618 21286 708 21320
rect 708 21286 776 21320
rect 776 21286 866 21320
rect 866 21286 934 21320
rect 934 21286 1024 21320
rect 1024 21286 1092 21320
rect 1092 21286 1182 21320
rect 1182 21286 1250 21320
rect 1250 21286 1340 21320
rect 1340 21286 1408 21320
rect 1408 21286 1498 21320
rect 1498 21286 1566 21320
rect 1566 21286 1656 21320
rect 1656 21286 1724 21320
rect 1724 21286 1814 21320
rect 1814 21286 1882 21320
rect 1882 21286 1972 21320
rect 1972 21286 2040 21320
rect 2040 21286 2130 21320
rect 2130 21286 2198 21320
rect 2198 21286 2288 21320
rect 2288 21286 2356 21320
rect 2356 21286 2446 21320
rect 2446 21286 2514 21320
rect 2514 21286 2604 21320
rect 2604 21286 2672 21320
rect 2672 21286 2762 21320
rect 2762 21286 2830 21320
rect 2830 21286 2920 21320
rect 2920 21286 2988 21320
rect 2988 21286 3078 21320
rect 3078 21286 3146 21320
rect 3146 21286 3236 21320
rect 3236 21286 3304 21320
rect 3304 21286 3394 21320
rect 3394 21286 3462 21320
rect 3462 21286 3552 21320
rect 3552 21286 3620 21320
rect 3620 21286 3710 21320
rect 3710 21286 3778 21320
rect 3778 21286 3868 21320
rect 3868 21286 3936 21320
rect 3936 21286 4026 21320
rect 4026 21286 4086 21320
rect -548 21226 4086 21286
rect 4240 21200 4310 21336
rect 5530 27380 5600 27520
rect 5752 27430 10386 27490
rect 5752 27396 5812 27430
rect 5812 27396 5902 27430
rect 5902 27396 5970 27430
rect 5970 27396 6060 27430
rect 6060 27396 6128 27430
rect 6128 27396 6218 27430
rect 6218 27396 6286 27430
rect 6286 27396 6376 27430
rect 6376 27396 6444 27430
rect 6444 27396 6534 27430
rect 6534 27396 6602 27430
rect 6602 27396 6692 27430
rect 6692 27396 6760 27430
rect 6760 27396 6850 27430
rect 6850 27396 6918 27430
rect 6918 27396 7008 27430
rect 7008 27396 7076 27430
rect 7076 27396 7166 27430
rect 7166 27396 7234 27430
rect 7234 27396 7324 27430
rect 7324 27396 7392 27430
rect 7392 27396 7482 27430
rect 7482 27396 7550 27430
rect 7550 27396 7640 27430
rect 7640 27396 7708 27430
rect 7708 27396 7798 27430
rect 7798 27396 7866 27430
rect 7866 27396 7956 27430
rect 7956 27396 8024 27430
rect 8024 27396 8114 27430
rect 8114 27396 8182 27430
rect 8182 27396 8272 27430
rect 8272 27396 8340 27430
rect 8340 27396 8430 27430
rect 8430 27396 8498 27430
rect 8498 27396 8588 27430
rect 8588 27396 8656 27430
rect 8656 27396 8746 27430
rect 8746 27396 8814 27430
rect 8814 27396 8904 27430
rect 8904 27396 8972 27430
rect 8972 27396 9062 27430
rect 9062 27396 9130 27430
rect 9130 27396 9220 27430
rect 9220 27396 9288 27430
rect 9288 27396 9378 27430
rect 9378 27396 9446 27430
rect 9446 27396 9536 27430
rect 9536 27396 9604 27430
rect 9604 27396 9694 27430
rect 9694 27396 9762 27430
rect 9762 27396 9852 27430
rect 9852 27396 9920 27430
rect 9920 27396 10010 27430
rect 10010 27396 10078 27430
rect 10078 27396 10168 27430
rect 10168 27396 10236 27430
rect 10236 27396 10326 27430
rect 10326 27396 10386 27430
rect 5752 27390 10386 27396
rect 5530 21336 5546 27380
rect 5546 21336 5584 27380
rect 5584 21336 5600 27380
rect 10540 27380 10610 27520
rect 5665 21378 5682 27338
rect 5682 21378 5716 27338
rect 5716 21378 5731 27338
rect 5823 21378 5840 27338
rect 5840 21378 5874 27338
rect 5874 21378 5889 27338
rect 5981 21378 5998 27338
rect 5998 21378 6032 27338
rect 6032 21378 6047 27338
rect 6139 21378 6156 27338
rect 6156 21378 6190 27338
rect 6190 21378 6205 27338
rect 6297 21378 6314 27338
rect 6314 21378 6348 27338
rect 6348 21378 6363 27338
rect 6455 21378 6472 27338
rect 6472 21378 6506 27338
rect 6506 21378 6521 27338
rect 6613 21378 6630 27338
rect 6630 21378 6664 27338
rect 6664 21378 6679 27338
rect 6771 21378 6788 27338
rect 6788 21378 6822 27338
rect 6822 21378 6837 27338
rect 6929 21378 6946 27338
rect 6946 21378 6980 27338
rect 6980 21378 6995 27338
rect 7087 21378 7104 27338
rect 7104 21378 7138 27338
rect 7138 21378 7153 27338
rect 7245 21378 7262 27338
rect 7262 21378 7296 27338
rect 7296 21378 7311 27338
rect 7403 21378 7420 27338
rect 7420 21378 7454 27338
rect 7454 21378 7469 27338
rect 7561 21378 7578 27338
rect 7578 21378 7612 27338
rect 7612 21378 7627 27338
rect 7719 21378 7736 27338
rect 7736 21378 7770 27338
rect 7770 21378 7785 27338
rect 7877 21378 7894 27338
rect 7894 21378 7928 27338
rect 7928 21378 7943 27338
rect 8035 21378 8052 27338
rect 8052 21378 8086 27338
rect 8086 21378 8101 27338
rect 8193 21378 8210 27338
rect 8210 21378 8244 27338
rect 8244 21378 8259 27338
rect 8351 21378 8368 27338
rect 8368 21378 8402 27338
rect 8402 21378 8417 27338
rect 8509 21378 8526 27338
rect 8526 21378 8560 27338
rect 8560 21378 8575 27338
rect 8667 21378 8684 27338
rect 8684 21378 8718 27338
rect 8718 21378 8733 27338
rect 8825 21378 8842 27338
rect 8842 21378 8876 27338
rect 8876 21378 8891 27338
rect 8983 21378 9000 27338
rect 9000 21378 9034 27338
rect 9034 21378 9049 27338
rect 9141 21378 9158 27338
rect 9158 21378 9192 27338
rect 9192 21378 9207 27338
rect 9299 21378 9316 27338
rect 9316 21378 9350 27338
rect 9350 21378 9365 27338
rect 9457 21378 9474 27338
rect 9474 21378 9508 27338
rect 9508 21378 9523 27338
rect 9615 21378 9632 27338
rect 9632 21378 9666 27338
rect 9666 21378 9681 27338
rect 9773 21378 9790 27338
rect 9790 21378 9824 27338
rect 9824 21378 9839 27338
rect 9931 21378 9948 27338
rect 9948 21378 9982 27338
rect 9982 21378 9997 27338
rect 10089 21378 10106 27338
rect 10106 21378 10140 27338
rect 10140 21378 10155 27338
rect 10247 21378 10264 27338
rect 10264 21378 10298 27338
rect 10298 21378 10313 27338
rect 10405 21378 10422 27338
rect 10422 21378 10456 27338
rect 10456 21378 10471 27338
rect 5530 21200 5600 21336
rect 10540 21336 10554 27380
rect 10554 21336 10592 27380
rect 10592 21336 10610 27380
rect 5752 21320 10386 21326
rect 5752 21286 5812 21320
rect 5812 21286 5902 21320
rect 5902 21286 5970 21320
rect 5970 21286 6060 21320
rect 6060 21286 6128 21320
rect 6128 21286 6218 21320
rect 6218 21286 6286 21320
rect 6286 21286 6376 21320
rect 6376 21286 6444 21320
rect 6444 21286 6534 21320
rect 6534 21286 6602 21320
rect 6602 21286 6692 21320
rect 6692 21286 6760 21320
rect 6760 21286 6850 21320
rect 6850 21286 6918 21320
rect 6918 21286 7008 21320
rect 7008 21286 7076 21320
rect 7076 21286 7166 21320
rect 7166 21286 7234 21320
rect 7234 21286 7324 21320
rect 7324 21286 7392 21320
rect 7392 21286 7482 21320
rect 7482 21286 7550 21320
rect 7550 21286 7640 21320
rect 7640 21286 7708 21320
rect 7708 21286 7798 21320
rect 7798 21286 7866 21320
rect 7866 21286 7956 21320
rect 7956 21286 8024 21320
rect 8024 21286 8114 21320
rect 8114 21286 8182 21320
rect 8182 21286 8272 21320
rect 8272 21286 8340 21320
rect 8340 21286 8430 21320
rect 8430 21286 8498 21320
rect 8498 21286 8588 21320
rect 8588 21286 8656 21320
rect 8656 21286 8746 21320
rect 8746 21286 8814 21320
rect 8814 21286 8904 21320
rect 8904 21286 8972 21320
rect 8972 21286 9062 21320
rect 9062 21286 9130 21320
rect 9130 21286 9220 21320
rect 9220 21286 9288 21320
rect 9288 21286 9378 21320
rect 9378 21286 9446 21320
rect 9446 21286 9536 21320
rect 9536 21286 9604 21320
rect 9604 21286 9694 21320
rect 9694 21286 9762 21320
rect 9762 21286 9852 21320
rect 9852 21286 9920 21320
rect 9920 21286 10010 21320
rect 10010 21286 10078 21320
rect 10078 21286 10168 21320
rect 10168 21286 10236 21320
rect 10236 21286 10326 21320
rect 10326 21286 10386 21320
rect 5752 21226 10386 21286
rect 10540 21200 10610 21336
rect -13370 19080 -13300 19220
rect -13148 19130 -8514 19190
rect -13148 19096 -13088 19130
rect -13088 19096 -12998 19130
rect -12998 19096 -12930 19130
rect -12930 19096 -12840 19130
rect -12840 19096 -12772 19130
rect -12772 19096 -12682 19130
rect -12682 19096 -12614 19130
rect -12614 19096 -12524 19130
rect -12524 19096 -12456 19130
rect -12456 19096 -12366 19130
rect -12366 19096 -12298 19130
rect -12298 19096 -12208 19130
rect -12208 19096 -12140 19130
rect -12140 19096 -12050 19130
rect -12050 19096 -11982 19130
rect -11982 19096 -11892 19130
rect -11892 19096 -11824 19130
rect -11824 19096 -11734 19130
rect -11734 19096 -11666 19130
rect -11666 19096 -11576 19130
rect -11576 19096 -11508 19130
rect -11508 19096 -11418 19130
rect -11418 19096 -11350 19130
rect -11350 19096 -11260 19130
rect -11260 19096 -11192 19130
rect -11192 19096 -11102 19130
rect -11102 19096 -11034 19130
rect -11034 19096 -10944 19130
rect -10944 19096 -10876 19130
rect -10876 19096 -10786 19130
rect -10786 19096 -10718 19130
rect -10718 19096 -10628 19130
rect -10628 19096 -10560 19130
rect -10560 19096 -10470 19130
rect -10470 19096 -10402 19130
rect -10402 19096 -10312 19130
rect -10312 19096 -10244 19130
rect -10244 19096 -10154 19130
rect -10154 19096 -10086 19130
rect -10086 19096 -9996 19130
rect -9996 19096 -9928 19130
rect -9928 19096 -9838 19130
rect -9838 19096 -9770 19130
rect -9770 19096 -9680 19130
rect -9680 19096 -9612 19130
rect -9612 19096 -9522 19130
rect -9522 19096 -9454 19130
rect -9454 19096 -9364 19130
rect -9364 19096 -9296 19130
rect -9296 19096 -9206 19130
rect -9206 19096 -9138 19130
rect -9138 19096 -9048 19130
rect -9048 19096 -8980 19130
rect -8980 19096 -8890 19130
rect -8890 19096 -8822 19130
rect -8822 19096 -8732 19130
rect -8732 19096 -8664 19130
rect -8664 19096 -8574 19130
rect -8574 19096 -8514 19130
rect -13148 19090 -8514 19096
rect -13370 13036 -13354 19080
rect -13354 13036 -13316 19080
rect -13316 13036 -13300 19080
rect -8360 19080 -8290 19220
rect -13235 13078 -13218 19038
rect -13218 13078 -13184 19038
rect -13184 13078 -13169 19038
rect -13077 13078 -13060 19038
rect -13060 13078 -13026 19038
rect -13026 13078 -13011 19038
rect -12919 13078 -12902 19038
rect -12902 13078 -12868 19038
rect -12868 13078 -12853 19038
rect -12761 13078 -12744 19038
rect -12744 13078 -12710 19038
rect -12710 13078 -12695 19038
rect -12603 13078 -12586 19038
rect -12586 13078 -12552 19038
rect -12552 13078 -12537 19038
rect -12445 13078 -12428 19038
rect -12428 13078 -12394 19038
rect -12394 13078 -12379 19038
rect -12287 13078 -12270 19038
rect -12270 13078 -12236 19038
rect -12236 13078 -12221 19038
rect -12129 13078 -12112 19038
rect -12112 13078 -12078 19038
rect -12078 13078 -12063 19038
rect -11971 13078 -11954 19038
rect -11954 13078 -11920 19038
rect -11920 13078 -11905 19038
rect -11813 13078 -11796 19038
rect -11796 13078 -11762 19038
rect -11762 13078 -11747 19038
rect -11655 13078 -11638 19038
rect -11638 13078 -11604 19038
rect -11604 13078 -11589 19038
rect -11497 13078 -11480 19038
rect -11480 13078 -11446 19038
rect -11446 13078 -11431 19038
rect -11339 13078 -11322 19038
rect -11322 13078 -11288 19038
rect -11288 13078 -11273 19038
rect -11181 13078 -11164 19038
rect -11164 13078 -11130 19038
rect -11130 13078 -11115 19038
rect -11023 13078 -11006 19038
rect -11006 13078 -10972 19038
rect -10972 13078 -10957 19038
rect -10865 13078 -10848 19038
rect -10848 13078 -10814 19038
rect -10814 13078 -10799 19038
rect -10707 13078 -10690 19038
rect -10690 13078 -10656 19038
rect -10656 13078 -10641 19038
rect -10549 13078 -10532 19038
rect -10532 13078 -10498 19038
rect -10498 13078 -10483 19038
rect -10391 13078 -10374 19038
rect -10374 13078 -10340 19038
rect -10340 13078 -10325 19038
rect -10233 13078 -10216 19038
rect -10216 13078 -10182 19038
rect -10182 13078 -10167 19038
rect -10075 13078 -10058 19038
rect -10058 13078 -10024 19038
rect -10024 13078 -10009 19038
rect -9917 13078 -9900 19038
rect -9900 13078 -9866 19038
rect -9866 13078 -9851 19038
rect -9759 13078 -9742 19038
rect -9742 13078 -9708 19038
rect -9708 13078 -9693 19038
rect -9601 13078 -9584 19038
rect -9584 13078 -9550 19038
rect -9550 13078 -9535 19038
rect -9443 13078 -9426 19038
rect -9426 13078 -9392 19038
rect -9392 13078 -9377 19038
rect -9285 13078 -9268 19038
rect -9268 13078 -9234 19038
rect -9234 13078 -9219 19038
rect -9127 13078 -9110 19038
rect -9110 13078 -9076 19038
rect -9076 13078 -9061 19038
rect -8969 13078 -8952 19038
rect -8952 13078 -8918 19038
rect -8918 13078 -8903 19038
rect -8811 13078 -8794 19038
rect -8794 13078 -8760 19038
rect -8760 13078 -8745 19038
rect -8653 13078 -8636 19038
rect -8636 13078 -8602 19038
rect -8602 13078 -8587 19038
rect -8495 13078 -8478 19038
rect -8478 13078 -8444 19038
rect -8444 13078 -8429 19038
rect -13370 12900 -13300 13036
rect -8360 13036 -8346 19080
rect -8346 13036 -8308 19080
rect -8308 13036 -8290 19080
rect -13148 13020 -8514 13026
rect -13148 12986 -13088 13020
rect -13088 12986 -12998 13020
rect -12998 12986 -12930 13020
rect -12930 12986 -12840 13020
rect -12840 12986 -12772 13020
rect -12772 12986 -12682 13020
rect -12682 12986 -12614 13020
rect -12614 12986 -12524 13020
rect -12524 12986 -12456 13020
rect -12456 12986 -12366 13020
rect -12366 12986 -12298 13020
rect -12298 12986 -12208 13020
rect -12208 12986 -12140 13020
rect -12140 12986 -12050 13020
rect -12050 12986 -11982 13020
rect -11982 12986 -11892 13020
rect -11892 12986 -11824 13020
rect -11824 12986 -11734 13020
rect -11734 12986 -11666 13020
rect -11666 12986 -11576 13020
rect -11576 12986 -11508 13020
rect -11508 12986 -11418 13020
rect -11418 12986 -11350 13020
rect -11350 12986 -11260 13020
rect -11260 12986 -11192 13020
rect -11192 12986 -11102 13020
rect -11102 12986 -11034 13020
rect -11034 12986 -10944 13020
rect -10944 12986 -10876 13020
rect -10876 12986 -10786 13020
rect -10786 12986 -10718 13020
rect -10718 12986 -10628 13020
rect -10628 12986 -10560 13020
rect -10560 12986 -10470 13020
rect -10470 12986 -10402 13020
rect -10402 12986 -10312 13020
rect -10312 12986 -10244 13020
rect -10244 12986 -10154 13020
rect -10154 12986 -10086 13020
rect -10086 12986 -9996 13020
rect -9996 12986 -9928 13020
rect -9928 12986 -9838 13020
rect -9838 12986 -9770 13020
rect -9770 12986 -9680 13020
rect -9680 12986 -9612 13020
rect -9612 12986 -9522 13020
rect -9522 12986 -9454 13020
rect -9454 12986 -9364 13020
rect -9364 12986 -9296 13020
rect -9296 12986 -9206 13020
rect -9206 12986 -9138 13020
rect -9138 12986 -9048 13020
rect -9048 12986 -8980 13020
rect -8980 12986 -8890 13020
rect -8890 12986 -8822 13020
rect -8822 12986 -8732 13020
rect -8732 12986 -8664 13020
rect -8664 12986 -8574 13020
rect -8574 12986 -8514 13020
rect -13148 12926 -8514 12986
rect -8360 12900 -8290 13036
rect -7070 19080 -7000 19220
rect -6848 19130 -2214 19190
rect -6848 19096 -6788 19130
rect -6788 19096 -6698 19130
rect -6698 19096 -6630 19130
rect -6630 19096 -6540 19130
rect -6540 19096 -6472 19130
rect -6472 19096 -6382 19130
rect -6382 19096 -6314 19130
rect -6314 19096 -6224 19130
rect -6224 19096 -6156 19130
rect -6156 19096 -6066 19130
rect -6066 19096 -5998 19130
rect -5998 19096 -5908 19130
rect -5908 19096 -5840 19130
rect -5840 19096 -5750 19130
rect -5750 19096 -5682 19130
rect -5682 19096 -5592 19130
rect -5592 19096 -5524 19130
rect -5524 19096 -5434 19130
rect -5434 19096 -5366 19130
rect -5366 19096 -5276 19130
rect -5276 19096 -5208 19130
rect -5208 19096 -5118 19130
rect -5118 19096 -5050 19130
rect -5050 19096 -4960 19130
rect -4960 19096 -4892 19130
rect -4892 19096 -4802 19130
rect -4802 19096 -4734 19130
rect -4734 19096 -4644 19130
rect -4644 19096 -4576 19130
rect -4576 19096 -4486 19130
rect -4486 19096 -4418 19130
rect -4418 19096 -4328 19130
rect -4328 19096 -4260 19130
rect -4260 19096 -4170 19130
rect -4170 19096 -4102 19130
rect -4102 19096 -4012 19130
rect -4012 19096 -3944 19130
rect -3944 19096 -3854 19130
rect -3854 19096 -3786 19130
rect -3786 19096 -3696 19130
rect -3696 19096 -3628 19130
rect -3628 19096 -3538 19130
rect -3538 19096 -3470 19130
rect -3470 19096 -3380 19130
rect -3380 19096 -3312 19130
rect -3312 19096 -3222 19130
rect -3222 19096 -3154 19130
rect -3154 19096 -3064 19130
rect -3064 19096 -2996 19130
rect -2996 19096 -2906 19130
rect -2906 19096 -2838 19130
rect -2838 19096 -2748 19130
rect -2748 19096 -2680 19130
rect -2680 19096 -2590 19130
rect -2590 19096 -2522 19130
rect -2522 19096 -2432 19130
rect -2432 19096 -2364 19130
rect -2364 19096 -2274 19130
rect -2274 19096 -2214 19130
rect -6848 19090 -2214 19096
rect -7070 13036 -7054 19080
rect -7054 13036 -7016 19080
rect -7016 13036 -7000 19080
rect -2060 19080 -1990 19220
rect -6935 13078 -6918 19038
rect -6918 13078 -6884 19038
rect -6884 13078 -6869 19038
rect -6777 13078 -6760 19038
rect -6760 13078 -6726 19038
rect -6726 13078 -6711 19038
rect -6619 13078 -6602 19038
rect -6602 13078 -6568 19038
rect -6568 13078 -6553 19038
rect -6461 13078 -6444 19038
rect -6444 13078 -6410 19038
rect -6410 13078 -6395 19038
rect -6303 13078 -6286 19038
rect -6286 13078 -6252 19038
rect -6252 13078 -6237 19038
rect -6145 13078 -6128 19038
rect -6128 13078 -6094 19038
rect -6094 13078 -6079 19038
rect -5987 13078 -5970 19038
rect -5970 13078 -5936 19038
rect -5936 13078 -5921 19038
rect -5829 13078 -5812 19038
rect -5812 13078 -5778 19038
rect -5778 13078 -5763 19038
rect -5671 13078 -5654 19038
rect -5654 13078 -5620 19038
rect -5620 13078 -5605 19038
rect -5513 13078 -5496 19038
rect -5496 13078 -5462 19038
rect -5462 13078 -5447 19038
rect -5355 13078 -5338 19038
rect -5338 13078 -5304 19038
rect -5304 13078 -5289 19038
rect -5197 13078 -5180 19038
rect -5180 13078 -5146 19038
rect -5146 13078 -5131 19038
rect -5039 13078 -5022 19038
rect -5022 13078 -4988 19038
rect -4988 13078 -4973 19038
rect -4881 13078 -4864 19038
rect -4864 13078 -4830 19038
rect -4830 13078 -4815 19038
rect -4723 13078 -4706 19038
rect -4706 13078 -4672 19038
rect -4672 13078 -4657 19038
rect -4565 13078 -4548 19038
rect -4548 13078 -4514 19038
rect -4514 13078 -4499 19038
rect -4407 13078 -4390 19038
rect -4390 13078 -4356 19038
rect -4356 13078 -4341 19038
rect -4249 13078 -4232 19038
rect -4232 13078 -4198 19038
rect -4198 13078 -4183 19038
rect -4091 13078 -4074 19038
rect -4074 13078 -4040 19038
rect -4040 13078 -4025 19038
rect -3933 13078 -3916 19038
rect -3916 13078 -3882 19038
rect -3882 13078 -3867 19038
rect -3775 13078 -3758 19038
rect -3758 13078 -3724 19038
rect -3724 13078 -3709 19038
rect -3617 13078 -3600 19038
rect -3600 13078 -3566 19038
rect -3566 13078 -3551 19038
rect -3459 13078 -3442 19038
rect -3442 13078 -3408 19038
rect -3408 13078 -3393 19038
rect -3301 13078 -3284 19038
rect -3284 13078 -3250 19038
rect -3250 13078 -3235 19038
rect -3143 13078 -3126 19038
rect -3126 13078 -3092 19038
rect -3092 13078 -3077 19038
rect -2985 13078 -2968 19038
rect -2968 13078 -2934 19038
rect -2934 13078 -2919 19038
rect -2827 13078 -2810 19038
rect -2810 13078 -2776 19038
rect -2776 13078 -2761 19038
rect -2669 13078 -2652 19038
rect -2652 13078 -2618 19038
rect -2618 13078 -2603 19038
rect -2511 13078 -2494 19038
rect -2494 13078 -2460 19038
rect -2460 13078 -2445 19038
rect -2353 13078 -2336 19038
rect -2336 13078 -2302 19038
rect -2302 13078 -2287 19038
rect -2195 13078 -2178 19038
rect -2178 13078 -2144 19038
rect -2144 13078 -2129 19038
rect -7070 12900 -7000 13036
rect -2060 13036 -2046 19080
rect -2046 13036 -2008 19080
rect -2008 13036 -1990 19080
rect -6848 13020 -2214 13026
rect -6848 12986 -6788 13020
rect -6788 12986 -6698 13020
rect -6698 12986 -6630 13020
rect -6630 12986 -6540 13020
rect -6540 12986 -6472 13020
rect -6472 12986 -6382 13020
rect -6382 12986 -6314 13020
rect -6314 12986 -6224 13020
rect -6224 12986 -6156 13020
rect -6156 12986 -6066 13020
rect -6066 12986 -5998 13020
rect -5998 12986 -5908 13020
rect -5908 12986 -5840 13020
rect -5840 12986 -5750 13020
rect -5750 12986 -5682 13020
rect -5682 12986 -5592 13020
rect -5592 12986 -5524 13020
rect -5524 12986 -5434 13020
rect -5434 12986 -5366 13020
rect -5366 12986 -5276 13020
rect -5276 12986 -5208 13020
rect -5208 12986 -5118 13020
rect -5118 12986 -5050 13020
rect -5050 12986 -4960 13020
rect -4960 12986 -4892 13020
rect -4892 12986 -4802 13020
rect -4802 12986 -4734 13020
rect -4734 12986 -4644 13020
rect -4644 12986 -4576 13020
rect -4576 12986 -4486 13020
rect -4486 12986 -4418 13020
rect -4418 12986 -4328 13020
rect -4328 12986 -4260 13020
rect -4260 12986 -4170 13020
rect -4170 12986 -4102 13020
rect -4102 12986 -4012 13020
rect -4012 12986 -3944 13020
rect -3944 12986 -3854 13020
rect -3854 12986 -3786 13020
rect -3786 12986 -3696 13020
rect -3696 12986 -3628 13020
rect -3628 12986 -3538 13020
rect -3538 12986 -3470 13020
rect -3470 12986 -3380 13020
rect -3380 12986 -3312 13020
rect -3312 12986 -3222 13020
rect -3222 12986 -3154 13020
rect -3154 12986 -3064 13020
rect -3064 12986 -2996 13020
rect -2996 12986 -2906 13020
rect -2906 12986 -2838 13020
rect -2838 12986 -2748 13020
rect -2748 12986 -2680 13020
rect -2680 12986 -2590 13020
rect -2590 12986 -2522 13020
rect -2522 12986 -2432 13020
rect -2432 12986 -2364 13020
rect -2364 12986 -2274 13020
rect -2274 12986 -2214 13020
rect -6848 12926 -2214 12986
rect -2060 12900 -1990 13036
rect -770 19080 -700 19220
rect -548 19130 4086 19190
rect -548 19096 -488 19130
rect -488 19096 -398 19130
rect -398 19096 -330 19130
rect -330 19096 -240 19130
rect -240 19096 -172 19130
rect -172 19096 -82 19130
rect -82 19096 -14 19130
rect -14 19096 76 19130
rect 76 19096 144 19130
rect 144 19096 234 19130
rect 234 19096 302 19130
rect 302 19096 392 19130
rect 392 19096 460 19130
rect 460 19096 550 19130
rect 550 19096 618 19130
rect 618 19096 708 19130
rect 708 19096 776 19130
rect 776 19096 866 19130
rect 866 19096 934 19130
rect 934 19096 1024 19130
rect 1024 19096 1092 19130
rect 1092 19096 1182 19130
rect 1182 19096 1250 19130
rect 1250 19096 1340 19130
rect 1340 19096 1408 19130
rect 1408 19096 1498 19130
rect 1498 19096 1566 19130
rect 1566 19096 1656 19130
rect 1656 19096 1724 19130
rect 1724 19096 1814 19130
rect 1814 19096 1882 19130
rect 1882 19096 1972 19130
rect 1972 19096 2040 19130
rect 2040 19096 2130 19130
rect 2130 19096 2198 19130
rect 2198 19096 2288 19130
rect 2288 19096 2356 19130
rect 2356 19096 2446 19130
rect 2446 19096 2514 19130
rect 2514 19096 2604 19130
rect 2604 19096 2672 19130
rect 2672 19096 2762 19130
rect 2762 19096 2830 19130
rect 2830 19096 2920 19130
rect 2920 19096 2988 19130
rect 2988 19096 3078 19130
rect 3078 19096 3146 19130
rect 3146 19096 3236 19130
rect 3236 19096 3304 19130
rect 3304 19096 3394 19130
rect 3394 19096 3462 19130
rect 3462 19096 3552 19130
rect 3552 19096 3620 19130
rect 3620 19096 3710 19130
rect 3710 19096 3778 19130
rect 3778 19096 3868 19130
rect 3868 19096 3936 19130
rect 3936 19096 4026 19130
rect 4026 19096 4086 19130
rect -548 19090 4086 19096
rect -770 13036 -754 19080
rect -754 13036 -716 19080
rect -716 13036 -700 19080
rect 4240 19080 4310 19220
rect -635 13078 -618 19038
rect -618 13078 -584 19038
rect -584 13078 -569 19038
rect -477 13078 -460 19038
rect -460 13078 -426 19038
rect -426 13078 -411 19038
rect -319 13078 -302 19038
rect -302 13078 -268 19038
rect -268 13078 -253 19038
rect -161 13078 -144 19038
rect -144 13078 -110 19038
rect -110 13078 -95 19038
rect -3 13078 14 19038
rect 14 13078 48 19038
rect 48 13078 63 19038
rect 155 13078 172 19038
rect 172 13078 206 19038
rect 206 13078 221 19038
rect 313 13078 330 19038
rect 330 13078 364 19038
rect 364 13078 379 19038
rect 471 13078 488 19038
rect 488 13078 522 19038
rect 522 13078 537 19038
rect 629 13078 646 19038
rect 646 13078 680 19038
rect 680 13078 695 19038
rect 787 13078 804 19038
rect 804 13078 838 19038
rect 838 13078 853 19038
rect 945 13078 962 19038
rect 962 13078 996 19038
rect 996 13078 1011 19038
rect 1103 13078 1120 19038
rect 1120 13078 1154 19038
rect 1154 13078 1169 19038
rect 1261 13078 1278 19038
rect 1278 13078 1312 19038
rect 1312 13078 1327 19038
rect 1419 13078 1436 19038
rect 1436 13078 1470 19038
rect 1470 13078 1485 19038
rect 1577 13078 1594 19038
rect 1594 13078 1628 19038
rect 1628 13078 1643 19038
rect 1735 13078 1752 19038
rect 1752 13078 1786 19038
rect 1786 13078 1801 19038
rect 1893 13078 1910 19038
rect 1910 13078 1944 19038
rect 1944 13078 1959 19038
rect 2051 13078 2068 19038
rect 2068 13078 2102 19038
rect 2102 13078 2117 19038
rect 2209 13078 2226 19038
rect 2226 13078 2260 19038
rect 2260 13078 2275 19038
rect 2367 13078 2384 19038
rect 2384 13078 2418 19038
rect 2418 13078 2433 19038
rect 2525 13078 2542 19038
rect 2542 13078 2576 19038
rect 2576 13078 2591 19038
rect 2683 13078 2700 19038
rect 2700 13078 2734 19038
rect 2734 13078 2749 19038
rect 2841 13078 2858 19038
rect 2858 13078 2892 19038
rect 2892 13078 2907 19038
rect 2999 13078 3016 19038
rect 3016 13078 3050 19038
rect 3050 13078 3065 19038
rect 3157 13078 3174 19038
rect 3174 13078 3208 19038
rect 3208 13078 3223 19038
rect 3315 13078 3332 19038
rect 3332 13078 3366 19038
rect 3366 13078 3381 19038
rect 3473 13078 3490 19038
rect 3490 13078 3524 19038
rect 3524 13078 3539 19038
rect 3631 13078 3648 19038
rect 3648 13078 3682 19038
rect 3682 13078 3697 19038
rect 3789 13078 3806 19038
rect 3806 13078 3840 19038
rect 3840 13078 3855 19038
rect 3947 13078 3964 19038
rect 3964 13078 3998 19038
rect 3998 13078 4013 19038
rect 4105 13078 4122 19038
rect 4122 13078 4156 19038
rect 4156 13078 4171 19038
rect -770 12900 -700 13036
rect 4240 13036 4254 19080
rect 4254 13036 4292 19080
rect 4292 13036 4310 19080
rect -548 13020 4086 13026
rect -548 12986 -488 13020
rect -488 12986 -398 13020
rect -398 12986 -330 13020
rect -330 12986 -240 13020
rect -240 12986 -172 13020
rect -172 12986 -82 13020
rect -82 12986 -14 13020
rect -14 12986 76 13020
rect 76 12986 144 13020
rect 144 12986 234 13020
rect 234 12986 302 13020
rect 302 12986 392 13020
rect 392 12986 460 13020
rect 460 12986 550 13020
rect 550 12986 618 13020
rect 618 12986 708 13020
rect 708 12986 776 13020
rect 776 12986 866 13020
rect 866 12986 934 13020
rect 934 12986 1024 13020
rect 1024 12986 1092 13020
rect 1092 12986 1182 13020
rect 1182 12986 1250 13020
rect 1250 12986 1340 13020
rect 1340 12986 1408 13020
rect 1408 12986 1498 13020
rect 1498 12986 1566 13020
rect 1566 12986 1656 13020
rect 1656 12986 1724 13020
rect 1724 12986 1814 13020
rect 1814 12986 1882 13020
rect 1882 12986 1972 13020
rect 1972 12986 2040 13020
rect 2040 12986 2130 13020
rect 2130 12986 2198 13020
rect 2198 12986 2288 13020
rect 2288 12986 2356 13020
rect 2356 12986 2446 13020
rect 2446 12986 2514 13020
rect 2514 12986 2604 13020
rect 2604 12986 2672 13020
rect 2672 12986 2762 13020
rect 2762 12986 2830 13020
rect 2830 12986 2920 13020
rect 2920 12986 2988 13020
rect 2988 12986 3078 13020
rect 3078 12986 3146 13020
rect 3146 12986 3236 13020
rect 3236 12986 3304 13020
rect 3304 12986 3394 13020
rect 3394 12986 3462 13020
rect 3462 12986 3552 13020
rect 3552 12986 3620 13020
rect 3620 12986 3710 13020
rect 3710 12986 3778 13020
rect 3778 12986 3868 13020
rect 3868 12986 3936 13020
rect 3936 12986 4026 13020
rect 4026 12986 4086 13020
rect -548 12926 4086 12986
rect 4240 12900 4310 13036
rect 5530 19080 5600 19220
rect 5752 19130 10386 19190
rect 5752 19096 5812 19130
rect 5812 19096 5902 19130
rect 5902 19096 5970 19130
rect 5970 19096 6060 19130
rect 6060 19096 6128 19130
rect 6128 19096 6218 19130
rect 6218 19096 6286 19130
rect 6286 19096 6376 19130
rect 6376 19096 6444 19130
rect 6444 19096 6534 19130
rect 6534 19096 6602 19130
rect 6602 19096 6692 19130
rect 6692 19096 6760 19130
rect 6760 19096 6850 19130
rect 6850 19096 6918 19130
rect 6918 19096 7008 19130
rect 7008 19096 7076 19130
rect 7076 19096 7166 19130
rect 7166 19096 7234 19130
rect 7234 19096 7324 19130
rect 7324 19096 7392 19130
rect 7392 19096 7482 19130
rect 7482 19096 7550 19130
rect 7550 19096 7640 19130
rect 7640 19096 7708 19130
rect 7708 19096 7798 19130
rect 7798 19096 7866 19130
rect 7866 19096 7956 19130
rect 7956 19096 8024 19130
rect 8024 19096 8114 19130
rect 8114 19096 8182 19130
rect 8182 19096 8272 19130
rect 8272 19096 8340 19130
rect 8340 19096 8430 19130
rect 8430 19096 8498 19130
rect 8498 19096 8588 19130
rect 8588 19096 8656 19130
rect 8656 19096 8746 19130
rect 8746 19096 8814 19130
rect 8814 19096 8904 19130
rect 8904 19096 8972 19130
rect 8972 19096 9062 19130
rect 9062 19096 9130 19130
rect 9130 19096 9220 19130
rect 9220 19096 9288 19130
rect 9288 19096 9378 19130
rect 9378 19096 9446 19130
rect 9446 19096 9536 19130
rect 9536 19096 9604 19130
rect 9604 19096 9694 19130
rect 9694 19096 9762 19130
rect 9762 19096 9852 19130
rect 9852 19096 9920 19130
rect 9920 19096 10010 19130
rect 10010 19096 10078 19130
rect 10078 19096 10168 19130
rect 10168 19096 10236 19130
rect 10236 19096 10326 19130
rect 10326 19096 10386 19130
rect 5752 19090 10386 19096
rect 5530 13036 5546 19080
rect 5546 13036 5584 19080
rect 5584 13036 5600 19080
rect 10540 19080 10610 19220
rect 5665 13078 5682 19038
rect 5682 13078 5716 19038
rect 5716 13078 5731 19038
rect 5823 13078 5840 19038
rect 5840 13078 5874 19038
rect 5874 13078 5889 19038
rect 5981 13078 5998 19038
rect 5998 13078 6032 19038
rect 6032 13078 6047 19038
rect 6139 13078 6156 19038
rect 6156 13078 6190 19038
rect 6190 13078 6205 19038
rect 6297 13078 6314 19038
rect 6314 13078 6348 19038
rect 6348 13078 6363 19038
rect 6455 13078 6472 19038
rect 6472 13078 6506 19038
rect 6506 13078 6521 19038
rect 6613 13078 6630 19038
rect 6630 13078 6664 19038
rect 6664 13078 6679 19038
rect 6771 13078 6788 19038
rect 6788 13078 6822 19038
rect 6822 13078 6837 19038
rect 6929 13078 6946 19038
rect 6946 13078 6980 19038
rect 6980 13078 6995 19038
rect 7087 13078 7104 19038
rect 7104 13078 7138 19038
rect 7138 13078 7153 19038
rect 7245 13078 7262 19038
rect 7262 13078 7296 19038
rect 7296 13078 7311 19038
rect 7403 13078 7420 19038
rect 7420 13078 7454 19038
rect 7454 13078 7469 19038
rect 7561 13078 7578 19038
rect 7578 13078 7612 19038
rect 7612 13078 7627 19038
rect 7719 13078 7736 19038
rect 7736 13078 7770 19038
rect 7770 13078 7785 19038
rect 7877 13078 7894 19038
rect 7894 13078 7928 19038
rect 7928 13078 7943 19038
rect 8035 13078 8052 19038
rect 8052 13078 8086 19038
rect 8086 13078 8101 19038
rect 8193 13078 8210 19038
rect 8210 13078 8244 19038
rect 8244 13078 8259 19038
rect 8351 13078 8368 19038
rect 8368 13078 8402 19038
rect 8402 13078 8417 19038
rect 8509 13078 8526 19038
rect 8526 13078 8560 19038
rect 8560 13078 8575 19038
rect 8667 13078 8684 19038
rect 8684 13078 8718 19038
rect 8718 13078 8733 19038
rect 8825 13078 8842 19038
rect 8842 13078 8876 19038
rect 8876 13078 8891 19038
rect 8983 13078 9000 19038
rect 9000 13078 9034 19038
rect 9034 13078 9049 19038
rect 9141 13078 9158 19038
rect 9158 13078 9192 19038
rect 9192 13078 9207 19038
rect 9299 13078 9316 19038
rect 9316 13078 9350 19038
rect 9350 13078 9365 19038
rect 9457 13078 9474 19038
rect 9474 13078 9508 19038
rect 9508 13078 9523 19038
rect 9615 13078 9632 19038
rect 9632 13078 9666 19038
rect 9666 13078 9681 19038
rect 9773 13078 9790 19038
rect 9790 13078 9824 19038
rect 9824 13078 9839 19038
rect 9931 13078 9948 19038
rect 9948 13078 9982 19038
rect 9982 13078 9997 19038
rect 10089 13078 10106 19038
rect 10106 13078 10140 19038
rect 10140 13078 10155 19038
rect 10247 13078 10264 19038
rect 10264 13078 10298 19038
rect 10298 13078 10313 19038
rect 10405 13078 10422 19038
rect 10422 13078 10456 19038
rect 10456 13078 10471 19038
rect 5530 12900 5600 13036
rect 10540 13036 10554 19080
rect 10554 13036 10592 19080
rect 10592 13036 10610 19080
rect 5752 13020 10386 13026
rect 5752 12986 5812 13020
rect 5812 12986 5902 13020
rect 5902 12986 5970 13020
rect 5970 12986 6060 13020
rect 6060 12986 6128 13020
rect 6128 12986 6218 13020
rect 6218 12986 6286 13020
rect 6286 12986 6376 13020
rect 6376 12986 6444 13020
rect 6444 12986 6534 13020
rect 6534 12986 6602 13020
rect 6602 12986 6692 13020
rect 6692 12986 6760 13020
rect 6760 12986 6850 13020
rect 6850 12986 6918 13020
rect 6918 12986 7008 13020
rect 7008 12986 7076 13020
rect 7076 12986 7166 13020
rect 7166 12986 7234 13020
rect 7234 12986 7324 13020
rect 7324 12986 7392 13020
rect 7392 12986 7482 13020
rect 7482 12986 7550 13020
rect 7550 12986 7640 13020
rect 7640 12986 7708 13020
rect 7708 12986 7798 13020
rect 7798 12986 7866 13020
rect 7866 12986 7956 13020
rect 7956 12986 8024 13020
rect 8024 12986 8114 13020
rect 8114 12986 8182 13020
rect 8182 12986 8272 13020
rect 8272 12986 8340 13020
rect 8340 12986 8430 13020
rect 8430 12986 8498 13020
rect 8498 12986 8588 13020
rect 8588 12986 8656 13020
rect 8656 12986 8746 13020
rect 8746 12986 8814 13020
rect 8814 12986 8904 13020
rect 8904 12986 8972 13020
rect 8972 12986 9062 13020
rect 9062 12986 9130 13020
rect 9130 12986 9220 13020
rect 9220 12986 9288 13020
rect 9288 12986 9378 13020
rect 9378 12986 9446 13020
rect 9446 12986 9536 13020
rect 9536 12986 9604 13020
rect 9604 12986 9694 13020
rect 9694 12986 9762 13020
rect 9762 12986 9852 13020
rect 9852 12986 9920 13020
rect 9920 12986 10010 13020
rect 10010 12986 10078 13020
rect 10078 12986 10168 13020
rect 10168 12986 10236 13020
rect 10236 12986 10326 13020
rect 10326 12986 10386 13020
rect 5752 12926 10386 12986
rect 10540 12900 10610 13036
rect -13370 12080 -13300 12220
rect -13148 12130 -8514 12190
rect -13148 12096 -13088 12130
rect -13088 12096 -12998 12130
rect -12998 12096 -12930 12130
rect -12930 12096 -12840 12130
rect -12840 12096 -12772 12130
rect -12772 12096 -12682 12130
rect -12682 12096 -12614 12130
rect -12614 12096 -12524 12130
rect -12524 12096 -12456 12130
rect -12456 12096 -12366 12130
rect -12366 12096 -12298 12130
rect -12298 12096 -12208 12130
rect -12208 12096 -12140 12130
rect -12140 12096 -12050 12130
rect -12050 12096 -11982 12130
rect -11982 12096 -11892 12130
rect -11892 12096 -11824 12130
rect -11824 12096 -11734 12130
rect -11734 12096 -11666 12130
rect -11666 12096 -11576 12130
rect -11576 12096 -11508 12130
rect -11508 12096 -11418 12130
rect -11418 12096 -11350 12130
rect -11350 12096 -11260 12130
rect -11260 12096 -11192 12130
rect -11192 12096 -11102 12130
rect -11102 12096 -11034 12130
rect -11034 12096 -10944 12130
rect -10944 12096 -10876 12130
rect -10876 12096 -10786 12130
rect -10786 12096 -10718 12130
rect -10718 12096 -10628 12130
rect -10628 12096 -10560 12130
rect -10560 12096 -10470 12130
rect -10470 12096 -10402 12130
rect -10402 12096 -10312 12130
rect -10312 12096 -10244 12130
rect -10244 12096 -10154 12130
rect -10154 12096 -10086 12130
rect -10086 12096 -9996 12130
rect -9996 12096 -9928 12130
rect -9928 12096 -9838 12130
rect -9838 12096 -9770 12130
rect -9770 12096 -9680 12130
rect -9680 12096 -9612 12130
rect -9612 12096 -9522 12130
rect -9522 12096 -9454 12130
rect -9454 12096 -9364 12130
rect -9364 12096 -9296 12130
rect -9296 12096 -9206 12130
rect -9206 12096 -9138 12130
rect -9138 12096 -9048 12130
rect -9048 12096 -8980 12130
rect -8980 12096 -8890 12130
rect -8890 12096 -8822 12130
rect -8822 12096 -8732 12130
rect -8732 12096 -8664 12130
rect -8664 12096 -8574 12130
rect -8574 12096 -8514 12130
rect -13148 12090 -8514 12096
rect -13370 6036 -13354 12080
rect -13354 6036 -13316 12080
rect -13316 6036 -13300 12080
rect -8360 12080 -8290 12220
rect -13235 6078 -13218 12038
rect -13218 6078 -13184 12038
rect -13184 6078 -13169 12038
rect -13077 6078 -13060 12038
rect -13060 6078 -13026 12038
rect -13026 6078 -13011 12038
rect -12919 6078 -12902 12038
rect -12902 6078 -12868 12038
rect -12868 6078 -12853 12038
rect -12761 6078 -12744 12038
rect -12744 6078 -12710 12038
rect -12710 6078 -12695 12038
rect -12603 6078 -12586 12038
rect -12586 6078 -12552 12038
rect -12552 6078 -12537 12038
rect -12445 6078 -12428 12038
rect -12428 6078 -12394 12038
rect -12394 6078 -12379 12038
rect -12287 6078 -12270 12038
rect -12270 6078 -12236 12038
rect -12236 6078 -12221 12038
rect -12129 6078 -12112 12038
rect -12112 6078 -12078 12038
rect -12078 6078 -12063 12038
rect -11971 6078 -11954 12038
rect -11954 6078 -11920 12038
rect -11920 6078 -11905 12038
rect -11813 6078 -11796 12038
rect -11796 6078 -11762 12038
rect -11762 6078 -11747 12038
rect -11655 6078 -11638 12038
rect -11638 6078 -11604 12038
rect -11604 6078 -11589 12038
rect -11497 6078 -11480 12038
rect -11480 6078 -11446 12038
rect -11446 6078 -11431 12038
rect -11339 6078 -11322 12038
rect -11322 6078 -11288 12038
rect -11288 6078 -11273 12038
rect -11181 6078 -11164 12038
rect -11164 6078 -11130 12038
rect -11130 6078 -11115 12038
rect -11023 6078 -11006 12038
rect -11006 6078 -10972 12038
rect -10972 6078 -10957 12038
rect -10865 6078 -10848 12038
rect -10848 6078 -10814 12038
rect -10814 6078 -10799 12038
rect -10707 6078 -10690 12038
rect -10690 6078 -10656 12038
rect -10656 6078 -10641 12038
rect -10549 6078 -10532 12038
rect -10532 6078 -10498 12038
rect -10498 6078 -10483 12038
rect -10391 6078 -10374 12038
rect -10374 6078 -10340 12038
rect -10340 6078 -10325 12038
rect -10233 6078 -10216 12038
rect -10216 6078 -10182 12038
rect -10182 6078 -10167 12038
rect -10075 6078 -10058 12038
rect -10058 6078 -10024 12038
rect -10024 6078 -10009 12038
rect -9917 6078 -9900 12038
rect -9900 6078 -9866 12038
rect -9866 6078 -9851 12038
rect -9759 6078 -9742 12038
rect -9742 6078 -9708 12038
rect -9708 6078 -9693 12038
rect -9601 6078 -9584 12038
rect -9584 6078 -9550 12038
rect -9550 6078 -9535 12038
rect -9443 6078 -9426 12038
rect -9426 6078 -9392 12038
rect -9392 6078 -9377 12038
rect -9285 6078 -9268 12038
rect -9268 6078 -9234 12038
rect -9234 6078 -9219 12038
rect -9127 6078 -9110 12038
rect -9110 6078 -9076 12038
rect -9076 6078 -9061 12038
rect -8969 6078 -8952 12038
rect -8952 6078 -8918 12038
rect -8918 6078 -8903 12038
rect -8811 6078 -8794 12038
rect -8794 6078 -8760 12038
rect -8760 6078 -8745 12038
rect -8653 6078 -8636 12038
rect -8636 6078 -8602 12038
rect -8602 6078 -8587 12038
rect -8495 6078 -8478 12038
rect -8478 6078 -8444 12038
rect -8444 6078 -8429 12038
rect -13370 5900 -13300 6036
rect -8360 6036 -8346 12080
rect -8346 6036 -8308 12080
rect -8308 6036 -8290 12080
rect -13148 6020 -8514 6026
rect -13148 5986 -13088 6020
rect -13088 5986 -12998 6020
rect -12998 5986 -12930 6020
rect -12930 5986 -12840 6020
rect -12840 5986 -12772 6020
rect -12772 5986 -12682 6020
rect -12682 5986 -12614 6020
rect -12614 5986 -12524 6020
rect -12524 5986 -12456 6020
rect -12456 5986 -12366 6020
rect -12366 5986 -12298 6020
rect -12298 5986 -12208 6020
rect -12208 5986 -12140 6020
rect -12140 5986 -12050 6020
rect -12050 5986 -11982 6020
rect -11982 5986 -11892 6020
rect -11892 5986 -11824 6020
rect -11824 5986 -11734 6020
rect -11734 5986 -11666 6020
rect -11666 5986 -11576 6020
rect -11576 5986 -11508 6020
rect -11508 5986 -11418 6020
rect -11418 5986 -11350 6020
rect -11350 5986 -11260 6020
rect -11260 5986 -11192 6020
rect -11192 5986 -11102 6020
rect -11102 5986 -11034 6020
rect -11034 5986 -10944 6020
rect -10944 5986 -10876 6020
rect -10876 5986 -10786 6020
rect -10786 5986 -10718 6020
rect -10718 5986 -10628 6020
rect -10628 5986 -10560 6020
rect -10560 5986 -10470 6020
rect -10470 5986 -10402 6020
rect -10402 5986 -10312 6020
rect -10312 5986 -10244 6020
rect -10244 5986 -10154 6020
rect -10154 5986 -10086 6020
rect -10086 5986 -9996 6020
rect -9996 5986 -9928 6020
rect -9928 5986 -9838 6020
rect -9838 5986 -9770 6020
rect -9770 5986 -9680 6020
rect -9680 5986 -9612 6020
rect -9612 5986 -9522 6020
rect -9522 5986 -9454 6020
rect -9454 5986 -9364 6020
rect -9364 5986 -9296 6020
rect -9296 5986 -9206 6020
rect -9206 5986 -9138 6020
rect -9138 5986 -9048 6020
rect -9048 5986 -8980 6020
rect -8980 5986 -8890 6020
rect -8890 5986 -8822 6020
rect -8822 5986 -8732 6020
rect -8732 5986 -8664 6020
rect -8664 5986 -8574 6020
rect -8574 5986 -8514 6020
rect -13148 5926 -8514 5986
rect -8360 5900 -8290 6036
rect -7070 12080 -7000 12220
rect -6848 12130 -2214 12190
rect -6848 12096 -6788 12130
rect -6788 12096 -6698 12130
rect -6698 12096 -6630 12130
rect -6630 12096 -6540 12130
rect -6540 12096 -6472 12130
rect -6472 12096 -6382 12130
rect -6382 12096 -6314 12130
rect -6314 12096 -6224 12130
rect -6224 12096 -6156 12130
rect -6156 12096 -6066 12130
rect -6066 12096 -5998 12130
rect -5998 12096 -5908 12130
rect -5908 12096 -5840 12130
rect -5840 12096 -5750 12130
rect -5750 12096 -5682 12130
rect -5682 12096 -5592 12130
rect -5592 12096 -5524 12130
rect -5524 12096 -5434 12130
rect -5434 12096 -5366 12130
rect -5366 12096 -5276 12130
rect -5276 12096 -5208 12130
rect -5208 12096 -5118 12130
rect -5118 12096 -5050 12130
rect -5050 12096 -4960 12130
rect -4960 12096 -4892 12130
rect -4892 12096 -4802 12130
rect -4802 12096 -4734 12130
rect -4734 12096 -4644 12130
rect -4644 12096 -4576 12130
rect -4576 12096 -4486 12130
rect -4486 12096 -4418 12130
rect -4418 12096 -4328 12130
rect -4328 12096 -4260 12130
rect -4260 12096 -4170 12130
rect -4170 12096 -4102 12130
rect -4102 12096 -4012 12130
rect -4012 12096 -3944 12130
rect -3944 12096 -3854 12130
rect -3854 12096 -3786 12130
rect -3786 12096 -3696 12130
rect -3696 12096 -3628 12130
rect -3628 12096 -3538 12130
rect -3538 12096 -3470 12130
rect -3470 12096 -3380 12130
rect -3380 12096 -3312 12130
rect -3312 12096 -3222 12130
rect -3222 12096 -3154 12130
rect -3154 12096 -3064 12130
rect -3064 12096 -2996 12130
rect -2996 12096 -2906 12130
rect -2906 12096 -2838 12130
rect -2838 12096 -2748 12130
rect -2748 12096 -2680 12130
rect -2680 12096 -2590 12130
rect -2590 12096 -2522 12130
rect -2522 12096 -2432 12130
rect -2432 12096 -2364 12130
rect -2364 12096 -2274 12130
rect -2274 12096 -2214 12130
rect -6848 12090 -2214 12096
rect -7070 6036 -7054 12080
rect -7054 6036 -7016 12080
rect -7016 6036 -7000 12080
rect -2060 12080 -1990 12220
rect -6935 6078 -6918 12038
rect -6918 6078 -6884 12038
rect -6884 6078 -6869 12038
rect -6777 6078 -6760 12038
rect -6760 6078 -6726 12038
rect -6726 6078 -6711 12038
rect -6619 6078 -6602 12038
rect -6602 6078 -6568 12038
rect -6568 6078 -6553 12038
rect -6461 6078 -6444 12038
rect -6444 6078 -6410 12038
rect -6410 6078 -6395 12038
rect -6303 6078 -6286 12038
rect -6286 6078 -6252 12038
rect -6252 6078 -6237 12038
rect -6145 6078 -6128 12038
rect -6128 6078 -6094 12038
rect -6094 6078 -6079 12038
rect -5987 6078 -5970 12038
rect -5970 6078 -5936 12038
rect -5936 6078 -5921 12038
rect -5829 6078 -5812 12038
rect -5812 6078 -5778 12038
rect -5778 6078 -5763 12038
rect -5671 6078 -5654 12038
rect -5654 6078 -5620 12038
rect -5620 6078 -5605 12038
rect -5513 6078 -5496 12038
rect -5496 6078 -5462 12038
rect -5462 6078 -5447 12038
rect -5355 6078 -5338 12038
rect -5338 6078 -5304 12038
rect -5304 6078 -5289 12038
rect -5197 6078 -5180 12038
rect -5180 6078 -5146 12038
rect -5146 6078 -5131 12038
rect -5039 6078 -5022 12038
rect -5022 6078 -4988 12038
rect -4988 6078 -4973 12038
rect -4881 6078 -4864 12038
rect -4864 6078 -4830 12038
rect -4830 6078 -4815 12038
rect -4723 6078 -4706 12038
rect -4706 6078 -4672 12038
rect -4672 6078 -4657 12038
rect -4565 6078 -4548 12038
rect -4548 6078 -4514 12038
rect -4514 6078 -4499 12038
rect -4407 6078 -4390 12038
rect -4390 6078 -4356 12038
rect -4356 6078 -4341 12038
rect -4249 6078 -4232 12038
rect -4232 6078 -4198 12038
rect -4198 6078 -4183 12038
rect -4091 6078 -4074 12038
rect -4074 6078 -4040 12038
rect -4040 6078 -4025 12038
rect -3933 6078 -3916 12038
rect -3916 6078 -3882 12038
rect -3882 6078 -3867 12038
rect -3775 6078 -3758 12038
rect -3758 6078 -3724 12038
rect -3724 6078 -3709 12038
rect -3617 6078 -3600 12038
rect -3600 6078 -3566 12038
rect -3566 6078 -3551 12038
rect -3459 6078 -3442 12038
rect -3442 6078 -3408 12038
rect -3408 6078 -3393 12038
rect -3301 6078 -3284 12038
rect -3284 6078 -3250 12038
rect -3250 6078 -3235 12038
rect -3143 6078 -3126 12038
rect -3126 6078 -3092 12038
rect -3092 6078 -3077 12038
rect -2985 6078 -2968 12038
rect -2968 6078 -2934 12038
rect -2934 6078 -2919 12038
rect -2827 6078 -2810 12038
rect -2810 6078 -2776 12038
rect -2776 6078 -2761 12038
rect -2669 6078 -2652 12038
rect -2652 6078 -2618 12038
rect -2618 6078 -2603 12038
rect -2511 6078 -2494 12038
rect -2494 6078 -2460 12038
rect -2460 6078 -2445 12038
rect -2353 6078 -2336 12038
rect -2336 6078 -2302 12038
rect -2302 6078 -2287 12038
rect -2195 6078 -2178 12038
rect -2178 6078 -2144 12038
rect -2144 6078 -2129 12038
rect -7070 5900 -7000 6036
rect -2060 6036 -2046 12080
rect -2046 6036 -2008 12080
rect -2008 6036 -1990 12080
rect -6848 6020 -2214 6026
rect -6848 5986 -6788 6020
rect -6788 5986 -6698 6020
rect -6698 5986 -6630 6020
rect -6630 5986 -6540 6020
rect -6540 5986 -6472 6020
rect -6472 5986 -6382 6020
rect -6382 5986 -6314 6020
rect -6314 5986 -6224 6020
rect -6224 5986 -6156 6020
rect -6156 5986 -6066 6020
rect -6066 5986 -5998 6020
rect -5998 5986 -5908 6020
rect -5908 5986 -5840 6020
rect -5840 5986 -5750 6020
rect -5750 5986 -5682 6020
rect -5682 5986 -5592 6020
rect -5592 5986 -5524 6020
rect -5524 5986 -5434 6020
rect -5434 5986 -5366 6020
rect -5366 5986 -5276 6020
rect -5276 5986 -5208 6020
rect -5208 5986 -5118 6020
rect -5118 5986 -5050 6020
rect -5050 5986 -4960 6020
rect -4960 5986 -4892 6020
rect -4892 5986 -4802 6020
rect -4802 5986 -4734 6020
rect -4734 5986 -4644 6020
rect -4644 5986 -4576 6020
rect -4576 5986 -4486 6020
rect -4486 5986 -4418 6020
rect -4418 5986 -4328 6020
rect -4328 5986 -4260 6020
rect -4260 5986 -4170 6020
rect -4170 5986 -4102 6020
rect -4102 5986 -4012 6020
rect -4012 5986 -3944 6020
rect -3944 5986 -3854 6020
rect -3854 5986 -3786 6020
rect -3786 5986 -3696 6020
rect -3696 5986 -3628 6020
rect -3628 5986 -3538 6020
rect -3538 5986 -3470 6020
rect -3470 5986 -3380 6020
rect -3380 5986 -3312 6020
rect -3312 5986 -3222 6020
rect -3222 5986 -3154 6020
rect -3154 5986 -3064 6020
rect -3064 5986 -2996 6020
rect -2996 5986 -2906 6020
rect -2906 5986 -2838 6020
rect -2838 5986 -2748 6020
rect -2748 5986 -2680 6020
rect -2680 5986 -2590 6020
rect -2590 5986 -2522 6020
rect -2522 5986 -2432 6020
rect -2432 5986 -2364 6020
rect -2364 5986 -2274 6020
rect -2274 5986 -2214 6020
rect -6848 5926 -2214 5986
rect -2060 5900 -1990 6036
rect -770 12080 -700 12220
rect -548 12130 4086 12190
rect -548 12096 -488 12130
rect -488 12096 -398 12130
rect -398 12096 -330 12130
rect -330 12096 -240 12130
rect -240 12096 -172 12130
rect -172 12096 -82 12130
rect -82 12096 -14 12130
rect -14 12096 76 12130
rect 76 12096 144 12130
rect 144 12096 234 12130
rect 234 12096 302 12130
rect 302 12096 392 12130
rect 392 12096 460 12130
rect 460 12096 550 12130
rect 550 12096 618 12130
rect 618 12096 708 12130
rect 708 12096 776 12130
rect 776 12096 866 12130
rect 866 12096 934 12130
rect 934 12096 1024 12130
rect 1024 12096 1092 12130
rect 1092 12096 1182 12130
rect 1182 12096 1250 12130
rect 1250 12096 1340 12130
rect 1340 12096 1408 12130
rect 1408 12096 1498 12130
rect 1498 12096 1566 12130
rect 1566 12096 1656 12130
rect 1656 12096 1724 12130
rect 1724 12096 1814 12130
rect 1814 12096 1882 12130
rect 1882 12096 1972 12130
rect 1972 12096 2040 12130
rect 2040 12096 2130 12130
rect 2130 12096 2198 12130
rect 2198 12096 2288 12130
rect 2288 12096 2356 12130
rect 2356 12096 2446 12130
rect 2446 12096 2514 12130
rect 2514 12096 2604 12130
rect 2604 12096 2672 12130
rect 2672 12096 2762 12130
rect 2762 12096 2830 12130
rect 2830 12096 2920 12130
rect 2920 12096 2988 12130
rect 2988 12096 3078 12130
rect 3078 12096 3146 12130
rect 3146 12096 3236 12130
rect 3236 12096 3304 12130
rect 3304 12096 3394 12130
rect 3394 12096 3462 12130
rect 3462 12096 3552 12130
rect 3552 12096 3620 12130
rect 3620 12096 3710 12130
rect 3710 12096 3778 12130
rect 3778 12096 3868 12130
rect 3868 12096 3936 12130
rect 3936 12096 4026 12130
rect 4026 12096 4086 12130
rect -548 12090 4086 12096
rect -770 6036 -754 12080
rect -754 6036 -716 12080
rect -716 6036 -700 12080
rect 4240 12080 4310 12220
rect -635 6078 -618 12038
rect -618 6078 -584 12038
rect -584 6078 -569 12038
rect -477 6078 -460 12038
rect -460 6078 -426 12038
rect -426 6078 -411 12038
rect -319 6078 -302 12038
rect -302 6078 -268 12038
rect -268 6078 -253 12038
rect -161 6078 -144 12038
rect -144 6078 -110 12038
rect -110 6078 -95 12038
rect -3 6078 14 12038
rect 14 6078 48 12038
rect 48 6078 63 12038
rect 155 6078 172 12038
rect 172 6078 206 12038
rect 206 6078 221 12038
rect 313 6078 330 12038
rect 330 6078 364 12038
rect 364 6078 379 12038
rect 471 6078 488 12038
rect 488 6078 522 12038
rect 522 6078 537 12038
rect 629 6078 646 12038
rect 646 6078 680 12038
rect 680 6078 695 12038
rect 787 6078 804 12038
rect 804 6078 838 12038
rect 838 6078 853 12038
rect 945 6078 962 12038
rect 962 6078 996 12038
rect 996 6078 1011 12038
rect 1103 6078 1120 12038
rect 1120 6078 1154 12038
rect 1154 6078 1169 12038
rect 1261 6078 1278 12038
rect 1278 6078 1312 12038
rect 1312 6078 1327 12038
rect 1419 6078 1436 12038
rect 1436 6078 1470 12038
rect 1470 6078 1485 12038
rect 1577 6078 1594 12038
rect 1594 6078 1628 12038
rect 1628 6078 1643 12038
rect 1735 6078 1752 12038
rect 1752 6078 1786 12038
rect 1786 6078 1801 12038
rect 1893 6078 1910 12038
rect 1910 6078 1944 12038
rect 1944 6078 1959 12038
rect 2051 6078 2068 12038
rect 2068 6078 2102 12038
rect 2102 6078 2117 12038
rect 2209 6078 2226 12038
rect 2226 6078 2260 12038
rect 2260 6078 2275 12038
rect 2367 6078 2384 12038
rect 2384 6078 2418 12038
rect 2418 6078 2433 12038
rect 2525 6078 2542 12038
rect 2542 6078 2576 12038
rect 2576 6078 2591 12038
rect 2683 6078 2700 12038
rect 2700 6078 2734 12038
rect 2734 6078 2749 12038
rect 2841 6078 2858 12038
rect 2858 6078 2892 12038
rect 2892 6078 2907 12038
rect 2999 6078 3016 12038
rect 3016 6078 3050 12038
rect 3050 6078 3065 12038
rect 3157 6078 3174 12038
rect 3174 6078 3208 12038
rect 3208 6078 3223 12038
rect 3315 6078 3332 12038
rect 3332 6078 3366 12038
rect 3366 6078 3381 12038
rect 3473 6078 3490 12038
rect 3490 6078 3524 12038
rect 3524 6078 3539 12038
rect 3631 6078 3648 12038
rect 3648 6078 3682 12038
rect 3682 6078 3697 12038
rect 3789 6078 3806 12038
rect 3806 6078 3840 12038
rect 3840 6078 3855 12038
rect 3947 6078 3964 12038
rect 3964 6078 3998 12038
rect 3998 6078 4013 12038
rect 4105 6078 4122 12038
rect 4122 6078 4156 12038
rect 4156 6078 4171 12038
rect -770 5900 -700 6036
rect 4240 6036 4254 12080
rect 4254 6036 4292 12080
rect 4292 6036 4310 12080
rect -548 6020 4086 6026
rect -548 5986 -488 6020
rect -488 5986 -398 6020
rect -398 5986 -330 6020
rect -330 5986 -240 6020
rect -240 5986 -172 6020
rect -172 5986 -82 6020
rect -82 5986 -14 6020
rect -14 5986 76 6020
rect 76 5986 144 6020
rect 144 5986 234 6020
rect 234 5986 302 6020
rect 302 5986 392 6020
rect 392 5986 460 6020
rect 460 5986 550 6020
rect 550 5986 618 6020
rect 618 5986 708 6020
rect 708 5986 776 6020
rect 776 5986 866 6020
rect 866 5986 934 6020
rect 934 5986 1024 6020
rect 1024 5986 1092 6020
rect 1092 5986 1182 6020
rect 1182 5986 1250 6020
rect 1250 5986 1340 6020
rect 1340 5986 1408 6020
rect 1408 5986 1498 6020
rect 1498 5986 1566 6020
rect 1566 5986 1656 6020
rect 1656 5986 1724 6020
rect 1724 5986 1814 6020
rect 1814 5986 1882 6020
rect 1882 5986 1972 6020
rect 1972 5986 2040 6020
rect 2040 5986 2130 6020
rect 2130 5986 2198 6020
rect 2198 5986 2288 6020
rect 2288 5986 2356 6020
rect 2356 5986 2446 6020
rect 2446 5986 2514 6020
rect 2514 5986 2604 6020
rect 2604 5986 2672 6020
rect 2672 5986 2762 6020
rect 2762 5986 2830 6020
rect 2830 5986 2920 6020
rect 2920 5986 2988 6020
rect 2988 5986 3078 6020
rect 3078 5986 3146 6020
rect 3146 5986 3236 6020
rect 3236 5986 3304 6020
rect 3304 5986 3394 6020
rect 3394 5986 3462 6020
rect 3462 5986 3552 6020
rect 3552 5986 3620 6020
rect 3620 5986 3710 6020
rect 3710 5986 3778 6020
rect 3778 5986 3868 6020
rect 3868 5986 3936 6020
rect 3936 5986 4026 6020
rect 4026 5986 4086 6020
rect -548 5926 4086 5986
rect 4240 5900 4310 6036
rect 5530 12080 5600 12220
rect 5752 12130 10386 12190
rect 5752 12096 5812 12130
rect 5812 12096 5902 12130
rect 5902 12096 5970 12130
rect 5970 12096 6060 12130
rect 6060 12096 6128 12130
rect 6128 12096 6218 12130
rect 6218 12096 6286 12130
rect 6286 12096 6376 12130
rect 6376 12096 6444 12130
rect 6444 12096 6534 12130
rect 6534 12096 6602 12130
rect 6602 12096 6692 12130
rect 6692 12096 6760 12130
rect 6760 12096 6850 12130
rect 6850 12096 6918 12130
rect 6918 12096 7008 12130
rect 7008 12096 7076 12130
rect 7076 12096 7166 12130
rect 7166 12096 7234 12130
rect 7234 12096 7324 12130
rect 7324 12096 7392 12130
rect 7392 12096 7482 12130
rect 7482 12096 7550 12130
rect 7550 12096 7640 12130
rect 7640 12096 7708 12130
rect 7708 12096 7798 12130
rect 7798 12096 7866 12130
rect 7866 12096 7956 12130
rect 7956 12096 8024 12130
rect 8024 12096 8114 12130
rect 8114 12096 8182 12130
rect 8182 12096 8272 12130
rect 8272 12096 8340 12130
rect 8340 12096 8430 12130
rect 8430 12096 8498 12130
rect 8498 12096 8588 12130
rect 8588 12096 8656 12130
rect 8656 12096 8746 12130
rect 8746 12096 8814 12130
rect 8814 12096 8904 12130
rect 8904 12096 8972 12130
rect 8972 12096 9062 12130
rect 9062 12096 9130 12130
rect 9130 12096 9220 12130
rect 9220 12096 9288 12130
rect 9288 12096 9378 12130
rect 9378 12096 9446 12130
rect 9446 12096 9536 12130
rect 9536 12096 9604 12130
rect 9604 12096 9694 12130
rect 9694 12096 9762 12130
rect 9762 12096 9852 12130
rect 9852 12096 9920 12130
rect 9920 12096 10010 12130
rect 10010 12096 10078 12130
rect 10078 12096 10168 12130
rect 10168 12096 10236 12130
rect 10236 12096 10326 12130
rect 10326 12096 10386 12130
rect 5752 12090 10386 12096
rect 5530 6036 5546 12080
rect 5546 6036 5584 12080
rect 5584 6036 5600 12080
rect 10540 12080 10610 12220
rect 5665 6078 5682 12038
rect 5682 6078 5716 12038
rect 5716 6078 5731 12038
rect 5823 6078 5840 12038
rect 5840 6078 5874 12038
rect 5874 6078 5889 12038
rect 5981 6078 5998 12038
rect 5998 6078 6032 12038
rect 6032 6078 6047 12038
rect 6139 6078 6156 12038
rect 6156 6078 6190 12038
rect 6190 6078 6205 12038
rect 6297 6078 6314 12038
rect 6314 6078 6348 12038
rect 6348 6078 6363 12038
rect 6455 6078 6472 12038
rect 6472 6078 6506 12038
rect 6506 6078 6521 12038
rect 6613 6078 6630 12038
rect 6630 6078 6664 12038
rect 6664 6078 6679 12038
rect 6771 6078 6788 12038
rect 6788 6078 6822 12038
rect 6822 6078 6837 12038
rect 6929 6078 6946 12038
rect 6946 6078 6980 12038
rect 6980 6078 6995 12038
rect 7087 6078 7104 12038
rect 7104 6078 7138 12038
rect 7138 6078 7153 12038
rect 7245 6078 7262 12038
rect 7262 6078 7296 12038
rect 7296 6078 7311 12038
rect 7403 6078 7420 12038
rect 7420 6078 7454 12038
rect 7454 6078 7469 12038
rect 7561 6078 7578 12038
rect 7578 6078 7612 12038
rect 7612 6078 7627 12038
rect 7719 6078 7736 12038
rect 7736 6078 7770 12038
rect 7770 6078 7785 12038
rect 7877 6078 7894 12038
rect 7894 6078 7928 12038
rect 7928 6078 7943 12038
rect 8035 6078 8052 12038
rect 8052 6078 8086 12038
rect 8086 6078 8101 12038
rect 8193 6078 8210 12038
rect 8210 6078 8244 12038
rect 8244 6078 8259 12038
rect 8351 6078 8368 12038
rect 8368 6078 8402 12038
rect 8402 6078 8417 12038
rect 8509 6078 8526 12038
rect 8526 6078 8560 12038
rect 8560 6078 8575 12038
rect 8667 6078 8684 12038
rect 8684 6078 8718 12038
rect 8718 6078 8733 12038
rect 8825 6078 8842 12038
rect 8842 6078 8876 12038
rect 8876 6078 8891 12038
rect 8983 6078 9000 12038
rect 9000 6078 9034 12038
rect 9034 6078 9049 12038
rect 9141 6078 9158 12038
rect 9158 6078 9192 12038
rect 9192 6078 9207 12038
rect 9299 6078 9316 12038
rect 9316 6078 9350 12038
rect 9350 6078 9365 12038
rect 9457 6078 9474 12038
rect 9474 6078 9508 12038
rect 9508 6078 9523 12038
rect 9615 6078 9632 12038
rect 9632 6078 9666 12038
rect 9666 6078 9681 12038
rect 9773 6078 9790 12038
rect 9790 6078 9824 12038
rect 9824 6078 9839 12038
rect 9931 6078 9948 12038
rect 9948 6078 9982 12038
rect 9982 6078 9997 12038
rect 10089 6078 10106 12038
rect 10106 6078 10140 12038
rect 10140 6078 10155 12038
rect 10247 6078 10264 12038
rect 10264 6078 10298 12038
rect 10298 6078 10313 12038
rect 10405 6078 10422 12038
rect 10422 6078 10456 12038
rect 10456 6078 10471 12038
rect 5530 5900 5600 6036
rect 10540 6036 10554 12080
rect 10554 6036 10592 12080
rect 10592 6036 10610 12080
rect 5752 6020 10386 6026
rect 5752 5986 5812 6020
rect 5812 5986 5902 6020
rect 5902 5986 5970 6020
rect 5970 5986 6060 6020
rect 6060 5986 6128 6020
rect 6128 5986 6218 6020
rect 6218 5986 6286 6020
rect 6286 5986 6376 6020
rect 6376 5986 6444 6020
rect 6444 5986 6534 6020
rect 6534 5986 6602 6020
rect 6602 5986 6692 6020
rect 6692 5986 6760 6020
rect 6760 5986 6850 6020
rect 6850 5986 6918 6020
rect 6918 5986 7008 6020
rect 7008 5986 7076 6020
rect 7076 5986 7166 6020
rect 7166 5986 7234 6020
rect 7234 5986 7324 6020
rect 7324 5986 7392 6020
rect 7392 5986 7482 6020
rect 7482 5986 7550 6020
rect 7550 5986 7640 6020
rect 7640 5986 7708 6020
rect 7708 5986 7798 6020
rect 7798 5986 7866 6020
rect 7866 5986 7956 6020
rect 7956 5986 8024 6020
rect 8024 5986 8114 6020
rect 8114 5986 8182 6020
rect 8182 5986 8272 6020
rect 8272 5986 8340 6020
rect 8340 5986 8430 6020
rect 8430 5986 8498 6020
rect 8498 5986 8588 6020
rect 8588 5986 8656 6020
rect 8656 5986 8746 6020
rect 8746 5986 8814 6020
rect 8814 5986 8904 6020
rect 8904 5986 8972 6020
rect 8972 5986 9062 6020
rect 9062 5986 9130 6020
rect 9130 5986 9220 6020
rect 9220 5986 9288 6020
rect 9288 5986 9378 6020
rect 9378 5986 9446 6020
rect 9446 5986 9536 6020
rect 9536 5986 9604 6020
rect 9604 5986 9694 6020
rect 9694 5986 9762 6020
rect 9762 5986 9852 6020
rect 9852 5986 9920 6020
rect 9920 5986 10010 6020
rect 10010 5986 10078 6020
rect 10078 5986 10168 6020
rect 10168 5986 10236 6020
rect 10236 5986 10326 6020
rect 10326 5986 10386 6020
rect 5752 5926 10386 5986
rect 10540 5900 10610 6036
<< metal2 >>
rect -8300 49880 -7000 49900
rect -2000 49880 -700 50000
rect 4300 49880 5600 49900
rect -13370 49820 -13300 49880
rect -8360 49820 -7000 49880
rect -13168 49780 -13148 49790
rect -8514 49780 -8494 49790
rect -13168 49710 -13160 49780
rect -8500 49710 -8494 49780
rect -13168 49690 -13148 49710
rect -8514 49690 -8494 49710
rect -13235 49638 -13169 49658
rect -13235 43658 -13169 43678
rect -13077 49638 -13011 49658
rect -13077 43658 -13011 43678
rect -12919 49638 -12853 49658
rect -12919 43658 -12853 43678
rect -12761 49638 -12695 49658
rect -12761 43658 -12695 43678
rect -12603 49638 -12537 49658
rect -12603 43658 -12537 43678
rect -12445 49638 -12379 49658
rect -12445 43658 -12379 43678
rect -12287 49638 -12221 49658
rect -12287 43658 -12221 43678
rect -12129 49638 -12063 49658
rect -12129 43658 -12063 43678
rect -11971 49638 -11905 49658
rect -11971 43658 -11905 43678
rect -11813 49638 -11747 49658
rect -11813 43658 -11747 43678
rect -11655 49638 -11589 49658
rect -11655 43658 -11589 43678
rect -11497 49638 -11431 49658
rect -11497 43658 -11431 43678
rect -11339 49638 -11273 49658
rect -11339 43658 -11273 43678
rect -11181 49638 -11115 49658
rect -11181 43658 -11115 43678
rect -11023 49638 -10957 49658
rect -11023 43658 -10957 43678
rect -10865 49638 -10799 49658
rect -10865 43658 -10799 43678
rect -10707 49638 -10641 49658
rect -10707 43658 -10641 43678
rect -10549 49638 -10483 49658
rect -10549 43658 -10483 43678
rect -10391 49638 -10325 49658
rect -10391 43658 -10325 43678
rect -10233 49638 -10167 49658
rect -10233 43658 -10167 43678
rect -10075 49638 -10009 49658
rect -10075 43658 -10009 43678
rect -9917 49638 -9851 49658
rect -9917 43658 -9851 43678
rect -9759 49638 -9693 49658
rect -9759 43658 -9693 43678
rect -9601 49638 -9535 49658
rect -9601 43658 -9535 43678
rect -9443 49638 -9377 49658
rect -9443 43658 -9377 43678
rect -9285 49638 -9219 49658
rect -9285 43658 -9219 43678
rect -9127 49638 -9061 49658
rect -9127 43658 -9061 43678
rect -8969 49638 -8903 49658
rect -8969 43658 -8903 43678
rect -8811 49638 -8745 49658
rect -8811 43658 -8745 43678
rect -8653 49638 -8587 49658
rect -8653 43658 -8587 43678
rect -8495 49638 -8429 49658
rect -8495 43658 -8429 43678
rect -13168 43610 -13148 43626
rect -8514 43610 -8494 43626
rect -13168 43540 -13160 43610
rect -8510 43540 -8494 43610
rect -13168 43526 -13148 43540
rect -8514 43526 -8494 43540
rect -13370 43430 -13300 43500
rect -8290 49500 -7070 49820
rect -8290 48900 -7070 49300
rect -8290 48300 -7070 48700
rect -8290 47700 -7070 48100
rect -8290 47100 -7070 47500
rect -8290 46500 -7070 46900
rect -8290 45900 -7070 46300
rect -8290 45300 -7070 45700
rect -8290 44700 -7070 45100
rect -8290 44100 -7070 44500
rect -8290 43500 -7070 43900
rect -2060 49820 -700 49880
rect -6868 49780 -6848 49790
rect -2214 49780 -2194 49790
rect -6868 49710 -6860 49780
rect -2200 49710 -2194 49780
rect -6868 49690 -6848 49710
rect -2214 49690 -2194 49710
rect -6935 49638 -6869 49658
rect -6935 43658 -6869 43678
rect -6777 49638 -6711 49658
rect -6777 43658 -6711 43678
rect -6619 49638 -6553 49658
rect -6619 43658 -6553 43678
rect -6461 49638 -6395 49658
rect -6461 43658 -6395 43678
rect -6303 49638 -6237 49658
rect -6303 43658 -6237 43678
rect -6145 49638 -6079 49658
rect -6145 43658 -6079 43678
rect -5987 49638 -5921 49658
rect -5987 43658 -5921 43678
rect -5829 49638 -5763 49658
rect -5829 43658 -5763 43678
rect -5671 49638 -5605 49658
rect -5671 43658 -5605 43678
rect -5513 49638 -5447 49658
rect -5513 43658 -5447 43678
rect -5355 49638 -5289 49658
rect -5355 43658 -5289 43678
rect -5197 49638 -5131 49658
rect -5197 43658 -5131 43678
rect -5039 49638 -4973 49658
rect -5039 43658 -4973 43678
rect -4881 49638 -4815 49658
rect -4881 43658 -4815 43678
rect -4723 49638 -4657 49658
rect -4723 43658 -4657 43678
rect -4565 49638 -4499 49658
rect -4565 43658 -4499 43678
rect -4407 49638 -4341 49658
rect -4407 43658 -4341 43678
rect -4249 49638 -4183 49658
rect -4249 43658 -4183 43678
rect -4091 49638 -4025 49658
rect -4091 43658 -4025 43678
rect -3933 49638 -3867 49658
rect -3933 43658 -3867 43678
rect -3775 49638 -3709 49658
rect -3775 43658 -3709 43678
rect -3617 49638 -3551 49658
rect -3617 43658 -3551 43678
rect -3459 49638 -3393 49658
rect -3459 43658 -3393 43678
rect -3301 49638 -3235 49658
rect -3301 43658 -3235 43678
rect -3143 49638 -3077 49658
rect -3143 43658 -3077 43678
rect -2985 49638 -2919 49658
rect -2985 43658 -2919 43678
rect -2827 49638 -2761 49658
rect -2827 43658 -2761 43678
rect -2669 49638 -2603 49658
rect -2669 43658 -2603 43678
rect -2511 49638 -2445 49658
rect -2511 43658 -2445 43678
rect -2353 49638 -2287 49658
rect -2353 43658 -2287 43678
rect -2195 49638 -2129 49658
rect -2195 43658 -2129 43678
rect -6868 43610 -6848 43626
rect -2214 43610 -2194 43626
rect -6868 43540 -6860 43610
rect -2210 43540 -2194 43610
rect -6868 43526 -6848 43540
rect -2214 43526 -2194 43540
rect -8360 43430 -8290 43500
rect -7900 42900 -7400 43500
rect -7070 43430 -7000 43500
rect -1990 49600 -770 49820
rect -1990 49000 -770 49400
rect -1990 48400 -770 48800
rect -1990 47800 -770 48200
rect -1990 47200 -770 47600
rect -1990 46600 -770 47000
rect -1990 46000 -770 46400
rect -1990 45400 -770 45800
rect -1990 44800 -770 45200
rect -1990 44200 -770 44600
rect -1990 43600 -770 44000
rect -2060 43430 -1990 43500
rect -1600 42900 -1100 43600
rect 4240 49820 5600 49880
rect -568 49780 -548 49790
rect 4086 49780 4106 49790
rect -568 49710 -560 49780
rect 4100 49710 4106 49780
rect -568 49690 -548 49710
rect 4086 49690 4106 49710
rect -635 49638 -569 49658
rect -635 43658 -569 43678
rect -477 49638 -411 49658
rect -477 43658 -411 43678
rect -319 49638 -253 49658
rect -319 43658 -253 43678
rect -161 49638 -95 49658
rect -161 43658 -95 43678
rect -3 49638 63 49658
rect -3 43658 63 43678
rect 155 49638 221 49658
rect 155 43658 221 43678
rect 313 49638 379 49658
rect 313 43658 379 43678
rect 471 49638 537 49658
rect 471 43658 537 43678
rect 629 49638 695 49658
rect 629 43658 695 43678
rect 787 49638 853 49658
rect 787 43658 853 43678
rect 945 49638 1011 49658
rect 945 43658 1011 43678
rect 1103 49638 1169 49658
rect 1103 43658 1169 43678
rect 1261 49638 1327 49658
rect 1261 43658 1327 43678
rect 1419 49638 1485 49658
rect 1419 43658 1485 43678
rect 1577 49638 1643 49658
rect 1577 43658 1643 43678
rect 1735 49638 1801 49658
rect 1735 43658 1801 43678
rect 1893 49638 1959 49658
rect 1893 43658 1959 43678
rect 2051 49638 2117 49658
rect 2051 43658 2117 43678
rect 2209 49638 2275 49658
rect 2209 43658 2275 43678
rect 2367 49638 2433 49658
rect 2367 43658 2433 43678
rect 2525 49638 2591 49658
rect 2525 43658 2591 43678
rect 2683 49638 2749 49658
rect 2683 43658 2749 43678
rect 2841 49638 2907 49658
rect 2841 43658 2907 43678
rect 2999 49638 3065 49658
rect 2999 43658 3065 43678
rect 3157 49638 3223 49658
rect 3157 43658 3223 43678
rect 3315 49638 3381 49658
rect 3315 43658 3381 43678
rect 3473 49638 3539 49658
rect 3473 43658 3539 43678
rect 3631 49638 3697 49658
rect 3631 43658 3697 43678
rect 3789 49638 3855 49658
rect 3789 43658 3855 43678
rect 3947 49638 4013 49658
rect 3947 43658 4013 43678
rect 4105 49638 4171 49658
rect 4105 43658 4171 43678
rect -568 43610 -548 43626
rect 4086 43610 4106 43626
rect -568 43540 -560 43610
rect 4090 43540 4106 43610
rect -568 43526 -548 43540
rect 4086 43526 4106 43540
rect -770 43430 -700 43500
rect 4310 49500 5530 49820
rect 4310 48900 5530 49300
rect 4310 48300 5530 48700
rect 4310 47700 5530 48100
rect 4310 47100 5530 47500
rect 4310 46500 5530 46900
rect 4310 45900 5530 46300
rect 4310 45300 5530 45700
rect 4310 44700 5530 45100
rect 4310 44100 5530 44500
rect 4310 43500 5530 43900
rect 10540 49820 10610 49880
rect 5732 49780 5752 49790
rect 10386 49780 10406 49790
rect 5732 49710 5740 49780
rect 10400 49710 10406 49780
rect 5732 49690 5752 49710
rect 10386 49690 10406 49710
rect 5665 49638 5731 49658
rect 5665 43658 5731 43678
rect 5823 49638 5889 49658
rect 5823 43658 5889 43678
rect 5981 49638 6047 49658
rect 5981 43658 6047 43678
rect 6139 49638 6205 49658
rect 6139 43658 6205 43678
rect 6297 49638 6363 49658
rect 6297 43658 6363 43678
rect 6455 49638 6521 49658
rect 6455 43658 6521 43678
rect 6613 49638 6679 49658
rect 6613 43658 6679 43678
rect 6771 49638 6837 49658
rect 6771 43658 6837 43678
rect 6929 49638 6995 49658
rect 6929 43658 6995 43678
rect 7087 49638 7153 49658
rect 7087 43658 7153 43678
rect 7245 49638 7311 49658
rect 7245 43658 7311 43678
rect 7403 49638 7469 49658
rect 7403 43658 7469 43678
rect 7561 49638 7627 49658
rect 7561 43658 7627 43678
rect 7719 49638 7785 49658
rect 7719 43658 7785 43678
rect 7877 49638 7943 49658
rect 7877 43658 7943 43678
rect 8035 49638 8101 49658
rect 8035 43658 8101 43678
rect 8193 49638 8259 49658
rect 8193 43658 8259 43678
rect 8351 49638 8417 49658
rect 8351 43658 8417 43678
rect 8509 49638 8575 49658
rect 8509 43658 8575 43678
rect 8667 49638 8733 49658
rect 8667 43658 8733 43678
rect 8825 49638 8891 49658
rect 8825 43658 8891 43678
rect 8983 49638 9049 49658
rect 8983 43658 9049 43678
rect 9141 49638 9207 49658
rect 9141 43658 9207 43678
rect 9299 49638 9365 49658
rect 9299 43658 9365 43678
rect 9457 49638 9523 49658
rect 9457 43658 9523 43678
rect 9615 49638 9681 49658
rect 9615 43658 9681 43678
rect 9773 49638 9839 49658
rect 9773 43658 9839 43678
rect 9931 49638 9997 49658
rect 9931 43658 9997 43678
rect 10089 49638 10155 49658
rect 10089 43658 10155 43678
rect 10247 49638 10313 49658
rect 10247 43658 10313 43678
rect 10405 49638 10471 49658
rect 10405 43658 10471 43678
rect 5732 43610 5752 43626
rect 10386 43610 10406 43626
rect 5732 43540 5740 43610
rect 10390 43540 10406 43610
rect 5732 43526 5752 43540
rect 10386 43526 10406 43540
rect 4240 43430 4310 43500
rect 4700 42900 5200 43500
rect 5530 43430 5600 43500
rect 10540 43430 10610 43500
rect -8300 42880 -7000 42900
rect -2000 42880 -700 42900
rect 4300 42880 5600 42900
rect -13370 42820 -13300 42880
rect -8360 42820 -7000 42880
rect -13168 42780 -13148 42790
rect -8514 42780 -8494 42790
rect -13168 42710 -13160 42780
rect -8500 42710 -8494 42780
rect -13168 42690 -13148 42710
rect -8514 42690 -8494 42710
rect -13235 42638 -13169 42658
rect -13235 36658 -13169 36678
rect -13077 42638 -13011 42658
rect -13077 36658 -13011 36678
rect -12919 42638 -12853 42658
rect -12919 36658 -12853 36678
rect -12761 42638 -12695 42658
rect -12761 36658 -12695 36678
rect -12603 42638 -12537 42658
rect -12603 36658 -12537 36678
rect -12445 42638 -12379 42658
rect -12445 36658 -12379 36678
rect -12287 42638 -12221 42658
rect -12287 36658 -12221 36678
rect -12129 42638 -12063 42658
rect -12129 36658 -12063 36678
rect -11971 42638 -11905 42658
rect -11971 36658 -11905 36678
rect -11813 42638 -11747 42658
rect -11813 36658 -11747 36678
rect -11655 42638 -11589 42658
rect -11655 36658 -11589 36678
rect -11497 42638 -11431 42658
rect -11497 36658 -11431 36678
rect -11339 42638 -11273 42658
rect -11339 36658 -11273 36678
rect -11181 42638 -11115 42658
rect -11181 36658 -11115 36678
rect -11023 42638 -10957 42658
rect -11023 36658 -10957 36678
rect -10865 42638 -10799 42658
rect -10865 36658 -10799 36678
rect -10707 42638 -10641 42658
rect -10707 36658 -10641 36678
rect -10549 42638 -10483 42658
rect -10549 36658 -10483 36678
rect -10391 42638 -10325 42658
rect -10391 36658 -10325 36678
rect -10233 42638 -10167 42658
rect -10233 36658 -10167 36678
rect -10075 42638 -10009 42658
rect -10075 36658 -10009 36678
rect -9917 42638 -9851 42658
rect -9917 36658 -9851 36678
rect -9759 42638 -9693 42658
rect -9759 36658 -9693 36678
rect -9601 42638 -9535 42658
rect -9601 36658 -9535 36678
rect -9443 42638 -9377 42658
rect -9443 36658 -9377 36678
rect -9285 42638 -9219 42658
rect -9285 36658 -9219 36678
rect -9127 42638 -9061 42658
rect -9127 36658 -9061 36678
rect -8969 42638 -8903 42658
rect -8969 36658 -8903 36678
rect -8811 42638 -8745 42658
rect -8811 36658 -8745 36678
rect -8653 42638 -8587 42658
rect -8653 36658 -8587 36678
rect -8495 42638 -8429 42658
rect -8495 36658 -8429 36678
rect -13168 36610 -13148 36626
rect -8514 36610 -8494 36626
rect -13168 36540 -13160 36610
rect -8510 36540 -8494 36610
rect -13168 36526 -13148 36540
rect -8514 36526 -8494 36540
rect -13370 36430 -13300 36500
rect -8290 42500 -7070 42820
rect -8290 41900 -7070 42300
rect -8290 41300 -7070 41700
rect -8290 40700 -7070 41100
rect -8290 40100 -7070 40500
rect -8290 39500 -7070 39900
rect -8290 38900 -7070 39300
rect -8290 38300 -7070 38700
rect -8290 37700 -7070 38100
rect -8290 37100 -7070 37500
rect -8290 36500 -7070 36900
rect -2060 42820 -700 42880
rect -6868 42780 -6848 42790
rect -2214 42780 -2194 42790
rect -6868 42710 -6860 42780
rect -2200 42710 -2194 42780
rect -6868 42690 -6848 42710
rect -2214 42690 -2194 42710
rect -6935 42638 -6869 42658
rect -6935 36658 -6869 36678
rect -6777 42638 -6711 42658
rect -6777 36658 -6711 36678
rect -6619 42638 -6553 42658
rect -6619 36658 -6553 36678
rect -6461 42638 -6395 42658
rect -6461 36658 -6395 36678
rect -6303 42638 -6237 42658
rect -6303 36658 -6237 36678
rect -6145 42638 -6079 42658
rect -6145 36658 -6079 36678
rect -5987 42638 -5921 42658
rect -5987 36658 -5921 36678
rect -5829 42638 -5763 42658
rect -5829 36658 -5763 36678
rect -5671 42638 -5605 42658
rect -5671 36658 -5605 36678
rect -5513 42638 -5447 42658
rect -5513 36658 -5447 36678
rect -5355 42638 -5289 42658
rect -5355 36658 -5289 36678
rect -5197 42638 -5131 42658
rect -5197 36658 -5131 36678
rect -5039 42638 -4973 42658
rect -5039 36658 -4973 36678
rect -4881 42638 -4815 42658
rect -4881 36658 -4815 36678
rect -4723 42638 -4657 42658
rect -4723 36658 -4657 36678
rect -4565 42638 -4499 42658
rect -4565 36658 -4499 36678
rect -4407 42638 -4341 42658
rect -4407 36658 -4341 36678
rect -4249 42638 -4183 42658
rect -4249 36658 -4183 36678
rect -4091 42638 -4025 42658
rect -4091 36658 -4025 36678
rect -3933 42638 -3867 42658
rect -3933 36658 -3867 36678
rect -3775 42638 -3709 42658
rect -3775 36658 -3709 36678
rect -3617 42638 -3551 42658
rect -3617 36658 -3551 36678
rect -3459 42638 -3393 42658
rect -3459 36658 -3393 36678
rect -3301 42638 -3235 42658
rect -3301 36658 -3235 36678
rect -3143 42638 -3077 42658
rect -3143 36658 -3077 36678
rect -2985 42638 -2919 42658
rect -2985 36658 -2919 36678
rect -2827 42638 -2761 42658
rect -2827 36658 -2761 36678
rect -2669 42638 -2603 42658
rect -2669 36658 -2603 36678
rect -2511 42638 -2445 42658
rect -2511 36658 -2445 36678
rect -2353 42638 -2287 42658
rect -2353 36658 -2287 36678
rect -2195 42638 -2129 42658
rect -2195 36658 -2129 36678
rect -6868 36610 -6848 36626
rect -2214 36610 -2194 36626
rect -6868 36540 -6860 36610
rect -2210 36540 -2194 36610
rect -6868 36526 -6848 36540
rect -2214 36526 -2194 36540
rect -8360 36430 -8290 36500
rect -7070 36430 -7000 36500
rect -1990 42500 -770 42820
rect -1990 41900 -770 42300
rect -1990 41300 -770 41700
rect -1990 40700 -770 41100
rect -1990 40100 -770 40500
rect -1990 39500 -770 39900
rect -1990 38900 -770 39300
rect -1990 38300 -770 38700
rect -1990 37700 -770 38100
rect -1990 37100 -770 37500
rect -1990 36500 -770 36900
rect 4240 42820 5600 42880
rect -568 42780 -548 42790
rect 4086 42780 4106 42790
rect -568 42710 -560 42780
rect 4100 42710 4106 42780
rect -568 42690 -548 42710
rect 4086 42690 4106 42710
rect -635 42638 -569 42658
rect -635 36658 -569 36678
rect -477 42638 -411 42658
rect -477 36658 -411 36678
rect -319 42638 -253 42658
rect -319 36658 -253 36678
rect -161 42638 -95 42658
rect -161 36658 -95 36678
rect -3 42638 63 42658
rect -3 36658 63 36678
rect 155 42638 221 42658
rect 155 36658 221 36678
rect 313 42638 379 42658
rect 313 36658 379 36678
rect 471 42638 537 42658
rect 471 36658 537 36678
rect 629 42638 695 42658
rect 629 36658 695 36678
rect 787 42638 853 42658
rect 787 36658 853 36678
rect 945 42638 1011 42658
rect 945 36658 1011 36678
rect 1103 42638 1169 42658
rect 1103 36658 1169 36678
rect 1261 42638 1327 42658
rect 1261 36658 1327 36678
rect 1419 42638 1485 42658
rect 1419 36658 1485 36678
rect 1577 42638 1643 42658
rect 1577 36658 1643 36678
rect 1735 42638 1801 42658
rect 1735 36658 1801 36678
rect 1893 42638 1959 42658
rect 1893 36658 1959 36678
rect 2051 42638 2117 42658
rect 2051 36658 2117 36678
rect 2209 42638 2275 42658
rect 2209 36658 2275 36678
rect 2367 42638 2433 42658
rect 2367 36658 2433 36678
rect 2525 42638 2591 42658
rect 2525 36658 2591 36678
rect 2683 42638 2749 42658
rect 2683 36658 2749 36678
rect 2841 42638 2907 42658
rect 2841 36658 2907 36678
rect 2999 42638 3065 42658
rect 2999 36658 3065 36678
rect 3157 42638 3223 42658
rect 3157 36658 3223 36678
rect 3315 42638 3381 42658
rect 3315 36658 3381 36678
rect 3473 42638 3539 42658
rect 3473 36658 3539 36678
rect 3631 42638 3697 42658
rect 3631 36658 3697 36678
rect 3789 42638 3855 42658
rect 3789 36658 3855 36678
rect 3947 42638 4013 42658
rect 3947 36658 4013 36678
rect 4105 42638 4171 42658
rect 4105 36658 4171 36678
rect -568 36610 -548 36626
rect 4086 36610 4106 36626
rect -568 36540 -560 36610
rect 4090 36540 4106 36610
rect -568 36526 -548 36540
rect 4086 36526 4106 36540
rect -2060 36430 -1990 36500
rect -770 36430 -700 36500
rect 4310 42500 5530 42820
rect 4310 41900 5530 42300
rect 4310 41300 5530 41700
rect 4310 40700 5530 41100
rect 4310 40100 5530 40500
rect 4310 39500 5530 39900
rect 4310 38900 5530 39300
rect 4310 38300 5530 38700
rect 4310 37700 5530 38100
rect 4310 37100 5530 37500
rect 4310 36500 5530 36900
rect 10540 42820 10610 42880
rect 5732 42780 5752 42790
rect 10386 42780 10406 42790
rect 5732 42710 5740 42780
rect 10400 42710 10406 42780
rect 5732 42690 5752 42710
rect 10386 42690 10406 42710
rect 5665 42638 5731 42658
rect 5665 36658 5731 36678
rect 5823 42638 5889 42658
rect 5823 36658 5889 36678
rect 5981 42638 6047 42658
rect 5981 36658 6047 36678
rect 6139 42638 6205 42658
rect 6139 36658 6205 36678
rect 6297 42638 6363 42658
rect 6297 36658 6363 36678
rect 6455 42638 6521 42658
rect 6455 36658 6521 36678
rect 6613 42638 6679 42658
rect 6613 36658 6679 36678
rect 6771 42638 6837 42658
rect 6771 36658 6837 36678
rect 6929 42638 6995 42658
rect 6929 36658 6995 36678
rect 7087 42638 7153 42658
rect 7087 36658 7153 36678
rect 7245 42638 7311 42658
rect 7245 36658 7311 36678
rect 7403 42638 7469 42658
rect 7403 36658 7469 36678
rect 7561 42638 7627 42658
rect 7561 36658 7627 36678
rect 7719 42638 7785 42658
rect 7719 36658 7785 36678
rect 7877 42638 7943 42658
rect 7877 36658 7943 36678
rect 8035 42638 8101 42658
rect 8035 36658 8101 36678
rect 8193 42638 8259 42658
rect 8193 36658 8259 36678
rect 8351 42638 8417 42658
rect 8351 36658 8417 36678
rect 8509 42638 8575 42658
rect 8509 36658 8575 36678
rect 8667 42638 8733 42658
rect 8667 36658 8733 36678
rect 8825 42638 8891 42658
rect 8825 36658 8891 36678
rect 8983 42638 9049 42658
rect 8983 36658 9049 36678
rect 9141 42638 9207 42658
rect 9141 36658 9207 36678
rect 9299 42638 9365 42658
rect 9299 36658 9365 36678
rect 9457 42638 9523 42658
rect 9457 36658 9523 36678
rect 9615 42638 9681 42658
rect 9615 36658 9681 36678
rect 9773 42638 9839 42658
rect 9773 36658 9839 36678
rect 9931 42638 9997 42658
rect 9931 36658 9997 36678
rect 10089 42638 10155 42658
rect 10089 36658 10155 36678
rect 10247 42638 10313 42658
rect 10247 36658 10313 36678
rect 10405 42638 10471 42658
rect 10405 36658 10471 36678
rect 5732 36610 5752 36626
rect 10386 36610 10406 36626
rect 5732 36540 5740 36610
rect 10390 36540 10406 36610
rect 5732 36526 5752 36540
rect 10386 36526 10406 36540
rect 4240 36430 4310 36500
rect 5530 36430 5600 36500
rect 10540 36430 10610 36500
rect -8300 34580 -7000 34600
rect -2000 34580 -700 34700
rect 4300 34580 5600 34600
rect -13370 34520 -13300 34580
rect -8360 34520 -7000 34580
rect -13168 34480 -13148 34490
rect -8514 34480 -8494 34490
rect -13168 34410 -13160 34480
rect -8500 34410 -8494 34480
rect -13168 34390 -13148 34410
rect -8514 34390 -8494 34410
rect -13235 34338 -13169 34358
rect -13235 28358 -13169 28378
rect -13077 34338 -13011 34358
rect -13077 28358 -13011 28378
rect -12919 34338 -12853 34358
rect -12919 28358 -12853 28378
rect -12761 34338 -12695 34358
rect -12761 28358 -12695 28378
rect -12603 34338 -12537 34358
rect -12603 28358 -12537 28378
rect -12445 34338 -12379 34358
rect -12445 28358 -12379 28378
rect -12287 34338 -12221 34358
rect -12287 28358 -12221 28378
rect -12129 34338 -12063 34358
rect -12129 28358 -12063 28378
rect -11971 34338 -11905 34358
rect -11971 28358 -11905 28378
rect -11813 34338 -11747 34358
rect -11813 28358 -11747 28378
rect -11655 34338 -11589 34358
rect -11655 28358 -11589 28378
rect -11497 34338 -11431 34358
rect -11497 28358 -11431 28378
rect -11339 34338 -11273 34358
rect -11339 28358 -11273 28378
rect -11181 34338 -11115 34358
rect -11181 28358 -11115 28378
rect -11023 34338 -10957 34358
rect -11023 28358 -10957 28378
rect -10865 34338 -10799 34358
rect -10865 28358 -10799 28378
rect -10707 34338 -10641 34358
rect -10707 28358 -10641 28378
rect -10549 34338 -10483 34358
rect -10549 28358 -10483 28378
rect -10391 34338 -10325 34358
rect -10391 28358 -10325 28378
rect -10233 34338 -10167 34358
rect -10233 28358 -10167 28378
rect -10075 34338 -10009 34358
rect -10075 28358 -10009 28378
rect -9917 34338 -9851 34358
rect -9917 28358 -9851 28378
rect -9759 34338 -9693 34358
rect -9759 28358 -9693 28378
rect -9601 34338 -9535 34358
rect -9601 28358 -9535 28378
rect -9443 34338 -9377 34358
rect -9443 28358 -9377 28378
rect -9285 34338 -9219 34358
rect -9285 28358 -9219 28378
rect -9127 34338 -9061 34358
rect -9127 28358 -9061 28378
rect -8969 34338 -8903 34358
rect -8969 28358 -8903 28378
rect -8811 34338 -8745 34358
rect -8811 28358 -8745 28378
rect -8653 34338 -8587 34358
rect -8653 28358 -8587 28378
rect -8495 34338 -8429 34358
rect -8495 28358 -8429 28378
rect -13168 28310 -13148 28326
rect -8514 28310 -8494 28326
rect -13168 28240 -13160 28310
rect -8510 28240 -8494 28310
rect -13168 28226 -13148 28240
rect -8514 28226 -8494 28240
rect -13370 28130 -13300 28200
rect -8290 34200 -7070 34520
rect -8290 33600 -7070 34000
rect -8290 33000 -7070 33400
rect -8290 32400 -7070 32800
rect -8290 31800 -7070 32200
rect -8290 31200 -7070 31600
rect -8290 30600 -7070 31000
rect -8290 30000 -7070 30400
rect -8290 29400 -7070 29800
rect -8290 28800 -7070 29200
rect -8290 28200 -7070 28600
rect -2060 34520 -700 34580
rect -6868 34480 -6848 34490
rect -2214 34480 -2194 34490
rect -6868 34410 -6860 34480
rect -2200 34410 -2194 34480
rect -6868 34390 -6848 34410
rect -2214 34390 -2194 34410
rect -6935 34338 -6869 34358
rect -6935 28358 -6869 28378
rect -6777 34338 -6711 34358
rect -6777 28358 -6711 28378
rect -6619 34338 -6553 34358
rect -6619 28358 -6553 28378
rect -6461 34338 -6395 34358
rect -6461 28358 -6395 28378
rect -6303 34338 -6237 34358
rect -6303 28358 -6237 28378
rect -6145 34338 -6079 34358
rect -6145 28358 -6079 28378
rect -5987 34338 -5921 34358
rect -5987 28358 -5921 28378
rect -5829 34338 -5763 34358
rect -5829 28358 -5763 28378
rect -5671 34338 -5605 34358
rect -5671 28358 -5605 28378
rect -5513 34338 -5447 34358
rect -5513 28358 -5447 28378
rect -5355 34338 -5289 34358
rect -5355 28358 -5289 28378
rect -5197 34338 -5131 34358
rect -5197 28358 -5131 28378
rect -5039 34338 -4973 34358
rect -5039 28358 -4973 28378
rect -4881 34338 -4815 34358
rect -4881 28358 -4815 28378
rect -4723 34338 -4657 34358
rect -4723 28358 -4657 28378
rect -4565 34338 -4499 34358
rect -4565 28358 -4499 28378
rect -4407 34338 -4341 34358
rect -4407 28358 -4341 28378
rect -4249 34338 -4183 34358
rect -4249 28358 -4183 28378
rect -4091 34338 -4025 34358
rect -4091 28358 -4025 28378
rect -3933 34338 -3867 34358
rect -3933 28358 -3867 28378
rect -3775 34338 -3709 34358
rect -3775 28358 -3709 28378
rect -3617 34338 -3551 34358
rect -3617 28358 -3551 28378
rect -3459 34338 -3393 34358
rect -3459 28358 -3393 28378
rect -3301 34338 -3235 34358
rect -3301 28358 -3235 28378
rect -3143 34338 -3077 34358
rect -3143 28358 -3077 28378
rect -2985 34338 -2919 34358
rect -2985 28358 -2919 28378
rect -2827 34338 -2761 34358
rect -2827 28358 -2761 28378
rect -2669 34338 -2603 34358
rect -2669 28358 -2603 28378
rect -2511 34338 -2445 34358
rect -2511 28358 -2445 28378
rect -2353 34338 -2287 34358
rect -2353 28358 -2287 28378
rect -2195 34338 -2129 34358
rect -2195 28358 -2129 28378
rect -6868 28310 -6848 28326
rect -2214 28310 -2194 28326
rect -6868 28240 -6860 28310
rect -2210 28240 -2194 28310
rect -6868 28226 -6848 28240
rect -2214 28226 -2194 28240
rect -8360 28130 -8290 28200
rect -7900 27600 -7400 28200
rect -7070 28130 -7000 28200
rect -1990 34300 -770 34520
rect -1990 33700 -770 34100
rect -1990 33100 -770 33500
rect -1990 32500 -770 32900
rect -1990 31900 -770 32300
rect -1990 31300 -770 31700
rect -1990 30700 -770 31100
rect -1990 30100 -770 30500
rect -1990 29500 -770 29900
rect -1990 28900 -770 29300
rect -1990 28300 -770 28700
rect -2060 28130 -1990 28200
rect -1600 27600 -1100 28300
rect 4240 34520 5600 34580
rect -568 34480 -548 34490
rect 4086 34480 4106 34490
rect -568 34410 -560 34480
rect 4100 34410 4106 34480
rect -568 34390 -548 34410
rect 4086 34390 4106 34410
rect -635 34338 -569 34358
rect -635 28358 -569 28378
rect -477 34338 -411 34358
rect -477 28358 -411 28378
rect -319 34338 -253 34358
rect -319 28358 -253 28378
rect -161 34338 -95 34358
rect -161 28358 -95 28378
rect -3 34338 63 34358
rect -3 28358 63 28378
rect 155 34338 221 34358
rect 155 28358 221 28378
rect 313 34338 379 34358
rect 313 28358 379 28378
rect 471 34338 537 34358
rect 471 28358 537 28378
rect 629 34338 695 34358
rect 629 28358 695 28378
rect 787 34338 853 34358
rect 787 28358 853 28378
rect 945 34338 1011 34358
rect 945 28358 1011 28378
rect 1103 34338 1169 34358
rect 1103 28358 1169 28378
rect 1261 34338 1327 34358
rect 1261 28358 1327 28378
rect 1419 34338 1485 34358
rect 1419 28358 1485 28378
rect 1577 34338 1643 34358
rect 1577 28358 1643 28378
rect 1735 34338 1801 34358
rect 1735 28358 1801 28378
rect 1893 34338 1959 34358
rect 1893 28358 1959 28378
rect 2051 34338 2117 34358
rect 2051 28358 2117 28378
rect 2209 34338 2275 34358
rect 2209 28358 2275 28378
rect 2367 34338 2433 34358
rect 2367 28358 2433 28378
rect 2525 34338 2591 34358
rect 2525 28358 2591 28378
rect 2683 34338 2749 34358
rect 2683 28358 2749 28378
rect 2841 34338 2907 34358
rect 2841 28358 2907 28378
rect 2999 34338 3065 34358
rect 2999 28358 3065 28378
rect 3157 34338 3223 34358
rect 3157 28358 3223 28378
rect 3315 34338 3381 34358
rect 3315 28358 3381 28378
rect 3473 34338 3539 34358
rect 3473 28358 3539 28378
rect 3631 34338 3697 34358
rect 3631 28358 3697 28378
rect 3789 34338 3855 34358
rect 3789 28358 3855 28378
rect 3947 34338 4013 34358
rect 3947 28358 4013 28378
rect 4105 34338 4171 34358
rect 4105 28358 4171 28378
rect -568 28310 -548 28326
rect 4086 28310 4106 28326
rect -568 28240 -560 28310
rect 4090 28240 4106 28310
rect -568 28226 -548 28240
rect 4086 28226 4106 28240
rect -770 28130 -700 28200
rect 4310 34200 5530 34520
rect 4310 33600 5530 34000
rect 4310 33000 5530 33400
rect 4310 32400 5530 32800
rect 4310 31800 5530 32200
rect 4310 31200 5530 31600
rect 4310 30600 5530 31000
rect 4310 30000 5530 30400
rect 4310 29400 5530 29800
rect 4310 28800 5530 29200
rect 4310 28200 5530 28600
rect 10540 34520 10610 34580
rect 5732 34480 5752 34490
rect 10386 34480 10406 34490
rect 5732 34410 5740 34480
rect 10400 34410 10406 34480
rect 5732 34390 5752 34410
rect 10386 34390 10406 34410
rect 5665 34338 5731 34358
rect 5665 28358 5731 28378
rect 5823 34338 5889 34358
rect 5823 28358 5889 28378
rect 5981 34338 6047 34358
rect 5981 28358 6047 28378
rect 6139 34338 6205 34358
rect 6139 28358 6205 28378
rect 6297 34338 6363 34358
rect 6297 28358 6363 28378
rect 6455 34338 6521 34358
rect 6455 28358 6521 28378
rect 6613 34338 6679 34358
rect 6613 28358 6679 28378
rect 6771 34338 6837 34358
rect 6771 28358 6837 28378
rect 6929 34338 6995 34358
rect 6929 28358 6995 28378
rect 7087 34338 7153 34358
rect 7087 28358 7153 28378
rect 7245 34338 7311 34358
rect 7245 28358 7311 28378
rect 7403 34338 7469 34358
rect 7403 28358 7469 28378
rect 7561 34338 7627 34358
rect 7561 28358 7627 28378
rect 7719 34338 7785 34358
rect 7719 28358 7785 28378
rect 7877 34338 7943 34358
rect 7877 28358 7943 28378
rect 8035 34338 8101 34358
rect 8035 28358 8101 28378
rect 8193 34338 8259 34358
rect 8193 28358 8259 28378
rect 8351 34338 8417 34358
rect 8351 28358 8417 28378
rect 8509 34338 8575 34358
rect 8509 28358 8575 28378
rect 8667 34338 8733 34358
rect 8667 28358 8733 28378
rect 8825 34338 8891 34358
rect 8825 28358 8891 28378
rect 8983 34338 9049 34358
rect 8983 28358 9049 28378
rect 9141 34338 9207 34358
rect 9141 28358 9207 28378
rect 9299 34338 9365 34358
rect 9299 28358 9365 28378
rect 9457 34338 9523 34358
rect 9457 28358 9523 28378
rect 9615 34338 9681 34358
rect 9615 28358 9681 28378
rect 9773 34338 9839 34358
rect 9773 28358 9839 28378
rect 9931 34338 9997 34358
rect 9931 28358 9997 28378
rect 10089 34338 10155 34358
rect 10089 28358 10155 28378
rect 10247 34338 10313 34358
rect 10247 28358 10313 28378
rect 10405 34338 10471 34358
rect 10405 28358 10471 28378
rect 5732 28310 5752 28326
rect 10386 28310 10406 28326
rect 5732 28240 5740 28310
rect 10390 28240 10406 28310
rect 5732 28226 5752 28240
rect 10386 28226 10406 28240
rect 4240 28130 4310 28200
rect 4700 27600 5200 28200
rect 5530 28130 5600 28200
rect 10540 28130 10610 28200
rect -8300 27580 -7000 27600
rect -2000 27580 -700 27600
rect 4300 27580 5600 27600
rect -13370 27520 -13300 27580
rect -8360 27520 -7000 27580
rect -13168 27480 -13148 27490
rect -8514 27480 -8494 27490
rect -13168 27410 -13160 27480
rect -8500 27410 -8494 27480
rect -13168 27390 -13148 27410
rect -8514 27390 -8494 27410
rect -13235 27338 -13169 27358
rect -13235 21358 -13169 21378
rect -13077 27338 -13011 27358
rect -13077 21358 -13011 21378
rect -12919 27338 -12853 27358
rect -12919 21358 -12853 21378
rect -12761 27338 -12695 27358
rect -12761 21358 -12695 21378
rect -12603 27338 -12537 27358
rect -12603 21358 -12537 21378
rect -12445 27338 -12379 27358
rect -12445 21358 -12379 21378
rect -12287 27338 -12221 27358
rect -12287 21358 -12221 21378
rect -12129 27338 -12063 27358
rect -12129 21358 -12063 21378
rect -11971 27338 -11905 27358
rect -11971 21358 -11905 21378
rect -11813 27338 -11747 27358
rect -11813 21358 -11747 21378
rect -11655 27338 -11589 27358
rect -11655 21358 -11589 21378
rect -11497 27338 -11431 27358
rect -11497 21358 -11431 21378
rect -11339 27338 -11273 27358
rect -11339 21358 -11273 21378
rect -11181 27338 -11115 27358
rect -11181 21358 -11115 21378
rect -11023 27338 -10957 27358
rect -11023 21358 -10957 21378
rect -10865 27338 -10799 27358
rect -10865 21358 -10799 21378
rect -10707 27338 -10641 27358
rect -10707 21358 -10641 21378
rect -10549 27338 -10483 27358
rect -10549 21358 -10483 21378
rect -10391 27338 -10325 27358
rect -10391 21358 -10325 21378
rect -10233 27338 -10167 27358
rect -10233 21358 -10167 21378
rect -10075 27338 -10009 27358
rect -10075 21358 -10009 21378
rect -9917 27338 -9851 27358
rect -9917 21358 -9851 21378
rect -9759 27338 -9693 27358
rect -9759 21358 -9693 21378
rect -9601 27338 -9535 27358
rect -9601 21358 -9535 21378
rect -9443 27338 -9377 27358
rect -9443 21358 -9377 21378
rect -9285 27338 -9219 27358
rect -9285 21358 -9219 21378
rect -9127 27338 -9061 27358
rect -9127 21358 -9061 21378
rect -8969 27338 -8903 27358
rect -8969 21358 -8903 21378
rect -8811 27338 -8745 27358
rect -8811 21358 -8745 21378
rect -8653 27338 -8587 27358
rect -8653 21358 -8587 21378
rect -8495 27338 -8429 27358
rect -8495 21358 -8429 21378
rect -13168 21310 -13148 21326
rect -8514 21310 -8494 21326
rect -13168 21240 -13160 21310
rect -8510 21240 -8494 21310
rect -13168 21226 -13148 21240
rect -8514 21226 -8494 21240
rect -13370 21130 -13300 21200
rect -8290 27200 -7070 27520
rect -8290 26600 -7070 27000
rect -8290 26000 -7070 26400
rect -8290 25400 -7070 25800
rect -8290 24800 -7070 25200
rect -8290 24200 -7070 24600
rect -8290 23600 -7070 24000
rect -8290 23000 -7070 23400
rect -8290 22400 -7070 22800
rect -8290 21800 -7070 22200
rect -8290 21200 -7070 21600
rect -2060 27520 -700 27580
rect -6868 27480 -6848 27490
rect -2214 27480 -2194 27490
rect -6868 27410 -6860 27480
rect -2200 27410 -2194 27480
rect -6868 27390 -6848 27410
rect -2214 27390 -2194 27410
rect -6935 27338 -6869 27358
rect -6935 21358 -6869 21378
rect -6777 27338 -6711 27358
rect -6777 21358 -6711 21378
rect -6619 27338 -6553 27358
rect -6619 21358 -6553 21378
rect -6461 27338 -6395 27358
rect -6461 21358 -6395 21378
rect -6303 27338 -6237 27358
rect -6303 21358 -6237 21378
rect -6145 27338 -6079 27358
rect -6145 21358 -6079 21378
rect -5987 27338 -5921 27358
rect -5987 21358 -5921 21378
rect -5829 27338 -5763 27358
rect -5829 21358 -5763 21378
rect -5671 27338 -5605 27358
rect -5671 21358 -5605 21378
rect -5513 27338 -5447 27358
rect -5513 21358 -5447 21378
rect -5355 27338 -5289 27358
rect -5355 21358 -5289 21378
rect -5197 27338 -5131 27358
rect -5197 21358 -5131 21378
rect -5039 27338 -4973 27358
rect -5039 21358 -4973 21378
rect -4881 27338 -4815 27358
rect -4881 21358 -4815 21378
rect -4723 27338 -4657 27358
rect -4723 21358 -4657 21378
rect -4565 27338 -4499 27358
rect -4565 21358 -4499 21378
rect -4407 27338 -4341 27358
rect -4407 21358 -4341 21378
rect -4249 27338 -4183 27358
rect -4249 21358 -4183 21378
rect -4091 27338 -4025 27358
rect -4091 21358 -4025 21378
rect -3933 27338 -3867 27358
rect -3933 21358 -3867 21378
rect -3775 27338 -3709 27358
rect -3775 21358 -3709 21378
rect -3617 27338 -3551 27358
rect -3617 21358 -3551 21378
rect -3459 27338 -3393 27358
rect -3459 21358 -3393 21378
rect -3301 27338 -3235 27358
rect -3301 21358 -3235 21378
rect -3143 27338 -3077 27358
rect -3143 21358 -3077 21378
rect -2985 27338 -2919 27358
rect -2985 21358 -2919 21378
rect -2827 27338 -2761 27358
rect -2827 21358 -2761 21378
rect -2669 27338 -2603 27358
rect -2669 21358 -2603 21378
rect -2511 27338 -2445 27358
rect -2511 21358 -2445 21378
rect -2353 27338 -2287 27358
rect -2353 21358 -2287 21378
rect -2195 27338 -2129 27358
rect -2195 21358 -2129 21378
rect -6868 21310 -6848 21326
rect -2214 21310 -2194 21326
rect -6868 21240 -6860 21310
rect -2210 21240 -2194 21310
rect -6868 21226 -6848 21240
rect -2214 21226 -2194 21240
rect -8360 21130 -8290 21200
rect -7070 21130 -7000 21200
rect -1990 27200 -770 27520
rect -1990 26600 -770 27000
rect -1990 26000 -770 26400
rect -1990 25400 -770 25800
rect -1990 24800 -770 25200
rect -1990 24200 -770 24600
rect -1990 23600 -770 24000
rect -1990 23000 -770 23400
rect -1990 22400 -770 22800
rect -1990 21800 -770 22200
rect -1990 21200 -770 21600
rect 4240 27520 5600 27580
rect -568 27480 -548 27490
rect 4086 27480 4106 27490
rect -568 27410 -560 27480
rect 4100 27410 4106 27480
rect -568 27390 -548 27410
rect 4086 27390 4106 27410
rect -635 27338 -569 27358
rect -635 21358 -569 21378
rect -477 27338 -411 27358
rect -477 21358 -411 21378
rect -319 27338 -253 27358
rect -319 21358 -253 21378
rect -161 27338 -95 27358
rect -161 21358 -95 21378
rect -3 27338 63 27358
rect -3 21358 63 21378
rect 155 27338 221 27358
rect 155 21358 221 21378
rect 313 27338 379 27358
rect 313 21358 379 21378
rect 471 27338 537 27358
rect 471 21358 537 21378
rect 629 27338 695 27358
rect 629 21358 695 21378
rect 787 27338 853 27358
rect 787 21358 853 21378
rect 945 27338 1011 27358
rect 945 21358 1011 21378
rect 1103 27338 1169 27358
rect 1103 21358 1169 21378
rect 1261 27338 1327 27358
rect 1261 21358 1327 21378
rect 1419 27338 1485 27358
rect 1419 21358 1485 21378
rect 1577 27338 1643 27358
rect 1577 21358 1643 21378
rect 1735 27338 1801 27358
rect 1735 21358 1801 21378
rect 1893 27338 1959 27358
rect 1893 21358 1959 21378
rect 2051 27338 2117 27358
rect 2051 21358 2117 21378
rect 2209 27338 2275 27358
rect 2209 21358 2275 21378
rect 2367 27338 2433 27358
rect 2367 21358 2433 21378
rect 2525 27338 2591 27358
rect 2525 21358 2591 21378
rect 2683 27338 2749 27358
rect 2683 21358 2749 21378
rect 2841 27338 2907 27358
rect 2841 21358 2907 21378
rect 2999 27338 3065 27358
rect 2999 21358 3065 21378
rect 3157 27338 3223 27358
rect 3157 21358 3223 21378
rect 3315 27338 3381 27358
rect 3315 21358 3381 21378
rect 3473 27338 3539 27358
rect 3473 21358 3539 21378
rect 3631 27338 3697 27358
rect 3631 21358 3697 21378
rect 3789 27338 3855 27358
rect 3789 21358 3855 21378
rect 3947 27338 4013 27358
rect 3947 21358 4013 21378
rect 4105 27338 4171 27358
rect 4105 21358 4171 21378
rect -568 21310 -548 21326
rect 4086 21310 4106 21326
rect -568 21240 -560 21310
rect 4090 21240 4106 21310
rect -568 21226 -548 21240
rect 4086 21226 4106 21240
rect -2060 21130 -1990 21200
rect -770 21130 -700 21200
rect 4310 27200 5530 27520
rect 4310 26600 5530 27000
rect 4310 26000 5530 26400
rect 4310 25400 5530 25800
rect 4310 24800 5530 25200
rect 4310 24200 5530 24600
rect 4310 23600 5530 24000
rect 4310 23000 5530 23400
rect 4310 22400 5530 22800
rect 4310 21800 5530 22200
rect 4310 21200 5530 21600
rect 10540 27520 10610 27580
rect 5732 27480 5752 27490
rect 10386 27480 10406 27490
rect 5732 27410 5740 27480
rect 10400 27410 10406 27480
rect 5732 27390 5752 27410
rect 10386 27390 10406 27410
rect 5665 27338 5731 27358
rect 5665 21358 5731 21378
rect 5823 27338 5889 27358
rect 5823 21358 5889 21378
rect 5981 27338 6047 27358
rect 5981 21358 6047 21378
rect 6139 27338 6205 27358
rect 6139 21358 6205 21378
rect 6297 27338 6363 27358
rect 6297 21358 6363 21378
rect 6455 27338 6521 27358
rect 6455 21358 6521 21378
rect 6613 27338 6679 27358
rect 6613 21358 6679 21378
rect 6771 27338 6837 27358
rect 6771 21358 6837 21378
rect 6929 27338 6995 27358
rect 6929 21358 6995 21378
rect 7087 27338 7153 27358
rect 7087 21358 7153 21378
rect 7245 27338 7311 27358
rect 7245 21358 7311 21378
rect 7403 27338 7469 27358
rect 7403 21358 7469 21378
rect 7561 27338 7627 27358
rect 7561 21358 7627 21378
rect 7719 27338 7785 27358
rect 7719 21358 7785 21378
rect 7877 27338 7943 27358
rect 7877 21358 7943 21378
rect 8035 27338 8101 27358
rect 8035 21358 8101 21378
rect 8193 27338 8259 27358
rect 8193 21358 8259 21378
rect 8351 27338 8417 27358
rect 8351 21358 8417 21378
rect 8509 27338 8575 27358
rect 8509 21358 8575 21378
rect 8667 27338 8733 27358
rect 8667 21358 8733 21378
rect 8825 27338 8891 27358
rect 8825 21358 8891 21378
rect 8983 27338 9049 27358
rect 8983 21358 9049 21378
rect 9141 27338 9207 27358
rect 9141 21358 9207 21378
rect 9299 27338 9365 27358
rect 9299 21358 9365 21378
rect 9457 27338 9523 27358
rect 9457 21358 9523 21378
rect 9615 27338 9681 27358
rect 9615 21358 9681 21378
rect 9773 27338 9839 27358
rect 9773 21358 9839 21378
rect 9931 27338 9997 27358
rect 9931 21358 9997 21378
rect 10089 27338 10155 27358
rect 10089 21358 10155 21378
rect 10247 27338 10313 27358
rect 10247 21358 10313 21378
rect 10405 27338 10471 27358
rect 10405 21358 10471 21378
rect 5732 21310 5752 21326
rect 10386 21310 10406 21326
rect 5732 21240 5740 21310
rect 10390 21240 10406 21310
rect 5732 21226 5752 21240
rect 10386 21226 10406 21240
rect 4240 21130 4310 21200
rect 5530 21130 5600 21200
rect 10540 21130 10610 21200
rect -8300 19280 -7000 19300
rect -2000 19280 -700 19400
rect 4300 19280 5600 19300
rect -13370 19220 -13300 19280
rect -8360 19220 -7000 19280
rect -13168 19180 -13148 19190
rect -8514 19180 -8494 19190
rect -13168 19110 -13160 19180
rect -8500 19110 -8494 19180
rect -13168 19090 -13148 19110
rect -8514 19090 -8494 19110
rect -13235 19038 -13169 19058
rect -13235 13058 -13169 13078
rect -13077 19038 -13011 19058
rect -13077 13058 -13011 13078
rect -12919 19038 -12853 19058
rect -12919 13058 -12853 13078
rect -12761 19038 -12695 19058
rect -12761 13058 -12695 13078
rect -12603 19038 -12537 19058
rect -12603 13058 -12537 13078
rect -12445 19038 -12379 19058
rect -12445 13058 -12379 13078
rect -12287 19038 -12221 19058
rect -12287 13058 -12221 13078
rect -12129 19038 -12063 19058
rect -12129 13058 -12063 13078
rect -11971 19038 -11905 19058
rect -11971 13058 -11905 13078
rect -11813 19038 -11747 19058
rect -11813 13058 -11747 13078
rect -11655 19038 -11589 19058
rect -11655 13058 -11589 13078
rect -11497 19038 -11431 19058
rect -11497 13058 -11431 13078
rect -11339 19038 -11273 19058
rect -11339 13058 -11273 13078
rect -11181 19038 -11115 19058
rect -11181 13058 -11115 13078
rect -11023 19038 -10957 19058
rect -11023 13058 -10957 13078
rect -10865 19038 -10799 19058
rect -10865 13058 -10799 13078
rect -10707 19038 -10641 19058
rect -10707 13058 -10641 13078
rect -10549 19038 -10483 19058
rect -10549 13058 -10483 13078
rect -10391 19038 -10325 19058
rect -10391 13058 -10325 13078
rect -10233 19038 -10167 19058
rect -10233 13058 -10167 13078
rect -10075 19038 -10009 19058
rect -10075 13058 -10009 13078
rect -9917 19038 -9851 19058
rect -9917 13058 -9851 13078
rect -9759 19038 -9693 19058
rect -9759 13058 -9693 13078
rect -9601 19038 -9535 19058
rect -9601 13058 -9535 13078
rect -9443 19038 -9377 19058
rect -9443 13058 -9377 13078
rect -9285 19038 -9219 19058
rect -9285 13058 -9219 13078
rect -9127 19038 -9061 19058
rect -9127 13058 -9061 13078
rect -8969 19038 -8903 19058
rect -8969 13058 -8903 13078
rect -8811 19038 -8745 19058
rect -8811 13058 -8745 13078
rect -8653 19038 -8587 19058
rect -8653 13058 -8587 13078
rect -8495 19038 -8429 19058
rect -8495 13058 -8429 13078
rect -13168 13010 -13148 13026
rect -8514 13010 -8494 13026
rect -13168 12940 -13160 13010
rect -8510 12940 -8494 13010
rect -13168 12926 -13148 12940
rect -8514 12926 -8494 12940
rect -13370 12830 -13300 12900
rect -8290 18900 -7070 19220
rect -8290 18300 -7070 18700
rect -8290 17700 -7070 18100
rect -8290 17100 -7070 17500
rect -8290 16500 -7070 16900
rect -8290 15900 -7070 16300
rect -8290 15300 -7070 15700
rect -8290 14700 -7070 15100
rect -8290 14100 -7070 14500
rect -8290 13500 -7070 13900
rect -8290 12900 -7070 13300
rect -2060 19220 -700 19280
rect -6868 19180 -6848 19190
rect -2214 19180 -2194 19190
rect -6868 19110 -6860 19180
rect -2200 19110 -2194 19180
rect -6868 19090 -6848 19110
rect -2214 19090 -2194 19110
rect -6935 19038 -6869 19058
rect -6935 13058 -6869 13078
rect -6777 19038 -6711 19058
rect -6777 13058 -6711 13078
rect -6619 19038 -6553 19058
rect -6619 13058 -6553 13078
rect -6461 19038 -6395 19058
rect -6461 13058 -6395 13078
rect -6303 19038 -6237 19058
rect -6303 13058 -6237 13078
rect -6145 19038 -6079 19058
rect -6145 13058 -6079 13078
rect -5987 19038 -5921 19058
rect -5987 13058 -5921 13078
rect -5829 19038 -5763 19058
rect -5829 13058 -5763 13078
rect -5671 19038 -5605 19058
rect -5671 13058 -5605 13078
rect -5513 19038 -5447 19058
rect -5513 13058 -5447 13078
rect -5355 19038 -5289 19058
rect -5355 13058 -5289 13078
rect -5197 19038 -5131 19058
rect -5197 13058 -5131 13078
rect -5039 19038 -4973 19058
rect -5039 13058 -4973 13078
rect -4881 19038 -4815 19058
rect -4881 13058 -4815 13078
rect -4723 19038 -4657 19058
rect -4723 13058 -4657 13078
rect -4565 19038 -4499 19058
rect -4565 13058 -4499 13078
rect -4407 19038 -4341 19058
rect -4407 13058 -4341 13078
rect -4249 19038 -4183 19058
rect -4249 13058 -4183 13078
rect -4091 19038 -4025 19058
rect -4091 13058 -4025 13078
rect -3933 19038 -3867 19058
rect -3933 13058 -3867 13078
rect -3775 19038 -3709 19058
rect -3775 13058 -3709 13078
rect -3617 19038 -3551 19058
rect -3617 13058 -3551 13078
rect -3459 19038 -3393 19058
rect -3459 13058 -3393 13078
rect -3301 19038 -3235 19058
rect -3301 13058 -3235 13078
rect -3143 19038 -3077 19058
rect -3143 13058 -3077 13078
rect -2985 19038 -2919 19058
rect -2985 13058 -2919 13078
rect -2827 19038 -2761 19058
rect -2827 13058 -2761 13078
rect -2669 19038 -2603 19058
rect -2669 13058 -2603 13078
rect -2511 19038 -2445 19058
rect -2511 13058 -2445 13078
rect -2353 19038 -2287 19058
rect -2353 13058 -2287 13078
rect -2195 19038 -2129 19058
rect -2195 13058 -2129 13078
rect -6868 13010 -6848 13026
rect -2214 13010 -2194 13026
rect -6868 12940 -6860 13010
rect -2210 12940 -2194 13010
rect -6868 12926 -6848 12940
rect -2214 12926 -2194 12940
rect -8360 12830 -8290 12900
rect -7900 12300 -7400 12900
rect -7070 12830 -7000 12900
rect -1990 19000 -770 19220
rect -1990 18400 -770 18800
rect -1990 17800 -770 18200
rect -1990 17200 -770 17600
rect -1990 16600 -770 17000
rect -1990 16000 -770 16400
rect -1990 15400 -770 15800
rect -1990 14800 -770 15200
rect -1990 14200 -770 14600
rect -1990 13600 -770 14000
rect -1990 13000 -770 13400
rect -2060 12830 -1990 12900
rect -1600 12300 -1100 13000
rect 4240 19220 5600 19280
rect -568 19180 -548 19190
rect 4086 19180 4106 19190
rect -568 19110 -560 19180
rect 4100 19110 4106 19180
rect -568 19090 -548 19110
rect 4086 19090 4106 19110
rect -635 19038 -569 19058
rect -635 13058 -569 13078
rect -477 19038 -411 19058
rect -477 13058 -411 13078
rect -319 19038 -253 19058
rect -319 13058 -253 13078
rect -161 19038 -95 19058
rect -161 13058 -95 13078
rect -3 19038 63 19058
rect -3 13058 63 13078
rect 155 19038 221 19058
rect 155 13058 221 13078
rect 313 19038 379 19058
rect 313 13058 379 13078
rect 471 19038 537 19058
rect 471 13058 537 13078
rect 629 19038 695 19058
rect 629 13058 695 13078
rect 787 19038 853 19058
rect 787 13058 853 13078
rect 945 19038 1011 19058
rect 945 13058 1011 13078
rect 1103 19038 1169 19058
rect 1103 13058 1169 13078
rect 1261 19038 1327 19058
rect 1261 13058 1327 13078
rect 1419 19038 1485 19058
rect 1419 13058 1485 13078
rect 1577 19038 1643 19058
rect 1577 13058 1643 13078
rect 1735 19038 1801 19058
rect 1735 13058 1801 13078
rect 1893 19038 1959 19058
rect 1893 13058 1959 13078
rect 2051 19038 2117 19058
rect 2051 13058 2117 13078
rect 2209 19038 2275 19058
rect 2209 13058 2275 13078
rect 2367 19038 2433 19058
rect 2367 13058 2433 13078
rect 2525 19038 2591 19058
rect 2525 13058 2591 13078
rect 2683 19038 2749 19058
rect 2683 13058 2749 13078
rect 2841 19038 2907 19058
rect 2841 13058 2907 13078
rect 2999 19038 3065 19058
rect 2999 13058 3065 13078
rect 3157 19038 3223 19058
rect 3157 13058 3223 13078
rect 3315 19038 3381 19058
rect 3315 13058 3381 13078
rect 3473 19038 3539 19058
rect 3473 13058 3539 13078
rect 3631 19038 3697 19058
rect 3631 13058 3697 13078
rect 3789 19038 3855 19058
rect 3789 13058 3855 13078
rect 3947 19038 4013 19058
rect 3947 13058 4013 13078
rect 4105 19038 4171 19058
rect 4105 13058 4171 13078
rect -568 13010 -548 13026
rect 4086 13010 4106 13026
rect -568 12940 -560 13010
rect 4090 12940 4106 13010
rect -568 12926 -548 12940
rect 4086 12926 4106 12940
rect -770 12830 -700 12900
rect 4310 18900 5530 19220
rect 4310 18300 5530 18700
rect 4310 17700 5530 18100
rect 4310 17100 5530 17500
rect 4310 16500 5530 16900
rect 4310 15900 5530 16300
rect 4310 15300 5530 15700
rect 4310 14700 5530 15100
rect 4310 14100 5530 14500
rect 4310 13500 5530 13900
rect 4310 12900 5530 13300
rect 10540 19220 10610 19280
rect 5732 19180 5752 19190
rect 10386 19180 10406 19190
rect 5732 19110 5740 19180
rect 10400 19110 10406 19180
rect 5732 19090 5752 19110
rect 10386 19090 10406 19110
rect 5665 19038 5731 19058
rect 5665 13058 5731 13078
rect 5823 19038 5889 19058
rect 5823 13058 5889 13078
rect 5981 19038 6047 19058
rect 5981 13058 6047 13078
rect 6139 19038 6205 19058
rect 6139 13058 6205 13078
rect 6297 19038 6363 19058
rect 6297 13058 6363 13078
rect 6455 19038 6521 19058
rect 6455 13058 6521 13078
rect 6613 19038 6679 19058
rect 6613 13058 6679 13078
rect 6771 19038 6837 19058
rect 6771 13058 6837 13078
rect 6929 19038 6995 19058
rect 6929 13058 6995 13078
rect 7087 19038 7153 19058
rect 7087 13058 7153 13078
rect 7245 19038 7311 19058
rect 7245 13058 7311 13078
rect 7403 19038 7469 19058
rect 7403 13058 7469 13078
rect 7561 19038 7627 19058
rect 7561 13058 7627 13078
rect 7719 19038 7785 19058
rect 7719 13058 7785 13078
rect 7877 19038 7943 19058
rect 7877 13058 7943 13078
rect 8035 19038 8101 19058
rect 8035 13058 8101 13078
rect 8193 19038 8259 19058
rect 8193 13058 8259 13078
rect 8351 19038 8417 19058
rect 8351 13058 8417 13078
rect 8509 19038 8575 19058
rect 8509 13058 8575 13078
rect 8667 19038 8733 19058
rect 8667 13058 8733 13078
rect 8825 19038 8891 19058
rect 8825 13058 8891 13078
rect 8983 19038 9049 19058
rect 8983 13058 9049 13078
rect 9141 19038 9207 19058
rect 9141 13058 9207 13078
rect 9299 19038 9365 19058
rect 9299 13058 9365 13078
rect 9457 19038 9523 19058
rect 9457 13058 9523 13078
rect 9615 19038 9681 19058
rect 9615 13058 9681 13078
rect 9773 19038 9839 19058
rect 9773 13058 9839 13078
rect 9931 19038 9997 19058
rect 9931 13058 9997 13078
rect 10089 19038 10155 19058
rect 10089 13058 10155 13078
rect 10247 19038 10313 19058
rect 10247 13058 10313 13078
rect 10405 19038 10471 19058
rect 10405 13058 10471 13078
rect 5732 13010 5752 13026
rect 10386 13010 10406 13026
rect 5732 12940 5740 13010
rect 10390 12940 10406 13010
rect 5732 12926 5752 12940
rect 10386 12926 10406 12940
rect 4240 12830 4310 12900
rect 4700 12300 5200 12900
rect 5530 12830 5600 12900
rect 10540 12830 10610 12900
rect -8300 12280 -7000 12300
rect -2000 12280 -700 12300
rect 4300 12280 5600 12300
rect -13370 12220 -13300 12280
rect -8360 12220 -7000 12280
rect -13168 12180 -13148 12190
rect -8514 12180 -8494 12190
rect -13168 12110 -13160 12180
rect -8500 12110 -8494 12180
rect -13168 12090 -13148 12110
rect -8514 12090 -8494 12110
rect -13235 12038 -13169 12058
rect -13235 6058 -13169 6078
rect -13077 12038 -13011 12058
rect -13077 6058 -13011 6078
rect -12919 12038 -12853 12058
rect -12919 6058 -12853 6078
rect -12761 12038 -12695 12058
rect -12761 6058 -12695 6078
rect -12603 12038 -12537 12058
rect -12603 6058 -12537 6078
rect -12445 12038 -12379 12058
rect -12445 6058 -12379 6078
rect -12287 12038 -12221 12058
rect -12287 6058 -12221 6078
rect -12129 12038 -12063 12058
rect -12129 6058 -12063 6078
rect -11971 12038 -11905 12058
rect -11971 6058 -11905 6078
rect -11813 12038 -11747 12058
rect -11813 6058 -11747 6078
rect -11655 12038 -11589 12058
rect -11655 6058 -11589 6078
rect -11497 12038 -11431 12058
rect -11497 6058 -11431 6078
rect -11339 12038 -11273 12058
rect -11339 6058 -11273 6078
rect -11181 12038 -11115 12058
rect -11181 6058 -11115 6078
rect -11023 12038 -10957 12058
rect -11023 6058 -10957 6078
rect -10865 12038 -10799 12058
rect -10865 6058 -10799 6078
rect -10707 12038 -10641 12058
rect -10707 6058 -10641 6078
rect -10549 12038 -10483 12058
rect -10549 6058 -10483 6078
rect -10391 12038 -10325 12058
rect -10391 6058 -10325 6078
rect -10233 12038 -10167 12058
rect -10233 6058 -10167 6078
rect -10075 12038 -10009 12058
rect -10075 6058 -10009 6078
rect -9917 12038 -9851 12058
rect -9917 6058 -9851 6078
rect -9759 12038 -9693 12058
rect -9759 6058 -9693 6078
rect -9601 12038 -9535 12058
rect -9601 6058 -9535 6078
rect -9443 12038 -9377 12058
rect -9443 6058 -9377 6078
rect -9285 12038 -9219 12058
rect -9285 6058 -9219 6078
rect -9127 12038 -9061 12058
rect -9127 6058 -9061 6078
rect -8969 12038 -8903 12058
rect -8969 6058 -8903 6078
rect -8811 12038 -8745 12058
rect -8811 6058 -8745 6078
rect -8653 12038 -8587 12058
rect -8653 6058 -8587 6078
rect -8495 12038 -8429 12058
rect -8495 6058 -8429 6078
rect -13168 6010 -13148 6026
rect -8514 6010 -8494 6026
rect -13168 5940 -13160 6010
rect -8510 5940 -8494 6010
rect -13168 5926 -13148 5940
rect -8514 5926 -8494 5940
rect -13370 5830 -13300 5900
rect -8290 11900 -7070 12220
rect -8290 11300 -7070 11700
rect -8290 10700 -7070 11100
rect -8290 10100 -7070 10500
rect -8290 9500 -7070 9900
rect -8290 8900 -7070 9300
rect -8290 8300 -7070 8700
rect -8290 7700 -7070 8100
rect -8290 7100 -7070 7500
rect -8290 6500 -7070 6900
rect -8290 5900 -7070 6300
rect -2060 12220 -700 12280
rect -6868 12180 -6848 12190
rect -2214 12180 -2194 12190
rect -6868 12110 -6860 12180
rect -2200 12110 -2194 12180
rect -6868 12090 -6848 12110
rect -2214 12090 -2194 12110
rect -6935 12038 -6869 12058
rect -6935 6058 -6869 6078
rect -6777 12038 -6711 12058
rect -6777 6058 -6711 6078
rect -6619 12038 -6553 12058
rect -6619 6058 -6553 6078
rect -6461 12038 -6395 12058
rect -6461 6058 -6395 6078
rect -6303 12038 -6237 12058
rect -6303 6058 -6237 6078
rect -6145 12038 -6079 12058
rect -6145 6058 -6079 6078
rect -5987 12038 -5921 12058
rect -5987 6058 -5921 6078
rect -5829 12038 -5763 12058
rect -5829 6058 -5763 6078
rect -5671 12038 -5605 12058
rect -5671 6058 -5605 6078
rect -5513 12038 -5447 12058
rect -5513 6058 -5447 6078
rect -5355 12038 -5289 12058
rect -5355 6058 -5289 6078
rect -5197 12038 -5131 12058
rect -5197 6058 -5131 6078
rect -5039 12038 -4973 12058
rect -5039 6058 -4973 6078
rect -4881 12038 -4815 12058
rect -4881 6058 -4815 6078
rect -4723 12038 -4657 12058
rect -4723 6058 -4657 6078
rect -4565 12038 -4499 12058
rect -4565 6058 -4499 6078
rect -4407 12038 -4341 12058
rect -4407 6058 -4341 6078
rect -4249 12038 -4183 12058
rect -4249 6058 -4183 6078
rect -4091 12038 -4025 12058
rect -4091 6058 -4025 6078
rect -3933 12038 -3867 12058
rect -3933 6058 -3867 6078
rect -3775 12038 -3709 12058
rect -3775 6058 -3709 6078
rect -3617 12038 -3551 12058
rect -3617 6058 -3551 6078
rect -3459 12038 -3393 12058
rect -3459 6058 -3393 6078
rect -3301 12038 -3235 12058
rect -3301 6058 -3235 6078
rect -3143 12038 -3077 12058
rect -3143 6058 -3077 6078
rect -2985 12038 -2919 12058
rect -2985 6058 -2919 6078
rect -2827 12038 -2761 12058
rect -2827 6058 -2761 6078
rect -2669 12038 -2603 12058
rect -2669 6058 -2603 6078
rect -2511 12038 -2445 12058
rect -2511 6058 -2445 6078
rect -2353 12038 -2287 12058
rect -2353 6058 -2287 6078
rect -2195 12038 -2129 12058
rect -2195 6058 -2129 6078
rect -6868 6010 -6848 6026
rect -2214 6010 -2194 6026
rect -6868 5940 -6860 6010
rect -2210 5940 -2194 6010
rect -6868 5926 -6848 5940
rect -2214 5926 -2194 5940
rect -8360 5830 -8290 5900
rect -7070 5830 -7000 5900
rect -1990 11900 -770 12220
rect -1990 11300 -770 11700
rect -1990 10700 -770 11100
rect -1990 10100 -770 10500
rect -1990 9500 -770 9900
rect -1990 8900 -770 9300
rect -1990 8300 -770 8700
rect -1990 7700 -770 8100
rect -1990 7100 -770 7500
rect -1990 6500 -770 6900
rect -1990 5900 -770 6300
rect 4240 12220 5600 12280
rect -568 12180 -548 12190
rect 4086 12180 4106 12190
rect -568 12110 -560 12180
rect 4100 12110 4106 12180
rect -568 12090 -548 12110
rect 4086 12090 4106 12110
rect -635 12038 -569 12058
rect -635 6058 -569 6078
rect -477 12038 -411 12058
rect -477 6058 -411 6078
rect -319 12038 -253 12058
rect -319 6058 -253 6078
rect -161 12038 -95 12058
rect -161 6058 -95 6078
rect -3 12038 63 12058
rect -3 6058 63 6078
rect 155 12038 221 12058
rect 155 6058 221 6078
rect 313 12038 379 12058
rect 313 6058 379 6078
rect 471 12038 537 12058
rect 471 6058 537 6078
rect 629 12038 695 12058
rect 629 6058 695 6078
rect 787 12038 853 12058
rect 787 6058 853 6078
rect 945 12038 1011 12058
rect 945 6058 1011 6078
rect 1103 12038 1169 12058
rect 1103 6058 1169 6078
rect 1261 12038 1327 12058
rect 1261 6058 1327 6078
rect 1419 12038 1485 12058
rect 1419 6058 1485 6078
rect 1577 12038 1643 12058
rect 1577 6058 1643 6078
rect 1735 12038 1801 12058
rect 1735 6058 1801 6078
rect 1893 12038 1959 12058
rect 1893 6058 1959 6078
rect 2051 12038 2117 12058
rect 2051 6058 2117 6078
rect 2209 12038 2275 12058
rect 2209 6058 2275 6078
rect 2367 12038 2433 12058
rect 2367 6058 2433 6078
rect 2525 12038 2591 12058
rect 2525 6058 2591 6078
rect 2683 12038 2749 12058
rect 2683 6058 2749 6078
rect 2841 12038 2907 12058
rect 2841 6058 2907 6078
rect 2999 12038 3065 12058
rect 2999 6058 3065 6078
rect 3157 12038 3223 12058
rect 3157 6058 3223 6078
rect 3315 12038 3381 12058
rect 3315 6058 3381 6078
rect 3473 12038 3539 12058
rect 3473 6058 3539 6078
rect 3631 12038 3697 12058
rect 3631 6058 3697 6078
rect 3789 12038 3855 12058
rect 3789 6058 3855 6078
rect 3947 12038 4013 12058
rect 3947 6058 4013 6078
rect 4105 12038 4171 12058
rect 4105 6058 4171 6078
rect -568 6010 -548 6026
rect 4086 6010 4106 6026
rect -568 5940 -560 6010
rect 4090 5940 4106 6010
rect -568 5926 -548 5940
rect 4086 5926 4106 5940
rect -2060 5830 -1990 5900
rect -770 5830 -700 5900
rect 4310 11900 5530 12220
rect 4310 11300 5530 11700
rect 4310 10700 5530 11100
rect 4310 10100 5530 10500
rect 4310 9500 5530 9900
rect 4310 8900 5530 9300
rect 4310 8300 5530 8700
rect 4310 7700 5530 8100
rect 4310 7100 5530 7500
rect 4310 6500 5530 6900
rect 4310 5900 5530 6300
rect 10540 12220 10610 12280
rect 5732 12180 5752 12190
rect 10386 12180 10406 12190
rect 5732 12110 5740 12180
rect 10400 12110 10406 12180
rect 5732 12090 5752 12110
rect 10386 12090 10406 12110
rect 5665 12038 5731 12058
rect 5665 6058 5731 6078
rect 5823 12038 5889 12058
rect 5823 6058 5889 6078
rect 5981 12038 6047 12058
rect 5981 6058 6047 6078
rect 6139 12038 6205 12058
rect 6139 6058 6205 6078
rect 6297 12038 6363 12058
rect 6297 6058 6363 6078
rect 6455 12038 6521 12058
rect 6455 6058 6521 6078
rect 6613 12038 6679 12058
rect 6613 6058 6679 6078
rect 6771 12038 6837 12058
rect 6771 6058 6837 6078
rect 6929 12038 6995 12058
rect 6929 6058 6995 6078
rect 7087 12038 7153 12058
rect 7087 6058 7153 6078
rect 7245 12038 7311 12058
rect 7245 6058 7311 6078
rect 7403 12038 7469 12058
rect 7403 6058 7469 6078
rect 7561 12038 7627 12058
rect 7561 6058 7627 6078
rect 7719 12038 7785 12058
rect 7719 6058 7785 6078
rect 7877 12038 7943 12058
rect 7877 6058 7943 6078
rect 8035 12038 8101 12058
rect 8035 6058 8101 6078
rect 8193 12038 8259 12058
rect 8193 6058 8259 6078
rect 8351 12038 8417 12058
rect 8351 6058 8417 6078
rect 8509 12038 8575 12058
rect 8509 6058 8575 6078
rect 8667 12038 8733 12058
rect 8667 6058 8733 6078
rect 8825 12038 8891 12058
rect 8825 6058 8891 6078
rect 8983 12038 9049 12058
rect 8983 6058 9049 6078
rect 9141 12038 9207 12058
rect 9141 6058 9207 6078
rect 9299 12038 9365 12058
rect 9299 6058 9365 6078
rect 9457 12038 9523 12058
rect 9457 6058 9523 6078
rect 9615 12038 9681 12058
rect 9615 6058 9681 6078
rect 9773 12038 9839 12058
rect 9773 6058 9839 6078
rect 9931 12038 9997 12058
rect 9931 6058 9997 6078
rect 10089 12038 10155 12058
rect 10089 6058 10155 6078
rect 10247 12038 10313 12058
rect 10247 6058 10313 6078
rect 10405 12038 10471 12058
rect 10405 6058 10471 6078
rect 5732 6010 5752 6026
rect 10386 6010 10406 6026
rect 5732 5940 5740 6010
rect 10390 5940 10406 6010
rect 5732 5926 5752 5940
rect 10386 5926 10406 5940
rect 4240 5830 4310 5900
rect 5530 5830 5600 5900
rect 10540 5830 10610 5900
<< via2 >>
rect -13160 49710 -13148 49780
rect -13148 49710 -8514 49780
rect -8514 49710 -8500 49780
rect -13235 44285 -13169 46045
rect -13077 47285 -13011 49045
rect -12919 44285 -12853 46045
rect -12761 47285 -12695 49045
rect -12603 44285 -12537 46045
rect -12445 47285 -12379 49045
rect -12287 44285 -12221 46045
rect -12129 47285 -12063 49045
rect -11971 44285 -11905 46045
rect -11813 47285 -11747 49045
rect -11655 44285 -11589 46045
rect -11497 47285 -11431 49045
rect -11339 44285 -11273 46045
rect -11181 47285 -11115 49045
rect -11023 44285 -10957 46045
rect -10865 47285 -10799 49045
rect -10707 44285 -10641 46045
rect -10549 47285 -10483 49045
rect -10391 44285 -10325 46045
rect -10233 47285 -10167 49045
rect -10075 44285 -10009 46045
rect -9917 47285 -9851 49045
rect -9759 44285 -9693 46045
rect -9601 47285 -9535 49045
rect -9443 44285 -9377 46045
rect -9285 47285 -9219 49045
rect -9127 44285 -9061 46045
rect -8969 47285 -8903 49045
rect -8811 44285 -8745 46045
rect -8653 47285 -8587 49045
rect -8495 44285 -8429 46045
rect -13160 43540 -13148 43610
rect -13148 43540 -8514 43610
rect -8514 43540 -8510 43610
rect -6860 49710 -6848 49780
rect -6848 49710 -2214 49780
rect -2214 49710 -2200 49780
rect -6935 44285 -6869 46045
rect -6777 47285 -6711 49045
rect -6619 44285 -6553 46045
rect -6461 47285 -6395 49045
rect -6303 44285 -6237 46045
rect -6145 47285 -6079 49045
rect -5987 44285 -5921 46045
rect -5829 47285 -5763 49045
rect -5671 44285 -5605 46045
rect -5513 47285 -5447 49045
rect -5355 44285 -5289 46045
rect -5197 47285 -5131 49045
rect -5039 44285 -4973 46045
rect -4881 47285 -4815 49045
rect -4723 44285 -4657 46045
rect -4565 47285 -4499 49045
rect -4407 44285 -4341 46045
rect -4249 47285 -4183 49045
rect -4091 44285 -4025 46045
rect -3933 47285 -3867 49045
rect -3775 44285 -3709 46045
rect -3617 47285 -3551 49045
rect -3459 44285 -3393 46045
rect -3301 47285 -3235 49045
rect -3143 44285 -3077 46045
rect -2985 47285 -2919 49045
rect -2827 44285 -2761 46045
rect -2669 47285 -2603 49045
rect -2511 44285 -2445 46045
rect -2353 47285 -2287 49045
rect -2195 44285 -2129 46045
rect -6860 43540 -6848 43610
rect -6848 43540 -2214 43610
rect -2214 43540 -2210 43610
rect -560 49710 -548 49780
rect -548 49710 4086 49780
rect 4086 49710 4100 49780
rect -635 44285 -569 46045
rect -477 47285 -411 49045
rect -319 44285 -253 46045
rect -161 47285 -95 49045
rect -3 44285 63 46045
rect 155 47285 221 49045
rect 313 44285 379 46045
rect 471 47285 537 49045
rect 629 44285 695 46045
rect 787 47285 853 49045
rect 945 44285 1011 46045
rect 1103 47285 1169 49045
rect 1261 44285 1327 46045
rect 1419 47285 1485 49045
rect 1577 44285 1643 46045
rect 1735 47285 1801 49045
rect 1893 44285 1959 46045
rect 2051 47285 2117 49045
rect 2209 44285 2275 46045
rect 2367 47285 2433 49045
rect 2525 44285 2591 46045
rect 2683 47285 2749 49045
rect 2841 44285 2907 46045
rect 2999 47285 3065 49045
rect 3157 44285 3223 46045
rect 3315 47285 3381 49045
rect 3473 44285 3539 46045
rect 3631 47285 3697 49045
rect 3789 44285 3855 46045
rect 3947 47285 4013 49045
rect 4105 44285 4171 46045
rect -560 43540 -548 43610
rect -548 43540 4086 43610
rect 4086 43540 4090 43610
rect 5740 49710 5752 49780
rect 5752 49710 10386 49780
rect 10386 49710 10400 49780
rect 5665 44285 5731 46045
rect 5823 47285 5889 49045
rect 5981 44285 6047 46045
rect 6139 47285 6205 49045
rect 6297 44285 6363 46045
rect 6455 47285 6521 49045
rect 6613 44285 6679 46045
rect 6771 47285 6837 49045
rect 6929 44285 6995 46045
rect 7087 47285 7153 49045
rect 7245 44285 7311 46045
rect 7403 47285 7469 49045
rect 7561 44285 7627 46045
rect 7719 47285 7785 49045
rect 7877 44285 7943 46045
rect 8035 47285 8101 49045
rect 8193 44285 8259 46045
rect 8351 47285 8417 49045
rect 8509 44285 8575 46045
rect 8667 47285 8733 49045
rect 8825 44285 8891 46045
rect 8983 47285 9049 49045
rect 9141 44285 9207 46045
rect 9299 47285 9365 49045
rect 9457 44285 9523 46045
rect 9615 47285 9681 49045
rect 9773 44285 9839 46045
rect 9931 47285 9997 49045
rect 10089 44285 10155 46045
rect 10247 47285 10313 49045
rect 10405 44285 10471 46045
rect 5740 43540 5752 43610
rect 5752 43540 10386 43610
rect 10386 43540 10390 43610
rect -13160 42710 -13148 42780
rect -13148 42710 -8514 42780
rect -8514 42710 -8500 42780
rect -13235 37285 -13169 39045
rect -13077 40285 -13011 42045
rect -12919 37285 -12853 39045
rect -12761 40285 -12695 42045
rect -12603 37285 -12537 39045
rect -12445 40285 -12379 42045
rect -12287 37285 -12221 39045
rect -12129 40285 -12063 42045
rect -11971 37285 -11905 39045
rect -11813 40285 -11747 42045
rect -11655 37285 -11589 39045
rect -11497 40285 -11431 42045
rect -11339 37285 -11273 39045
rect -11181 40285 -11115 42045
rect -11023 37285 -10957 39045
rect -10865 40285 -10799 42045
rect -10707 37285 -10641 39045
rect -10549 40285 -10483 42045
rect -10391 37285 -10325 39045
rect -10233 40285 -10167 42045
rect -10075 37285 -10009 39045
rect -9917 40285 -9851 42045
rect -9759 37285 -9693 39045
rect -9601 40285 -9535 42045
rect -9443 37285 -9377 39045
rect -9285 40285 -9219 42045
rect -9127 37285 -9061 39045
rect -8969 40285 -8903 42045
rect -8811 37285 -8745 39045
rect -8653 40285 -8587 42045
rect -8495 37285 -8429 39045
rect -13160 36540 -13148 36610
rect -13148 36540 -8514 36610
rect -8514 36540 -8510 36610
rect -6860 42710 -6848 42780
rect -6848 42710 -2214 42780
rect -2214 42710 -2200 42780
rect -6935 37285 -6869 39045
rect -6777 40285 -6711 42045
rect -6619 37285 -6553 39045
rect -6461 40285 -6395 42045
rect -6303 37285 -6237 39045
rect -6145 40285 -6079 42045
rect -5987 37285 -5921 39045
rect -5829 40285 -5763 42045
rect -5671 37285 -5605 39045
rect -5513 40285 -5447 42045
rect -5355 37285 -5289 39045
rect -5197 40285 -5131 42045
rect -5039 37285 -4973 39045
rect -4881 40285 -4815 42045
rect -4723 37285 -4657 39045
rect -4565 40285 -4499 42045
rect -4407 37285 -4341 39045
rect -4249 40285 -4183 42045
rect -4091 37285 -4025 39045
rect -3933 40285 -3867 42045
rect -3775 37285 -3709 39045
rect -3617 40285 -3551 42045
rect -3459 37285 -3393 39045
rect -3301 40285 -3235 42045
rect -3143 37285 -3077 39045
rect -2985 40285 -2919 42045
rect -2827 37285 -2761 39045
rect -2669 40285 -2603 42045
rect -2511 37285 -2445 39045
rect -2353 40285 -2287 42045
rect -2195 37285 -2129 39045
rect -6860 36540 -6848 36610
rect -6848 36540 -2214 36610
rect -2214 36540 -2210 36610
rect -560 42710 -548 42780
rect -548 42710 4086 42780
rect 4086 42710 4100 42780
rect -635 37285 -569 39045
rect -477 40285 -411 42045
rect -319 37285 -253 39045
rect -161 40285 -95 42045
rect -3 37285 63 39045
rect 155 40285 221 42045
rect 313 37285 379 39045
rect 471 40285 537 42045
rect 629 37285 695 39045
rect 787 40285 853 42045
rect 945 37285 1011 39045
rect 1103 40285 1169 42045
rect 1261 37285 1327 39045
rect 1419 40285 1485 42045
rect 1577 37285 1643 39045
rect 1735 40285 1801 42045
rect 1893 37285 1959 39045
rect 2051 40285 2117 42045
rect 2209 37285 2275 39045
rect 2367 40285 2433 42045
rect 2525 37285 2591 39045
rect 2683 40285 2749 42045
rect 2841 37285 2907 39045
rect 2999 40285 3065 42045
rect 3157 37285 3223 39045
rect 3315 40285 3381 42045
rect 3473 37285 3539 39045
rect 3631 40285 3697 42045
rect 3789 37285 3855 39045
rect 3947 40285 4013 42045
rect 4105 37285 4171 39045
rect -560 36540 -548 36610
rect -548 36540 4086 36610
rect 4086 36540 4090 36610
rect 5740 42710 5752 42780
rect 5752 42710 10386 42780
rect 10386 42710 10400 42780
rect 5665 37285 5731 39045
rect 5823 40285 5889 42045
rect 5981 37285 6047 39045
rect 6139 40285 6205 42045
rect 6297 37285 6363 39045
rect 6455 40285 6521 42045
rect 6613 37285 6679 39045
rect 6771 40285 6837 42045
rect 6929 37285 6995 39045
rect 7087 40285 7153 42045
rect 7245 37285 7311 39045
rect 7403 40285 7469 42045
rect 7561 37285 7627 39045
rect 7719 40285 7785 42045
rect 7877 37285 7943 39045
rect 8035 40285 8101 42045
rect 8193 37285 8259 39045
rect 8351 40285 8417 42045
rect 8509 37285 8575 39045
rect 8667 40285 8733 42045
rect 8825 37285 8891 39045
rect 8983 40285 9049 42045
rect 9141 37285 9207 39045
rect 9299 40285 9365 42045
rect 9457 37285 9523 39045
rect 9615 40285 9681 42045
rect 9773 37285 9839 39045
rect 9931 40285 9997 42045
rect 10089 37285 10155 39045
rect 10247 40285 10313 42045
rect 10405 37285 10471 39045
rect 5740 36540 5752 36610
rect 5752 36540 10386 36610
rect 10386 36540 10390 36610
rect -13160 34410 -13148 34480
rect -13148 34410 -8514 34480
rect -8514 34410 -8500 34480
rect -13235 28985 -13169 30745
rect -13077 31985 -13011 33745
rect -12919 28985 -12853 30745
rect -12761 31985 -12695 33745
rect -12603 28985 -12537 30745
rect -12445 31985 -12379 33745
rect -12287 28985 -12221 30745
rect -12129 31985 -12063 33745
rect -11971 28985 -11905 30745
rect -11813 31985 -11747 33745
rect -11655 28985 -11589 30745
rect -11497 31985 -11431 33745
rect -11339 28985 -11273 30745
rect -11181 31985 -11115 33745
rect -11023 28985 -10957 30745
rect -10865 31985 -10799 33745
rect -10707 28985 -10641 30745
rect -10549 31985 -10483 33745
rect -10391 28985 -10325 30745
rect -10233 31985 -10167 33745
rect -10075 28985 -10009 30745
rect -9917 31985 -9851 33745
rect -9759 28985 -9693 30745
rect -9601 31985 -9535 33745
rect -9443 28985 -9377 30745
rect -9285 31985 -9219 33745
rect -9127 28985 -9061 30745
rect -8969 31985 -8903 33745
rect -8811 28985 -8745 30745
rect -8653 31985 -8587 33745
rect -8495 28985 -8429 30745
rect -13160 28240 -13148 28310
rect -13148 28240 -8514 28310
rect -8514 28240 -8510 28310
rect -6860 34410 -6848 34480
rect -6848 34410 -2214 34480
rect -2214 34410 -2200 34480
rect -6935 28985 -6869 30745
rect -6777 31985 -6711 33745
rect -6619 28985 -6553 30745
rect -6461 31985 -6395 33745
rect -6303 28985 -6237 30745
rect -6145 31985 -6079 33745
rect -5987 28985 -5921 30745
rect -5829 31985 -5763 33745
rect -5671 28985 -5605 30745
rect -5513 31985 -5447 33745
rect -5355 28985 -5289 30745
rect -5197 31985 -5131 33745
rect -5039 28985 -4973 30745
rect -4881 31985 -4815 33745
rect -4723 28985 -4657 30745
rect -4565 31985 -4499 33745
rect -4407 28985 -4341 30745
rect -4249 31985 -4183 33745
rect -4091 28985 -4025 30745
rect -3933 31985 -3867 33745
rect -3775 28985 -3709 30745
rect -3617 31985 -3551 33745
rect -3459 28985 -3393 30745
rect -3301 31985 -3235 33745
rect -3143 28985 -3077 30745
rect -2985 31985 -2919 33745
rect -2827 28985 -2761 30745
rect -2669 31985 -2603 33745
rect -2511 28985 -2445 30745
rect -2353 31985 -2287 33745
rect -2195 28985 -2129 30745
rect -6860 28240 -6848 28310
rect -6848 28240 -2214 28310
rect -2214 28240 -2210 28310
rect -560 34410 -548 34480
rect -548 34410 4086 34480
rect 4086 34410 4100 34480
rect -635 28985 -569 30745
rect -477 31985 -411 33745
rect -319 28985 -253 30745
rect -161 31985 -95 33745
rect -3 28985 63 30745
rect 155 31985 221 33745
rect 313 28985 379 30745
rect 471 31985 537 33745
rect 629 28985 695 30745
rect 787 31985 853 33745
rect 945 28985 1011 30745
rect 1103 31985 1169 33745
rect 1261 28985 1327 30745
rect 1419 31985 1485 33745
rect 1577 28985 1643 30745
rect 1735 31985 1801 33745
rect 1893 28985 1959 30745
rect 2051 31985 2117 33745
rect 2209 28985 2275 30745
rect 2367 31985 2433 33745
rect 2525 28985 2591 30745
rect 2683 31985 2749 33745
rect 2841 28985 2907 30745
rect 2999 31985 3065 33745
rect 3157 28985 3223 30745
rect 3315 31985 3381 33745
rect 3473 28985 3539 30745
rect 3631 31985 3697 33745
rect 3789 28985 3855 30745
rect 3947 31985 4013 33745
rect 4105 28985 4171 30745
rect -560 28240 -548 28310
rect -548 28240 4086 28310
rect 4086 28240 4090 28310
rect 5740 34410 5752 34480
rect 5752 34410 10386 34480
rect 10386 34410 10400 34480
rect 5665 28985 5731 30745
rect 5823 31985 5889 33745
rect 5981 28985 6047 30745
rect 6139 31985 6205 33745
rect 6297 28985 6363 30745
rect 6455 31985 6521 33745
rect 6613 28985 6679 30745
rect 6771 31985 6837 33745
rect 6929 28985 6995 30745
rect 7087 31985 7153 33745
rect 7245 28985 7311 30745
rect 7403 31985 7469 33745
rect 7561 28985 7627 30745
rect 7719 31985 7785 33745
rect 7877 28985 7943 30745
rect 8035 31985 8101 33745
rect 8193 28985 8259 30745
rect 8351 31985 8417 33745
rect 8509 28985 8575 30745
rect 8667 31985 8733 33745
rect 8825 28985 8891 30745
rect 8983 31985 9049 33745
rect 9141 28985 9207 30745
rect 9299 31985 9365 33745
rect 9457 28985 9523 30745
rect 9615 31985 9681 33745
rect 9773 28985 9839 30745
rect 9931 31985 9997 33745
rect 10089 28985 10155 30745
rect 10247 31985 10313 33745
rect 10405 28985 10471 30745
rect 5740 28240 5752 28310
rect 5752 28240 10386 28310
rect 10386 28240 10390 28310
rect -13160 27410 -13148 27480
rect -13148 27410 -8514 27480
rect -8514 27410 -8500 27480
rect -13235 21985 -13169 23745
rect -13077 24985 -13011 26745
rect -12919 21985 -12853 23745
rect -12761 24985 -12695 26745
rect -12603 21985 -12537 23745
rect -12445 24985 -12379 26745
rect -12287 21985 -12221 23745
rect -12129 24985 -12063 26745
rect -11971 21985 -11905 23745
rect -11813 24985 -11747 26745
rect -11655 21985 -11589 23745
rect -11497 24985 -11431 26745
rect -11339 21985 -11273 23745
rect -11181 24985 -11115 26745
rect -11023 21985 -10957 23745
rect -10865 24985 -10799 26745
rect -10707 21985 -10641 23745
rect -10549 24985 -10483 26745
rect -10391 21985 -10325 23745
rect -10233 24985 -10167 26745
rect -10075 21985 -10009 23745
rect -9917 24985 -9851 26745
rect -9759 21985 -9693 23745
rect -9601 24985 -9535 26745
rect -9443 21985 -9377 23745
rect -9285 24985 -9219 26745
rect -9127 21985 -9061 23745
rect -8969 24985 -8903 26745
rect -8811 21985 -8745 23745
rect -8653 24985 -8587 26745
rect -8495 21985 -8429 23745
rect -13160 21240 -13148 21310
rect -13148 21240 -8514 21310
rect -8514 21240 -8510 21310
rect -6860 27410 -6848 27480
rect -6848 27410 -2214 27480
rect -2214 27410 -2200 27480
rect -6935 21985 -6869 23745
rect -6777 24985 -6711 26745
rect -6619 21985 -6553 23745
rect -6461 24985 -6395 26745
rect -6303 21985 -6237 23745
rect -6145 24985 -6079 26745
rect -5987 21985 -5921 23745
rect -5829 24985 -5763 26745
rect -5671 21985 -5605 23745
rect -5513 24985 -5447 26745
rect -5355 21985 -5289 23745
rect -5197 24985 -5131 26745
rect -5039 21985 -4973 23745
rect -4881 24985 -4815 26745
rect -4723 21985 -4657 23745
rect -4565 24985 -4499 26745
rect -4407 21985 -4341 23745
rect -4249 24985 -4183 26745
rect -4091 21985 -4025 23745
rect -3933 24985 -3867 26745
rect -3775 21985 -3709 23745
rect -3617 24985 -3551 26745
rect -3459 21985 -3393 23745
rect -3301 24985 -3235 26745
rect -3143 21985 -3077 23745
rect -2985 24985 -2919 26745
rect -2827 21985 -2761 23745
rect -2669 24985 -2603 26745
rect -2511 21985 -2445 23745
rect -2353 24985 -2287 26745
rect -2195 21985 -2129 23745
rect -6860 21240 -6848 21310
rect -6848 21240 -2214 21310
rect -2214 21240 -2210 21310
rect -560 27410 -548 27480
rect -548 27410 4086 27480
rect 4086 27410 4100 27480
rect -635 21985 -569 23745
rect -477 24985 -411 26745
rect -319 21985 -253 23745
rect -161 24985 -95 26745
rect -3 21985 63 23745
rect 155 24985 221 26745
rect 313 21985 379 23745
rect 471 24985 537 26745
rect 629 21985 695 23745
rect 787 24985 853 26745
rect 945 21985 1011 23745
rect 1103 24985 1169 26745
rect 1261 21985 1327 23745
rect 1419 24985 1485 26745
rect 1577 21985 1643 23745
rect 1735 24985 1801 26745
rect 1893 21985 1959 23745
rect 2051 24985 2117 26745
rect 2209 21985 2275 23745
rect 2367 24985 2433 26745
rect 2525 21985 2591 23745
rect 2683 24985 2749 26745
rect 2841 21985 2907 23745
rect 2999 24985 3065 26745
rect 3157 21985 3223 23745
rect 3315 24985 3381 26745
rect 3473 21985 3539 23745
rect 3631 24985 3697 26745
rect 3789 21985 3855 23745
rect 3947 24985 4013 26745
rect 4105 21985 4171 23745
rect -560 21240 -548 21310
rect -548 21240 4086 21310
rect 4086 21240 4090 21310
rect 5740 27410 5752 27480
rect 5752 27410 10386 27480
rect 10386 27410 10400 27480
rect 5665 21985 5731 23745
rect 5823 24985 5889 26745
rect 5981 21985 6047 23745
rect 6139 24985 6205 26745
rect 6297 21985 6363 23745
rect 6455 24985 6521 26745
rect 6613 21985 6679 23745
rect 6771 24985 6837 26745
rect 6929 21985 6995 23745
rect 7087 24985 7153 26745
rect 7245 21985 7311 23745
rect 7403 24985 7469 26745
rect 7561 21985 7627 23745
rect 7719 24985 7785 26745
rect 7877 21985 7943 23745
rect 8035 24985 8101 26745
rect 8193 21985 8259 23745
rect 8351 24985 8417 26745
rect 8509 21985 8575 23745
rect 8667 24985 8733 26745
rect 8825 21985 8891 23745
rect 8983 24985 9049 26745
rect 9141 21985 9207 23745
rect 9299 24985 9365 26745
rect 9457 21985 9523 23745
rect 9615 24985 9681 26745
rect 9773 21985 9839 23745
rect 9931 24985 9997 26745
rect 10089 21985 10155 23745
rect 10247 24985 10313 26745
rect 10405 21985 10471 23745
rect 5740 21240 5752 21310
rect 5752 21240 10386 21310
rect 10386 21240 10390 21310
rect -13160 19110 -13148 19180
rect -13148 19110 -8514 19180
rect -8514 19110 -8500 19180
rect -13235 13685 -13169 15445
rect -13077 16685 -13011 18445
rect -12919 13685 -12853 15445
rect -12761 16685 -12695 18445
rect -12603 13685 -12537 15445
rect -12445 16685 -12379 18445
rect -12287 13685 -12221 15445
rect -12129 16685 -12063 18445
rect -11971 13685 -11905 15445
rect -11813 16685 -11747 18445
rect -11655 13685 -11589 15445
rect -11497 16685 -11431 18445
rect -11339 13685 -11273 15445
rect -11181 16685 -11115 18445
rect -11023 13685 -10957 15445
rect -10865 16685 -10799 18445
rect -10707 13685 -10641 15445
rect -10549 16685 -10483 18445
rect -10391 13685 -10325 15445
rect -10233 16685 -10167 18445
rect -10075 13685 -10009 15445
rect -9917 16685 -9851 18445
rect -9759 13685 -9693 15445
rect -9601 16685 -9535 18445
rect -9443 13685 -9377 15445
rect -9285 16685 -9219 18445
rect -9127 13685 -9061 15445
rect -8969 16685 -8903 18445
rect -8811 13685 -8745 15445
rect -8653 16685 -8587 18445
rect -8495 13685 -8429 15445
rect -13160 12940 -13148 13010
rect -13148 12940 -8514 13010
rect -8514 12940 -8510 13010
rect -6860 19110 -6848 19180
rect -6848 19110 -2214 19180
rect -2214 19110 -2200 19180
rect -6935 13685 -6869 15445
rect -6777 16685 -6711 18445
rect -6619 13685 -6553 15445
rect -6461 16685 -6395 18445
rect -6303 13685 -6237 15445
rect -6145 16685 -6079 18445
rect -5987 13685 -5921 15445
rect -5829 16685 -5763 18445
rect -5671 13685 -5605 15445
rect -5513 16685 -5447 18445
rect -5355 13685 -5289 15445
rect -5197 16685 -5131 18445
rect -5039 13685 -4973 15445
rect -4881 16685 -4815 18445
rect -4723 13685 -4657 15445
rect -4565 16685 -4499 18445
rect -4407 13685 -4341 15445
rect -4249 16685 -4183 18445
rect -4091 13685 -4025 15445
rect -3933 16685 -3867 18445
rect -3775 13685 -3709 15445
rect -3617 16685 -3551 18445
rect -3459 13685 -3393 15445
rect -3301 16685 -3235 18445
rect -3143 13685 -3077 15445
rect -2985 16685 -2919 18445
rect -2827 13685 -2761 15445
rect -2669 16685 -2603 18445
rect -2511 13685 -2445 15445
rect -2353 16685 -2287 18445
rect -2195 13685 -2129 15445
rect -6860 12940 -6848 13010
rect -6848 12940 -2214 13010
rect -2214 12940 -2210 13010
rect -560 19110 -548 19180
rect -548 19110 4086 19180
rect 4086 19110 4100 19180
rect -635 13685 -569 15445
rect -477 16685 -411 18445
rect -319 13685 -253 15445
rect -161 16685 -95 18445
rect -3 13685 63 15445
rect 155 16685 221 18445
rect 313 13685 379 15445
rect 471 16685 537 18445
rect 629 13685 695 15445
rect 787 16685 853 18445
rect 945 13685 1011 15445
rect 1103 16685 1169 18445
rect 1261 13685 1327 15445
rect 1419 16685 1485 18445
rect 1577 13685 1643 15445
rect 1735 16685 1801 18445
rect 1893 13685 1959 15445
rect 2051 16685 2117 18445
rect 2209 13685 2275 15445
rect 2367 16685 2433 18445
rect 2525 13685 2591 15445
rect 2683 16685 2749 18445
rect 2841 13685 2907 15445
rect 2999 16685 3065 18445
rect 3157 13685 3223 15445
rect 3315 16685 3381 18445
rect 3473 13685 3539 15445
rect 3631 16685 3697 18445
rect 3789 13685 3855 15445
rect 3947 16685 4013 18445
rect 4105 13685 4171 15445
rect -560 12940 -548 13010
rect -548 12940 4086 13010
rect 4086 12940 4090 13010
rect 5740 19110 5752 19180
rect 5752 19110 10386 19180
rect 10386 19110 10400 19180
rect 5665 13685 5731 15445
rect 5823 16685 5889 18445
rect 5981 13685 6047 15445
rect 6139 16685 6205 18445
rect 6297 13685 6363 15445
rect 6455 16685 6521 18445
rect 6613 13685 6679 15445
rect 6771 16685 6837 18445
rect 6929 13685 6995 15445
rect 7087 16685 7153 18445
rect 7245 13685 7311 15445
rect 7403 16685 7469 18445
rect 7561 13685 7627 15445
rect 7719 16685 7785 18445
rect 7877 13685 7943 15445
rect 8035 16685 8101 18445
rect 8193 13685 8259 15445
rect 8351 16685 8417 18445
rect 8509 13685 8575 15445
rect 8667 16685 8733 18445
rect 8825 13685 8891 15445
rect 8983 16685 9049 18445
rect 9141 13685 9207 15445
rect 9299 16685 9365 18445
rect 9457 13685 9523 15445
rect 9615 16685 9681 18445
rect 9773 13685 9839 15445
rect 9931 16685 9997 18445
rect 10089 13685 10155 15445
rect 10247 16685 10313 18445
rect 10405 13685 10471 15445
rect 5740 12940 5752 13010
rect 5752 12940 10386 13010
rect 10386 12940 10390 13010
rect -13160 12110 -13148 12180
rect -13148 12110 -8514 12180
rect -8514 12110 -8500 12180
rect -13235 6685 -13169 8445
rect -13077 9685 -13011 11445
rect -12919 6685 -12853 8445
rect -12761 9685 -12695 11445
rect -12603 6685 -12537 8445
rect -12445 9685 -12379 11445
rect -12287 6685 -12221 8445
rect -12129 9685 -12063 11445
rect -11971 6685 -11905 8445
rect -11813 9685 -11747 11445
rect -11655 6685 -11589 8445
rect -11497 9685 -11431 11445
rect -11339 6685 -11273 8445
rect -11181 9685 -11115 11445
rect -11023 6685 -10957 8445
rect -10865 9685 -10799 11445
rect -10707 6685 -10641 8445
rect -10549 9685 -10483 11445
rect -10391 6685 -10325 8445
rect -10233 9685 -10167 11445
rect -10075 6685 -10009 8445
rect -9917 9685 -9851 11445
rect -9759 6685 -9693 8445
rect -9601 9685 -9535 11445
rect -9443 6685 -9377 8445
rect -9285 9685 -9219 11445
rect -9127 6685 -9061 8445
rect -8969 9685 -8903 11445
rect -8811 6685 -8745 8445
rect -8653 9685 -8587 11445
rect -8495 6685 -8429 8445
rect -13160 5940 -13148 6010
rect -13148 5940 -8514 6010
rect -8514 5940 -8510 6010
rect -6860 12110 -6848 12180
rect -6848 12110 -2214 12180
rect -2214 12110 -2200 12180
rect -6935 6685 -6869 8445
rect -6777 9685 -6711 11445
rect -6619 6685 -6553 8445
rect -6461 9685 -6395 11445
rect -6303 6685 -6237 8445
rect -6145 9685 -6079 11445
rect -5987 6685 -5921 8445
rect -5829 9685 -5763 11445
rect -5671 6685 -5605 8445
rect -5513 9685 -5447 11445
rect -5355 6685 -5289 8445
rect -5197 9685 -5131 11445
rect -5039 6685 -4973 8445
rect -4881 9685 -4815 11445
rect -4723 6685 -4657 8445
rect -4565 9685 -4499 11445
rect -4407 6685 -4341 8445
rect -4249 9685 -4183 11445
rect -4091 6685 -4025 8445
rect -3933 9685 -3867 11445
rect -3775 6685 -3709 8445
rect -3617 9685 -3551 11445
rect -3459 6685 -3393 8445
rect -3301 9685 -3235 11445
rect -3143 6685 -3077 8445
rect -2985 9685 -2919 11445
rect -2827 6685 -2761 8445
rect -2669 9685 -2603 11445
rect -2511 6685 -2445 8445
rect -2353 9685 -2287 11445
rect -2195 6685 -2129 8445
rect -6860 5940 -6848 6010
rect -6848 5940 -2214 6010
rect -2214 5940 -2210 6010
rect -560 12110 -548 12180
rect -548 12110 4086 12180
rect 4086 12110 4100 12180
rect -635 6685 -569 8445
rect -477 9685 -411 11445
rect -319 6685 -253 8445
rect -161 9685 -95 11445
rect -3 6685 63 8445
rect 155 9685 221 11445
rect 313 6685 379 8445
rect 471 9685 537 11445
rect 629 6685 695 8445
rect 787 9685 853 11445
rect 945 6685 1011 8445
rect 1103 9685 1169 11445
rect 1261 6685 1327 8445
rect 1419 9685 1485 11445
rect 1577 6685 1643 8445
rect 1735 9685 1801 11445
rect 1893 6685 1959 8445
rect 2051 9685 2117 11445
rect 2209 6685 2275 8445
rect 2367 9685 2433 11445
rect 2525 6685 2591 8445
rect 2683 9685 2749 11445
rect 2841 6685 2907 8445
rect 2999 9685 3065 11445
rect 3157 6685 3223 8445
rect 3315 9685 3381 11445
rect 3473 6685 3539 8445
rect 3631 9685 3697 11445
rect 3789 6685 3855 8445
rect 3947 9685 4013 11445
rect 4105 6685 4171 8445
rect -560 5940 -548 6010
rect -548 5940 4086 6010
rect 4086 5940 4090 6010
rect 5740 12110 5752 12180
rect 5752 12110 10386 12180
rect 10386 12110 10400 12180
rect 5665 6685 5731 8445
rect 5823 9685 5889 11445
rect 5981 6685 6047 8445
rect 6139 9685 6205 11445
rect 6297 6685 6363 8445
rect 6455 9685 6521 11445
rect 6613 6685 6679 8445
rect 6771 9685 6837 11445
rect 6929 6685 6995 8445
rect 7087 9685 7153 11445
rect 7245 6685 7311 8445
rect 7403 9685 7469 11445
rect 7561 6685 7627 8445
rect 7719 9685 7785 11445
rect 7877 6685 7943 8445
rect 8035 9685 8101 11445
rect 8193 6685 8259 8445
rect 8351 9685 8417 11445
rect 8509 6685 8575 8445
rect 8667 9685 8733 11445
rect 8825 6685 8891 8445
rect 8983 9685 9049 11445
rect 9141 6685 9207 8445
rect 9299 9685 9365 11445
rect 9457 6685 9523 8445
rect 9615 9685 9681 11445
rect 9773 6685 9839 8445
rect 9931 9685 9997 11445
rect 10089 6685 10155 8445
rect 10247 9685 10313 11445
rect 10405 6685 10471 8445
rect 5740 5940 5752 6010
rect 5752 5940 10386 6010
rect 10386 5940 10390 6010
<< metal3 >>
rect -13300 49780 -8300 49900
rect -13300 49710 -13160 49780
rect -8500 49710 -8300 49780
rect -13300 49700 -8300 49710
rect -7000 49780 -2000 49900
rect -7000 49710 -6860 49780
rect -2200 49710 -2000 49780
rect -7000 49700 -2000 49710
rect -700 49780 4300 49900
rect -700 49710 -560 49780
rect 4100 49710 4300 49780
rect -700 49700 4300 49710
rect 5600 49780 10600 49900
rect 5600 49710 5740 49780
rect 10400 49710 10600 49780
rect 5600 49700 10600 49710
rect -13400 49100 -8290 49200
rect -13400 47300 -13300 49100
rect -12000 49045 -8290 49100
rect -12000 47300 -11813 49045
rect -13400 47285 -13077 47300
rect -13011 47285 -12761 47300
rect -12695 47285 -12445 47300
rect -12379 47285 -12129 47300
rect -12063 47285 -11813 47300
rect -11747 47285 -11497 49045
rect -11431 47285 -11181 49045
rect -11115 47285 -10865 49045
rect -10799 47285 -10549 49045
rect -10483 47285 -10233 49045
rect -10167 47285 -9917 49045
rect -9851 47285 -9601 49045
rect -9535 47285 -9285 49045
rect -9219 47285 -8969 49045
rect -8903 47285 -8653 49045
rect -8587 47285 -8290 49045
rect -13400 47200 -8290 47285
rect -7100 49100 -1990 49200
rect -7100 47300 -7000 49100
rect -5800 49045 -1990 49100
rect -7100 47285 -6777 47300
rect -6711 47285 -6461 47300
rect -6395 47285 -6145 47300
rect -6079 47285 -5829 47300
rect -5763 47285 -5513 49045
rect -5447 47285 -5197 49045
rect -5131 47285 -4881 49045
rect -4815 47285 -4565 49045
rect -4499 47285 -4249 49045
rect -4183 47285 -3933 49045
rect -3867 47285 -3617 49045
rect -3551 47285 -3301 49045
rect -3235 47285 -2985 49045
rect -2919 47285 -2669 49045
rect -2603 47285 -2353 49045
rect -2287 47285 -1990 49045
rect -7100 47200 -1990 47285
rect -800 49100 4310 49200
rect -800 47300 -700 49100
rect 600 49045 4310 49100
rect 600 47300 787 49045
rect -800 47285 -477 47300
rect -411 47285 -161 47300
rect -95 47285 155 47300
rect 221 47285 471 47300
rect 537 47285 787 47300
rect 853 47285 1103 49045
rect 1169 47285 1419 49045
rect 1485 47285 1735 49045
rect 1801 47285 2051 49045
rect 2117 47285 2367 49045
rect 2433 47285 2683 49045
rect 2749 47285 2999 49045
rect 3065 47285 3315 49045
rect 3381 47285 3631 49045
rect 3697 47285 3947 49045
rect 4013 47285 4310 49045
rect -800 47200 4310 47285
rect 5500 49100 10610 49200
rect 5500 47300 5600 49100
rect 6800 49045 10610 49100
rect 5500 47285 5823 47300
rect 5889 47285 6139 47300
rect 6205 47285 6455 47300
rect 6521 47285 6771 47300
rect 6837 47285 7087 49045
rect 7153 47285 7403 49045
rect 7469 47285 7719 49045
rect 7785 47285 8035 49045
rect 8101 47285 8351 49045
rect 8417 47285 8667 49045
rect 8733 47285 8983 49045
rect 9049 47285 9299 49045
rect 9365 47285 9615 49045
rect 9681 47285 9931 49045
rect 9997 47285 10247 49045
rect 10313 47285 10610 49045
rect 5500 47200 10610 47285
rect -13400 46100 -8290 46200
rect -13400 44300 -13300 46100
rect -12000 46045 -8290 46100
rect -12000 44300 -11971 46045
rect -13400 44285 -13235 44300
rect -13169 44285 -12919 44300
rect -12853 44285 -12603 44300
rect -12537 44285 -12287 44300
rect -12221 44285 -11971 44300
rect -11905 44285 -11655 46045
rect -11589 44285 -11339 46045
rect -11273 44285 -11023 46045
rect -10957 44285 -10707 46045
rect -10641 44285 -10391 46045
rect -10325 44285 -10075 46045
rect -10009 44285 -9759 46045
rect -9693 44285 -9443 46045
rect -9377 44285 -9127 46045
rect -9061 44285 -8811 46045
rect -8745 44285 -8495 46045
rect -8429 44285 -8290 46045
rect -13400 44200 -8290 44285
rect -7070 46100 -1800 46200
rect -7070 46045 -3200 46100
rect -7070 44285 -6935 46045
rect -6869 44285 -6619 46045
rect -6553 44285 -6303 46045
rect -6237 44285 -5987 46045
rect -5921 44285 -5671 46045
rect -5605 44285 -5355 46045
rect -5289 44285 -5039 46045
rect -4973 44285 -4723 46045
rect -4657 44285 -4407 46045
rect -4341 44285 -4091 46045
rect -4025 44285 -3775 46045
rect -3709 44285 -3459 46045
rect -3393 44300 -3200 46045
rect -1900 44300 -1800 46100
rect -3393 44285 -3143 44300
rect -3077 44285 -2827 44300
rect -2761 44285 -2511 44300
rect -2445 44285 -2195 44300
rect -2129 44285 -1800 44300
rect -7070 44200 -1800 44285
rect -800 46100 4310 46200
rect -800 44300 -700 46100
rect 600 46045 4310 46100
rect 600 44300 629 46045
rect -800 44285 -635 44300
rect -569 44285 -319 44300
rect -253 44285 -3 44300
rect 63 44285 313 44300
rect 379 44285 629 44300
rect 695 44285 945 46045
rect 1011 44285 1261 46045
rect 1327 44285 1577 46045
rect 1643 44285 1893 46045
rect 1959 44285 2209 46045
rect 2275 44285 2525 46045
rect 2591 44285 2841 46045
rect 2907 44285 3157 46045
rect 3223 44285 3473 46045
rect 3539 44285 3789 46045
rect 3855 44285 4105 46045
rect 4171 44285 4310 46045
rect -800 44200 4310 44285
rect 5530 46100 10800 46200
rect 5530 46045 9400 46100
rect 5530 44285 5665 46045
rect 5731 44285 5981 46045
rect 6047 44285 6297 46045
rect 6363 44285 6613 46045
rect 6679 44285 6929 46045
rect 6995 44285 7245 46045
rect 7311 44285 7561 46045
rect 7627 44285 7877 46045
rect 7943 44285 8193 46045
rect 8259 44285 8509 46045
rect 8575 44285 8825 46045
rect 8891 44285 9141 46045
rect 9207 44300 9400 46045
rect 10700 44300 10800 46100
rect 9207 44285 9457 44300
rect 9523 44285 9773 44300
rect 9839 44285 10089 44300
rect 10155 44285 10405 44300
rect 10471 44285 10800 44300
rect 5530 44200 10800 44285
rect -11700 43800 -9800 43900
rect -11700 43700 -11500 43800
rect -13400 43610 -11500 43700
rect -10000 43700 -9800 43800
rect 900 43800 2800 43900
rect 900 43700 1100 43800
rect -10000 43610 -7400 43700
rect -13400 43540 -13160 43610
rect -8510 43580 -7400 43610
rect -8510 43540 -7780 43580
rect -13400 43500 -11500 43540
rect -10000 43500 -7780 43540
rect -13400 43420 -7780 43500
rect -7420 43420 -7400 43580
rect -13400 43400 -7400 43420
rect -7200 43610 -1100 43700
rect -7200 43540 -6860 43610
rect -2210 43580 -1100 43610
rect -2210 43540 -1480 43580
rect -7200 43420 -1480 43540
rect -1120 43420 -1100 43580
rect -7200 43400 -1100 43420
rect -900 43610 1100 43700
rect 2600 43700 2800 43800
rect 2600 43610 5200 43700
rect -900 43540 -560 43610
rect 4090 43580 5200 43610
rect 4090 43540 4820 43580
rect -900 43500 1100 43540
rect 2600 43500 4820 43540
rect -900 43420 4820 43500
rect 5180 43420 5200 43580
rect -900 43400 5200 43420
rect 5400 43610 10600 43700
rect 5400 43540 5740 43610
rect 10390 43540 10600 43610
rect 5400 43400 10600 43540
rect -7200 43200 -6900 43400
rect -5400 43300 -2800 43400
rect -900 43300 -700 43400
rect 5400 43300 5700 43400
rect 7200 43300 9800 43400
rect -8300 43000 -6900 43200
rect -2000 43100 -700 43300
rect 4300 43100 5700 43300
rect -11700 42900 -9800 43000
rect -8300 42900 -8000 43000
rect -5400 42900 -2800 43000
rect -2000 42900 -1700 43100
rect 900 42900 2800 43000
rect 4300 42900 4600 43100
rect 7200 42900 9800 43000
rect -13400 42780 -11500 42900
rect -10000 42780 -8000 42900
rect -13400 42710 -13160 42780
rect -8500 42710 -8000 42780
rect -13400 42600 -11500 42710
rect -10000 42600 -8000 42710
rect -7800 42880 -1700 42900
rect -7800 42720 -7780 42880
rect -7420 42780 -1700 42880
rect -7420 42720 -6860 42780
rect -7800 42710 -6860 42720
rect -2200 42710 -1700 42780
rect -7800 42600 -1700 42710
rect -1500 42880 1100 42900
rect -1500 42720 -1480 42880
rect -1120 42780 1100 42880
rect 2600 42780 4600 42900
rect -1120 42720 -560 42780
rect -1500 42710 -560 42720
rect 4100 42710 4600 42780
rect -1500 42600 1100 42710
rect 2600 42600 4600 42710
rect 4800 42880 10600 42900
rect 4800 42720 4820 42880
rect 5180 42780 10600 42880
rect 5180 42720 5740 42780
rect 4800 42710 5740 42720
rect 10400 42710 10600 42780
rect 4800 42600 10600 42710
rect -11700 42500 -9800 42600
rect 900 42500 2800 42600
rect -13370 42100 -8290 42200
rect -13370 42045 -11400 42100
rect -10100 42045 -8290 42100
rect -13370 40285 -13077 42045
rect -13011 40285 -12761 42045
rect -12695 40285 -12445 42045
rect -12379 40285 -12129 42045
rect -12063 40285 -11813 42045
rect -11747 40285 -11497 42045
rect -11431 40300 -11400 42045
rect -10100 40300 -9917 42045
rect -11431 40285 -11181 40300
rect -11115 40285 -10865 40300
rect -10799 40285 -10549 40300
rect -10483 40285 -10233 40300
rect -10167 40285 -9917 40300
rect -9851 40285 -9601 42045
rect -9535 40285 -9285 42045
rect -9219 40285 -8969 42045
rect -8903 40285 -8653 42045
rect -8587 40285 -8290 42045
rect -13370 40200 -8290 40285
rect -7100 42100 -1990 42200
rect -7100 40300 -7000 42100
rect -5700 42045 -1990 42100
rect -5700 40300 -5513 42045
rect -7100 40285 -6777 40300
rect -6711 40285 -6461 40300
rect -6395 40285 -6145 40300
rect -6079 40285 -5829 40300
rect -5763 40285 -5513 40300
rect -5447 40285 -5197 42045
rect -5131 40285 -4881 42045
rect -4815 40285 -4565 42045
rect -4499 40285 -4249 42045
rect -4183 40285 -3933 42045
rect -3867 40285 -3617 42045
rect -3551 40285 -3301 42045
rect -3235 40285 -2985 42045
rect -2919 40285 -2669 42045
rect -2603 40285 -2353 42045
rect -2287 40285 -1990 42045
rect -7100 40200 -1990 40285
rect -770 42100 4310 42200
rect -770 42045 1200 42100
rect 2500 42045 4310 42100
rect -770 40285 -477 42045
rect -411 40285 -161 42045
rect -95 40285 155 42045
rect 221 40285 471 42045
rect 537 40285 787 42045
rect 853 40285 1103 42045
rect 1169 40300 1200 42045
rect 2500 40300 2683 42045
rect 1169 40285 1419 40300
rect 1485 40285 1735 40300
rect 1801 40285 2051 40300
rect 2117 40285 2367 40300
rect 2433 40285 2683 40300
rect 2749 40285 2999 42045
rect 3065 40285 3315 42045
rect 3381 40285 3631 42045
rect 3697 40285 3947 42045
rect 4013 40285 4310 42045
rect -770 40200 4310 40285
rect 5500 42100 10610 42200
rect 5500 40300 5600 42100
rect 6900 42045 10610 42100
rect 6900 40300 7087 42045
rect 5500 40285 5823 40300
rect 5889 40285 6139 40300
rect 6205 40285 6455 40300
rect 6521 40285 6771 40300
rect 6837 40285 7087 40300
rect 7153 40285 7403 42045
rect 7469 40285 7719 42045
rect 7785 40285 8035 42045
rect 8101 40285 8351 42045
rect 8417 40285 8667 42045
rect 8733 40285 8983 42045
rect 9049 40285 9299 42045
rect 9365 40285 9615 42045
rect 9681 40285 9931 42045
rect 9997 40285 10247 42045
rect 10313 40285 10610 42045
rect 5500 40200 10610 40285
rect -13370 39100 -8100 39200
rect -13370 39045 -9500 39100
rect -13370 37285 -13235 39045
rect -13169 37285 -12919 39045
rect -12853 37285 -12603 39045
rect -12537 37285 -12287 39045
rect -12221 37285 -11971 39045
rect -11905 37285 -11655 39045
rect -11589 37285 -11339 39045
rect -11273 37285 -11023 39045
rect -10957 37285 -10707 39045
rect -10641 37285 -10391 39045
rect -10325 37285 -10075 39045
rect -10009 37285 -9759 39045
rect -9693 37300 -9500 39045
rect -8200 37300 -8100 39100
rect -9693 37285 -9443 37300
rect -9377 37285 -9127 37300
rect -9061 37285 -8811 37300
rect -8745 37285 -8495 37300
rect -8429 37285 -8100 37300
rect -13370 37200 -8100 37285
rect -7070 39100 -1990 39200
rect -7070 39045 -5100 39100
rect -3800 39045 -1990 39100
rect -7070 37285 -6935 39045
rect -6869 37285 -6619 39045
rect -6553 37285 -6303 39045
rect -6237 37285 -5987 39045
rect -5921 37285 -5671 39045
rect -5605 37285 -5355 39045
rect -5289 37300 -5100 39045
rect -3800 37300 -3775 39045
rect -5289 37285 -5039 37300
rect -4973 37285 -4723 37300
rect -4657 37285 -4407 37300
rect -4341 37285 -4091 37300
rect -4025 37285 -3775 37300
rect -3709 37285 -3459 39045
rect -3393 37285 -3143 39045
rect -3077 37285 -2827 39045
rect -2761 37285 -2511 39045
rect -2445 37285 -2195 39045
rect -2129 37285 -1990 39045
rect -7070 37200 -1990 37285
rect -770 39100 4500 39200
rect -770 39045 3100 39100
rect -770 37285 -635 39045
rect -569 37285 -319 39045
rect -253 37285 -3 39045
rect 63 37285 313 39045
rect 379 37285 629 39045
rect 695 37285 945 39045
rect 1011 37285 1261 39045
rect 1327 37285 1577 39045
rect 1643 37285 1893 39045
rect 1959 37285 2209 39045
rect 2275 37285 2525 39045
rect 2591 37285 2841 39045
rect 2907 37300 3100 39045
rect 4400 37300 4500 39100
rect 2907 37285 3157 37300
rect 3223 37285 3473 37300
rect 3539 37285 3789 37300
rect 3855 37285 4105 37300
rect 4171 37285 4500 37300
rect -770 37200 4500 37285
rect 5500 39100 10800 39200
rect 5500 39045 7500 39100
rect 8800 39045 10800 39100
rect 5500 37285 5665 39045
rect 5731 37285 5981 39045
rect 6047 37285 6297 39045
rect 6363 37285 6613 39045
rect 6679 37285 6929 39045
rect 6995 37285 7245 39045
rect 7311 37300 7500 39045
rect 8800 37300 8825 39045
rect 7311 37285 7561 37300
rect 7627 37285 7877 37300
rect 7943 37285 8193 37300
rect 8259 37285 8509 37300
rect 8575 37285 8825 37300
rect 8891 37285 9141 39045
rect 9207 37285 9457 39045
rect 9523 37285 9773 39045
rect 9839 37285 10089 39045
rect 10155 37285 10405 39045
rect 10471 37285 10800 39045
rect 5500 37200 10800 37285
rect -13300 36610 -8300 36630
rect -13300 36540 -13160 36610
rect -8510 36540 -8300 36610
rect -13300 36430 -8300 36540
rect -7000 36610 -2000 36630
rect -7000 36540 -6860 36610
rect -2210 36540 -2000 36610
rect -7000 36430 -2000 36540
rect -700 36610 4300 36630
rect -700 36540 -560 36610
rect 4090 36540 4300 36610
rect -700 36430 4300 36540
rect 5600 36610 10600 36630
rect 5600 36540 5740 36610
rect 10390 36540 10600 36610
rect 5600 36430 10600 36540
rect -13300 34480 -8300 34600
rect -13300 34410 -13160 34480
rect -8500 34410 -8300 34480
rect -13300 34400 -8300 34410
rect -7000 34480 -2000 34600
rect -7000 34410 -6860 34480
rect -2200 34410 -2000 34480
rect -7000 34400 -2000 34410
rect -700 34480 4300 34600
rect -700 34410 -560 34480
rect 4100 34410 4300 34480
rect -700 34400 4300 34410
rect 5600 34480 10600 34600
rect 5600 34410 5740 34480
rect 10400 34410 10600 34480
rect 5600 34400 10600 34410
rect -13400 33800 -8290 33900
rect -13400 32000 -13300 33800
rect -12000 33745 -8290 33800
rect -12000 32000 -11813 33745
rect -13400 31985 -13077 32000
rect -13011 31985 -12761 32000
rect -12695 31985 -12445 32000
rect -12379 31985 -12129 32000
rect -12063 31985 -11813 32000
rect -11747 31985 -11497 33745
rect -11431 31985 -11181 33745
rect -11115 31985 -10865 33745
rect -10799 31985 -10549 33745
rect -10483 31985 -10233 33745
rect -10167 31985 -9917 33745
rect -9851 31985 -9601 33745
rect -9535 31985 -9285 33745
rect -9219 31985 -8969 33745
rect -8903 31985 -8653 33745
rect -8587 31985 -8290 33745
rect -13400 31900 -8290 31985
rect -7100 33800 -1990 33900
rect -7100 32000 -7000 33800
rect -5800 33745 -1990 33800
rect -7100 31985 -6777 32000
rect -6711 31985 -6461 32000
rect -6395 31985 -6145 32000
rect -6079 31985 -5829 32000
rect -5763 31985 -5513 33745
rect -5447 31985 -5197 33745
rect -5131 31985 -4881 33745
rect -4815 31985 -4565 33745
rect -4499 31985 -4249 33745
rect -4183 31985 -3933 33745
rect -3867 31985 -3617 33745
rect -3551 31985 -3301 33745
rect -3235 31985 -2985 33745
rect -2919 31985 -2669 33745
rect -2603 31985 -2353 33745
rect -2287 31985 -1990 33745
rect -7100 31900 -1990 31985
rect -800 33800 4310 33900
rect -800 32000 -700 33800
rect 600 33745 4310 33800
rect 600 32000 787 33745
rect -800 31985 -477 32000
rect -411 31985 -161 32000
rect -95 31985 155 32000
rect 221 31985 471 32000
rect 537 31985 787 32000
rect 853 31985 1103 33745
rect 1169 31985 1419 33745
rect 1485 31985 1735 33745
rect 1801 31985 2051 33745
rect 2117 31985 2367 33745
rect 2433 31985 2683 33745
rect 2749 31985 2999 33745
rect 3065 31985 3315 33745
rect 3381 31985 3631 33745
rect 3697 31985 3947 33745
rect 4013 31985 4310 33745
rect -800 31900 4310 31985
rect 5500 33800 10610 33900
rect 5500 32000 5600 33800
rect 6800 33745 10610 33800
rect 5500 31985 5823 32000
rect 5889 31985 6139 32000
rect 6205 31985 6455 32000
rect 6521 31985 6771 32000
rect 6837 31985 7087 33745
rect 7153 31985 7403 33745
rect 7469 31985 7719 33745
rect 7785 31985 8035 33745
rect 8101 31985 8351 33745
rect 8417 31985 8667 33745
rect 8733 31985 8983 33745
rect 9049 31985 9299 33745
rect 9365 31985 9615 33745
rect 9681 31985 9931 33745
rect 9997 31985 10247 33745
rect 10313 31985 10610 33745
rect 5500 31900 10610 31985
rect -13400 30800 -8290 30900
rect -13400 29000 -13300 30800
rect -12000 30745 -8290 30800
rect -12000 29000 -11971 30745
rect -13400 28985 -13235 29000
rect -13169 28985 -12919 29000
rect -12853 28985 -12603 29000
rect -12537 28985 -12287 29000
rect -12221 28985 -11971 29000
rect -11905 28985 -11655 30745
rect -11589 28985 -11339 30745
rect -11273 28985 -11023 30745
rect -10957 28985 -10707 30745
rect -10641 28985 -10391 30745
rect -10325 28985 -10075 30745
rect -10009 28985 -9759 30745
rect -9693 28985 -9443 30745
rect -9377 28985 -9127 30745
rect -9061 28985 -8811 30745
rect -8745 28985 -8495 30745
rect -8429 28985 -8290 30745
rect -13400 28900 -8290 28985
rect -7070 30800 -1800 30900
rect -7070 30745 -3200 30800
rect -7070 28985 -6935 30745
rect -6869 28985 -6619 30745
rect -6553 28985 -6303 30745
rect -6237 28985 -5987 30745
rect -5921 28985 -5671 30745
rect -5605 28985 -5355 30745
rect -5289 28985 -5039 30745
rect -4973 28985 -4723 30745
rect -4657 28985 -4407 30745
rect -4341 28985 -4091 30745
rect -4025 28985 -3775 30745
rect -3709 28985 -3459 30745
rect -3393 29000 -3200 30745
rect -1900 29000 -1800 30800
rect -3393 28985 -3143 29000
rect -3077 28985 -2827 29000
rect -2761 28985 -2511 29000
rect -2445 28985 -2195 29000
rect -2129 28985 -1800 29000
rect -7070 28900 -1800 28985
rect -800 30800 4310 30900
rect -800 29000 -700 30800
rect 600 30745 4310 30800
rect 600 29000 629 30745
rect -800 28985 -635 29000
rect -569 28985 -319 29000
rect -253 28985 -3 29000
rect 63 28985 313 29000
rect 379 28985 629 29000
rect 695 28985 945 30745
rect 1011 28985 1261 30745
rect 1327 28985 1577 30745
rect 1643 28985 1893 30745
rect 1959 28985 2209 30745
rect 2275 28985 2525 30745
rect 2591 28985 2841 30745
rect 2907 28985 3157 30745
rect 3223 28985 3473 30745
rect 3539 28985 3789 30745
rect 3855 28985 4105 30745
rect 4171 28985 4310 30745
rect -800 28900 4310 28985
rect 5530 30800 10800 30900
rect 5530 30745 9400 30800
rect 5530 28985 5665 30745
rect 5731 28985 5981 30745
rect 6047 28985 6297 30745
rect 6363 28985 6613 30745
rect 6679 28985 6929 30745
rect 6995 28985 7245 30745
rect 7311 28985 7561 30745
rect 7627 28985 7877 30745
rect 7943 28985 8193 30745
rect 8259 28985 8509 30745
rect 8575 28985 8825 30745
rect 8891 28985 9141 30745
rect 9207 29000 9400 30745
rect 10700 29000 10800 30800
rect 9207 28985 9457 29000
rect 9523 28985 9773 29000
rect 9839 28985 10089 29000
rect 10155 28985 10405 29000
rect 10471 28985 10800 29000
rect 5530 28900 10800 28985
rect -11700 28500 -9800 28600
rect -11700 28400 -11500 28500
rect -13400 28310 -11500 28400
rect -10000 28400 -9800 28500
rect 900 28500 2800 28600
rect 900 28400 1100 28500
rect -10000 28310 -7400 28400
rect -13400 28240 -13160 28310
rect -8510 28280 -7400 28310
rect -8510 28240 -7780 28280
rect -13400 28200 -11500 28240
rect -10000 28200 -7780 28240
rect -13400 28120 -7780 28200
rect -7420 28120 -7400 28280
rect -13400 28100 -7400 28120
rect -7200 28310 -1100 28400
rect -7200 28240 -6860 28310
rect -2210 28280 -1100 28310
rect -2210 28240 -1480 28280
rect -7200 28120 -1480 28240
rect -1120 28120 -1100 28280
rect -7200 28100 -1100 28120
rect -900 28310 1100 28400
rect 2600 28400 2800 28500
rect 2600 28310 5200 28400
rect -900 28240 -560 28310
rect 4090 28280 5200 28310
rect 4090 28240 4820 28280
rect -900 28200 1100 28240
rect 2600 28200 4820 28240
rect -900 28120 4820 28200
rect 5180 28120 5200 28280
rect -900 28100 5200 28120
rect 5400 28310 10600 28400
rect 5400 28240 5740 28310
rect 10390 28240 10600 28310
rect 5400 28100 10600 28240
rect -7200 27900 -6900 28100
rect -5400 28000 -2800 28100
rect -900 28000 -700 28100
rect 5400 28000 5700 28100
rect 7200 28000 9800 28100
rect -8300 27700 -6900 27900
rect -2000 27800 -700 28000
rect 4300 27800 5700 28000
rect -11700 27600 -9800 27700
rect -8300 27600 -8000 27700
rect -5400 27600 -2800 27700
rect -2000 27600 -1700 27800
rect 900 27600 2800 27700
rect 4300 27600 4600 27800
rect 7200 27600 9800 27700
rect -13400 27480 -11500 27600
rect -10000 27480 -8000 27600
rect -13400 27410 -13160 27480
rect -8500 27410 -8000 27480
rect -13400 27300 -11500 27410
rect -10000 27300 -8000 27410
rect -7800 27580 -1700 27600
rect -7800 27420 -7780 27580
rect -7420 27480 -1700 27580
rect -7420 27420 -6860 27480
rect -7800 27410 -6860 27420
rect -2200 27410 -1700 27480
rect -7800 27300 -1700 27410
rect -1500 27580 1100 27600
rect -1500 27420 -1480 27580
rect -1120 27480 1100 27580
rect 2600 27480 4600 27600
rect -1120 27420 -560 27480
rect -1500 27410 -560 27420
rect 4100 27410 4600 27480
rect -1500 27300 1100 27410
rect 2600 27300 4600 27410
rect 4800 27580 10600 27600
rect 4800 27420 4820 27580
rect 5180 27480 10600 27580
rect 5180 27420 5740 27480
rect 4800 27410 5740 27420
rect 10400 27410 10600 27480
rect 4800 27300 10600 27410
rect -11700 27200 -9800 27300
rect 900 27200 2800 27300
rect -13370 26800 -8290 26900
rect -13370 26745 -11400 26800
rect -10100 26745 -8290 26800
rect -13370 24985 -13077 26745
rect -13011 24985 -12761 26745
rect -12695 24985 -12445 26745
rect -12379 24985 -12129 26745
rect -12063 24985 -11813 26745
rect -11747 24985 -11497 26745
rect -11431 25000 -11400 26745
rect -10100 25000 -9917 26745
rect -11431 24985 -11181 25000
rect -11115 24985 -10865 25000
rect -10799 24985 -10549 25000
rect -10483 24985 -10233 25000
rect -10167 24985 -9917 25000
rect -9851 24985 -9601 26745
rect -9535 24985 -9285 26745
rect -9219 24985 -8969 26745
rect -8903 24985 -8653 26745
rect -8587 24985 -8290 26745
rect -13370 24900 -8290 24985
rect -7100 26800 -1990 26900
rect -7100 25000 -7000 26800
rect -5700 26745 -1990 26800
rect -5700 25000 -5513 26745
rect -7100 24985 -6777 25000
rect -6711 24985 -6461 25000
rect -6395 24985 -6145 25000
rect -6079 24985 -5829 25000
rect -5763 24985 -5513 25000
rect -5447 24985 -5197 26745
rect -5131 24985 -4881 26745
rect -4815 24985 -4565 26745
rect -4499 24985 -4249 26745
rect -4183 24985 -3933 26745
rect -3867 24985 -3617 26745
rect -3551 24985 -3301 26745
rect -3235 24985 -2985 26745
rect -2919 24985 -2669 26745
rect -2603 24985 -2353 26745
rect -2287 24985 -1990 26745
rect -7100 24900 -1990 24985
rect -770 26800 4310 26900
rect -770 26745 1200 26800
rect 2500 26745 4310 26800
rect -770 24985 -477 26745
rect -411 24985 -161 26745
rect -95 24985 155 26745
rect 221 24985 471 26745
rect 537 24985 787 26745
rect 853 24985 1103 26745
rect 1169 25000 1200 26745
rect 2500 25000 2683 26745
rect 1169 24985 1419 25000
rect 1485 24985 1735 25000
rect 1801 24985 2051 25000
rect 2117 24985 2367 25000
rect 2433 24985 2683 25000
rect 2749 24985 2999 26745
rect 3065 24985 3315 26745
rect 3381 24985 3631 26745
rect 3697 24985 3947 26745
rect 4013 24985 4310 26745
rect -770 24900 4310 24985
rect 5500 26800 10610 26900
rect 5500 25000 5600 26800
rect 6900 26745 10610 26800
rect 6900 25000 7087 26745
rect 5500 24985 5823 25000
rect 5889 24985 6139 25000
rect 6205 24985 6455 25000
rect 6521 24985 6771 25000
rect 6837 24985 7087 25000
rect 7153 24985 7403 26745
rect 7469 24985 7719 26745
rect 7785 24985 8035 26745
rect 8101 24985 8351 26745
rect 8417 24985 8667 26745
rect 8733 24985 8983 26745
rect 9049 24985 9299 26745
rect 9365 24985 9615 26745
rect 9681 24985 9931 26745
rect 9997 24985 10247 26745
rect 10313 24985 10610 26745
rect 5500 24900 10610 24985
rect -13370 23800 -8100 23900
rect -13370 23745 -9500 23800
rect -13370 21985 -13235 23745
rect -13169 21985 -12919 23745
rect -12853 21985 -12603 23745
rect -12537 21985 -12287 23745
rect -12221 21985 -11971 23745
rect -11905 21985 -11655 23745
rect -11589 21985 -11339 23745
rect -11273 21985 -11023 23745
rect -10957 21985 -10707 23745
rect -10641 21985 -10391 23745
rect -10325 21985 -10075 23745
rect -10009 21985 -9759 23745
rect -9693 22000 -9500 23745
rect -8200 22000 -8100 23800
rect -9693 21985 -9443 22000
rect -9377 21985 -9127 22000
rect -9061 21985 -8811 22000
rect -8745 21985 -8495 22000
rect -8429 21985 -8100 22000
rect -13370 21900 -8100 21985
rect -7070 23800 -1990 23900
rect -7070 23745 -5100 23800
rect -3800 23745 -1990 23800
rect -7070 21985 -6935 23745
rect -6869 21985 -6619 23745
rect -6553 21985 -6303 23745
rect -6237 21985 -5987 23745
rect -5921 21985 -5671 23745
rect -5605 21985 -5355 23745
rect -5289 22000 -5100 23745
rect -3800 22000 -3775 23745
rect -5289 21985 -5039 22000
rect -4973 21985 -4723 22000
rect -4657 21985 -4407 22000
rect -4341 21985 -4091 22000
rect -4025 21985 -3775 22000
rect -3709 21985 -3459 23745
rect -3393 21985 -3143 23745
rect -3077 21985 -2827 23745
rect -2761 21985 -2511 23745
rect -2445 21985 -2195 23745
rect -2129 21985 -1990 23745
rect -7070 21900 -1990 21985
rect -770 23800 4500 23900
rect -770 23745 3100 23800
rect -770 21985 -635 23745
rect -569 21985 -319 23745
rect -253 21985 -3 23745
rect 63 21985 313 23745
rect 379 21985 629 23745
rect 695 21985 945 23745
rect 1011 21985 1261 23745
rect 1327 21985 1577 23745
rect 1643 21985 1893 23745
rect 1959 21985 2209 23745
rect 2275 21985 2525 23745
rect 2591 21985 2841 23745
rect 2907 22000 3100 23745
rect 4400 22000 4500 23800
rect 2907 21985 3157 22000
rect 3223 21985 3473 22000
rect 3539 21985 3789 22000
rect 3855 21985 4105 22000
rect 4171 21985 4500 22000
rect -770 21900 4500 21985
rect 5500 23800 10800 23900
rect 5500 23745 7500 23800
rect 8800 23745 10800 23800
rect 5500 21985 5665 23745
rect 5731 21985 5981 23745
rect 6047 21985 6297 23745
rect 6363 21985 6613 23745
rect 6679 21985 6929 23745
rect 6995 21985 7245 23745
rect 7311 22000 7500 23745
rect 8800 22000 8825 23745
rect 7311 21985 7561 22000
rect 7627 21985 7877 22000
rect 7943 21985 8193 22000
rect 8259 21985 8509 22000
rect 8575 21985 8825 22000
rect 8891 21985 9141 23745
rect 9207 21985 9457 23745
rect 9523 21985 9773 23745
rect 9839 21985 10089 23745
rect 10155 21985 10405 23745
rect 10471 21985 10800 23745
rect 5500 21900 10800 21985
rect -13300 21310 -8300 21330
rect -13300 21240 -13160 21310
rect -8510 21240 -8300 21310
rect -13300 21130 -8300 21240
rect -7000 21310 -2000 21330
rect -7000 21240 -6860 21310
rect -2210 21240 -2000 21310
rect -7000 21130 -2000 21240
rect -700 21310 4300 21330
rect -700 21240 -560 21310
rect 4090 21240 4300 21310
rect -700 21130 4300 21240
rect 5600 21310 10600 21330
rect 5600 21240 5740 21310
rect 10390 21240 10600 21310
rect 5600 21130 10600 21240
rect -13300 19180 -8300 19300
rect -13300 19110 -13160 19180
rect -8500 19110 -8300 19180
rect -13300 19100 -8300 19110
rect -7000 19180 -2000 19300
rect -7000 19110 -6860 19180
rect -2200 19110 -2000 19180
rect -7000 19100 -2000 19110
rect -700 19180 4300 19300
rect -700 19110 -560 19180
rect 4100 19110 4300 19180
rect -700 19100 4300 19110
rect 5600 19180 10600 19300
rect 5600 19110 5740 19180
rect 10400 19110 10600 19180
rect 5600 19100 10600 19110
rect -13400 18500 -8290 18600
rect -13400 16700 -13300 18500
rect -12000 18445 -8290 18500
rect -12000 16700 -11813 18445
rect -13400 16685 -13077 16700
rect -13011 16685 -12761 16700
rect -12695 16685 -12445 16700
rect -12379 16685 -12129 16700
rect -12063 16685 -11813 16700
rect -11747 16685 -11497 18445
rect -11431 16685 -11181 18445
rect -11115 16685 -10865 18445
rect -10799 16685 -10549 18445
rect -10483 16685 -10233 18445
rect -10167 16685 -9917 18445
rect -9851 16685 -9601 18445
rect -9535 16685 -9285 18445
rect -9219 16685 -8969 18445
rect -8903 16685 -8653 18445
rect -8587 16685 -8290 18445
rect -13400 16600 -8290 16685
rect -7100 18500 -1990 18600
rect -7100 16700 -7000 18500
rect -5800 18445 -1990 18500
rect -7100 16685 -6777 16700
rect -6711 16685 -6461 16700
rect -6395 16685 -6145 16700
rect -6079 16685 -5829 16700
rect -5763 16685 -5513 18445
rect -5447 16685 -5197 18445
rect -5131 16685 -4881 18445
rect -4815 16685 -4565 18445
rect -4499 16685 -4249 18445
rect -4183 16685 -3933 18445
rect -3867 16685 -3617 18445
rect -3551 16685 -3301 18445
rect -3235 16685 -2985 18445
rect -2919 16685 -2669 18445
rect -2603 16685 -2353 18445
rect -2287 16685 -1990 18445
rect -7100 16600 -1990 16685
rect -800 18500 4310 18600
rect -800 16700 -700 18500
rect 600 18445 4310 18500
rect 600 16700 787 18445
rect -800 16685 -477 16700
rect -411 16685 -161 16700
rect -95 16685 155 16700
rect 221 16685 471 16700
rect 537 16685 787 16700
rect 853 16685 1103 18445
rect 1169 16685 1419 18445
rect 1485 16685 1735 18445
rect 1801 16685 2051 18445
rect 2117 16685 2367 18445
rect 2433 16685 2683 18445
rect 2749 16685 2999 18445
rect 3065 16685 3315 18445
rect 3381 16685 3631 18445
rect 3697 16685 3947 18445
rect 4013 16685 4310 18445
rect -800 16600 4310 16685
rect 5500 18500 10610 18600
rect 5500 16700 5600 18500
rect 6800 18445 10610 18500
rect 5500 16685 5823 16700
rect 5889 16685 6139 16700
rect 6205 16685 6455 16700
rect 6521 16685 6771 16700
rect 6837 16685 7087 18445
rect 7153 16685 7403 18445
rect 7469 16685 7719 18445
rect 7785 16685 8035 18445
rect 8101 16685 8351 18445
rect 8417 16685 8667 18445
rect 8733 16685 8983 18445
rect 9049 16685 9299 18445
rect 9365 16685 9615 18445
rect 9681 16685 9931 18445
rect 9997 16685 10247 18445
rect 10313 16685 10610 18445
rect 5500 16600 10610 16685
rect -13400 15500 -8290 15600
rect -13400 13700 -13300 15500
rect -12000 15445 -8290 15500
rect -12000 13700 -11971 15445
rect -13400 13685 -13235 13700
rect -13169 13685 -12919 13700
rect -12853 13685 -12603 13700
rect -12537 13685 -12287 13700
rect -12221 13685 -11971 13700
rect -11905 13685 -11655 15445
rect -11589 13685 -11339 15445
rect -11273 13685 -11023 15445
rect -10957 13685 -10707 15445
rect -10641 13685 -10391 15445
rect -10325 13685 -10075 15445
rect -10009 13685 -9759 15445
rect -9693 13685 -9443 15445
rect -9377 13685 -9127 15445
rect -9061 13685 -8811 15445
rect -8745 13685 -8495 15445
rect -8429 13685 -8290 15445
rect -13400 13600 -8290 13685
rect -7070 15500 -1800 15600
rect -7070 15445 -3200 15500
rect -7070 13685 -6935 15445
rect -6869 13685 -6619 15445
rect -6553 13685 -6303 15445
rect -6237 13685 -5987 15445
rect -5921 13685 -5671 15445
rect -5605 13685 -5355 15445
rect -5289 13685 -5039 15445
rect -4973 13685 -4723 15445
rect -4657 13685 -4407 15445
rect -4341 13685 -4091 15445
rect -4025 13685 -3775 15445
rect -3709 13685 -3459 15445
rect -3393 13700 -3200 15445
rect -1900 13700 -1800 15500
rect -3393 13685 -3143 13700
rect -3077 13685 -2827 13700
rect -2761 13685 -2511 13700
rect -2445 13685 -2195 13700
rect -2129 13685 -1800 13700
rect -7070 13600 -1800 13685
rect -800 15500 4310 15600
rect -800 13700 -700 15500
rect 600 15445 4310 15500
rect 600 13700 629 15445
rect -800 13685 -635 13700
rect -569 13685 -319 13700
rect -253 13685 -3 13700
rect 63 13685 313 13700
rect 379 13685 629 13700
rect 695 13685 945 15445
rect 1011 13685 1261 15445
rect 1327 13685 1577 15445
rect 1643 13685 1893 15445
rect 1959 13685 2209 15445
rect 2275 13685 2525 15445
rect 2591 13685 2841 15445
rect 2907 13685 3157 15445
rect 3223 13685 3473 15445
rect 3539 13685 3789 15445
rect 3855 13685 4105 15445
rect 4171 13685 4310 15445
rect -800 13600 4310 13685
rect 5530 15500 10800 15600
rect 5530 15445 9400 15500
rect 5530 13685 5665 15445
rect 5731 13685 5981 15445
rect 6047 13685 6297 15445
rect 6363 13685 6613 15445
rect 6679 13685 6929 15445
rect 6995 13685 7245 15445
rect 7311 13685 7561 15445
rect 7627 13685 7877 15445
rect 7943 13685 8193 15445
rect 8259 13685 8509 15445
rect 8575 13685 8825 15445
rect 8891 13685 9141 15445
rect 9207 13700 9400 15445
rect 10700 13700 10800 15500
rect 9207 13685 9457 13700
rect 9523 13685 9773 13700
rect 9839 13685 10089 13700
rect 10155 13685 10405 13700
rect 10471 13685 10800 13700
rect 5530 13600 10800 13685
rect -11700 13200 -9800 13300
rect -11700 13100 -11500 13200
rect -13400 13010 -11500 13100
rect -10000 13100 -9800 13200
rect 900 13200 2800 13300
rect 900 13100 1100 13200
rect -10000 13010 -7400 13100
rect -13400 12940 -13160 13010
rect -8510 12980 -7400 13010
rect -8510 12940 -7780 12980
rect -13400 12900 -11500 12940
rect -10000 12900 -7780 12940
rect -13400 12820 -7780 12900
rect -7420 12820 -7400 12980
rect -13400 12800 -7400 12820
rect -7200 13010 -1100 13100
rect -7200 12940 -6860 13010
rect -2210 12980 -1100 13010
rect -2210 12940 -1480 12980
rect -7200 12820 -1480 12940
rect -1120 12820 -1100 12980
rect -7200 12800 -1100 12820
rect -900 13010 1100 13100
rect 2600 13100 2800 13200
rect 2600 13010 5200 13100
rect -900 12940 -560 13010
rect 4090 12980 5200 13010
rect 4090 12940 4820 12980
rect -900 12900 1100 12940
rect 2600 12900 4820 12940
rect -900 12820 4820 12900
rect 5180 12820 5200 12980
rect -900 12800 5200 12820
rect 5400 13010 10600 13100
rect 5400 12940 5740 13010
rect 10390 12940 10600 13010
rect 5400 12800 10600 12940
rect -7200 12600 -6900 12800
rect -5400 12700 -2800 12800
rect -900 12700 -700 12800
rect 5400 12700 5700 12800
rect 7200 12700 9800 12800
rect -8300 12400 -6900 12600
rect -2000 12500 -700 12700
rect 4300 12500 5700 12700
rect -11700 12300 -9800 12400
rect -8300 12300 -8000 12400
rect -5400 12300 -2800 12400
rect -2000 12300 -1700 12500
rect 900 12300 2800 12400
rect 4300 12300 4600 12500
rect 7200 12300 9800 12400
rect -13400 12180 -11500 12300
rect -10000 12180 -8000 12300
rect -13400 12110 -13160 12180
rect -8500 12110 -8000 12180
rect -13400 12000 -11500 12110
rect -10000 12000 -8000 12110
rect -7800 12280 -1700 12300
rect -7800 12120 -7780 12280
rect -7420 12180 -1700 12280
rect -7420 12120 -6860 12180
rect -7800 12110 -6860 12120
rect -2200 12110 -1700 12180
rect -7800 12000 -1700 12110
rect -1500 12280 1100 12300
rect -1500 12120 -1480 12280
rect -1120 12180 1100 12280
rect 2600 12180 4600 12300
rect -1120 12120 -560 12180
rect -1500 12110 -560 12120
rect 4100 12110 4600 12180
rect -1500 12000 1100 12110
rect 2600 12000 4600 12110
rect 4800 12280 10600 12300
rect 4800 12120 4820 12280
rect 5180 12180 10600 12280
rect 5180 12120 5740 12180
rect 4800 12110 5740 12120
rect 10400 12110 10600 12180
rect 4800 12000 10600 12110
rect -11700 11900 -9800 12000
rect 900 11900 2800 12000
rect -13370 11500 -8290 11600
rect -13370 11445 -11400 11500
rect -10100 11445 -8290 11500
rect -13370 9685 -13077 11445
rect -13011 9685 -12761 11445
rect -12695 9685 -12445 11445
rect -12379 9685 -12129 11445
rect -12063 9685 -11813 11445
rect -11747 9685 -11497 11445
rect -11431 9700 -11400 11445
rect -10100 9700 -9917 11445
rect -11431 9685 -11181 9700
rect -11115 9685 -10865 9700
rect -10799 9685 -10549 9700
rect -10483 9685 -10233 9700
rect -10167 9685 -9917 9700
rect -9851 9685 -9601 11445
rect -9535 9685 -9285 11445
rect -9219 9685 -8969 11445
rect -8903 9685 -8653 11445
rect -8587 9685 -8290 11445
rect -13370 9600 -8290 9685
rect -7100 11500 -1990 11600
rect -7100 9700 -7000 11500
rect -5700 11445 -1990 11500
rect -5700 9700 -5513 11445
rect -7100 9685 -6777 9700
rect -6711 9685 -6461 9700
rect -6395 9685 -6145 9700
rect -6079 9685 -5829 9700
rect -5763 9685 -5513 9700
rect -5447 9685 -5197 11445
rect -5131 9685 -4881 11445
rect -4815 9685 -4565 11445
rect -4499 9685 -4249 11445
rect -4183 9685 -3933 11445
rect -3867 9685 -3617 11445
rect -3551 9685 -3301 11445
rect -3235 9685 -2985 11445
rect -2919 9685 -2669 11445
rect -2603 9685 -2353 11445
rect -2287 9685 -1990 11445
rect -7100 9600 -1990 9685
rect -770 11500 4310 11600
rect -770 11445 1200 11500
rect 2500 11445 4310 11500
rect -770 9685 -477 11445
rect -411 9685 -161 11445
rect -95 9685 155 11445
rect 221 9685 471 11445
rect 537 9685 787 11445
rect 853 9685 1103 11445
rect 1169 9700 1200 11445
rect 2500 9700 2683 11445
rect 1169 9685 1419 9700
rect 1485 9685 1735 9700
rect 1801 9685 2051 9700
rect 2117 9685 2367 9700
rect 2433 9685 2683 9700
rect 2749 9685 2999 11445
rect 3065 9685 3315 11445
rect 3381 9685 3631 11445
rect 3697 9685 3947 11445
rect 4013 9685 4310 11445
rect -770 9600 4310 9685
rect 5500 11500 10610 11600
rect 5500 9700 5600 11500
rect 6900 11445 10610 11500
rect 6900 9700 7087 11445
rect 5500 9685 5823 9700
rect 5889 9685 6139 9700
rect 6205 9685 6455 9700
rect 6521 9685 6771 9700
rect 6837 9685 7087 9700
rect 7153 9685 7403 11445
rect 7469 9685 7719 11445
rect 7785 9685 8035 11445
rect 8101 9685 8351 11445
rect 8417 9685 8667 11445
rect 8733 9685 8983 11445
rect 9049 9685 9299 11445
rect 9365 9685 9615 11445
rect 9681 9685 9931 11445
rect 9997 9685 10247 11445
rect 10313 9685 10610 11445
rect 5500 9600 10610 9685
rect -13370 8500 -8100 8600
rect -13370 8445 -9500 8500
rect -13370 6685 -13235 8445
rect -13169 6685 -12919 8445
rect -12853 6685 -12603 8445
rect -12537 6685 -12287 8445
rect -12221 6685 -11971 8445
rect -11905 6685 -11655 8445
rect -11589 6685 -11339 8445
rect -11273 6685 -11023 8445
rect -10957 6685 -10707 8445
rect -10641 6685 -10391 8445
rect -10325 6685 -10075 8445
rect -10009 6685 -9759 8445
rect -9693 6700 -9500 8445
rect -8200 6700 -8100 8500
rect -9693 6685 -9443 6700
rect -9377 6685 -9127 6700
rect -9061 6685 -8811 6700
rect -8745 6685 -8495 6700
rect -8429 6685 -8100 6700
rect -13370 6600 -8100 6685
rect -7070 8500 -1990 8600
rect -7070 8445 -5100 8500
rect -3800 8445 -1990 8500
rect -7070 6685 -6935 8445
rect -6869 6685 -6619 8445
rect -6553 6685 -6303 8445
rect -6237 6685 -5987 8445
rect -5921 6685 -5671 8445
rect -5605 6685 -5355 8445
rect -5289 6700 -5100 8445
rect -3800 6700 -3775 8445
rect -5289 6685 -5039 6700
rect -4973 6685 -4723 6700
rect -4657 6685 -4407 6700
rect -4341 6685 -4091 6700
rect -4025 6685 -3775 6700
rect -3709 6685 -3459 8445
rect -3393 6685 -3143 8445
rect -3077 6685 -2827 8445
rect -2761 6685 -2511 8445
rect -2445 6685 -2195 8445
rect -2129 6685 -1990 8445
rect -7070 6600 -1990 6685
rect -770 8500 4500 8600
rect -770 8445 3100 8500
rect -770 6685 -635 8445
rect -569 6685 -319 8445
rect -253 6685 -3 8445
rect 63 6685 313 8445
rect 379 6685 629 8445
rect 695 6685 945 8445
rect 1011 6685 1261 8445
rect 1327 6685 1577 8445
rect 1643 6685 1893 8445
rect 1959 6685 2209 8445
rect 2275 6685 2525 8445
rect 2591 6685 2841 8445
rect 2907 6700 3100 8445
rect 4400 6700 4500 8500
rect 2907 6685 3157 6700
rect 3223 6685 3473 6700
rect 3539 6685 3789 6700
rect 3855 6685 4105 6700
rect 4171 6685 4500 6700
rect -770 6600 4500 6685
rect 5500 8500 10800 8600
rect 5500 8445 7500 8500
rect 8800 8445 10800 8500
rect 5500 6685 5665 8445
rect 5731 6685 5981 8445
rect 6047 6685 6297 8445
rect 6363 6685 6613 8445
rect 6679 6685 6929 8445
rect 6995 6685 7245 8445
rect 7311 6700 7500 8445
rect 8800 6700 8825 8445
rect 7311 6685 7561 6700
rect 7627 6685 7877 6700
rect 7943 6685 8193 6700
rect 8259 6685 8509 6700
rect 8575 6685 8825 6700
rect 8891 6685 9141 8445
rect 9207 6685 9457 8445
rect 9523 6685 9773 8445
rect 9839 6685 10089 8445
rect 10155 6685 10405 8445
rect 10471 6685 10800 8445
rect 5500 6600 10800 6685
rect -13300 6010 -8300 6030
rect -13300 5940 -13160 6010
rect -8510 5940 -8300 6010
rect -13300 5830 -8300 5940
rect -7000 6010 -2000 6030
rect -7000 5940 -6860 6010
rect -2210 5940 -2000 6010
rect -7000 5830 -2000 5940
rect -700 6010 4300 6030
rect -700 5940 -560 6010
rect 4090 5940 4300 6010
rect -700 5830 4300 5940
rect 5600 6010 10600 6030
rect 5600 5940 5740 6010
rect 10390 5940 10600 6010
rect 5600 5830 10600 5940
<< via3 >>
rect -13300 49045 -12000 49100
rect -13300 47300 -13077 49045
rect -13077 47300 -13011 49045
rect -13011 47300 -12761 49045
rect -12761 47300 -12695 49045
rect -12695 47300 -12445 49045
rect -12445 47300 -12379 49045
rect -12379 47300 -12129 49045
rect -12129 47300 -12063 49045
rect -12063 47300 -12000 49045
rect -7000 49045 -5800 49100
rect -7000 47300 -6777 49045
rect -6777 47300 -6711 49045
rect -6711 47300 -6461 49045
rect -6461 47300 -6395 49045
rect -6395 47300 -6145 49045
rect -6145 47300 -6079 49045
rect -6079 47300 -5829 49045
rect -5829 47300 -5800 49045
rect -700 49045 600 49100
rect -700 47300 -477 49045
rect -477 47300 -411 49045
rect -411 47300 -161 49045
rect -161 47300 -95 49045
rect -95 47300 155 49045
rect 155 47300 221 49045
rect 221 47300 471 49045
rect 471 47300 537 49045
rect 537 47300 600 49045
rect 5600 49045 6800 49100
rect 5600 47300 5823 49045
rect 5823 47300 5889 49045
rect 5889 47300 6139 49045
rect 6139 47300 6205 49045
rect 6205 47300 6455 49045
rect 6455 47300 6521 49045
rect 6521 47300 6771 49045
rect 6771 47300 6800 49045
rect -13300 46045 -12000 46100
rect -13300 44300 -13235 46045
rect -13235 44300 -13169 46045
rect -13169 44300 -12919 46045
rect -12919 44300 -12853 46045
rect -12853 44300 -12603 46045
rect -12603 44300 -12537 46045
rect -12537 44300 -12287 46045
rect -12287 44300 -12221 46045
rect -12221 44300 -12000 46045
rect -3200 46045 -1900 46100
rect -3200 44300 -3143 46045
rect -3143 44300 -3077 46045
rect -3077 44300 -2827 46045
rect -2827 44300 -2761 46045
rect -2761 44300 -2511 46045
rect -2511 44300 -2445 46045
rect -2445 44300 -2195 46045
rect -2195 44300 -2129 46045
rect -2129 44300 -1900 46045
rect -700 46045 600 46100
rect -700 44300 -635 46045
rect -635 44300 -569 46045
rect -569 44300 -319 46045
rect -319 44300 -253 46045
rect -253 44300 -3 46045
rect -3 44300 63 46045
rect 63 44300 313 46045
rect 313 44300 379 46045
rect 379 44300 600 46045
rect 9400 46045 10700 46100
rect 9400 44300 9457 46045
rect 9457 44300 9523 46045
rect 9523 44300 9773 46045
rect 9773 44300 9839 46045
rect 9839 44300 10089 46045
rect 10089 44300 10155 46045
rect 10155 44300 10405 46045
rect 10405 44300 10471 46045
rect 10471 44300 10700 46045
rect -11500 43610 -10000 43800
rect -11500 43540 -10000 43610
rect -11500 43500 -10000 43540
rect -7780 43420 -7420 43580
rect -1480 43420 -1120 43580
rect 1100 43610 2600 43800
rect 1100 43540 2600 43610
rect 1100 43500 2600 43540
rect 4820 43420 5180 43580
rect -11500 42780 -10000 42900
rect -11500 42710 -10000 42780
rect -11500 42600 -10000 42710
rect -7780 42720 -7420 42880
rect -1480 42720 -1120 42880
rect 1100 42780 2600 42900
rect 1100 42710 2600 42780
rect 1100 42600 2600 42710
rect 4820 42720 5180 42880
rect -11400 42045 -10100 42100
rect -11400 40300 -11181 42045
rect -11181 40300 -11115 42045
rect -11115 40300 -10865 42045
rect -10865 40300 -10799 42045
rect -10799 40300 -10549 42045
rect -10549 40300 -10483 42045
rect -10483 40300 -10233 42045
rect -10233 40300 -10167 42045
rect -10167 40300 -10100 42045
rect -7000 42045 -5700 42100
rect -7000 40300 -6777 42045
rect -6777 40300 -6711 42045
rect -6711 40300 -6461 42045
rect -6461 40300 -6395 42045
rect -6395 40300 -6145 42045
rect -6145 40300 -6079 42045
rect -6079 40300 -5829 42045
rect -5829 40300 -5763 42045
rect -5763 40300 -5700 42045
rect 1200 42045 2500 42100
rect 1200 40300 1419 42045
rect 1419 40300 1485 42045
rect 1485 40300 1735 42045
rect 1735 40300 1801 42045
rect 1801 40300 2051 42045
rect 2051 40300 2117 42045
rect 2117 40300 2367 42045
rect 2367 40300 2433 42045
rect 2433 40300 2500 42045
rect 5600 42045 6900 42100
rect 5600 40300 5823 42045
rect 5823 40300 5889 42045
rect 5889 40300 6139 42045
rect 6139 40300 6205 42045
rect 6205 40300 6455 42045
rect 6455 40300 6521 42045
rect 6521 40300 6771 42045
rect 6771 40300 6837 42045
rect 6837 40300 6900 42045
rect -9500 39045 -8200 39100
rect -9500 37300 -9443 39045
rect -9443 37300 -9377 39045
rect -9377 37300 -9127 39045
rect -9127 37300 -9061 39045
rect -9061 37300 -8811 39045
rect -8811 37300 -8745 39045
rect -8745 37300 -8495 39045
rect -8495 37300 -8429 39045
rect -8429 37300 -8200 39045
rect -5100 39045 -3800 39100
rect -5100 37300 -5039 39045
rect -5039 37300 -4973 39045
rect -4973 37300 -4723 39045
rect -4723 37300 -4657 39045
rect -4657 37300 -4407 39045
rect -4407 37300 -4341 39045
rect -4341 37300 -4091 39045
rect -4091 37300 -4025 39045
rect -4025 37300 -3800 39045
rect 3100 39045 4400 39100
rect 3100 37300 3157 39045
rect 3157 37300 3223 39045
rect 3223 37300 3473 39045
rect 3473 37300 3539 39045
rect 3539 37300 3789 39045
rect 3789 37300 3855 39045
rect 3855 37300 4105 39045
rect 4105 37300 4171 39045
rect 4171 37300 4400 39045
rect 7500 39045 8800 39100
rect 7500 37300 7561 39045
rect 7561 37300 7627 39045
rect 7627 37300 7877 39045
rect 7877 37300 7943 39045
rect 7943 37300 8193 39045
rect 8193 37300 8259 39045
rect 8259 37300 8509 39045
rect 8509 37300 8575 39045
rect 8575 37300 8800 39045
rect -13300 33745 -12000 33800
rect -13300 32000 -13077 33745
rect -13077 32000 -13011 33745
rect -13011 32000 -12761 33745
rect -12761 32000 -12695 33745
rect -12695 32000 -12445 33745
rect -12445 32000 -12379 33745
rect -12379 32000 -12129 33745
rect -12129 32000 -12063 33745
rect -12063 32000 -12000 33745
rect -7000 33745 -5800 33800
rect -7000 32000 -6777 33745
rect -6777 32000 -6711 33745
rect -6711 32000 -6461 33745
rect -6461 32000 -6395 33745
rect -6395 32000 -6145 33745
rect -6145 32000 -6079 33745
rect -6079 32000 -5829 33745
rect -5829 32000 -5800 33745
rect -700 33745 600 33800
rect -700 32000 -477 33745
rect -477 32000 -411 33745
rect -411 32000 -161 33745
rect -161 32000 -95 33745
rect -95 32000 155 33745
rect 155 32000 221 33745
rect 221 32000 471 33745
rect 471 32000 537 33745
rect 537 32000 600 33745
rect 5600 33745 6800 33800
rect 5600 32000 5823 33745
rect 5823 32000 5889 33745
rect 5889 32000 6139 33745
rect 6139 32000 6205 33745
rect 6205 32000 6455 33745
rect 6455 32000 6521 33745
rect 6521 32000 6771 33745
rect 6771 32000 6800 33745
rect -13300 30745 -12000 30800
rect -13300 29000 -13235 30745
rect -13235 29000 -13169 30745
rect -13169 29000 -12919 30745
rect -12919 29000 -12853 30745
rect -12853 29000 -12603 30745
rect -12603 29000 -12537 30745
rect -12537 29000 -12287 30745
rect -12287 29000 -12221 30745
rect -12221 29000 -12000 30745
rect -3200 30745 -1900 30800
rect -3200 29000 -3143 30745
rect -3143 29000 -3077 30745
rect -3077 29000 -2827 30745
rect -2827 29000 -2761 30745
rect -2761 29000 -2511 30745
rect -2511 29000 -2445 30745
rect -2445 29000 -2195 30745
rect -2195 29000 -2129 30745
rect -2129 29000 -1900 30745
rect -700 30745 600 30800
rect -700 29000 -635 30745
rect -635 29000 -569 30745
rect -569 29000 -319 30745
rect -319 29000 -253 30745
rect -253 29000 -3 30745
rect -3 29000 63 30745
rect 63 29000 313 30745
rect 313 29000 379 30745
rect 379 29000 600 30745
rect 9400 30745 10700 30800
rect 9400 29000 9457 30745
rect 9457 29000 9523 30745
rect 9523 29000 9773 30745
rect 9773 29000 9839 30745
rect 9839 29000 10089 30745
rect 10089 29000 10155 30745
rect 10155 29000 10405 30745
rect 10405 29000 10471 30745
rect 10471 29000 10700 30745
rect -11500 28310 -10000 28500
rect -11500 28240 -10000 28310
rect -11500 28200 -10000 28240
rect -7780 28120 -7420 28280
rect -1480 28120 -1120 28280
rect 1100 28310 2600 28500
rect 1100 28240 2600 28310
rect 1100 28200 2600 28240
rect 4820 28120 5180 28280
rect -11500 27480 -10000 27600
rect -11500 27410 -10000 27480
rect -11500 27300 -10000 27410
rect -7780 27420 -7420 27580
rect -1480 27420 -1120 27580
rect 1100 27480 2600 27600
rect 1100 27410 2600 27480
rect 1100 27300 2600 27410
rect 4820 27420 5180 27580
rect -11400 26745 -10100 26800
rect -11400 25000 -11181 26745
rect -11181 25000 -11115 26745
rect -11115 25000 -10865 26745
rect -10865 25000 -10799 26745
rect -10799 25000 -10549 26745
rect -10549 25000 -10483 26745
rect -10483 25000 -10233 26745
rect -10233 25000 -10167 26745
rect -10167 25000 -10100 26745
rect -7000 26745 -5700 26800
rect -7000 25000 -6777 26745
rect -6777 25000 -6711 26745
rect -6711 25000 -6461 26745
rect -6461 25000 -6395 26745
rect -6395 25000 -6145 26745
rect -6145 25000 -6079 26745
rect -6079 25000 -5829 26745
rect -5829 25000 -5763 26745
rect -5763 25000 -5700 26745
rect 1200 26745 2500 26800
rect 1200 25000 1419 26745
rect 1419 25000 1485 26745
rect 1485 25000 1735 26745
rect 1735 25000 1801 26745
rect 1801 25000 2051 26745
rect 2051 25000 2117 26745
rect 2117 25000 2367 26745
rect 2367 25000 2433 26745
rect 2433 25000 2500 26745
rect 5600 26745 6900 26800
rect 5600 25000 5823 26745
rect 5823 25000 5889 26745
rect 5889 25000 6139 26745
rect 6139 25000 6205 26745
rect 6205 25000 6455 26745
rect 6455 25000 6521 26745
rect 6521 25000 6771 26745
rect 6771 25000 6837 26745
rect 6837 25000 6900 26745
rect -9500 23745 -8200 23800
rect -9500 22000 -9443 23745
rect -9443 22000 -9377 23745
rect -9377 22000 -9127 23745
rect -9127 22000 -9061 23745
rect -9061 22000 -8811 23745
rect -8811 22000 -8745 23745
rect -8745 22000 -8495 23745
rect -8495 22000 -8429 23745
rect -8429 22000 -8200 23745
rect -5100 23745 -3800 23800
rect -5100 22000 -5039 23745
rect -5039 22000 -4973 23745
rect -4973 22000 -4723 23745
rect -4723 22000 -4657 23745
rect -4657 22000 -4407 23745
rect -4407 22000 -4341 23745
rect -4341 22000 -4091 23745
rect -4091 22000 -4025 23745
rect -4025 22000 -3800 23745
rect 3100 23745 4400 23800
rect 3100 22000 3157 23745
rect 3157 22000 3223 23745
rect 3223 22000 3473 23745
rect 3473 22000 3539 23745
rect 3539 22000 3789 23745
rect 3789 22000 3855 23745
rect 3855 22000 4105 23745
rect 4105 22000 4171 23745
rect 4171 22000 4400 23745
rect 7500 23745 8800 23800
rect 7500 22000 7561 23745
rect 7561 22000 7627 23745
rect 7627 22000 7877 23745
rect 7877 22000 7943 23745
rect 7943 22000 8193 23745
rect 8193 22000 8259 23745
rect 8259 22000 8509 23745
rect 8509 22000 8575 23745
rect 8575 22000 8800 23745
rect -13300 18445 -12000 18500
rect -13300 16700 -13077 18445
rect -13077 16700 -13011 18445
rect -13011 16700 -12761 18445
rect -12761 16700 -12695 18445
rect -12695 16700 -12445 18445
rect -12445 16700 -12379 18445
rect -12379 16700 -12129 18445
rect -12129 16700 -12063 18445
rect -12063 16700 -12000 18445
rect -7000 18445 -5800 18500
rect -7000 16700 -6777 18445
rect -6777 16700 -6711 18445
rect -6711 16700 -6461 18445
rect -6461 16700 -6395 18445
rect -6395 16700 -6145 18445
rect -6145 16700 -6079 18445
rect -6079 16700 -5829 18445
rect -5829 16700 -5800 18445
rect -700 18445 600 18500
rect -700 16700 -477 18445
rect -477 16700 -411 18445
rect -411 16700 -161 18445
rect -161 16700 -95 18445
rect -95 16700 155 18445
rect 155 16700 221 18445
rect 221 16700 471 18445
rect 471 16700 537 18445
rect 537 16700 600 18445
rect 5600 18445 6800 18500
rect 5600 16700 5823 18445
rect 5823 16700 5889 18445
rect 5889 16700 6139 18445
rect 6139 16700 6205 18445
rect 6205 16700 6455 18445
rect 6455 16700 6521 18445
rect 6521 16700 6771 18445
rect 6771 16700 6800 18445
rect -13300 15445 -12000 15500
rect -13300 13700 -13235 15445
rect -13235 13700 -13169 15445
rect -13169 13700 -12919 15445
rect -12919 13700 -12853 15445
rect -12853 13700 -12603 15445
rect -12603 13700 -12537 15445
rect -12537 13700 -12287 15445
rect -12287 13700 -12221 15445
rect -12221 13700 -12000 15445
rect -3200 15445 -1900 15500
rect -3200 13700 -3143 15445
rect -3143 13700 -3077 15445
rect -3077 13700 -2827 15445
rect -2827 13700 -2761 15445
rect -2761 13700 -2511 15445
rect -2511 13700 -2445 15445
rect -2445 13700 -2195 15445
rect -2195 13700 -2129 15445
rect -2129 13700 -1900 15445
rect -700 15445 600 15500
rect -700 13700 -635 15445
rect -635 13700 -569 15445
rect -569 13700 -319 15445
rect -319 13700 -253 15445
rect -253 13700 -3 15445
rect -3 13700 63 15445
rect 63 13700 313 15445
rect 313 13700 379 15445
rect 379 13700 600 15445
rect 9400 15445 10700 15500
rect 9400 13700 9457 15445
rect 9457 13700 9523 15445
rect 9523 13700 9773 15445
rect 9773 13700 9839 15445
rect 9839 13700 10089 15445
rect 10089 13700 10155 15445
rect 10155 13700 10405 15445
rect 10405 13700 10471 15445
rect 10471 13700 10700 15445
rect -11500 13010 -10000 13200
rect -11500 12940 -10000 13010
rect -11500 12900 -10000 12940
rect -7780 12820 -7420 12980
rect -1480 12820 -1120 12980
rect 1100 13010 2600 13200
rect 1100 12940 2600 13010
rect 1100 12900 2600 12940
rect 4820 12820 5180 12980
rect -11500 12180 -10000 12300
rect -11500 12110 -10000 12180
rect -11500 12000 -10000 12110
rect -7780 12120 -7420 12280
rect -1480 12120 -1120 12280
rect 1100 12180 2600 12300
rect 1100 12110 2600 12180
rect 1100 12000 2600 12110
rect 4820 12120 5180 12280
rect -11400 11445 -10100 11500
rect -11400 9700 -11181 11445
rect -11181 9700 -11115 11445
rect -11115 9700 -10865 11445
rect -10865 9700 -10799 11445
rect -10799 9700 -10549 11445
rect -10549 9700 -10483 11445
rect -10483 9700 -10233 11445
rect -10233 9700 -10167 11445
rect -10167 9700 -10100 11445
rect -7000 11445 -5700 11500
rect -7000 9700 -6777 11445
rect -6777 9700 -6711 11445
rect -6711 9700 -6461 11445
rect -6461 9700 -6395 11445
rect -6395 9700 -6145 11445
rect -6145 9700 -6079 11445
rect -6079 9700 -5829 11445
rect -5829 9700 -5763 11445
rect -5763 9700 -5700 11445
rect 1200 11445 2500 11500
rect 1200 9700 1419 11445
rect 1419 9700 1485 11445
rect 1485 9700 1735 11445
rect 1735 9700 1801 11445
rect 1801 9700 2051 11445
rect 2051 9700 2117 11445
rect 2117 9700 2367 11445
rect 2367 9700 2433 11445
rect 2433 9700 2500 11445
rect 5600 11445 6900 11500
rect 5600 9700 5823 11445
rect 5823 9700 5889 11445
rect 5889 9700 6139 11445
rect 6139 9700 6205 11445
rect 6205 9700 6455 11445
rect 6455 9700 6521 11445
rect 6521 9700 6771 11445
rect 6771 9700 6837 11445
rect 6837 9700 6900 11445
rect -9500 8445 -8200 8500
rect -9500 6700 -9443 8445
rect -9443 6700 -9377 8445
rect -9377 6700 -9127 8445
rect -9127 6700 -9061 8445
rect -9061 6700 -8811 8445
rect -8811 6700 -8745 8445
rect -8745 6700 -8495 8445
rect -8495 6700 -8429 8445
rect -8429 6700 -8200 8445
rect -5100 8445 -3800 8500
rect -5100 6700 -5039 8445
rect -5039 6700 -4973 8445
rect -4973 6700 -4723 8445
rect -4723 6700 -4657 8445
rect -4657 6700 -4407 8445
rect -4407 6700 -4341 8445
rect -4341 6700 -4091 8445
rect -4091 6700 -4025 8445
rect -4025 6700 -3800 8445
rect 3100 8445 4400 8500
rect 3100 6700 3157 8445
rect 3157 6700 3223 8445
rect 3223 6700 3473 8445
rect 3473 6700 3539 8445
rect 3539 6700 3789 8445
rect 3789 6700 3855 8445
rect 3855 6700 4105 8445
rect 4105 6700 4171 8445
rect 4171 6700 4400 8445
rect 7500 8445 8800 8500
rect 7500 6700 7561 8445
rect 7561 6700 7627 8445
rect 7627 6700 7877 8445
rect 7877 6700 7943 8445
rect 7943 6700 8193 8445
rect 8193 6700 8259 8445
rect 8259 6700 8509 8445
rect 8509 6700 8575 8445
rect 8575 6700 8800 8445
<< metal4 >>
rect -13400 51700 -11900 51800
rect -13400 50500 -13300 51700
rect -12000 50500 -11900 51700
rect -13400 49100 -11900 50500
rect -5200 51700 -3700 51800
rect -5200 50500 -5100 51700
rect -3800 50500 -3700 51700
rect -13400 47300 -13300 49100
rect -12000 47300 -11900 49100
rect -13400 47200 -11900 47300
rect -9600 49900 -8100 50000
rect -9600 48700 -9500 49900
rect -8200 48700 -8100 49900
rect -13400 46100 -11900 46200
rect -13400 44300 -13300 46100
rect -12000 44300 -11900 46100
rect -13400 36800 -11900 44300
rect -11600 43800 -9900 43900
rect -11600 43500 -11500 43800
rect -10000 43500 -9900 43800
rect -11600 43400 -9900 43500
rect -11600 42900 -9900 43000
rect -11600 42600 -11500 42900
rect -10000 42600 -9900 42900
rect -11600 42500 -9900 42600
rect -13400 35600 -13300 36800
rect -12000 35600 -11900 36800
rect -13400 33800 -11900 35600
rect -13400 32000 -13300 33800
rect -12000 32000 -11900 33800
rect -11500 42100 -10000 42200
rect -11500 40300 -11400 42100
rect -10100 40300 -10000 42100
rect -11500 34600 -10000 40300
rect -9600 39100 -8100 48700
rect -7100 49900 -5600 50000
rect -7100 47300 -7000 49900
rect -5700 48700 -5600 49900
rect -5800 47300 -5600 48700
rect -7100 47200 -5600 47300
rect -7800 43580 -7400 43600
rect -7800 43420 -7780 43580
rect -7420 43420 -7400 43580
rect -7800 42880 -7400 43420
rect -7800 42720 -7780 42880
rect -7420 42720 -7400 42880
rect -7800 42700 -7400 42720
rect -9600 37300 -9500 39100
rect -8200 37300 -8100 39100
rect -9600 37200 -8100 37300
rect -7100 42100 -5600 42200
rect -7100 40300 -7000 42100
rect -5700 40300 -5600 42100
rect -7100 36800 -5600 40300
rect -5200 39100 -3700 50500
rect -800 51700 700 51800
rect -800 50500 -700 51700
rect 600 50500 700 51700
rect -800 49100 700 50500
rect 7400 51700 8900 51800
rect 7400 50500 7500 51700
rect 8800 50500 8900 51700
rect -800 47300 -700 49100
rect 600 47300 700 49100
rect -800 47200 700 47300
rect 3000 49900 4500 50000
rect 3000 48700 3100 49900
rect 4400 48700 4500 49900
rect -5200 37300 -5100 39100
rect -3800 37300 -3700 39100
rect -5200 37200 -3700 37300
rect -3300 46100 -1800 46200
rect -3300 44300 -3200 46100
rect -1900 44300 -1800 46100
rect -7100 35600 -7000 36800
rect -5700 35600 -5600 36800
rect -7100 35500 -5600 35600
rect -5200 36800 -3700 36900
rect -5200 35600 -5100 36800
rect -3800 35600 -3700 36800
rect -11500 33400 -11400 34600
rect -10100 33400 -10000 34600
rect -11500 33300 -10000 33400
rect -9600 34600 -8100 34700
rect -9600 33400 -9500 34600
rect -8200 33400 -8100 34600
rect -13400 31900 -11900 32000
rect -13400 30800 -11900 30900
rect -13400 29000 -13300 30800
rect -12000 29000 -11900 30800
rect -13400 21500 -11900 29000
rect -11600 28500 -9900 28600
rect -11600 28200 -11500 28500
rect -10000 28200 -9900 28500
rect -11600 28100 -9900 28200
rect -11600 27600 -9900 27700
rect -11600 27300 -11500 27600
rect -10000 27300 -9900 27600
rect -11600 27200 -9900 27300
rect -13400 20300 -13300 21500
rect -12000 20300 -11900 21500
rect -13400 18500 -11900 20300
rect -13400 16700 -13300 18500
rect -12000 16700 -11900 18500
rect -11500 26800 -10000 26900
rect -11500 25000 -11400 26800
rect -10100 25000 -10000 26800
rect -11500 19300 -10000 25000
rect -9600 23800 -8100 33400
rect -7100 34600 -5600 34700
rect -7100 32000 -7000 34600
rect -5700 33400 -5600 34600
rect -5800 32000 -5600 33400
rect -7100 31900 -5600 32000
rect -7800 28280 -7400 28300
rect -7800 28120 -7780 28280
rect -7420 28120 -7400 28280
rect -7800 27580 -7400 28120
rect -7800 27420 -7780 27580
rect -7420 27420 -7400 27580
rect -7800 27400 -7400 27420
rect -9600 22000 -9500 23800
rect -8200 22000 -8100 23800
rect -9600 21900 -8100 22000
rect -7100 26800 -5600 26900
rect -7100 25000 -7000 26800
rect -5700 25000 -5600 26800
rect -7100 21500 -5600 25000
rect -5200 23800 -3700 35600
rect -3300 34600 -1800 44300
rect -800 46100 700 46200
rect -800 44300 -700 46100
rect 600 44300 700 46100
rect -1500 43580 -1100 43600
rect -1500 43420 -1480 43580
rect -1120 43420 -1100 43580
rect -1500 42880 -1100 43420
rect -1500 42720 -1480 42880
rect -1120 42720 -1100 42880
rect -1500 42700 -1100 42720
rect -3300 33400 -3200 34600
rect -1900 33400 -1800 34600
rect -3300 33300 -1800 33400
rect -800 36800 700 44300
rect 1000 43800 2700 43900
rect 1000 43500 1100 43800
rect 2600 43500 2700 43800
rect 1000 43400 2700 43500
rect 1000 42900 2700 43000
rect 1000 42600 1100 42900
rect 2600 42600 2700 42900
rect 1000 42500 2700 42600
rect -800 35600 -700 36800
rect 600 35600 700 36800
rect -800 33800 700 35600
rect -800 32000 -700 33800
rect 600 32000 700 33800
rect 1100 42100 2600 42200
rect 1100 40300 1200 42100
rect 2500 40300 2600 42100
rect 1100 34600 2600 40300
rect 3000 39100 4500 48700
rect 5500 49900 7000 50000
rect 5500 47300 5600 49900
rect 6900 48700 7000 49900
rect 6800 47300 7000 48700
rect 5500 47200 7000 47300
rect 4800 43580 5200 43600
rect 4800 43420 4820 43580
rect 5180 43420 5200 43580
rect 4800 42880 5200 43420
rect 4800 42720 4820 42880
rect 5180 42720 5200 42880
rect 4800 42700 5200 42720
rect 3000 37300 3100 39100
rect 4400 37300 4500 39100
rect 3000 37200 4500 37300
rect 5500 42100 7000 42200
rect 5500 40300 5600 42100
rect 6900 40300 7000 42100
rect 5500 36800 7000 40300
rect 7400 39100 8900 50500
rect 7400 37300 7500 39100
rect 8800 37300 8900 39100
rect 7400 37200 8900 37300
rect 9300 46100 10800 46200
rect 9300 44300 9400 46100
rect 10700 44300 10800 46100
rect 5500 35600 5600 36800
rect 6900 35600 7000 36800
rect 5500 35500 7000 35600
rect 7400 36800 8900 36900
rect 7400 35600 7500 36800
rect 8800 35600 8900 36800
rect 1100 33400 1200 34600
rect 2500 33400 2600 34600
rect 1100 33300 2600 33400
rect 3000 34600 4500 34700
rect 3000 33400 3100 34600
rect 4400 33400 4500 34600
rect -800 31900 700 32000
rect -5200 22000 -5100 23800
rect -3800 22000 -3700 23800
rect -5200 21900 -3700 22000
rect -3300 30800 -1800 30900
rect -3300 29000 -3200 30800
rect -1900 29000 -1800 30800
rect -7100 20300 -7000 21500
rect -5700 20300 -5600 21500
rect -7100 20200 -5600 20300
rect -5200 21500 -3700 21600
rect -5200 20300 -5100 21500
rect -3800 20300 -3700 21500
rect -11500 18100 -11400 19300
rect -10100 18100 -10000 19300
rect -11500 18000 -10000 18100
rect -9600 19300 -8100 19400
rect -9600 18100 -9500 19300
rect -8200 18100 -8100 19300
rect -13400 16600 -11900 16700
rect -13400 15500 -11900 15600
rect -13400 13700 -13300 15500
rect -12000 13700 -11900 15500
rect -13400 7200 -11900 13700
rect -11600 13200 -9900 13300
rect -11600 12900 -11500 13200
rect -10000 12900 -9900 13200
rect -11600 12800 -9900 12900
rect -11600 12300 -9900 12400
rect -11600 12000 -11500 12300
rect -10000 12000 -9900 12300
rect -11600 11900 -9900 12000
rect -13400 6000 -13300 7200
rect -12000 6000 -11900 7200
rect -13400 5900 -11900 6000
rect -11500 11500 -10000 11600
rect -11500 9700 -11400 11500
rect -10100 9700 -10000 11500
rect -11500 5400 -10000 9700
rect -9600 8500 -8100 18100
rect -7100 19300 -5600 19400
rect -7100 16700 -7000 19300
rect -5700 18100 -5600 19300
rect -5800 16700 -5600 18100
rect -7100 16600 -5600 16700
rect -7800 12980 -7400 13000
rect -7800 12820 -7780 12980
rect -7420 12820 -7400 12980
rect -7800 12280 -7400 12820
rect -7800 12120 -7780 12280
rect -7420 12120 -7400 12280
rect -7800 12100 -7400 12120
rect -9600 6700 -9500 8500
rect -8200 6700 -8100 8500
rect -9600 6600 -8100 6700
rect -7100 11500 -5600 11600
rect -7100 9700 -7000 11500
rect -5700 9700 -5600 11500
rect -7100 7200 -5600 9700
rect -7100 6000 -7000 7200
rect -5700 6000 -5600 7200
rect -5200 8500 -3700 20300
rect -3300 19300 -1800 29000
rect -800 30800 700 30900
rect -800 29000 -700 30800
rect 600 29000 700 30800
rect -1500 28280 -1100 28300
rect -1500 28120 -1480 28280
rect -1120 28120 -1100 28280
rect -1500 27580 -1100 28120
rect -1500 27420 -1480 27580
rect -1120 27420 -1100 27580
rect -1500 27400 -1100 27420
rect -3300 18100 -3200 19300
rect -1900 18100 -1800 19300
rect -3300 18000 -1800 18100
rect -800 21500 700 29000
rect 1000 28500 2700 28600
rect 1000 28200 1100 28500
rect 2600 28200 2700 28500
rect 1000 28100 2700 28200
rect 1000 27600 2700 27700
rect 1000 27300 1100 27600
rect 2600 27300 2700 27600
rect 1000 27200 2700 27300
rect -800 20300 -700 21500
rect 600 20300 700 21500
rect -800 18500 700 20300
rect -800 16700 -700 18500
rect 600 16700 700 18500
rect 1100 26800 2600 26900
rect 1100 25000 1200 26800
rect 2500 25000 2600 26800
rect 1100 19300 2600 25000
rect 3000 23800 4500 33400
rect 5500 34600 7000 34700
rect 5500 32000 5600 34600
rect 6900 33400 7000 34600
rect 6800 32000 7000 33400
rect 5500 31900 7000 32000
rect 4800 28280 5200 28300
rect 4800 28120 4820 28280
rect 5180 28120 5200 28280
rect 4800 27580 5200 28120
rect 4800 27420 4820 27580
rect 5180 27420 5200 27580
rect 4800 27400 5200 27420
rect 3000 22000 3100 23800
rect 4400 22000 4500 23800
rect 3000 21900 4500 22000
rect 5500 26800 7000 26900
rect 5500 25000 5600 26800
rect 6900 25000 7000 26800
rect 5500 21500 7000 25000
rect 7400 23800 8900 35600
rect 9300 34600 10800 44300
rect 9300 33400 9400 34600
rect 10700 33400 10800 34600
rect 9300 33300 10800 33400
rect 7400 22000 7500 23800
rect 8800 22000 8900 23800
rect 7400 21900 8900 22000
rect 9300 30800 10800 30900
rect 9300 29000 9400 30800
rect 10700 29000 10800 30800
rect 5500 20300 5600 21500
rect 6900 20300 7000 21500
rect 5500 20200 7000 20300
rect 7400 21500 8900 21600
rect 7400 20300 7500 21500
rect 8800 20300 8900 21500
rect 1100 18100 1200 19300
rect 2500 18100 2600 19300
rect 1100 18000 2600 18100
rect 3000 19300 4500 19400
rect 3000 18100 3100 19300
rect 4400 18100 4500 19300
rect -800 16600 700 16700
rect -5200 6700 -5100 8500
rect -3800 6700 -3700 8500
rect -5200 6600 -3700 6700
rect -3300 15500 -1800 15600
rect -3300 13700 -3200 15500
rect -1900 13700 -1800 15500
rect -7100 5900 -5600 6000
rect -11500 4200 -11400 5400
rect -10100 4200 -10000 5400
rect -11500 4100 -10000 4200
rect -3300 5400 -1800 13700
rect -800 15500 700 15600
rect -800 13700 -700 15500
rect 600 13700 700 15500
rect -1500 12980 -1100 13000
rect -1500 12820 -1480 12980
rect -1120 12820 -1100 12980
rect -1500 12280 -1100 12820
rect -1500 12120 -1480 12280
rect -1120 12120 -1100 12280
rect -1500 12100 -1100 12120
rect -800 7200 700 13700
rect 1000 13200 2700 13300
rect 1000 12900 1100 13200
rect 2600 12900 2700 13200
rect 1000 12800 2700 12900
rect 1000 12300 2700 12400
rect 1000 12000 1100 12300
rect 2600 12000 2700 12300
rect 1000 11900 2700 12000
rect -800 6000 -700 7200
rect 600 6000 700 7200
rect -800 5900 700 6000
rect 1100 11500 2600 11600
rect 1100 9700 1200 11500
rect 2500 9700 2600 11500
rect -3300 4200 -3200 5400
rect -1900 4200 -1800 5400
rect -3300 4100 -1800 4200
rect 1100 5400 2600 9700
rect 3000 8500 4500 18100
rect 5500 19300 7000 19400
rect 5500 16700 5600 19300
rect 6900 18100 7000 19300
rect 6800 16700 7000 18100
rect 5500 16600 7000 16700
rect 4800 12980 5200 13000
rect 4800 12820 4820 12980
rect 5180 12820 5200 12980
rect 4800 12280 5200 12820
rect 4800 12120 4820 12280
rect 5180 12120 5200 12280
rect 4800 12100 5200 12120
rect 3000 6700 3100 8500
rect 4400 6700 4500 8500
rect 3000 6600 4500 6700
rect 5500 11500 7000 11600
rect 5500 9700 5600 11500
rect 6900 9700 7000 11500
rect 5500 7200 7000 9700
rect 5500 6000 5600 7200
rect 6900 6000 7000 7200
rect 7400 8500 8900 20300
rect 9300 19300 10800 29000
rect 9300 18100 9400 19300
rect 10700 18100 10800 19300
rect 9300 18000 10800 18100
rect 7400 6700 7500 8500
rect 8800 6700 8900 8500
rect 7400 6600 8900 6700
rect 9300 15500 10800 15600
rect 9300 13700 9400 15500
rect 10700 13700 10800 15500
rect 5500 5900 7000 6000
rect 1100 4200 1200 5400
rect 2500 4200 2600 5400
rect 1100 4100 2600 4200
rect 9300 5400 10800 13700
rect 9300 4200 9400 5400
rect 10700 4200 10800 5400
rect 9300 4100 10800 4200
<< via4 >>
rect -13300 50500 -12000 51700
rect -5100 50500 -3800 51700
rect -9500 48700 -8200 49900
rect -11500 43500 -10000 43800
rect -11500 42600 -10000 42900
rect -13300 35600 -12000 36800
rect -7000 49100 -5700 49900
rect -7000 48700 -5800 49100
rect -5800 48700 -5700 49100
rect -700 50500 600 51700
rect 7500 50500 8800 51700
rect 3100 48700 4400 49900
rect -7000 35600 -5700 36800
rect -5100 35600 -3800 36800
rect -11400 33400 -10100 34600
rect -9500 33400 -8200 34600
rect -11500 28200 -10000 28500
rect -11500 27300 -10000 27600
rect -13300 20300 -12000 21500
rect -7000 33800 -5700 34600
rect -7000 33400 -5800 33800
rect -5800 33400 -5700 33800
rect -3200 33400 -1900 34600
rect 1100 43500 2600 43800
rect 1100 42600 2600 42900
rect -700 35600 600 36800
rect 5600 49100 6900 49900
rect 5600 48700 6800 49100
rect 6800 48700 6900 49100
rect 5600 35600 6900 36800
rect 7500 35600 8800 36800
rect 1200 33400 2500 34600
rect 3100 33400 4400 34600
rect -7000 20300 -5700 21500
rect -5100 20300 -3800 21500
rect -11400 18100 -10100 19300
rect -9500 18100 -8200 19300
rect -11500 12900 -10000 13200
rect -11500 12000 -10000 12300
rect -13300 6000 -12000 7200
rect -7000 18500 -5700 19300
rect -7000 18100 -5800 18500
rect -5800 18100 -5700 18500
rect -7000 6000 -5700 7200
rect -3200 18100 -1900 19300
rect 1100 28200 2600 28500
rect 1100 27300 2600 27600
rect -700 20300 600 21500
rect 5600 33800 6900 34600
rect 5600 33400 6800 33800
rect 6800 33400 6900 33800
rect 9400 33400 10700 34600
rect 5600 20300 6900 21500
rect 7500 20300 8800 21500
rect 1200 18100 2500 19300
rect 3100 18100 4400 19300
rect -11400 4200 -10100 5400
rect 1100 12900 2600 13200
rect 1100 12000 2600 12300
rect -700 6000 600 7200
rect -3200 4200 -1900 5400
rect 5600 18500 6900 19300
rect 5600 18100 6800 18500
rect 6800 18100 6900 18500
rect 5600 6000 6900 7200
rect 9400 18100 10700 19300
rect 1200 4200 2500 5400
rect 9400 4200 10700 5400
<< metal5 >>
rect -13400 51800 -11900 52200
rect -13400 51700 8900 51800
rect -13400 50500 -13300 51700
rect -12000 50500 -5100 51700
rect -3800 50500 -700 51700
rect 600 50500 7500 51700
rect 8800 50500 8900 51700
rect -13400 50400 8900 50500
rect 9300 50000 10800 52200
rect -9600 49900 10800 50000
rect -9600 48700 -9500 49900
rect -8200 48700 -7000 49900
rect -5700 48700 3100 49900
rect 4400 48700 5600 49900
rect 6900 48700 10800 49900
rect -9600 48600 10800 48700
rect -13500 43800 10700 43900
rect -13500 43500 -11500 43800
rect -10000 43500 1100 43800
rect 2600 43500 10700 43800
rect -13500 43400 10700 43500
rect -13500 42900 10700 43000
rect -13500 42600 -11500 42900
rect -10000 42600 1100 42900
rect 2600 42600 10700 42900
rect -13500 42500 10700 42600
rect -13400 36800 10800 36900
rect -13400 35600 -13300 36800
rect -12000 35600 -7000 36800
rect -5700 35600 -5100 36800
rect -3800 35600 -700 36800
rect 600 35600 5600 36800
rect 6900 35600 7500 36800
rect 8800 35600 10800 36800
rect -13400 35500 10800 35600
rect -13400 34600 10800 34700
rect -13400 33400 -11400 34600
rect -10100 33400 -9500 34600
rect -8200 33400 -7000 34600
rect -5700 33400 -3200 34600
rect -1900 33400 1200 34600
rect 2500 33400 3100 34600
rect 4400 33400 5600 34600
rect 6900 33400 9400 34600
rect 10700 33400 10800 34600
rect -13400 33300 10800 33400
rect -13500 28500 10700 28600
rect -13500 28200 -11500 28500
rect -10000 28200 1100 28500
rect 2600 28200 10700 28500
rect -13500 28100 10700 28200
rect -13500 27600 10700 27700
rect -13500 27300 -11500 27600
rect -10000 27300 1100 27600
rect 2600 27300 10700 27600
rect -13500 27200 10700 27300
rect -13400 21500 10800 21600
rect -13400 20300 -13300 21500
rect -12000 20300 -7000 21500
rect -5700 20300 -5100 21500
rect -3800 20300 -700 21500
rect 600 20300 5600 21500
rect 6900 20300 7500 21500
rect 8800 20300 10800 21500
rect -13400 20200 10800 20300
rect -13400 19300 10800 19400
rect -13400 18100 -11400 19300
rect -10100 18100 -9500 19300
rect -8200 18100 -7000 19300
rect -5700 18100 -3200 19300
rect -1900 18100 1200 19300
rect 2500 18100 3100 19300
rect 4400 18100 5600 19300
rect 6900 18100 9400 19300
rect 10700 18100 10800 19300
rect -13400 18000 10800 18100
rect -13500 13200 10700 13300
rect -13500 12900 -11500 13200
rect -10000 12900 1100 13200
rect 2600 12900 10700 13200
rect -13500 12800 10700 12900
rect -13500 12300 10700 12400
rect -13500 12000 -11500 12300
rect -10000 12000 1100 12300
rect 2600 12000 10700 12300
rect -13500 11900 10700 12000
rect -13400 7200 7000 7300
rect -13400 6000 -13300 7200
rect -12000 6000 -7000 7200
rect -5700 6000 -700 7200
rect 600 6000 5600 7200
rect 6900 6000 7000 7200
rect -13400 5900 7000 6000
rect -13400 3700 -11900 5900
rect -11500 5400 10800 5500
rect -11500 4200 -11400 5400
rect -10100 4200 -3200 5400
rect -1900 4200 1200 5400
rect 2500 4200 9400 5400
rect 10700 4200 10800 5400
rect -11500 4100 10800 4200
rect 9300 3700 10800 4100
<< comment >>
rect -13400 50100 -13300 50300
rect -9600 50200 -9400 50300
rect -7100 50200 -6900 50300
rect -5200 50200 -5100 50400
rect -13400 50000 -13200 50100
rect -9600 50012 -9500 50200
rect -7100 50012 -7000 50200
rect -5200 50100 -5000 50200
rect -700 50100 -600 50300
rect 3000 50200 3200 50300
rect 5500 50200 5700 50300
rect 7400 50200 7500 50400
rect -700 50000 -500 50100
rect 3000 50012 3100 50200
rect 5500 50012 5600 50200
rect 7400 50100 7600 50200
rect -14500 49800 -14400 49900
rect -14600 49600 -14500 49800
rect -14400 49600 -14300 49700
rect -14600 49500 -14300 49600
rect -14400 49400 -14300 49500
rect -13400 36200 -13300 36400
rect -11500 36300 -11300 36400
rect -13400 36100 -13200 36200
rect -11500 36112 -11400 36300
rect -7100 36200 -7000 36400
rect -3300 36300 -3100 36400
rect -7100 36100 -6900 36200
rect -3300 36112 -3200 36300
rect -800 36200 -700 36400
rect 1100 36300 1300 36400
rect -800 36100 -600 36200
rect 1100 36112 1200 36300
rect 5500 36200 5600 36400
rect 9300 36300 9500 36400
rect 5500 36100 5700 36200
rect 9300 36112 9400 36300
rect -14700 35100 -14400 35200
rect -14500 35000 -14400 35100
rect -14600 34900 -14400 35000
rect -14500 34800 -14400 34900
rect -14700 34700 -14400 34800
rect -13400 34800 -13300 35000
rect -9600 34900 -9400 35000
rect -7100 34900 -6900 35000
rect -5200 34900 -5100 35100
rect -13400 34700 -13200 34800
rect -9600 34712 -9500 34900
rect -7100 34712 -7000 34900
rect -5200 34800 -5000 34900
rect -700 34800 -600 35000
rect 3000 34900 3200 35000
rect 5500 34900 5700 35000
rect 7400 34900 7500 35100
rect -700 34700 -500 34800
rect 3000 34712 3100 34900
rect 5500 34712 5600 34900
rect 7400 34800 7600 34900
rect -13400 20900 -13300 21100
rect -11500 21000 -11300 21100
rect -13400 20800 -13200 20900
rect -11500 20812 -11400 21000
rect -7100 20900 -7000 21100
rect -3300 21000 -3100 21100
rect -7100 20800 -6900 20900
rect -3300 20812 -3200 21000
rect -800 20900 -700 21100
rect 1100 21000 1300 21100
rect -800 20800 -600 20900
rect 1100 20812 1200 21000
rect 5500 20900 5600 21100
rect 9300 21000 9500 21100
rect 5500 20800 5700 20900
rect 9300 20812 9400 21000
rect -13400 19500 -13300 19700
rect -9600 19600 -9400 19700
rect -7100 19600 -6900 19700
rect -5200 19600 -5100 19800
rect -13400 19400 -13200 19500
rect -9600 19412 -9500 19600
rect -7100 19412 -7000 19600
rect -5200 19500 -5000 19600
rect -700 19500 -600 19700
rect 3000 19600 3200 19700
rect 5500 19600 5700 19700
rect 7400 19600 7500 19800
rect -700 19400 -500 19500
rect 3000 19412 3100 19600
rect 5500 19412 5600 19600
rect 7400 19500 7600 19600
rect -14600 19300 -14300 19400
rect -14400 19200 -14300 19300
rect -14500 19100 -14300 19200
rect -14600 19000 -14500 19100
rect -14600 18900 -14300 19000
rect -13400 5600 -13300 5800
rect -11500 5700 -11300 5800
rect -13400 5500 -13200 5600
rect -11500 5512 -11400 5700
rect -7100 5600 -7000 5800
rect -3300 5700 -3100 5800
rect -7100 5500 -6900 5600
rect -3300 5512 -3200 5700
rect -800 5600 -700 5800
rect 1100 5700 1300 5800
rect -800 5500 -600 5600
rect 1100 5512 1200 5700
rect 5500 5600 5600 5800
rect 9300 5700 9500 5800
rect 5500 5500 5700 5600
rect 9300 5512 9400 5700
rect -14300 4500 -14200 4600
rect -14400 4400 -14200 4500
rect -14300 4200 -14200 4400
rect -14400 4100 -14100 4200
<< labels >>
rlabel metal5 -13400 3700 -11900 4100 1 SD1L
rlabel metal5 9300 3700 10800 4100 1 SD1R
rlabel metal5 -13400 18000 -13100 19400 1 SD2R
rlabel metal5 -13400 20200 -13100 21600 1 SD2L
rlabel metal5 -13400 33300 -13100 34700 1 SD3R
rlabel metal5 -13400 35500 -13100 36900 1 SD3L
rlabel metal5 -13400 51800 -11900 52200 1 SD4L
rlabel metal5 9300 51800 10800 52200 1 SD4R
rlabel metal5 -13500 12800 -13400 13300 1 G12L
rlabel metal5 -13500 11900 -13400 12400 1 G12R
rlabel metal5 -13500 27200 -13400 27700 1 G23R
rlabel metal5 -13500 28100 -13400 28600 1 G23L
rlabel metal5 -13500 42500 -13400 43000 1 G34R
rlabel metal5 -13500 43400 -13400 43900 1 G34L
<< end >>
