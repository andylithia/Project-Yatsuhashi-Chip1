magic
tech sky130B
timestamp 1658699409
<< metal4 >>
rect 1700 -2750 2200 -150
rect 1700 -2900 1750 -2750
rect 1900 -2900 1950 -2750
rect 2100 -2900 2200 -2750
rect 1700 -2950 2200 -2900
rect 1700 -3100 1800 -2950
rect 1950 -3100 2000 -2950
rect 2150 -3100 2200 -2950
rect 1700 -3200 2200 -3100
<< via4 >>
rect 1750 -2900 1900 -2750
rect 1950 -2900 2100 -2750
rect 1800 -3100 1950 -2950
rect 2000 -3100 2150 -2950
<< metal5 >>
rect 100 -800 6600 -300
rect 100 -1600 5800 -1100
rect 100 -6300 600 -1600
rect 900 -2400 5000 -1900
rect 900 -5500 1400 -2400
rect 1700 -2750 2200 -2700
rect 1700 -2900 1750 -2750
rect 1900 -2900 1950 -2750
rect 2100 -2900 2200 -2750
rect 1700 -2950 2200 -2900
rect 1700 -3100 1800 -2950
rect 1950 -3100 2000 -2950
rect 2150 -3100 2200 -2950
rect 1700 -4600 2200 -3100
rect 4500 -4600 5000 -2400
rect 1700 -5200 5000 -4600
rect 5300 -5500 5800 -1600
rect 900 -6000 5800 -5500
rect 6100 -6300 6600 -800
rect 100 -6800 6600 -6300
<< labels >>
rlabel metal4 1700 -300 2200 -150 1 B
rlabel metal5 100 -800 350 -300 1 A
<< end >>
