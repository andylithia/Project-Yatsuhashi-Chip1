magic
tech sky130B
magscale 1 2
timestamp 1659840519
<< error_p >>
rect 3188 3291 3246 3297
rect 3306 3291 3364 3297
rect 3424 3291 3482 3297
rect 3542 3291 3600 3297
rect 3660 3291 3718 3297
rect 3778 3291 3836 3297
rect 3896 3291 3954 3297
rect 4014 3291 4072 3297
rect 3188 3257 3200 3291
rect 3306 3257 3318 3291
rect 3424 3257 3436 3291
rect 3542 3257 3554 3291
rect 3660 3257 3672 3291
rect 3778 3257 3790 3291
rect 3896 3257 3908 3291
rect 4014 3257 4026 3291
rect 3188 3251 3246 3257
rect 3306 3251 3364 3257
rect 3424 3251 3482 3257
rect 3542 3251 3600 3257
rect 3660 3251 3718 3257
rect 3778 3251 3836 3257
rect 3896 3251 3954 3257
rect 4014 3251 4072 3257
rect 3188 2419 3246 2425
rect 3188 2385 3200 2419
rect 3188 2379 3246 2385
<< nwell >>
rect 2047 2247 5213 3757
<< pmos >>
rect 2243 3338 2303 3538
rect 2361 3338 2421 3538
rect 2479 3338 2539 3538
rect 2597 3338 2657 3538
rect 2715 3338 2775 3538
rect 2833 3338 2893 3538
rect 2951 3338 3011 3538
rect 3069 3338 3129 3538
rect 3187 3338 3247 3538
rect 3305 3338 3365 3538
rect 3423 3338 3483 3538
rect 3541 3338 3601 3538
rect 3659 3338 3719 3538
rect 3777 3338 3837 3538
rect 3895 3338 3955 3538
rect 4013 3338 4073 3538
rect 4131 3338 4191 3538
rect 4249 3338 4309 3538
rect 4367 3338 4427 3538
rect 4485 3338 4545 3538
rect 4603 3338 4663 3538
rect 4721 3338 4781 3538
rect 4839 3338 4899 3538
rect 4957 3338 5017 3538
rect 2243 2902 2303 3102
rect 2361 2902 2421 3102
rect 2479 2902 2539 3102
rect 2597 2902 2657 3102
rect 2715 2902 2775 3102
rect 2833 2902 2893 3102
rect 2951 2902 3011 3102
rect 3069 2902 3129 3102
rect 3187 2902 3247 3102
rect 3305 2902 3365 3102
rect 3423 2902 3483 3102
rect 3541 2902 3601 3102
rect 3659 2902 3719 3102
rect 3777 2902 3837 3102
rect 3895 2902 3955 3102
rect 4013 2902 4073 3102
rect 4131 2902 4191 3102
rect 4249 2902 4309 3102
rect 4367 2902 4427 3102
rect 4485 2902 4545 3102
rect 4603 2902 4663 3102
rect 4721 2902 4781 3102
rect 4839 2902 4899 3102
rect 4957 2902 5017 3102
rect 2243 2466 2303 2666
rect 2361 2466 2421 2666
rect 2479 2466 2539 2666
rect 2597 2466 2657 2666
rect 2715 2466 2775 2666
rect 2833 2466 2893 2666
rect 2951 2466 3011 2666
rect 3069 2466 3129 2666
rect 3187 2466 3247 2666
rect 3305 2466 3365 2666
rect 3423 2466 3483 2666
rect 3541 2466 3601 2666
rect 3659 2466 3719 2666
rect 3777 2466 3837 2666
rect 3895 2466 3955 2666
rect 4013 2466 4073 2666
rect 4131 2466 4191 2666
rect 4249 2466 4309 2666
rect 4367 2466 4427 2666
rect 4485 2466 4545 2666
rect 4603 2466 4663 2666
rect 4721 2466 4781 2666
rect 4839 2466 4899 2666
rect 4957 2466 5017 2666
<< pdiff >>
rect 2185 3526 2243 3538
rect 2185 3350 2197 3526
rect 2231 3350 2243 3526
rect 2185 3338 2243 3350
rect 2303 3526 2361 3538
rect 2303 3350 2315 3526
rect 2349 3350 2361 3526
rect 2303 3338 2361 3350
rect 2421 3526 2479 3538
rect 2421 3350 2433 3526
rect 2467 3350 2479 3526
rect 2421 3338 2479 3350
rect 2539 3526 2597 3538
rect 2539 3350 2551 3526
rect 2585 3350 2597 3526
rect 2539 3338 2597 3350
rect 2657 3526 2715 3538
rect 2657 3350 2669 3526
rect 2703 3350 2715 3526
rect 2657 3338 2715 3350
rect 2775 3526 2833 3538
rect 2775 3350 2787 3526
rect 2821 3350 2833 3526
rect 2775 3338 2833 3350
rect 2893 3526 2951 3538
rect 2893 3350 2905 3526
rect 2939 3350 2951 3526
rect 2893 3338 2951 3350
rect 3011 3526 3069 3538
rect 3011 3350 3023 3526
rect 3057 3350 3069 3526
rect 3011 3338 3069 3350
rect 3129 3526 3187 3538
rect 3129 3350 3141 3526
rect 3175 3350 3187 3526
rect 3129 3338 3187 3350
rect 3247 3526 3305 3538
rect 3247 3350 3259 3526
rect 3293 3350 3305 3526
rect 3247 3338 3305 3350
rect 3365 3526 3423 3538
rect 3365 3350 3377 3526
rect 3411 3350 3423 3526
rect 3365 3338 3423 3350
rect 3483 3526 3541 3538
rect 3483 3350 3495 3526
rect 3529 3350 3541 3526
rect 3483 3338 3541 3350
rect 3601 3526 3659 3538
rect 3601 3350 3613 3526
rect 3647 3350 3659 3526
rect 3601 3338 3659 3350
rect 3719 3526 3777 3538
rect 3719 3350 3731 3526
rect 3765 3350 3777 3526
rect 3719 3338 3777 3350
rect 3837 3526 3895 3538
rect 3837 3350 3849 3526
rect 3883 3350 3895 3526
rect 3837 3338 3895 3350
rect 3955 3526 4013 3538
rect 3955 3350 3967 3526
rect 4001 3350 4013 3526
rect 3955 3338 4013 3350
rect 4073 3526 4131 3538
rect 4073 3350 4085 3526
rect 4119 3350 4131 3526
rect 4073 3338 4131 3350
rect 4191 3526 4249 3538
rect 4191 3350 4203 3526
rect 4237 3350 4249 3526
rect 4191 3338 4249 3350
rect 4309 3526 4367 3538
rect 4309 3350 4321 3526
rect 4355 3350 4367 3526
rect 4309 3338 4367 3350
rect 4427 3526 4485 3538
rect 4427 3350 4439 3526
rect 4473 3350 4485 3526
rect 4427 3338 4485 3350
rect 4545 3526 4603 3538
rect 4545 3350 4557 3526
rect 4591 3350 4603 3526
rect 4545 3338 4603 3350
rect 4663 3526 4721 3538
rect 4663 3350 4675 3526
rect 4709 3350 4721 3526
rect 4663 3338 4721 3350
rect 4781 3526 4839 3538
rect 4781 3350 4793 3526
rect 4827 3350 4839 3526
rect 4781 3338 4839 3350
rect 4899 3526 4957 3538
rect 4899 3350 4911 3526
rect 4945 3350 4957 3526
rect 4899 3338 4957 3350
rect 5017 3526 5075 3538
rect 5017 3350 5029 3526
rect 5063 3350 5075 3526
rect 5017 3338 5075 3350
rect 2185 3090 2243 3102
rect 2185 2914 2197 3090
rect 2231 2914 2243 3090
rect 2185 2902 2243 2914
rect 2303 3090 2361 3102
rect 2303 2914 2315 3090
rect 2349 2914 2361 3090
rect 2303 2902 2361 2914
rect 2421 3090 2479 3102
rect 2421 2914 2433 3090
rect 2467 2914 2479 3090
rect 2421 2902 2479 2914
rect 2539 3090 2597 3102
rect 2539 2914 2551 3090
rect 2585 2914 2597 3090
rect 2539 2902 2597 2914
rect 2657 3090 2715 3102
rect 2657 2914 2669 3090
rect 2703 2914 2715 3090
rect 2657 2902 2715 2914
rect 2775 3090 2833 3102
rect 2775 2914 2787 3090
rect 2821 2914 2833 3090
rect 2775 2902 2833 2914
rect 2893 3090 2951 3102
rect 2893 2914 2905 3090
rect 2939 2914 2951 3090
rect 2893 2902 2951 2914
rect 3011 3090 3069 3102
rect 3011 2914 3023 3090
rect 3057 2914 3069 3090
rect 3011 2902 3069 2914
rect 3129 3090 3187 3102
rect 3129 2914 3141 3090
rect 3175 2914 3187 3090
rect 3129 2902 3187 2914
rect 3247 3090 3305 3102
rect 3247 2914 3259 3090
rect 3293 2914 3305 3090
rect 3247 2902 3305 2914
rect 3365 3090 3423 3102
rect 3365 2914 3377 3090
rect 3411 2914 3423 3090
rect 3365 2902 3423 2914
rect 3483 3090 3541 3102
rect 3483 2914 3495 3090
rect 3529 2914 3541 3090
rect 3483 2902 3541 2914
rect 3601 3090 3659 3102
rect 3601 2914 3613 3090
rect 3647 2914 3659 3090
rect 3601 2902 3659 2914
rect 3719 3090 3777 3102
rect 3719 2914 3731 3090
rect 3765 2914 3777 3090
rect 3719 2902 3777 2914
rect 3837 3090 3895 3102
rect 3837 2914 3849 3090
rect 3883 2914 3895 3090
rect 3837 2902 3895 2914
rect 3955 3090 4013 3102
rect 3955 2914 3967 3090
rect 4001 2914 4013 3090
rect 3955 2902 4013 2914
rect 4073 3090 4131 3102
rect 4073 2914 4085 3090
rect 4119 2914 4131 3090
rect 4073 2902 4131 2914
rect 4191 3090 4249 3102
rect 4191 2914 4203 3090
rect 4237 2914 4249 3090
rect 4191 2902 4249 2914
rect 4309 3090 4367 3102
rect 4309 2914 4321 3090
rect 4355 2914 4367 3090
rect 4309 2902 4367 2914
rect 4427 3090 4485 3102
rect 4427 2914 4439 3090
rect 4473 2914 4485 3090
rect 4427 2902 4485 2914
rect 4545 3090 4603 3102
rect 4545 2914 4557 3090
rect 4591 2914 4603 3090
rect 4545 2902 4603 2914
rect 4663 3090 4721 3102
rect 4663 2914 4675 3090
rect 4709 2914 4721 3090
rect 4663 2902 4721 2914
rect 4781 3090 4839 3102
rect 4781 2914 4793 3090
rect 4827 2914 4839 3090
rect 4781 2902 4839 2914
rect 4899 3090 4957 3102
rect 4899 2914 4911 3090
rect 4945 2914 4957 3090
rect 4899 2902 4957 2914
rect 5017 3090 5075 3102
rect 5017 2914 5029 3090
rect 5063 2914 5075 3090
rect 5017 2902 5075 2914
rect 2185 2654 2243 2666
rect 2185 2478 2197 2654
rect 2231 2478 2243 2654
rect 2185 2466 2243 2478
rect 2303 2654 2361 2666
rect 2303 2478 2315 2654
rect 2349 2478 2361 2654
rect 2303 2466 2361 2478
rect 2421 2654 2479 2666
rect 2421 2478 2433 2654
rect 2467 2478 2479 2654
rect 2421 2466 2479 2478
rect 2539 2654 2597 2666
rect 2539 2478 2551 2654
rect 2585 2478 2597 2654
rect 2539 2466 2597 2478
rect 2657 2654 2715 2666
rect 2657 2478 2669 2654
rect 2703 2478 2715 2654
rect 2657 2466 2715 2478
rect 2775 2654 2833 2666
rect 2775 2478 2787 2654
rect 2821 2478 2833 2654
rect 2775 2466 2833 2478
rect 2893 2654 2951 2666
rect 2893 2478 2905 2654
rect 2939 2478 2951 2654
rect 2893 2466 2951 2478
rect 3011 2654 3069 2666
rect 3011 2478 3023 2654
rect 3057 2478 3069 2654
rect 3011 2466 3069 2478
rect 3129 2654 3187 2666
rect 3129 2478 3141 2654
rect 3175 2478 3187 2654
rect 3129 2466 3187 2478
rect 3247 2654 3305 2666
rect 3247 2478 3259 2654
rect 3293 2478 3305 2654
rect 3247 2466 3305 2478
rect 3365 2654 3423 2666
rect 3365 2478 3377 2654
rect 3411 2478 3423 2654
rect 3365 2466 3423 2478
rect 3483 2654 3541 2666
rect 3483 2478 3495 2654
rect 3529 2478 3541 2654
rect 3483 2466 3541 2478
rect 3601 2654 3659 2666
rect 3601 2478 3613 2654
rect 3647 2478 3659 2654
rect 3601 2466 3659 2478
rect 3719 2654 3777 2666
rect 3719 2478 3731 2654
rect 3765 2478 3777 2654
rect 3719 2466 3777 2478
rect 3837 2654 3895 2666
rect 3837 2478 3849 2654
rect 3883 2478 3895 2654
rect 3837 2466 3895 2478
rect 3955 2654 4013 2666
rect 3955 2478 3967 2654
rect 4001 2478 4013 2654
rect 3955 2466 4013 2478
rect 4073 2654 4131 2666
rect 4073 2478 4085 2654
rect 4119 2478 4131 2654
rect 4073 2466 4131 2478
rect 4191 2654 4249 2666
rect 4191 2478 4203 2654
rect 4237 2478 4249 2654
rect 4191 2466 4249 2478
rect 4309 2654 4367 2666
rect 4309 2478 4321 2654
rect 4355 2478 4367 2654
rect 4309 2466 4367 2478
rect 4427 2654 4485 2666
rect 4427 2478 4439 2654
rect 4473 2478 4485 2654
rect 4427 2466 4485 2478
rect 4545 2654 4603 2666
rect 4545 2478 4557 2654
rect 4591 2478 4603 2654
rect 4545 2466 4603 2478
rect 4663 2654 4721 2666
rect 4663 2478 4675 2654
rect 4709 2478 4721 2654
rect 4663 2466 4721 2478
rect 4781 2654 4839 2666
rect 4781 2478 4793 2654
rect 4827 2478 4839 2654
rect 4781 2466 4839 2478
rect 4899 2654 4957 2666
rect 4899 2478 4911 2654
rect 4945 2478 4957 2654
rect 4899 2466 4957 2478
rect 5017 2654 5075 2666
rect 5017 2478 5029 2654
rect 5063 2478 5075 2654
rect 5017 2466 5075 2478
<< pdiffc >>
rect 2197 3350 2231 3526
rect 2315 3350 2349 3526
rect 2433 3350 2467 3526
rect 2551 3350 2585 3526
rect 2669 3350 2703 3526
rect 2787 3350 2821 3526
rect 2905 3350 2939 3526
rect 3023 3350 3057 3526
rect 3141 3350 3175 3526
rect 3259 3350 3293 3526
rect 3377 3350 3411 3526
rect 3495 3350 3529 3526
rect 3613 3350 3647 3526
rect 3731 3350 3765 3526
rect 3849 3350 3883 3526
rect 3967 3350 4001 3526
rect 4085 3350 4119 3526
rect 4203 3350 4237 3526
rect 4321 3350 4355 3526
rect 4439 3350 4473 3526
rect 4557 3350 4591 3526
rect 4675 3350 4709 3526
rect 4793 3350 4827 3526
rect 4911 3350 4945 3526
rect 5029 3350 5063 3526
rect 2197 2914 2231 3090
rect 2315 2914 2349 3090
rect 2433 2914 2467 3090
rect 2551 2914 2585 3090
rect 2669 2914 2703 3090
rect 2787 2914 2821 3090
rect 2905 2914 2939 3090
rect 3023 2914 3057 3090
rect 3141 2914 3175 3090
rect 3259 2914 3293 3090
rect 3377 2914 3411 3090
rect 3495 2914 3529 3090
rect 3613 2914 3647 3090
rect 3731 2914 3765 3090
rect 3849 2914 3883 3090
rect 3967 2914 4001 3090
rect 4085 2914 4119 3090
rect 4203 2914 4237 3090
rect 4321 2914 4355 3090
rect 4439 2914 4473 3090
rect 4557 2914 4591 3090
rect 4675 2914 4709 3090
rect 4793 2914 4827 3090
rect 4911 2914 4945 3090
rect 5029 2914 5063 3090
rect 2197 2478 2231 2654
rect 2315 2478 2349 2654
rect 2433 2478 2467 2654
rect 2551 2478 2585 2654
rect 2669 2478 2703 2654
rect 2787 2478 2821 2654
rect 2905 2478 2939 2654
rect 3023 2478 3057 2654
rect 3141 2478 3175 2654
rect 3259 2478 3293 2654
rect 3377 2478 3411 2654
rect 3495 2478 3529 2654
rect 3613 2478 3647 2654
rect 3731 2478 3765 2654
rect 3849 2478 3883 2654
rect 3967 2478 4001 2654
rect 4085 2478 4119 2654
rect 4203 2478 4237 2654
rect 4321 2478 4355 2654
rect 4439 2478 4473 2654
rect 4557 2478 4591 2654
rect 4675 2478 4709 2654
rect 4793 2478 4827 2654
rect 4911 2478 4945 2654
rect 5029 2478 5063 2654
<< nsubdiff >>
rect 2083 3687 2179 3721
rect 5081 3687 5177 3721
rect 2083 3625 2117 3687
rect 5143 3625 5177 3687
rect 2083 2317 2117 2379
rect 5143 2317 5177 2379
rect 2083 2283 2179 2317
rect 5081 2283 5177 2317
<< nsubdiffcont >>
rect 2179 3687 5081 3721
rect 2083 2379 2117 3625
rect 5143 2379 5177 3625
rect 2179 2283 5081 2317
<< poly >>
rect 2243 3538 2303 3569
rect 2361 3538 2421 3569
rect 2479 3538 2539 3569
rect 2597 3538 2657 3569
rect 2715 3538 2775 3569
rect 2833 3538 2893 3569
rect 2951 3538 3011 3569
rect 3069 3538 3129 3569
rect 3187 3538 3247 3569
rect 3305 3538 3365 3569
rect 3423 3538 3483 3569
rect 3541 3538 3601 3569
rect 3659 3538 3719 3569
rect 3777 3538 3837 3569
rect 3895 3538 3955 3569
rect 4013 3538 4073 3569
rect 4131 3538 4191 3569
rect 4249 3538 4309 3569
rect 4367 3538 4427 3569
rect 4485 3538 4545 3569
rect 4603 3538 4663 3569
rect 4721 3538 4781 3569
rect 4839 3538 4899 3569
rect 4957 3538 5017 3569
rect 2243 3307 2303 3338
rect 2361 3307 2421 3338
rect 2479 3307 2539 3338
rect 2597 3307 2657 3338
rect 2715 3307 2775 3338
rect 2833 3307 2893 3338
rect 2951 3307 3011 3338
rect 3069 3307 3129 3338
rect 3187 3307 3247 3338
rect 3305 3307 3365 3338
rect 3423 3307 3483 3338
rect 3541 3307 3601 3338
rect 3659 3307 3719 3338
rect 3777 3307 3837 3338
rect 3895 3307 3955 3338
rect 4013 3307 4073 3338
rect 4131 3307 4191 3338
rect 4249 3307 4309 3338
rect 4367 3307 4427 3338
rect 4485 3307 4545 3338
rect 4603 3307 4663 3338
rect 4721 3307 4781 3338
rect 4839 3307 4899 3338
rect 4957 3307 5017 3338
rect 2240 3291 2306 3307
rect 2240 3257 2256 3291
rect 2290 3257 2306 3291
rect 2240 3241 2306 3257
rect 2358 3291 2424 3307
rect 2358 3257 2374 3291
rect 2408 3257 2424 3291
rect 2358 3241 2424 3257
rect 2476 3291 2542 3307
rect 2476 3257 2492 3291
rect 2526 3257 2542 3291
rect 2476 3241 2542 3257
rect 2594 3291 2660 3307
rect 2594 3257 2610 3291
rect 2644 3257 2660 3291
rect 2594 3241 2660 3257
rect 2712 3291 2778 3307
rect 2712 3257 2728 3291
rect 2762 3257 2778 3291
rect 2712 3241 2778 3257
rect 2830 3291 2896 3307
rect 2830 3257 2846 3291
rect 2880 3257 2896 3291
rect 2830 3241 2896 3257
rect 2948 3291 3014 3307
rect 2948 3257 2964 3291
rect 2998 3257 3014 3291
rect 2948 3241 3014 3257
rect 3066 3291 3132 3307
rect 3066 3257 3082 3291
rect 3116 3257 3132 3291
rect 3066 3241 3132 3257
rect 3184 3291 3250 3307
rect 3184 3257 3200 3291
rect 3234 3257 3250 3291
rect 3184 3241 3250 3257
rect 3302 3291 3368 3307
rect 3302 3257 3318 3291
rect 3352 3257 3368 3291
rect 3302 3241 3368 3257
rect 3420 3291 3486 3307
rect 3420 3257 3436 3291
rect 3470 3257 3486 3291
rect 3420 3241 3486 3257
rect 3538 3291 3604 3307
rect 3538 3257 3554 3291
rect 3588 3257 3604 3291
rect 3538 3241 3604 3257
rect 3656 3291 3722 3307
rect 3656 3257 3672 3291
rect 3706 3257 3722 3291
rect 3656 3241 3722 3257
rect 3774 3291 3840 3307
rect 3774 3257 3790 3291
rect 3824 3257 3840 3291
rect 3774 3241 3840 3257
rect 3892 3291 3958 3307
rect 3892 3257 3908 3291
rect 3942 3257 3958 3291
rect 3892 3241 3958 3257
rect 4010 3291 4076 3307
rect 4010 3257 4026 3291
rect 4060 3257 4076 3291
rect 4010 3241 4076 3257
rect 4128 3291 4194 3307
rect 4128 3257 4144 3291
rect 4178 3257 4194 3291
rect 4128 3241 4194 3257
rect 4246 3291 4312 3307
rect 4246 3257 4262 3291
rect 4296 3257 4312 3291
rect 4246 3241 4312 3257
rect 4364 3291 4430 3307
rect 4364 3257 4380 3291
rect 4414 3257 4430 3291
rect 4364 3241 4430 3257
rect 4482 3291 4548 3307
rect 4482 3257 4498 3291
rect 4532 3257 4548 3291
rect 4482 3241 4548 3257
rect 4600 3291 4666 3307
rect 4600 3257 4616 3291
rect 4650 3257 4666 3291
rect 4600 3241 4666 3257
rect 4718 3291 4784 3307
rect 4718 3257 4734 3291
rect 4768 3257 4784 3291
rect 4718 3241 4784 3257
rect 4836 3291 4902 3307
rect 4836 3257 4852 3291
rect 4886 3257 4902 3291
rect 4836 3241 4902 3257
rect 4954 3291 5020 3307
rect 4954 3257 4970 3291
rect 5004 3257 5020 3291
rect 4954 3241 5020 3257
rect 2243 3102 2303 3133
rect 2361 3102 2421 3133
rect 2479 3102 2539 3133
rect 2597 3102 2657 3133
rect 2715 3102 2775 3133
rect 2833 3102 2893 3133
rect 2951 3102 3011 3133
rect 3069 3102 3129 3133
rect 3187 3102 3247 3133
rect 3305 3102 3365 3133
rect 3423 3102 3483 3133
rect 3541 3102 3601 3133
rect 3659 3102 3719 3133
rect 3777 3102 3837 3133
rect 3895 3102 3955 3133
rect 4013 3102 4073 3133
rect 4131 3102 4191 3133
rect 4249 3102 4309 3133
rect 4367 3102 4427 3133
rect 4485 3102 4545 3133
rect 4603 3102 4663 3133
rect 4721 3102 4781 3133
rect 4839 3102 4899 3133
rect 4957 3102 5017 3133
rect 2243 2871 2303 2902
rect 2361 2871 2421 2902
rect 2479 2871 2539 2902
rect 2597 2871 2657 2902
rect 2715 2871 2775 2902
rect 2833 2871 2893 2902
rect 2951 2871 3011 2902
rect 3069 2871 3129 2902
rect 3187 2871 3247 2902
rect 3305 2871 3365 2902
rect 3423 2871 3483 2902
rect 3541 2871 3601 2902
rect 3659 2871 3719 2902
rect 3777 2871 3837 2902
rect 3895 2871 3955 2902
rect 4013 2871 4073 2902
rect 4131 2871 4191 2902
rect 4249 2871 4309 2902
rect 4367 2871 4427 2902
rect 4485 2871 4545 2902
rect 4603 2871 4663 2902
rect 4721 2871 4781 2902
rect 4839 2871 4899 2902
rect 4957 2871 5017 2902
rect 2240 2855 2306 2871
rect 2240 2821 2256 2855
rect 2290 2821 2306 2855
rect 2240 2805 2306 2821
rect 2358 2855 2424 2871
rect 2358 2821 2374 2855
rect 2408 2821 2424 2855
rect 2358 2805 2424 2821
rect 2476 2855 2542 2871
rect 2476 2821 2492 2855
rect 2526 2821 2542 2855
rect 2476 2805 2542 2821
rect 2594 2855 2660 2871
rect 2594 2821 2610 2855
rect 2644 2821 2660 2855
rect 2594 2805 2660 2821
rect 2712 2855 2778 2871
rect 2712 2821 2728 2855
rect 2762 2821 2778 2855
rect 2712 2805 2778 2821
rect 2830 2855 2896 2871
rect 2830 2821 2846 2855
rect 2880 2821 2896 2855
rect 2830 2805 2896 2821
rect 2948 2855 3014 2871
rect 2948 2821 2964 2855
rect 2998 2821 3014 2855
rect 2948 2805 3014 2821
rect 3066 2855 3132 2871
rect 3066 2821 3082 2855
rect 3116 2821 3132 2855
rect 3066 2805 3132 2821
rect 3184 2855 3250 2871
rect 3184 2821 3200 2855
rect 3234 2821 3250 2855
rect 3184 2805 3250 2821
rect 3302 2855 3368 2871
rect 3302 2821 3318 2855
rect 3352 2821 3368 2855
rect 3302 2805 3368 2821
rect 3420 2855 3486 2871
rect 3420 2821 3436 2855
rect 3470 2821 3486 2855
rect 3420 2805 3486 2821
rect 3538 2855 3604 2871
rect 3538 2821 3554 2855
rect 3588 2821 3604 2855
rect 3538 2805 3604 2821
rect 3656 2855 3722 2871
rect 3656 2821 3672 2855
rect 3706 2821 3722 2855
rect 3656 2805 3722 2821
rect 3774 2855 3840 2871
rect 3774 2821 3790 2855
rect 3824 2821 3840 2855
rect 3774 2805 3840 2821
rect 3892 2855 3958 2871
rect 3892 2821 3908 2855
rect 3942 2821 3958 2855
rect 3892 2805 3958 2821
rect 4010 2855 4076 2871
rect 4010 2821 4026 2855
rect 4060 2821 4076 2855
rect 4010 2805 4076 2821
rect 4128 2855 4194 2871
rect 4128 2821 4144 2855
rect 4178 2821 4194 2855
rect 4128 2805 4194 2821
rect 4246 2855 4312 2871
rect 4246 2821 4262 2855
rect 4296 2821 4312 2855
rect 4246 2805 4312 2821
rect 4364 2855 4430 2871
rect 4364 2821 4380 2855
rect 4414 2821 4430 2855
rect 4364 2805 4430 2821
rect 4482 2855 4548 2871
rect 4482 2821 4498 2855
rect 4532 2821 4548 2855
rect 4482 2805 4548 2821
rect 4600 2855 4666 2871
rect 4600 2821 4616 2855
rect 4650 2821 4666 2855
rect 4600 2805 4666 2821
rect 4718 2855 4784 2871
rect 4718 2821 4734 2855
rect 4768 2821 4784 2855
rect 4718 2805 4784 2821
rect 4836 2855 4902 2871
rect 4836 2821 4852 2855
rect 4886 2821 4902 2855
rect 4836 2805 4902 2821
rect 4954 2855 5020 2871
rect 4954 2821 4970 2855
rect 5004 2821 5020 2855
rect 4954 2805 5020 2821
rect 2243 2666 2303 2697
rect 2361 2666 2421 2697
rect 2479 2666 2539 2697
rect 2597 2666 2657 2697
rect 2715 2666 2775 2697
rect 2833 2666 2893 2697
rect 2951 2666 3011 2697
rect 3069 2666 3129 2697
rect 3187 2666 3247 2697
rect 3305 2666 3365 2697
rect 3423 2666 3483 2697
rect 3541 2666 3601 2697
rect 3659 2666 3719 2697
rect 3777 2666 3837 2697
rect 3895 2666 3955 2697
rect 4013 2666 4073 2697
rect 4131 2666 4191 2697
rect 4249 2666 4309 2697
rect 4367 2666 4427 2697
rect 4485 2666 4545 2697
rect 4603 2666 4663 2697
rect 4721 2666 4781 2697
rect 4839 2666 4899 2697
rect 4957 2666 5017 2697
rect 2243 2435 2303 2466
rect 2361 2435 2421 2466
rect 2479 2435 2539 2466
rect 2597 2435 2657 2466
rect 2715 2435 2775 2466
rect 2833 2435 2893 2466
rect 2951 2435 3011 2466
rect 3069 2435 3129 2466
rect 3187 2435 3247 2466
rect 3305 2435 3365 2466
rect 3423 2435 3483 2466
rect 3541 2435 3601 2466
rect 3659 2435 3719 2466
rect 3777 2435 3837 2466
rect 3895 2435 3955 2466
rect 4013 2435 4073 2466
rect 4131 2435 4191 2466
rect 4249 2435 4309 2466
rect 4367 2435 4427 2466
rect 4485 2435 4545 2466
rect 4603 2435 4663 2466
rect 4721 2435 4781 2466
rect 4839 2435 4899 2466
rect 4957 2435 5017 2466
rect 2240 2419 2306 2435
rect 2240 2385 2256 2419
rect 2290 2385 2306 2419
rect 2240 2369 2306 2385
rect 2358 2419 2424 2435
rect 2358 2385 2374 2419
rect 2408 2385 2424 2419
rect 2358 2369 2424 2385
rect 2476 2419 2542 2435
rect 2476 2385 2492 2419
rect 2526 2385 2542 2419
rect 2476 2369 2542 2385
rect 2594 2419 2660 2435
rect 2594 2385 2610 2419
rect 2644 2385 2660 2419
rect 2594 2369 2660 2385
rect 2712 2419 2778 2435
rect 2712 2385 2728 2419
rect 2762 2385 2778 2419
rect 2712 2369 2778 2385
rect 2830 2419 2896 2435
rect 2830 2385 2846 2419
rect 2880 2385 2896 2419
rect 2830 2369 2896 2385
rect 2948 2419 3014 2435
rect 2948 2385 2964 2419
rect 2998 2385 3014 2419
rect 2948 2369 3014 2385
rect 3066 2419 3132 2435
rect 3066 2385 3082 2419
rect 3116 2385 3132 2419
rect 3066 2369 3132 2385
rect 3184 2419 3250 2435
rect 3184 2385 3200 2419
rect 3234 2385 3250 2419
rect 3184 2369 3250 2385
rect 3302 2419 3368 2435
rect 3302 2385 3318 2419
rect 3352 2385 3368 2419
rect 3302 2369 3368 2385
rect 3420 2419 3486 2435
rect 3420 2385 3436 2419
rect 3470 2385 3486 2419
rect 3420 2369 3486 2385
rect 3538 2419 3604 2435
rect 3538 2385 3554 2419
rect 3588 2385 3604 2419
rect 3538 2369 3604 2385
rect 3656 2419 3722 2435
rect 3656 2385 3672 2419
rect 3706 2385 3722 2419
rect 3656 2369 3722 2385
rect 3774 2419 3840 2435
rect 3774 2385 3790 2419
rect 3824 2385 3840 2419
rect 3774 2369 3840 2385
rect 3892 2419 3958 2435
rect 3892 2385 3908 2419
rect 3942 2385 3958 2419
rect 3892 2369 3958 2385
rect 4010 2419 4076 2435
rect 4010 2385 4026 2419
rect 4060 2385 4076 2419
rect 4010 2369 4076 2385
rect 4128 2419 4194 2435
rect 4128 2385 4144 2419
rect 4178 2385 4194 2419
rect 4128 2369 4194 2385
rect 4246 2419 4312 2435
rect 4246 2385 4262 2419
rect 4296 2385 4312 2419
rect 4246 2369 4312 2385
rect 4364 2419 4430 2435
rect 4364 2385 4380 2419
rect 4414 2385 4430 2419
rect 4364 2369 4430 2385
rect 4482 2419 4548 2435
rect 4482 2385 4498 2419
rect 4532 2385 4548 2419
rect 4482 2369 4548 2385
rect 4600 2419 4666 2435
rect 4600 2385 4616 2419
rect 4650 2385 4666 2419
rect 4600 2369 4666 2385
rect 4718 2419 4784 2435
rect 4718 2385 4734 2419
rect 4768 2385 4784 2419
rect 4718 2369 4784 2385
rect 4836 2419 4902 2435
rect 4836 2385 4852 2419
rect 4886 2385 4902 2419
rect 4836 2369 4902 2385
rect 4954 2419 5020 2435
rect 4954 2385 4970 2419
rect 5004 2385 5020 2419
rect 4954 2369 5020 2385
<< polycont >>
rect 2256 3257 2290 3291
rect 2374 3257 2408 3291
rect 2492 3257 2526 3291
rect 2610 3257 2644 3291
rect 2728 3257 2762 3291
rect 2846 3257 2880 3291
rect 2964 3257 2998 3291
rect 3082 3257 3116 3291
rect 3200 3257 3234 3291
rect 3318 3257 3352 3291
rect 3436 3257 3470 3291
rect 3554 3257 3588 3291
rect 3672 3257 3706 3291
rect 3790 3257 3824 3291
rect 3908 3257 3942 3291
rect 4026 3257 4060 3291
rect 4144 3257 4178 3291
rect 4262 3257 4296 3291
rect 4380 3257 4414 3291
rect 4498 3257 4532 3291
rect 4616 3257 4650 3291
rect 4734 3257 4768 3291
rect 4852 3257 4886 3291
rect 4970 3257 5004 3291
rect 2256 2821 2290 2855
rect 2374 2821 2408 2855
rect 2492 2821 2526 2855
rect 2610 2821 2644 2855
rect 2728 2821 2762 2855
rect 2846 2821 2880 2855
rect 2964 2821 2998 2855
rect 3082 2821 3116 2855
rect 3200 2821 3234 2855
rect 3318 2821 3352 2855
rect 3436 2821 3470 2855
rect 3554 2821 3588 2855
rect 3672 2821 3706 2855
rect 3790 2821 3824 2855
rect 3908 2821 3942 2855
rect 4026 2821 4060 2855
rect 4144 2821 4178 2855
rect 4262 2821 4296 2855
rect 4380 2821 4414 2855
rect 4498 2821 4532 2855
rect 4616 2821 4650 2855
rect 4734 2821 4768 2855
rect 4852 2821 4886 2855
rect 4970 2821 5004 2855
rect 2256 2385 2290 2419
rect 2374 2385 2408 2419
rect 2492 2385 2526 2419
rect 2610 2385 2644 2419
rect 2728 2385 2762 2419
rect 2846 2385 2880 2419
rect 2964 2385 2998 2419
rect 3082 2385 3116 2419
rect 3200 2385 3234 2419
rect 3318 2385 3352 2419
rect 3436 2385 3470 2419
rect 3554 2385 3588 2419
rect 3672 2385 3706 2419
rect 3790 2385 3824 2419
rect 3908 2385 3942 2419
rect 4026 2385 4060 2419
rect 4144 2385 4178 2419
rect 4262 2385 4296 2419
rect 4380 2385 4414 2419
rect 4498 2385 4532 2419
rect 4616 2385 4650 2419
rect 4734 2385 4768 2419
rect 4852 2385 4886 2419
rect 4970 2385 5004 2419
<< locali >>
rect 2083 3687 2179 3721
rect 5081 3687 5177 3721
rect 2083 3625 2117 3687
rect 5143 3625 5177 3687
rect 2197 3526 2231 3542
rect 2197 3334 2231 3350
rect 2315 3526 2349 3542
rect 2315 3334 2349 3350
rect 2433 3526 2467 3542
rect 2433 3334 2467 3350
rect 2551 3526 2585 3542
rect 2551 3334 2585 3350
rect 2669 3526 2703 3542
rect 2669 3334 2703 3350
rect 2787 3526 2821 3542
rect 2787 3334 2821 3350
rect 2905 3526 2939 3542
rect 2905 3334 2939 3350
rect 3023 3526 3057 3542
rect 3023 3334 3057 3350
rect 3141 3526 3175 3542
rect 3141 3334 3175 3350
rect 3259 3526 3293 3542
rect 3259 3334 3293 3350
rect 3377 3526 3411 3542
rect 3377 3334 3411 3350
rect 3495 3526 3529 3542
rect 3495 3334 3529 3350
rect 3613 3526 3647 3542
rect 3613 3334 3647 3350
rect 3731 3526 3765 3542
rect 3731 3334 3765 3350
rect 3849 3526 3883 3542
rect 3849 3334 3883 3350
rect 3967 3526 4001 3542
rect 3967 3334 4001 3350
rect 4085 3526 4119 3542
rect 4085 3334 4119 3350
rect 4203 3526 4237 3542
rect 4203 3334 4237 3350
rect 4321 3526 4355 3542
rect 4321 3334 4355 3350
rect 4439 3526 4473 3542
rect 4439 3334 4473 3350
rect 4557 3526 4591 3542
rect 4557 3334 4591 3350
rect 4675 3526 4709 3542
rect 4675 3334 4709 3350
rect 4793 3526 4827 3542
rect 4793 3334 4827 3350
rect 4911 3526 4945 3542
rect 4911 3334 4945 3350
rect 5029 3526 5063 3542
rect 5029 3334 5063 3350
rect 2240 3257 2256 3291
rect 2290 3257 2306 3291
rect 2358 3257 2374 3291
rect 2408 3257 2424 3291
rect 2476 3257 2492 3291
rect 2526 3257 2542 3291
rect 2594 3257 2610 3291
rect 2644 3257 2660 3291
rect 2712 3257 2728 3291
rect 2762 3257 2778 3291
rect 2830 3257 2846 3291
rect 2880 3257 2896 3291
rect 2948 3257 2964 3291
rect 2998 3257 3014 3291
rect 3066 3257 3082 3291
rect 3116 3257 3132 3291
rect 3184 3257 3200 3291
rect 3234 3257 3250 3291
rect 3302 3257 3318 3291
rect 3352 3257 3368 3291
rect 3420 3257 3436 3291
rect 3470 3257 3486 3291
rect 3538 3257 3554 3291
rect 3588 3257 3604 3291
rect 3656 3257 3672 3291
rect 3706 3257 3722 3291
rect 3774 3257 3790 3291
rect 3824 3257 3840 3291
rect 3892 3257 3908 3291
rect 3942 3257 3958 3291
rect 4010 3257 4026 3291
rect 4060 3257 4076 3291
rect 4128 3257 4144 3291
rect 4178 3257 4194 3291
rect 4246 3257 4262 3291
rect 4296 3257 4312 3291
rect 4364 3257 4380 3291
rect 4414 3257 4430 3291
rect 4482 3257 4498 3291
rect 4532 3257 4548 3291
rect 4600 3257 4616 3291
rect 4650 3257 4666 3291
rect 4718 3257 4734 3291
rect 4768 3257 4784 3291
rect 4836 3257 4852 3291
rect 4886 3257 4902 3291
rect 4954 3257 4970 3291
rect 5004 3257 5020 3291
rect 2197 3090 2231 3106
rect 2197 2898 2231 2914
rect 2315 3090 2349 3106
rect 2315 2898 2349 2914
rect 2433 3090 2467 3106
rect 2433 2898 2467 2914
rect 2551 3090 2585 3106
rect 2551 2898 2585 2914
rect 2669 3090 2703 3106
rect 2669 2898 2703 2914
rect 2787 3090 2821 3106
rect 2787 2898 2821 2914
rect 2905 3090 2939 3106
rect 2905 2898 2939 2914
rect 3023 3090 3057 3106
rect 3023 2898 3057 2914
rect 3141 3090 3175 3106
rect 3141 2898 3175 2914
rect 3259 3090 3293 3106
rect 3259 2898 3293 2914
rect 3377 3090 3411 3106
rect 3377 2898 3411 2914
rect 3495 3090 3529 3106
rect 3495 2898 3529 2914
rect 3613 3090 3647 3106
rect 3613 2898 3647 2914
rect 3731 3090 3765 3106
rect 3731 2898 3765 2914
rect 3849 3090 3883 3106
rect 3849 2898 3883 2914
rect 3967 3090 4001 3106
rect 3967 2898 4001 2914
rect 4085 3090 4119 3106
rect 4085 2898 4119 2914
rect 4203 3090 4237 3106
rect 4203 2898 4237 2914
rect 4321 3090 4355 3106
rect 4321 2898 4355 2914
rect 4439 3090 4473 3106
rect 4439 2898 4473 2914
rect 4557 3090 4591 3106
rect 4557 2898 4591 2914
rect 4675 3090 4709 3106
rect 4675 2898 4709 2914
rect 4793 3090 4827 3106
rect 4793 2898 4827 2914
rect 4911 3090 4945 3106
rect 4911 2898 4945 2914
rect 5029 3090 5063 3106
rect 5029 2898 5063 2914
rect 2240 2821 2256 2855
rect 2290 2821 2306 2855
rect 2358 2821 2374 2855
rect 2408 2821 2424 2855
rect 2476 2821 2492 2855
rect 2526 2821 2542 2855
rect 2594 2821 2610 2855
rect 2644 2821 2660 2855
rect 2712 2821 2728 2855
rect 2762 2821 2778 2855
rect 2830 2821 2846 2855
rect 2880 2821 2896 2855
rect 2948 2821 2964 2855
rect 2998 2821 3014 2855
rect 3066 2821 3082 2855
rect 3116 2821 3132 2855
rect 3184 2821 3200 2855
rect 3234 2821 3250 2855
rect 3302 2821 3318 2855
rect 3352 2821 3368 2855
rect 3420 2821 3436 2855
rect 3470 2821 3486 2855
rect 3538 2821 3554 2855
rect 3588 2821 3604 2855
rect 3656 2821 3672 2855
rect 3706 2821 3722 2855
rect 3774 2821 3790 2855
rect 3824 2821 3840 2855
rect 3892 2821 3908 2855
rect 3942 2821 3958 2855
rect 4010 2821 4026 2855
rect 4060 2821 4076 2855
rect 4128 2821 4144 2855
rect 4178 2821 4194 2855
rect 4246 2821 4262 2855
rect 4296 2821 4312 2855
rect 4364 2821 4380 2855
rect 4414 2821 4430 2855
rect 4482 2821 4498 2855
rect 4532 2821 4548 2855
rect 4600 2821 4616 2855
rect 4650 2821 4666 2855
rect 4718 2821 4734 2855
rect 4768 2821 4784 2855
rect 4836 2821 4852 2855
rect 4886 2821 4902 2855
rect 4954 2821 4970 2855
rect 5004 2821 5020 2855
rect 2197 2654 2231 2670
rect 2197 2462 2231 2478
rect 2315 2654 2349 2670
rect 2315 2462 2349 2478
rect 2433 2654 2467 2670
rect 2433 2462 2467 2478
rect 2551 2654 2585 2670
rect 2551 2462 2585 2478
rect 2669 2654 2703 2670
rect 2669 2462 2703 2478
rect 2787 2654 2821 2670
rect 2787 2462 2821 2478
rect 2905 2654 2939 2670
rect 2905 2462 2939 2478
rect 3023 2654 3057 2670
rect 3023 2462 3057 2478
rect 3141 2654 3175 2670
rect 3141 2462 3175 2478
rect 3259 2654 3293 2670
rect 3259 2462 3293 2478
rect 3377 2654 3411 2670
rect 3377 2462 3411 2478
rect 3495 2654 3529 2670
rect 3495 2462 3529 2478
rect 3613 2654 3647 2670
rect 3613 2462 3647 2478
rect 3731 2654 3765 2670
rect 3731 2462 3765 2478
rect 3849 2654 3883 2670
rect 3849 2462 3883 2478
rect 3967 2654 4001 2670
rect 3967 2462 4001 2478
rect 4085 2654 4119 2670
rect 4085 2462 4119 2478
rect 4203 2654 4237 2670
rect 4203 2462 4237 2478
rect 4321 2654 4355 2670
rect 4321 2462 4355 2478
rect 4439 2654 4473 2670
rect 4439 2462 4473 2478
rect 4557 2654 4591 2670
rect 4557 2462 4591 2478
rect 4675 2654 4709 2670
rect 4675 2462 4709 2478
rect 4793 2654 4827 2670
rect 4793 2462 4827 2478
rect 4911 2654 4945 2670
rect 4911 2462 4945 2478
rect 5029 2654 5063 2670
rect 5029 2462 5063 2478
rect 2240 2385 2256 2419
rect 2290 2385 2306 2419
rect 2358 2385 2374 2419
rect 2408 2385 2424 2419
rect 2476 2385 2492 2419
rect 2526 2385 2542 2419
rect 2594 2385 2610 2419
rect 2644 2385 2660 2419
rect 2712 2385 2728 2419
rect 2762 2385 2778 2419
rect 2830 2385 2846 2419
rect 2880 2385 2896 2419
rect 2948 2385 2964 2419
rect 2998 2385 3014 2419
rect 3066 2385 3082 2419
rect 3116 2385 3132 2419
rect 3184 2385 3200 2419
rect 3234 2385 3250 2419
rect 3302 2385 3318 2419
rect 3352 2385 3368 2419
rect 3420 2385 3436 2419
rect 3470 2385 3486 2419
rect 3538 2385 3554 2419
rect 3588 2385 3604 2419
rect 3656 2385 3672 2419
rect 3706 2385 3722 2419
rect 3774 2385 3790 2419
rect 3824 2385 3840 2419
rect 3892 2385 3908 2419
rect 3942 2385 3958 2419
rect 4010 2385 4026 2419
rect 4060 2385 4076 2419
rect 4128 2385 4144 2419
rect 4178 2385 4194 2419
rect 4246 2385 4262 2419
rect 4296 2385 4312 2419
rect 4364 2385 4380 2419
rect 4414 2385 4430 2419
rect 4482 2385 4498 2419
rect 4532 2385 4548 2419
rect 4600 2385 4616 2419
rect 4650 2385 4666 2419
rect 4718 2385 4734 2419
rect 4768 2385 4784 2419
rect 4836 2385 4852 2419
rect 4886 2385 4902 2419
rect 4954 2385 4970 2419
rect 5004 2385 5020 2419
rect 2083 2317 2117 2379
rect 5143 2317 5177 2379
rect 2083 2283 2179 2317
rect 5081 2283 5177 2317
<< viali >>
rect 2197 3350 2231 3526
rect 2315 3350 2349 3526
rect 2433 3350 2467 3526
rect 2551 3350 2585 3526
rect 2669 3350 2703 3526
rect 2787 3350 2821 3526
rect 2905 3350 2939 3526
rect 3023 3350 3057 3526
rect 3141 3350 3175 3526
rect 3259 3350 3293 3526
rect 3377 3350 3411 3526
rect 3495 3350 3529 3526
rect 3613 3350 3647 3526
rect 3731 3350 3765 3526
rect 3849 3350 3883 3526
rect 3967 3350 4001 3526
rect 4085 3350 4119 3526
rect 4203 3350 4237 3526
rect 4321 3350 4355 3526
rect 4439 3350 4473 3526
rect 4557 3350 4591 3526
rect 4675 3350 4709 3526
rect 4793 3350 4827 3526
rect 4911 3350 4945 3526
rect 5029 3350 5063 3526
rect 2256 3257 2290 3291
rect 2374 3257 2408 3291
rect 2492 3257 2526 3291
rect 2610 3257 2644 3291
rect 2728 3257 2762 3291
rect 2846 3257 2880 3291
rect 2964 3257 2998 3291
rect 3082 3257 3116 3291
rect 3200 3257 3234 3291
rect 3318 3257 3352 3291
rect 3436 3257 3470 3291
rect 3554 3257 3588 3291
rect 3672 3257 3706 3291
rect 3790 3257 3824 3291
rect 3908 3257 3942 3291
rect 4026 3257 4060 3291
rect 4144 3257 4178 3291
rect 4262 3257 4296 3291
rect 4380 3257 4414 3291
rect 4498 3257 4532 3291
rect 4616 3257 4650 3291
rect 4734 3257 4768 3291
rect 4852 3257 4886 3291
rect 4970 3257 5004 3291
rect 2197 2914 2231 3090
rect 2315 2914 2349 3090
rect 2433 2914 2467 3090
rect 2551 2914 2585 3090
rect 2669 2914 2703 3090
rect 2787 2914 2821 3090
rect 2905 2914 2939 3090
rect 3023 2914 3057 3090
rect 3141 2914 3175 3090
rect 3259 2914 3293 3090
rect 3377 2914 3411 3090
rect 3495 2914 3529 3090
rect 3613 2914 3647 3090
rect 3731 2914 3765 3090
rect 3849 2914 3883 3090
rect 3967 2914 4001 3090
rect 4085 2914 4119 3090
rect 4203 2914 4237 3090
rect 4321 2914 4355 3090
rect 4439 2914 4473 3090
rect 4557 2914 4591 3090
rect 4675 2914 4709 3090
rect 4793 2914 4827 3090
rect 4911 2914 4945 3090
rect 5029 2914 5063 3090
rect 2256 2821 2290 2855
rect 2374 2821 2408 2855
rect 2492 2821 2526 2855
rect 2610 2821 2644 2855
rect 2728 2821 2762 2855
rect 2846 2821 2880 2855
rect 2964 2821 2998 2855
rect 3082 2821 3116 2855
rect 3200 2821 3234 2855
rect 3318 2821 3352 2855
rect 3436 2821 3470 2855
rect 3554 2821 3588 2855
rect 3672 2821 3706 2855
rect 3790 2821 3824 2855
rect 3908 2821 3942 2855
rect 4026 2821 4060 2855
rect 4144 2821 4178 2855
rect 4262 2821 4296 2855
rect 4380 2821 4414 2855
rect 4498 2821 4532 2855
rect 4616 2821 4650 2855
rect 4734 2821 4768 2855
rect 4852 2821 4886 2855
rect 4970 2821 5004 2855
rect 2197 2478 2231 2654
rect 2315 2478 2349 2654
rect 2433 2478 2467 2654
rect 2551 2478 2585 2654
rect 2669 2478 2703 2654
rect 2787 2478 2821 2654
rect 2905 2478 2939 2654
rect 3023 2478 3057 2654
rect 3141 2478 3175 2654
rect 3259 2478 3293 2654
rect 3377 2478 3411 2654
rect 3495 2478 3529 2654
rect 3613 2478 3647 2654
rect 3731 2478 3765 2654
rect 3849 2478 3883 2654
rect 3967 2478 4001 2654
rect 4085 2478 4119 2654
rect 4203 2478 4237 2654
rect 4321 2478 4355 2654
rect 4439 2478 4473 2654
rect 4557 2478 4591 2654
rect 4675 2478 4709 2654
rect 4793 2478 4827 2654
rect 4911 2478 4945 2654
rect 5029 2478 5063 2654
rect 2256 2385 2290 2419
rect 2374 2385 2408 2419
rect 2492 2385 2526 2419
rect 2610 2385 2644 2419
rect 2728 2385 2762 2419
rect 2846 2385 2880 2419
rect 2964 2385 2998 2419
rect 3082 2385 3116 2419
rect 3200 2385 3234 2419
rect 3318 2385 3352 2419
rect 3436 2385 3470 2419
rect 3554 2385 3588 2419
rect 3672 2385 3706 2419
rect 3790 2385 3824 2419
rect 3908 2385 3942 2419
rect 4026 2385 4060 2419
rect 4144 2385 4178 2419
rect 4262 2385 4296 2419
rect 4380 2385 4414 2419
rect 4498 2385 4532 2419
rect 4616 2385 4650 2419
rect 4734 2385 4768 2419
rect 4852 2385 4886 2419
rect 4970 2385 5004 2419
<< metal1 >>
rect 2191 3526 2237 3538
rect 2191 3350 2197 3526
rect 2231 3350 2237 3526
rect 2191 3338 2237 3350
rect 2309 3526 2355 3538
rect 2309 3350 2315 3526
rect 2349 3350 2355 3526
rect 2309 3338 2355 3350
rect 2427 3526 2473 3538
rect 2427 3350 2433 3526
rect 2467 3350 2473 3526
rect 2427 3338 2473 3350
rect 2545 3526 2591 3538
rect 2545 3350 2551 3526
rect 2585 3350 2591 3526
rect 2545 3338 2591 3350
rect 2663 3526 2709 3538
rect 2663 3350 2669 3526
rect 2703 3350 2709 3526
rect 2663 3338 2709 3350
rect 2781 3526 2827 3538
rect 2781 3350 2787 3526
rect 2821 3350 2827 3526
rect 2781 3338 2827 3350
rect 2899 3526 2945 3538
rect 2899 3350 2905 3526
rect 2939 3350 2945 3526
rect 2899 3338 2945 3350
rect 3017 3526 3063 3538
rect 3017 3350 3023 3526
rect 3057 3350 3063 3526
rect 3017 3338 3063 3350
rect 3135 3526 3181 3538
rect 3135 3350 3141 3526
rect 3175 3350 3181 3526
rect 3135 3338 3181 3350
rect 3253 3526 3299 3538
rect 3253 3350 3259 3526
rect 3293 3350 3299 3526
rect 3253 3338 3299 3350
rect 3371 3526 3417 3538
rect 3371 3350 3377 3526
rect 3411 3350 3417 3526
rect 3371 3338 3417 3350
rect 3489 3526 3535 3538
rect 3489 3350 3495 3526
rect 3529 3350 3535 3526
rect 3489 3338 3535 3350
rect 3607 3526 3653 3538
rect 3607 3350 3613 3526
rect 3647 3350 3653 3526
rect 3607 3338 3653 3350
rect 3725 3526 3771 3538
rect 3725 3350 3731 3526
rect 3765 3350 3771 3526
rect 3725 3338 3771 3350
rect 3843 3526 3889 3538
rect 3843 3350 3849 3526
rect 3883 3350 3889 3526
rect 3843 3338 3889 3350
rect 3961 3526 4007 3538
rect 3961 3350 3967 3526
rect 4001 3350 4007 3526
rect 3961 3338 4007 3350
rect 4079 3526 4125 3538
rect 4079 3350 4085 3526
rect 4119 3350 4125 3526
rect 4079 3338 4125 3350
rect 4197 3526 4243 3538
rect 4197 3350 4203 3526
rect 4237 3350 4243 3526
rect 4197 3338 4243 3350
rect 4315 3526 4361 3538
rect 4315 3350 4321 3526
rect 4355 3350 4361 3526
rect 4315 3338 4361 3350
rect 4433 3526 4479 3538
rect 4433 3350 4439 3526
rect 4473 3350 4479 3526
rect 4433 3338 4479 3350
rect 4551 3526 4597 3538
rect 4551 3350 4557 3526
rect 4591 3350 4597 3526
rect 4551 3338 4597 3350
rect 4669 3526 4715 3538
rect 4669 3350 4675 3526
rect 4709 3350 4715 3526
rect 4669 3338 4715 3350
rect 4787 3526 4833 3538
rect 4787 3350 4793 3526
rect 4827 3350 4833 3526
rect 4787 3338 4833 3350
rect 4905 3526 4951 3538
rect 4905 3350 4911 3526
rect 4945 3350 4951 3526
rect 4905 3338 4951 3350
rect 5023 3526 5069 3538
rect 5023 3350 5029 3526
rect 5063 3350 5069 3526
rect 2191 3307 2240 3338
rect 5023 3307 5069 3350
rect 2191 3291 2306 3307
rect 2191 3257 2256 3291
rect 2290 3257 2306 3291
rect 2191 3241 2306 3257
rect 2358 3291 3132 3307
rect 2358 3257 2374 3291
rect 2408 3257 2492 3291
rect 2526 3257 2610 3291
rect 2644 3257 2728 3291
rect 2762 3257 2846 3291
rect 2880 3257 2964 3291
rect 2998 3257 3082 3291
rect 3116 3257 3132 3291
rect 2358 3241 3132 3257
rect 3188 3291 3246 3297
rect 3188 3257 3200 3291
rect 3234 3257 3246 3291
rect 3188 3251 3246 3257
rect 3306 3291 3364 3297
rect 3306 3257 3318 3291
rect 3352 3257 3364 3291
rect 3306 3251 3364 3257
rect 3424 3291 3482 3297
rect 3424 3257 3436 3291
rect 3470 3257 3482 3291
rect 3424 3251 3482 3257
rect 3542 3291 3600 3297
rect 3542 3257 3554 3291
rect 3588 3257 3600 3291
rect 3542 3251 3600 3257
rect 3660 3291 3718 3297
rect 3660 3257 3672 3291
rect 3706 3257 3718 3291
rect 3660 3251 3718 3257
rect 3778 3291 3836 3297
rect 3778 3257 3790 3291
rect 3824 3257 3836 3291
rect 3778 3251 3836 3257
rect 3896 3291 3954 3297
rect 3896 3257 3908 3291
rect 3942 3257 3954 3291
rect 3896 3251 3954 3257
rect 4014 3291 4072 3297
rect 4014 3257 4026 3291
rect 4060 3257 4072 3291
rect 4014 3251 4072 3257
rect 4128 3291 4902 3307
rect 4128 3257 4144 3291
rect 4178 3257 4262 3291
rect 4296 3257 4380 3291
rect 4414 3257 4498 3291
rect 4532 3257 4616 3291
rect 4650 3257 4734 3291
rect 4768 3257 4852 3291
rect 4886 3257 4902 3291
rect 4128 3241 4902 3257
rect 4954 3291 5069 3307
rect 4954 3257 4970 3291
rect 5004 3257 5069 3291
rect 4954 3241 5069 3257
rect 2191 3090 2237 3102
rect 2191 2914 2197 3090
rect 2231 2914 2237 3090
rect 2191 2902 2237 2914
rect 2309 3090 2355 3102
rect 2309 2914 2315 3090
rect 2349 2914 2355 3090
rect 2309 2902 2355 2914
rect 2427 3090 2473 3102
rect 2427 2914 2433 3090
rect 2467 2914 2473 3090
rect 2427 2902 2473 2914
rect 2545 3090 2591 3102
rect 2545 2914 2551 3090
rect 2585 2914 2591 3090
rect 2545 2902 2591 2914
rect 2663 3090 2709 3102
rect 2663 2914 2669 3090
rect 2703 2914 2709 3090
rect 2663 2902 2709 2914
rect 2781 3090 2827 3102
rect 2781 2914 2787 3090
rect 2821 2914 2827 3090
rect 2781 2902 2827 2914
rect 2899 3090 2945 3102
rect 2899 2914 2905 3090
rect 2939 2914 2945 3090
rect 2899 2902 2945 2914
rect 3017 3090 3063 3102
rect 3017 2914 3023 3090
rect 3057 2914 3063 3090
rect 3017 2902 3063 2914
rect 3135 3090 3181 3102
rect 3135 2914 3141 3090
rect 3175 2914 3181 3090
rect 3135 2902 3181 2914
rect 3253 3090 3299 3102
rect 3253 2914 3259 3090
rect 3293 2914 3299 3090
rect 3253 2902 3299 2914
rect 3371 3090 3417 3102
rect 3371 2914 3377 3090
rect 3411 2914 3417 3090
rect 3371 2902 3417 2914
rect 3489 3090 3535 3102
rect 3489 2914 3495 3090
rect 3529 2914 3535 3090
rect 3489 2902 3535 2914
rect 3607 3090 3653 3102
rect 3607 2914 3613 3090
rect 3647 2914 3653 3090
rect 3607 2902 3653 2914
rect 3725 3090 3771 3102
rect 3725 2914 3731 3090
rect 3765 2914 3771 3090
rect 3725 2902 3771 2914
rect 3843 3090 3889 3102
rect 3843 2914 3849 3090
rect 3883 2914 3889 3090
rect 3843 2902 3889 2914
rect 3961 3090 4007 3102
rect 3961 2914 3967 3090
rect 4001 2914 4007 3090
rect 3961 2902 4007 2914
rect 4079 3090 4125 3102
rect 4079 2914 4085 3090
rect 4119 2914 4125 3090
rect 4079 2902 4125 2914
rect 4197 3090 4243 3102
rect 4197 2914 4203 3090
rect 4237 2914 4243 3090
rect 4197 2902 4243 2914
rect 4315 3090 4361 3102
rect 4315 2914 4321 3090
rect 4355 2914 4361 3090
rect 4315 2902 4361 2914
rect 4433 3090 4479 3102
rect 4433 2914 4439 3090
rect 4473 2914 4479 3090
rect 4433 2902 4479 2914
rect 4551 3090 4597 3102
rect 4551 2914 4557 3090
rect 4591 2914 4597 3090
rect 4551 2902 4597 2914
rect 4669 3090 4715 3102
rect 4669 2914 4675 3090
rect 4709 2914 4715 3090
rect 4669 2902 4715 2914
rect 4787 3090 4833 3102
rect 4787 2914 4793 3090
rect 4827 2914 4833 3090
rect 4787 2902 4833 2914
rect 4905 3090 4951 3102
rect 4905 2914 4911 3090
rect 4945 2914 4951 3090
rect 4905 2902 4951 2914
rect 5023 3090 5069 3102
rect 5023 2914 5029 3090
rect 5063 2914 5069 3090
rect 2191 2871 2240 2902
rect 5023 2871 5069 2914
rect 2191 2855 2542 2871
rect 2191 2821 2256 2855
rect 2290 2821 2374 2855
rect 2408 2821 2492 2855
rect 2526 2821 2542 2855
rect 2191 2805 2542 2821
rect 2594 2855 2778 2871
rect 2594 2821 2610 2855
rect 2644 2821 2728 2855
rect 2762 2821 2778 2855
rect 2594 2805 2778 2821
rect 2830 2855 3250 2871
rect 3305 2870 3368 2871
rect 2830 2821 2846 2855
rect 2880 2821 2964 2855
rect 2998 2821 3082 2855
rect 3116 2821 3200 2855
rect 3234 2821 3250 2855
rect 2830 2805 3250 2821
rect 3294 2860 3486 2870
rect 3294 2805 3305 2860
rect 3365 2855 3486 2860
rect 3365 2821 3436 2855
rect 3470 2821 3486 2855
rect 3295 2740 3305 2805
rect 3365 2805 3486 2821
rect 3531 2860 3611 2870
rect 3365 2740 3375 2805
rect 3295 2730 3375 2740
rect 3531 2740 3541 2860
rect 3601 2740 3611 2860
rect 3656 2855 4076 2871
rect 3656 2821 3672 2855
rect 3706 2821 3790 2855
rect 3824 2821 3908 2855
rect 3942 2821 4026 2855
rect 4060 2821 4076 2855
rect 3656 2805 4076 2821
rect 4129 2855 4549 2871
rect 4129 2821 4144 2855
rect 4178 2821 4262 2855
rect 4296 2821 4380 2855
rect 4414 2821 4498 2855
rect 4532 2821 4549 2855
rect 4129 2805 4549 2821
rect 4600 2855 4784 2871
rect 4600 2821 4616 2855
rect 4650 2821 4734 2855
rect 4768 2821 4784 2855
rect 4600 2805 4784 2821
rect 4836 2855 5069 2871
rect 4836 2821 4852 2855
rect 4886 2821 4970 2855
rect 5004 2821 5069 2855
rect 4836 2805 5069 2821
rect 3531 2730 3611 2740
rect 2191 2654 2237 2666
rect 2191 2478 2197 2654
rect 2231 2478 2237 2654
rect 2191 2466 2237 2478
rect 2309 2654 2355 2666
rect 2309 2478 2315 2654
rect 2349 2478 2355 2654
rect 2309 2466 2355 2478
rect 2427 2654 2473 2666
rect 2427 2478 2433 2654
rect 2467 2478 2473 2654
rect 2427 2466 2473 2478
rect 2545 2654 2591 2666
rect 2545 2478 2551 2654
rect 2585 2478 2591 2654
rect 2545 2466 2591 2478
rect 2663 2654 2709 2666
rect 2663 2478 2669 2654
rect 2703 2478 2709 2654
rect 2663 2466 2709 2478
rect 2781 2654 2827 2666
rect 2781 2478 2787 2654
rect 2821 2478 2827 2654
rect 2781 2466 2827 2478
rect 2899 2654 2945 2666
rect 2899 2478 2905 2654
rect 2939 2478 2945 2654
rect 2899 2466 2945 2478
rect 3017 2654 3063 2666
rect 3017 2478 3023 2654
rect 3057 2478 3063 2654
rect 3017 2466 3063 2478
rect 3135 2654 3181 2666
rect 3135 2478 3141 2654
rect 3175 2478 3181 2654
rect 3135 2466 3181 2478
rect 3253 2654 3299 2666
rect 3253 2478 3259 2654
rect 3293 2478 3299 2654
rect 3253 2466 3299 2478
rect 3371 2654 3417 2666
rect 3371 2478 3377 2654
rect 3411 2478 3417 2654
rect 3371 2466 3417 2478
rect 3489 2654 3535 2666
rect 3489 2478 3495 2654
rect 3529 2478 3535 2654
rect 3489 2466 3535 2478
rect 3607 2654 3653 2666
rect 3607 2478 3613 2654
rect 3647 2478 3653 2654
rect 3607 2466 3653 2478
rect 3725 2654 3771 2666
rect 3725 2478 3731 2654
rect 3765 2478 3771 2654
rect 3725 2466 3771 2478
rect 3843 2654 3889 2666
rect 3843 2478 3849 2654
rect 3883 2478 3889 2654
rect 3843 2466 3889 2478
rect 3961 2654 4007 2666
rect 3961 2478 3967 2654
rect 4001 2478 4007 2654
rect 3961 2466 4007 2478
rect 4079 2654 4125 2666
rect 4079 2478 4085 2654
rect 4119 2478 4125 2654
rect 4079 2466 4125 2478
rect 4197 2654 4243 2666
rect 4197 2478 4203 2654
rect 4237 2478 4243 2654
rect 4197 2466 4243 2478
rect 4315 2654 4361 2666
rect 4315 2478 4321 2654
rect 4355 2478 4361 2654
rect 4315 2466 4361 2478
rect 4433 2654 4479 2666
rect 4433 2478 4439 2654
rect 4473 2478 4479 2654
rect 4433 2466 4479 2478
rect 4551 2654 4597 2666
rect 4551 2478 4557 2654
rect 4591 2478 4597 2654
rect 4551 2466 4597 2478
rect 4669 2654 4715 2666
rect 4669 2478 4675 2654
rect 4709 2478 4715 2654
rect 4669 2466 4715 2478
rect 4787 2654 4833 2666
rect 4787 2478 4793 2654
rect 4827 2478 4833 2654
rect 4787 2466 4833 2478
rect 4905 2654 4951 2666
rect 4905 2478 4911 2654
rect 4945 2478 4951 2654
rect 4905 2466 4951 2478
rect 5023 2654 5069 2666
rect 5023 2478 5029 2654
rect 5063 2478 5069 2654
rect 2190 2435 2240 2466
rect 5023 2435 5069 2478
rect 2190 2419 2306 2435
rect 2190 2385 2256 2419
rect 2290 2385 2306 2419
rect 2190 2369 2306 2385
rect 2358 2419 3132 2435
rect 2358 2385 2374 2419
rect 2408 2385 2492 2419
rect 2526 2385 2610 2419
rect 2644 2385 2728 2419
rect 2762 2385 2846 2419
rect 2880 2385 2964 2419
rect 2998 2385 3082 2419
rect 3116 2385 3132 2419
rect 2358 2369 3132 2385
rect 3188 2419 3246 2425
rect 3188 2385 3200 2419
rect 3234 2385 3246 2419
rect 3188 2379 3246 2385
rect 3302 2419 4076 2435
rect 3302 2385 3318 2419
rect 3352 2385 3436 2419
rect 3470 2385 3554 2419
rect 3588 2385 3672 2419
rect 3706 2385 3790 2419
rect 3824 2385 3908 2419
rect 3942 2385 4026 2419
rect 4060 2385 4076 2419
rect 3302 2369 4076 2385
rect 4128 2419 4902 2435
rect 4128 2385 4144 2419
rect 4178 2385 4262 2419
rect 4296 2385 4380 2419
rect 4414 2385 4498 2419
rect 4532 2385 4616 2419
rect 4650 2385 4734 2419
rect 4768 2385 4852 2419
rect 4886 2385 4902 2419
rect 4128 2369 4902 2385
rect 4954 2419 5069 2435
rect 4954 2385 4970 2419
rect 5004 2385 5069 2419
rect 4954 2369 5069 2385
<< via1 >>
rect 3305 2855 3365 2860
rect 3305 2821 3318 2855
rect 3318 2821 3352 2855
rect 3352 2821 3365 2855
rect 3305 2740 3365 2821
rect 3541 2855 3601 2860
rect 3541 2821 3554 2855
rect 3554 2821 3588 2855
rect 3588 2821 3601 2855
rect 3541 2740 3601 2821
<< metal2 >>
rect 3302 2870 3368 2871
rect 3295 2860 3375 2870
rect 3295 2740 3305 2860
rect 3365 2740 3375 2860
rect 3295 2730 3375 2740
rect 3531 2860 3611 2870
rect 3531 2740 3541 2860
rect 3601 2740 3611 2860
rect 3531 2730 3611 2740
<< via2 >>
rect 3305 2740 3365 2860
rect 3541 2740 3601 2860
<< metal3 >>
rect 3295 2860 3375 2870
rect 3295 2740 3305 2860
rect 3365 2740 3375 2860
rect 3295 2730 3375 2740
rect 3531 2860 3611 2870
rect 3531 2740 3541 2860
rect 3601 2740 3611 2860
rect 3531 2730 3611 2740
<< end >>
